VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO decred_hash_macro
  CLASS BLOCK ;
  FOREIGN decred_hash_macro ;
  ORIGIN 0.000 0.000 ;
  SIZE 1200.000 BY 1000.000 ;
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 655.130 996.000 655.410 1000.000 ;
    END
  END CLK
  PIN DATA_AVAILABLE
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 724.130 0.000 724.410 4.000 ;
    END
  END DATA_AVAILABLE
  PIN DATA_FROM_HASH[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.450 0.000 122.730 4.000 ;
    END
  END DATA_FROM_HASH[0]
  PIN DATA_FROM_HASH[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.850 0.000 3.130 4.000 ;
    END
  END DATA_FROM_HASH[1]
  PIN DATA_FROM_HASH[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 896.170 996.000 896.450 1000.000 ;
    END
  END DATA_FROM_HASH[2]
  PIN DATA_FROM_HASH[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1084.770 0.000 1085.050 4.000 ;
    END
  END DATA_FROM_HASH[3]
  PIN DATA_FROM_HASH[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 194.520 1200.000 195.120 ;
    END
  END DATA_FROM_HASH[4]
  PIN DATA_FROM_HASH[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.490 0.000 363.770 4.000 ;
    END
  END DATA_FROM_HASH[5]
  PIN DATA_FROM_HASH[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.970 996.000 174.250 1000.000 ;
    END
  END DATA_FROM_HASH[6]
  PIN DATA_FROM_HASH[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 715.400 4.000 716.000 ;
    END
  END DATA_FROM_HASH[7]
  PIN DATA_TO_HASH[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 414.090 996.000 414.370 1000.000 ;
    END
  END DATA_TO_HASH[0]
  PIN DATA_TO_HASH[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 359.080 4.000 359.680 ;
    END
  END DATA_TO_HASH[1]
  PIN DATA_TO_HASH[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 372.680 1200.000 373.280 ;
    END
  END DATA_TO_HASH[2]
  PIN DATA_TO_HASH[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 16.360 1200.000 16.960 ;
    END
  END DATA_TO_HASH[3]
  PIN DATA_TO_HASH[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 892.200 4.000 892.800 ;
    END
  END DATA_TO_HASH[4]
  PIN DATA_TO_HASH[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.970 0.000 243.250 4.000 ;
    END
  END DATA_TO_HASH[5]
  PIN DATA_TO_HASH[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1015.770 996.000 1016.050 1000.000 ;
    END
  END DATA_TO_HASH[6]
  PIN DATA_TO_HASH[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.490 996.000 294.770 1000.000 ;
    END
  END DATA_TO_HASH[7]
  PIN HASH_ADDR[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 775.650 996.000 775.930 1000.000 ;
    END
  END HASH_ADDR[0]
  PIN HASH_ADDR[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.450 996.000 53.730 1000.000 ;
    END
  END HASH_ADDR[1]
  PIN HASH_ADDR[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1136.290 996.000 1136.570 1000.000 ;
    END
  END HASH_ADDR[2]
  PIN HASH_ADDR[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 965.170 0.000 965.450 4.000 ;
    END
  END HASH_ADDR[3]
  PIN HASH_ADDR[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 180.920 4.000 181.520 ;
    END
  END HASH_ADDR[4]
  PIN HASH_ADDR[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 905.800 1200.000 906.400 ;
    END
  END HASH_ADDR[5]
  PIN HASH_EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 484.010 0.000 484.290 4.000 ;
    END
  END HASH_EN
  PIN MACRO_RD_SELECT
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 603.610 0.000 603.890 4.000 ;
    END
  END MACRO_RD_SELECT
  PIN MACRO_WR_SELECT
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 550.840 1200.000 551.440 ;
    END
  END MACRO_WR_SELECT
  PIN THREAD_COUNT[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 727.640 1200.000 728.240 ;
    END
  END THREAD_COUNT[0]
  PIN THREAD_COUNT[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 537.240 4.000 537.840 ;
    END
  END THREAD_COUNT[1]
  PIN THREAD_COUNT[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 534.610 996.000 534.890 1000.000 ;
    END
  END THREAD_COUNT[2]
  PIN THREAD_COUNT[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 844.650 0.000 844.930 4.000 ;
    END
  END THREAD_COUNT[3]
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1096.240 10.640 1097.840 987.600 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 987.600 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 987.600 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 987.600 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 987.600 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 987.600 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 987.600 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 987.600 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1173.040 10.640 1174.640 987.600 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1019.440 10.640 1021.040 987.600 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 987.600 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 987.600 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 987.600 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 987.600 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 987.600 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 987.600 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 0.425 1194.160 987.445 ;
      LAYER met1 ;
        RECT 2.830 0.040 1194.160 987.600 ;
      LAYER met2 ;
        RECT 0.090 995.720 53.170 996.000 ;
        RECT 54.010 995.720 173.690 996.000 ;
        RECT 174.530 995.720 294.210 996.000 ;
        RECT 295.050 995.720 413.810 996.000 ;
        RECT 414.650 995.720 534.330 996.000 ;
        RECT 535.170 995.720 654.850 996.000 ;
        RECT 655.690 995.720 775.370 996.000 ;
        RECT 776.210 995.720 895.890 996.000 ;
        RECT 896.730 995.720 1015.490 996.000 ;
        RECT 1016.330 995.720 1136.010 996.000 ;
        RECT 1136.850 995.720 1192.220 996.000 ;
        RECT 0.090 4.280 1192.220 995.720 ;
        RECT 0.090 0.010 2.570 4.280 ;
        RECT 3.410 0.010 122.170 4.280 ;
        RECT 123.010 0.010 242.690 4.280 ;
        RECT 243.530 0.010 363.210 4.280 ;
        RECT 364.050 0.010 483.730 4.280 ;
        RECT 484.570 0.010 603.330 4.280 ;
        RECT 604.170 0.010 723.850 4.280 ;
        RECT 724.690 0.010 844.370 4.280 ;
        RECT 845.210 0.010 964.890 4.280 ;
        RECT 965.730 0.010 1084.490 4.280 ;
        RECT 1085.330 0.010 1192.220 4.280 ;
      LAYER met3 ;
        RECT 0.065 906.800 1196.000 987.525 ;
        RECT 0.065 905.400 1195.600 906.800 ;
        RECT 0.065 893.200 1196.000 905.400 ;
        RECT 4.400 891.800 1196.000 893.200 ;
        RECT 0.065 728.640 1196.000 891.800 ;
        RECT 0.065 727.240 1195.600 728.640 ;
        RECT 0.065 716.400 1196.000 727.240 ;
        RECT 4.400 715.000 1196.000 716.400 ;
        RECT 0.065 551.840 1196.000 715.000 ;
        RECT 0.065 550.440 1195.600 551.840 ;
        RECT 0.065 538.240 1196.000 550.440 ;
        RECT 4.400 536.840 1196.000 538.240 ;
        RECT 0.065 373.680 1196.000 536.840 ;
        RECT 0.065 372.280 1195.600 373.680 ;
        RECT 0.065 360.080 1196.000 372.280 ;
        RECT 4.400 358.680 1196.000 360.080 ;
        RECT 0.065 195.520 1196.000 358.680 ;
        RECT 0.065 194.120 1195.600 195.520 ;
        RECT 0.065 181.920 1196.000 194.120 ;
        RECT 4.400 180.520 1196.000 181.920 ;
        RECT 0.065 17.360 1196.000 180.520 ;
        RECT 0.065 15.960 1195.600 17.360 ;
        RECT 0.065 0.175 1196.000 15.960 ;
      LAYER met4 ;
        RECT 14.095 10.240 20.640 985.825 ;
        RECT 23.040 10.240 97.440 985.825 ;
        RECT 99.840 10.240 174.240 985.825 ;
        RECT 176.640 10.240 251.040 985.825 ;
        RECT 253.440 10.240 327.840 985.825 ;
        RECT 330.240 10.240 404.640 985.825 ;
        RECT 407.040 10.240 481.440 985.825 ;
        RECT 483.840 10.240 558.240 985.825 ;
        RECT 560.640 10.240 635.040 985.825 ;
        RECT 637.440 10.240 711.840 985.825 ;
        RECT 714.240 10.240 788.640 985.825 ;
        RECT 791.040 10.240 865.440 985.825 ;
        RECT 867.840 10.240 942.240 985.825 ;
        RECT 944.640 10.240 1019.040 985.825 ;
        RECT 1021.440 10.240 1095.840 985.825 ;
        RECT 1098.240 10.240 1172.640 985.825 ;
        RECT 1175.040 10.240 1178.225 985.825 ;
        RECT 14.095 1.535 1178.225 10.240 ;
      LAYER met5 ;
        RECT 307.860 85.900 947.940 607.700 ;
  END
END decred_hash_macro
END LIBRARY


magic
tech sky130A
magscale 1 2
timestamp 1608864223
<< locali >>
rect 7941 35479 7975 35785
rect 12265 35479 12299 35785
rect 35633 26911 35667 27013
rect 17877 23647 17911 23749
rect 24777 21879 24811 22117
rect 29653 20383 29687 20553
rect 28457 19703 28491 19873
rect 9229 18207 9263 18377
rect 12449 18207 12483 18377
rect 12391 18173 12483 18207
rect 29285 13923 29319 14025
rect 32137 12155 32171 12393
rect 32229 11203 32263 11305
rect 32229 11067 32263 11169
rect 29101 10659 29135 10761
rect 34805 10115 34839 10217
rect 16957 9911 16991 10013
rect 34805 9911 34839 10081
<< viali >>
rect 8309 38505 8343 38539
rect 29837 38505 29871 38539
rect 9045 38369 9079 38403
rect 10701 38369 10735 38403
rect 11345 38369 11379 38403
rect 12633 38369 12667 38403
rect 30021 38369 30055 38403
rect 30205 38369 30239 38403
rect 6929 38301 6963 38335
rect 7205 38301 7239 38335
rect 9137 38165 9171 38199
rect 10793 38165 10827 38199
rect 11437 38165 11471 38199
rect 12725 38165 12759 38199
rect 6193 37961 6227 37995
rect 14013 37961 14047 37995
rect 20821 37961 20855 37995
rect 36461 37961 36495 37995
rect 29837 37893 29871 37927
rect 8125 37825 8159 37859
rect 10057 37825 10091 37859
rect 14565 37825 14599 37859
rect 25605 37825 25639 37859
rect 26341 37825 26375 37859
rect 35173 37825 35207 37859
rect 4629 37757 4663 37791
rect 4905 37757 4939 37791
rect 6837 37757 6871 37791
rect 7849 37757 7883 37791
rect 9505 37757 9539 37791
rect 9965 37757 9999 37791
rect 10609 37757 10643 37791
rect 10977 37757 11011 37791
rect 11437 37757 11471 37791
rect 12449 37757 12483 37791
rect 12725 37757 12759 37791
rect 14841 37757 14875 37791
rect 19257 37757 19291 37791
rect 19533 37757 19567 37791
rect 21465 37757 21499 37791
rect 21741 37757 21775 37791
rect 23949 37757 23983 37791
rect 24225 37757 24259 37791
rect 26065 37757 26099 37791
rect 29837 37757 29871 37791
rect 30481 37757 30515 37791
rect 30757 37757 30791 37791
rect 34897 37757 34931 37791
rect 23121 37689 23155 37723
rect 6929 37621 6963 37655
rect 15945 37621 15979 37655
rect 19073 37621 19107 37655
rect 27445 37621 27479 37655
rect 1685 37417 1719 37451
rect 22293 37417 22327 37451
rect 24409 37417 24443 37451
rect 25329 37417 25363 37451
rect 9045 37349 9079 37383
rect 35265 37349 35299 37383
rect 1777 37281 1811 37315
rect 4997 37281 5031 37315
rect 5089 37281 5123 37315
rect 5917 37281 5951 37315
rect 8217 37281 8251 37315
rect 8309 37281 8343 37315
rect 8677 37281 8711 37315
rect 9689 37281 9723 37315
rect 11069 37281 11103 37315
rect 13369 37281 13403 37315
rect 13737 37281 13771 37315
rect 14105 37281 14139 37315
rect 14381 37281 14415 37315
rect 15301 37281 15335 37315
rect 15945 37281 15979 37315
rect 16037 37281 16071 37315
rect 17233 37281 17267 37315
rect 17509 37281 17543 37315
rect 18889 37281 18923 37315
rect 23305 37281 23339 37315
rect 25513 37281 25547 37315
rect 25789 37281 25823 37315
rect 26525 37281 26559 37315
rect 26801 37281 26835 37315
rect 28641 37281 28675 37315
rect 33517 37281 33551 37315
rect 33885 37281 33919 37315
rect 5641 37213 5675 37247
rect 10793 37213 10827 37247
rect 20913 37213 20947 37247
rect 21189 37213 21223 37247
rect 23029 37213 23063 37247
rect 28917 37213 28951 37247
rect 33609 37213 33643 37247
rect 1961 37145 1995 37179
rect 12357 37145 12391 37179
rect 7205 37077 7239 37111
rect 9781 37077 9815 37111
rect 13185 37077 13219 37111
rect 15393 37077 15427 37111
rect 27905 37077 27939 37111
rect 30021 37077 30055 37111
rect 8677 36873 8711 36907
rect 15853 36873 15887 36907
rect 24593 36805 24627 36839
rect 31493 36805 31527 36839
rect 5549 36737 5583 36771
rect 10977 36737 11011 36771
rect 18061 36737 18095 36771
rect 20177 36737 20211 36771
rect 25973 36737 26007 36771
rect 27077 36737 27111 36771
rect 27353 36737 27387 36771
rect 28733 36737 28767 36771
rect 29561 36737 29595 36771
rect 5365 36669 5399 36703
rect 5733 36669 5767 36703
rect 6101 36669 6135 36703
rect 7205 36669 7239 36703
rect 7941 36669 7975 36703
rect 8861 36669 8895 36703
rect 9321 36669 9355 36703
rect 10057 36669 10091 36703
rect 10149 36669 10183 36703
rect 10793 36669 10827 36703
rect 11713 36669 11747 36703
rect 12725 36669 12759 36703
rect 14013 36669 14047 36703
rect 14197 36669 14231 36703
rect 14289 36669 14323 36703
rect 14473 36669 14507 36703
rect 14841 36669 14875 36703
rect 15393 36669 15427 36703
rect 15669 36669 15703 36703
rect 18337 36669 18371 36703
rect 20453 36669 20487 36703
rect 22477 36669 22511 36703
rect 22845 36669 22879 36703
rect 24777 36669 24811 36703
rect 25329 36669 25363 36703
rect 25881 36669 25915 36703
rect 29285 36669 29319 36703
rect 31401 36669 31435 36703
rect 13461 36601 13495 36635
rect 15577 36601 15611 36635
rect 19717 36601 19751 36635
rect 7389 36533 7423 36567
rect 8033 36533 8067 36567
rect 11805 36533 11839 36567
rect 12909 36533 12943 36567
rect 21557 36533 21591 36567
rect 22385 36533 22419 36567
rect 25237 36533 25271 36567
rect 30665 36533 30699 36567
rect 7481 36329 7515 36363
rect 25513 36329 25547 36363
rect 14197 36261 14231 36295
rect 20361 36261 20395 36295
rect 4813 36193 4847 36227
rect 5365 36193 5399 36227
rect 6745 36193 6779 36227
rect 7389 36193 7423 36227
rect 8125 36193 8159 36227
rect 8861 36193 8895 36227
rect 9965 36193 9999 36227
rect 10333 36193 10367 36227
rect 10701 36193 10735 36227
rect 11621 36193 11655 36227
rect 11805 36193 11839 36227
rect 12357 36193 12391 36227
rect 12541 36193 12575 36227
rect 13737 36193 13771 36227
rect 13921 36193 13955 36227
rect 15301 36193 15335 36227
rect 18705 36193 18739 36227
rect 20913 36193 20947 36227
rect 22661 36193 22695 36227
rect 23121 36193 23155 36227
rect 30021 36193 30055 36227
rect 32137 36193 32171 36227
rect 34253 36193 34287 36227
rect 5457 36125 5491 36159
rect 7481 36125 7515 36159
rect 8217 36125 8251 36159
rect 15393 36125 15427 36159
rect 16405 36125 16439 36159
rect 16681 36125 16715 36159
rect 18981 36125 19015 36159
rect 24133 36125 24167 36159
rect 24409 36125 24443 36159
rect 27353 36125 27387 36159
rect 27629 36125 27663 36159
rect 29745 36125 29779 36159
rect 32413 36125 32447 36159
rect 34529 36125 34563 36159
rect 4905 36057 4939 36091
rect 10609 36057 10643 36091
rect 12725 36057 12759 36091
rect 23029 36057 23063 36091
rect 9045 35989 9079 36023
rect 17969 35989 18003 36023
rect 21005 35989 21039 36023
rect 28733 35989 28767 36023
rect 31125 35989 31159 36023
rect 33517 35989 33551 36023
rect 35633 35989 35667 36023
rect 7941 35785 7975 35819
rect 9413 35785 9447 35819
rect 12265 35785 12299 35819
rect 16681 35785 16715 35819
rect 18337 35785 18371 35819
rect 19073 35785 19107 35819
rect 20821 35785 20855 35819
rect 22661 35785 22695 35819
rect 29745 35785 29779 35819
rect 32413 35785 32447 35819
rect 33241 35785 33275 35819
rect 5825 35717 5859 35751
rect 5181 35649 5215 35683
rect 1777 35581 1811 35615
rect 3801 35581 3835 35615
rect 5365 35581 5399 35615
rect 5917 35581 5951 35615
rect 6837 35581 6871 35615
rect 11069 35717 11103 35751
rect 8033 35649 8067 35683
rect 11253 35649 11287 35683
rect 8309 35581 8343 35615
rect 10609 35581 10643 35615
rect 11161 35581 11195 35615
rect 1961 35445 1995 35479
rect 3985 35445 4019 35479
rect 7021 35445 7055 35479
rect 7941 35445 7975 35479
rect 24409 35717 24443 35751
rect 27169 35717 27203 35751
rect 29285 35717 29319 35751
rect 13277 35649 13311 35683
rect 14289 35649 14323 35683
rect 15577 35649 15611 35683
rect 21281 35649 21315 35683
rect 21557 35649 21591 35683
rect 24593 35649 24627 35683
rect 31125 35649 31159 35683
rect 12449 35581 12483 35615
rect 13001 35581 13035 35615
rect 14381 35581 14415 35615
rect 15301 35581 15335 35615
rect 18061 35581 18095 35615
rect 18153 35581 18187 35615
rect 19257 35581 19291 35615
rect 19993 35581 20027 35615
rect 20177 35581 20211 35615
rect 20545 35581 20579 35615
rect 23949 35581 23983 35615
rect 24501 35581 24535 35615
rect 25513 35581 25547 35615
rect 26157 35581 26191 35615
rect 26341 35581 26375 35615
rect 27353 35581 27387 35615
rect 27537 35581 27571 35615
rect 27721 35581 27755 35615
rect 29561 35581 29595 35615
rect 30849 35581 30883 35615
rect 32965 35581 32999 35615
rect 33057 35581 33091 35615
rect 14841 35513 14875 35547
rect 26433 35513 26467 35547
rect 29469 35513 29503 35547
rect 12265 35445 12299 35479
rect 12541 35445 12575 35479
rect 11805 35241 11839 35275
rect 6377 35173 6411 35207
rect 11161 35173 11195 35207
rect 23857 35173 23891 35207
rect 34437 35173 34471 35207
rect 4077 35105 4111 35139
rect 4997 35105 5031 35139
rect 7297 35105 7331 35139
rect 7481 35105 7515 35139
rect 8033 35105 8067 35139
rect 8217 35105 8251 35139
rect 8953 35105 8987 35139
rect 10425 35105 10459 35139
rect 10885 35105 10919 35139
rect 11621 35105 11655 35139
rect 13093 35105 13127 35139
rect 15577 35105 15611 35139
rect 18061 35105 18095 35139
rect 22385 35105 22419 35139
rect 22569 35105 22603 35139
rect 23121 35105 23155 35139
rect 23213 35105 23247 35139
rect 23397 35105 23431 35139
rect 24317 35105 24351 35139
rect 24777 35105 24811 35139
rect 25513 35105 25547 35139
rect 26341 35105 26375 35139
rect 26801 35105 26835 35139
rect 27077 35105 27111 35139
rect 27261 35105 27295 35139
rect 30757 35105 30791 35139
rect 30849 35105 30883 35139
rect 32781 35105 32815 35139
rect 33057 35105 33091 35139
rect 1409 35037 1443 35071
rect 1685 35037 1719 35071
rect 4721 35037 4755 35071
rect 9045 35037 9079 35071
rect 10241 35037 10275 35071
rect 12817 35037 12851 35071
rect 15301 35037 15335 35071
rect 17785 35037 17819 35071
rect 21557 35037 21591 35071
rect 22109 35037 22143 35071
rect 25053 35037 25087 35071
rect 26617 35037 26651 35071
rect 28641 35037 28675 35071
rect 28917 35037 28951 35071
rect 31309 35037 31343 35071
rect 8401 34969 8435 35003
rect 2789 34901 2823 34935
rect 4169 34901 4203 34935
rect 14197 34901 14231 34935
rect 16865 34901 16899 34935
rect 19165 34901 19199 34935
rect 25605 34901 25639 34935
rect 26157 34901 26191 34935
rect 30021 34901 30055 34935
rect 2145 34697 2179 34731
rect 11437 34697 11471 34731
rect 16221 34697 16255 34731
rect 17233 34697 17267 34731
rect 22109 34697 22143 34731
rect 23305 34697 23339 34731
rect 32965 34697 32999 34731
rect 5825 34629 5859 34663
rect 12449 34629 12483 34663
rect 2881 34561 2915 34595
rect 5181 34561 5215 34595
rect 9045 34561 9079 34595
rect 12817 34561 12851 34595
rect 14841 34561 14875 34595
rect 16957 34561 16991 34595
rect 18889 34561 18923 34595
rect 24501 34561 24535 34595
rect 25605 34561 25639 34595
rect 29561 34561 29595 34595
rect 31677 34561 31711 34595
rect 34897 34561 34931 34595
rect 1777 34493 1811 34527
rect 1961 34493 1995 34527
rect 3157 34493 3191 34527
rect 5365 34493 5399 34527
rect 5917 34493 5951 34527
rect 6929 34493 6963 34527
rect 7389 34493 7423 34527
rect 8217 34493 8251 34527
rect 8953 34493 8987 34527
rect 9965 34493 9999 34527
rect 10241 34493 10275 34527
rect 10701 34493 10735 34527
rect 10793 34493 10827 34527
rect 11345 34493 11379 34527
rect 12909 34493 12943 34527
rect 13369 34493 13403 34527
rect 13829 34493 13863 34527
rect 14381 34493 14415 34527
rect 15117 34493 15151 34527
rect 17049 34493 17083 34527
rect 18981 34493 19015 34527
rect 19901 34493 19935 34527
rect 20177 34493 20211 34527
rect 22293 34493 22327 34527
rect 22753 34493 22787 34527
rect 23489 34493 23523 34527
rect 24225 34493 24259 34527
rect 26801 34493 26835 34527
rect 27077 34493 27111 34527
rect 29285 34493 29319 34527
rect 31401 34493 31435 34527
rect 33701 34493 33735 34527
rect 33793 34493 33827 34527
rect 34253 34493 34287 34527
rect 34989 34493 35023 34527
rect 1869 34425 1903 34459
rect 4537 34425 4571 34459
rect 7665 34425 7699 34459
rect 19441 34425 19475 34459
rect 21557 34425 21591 34459
rect 35449 34425 35483 34459
rect 8309 34357 8343 34391
rect 9781 34357 9815 34391
rect 28365 34357 28399 34391
rect 30665 34357 30699 34391
rect 8309 34153 8343 34187
rect 10057 34153 10091 34187
rect 14197 34153 14231 34187
rect 31493 34153 31527 34187
rect 2053 34085 2087 34119
rect 4077 34085 4111 34119
rect 9965 34085 9999 34119
rect 10149 34085 10183 34119
rect 12633 34085 12667 34119
rect 28917 34085 28951 34119
rect 34989 34085 35023 34119
rect 2605 34017 2639 34051
rect 2697 34017 2731 34051
rect 2881 34017 2915 34051
rect 3157 34017 3191 34051
rect 3341 34017 3375 34051
rect 4905 34017 4939 34051
rect 5825 34017 5859 34051
rect 6469 34017 6503 34051
rect 6561 34017 6595 34051
rect 6745 34017 6779 34051
rect 7021 34017 7055 34051
rect 7205 34017 7239 34051
rect 8217 34017 8251 34051
rect 8493 34017 8527 34051
rect 8861 34017 8895 34051
rect 10517 34017 10551 34051
rect 13369 34017 13403 34051
rect 13921 34017 13955 34051
rect 16865 34017 16899 34051
rect 18981 34017 19015 34051
rect 21925 34017 21959 34051
rect 24225 34017 24259 34051
rect 25237 34017 25271 34051
rect 26801 34017 26835 34051
rect 27261 34017 27295 34051
rect 27721 34017 27755 34051
rect 27905 34017 27939 34051
rect 27997 34017 28031 34051
rect 29101 34017 29135 34051
rect 32229 34017 32263 34051
rect 33333 34017 33367 34051
rect 35449 34017 35483 34051
rect 35541 34017 35575 34051
rect 4629 33949 4663 33983
rect 5089 33949 5123 33983
rect 5917 33949 5951 33983
rect 9781 33949 9815 33983
rect 10977 33949 11011 33983
rect 11253 33949 11287 33983
rect 13829 33949 13863 33983
rect 16589 33949 16623 33983
rect 18705 33949 18739 33983
rect 22017 33949 22051 33983
rect 22293 33949 22327 33983
rect 24133 33949 24167 33983
rect 25145 33949 25179 33983
rect 29377 33949 29411 33983
rect 29929 33949 29963 33983
rect 30205 33949 30239 33983
rect 32137 33949 32171 33983
rect 32689 33949 32723 33983
rect 33609 33949 33643 33983
rect 5641 33881 5675 33915
rect 26617 33881 26651 33915
rect 18153 33813 18187 33847
rect 20269 33813 20303 33847
rect 21741 33813 21775 33847
rect 23581 33813 23615 33847
rect 24409 33813 24443 33847
rect 25421 33813 25455 33847
rect 28181 33813 28215 33847
rect 35725 33813 35759 33847
rect 4905 33609 4939 33643
rect 9229 33609 9263 33643
rect 19993 33609 20027 33643
rect 23857 33609 23891 33643
rect 31585 33609 31619 33643
rect 33701 33609 33735 33643
rect 3801 33473 3835 33507
rect 5549 33473 5583 33507
rect 6929 33473 6963 33507
rect 8769 33473 8803 33507
rect 9965 33473 9999 33507
rect 14841 33473 14875 33507
rect 19717 33473 19751 33507
rect 20729 33473 20763 33507
rect 21741 33473 21775 33507
rect 22293 33473 22327 33507
rect 24593 33473 24627 33507
rect 24869 33473 24903 33507
rect 29285 33473 29319 33507
rect 29561 33473 29595 33507
rect 32321 33473 32355 33507
rect 32597 33473 32631 33507
rect 35173 33473 35207 33507
rect 2789 33405 2823 33439
rect 3341 33405 3375 33439
rect 3709 33405 3743 33439
rect 4261 33405 4295 33439
rect 4721 33405 4755 33439
rect 5733 33405 5767 33439
rect 7113 33405 7147 33439
rect 7481 33405 7515 33439
rect 7849 33405 7883 33439
rect 8125 33405 8159 33439
rect 8953 33405 8987 33439
rect 9045 33405 9079 33439
rect 10517 33405 10551 33439
rect 10609 33405 10643 33439
rect 10793 33405 10827 33439
rect 11069 33405 11103 33439
rect 11253 33405 11287 33439
rect 13645 33405 13679 33439
rect 13921 33405 13955 33439
rect 14105 33405 14139 33439
rect 15117 33405 15151 33439
rect 17049 33405 17083 33439
rect 19441 33405 19475 33439
rect 19809 33405 19843 33439
rect 20821 33405 20855 33439
rect 21833 33405 21867 33439
rect 23673 33405 23707 33439
rect 26709 33405 26743 33439
rect 26985 33405 27019 33439
rect 31401 33405 31435 33439
rect 34897 33405 34931 33439
rect 5917 33337 5951 33371
rect 6285 33337 6319 33371
rect 13093 33337 13127 33371
rect 21281 33337 21315 33371
rect 36553 33337 36587 33371
rect 5825 33269 5859 33303
rect 16221 33269 16255 33303
rect 17141 33269 17175 33303
rect 19257 33269 19291 33303
rect 25973 33269 26007 33303
rect 28089 33269 28123 33303
rect 30849 33269 30883 33303
rect 9321 33065 9355 33099
rect 14749 33065 14783 33099
rect 24777 33065 24811 33099
rect 30481 33065 30515 33099
rect 3065 32997 3099 33031
rect 4445 32997 4479 33031
rect 11161 32997 11195 33031
rect 11521 32997 11555 33031
rect 1409 32929 1443 32963
rect 4353 32929 4387 32963
rect 4721 32929 4755 32963
rect 4997 32929 5031 32963
rect 5365 32929 5399 32963
rect 5733 32929 5767 32963
rect 8585 32929 8619 32963
rect 9505 32929 9539 32963
rect 10517 32929 10551 32963
rect 11345 32929 11379 32963
rect 11437 32929 11471 32963
rect 13921 32929 13955 32963
rect 14473 32929 14507 32963
rect 15669 32929 15703 32963
rect 15761 32929 15795 32963
rect 16129 32929 16163 32963
rect 16865 32929 16899 32963
rect 20913 32929 20947 32963
rect 21189 32929 21223 32963
rect 22569 32929 22603 32963
rect 23489 32929 23523 32963
rect 25421 32929 25455 32963
rect 28825 32929 28859 32963
rect 29377 32929 29411 32963
rect 30297 32929 30331 32963
rect 32137 32929 32171 32963
rect 32873 32929 32907 32963
rect 33701 32929 33735 32963
rect 33885 32929 33919 32963
rect 34989 32929 35023 32963
rect 38853 32929 38887 32963
rect 1685 32861 1719 32895
rect 6469 32861 6503 32895
rect 6745 32861 6779 32895
rect 9689 32861 9723 32895
rect 10241 32861 10275 32895
rect 10701 32861 10735 32895
rect 11897 32861 11931 32895
rect 14565 32861 14599 32895
rect 16589 32861 16623 32895
rect 18705 32861 18739 32895
rect 18981 32861 19015 32895
rect 23213 32861 23247 32895
rect 25329 32861 25363 32895
rect 27169 32861 27203 32895
rect 27445 32861 27479 32895
rect 29285 32861 29319 32895
rect 32965 32861 32999 32895
rect 34713 32861 34747 32895
rect 32413 32793 32447 32827
rect 8033 32725 8067 32759
rect 8769 32725 8803 32759
rect 17969 32725 18003 32759
rect 20085 32725 20119 32759
rect 25605 32725 25639 32759
rect 29561 32725 29595 32759
rect 33977 32725 34011 32759
rect 36277 32725 36311 32759
rect 38945 32725 38979 32759
rect 5549 32521 5583 32555
rect 15761 32521 15795 32555
rect 17693 32521 17727 32555
rect 22845 32521 22879 32555
rect 29561 32521 29595 32555
rect 3249 32453 3283 32487
rect 7205 32453 7239 32487
rect 18981 32453 19015 32487
rect 28089 32453 28123 32487
rect 34069 32453 34103 32487
rect 6285 32385 6319 32419
rect 9965 32385 9999 32419
rect 13185 32385 13219 32419
rect 13461 32385 13495 32419
rect 20453 32385 20487 32419
rect 22569 32385 22603 32419
rect 23673 32385 23707 32419
rect 23949 32385 23983 32419
rect 29285 32385 29319 32419
rect 33333 32385 33367 32419
rect 2145 32317 2179 32351
rect 3341 32317 3375 32351
rect 3893 32317 3927 32351
rect 4169 32317 4203 32351
rect 4445 32317 4479 32351
rect 5089 32317 5123 32351
rect 5733 32317 5767 32351
rect 5825 32317 5859 32351
rect 7113 32317 7147 32351
rect 8309 32317 8343 32351
rect 8585 32317 8619 32351
rect 8769 32317 8803 32351
rect 9873 32317 9907 32351
rect 10333 32317 10367 32351
rect 10609 32317 10643 32351
rect 11069 32317 11103 32351
rect 11253 32317 11287 32351
rect 15669 32317 15703 32351
rect 16037 32317 16071 32351
rect 16405 32317 16439 32351
rect 17141 32317 17175 32351
rect 17877 32317 17911 32351
rect 18061 32317 18095 32351
rect 18521 32317 18555 32351
rect 18889 32317 18923 32351
rect 20729 32317 20763 32351
rect 22109 32317 22143 32351
rect 22661 32317 22695 32351
rect 25789 32317 25823 32351
rect 26065 32317 26099 32351
rect 28273 32317 28307 32351
rect 28733 32317 28767 32351
rect 29377 32317 29411 32351
rect 30573 32317 30607 32351
rect 30849 32317 30883 32351
rect 32965 32317 32999 32351
rect 33609 32317 33643 32351
rect 34161 32317 34195 32351
rect 35449 32317 35483 32351
rect 36277 32317 36311 32351
rect 38669 32317 38703 32351
rect 1961 32249 1995 32283
rect 2329 32249 2363 32283
rect 2697 32249 2731 32283
rect 7757 32249 7791 32283
rect 14841 32249 14875 32283
rect 32229 32249 32263 32283
rect 35265 32249 35299 32283
rect 35817 32249 35851 32283
rect 2237 32181 2271 32215
rect 25053 32181 25087 32215
rect 27169 32181 27203 32215
rect 32781 32181 32815 32215
rect 36369 32181 36403 32215
rect 38761 32181 38795 32215
rect 2329 31977 2363 32011
rect 4261 31977 4295 32011
rect 11253 31977 11287 32011
rect 13093 31977 13127 32011
rect 15393 31977 15427 32011
rect 19625 31977 19659 32011
rect 26893 31977 26927 32011
rect 31125 31977 31159 32011
rect 16865 31909 16899 31943
rect 18521 31909 18555 31943
rect 18705 31909 18739 31943
rect 19073 31909 19107 31943
rect 33793 31909 33827 31943
rect 2513 31841 2547 31875
rect 3065 31841 3099 31875
rect 3249 31841 3283 31875
rect 4077 31841 4111 31875
rect 5549 31841 5583 31875
rect 6653 31841 6687 31875
rect 7113 31841 7147 31875
rect 7849 31841 7883 31875
rect 8217 31841 8251 31875
rect 8585 31841 8619 31875
rect 9045 31841 9079 31875
rect 10149 31841 10183 31875
rect 11989 31841 12023 31875
rect 13001 31841 13035 31875
rect 13737 31841 13771 31875
rect 14013 31841 14047 31875
rect 14565 31841 14599 31875
rect 15485 31841 15519 31875
rect 16037 31841 16071 31875
rect 17693 31841 17727 31875
rect 17877 31841 17911 31875
rect 18613 31841 18647 31875
rect 19533 31841 19567 31875
rect 19993 31841 20027 31875
rect 21005 31841 21039 31875
rect 21557 31841 21591 31875
rect 22661 31841 22695 31875
rect 25145 31841 25179 31875
rect 25697 31841 25731 31875
rect 27077 31841 27111 31875
rect 29377 31841 29411 31875
rect 29929 31841 29963 31875
rect 30297 31841 30331 31875
rect 30941 31841 30975 31875
rect 32137 31841 32171 31875
rect 32413 31841 32447 31875
rect 34529 31841 34563 31875
rect 36645 31841 36679 31875
rect 37749 31841 37783 31875
rect 38761 31841 38795 31875
rect 7665 31773 7699 31807
rect 9873 31773 9907 31807
rect 12081 31773 12115 31807
rect 16129 31773 16163 31807
rect 17417 31773 17451 31807
rect 18337 31773 18371 31807
rect 20913 31773 20947 31807
rect 22385 31773 22419 31807
rect 25513 31773 25547 31807
rect 27261 31773 27295 31807
rect 27537 31773 27571 31807
rect 28917 31773 28951 31807
rect 34805 31773 34839 31807
rect 30297 31705 30331 31739
rect 5641 31637 5675 31671
rect 6469 31637 6503 31671
rect 14657 31637 14691 31671
rect 21189 31637 21223 31671
rect 23949 31637 23983 31671
rect 36093 31637 36127 31671
rect 36737 31637 36771 31671
rect 37933 31637 37967 31671
rect 38945 31637 38979 31671
rect 2973 31433 3007 31467
rect 9505 31433 9539 31467
rect 17417 31433 17451 31467
rect 18337 31433 18371 31467
rect 27353 31433 27387 31467
rect 36737 31433 36771 31467
rect 12449 31365 12483 31399
rect 12541 31365 12575 31399
rect 20545 31365 20579 31399
rect 22477 31365 22511 31399
rect 23949 31365 23983 31399
rect 29377 31365 29411 31399
rect 30757 31365 30791 31399
rect 33149 31365 33183 31399
rect 35725 31365 35759 31399
rect 1409 31297 1443 31331
rect 6193 31297 6227 31331
rect 7573 31297 7607 31331
rect 11437 31297 11471 31331
rect 16037 31297 16071 31331
rect 19809 31297 19843 31331
rect 24317 31297 24351 31331
rect 1685 31229 1719 31263
rect 3709 31229 3743 31263
rect 4261 31229 4295 31263
rect 4537 31229 4571 31263
rect 5457 31229 5491 31263
rect 6101 31229 6135 31263
rect 7297 31229 7331 31263
rect 8953 31229 8987 31263
rect 9413 31229 9447 31263
rect 9965 31229 9999 31263
rect 11713 31229 11747 31263
rect 11897 31229 11931 31263
rect 12909 31229 12943 31263
rect 13645 31229 13679 31263
rect 13921 31229 13955 31263
rect 14381 31229 14415 31263
rect 15117 31229 15151 31263
rect 15209 31229 15243 31263
rect 15577 31229 15611 31263
rect 16221 31229 16255 31263
rect 17233 31229 17267 31263
rect 18153 31229 18187 31263
rect 19165 31229 19199 31263
rect 19717 31229 19751 31263
rect 20453 31229 20487 31263
rect 21189 31229 21223 31263
rect 21649 31229 21683 31263
rect 22385 31229 22419 31263
rect 22661 31229 22695 31263
rect 23857 31229 23891 31263
rect 24133 31229 24167 31263
rect 26249 31229 26283 31263
rect 26433 31229 26467 31263
rect 26801 31229 26835 31263
rect 27261 31229 27295 31263
rect 27997 31229 28031 31263
rect 28641 31229 28675 31263
rect 29469 31229 29503 31263
rect 29837 31229 29871 31263
rect 30481 31229 30515 31263
rect 31125 31229 31159 31263
rect 31493 31229 31527 31263
rect 32413 31229 32447 31263
rect 32781 31229 32815 31263
rect 33149 31229 33183 31263
rect 33977 31229 34011 31263
rect 34897 31229 34931 31263
rect 35265 31229 35299 31263
rect 35817 31229 35851 31263
rect 36645 31229 36679 31263
rect 37473 31229 37507 31263
rect 37749 31229 37783 31263
rect 10885 31161 10919 31195
rect 16405 31161 16439 31195
rect 16773 31161 16807 31195
rect 33793 31161 33827 31195
rect 36461 31161 36495 31195
rect 3617 31093 3651 31127
rect 5549 31093 5583 31127
rect 16313 31093 16347 31127
rect 18981 31093 19015 31127
rect 21741 31093 21775 31127
rect 22845 31093 22879 31127
rect 28457 31093 28491 31127
rect 34069 31093 34103 31127
rect 38853 31093 38887 31127
rect 2513 30889 2547 30923
rect 18613 30889 18647 30923
rect 34253 30889 34287 30923
rect 7205 30821 7239 30855
rect 30021 30821 30055 30855
rect 1777 30753 1811 30787
rect 2697 30753 2731 30787
rect 3249 30753 3283 30787
rect 3433 30753 3467 30787
rect 4077 30753 4111 30787
rect 5365 30753 5399 30787
rect 7665 30753 7699 30787
rect 7849 30753 7883 30787
rect 8033 30753 8067 30787
rect 8677 30753 8711 30787
rect 9689 30753 9723 30787
rect 10425 30753 10459 30787
rect 11989 30753 12023 30787
rect 13369 30753 13403 30787
rect 14105 30753 14139 30787
rect 14565 30753 14599 30787
rect 15301 30753 15335 30787
rect 16221 30753 16255 30787
rect 16957 30753 16991 30787
rect 17417 30753 17451 30787
rect 18521 30753 18555 30787
rect 19165 30753 19199 30787
rect 19441 30753 19475 30787
rect 19901 30753 19935 30787
rect 21557 30753 21591 30787
rect 23673 30753 23707 30787
rect 23949 30753 23983 30787
rect 24225 30753 24259 30787
rect 24593 30753 24627 30787
rect 25329 30753 25363 30787
rect 27169 30753 27203 30787
rect 27721 30753 27755 30787
rect 28825 30753 28859 30787
rect 29469 30753 29503 30787
rect 29837 30753 29871 30787
rect 30573 30753 30607 30787
rect 31217 30753 31251 30787
rect 32689 30753 32723 30787
rect 33057 30753 33091 30787
rect 34161 30753 34195 30787
rect 34897 30753 34931 30787
rect 36645 30753 36679 30787
rect 36921 30753 36955 30787
rect 37749 30753 37783 30787
rect 38117 30753 38151 30787
rect 38485 30753 38519 30787
rect 5089 30685 5123 30719
rect 6745 30685 6779 30719
rect 11713 30685 11747 30719
rect 14197 30685 14231 30719
rect 21281 30685 21315 30719
rect 23857 30685 23891 30719
rect 26893 30685 26927 30719
rect 29009 30685 29043 30719
rect 31309 30685 31343 30719
rect 32229 30685 32263 30719
rect 32965 30685 32999 30719
rect 34989 30685 35023 30719
rect 36093 30685 36127 30719
rect 37105 30685 37139 30719
rect 38853 30685 38887 30719
rect 16313 30617 16347 30651
rect 27629 30617 27663 30651
rect 30757 30617 30791 30651
rect 1869 30549 1903 30583
rect 4261 30549 4295 30583
rect 8861 30549 8895 30583
rect 9873 30549 9907 30583
rect 10609 30549 10643 30583
rect 15485 30549 15519 30583
rect 17601 30549 17635 30583
rect 22661 30549 22695 30583
rect 25421 30549 25455 30583
rect 28641 30549 28675 30583
rect 19625 30345 19659 30379
rect 26525 30345 26559 30379
rect 32229 30345 32263 30379
rect 37473 30345 37507 30379
rect 3709 30277 3743 30311
rect 7665 30277 7699 30311
rect 10333 30277 10367 30311
rect 12541 30277 12575 30311
rect 17417 30277 17451 30311
rect 38117 30277 38151 30311
rect 4813 30209 4847 30243
rect 6285 30209 6319 30243
rect 9689 30209 9723 30243
rect 13737 30209 13771 30243
rect 15577 30209 15611 30243
rect 21741 30209 21775 30243
rect 24961 30209 24995 30243
rect 27077 30209 27111 30243
rect 29469 30209 29503 30243
rect 30849 30209 30883 30243
rect 31125 30209 31159 30243
rect 34253 30209 34287 30243
rect 36185 30209 36219 30243
rect 38853 30209 38887 30243
rect 1685 30141 1719 30175
rect 1777 30141 1811 30175
rect 2421 30141 2455 30175
rect 2789 30141 2823 30175
rect 3157 30141 3191 30175
rect 3525 30141 3559 30175
rect 4537 30141 4571 30175
rect 4721 30141 4755 30175
rect 5825 30141 5859 30175
rect 6009 30141 6043 30175
rect 7021 30141 7055 30175
rect 7205 30141 7239 30175
rect 7757 30141 7791 30175
rect 8401 30141 8435 30175
rect 9321 30141 9355 30175
rect 10057 30141 10091 30175
rect 10333 30141 10367 30175
rect 11345 30141 11379 30175
rect 11529 30141 11563 30175
rect 12541 30141 12575 30175
rect 13001 30141 13035 30175
rect 13921 30141 13955 30175
rect 14289 30141 14323 30175
rect 14473 30141 14507 30175
rect 14933 30141 14967 30175
rect 16129 30141 16163 30175
rect 16405 30141 16439 30175
rect 16589 30141 16623 30175
rect 17325 30141 17359 30175
rect 18061 30141 18095 30175
rect 18337 30141 18371 30175
rect 20177 30141 20211 30175
rect 20637 30141 20671 30175
rect 21005 30141 21039 30175
rect 22201 30141 22235 30175
rect 22385 30141 22419 30175
rect 22569 30141 22603 30175
rect 23949 30141 23983 30175
rect 24133 30141 24167 30175
rect 25237 30141 25271 30175
rect 27353 30141 27387 30175
rect 29837 30141 29871 30175
rect 30205 30141 30239 30175
rect 30389 30141 30423 30175
rect 33241 30141 33275 30175
rect 33977 30141 34011 30175
rect 34897 30141 34931 30175
rect 35081 30141 35115 30175
rect 35909 30141 35943 30175
rect 38117 30141 38151 30175
rect 38761 30141 38795 30175
rect 21281 30073 21315 30107
rect 28733 30073 28767 30107
rect 35449 30073 35483 30107
rect 8585 30005 8619 30039
rect 9137 30005 9171 30039
rect 11161 30005 11195 30039
rect 23765 30005 23799 30039
rect 33333 30005 33367 30039
rect 17141 29801 17175 29835
rect 25237 29801 25271 29835
rect 31033 29801 31067 29835
rect 34989 29801 35023 29835
rect 35909 29801 35943 29835
rect 22017 29733 22051 29767
rect 27997 29733 28031 29767
rect 30573 29733 30607 29767
rect 4077 29665 4111 29699
rect 4629 29665 4663 29699
rect 6009 29665 6043 29699
rect 6561 29665 6595 29699
rect 7205 29665 7239 29699
rect 7573 29665 7607 29699
rect 7757 29665 7791 29699
rect 8401 29665 8435 29699
rect 10057 29665 10091 29699
rect 12633 29665 12667 29699
rect 12725 29665 12759 29699
rect 13369 29665 13403 29699
rect 13829 29665 13863 29699
rect 14289 29665 14323 29699
rect 15301 29665 15335 29699
rect 15945 29665 15979 29699
rect 16129 29665 16163 29699
rect 17049 29665 17083 29699
rect 17785 29665 17819 29699
rect 19073 29665 19107 29699
rect 19441 29665 19475 29699
rect 20177 29665 20211 29699
rect 21281 29665 21315 29699
rect 21741 29665 21775 29699
rect 23305 29665 23339 29699
rect 23581 29665 23615 29699
rect 24041 29665 24075 29699
rect 24225 29665 24259 29699
rect 25237 29665 25271 29699
rect 25421 29665 25455 29699
rect 27261 29665 27295 29699
rect 27813 29665 27847 29699
rect 28457 29665 28491 29699
rect 29469 29665 29503 29699
rect 30021 29665 30055 29699
rect 30297 29665 30331 29699
rect 31217 29665 31251 29699
rect 31309 29665 31343 29699
rect 32505 29665 32539 29699
rect 32689 29665 32723 29699
rect 33885 29665 33919 29699
rect 35817 29665 35851 29699
rect 36737 29665 36771 29699
rect 37013 29665 37047 29699
rect 37933 29665 37967 29699
rect 38117 29665 38151 29699
rect 38301 29665 38335 29699
rect 38945 29665 38979 29699
rect 1409 29597 1443 29631
rect 1685 29597 1719 29631
rect 4905 29597 4939 29631
rect 5825 29597 5859 29631
rect 9781 29597 9815 29631
rect 12541 29597 12575 29631
rect 18061 29597 18095 29631
rect 18797 29597 18831 29631
rect 21097 29597 21131 29631
rect 23489 29597 23523 29631
rect 27077 29597 27111 29631
rect 33057 29597 33091 29631
rect 33609 29597 33643 29631
rect 4353 29529 4387 29563
rect 6469 29529 6503 29563
rect 11345 29529 11379 29563
rect 14473 29529 14507 29563
rect 15393 29529 15427 29563
rect 19441 29529 19475 29563
rect 31493 29529 31527 29563
rect 2973 29461 3007 29495
rect 8585 29461 8619 29495
rect 20269 29461 20303 29495
rect 28641 29461 28675 29495
rect 36553 29461 36587 29495
rect 39037 29461 39071 29495
rect 1869 29257 1903 29291
rect 5733 29257 5767 29291
rect 6193 29257 6227 29291
rect 14657 29257 14691 29291
rect 16773 29257 16807 29291
rect 17417 29257 17451 29291
rect 29745 29257 29779 29291
rect 3157 29189 3191 29223
rect 9873 29189 9907 29223
rect 21741 29189 21775 29223
rect 26433 29189 26467 29223
rect 33241 29189 33275 29223
rect 35725 29189 35759 29223
rect 36645 29189 36679 29223
rect 4905 29121 4939 29155
rect 8309 29121 8343 29155
rect 15393 29121 15427 29155
rect 16129 29121 16163 29155
rect 20085 29121 20119 29155
rect 22293 29121 22327 29155
rect 24133 29121 24167 29155
rect 28089 29121 28123 29155
rect 30297 29121 30331 29155
rect 38025 29121 38059 29155
rect 1777 29053 1811 29087
rect 2421 29053 2455 29087
rect 3065 29053 3099 29087
rect 3249 29053 3283 29087
rect 4169 29053 4203 29087
rect 4537 29053 4571 29087
rect 4813 29053 4847 29087
rect 5917 29053 5951 29087
rect 6009 29053 6043 29087
rect 6843 29053 6877 29087
rect 7573 29053 7607 29087
rect 8861 29053 8895 29087
rect 9137 29053 9171 29087
rect 9321 29053 9355 29087
rect 9965 29053 9999 29087
rect 10517 29053 10551 29087
rect 10609 29053 10643 29087
rect 11345 29053 11379 29087
rect 12449 29053 12483 29087
rect 12725 29053 12759 29087
rect 14565 29053 14599 29087
rect 16589 29053 16623 29087
rect 17325 29053 17359 29087
rect 18061 29053 18095 29087
rect 18889 29053 18923 29087
rect 19073 29053 19107 29087
rect 20453 29053 20487 29087
rect 20729 29053 20763 29087
rect 21557 29053 21591 29087
rect 22109 29053 22143 29087
rect 23673 29053 23707 29087
rect 24225 29053 24259 29087
rect 24501 29053 24535 29087
rect 24869 29053 24903 29087
rect 25605 29053 25639 29087
rect 25973 29053 26007 29087
rect 26433 29053 26467 29087
rect 27261 29053 27295 29087
rect 27537 29053 27571 29087
rect 27997 29053 28031 29087
rect 28917 29053 28951 29087
rect 29561 29053 29595 29087
rect 30573 29053 30607 29087
rect 31953 29053 31987 29087
rect 32413 29053 32447 29087
rect 32781 29053 32815 29087
rect 33241 29053 33275 29087
rect 33977 29053 34011 29087
rect 34897 29053 34931 29087
rect 35265 29053 35299 29087
rect 35725 29053 35759 29087
rect 36461 29053 36495 29087
rect 37473 29053 37507 29087
rect 37933 29053 37967 29087
rect 38117 29053 38151 29087
rect 38669 29053 38703 29087
rect 14105 28985 14139 29019
rect 15669 28985 15703 29019
rect 15761 28985 15795 29019
rect 21005 28985 21039 29019
rect 7021 28917 7055 28951
rect 7757 28917 7791 28951
rect 11529 28917 11563 28951
rect 15577 28917 15611 28951
rect 18337 28917 18371 28951
rect 28733 28917 28767 28951
rect 34161 28917 34195 28951
rect 3341 28713 3375 28747
rect 7665 28713 7699 28747
rect 13461 28713 13495 28747
rect 23489 28713 23523 28747
rect 25881 28713 25915 28747
rect 2145 28645 2179 28679
rect 4261 28645 4295 28679
rect 7113 28645 7147 28679
rect 31033 28645 31067 28679
rect 35265 28645 35299 28679
rect 36829 28645 36863 28679
rect 2237 28577 2271 28611
rect 3157 28577 3191 28611
rect 4169 28577 4203 28611
rect 4353 28577 4387 28611
rect 7849 28577 7883 28611
rect 8585 28577 8619 28611
rect 8953 28577 8987 28611
rect 9781 28577 9815 28611
rect 10609 28577 10643 28611
rect 10793 28577 10827 28611
rect 11529 28577 11563 28611
rect 11989 28577 12023 28611
rect 12357 28577 12391 28611
rect 12725 28577 12759 28611
rect 13553 28577 13587 28611
rect 13921 28577 13955 28611
rect 14197 28577 14231 28611
rect 15301 28577 15335 28611
rect 17601 28577 17635 28611
rect 18521 28577 18555 28611
rect 21373 28577 21407 28611
rect 21925 28577 21959 28611
rect 23305 28577 23339 28611
rect 24041 28577 24075 28611
rect 24409 28577 24443 28611
rect 24777 28577 24811 28611
rect 25697 28577 25731 28611
rect 26801 28577 26835 28611
rect 27261 28577 27295 28611
rect 28089 28577 28123 28611
rect 29929 28577 29963 28611
rect 30389 28577 30423 28611
rect 30757 28577 30791 28611
rect 32321 28577 32355 28611
rect 32965 28577 32999 28611
rect 35725 28577 35759 28611
rect 36369 28577 36403 28611
rect 36553 28577 36587 28611
rect 38301 28577 38335 28611
rect 38485 28577 38519 28611
rect 38669 28577 38703 28611
rect 5457 28509 5491 28543
rect 5733 28509 5767 28543
rect 8217 28509 8251 28543
rect 9137 28509 9171 28543
rect 15577 28509 15611 28543
rect 18245 28509 18279 28543
rect 22201 28509 22235 28543
rect 24685 28509 24719 28543
rect 27813 28509 27847 28543
rect 33609 28509 33643 28543
rect 33885 28509 33919 28543
rect 37841 28509 37875 28543
rect 10885 28441 10919 28475
rect 12725 28441 12759 28475
rect 21649 28441 21683 28475
rect 32413 28441 32447 28475
rect 1961 28373 1995 28407
rect 2421 28373 2455 28407
rect 4537 28373 4571 28407
rect 11345 28373 11379 28407
rect 16681 28373 16715 28407
rect 17693 28373 17727 28407
rect 19809 28373 19843 28407
rect 26617 28373 26651 28407
rect 29377 28373 29411 28407
rect 33057 28373 33091 28407
rect 9965 28169 9999 28203
rect 15485 28169 15519 28203
rect 16129 28169 16163 28203
rect 32781 28169 32815 28203
rect 35081 28169 35115 28203
rect 37381 28169 37415 28203
rect 5457 28101 5491 28135
rect 7021 28101 7055 28135
rect 16681 28101 16715 28135
rect 20729 28101 20763 28135
rect 22293 28101 22327 28135
rect 28089 28101 28123 28135
rect 30573 28101 30607 28135
rect 38761 28101 38795 28135
rect 3249 28033 3283 28067
rect 4629 28033 4663 28067
rect 8033 28033 8067 28067
rect 14289 28033 14323 28067
rect 18521 28033 18555 28067
rect 19349 28033 19383 28067
rect 22845 28033 22879 28067
rect 25881 28033 25915 28067
rect 38117 28033 38151 28067
rect 1961 27965 1995 27999
rect 2605 27965 2639 27999
rect 2973 27965 3007 27999
rect 3341 27965 3375 27999
rect 4077 27965 4111 27999
rect 4537 27965 4571 27999
rect 5365 27965 5399 27999
rect 5825 27965 5859 27999
rect 6009 27965 6043 27999
rect 6837 27965 6871 27999
rect 7757 27965 7791 27999
rect 9873 27965 9907 27999
rect 10241 27965 10275 27999
rect 10885 27965 10919 27999
rect 11529 27965 11563 27999
rect 12449 27965 12483 27999
rect 13645 27965 13679 27999
rect 14013 27965 14047 27999
rect 15393 27965 15427 27999
rect 16313 27965 16347 27999
rect 16405 27965 16439 27999
rect 17049 27965 17083 27999
rect 17233 27965 17267 27999
rect 18153 27965 18187 27999
rect 18889 27965 18923 27999
rect 19625 27965 19659 27999
rect 22017 27965 22051 27999
rect 22569 27965 22603 27999
rect 23765 27965 23799 27999
rect 24317 27965 24351 27999
rect 24593 27965 24627 27999
rect 24869 27965 24903 27999
rect 26157 27965 26191 27999
rect 28273 27965 28307 27999
rect 28549 27965 28583 27999
rect 29653 27965 29687 27999
rect 30205 27965 30239 27999
rect 30573 27965 30607 27999
rect 31217 27965 31251 27999
rect 31953 27965 31987 27999
rect 32229 27965 32263 27999
rect 32965 27965 32999 27999
rect 33241 27965 33275 27999
rect 33609 27965 33643 27999
rect 34161 27965 34195 27999
rect 34989 27965 35023 27999
rect 35817 27965 35851 27999
rect 36093 27965 36127 27999
rect 38485 27965 38519 27999
rect 38761 27965 38795 27999
rect 12541 27897 12575 27931
rect 27537 27897 27571 27931
rect 34345 27897 34379 27931
rect 2053 27829 2087 27863
rect 9321 27829 9355 27863
rect 11621 27829 11655 27863
rect 13553 27829 13587 27863
rect 23949 27829 23983 27863
rect 31309 27829 31343 27863
rect 2973 27625 3007 27659
rect 17601 27625 17635 27659
rect 19073 27625 19107 27659
rect 20085 27625 20119 27659
rect 21097 27625 21131 27659
rect 33885 27625 33919 27659
rect 35633 27625 35667 27659
rect 36553 27625 36587 27659
rect 23857 27557 23891 27591
rect 29377 27557 29411 27591
rect 30941 27557 30975 27591
rect 36737 27557 36771 27591
rect 37105 27557 37139 27591
rect 1409 27489 1443 27523
rect 1685 27489 1719 27523
rect 4353 27489 4387 27523
rect 6193 27489 6227 27523
rect 7021 27489 7055 27523
rect 7665 27489 7699 27523
rect 8677 27489 8711 27523
rect 9137 27489 9171 27523
rect 10149 27489 10183 27523
rect 10425 27489 10459 27523
rect 11069 27489 11103 27523
rect 11345 27489 11379 27523
rect 13369 27489 13403 27523
rect 13921 27489 13955 27523
rect 15577 27489 15611 27523
rect 15669 27489 15703 27523
rect 19073 27489 19107 27523
rect 19257 27489 19291 27523
rect 19993 27489 20027 27523
rect 20913 27489 20947 27523
rect 22109 27489 22143 27523
rect 22293 27489 22327 27523
rect 22477 27489 22511 27523
rect 23121 27489 23155 27523
rect 24409 27489 24443 27523
rect 24777 27489 24811 27523
rect 25145 27489 25179 27523
rect 26617 27489 26651 27523
rect 27077 27489 27111 27523
rect 29837 27489 29871 27523
rect 30297 27489 30331 27523
rect 30757 27489 30791 27523
rect 31401 27489 31435 27523
rect 32321 27489 32355 27523
rect 32505 27489 32539 27523
rect 32965 27489 32999 27523
rect 33793 27489 33827 27523
rect 34345 27489 34379 27523
rect 35357 27489 35391 27523
rect 35541 27489 35575 27523
rect 36645 27489 36679 27523
rect 37749 27489 37783 27523
rect 38301 27489 38335 27523
rect 38945 27489 38979 27523
rect 4077 27421 4111 27455
rect 8769 27421 8803 27455
rect 10241 27421 10275 27455
rect 12725 27421 12759 27455
rect 14013 27421 14047 27455
rect 16221 27421 16255 27455
rect 16497 27421 16531 27455
rect 23489 27421 23523 27455
rect 25605 27421 25639 27455
rect 27721 27421 27755 27455
rect 27997 27421 28031 27455
rect 34621 27421 34655 27455
rect 36369 27421 36403 27455
rect 7849 27353 7883 27387
rect 13461 27353 13495 27387
rect 21925 27353 21959 27387
rect 26617 27353 26651 27387
rect 31493 27353 31527 27387
rect 39037 27353 39071 27387
rect 5641 27285 5675 27319
rect 6377 27285 6411 27319
rect 7113 27285 7147 27319
rect 23259 27285 23293 27319
rect 23397 27285 23431 27319
rect 32229 27285 32263 27319
rect 37841 27285 37875 27319
rect 2329 27081 2363 27115
rect 9689 27081 9723 27115
rect 11345 27081 11379 27115
rect 12541 27081 12575 27115
rect 14841 27081 14875 27115
rect 21097 27081 21131 27115
rect 24501 27081 24535 27115
rect 29377 27081 29411 27115
rect 31033 27081 31067 27115
rect 33149 27081 33183 27115
rect 38853 27081 38887 27115
rect 5641 27013 5675 27047
rect 8493 27013 8527 27047
rect 14105 27013 14139 27047
rect 24133 27013 24167 27047
rect 35081 27013 35115 27047
rect 35633 27013 35667 27047
rect 4445 26945 4479 26979
rect 13369 26945 13403 26979
rect 17049 26945 17083 26979
rect 18981 26945 19015 26979
rect 24225 26945 24259 26979
rect 27721 26945 27755 26979
rect 37749 26945 37783 26979
rect 2421 26877 2455 26911
rect 2881 26877 2915 26911
rect 3065 26877 3099 26911
rect 3893 26877 3927 26911
rect 4077 26877 4111 26911
rect 4905 26877 4939 26911
rect 5549 26877 5583 26911
rect 6285 26877 6319 26911
rect 6837 26877 6871 26911
rect 7389 26877 7423 26911
rect 7665 26877 7699 26911
rect 7849 26877 7883 26911
rect 8677 26877 8711 26911
rect 9137 26877 9171 26911
rect 9873 26877 9907 26911
rect 10241 26877 10275 26911
rect 10517 26877 10551 26911
rect 11253 26877 11287 26911
rect 12449 26877 12483 26911
rect 13553 26877 13587 26911
rect 14013 26877 14047 26911
rect 14749 26877 14783 26911
rect 15393 26877 15427 26911
rect 16129 26877 16163 26911
rect 16497 26877 16531 26911
rect 16957 26877 16991 26911
rect 18889 26877 18923 26911
rect 19073 26877 19107 26911
rect 19533 26877 19567 26911
rect 20085 26877 20119 26911
rect 20453 26877 20487 26911
rect 21005 26877 21039 26911
rect 21741 26877 21775 26911
rect 22109 26877 22143 26911
rect 22293 26877 22327 26911
rect 22661 26877 22695 26911
rect 24004 26877 24038 26911
rect 25605 26877 25639 26911
rect 27537 26877 27571 26911
rect 28089 26877 28123 26911
rect 28549 26877 28583 26911
rect 29561 26877 29595 26911
rect 29837 26877 29871 26911
rect 30849 26877 30883 26911
rect 31585 26877 31619 26911
rect 31861 26877 31895 26911
rect 33701 26877 33735 26911
rect 33885 26877 33919 26911
rect 34897 26877 34931 26911
rect 35633 26877 35667 26911
rect 35725 26877 35759 26911
rect 36277 26877 36311 26911
rect 37473 26877 37507 26911
rect 23857 26809 23891 26843
rect 4997 26741 5031 26775
rect 15577 26741 15611 26775
rect 25697 26741 25731 26775
rect 28641 26741 28675 26775
rect 33977 26741 34011 26775
rect 35817 26741 35851 26775
rect 8309 26537 8343 26571
rect 14565 26537 14599 26571
rect 21097 26537 21131 26571
rect 25605 26537 25639 26571
rect 26617 26537 26651 26571
rect 37933 26537 37967 26571
rect 1961 26469 1995 26503
rect 10425 26469 10459 26503
rect 19809 26469 19843 26503
rect 20361 26469 20395 26503
rect 2421 26401 2455 26435
rect 2789 26401 2823 26435
rect 2881 26401 2915 26435
rect 4077 26401 4111 26435
rect 4813 26401 4847 26435
rect 4905 26401 4939 26435
rect 5733 26401 5767 26435
rect 8217 26401 8251 26435
rect 8585 26401 8619 26435
rect 9689 26401 9723 26435
rect 11253 26401 11287 26435
rect 11437 26401 11471 26435
rect 11897 26401 11931 26435
rect 13001 26401 13035 26435
rect 13553 26401 13587 26435
rect 13645 26401 13679 26435
rect 14381 26401 14415 26435
rect 15761 26401 15795 26435
rect 16129 26401 16163 26435
rect 16221 26401 16255 26435
rect 17049 26401 17083 26435
rect 17417 26401 17451 26435
rect 18245 26401 18279 26435
rect 18337 26401 18371 26435
rect 18705 26401 18739 26435
rect 19901 26401 19935 26435
rect 20913 26401 20947 26435
rect 21833 26401 21867 26435
rect 22569 26401 22603 26435
rect 22845 26401 22879 26435
rect 23305 26401 23339 26435
rect 23673 26401 23707 26435
rect 24225 26401 24259 26435
rect 25421 26401 25455 26435
rect 26525 26401 26559 26435
rect 27077 26401 27111 26435
rect 30113 26401 30147 26435
rect 30665 26401 30699 26435
rect 32321 26401 32355 26435
rect 33517 26401 33551 26435
rect 35541 26401 35575 26435
rect 35817 26401 35851 26435
rect 38025 26401 38059 26435
rect 38393 26401 38427 26435
rect 5457 26333 5491 26367
rect 7113 26333 7147 26367
rect 10977 26333 11011 26367
rect 15301 26333 15335 26367
rect 17141 26333 17175 26367
rect 18061 26333 18095 26367
rect 22109 26333 22143 26367
rect 24593 26333 24627 26367
rect 27813 26333 27847 26367
rect 28089 26333 28123 26367
rect 30757 26333 30791 26367
rect 33241 26333 33275 26367
rect 9781 26265 9815 26299
rect 11989 26265 12023 26299
rect 13093 26265 13127 26299
rect 24501 26265 24535 26299
rect 30021 26265 30055 26299
rect 32505 26265 32539 26299
rect 4261 26197 4295 26231
rect 19625 26197 19659 26231
rect 24363 26197 24397 26231
rect 24869 26197 24903 26231
rect 29193 26197 29227 26231
rect 34621 26197 34655 26231
rect 36921 26197 36955 26231
rect 4169 25993 4203 26027
rect 25605 25993 25639 26027
rect 33241 25993 33275 26027
rect 36277 25993 36311 26027
rect 39037 25993 39071 26027
rect 11805 25925 11839 25959
rect 14657 25925 14691 25959
rect 15577 25925 15611 25959
rect 23949 25925 23983 25959
rect 31861 25925 31895 25959
rect 12449 25857 12483 25891
rect 21373 25857 21407 25891
rect 22109 25857 22143 25891
rect 24685 25857 24719 25891
rect 26433 25857 26467 25891
rect 29653 25857 29687 25891
rect 34897 25857 34931 25891
rect 37473 25857 37507 25891
rect 37749 25857 37783 25891
rect 2605 25789 2639 25823
rect 2881 25789 2915 25823
rect 4721 25789 4755 25823
rect 5733 25789 5767 25823
rect 7113 25789 7147 25823
rect 8125 25789 8159 25823
rect 8677 25789 8711 25823
rect 8861 25789 8895 25823
rect 9413 25789 9447 25823
rect 10701 25789 10735 25823
rect 10885 25789 10919 25823
rect 11253 25789 11287 25823
rect 11621 25789 11655 25823
rect 12725 25789 12759 25823
rect 13829 25789 13863 25823
rect 14289 25789 14323 25823
rect 14565 25789 14599 25823
rect 15301 25789 15335 25823
rect 15853 25789 15887 25823
rect 16129 25789 16163 25823
rect 16957 25789 16991 25823
rect 17141 25789 17175 25823
rect 18613 25789 18647 25823
rect 18705 25789 18739 25823
rect 19165 25789 19199 25823
rect 19809 25789 19843 25823
rect 20453 25789 20487 25823
rect 20637 25789 20671 25823
rect 21189 25789 21223 25823
rect 22385 25789 22419 25823
rect 22937 25789 22971 25823
rect 23673 25789 23707 25823
rect 24593 25789 24627 25823
rect 25421 25789 25455 25823
rect 26709 25789 26743 25823
rect 28549 25789 28583 25823
rect 29377 25789 29411 25823
rect 31677 25789 31711 25823
rect 32229 25789 32263 25823
rect 32505 25789 32539 25823
rect 33149 25789 33183 25823
rect 33885 25789 33919 25823
rect 35173 25789 35207 25823
rect 12633 25721 12667 25755
rect 13185 25721 13219 25755
rect 17509 25721 17543 25755
rect 19533 25721 19567 25755
rect 23121 25721 23155 25755
rect 28089 25721 28123 25755
rect 31033 25721 31067 25755
rect 4905 25653 4939 25687
rect 5917 25653 5951 25687
rect 7297 25653 7331 25687
rect 8125 25653 8159 25687
rect 9505 25653 9539 25687
rect 28641 25653 28675 25687
rect 2973 25449 3007 25483
rect 4169 25449 4203 25483
rect 15393 25449 15427 25483
rect 18705 25449 18739 25483
rect 19533 25449 19567 25483
rect 23489 25449 23523 25483
rect 26617 25449 26651 25483
rect 33517 25449 33551 25483
rect 7757 25381 7791 25415
rect 8125 25381 8159 25415
rect 11529 25381 11563 25415
rect 19257 25381 19291 25415
rect 29285 25381 29319 25415
rect 34529 25381 34563 25415
rect 35081 25381 35115 25415
rect 38209 25381 38243 25415
rect 1409 25313 1443 25347
rect 4353 25313 4387 25347
rect 4537 25313 4571 25347
rect 5641 25313 5675 25347
rect 5825 25313 5859 25347
rect 6101 25313 6135 25347
rect 6837 25313 6871 25347
rect 7573 25313 7607 25347
rect 7665 25313 7699 25347
rect 8585 25313 8619 25347
rect 9873 25313 9907 25347
rect 12817 25313 12851 25347
rect 13277 25313 13311 25347
rect 13553 25313 13587 25347
rect 14565 25313 14599 25347
rect 15393 25313 15427 25347
rect 15853 25313 15887 25347
rect 16129 25313 16163 25347
rect 17141 25313 17175 25347
rect 19441 25313 19475 25347
rect 20913 25313 20947 25347
rect 21649 25313 21683 25347
rect 21741 25313 21775 25347
rect 22293 25313 22327 25347
rect 22569 25313 22603 25347
rect 23305 25313 23339 25347
rect 24777 25313 24811 25347
rect 25145 25313 25179 25347
rect 25789 25313 25823 25347
rect 26617 25313 26651 25347
rect 27077 25313 27111 25347
rect 27353 25313 27387 25347
rect 28641 25313 28675 25347
rect 29929 25313 29963 25347
rect 30297 25313 30331 25347
rect 30941 25313 30975 25347
rect 32321 25313 32355 25347
rect 32505 25313 32539 25347
rect 32689 25313 32723 25347
rect 33333 25313 33367 25347
rect 34713 25313 34747 25347
rect 35541 25313 35575 25347
rect 36001 25313 36035 25347
rect 36553 25313 36587 25347
rect 36737 25313 36771 25347
rect 38301 25313 38335 25347
rect 1685 25245 1719 25279
rect 5549 25245 5583 25279
rect 7389 25245 7423 25279
rect 8677 25245 8711 25279
rect 10149 25245 10183 25279
rect 12633 25245 12667 25279
rect 17417 25245 17451 25279
rect 21005 25245 21039 25279
rect 24961 25245 24995 25279
rect 30021 25245 30055 25279
rect 30389 25245 30423 25279
rect 38761 25245 38795 25279
rect 31125 25177 31159 25211
rect 36921 25177 36955 25211
rect 14657 25109 14691 25143
rect 25881 25109 25915 25143
rect 28733 25109 28767 25143
rect 38025 25109 38059 25143
rect 1685 24905 1719 24939
rect 5641 24905 5675 24939
rect 15209 24905 15243 24939
rect 18521 24905 18555 24939
rect 23029 24905 23063 24939
rect 26525 24905 26559 24939
rect 13829 24837 13863 24871
rect 16129 24837 16163 24871
rect 30021 24837 30055 24871
rect 3065 24769 3099 24803
rect 4077 24769 4111 24803
rect 4353 24769 4387 24803
rect 10425 24769 10459 24803
rect 12541 24769 12575 24803
rect 16773 24769 16807 24803
rect 18061 24769 18095 24803
rect 20453 24769 20487 24803
rect 22293 24769 22327 24803
rect 25421 24769 25455 24803
rect 27997 24769 28031 24803
rect 31769 24769 31803 24803
rect 35449 24769 35483 24803
rect 37289 24769 37323 24803
rect 38669 24769 38703 24803
rect 1593 24701 1627 24735
rect 2237 24701 2271 24735
rect 2973 24701 3007 24735
rect 7113 24701 7147 24735
rect 7481 24701 7515 24735
rect 8033 24701 8067 24735
rect 8309 24701 8343 24735
rect 8493 24701 8527 24735
rect 9505 24701 9539 24735
rect 9781 24701 9815 24735
rect 9965 24701 9999 24735
rect 11069 24701 11103 24735
rect 11253 24701 11287 24735
rect 11437 24701 11471 24735
rect 12449 24701 12483 24735
rect 14013 24701 14047 24735
rect 14197 24701 14231 24735
rect 14381 24701 14415 24735
rect 15025 24701 15059 24735
rect 16313 24701 16347 24735
rect 16681 24701 16715 24735
rect 17325 24701 17359 24735
rect 18337 24701 18371 24735
rect 19809 24701 19843 24735
rect 20545 24701 20579 24735
rect 20821 24701 20855 24735
rect 21189 24701 21223 24735
rect 21465 24701 21499 24735
rect 22201 24701 22235 24735
rect 22845 24701 22879 24735
rect 24041 24701 24075 24735
rect 25145 24701 25179 24735
rect 28273 24701 28307 24735
rect 28457 24701 28491 24735
rect 29561 24701 29595 24735
rect 30113 24701 30147 24735
rect 30297 24701 30331 24735
rect 31309 24701 31343 24735
rect 31677 24701 31711 24735
rect 32321 24701 32355 24735
rect 32597 24701 32631 24735
rect 35541 24701 35575 24735
rect 35909 24701 35943 24735
rect 36093 24701 36127 24735
rect 36553 24701 36587 24735
rect 37565 24701 37599 24735
rect 7205 24633 7239 24667
rect 18245 24633 18279 24667
rect 27445 24633 27479 24667
rect 30849 24633 30883 24667
rect 34897 24633 34931 24667
rect 2329 24565 2363 24599
rect 17417 24565 17451 24599
rect 24225 24565 24259 24599
rect 33701 24565 33735 24599
rect 36737 24565 36771 24599
rect 15945 24361 15979 24395
rect 20269 24361 20303 24395
rect 27169 24361 27203 24395
rect 30389 24361 30423 24395
rect 37841 24361 37875 24395
rect 1869 24293 1903 24327
rect 23029 24293 23063 24327
rect 28641 24293 28675 24327
rect 2421 24225 2455 24259
rect 2697 24225 2731 24259
rect 2881 24225 2915 24259
rect 3341 24225 3375 24259
rect 4353 24225 4387 24259
rect 4813 24225 4847 24259
rect 5917 24225 5951 24259
rect 6285 24225 6319 24259
rect 7021 24225 7055 24259
rect 7573 24225 7607 24259
rect 7757 24225 7791 24259
rect 8585 24225 8619 24259
rect 10149 24225 10183 24259
rect 10333 24225 10367 24259
rect 10517 24225 10551 24259
rect 11161 24225 11195 24259
rect 12725 24225 12759 24259
rect 13093 24225 13127 24259
rect 14289 24225 14323 24259
rect 14565 24225 14599 24259
rect 15301 24225 15335 24259
rect 16137 24225 16171 24259
rect 16313 24225 16347 24259
rect 16957 24225 16991 24259
rect 18245 24225 18279 24259
rect 18429 24225 18463 24259
rect 18613 24225 18647 24259
rect 19257 24225 19291 24259
rect 20085 24225 20119 24259
rect 21373 24225 21407 24259
rect 21649 24225 21683 24259
rect 22293 24225 22327 24259
rect 23673 24225 23707 24259
rect 23765 24225 23799 24259
rect 24041 24225 24075 24259
rect 24133 24225 24167 24259
rect 24869 24225 24903 24259
rect 25605 24225 25639 24259
rect 25789 24225 25823 24259
rect 27353 24225 27387 24259
rect 27629 24225 27663 24259
rect 27905 24225 27939 24259
rect 29285 24225 29319 24259
rect 29653 24225 29687 24259
rect 29837 24225 29871 24259
rect 30481 24225 30515 24259
rect 30757 24225 30791 24259
rect 32505 24225 32539 24259
rect 33057 24225 33091 24259
rect 33333 24225 33367 24259
rect 33609 24225 33643 24259
rect 34069 24225 34103 24259
rect 35081 24225 35115 24259
rect 36921 24225 36955 24259
rect 37841 24225 37875 24259
rect 38301 24225 38335 24259
rect 38577 24225 38611 24259
rect 5457 24157 5491 24191
rect 6193 24157 6227 24191
rect 8125 24157 8159 24191
rect 12265 24157 12299 24191
rect 13737 24157 13771 24191
rect 14749 24157 14783 24191
rect 17049 24157 17083 24191
rect 29377 24157 29411 24191
rect 32597 24157 32631 24191
rect 34805 24157 34839 24191
rect 4169 24089 4203 24123
rect 9965 24089 9999 24123
rect 11345 24089 11379 24123
rect 13001 24089 13035 24123
rect 16497 24089 16531 24123
rect 18061 24089 18095 24123
rect 21189 24089 21223 24123
rect 25145 24089 25179 24123
rect 37013 24089 37047 24123
rect 3433 24021 3467 24055
rect 8769 24021 8803 24055
rect 15393 24021 15427 24055
rect 19441 24021 19475 24055
rect 22477 24021 22511 24055
rect 36369 24021 36403 24055
rect 14013 23817 14047 23851
rect 17141 23817 17175 23851
rect 22937 23817 22971 23851
rect 24133 23817 24167 23851
rect 30113 23817 30147 23851
rect 35909 23817 35943 23851
rect 5641 23749 5675 23783
rect 8493 23749 8527 23783
rect 15577 23749 15611 23783
rect 17877 23749 17911 23783
rect 18337 23749 18371 23783
rect 25973 23749 26007 23783
rect 2789 23681 2823 23715
rect 3433 23681 3467 23715
rect 3709 23681 3743 23715
rect 6929 23681 6963 23715
rect 7481 23681 7515 23715
rect 10885 23681 10919 23715
rect 11897 23681 11931 23715
rect 22293 23681 22327 23715
rect 25329 23681 25363 23715
rect 32045 23681 32079 23715
rect 37013 23681 37047 23715
rect 37289 23681 37323 23715
rect 2053 23613 2087 23647
rect 2421 23613 2455 23647
rect 2697 23613 2731 23647
rect 5733 23613 5767 23647
rect 6285 23613 6319 23647
rect 7757 23613 7791 23647
rect 7941 23613 7975 23647
rect 8401 23613 8435 23647
rect 8861 23613 8895 23647
rect 9597 23613 9631 23647
rect 9873 23613 9907 23647
rect 10333 23613 10367 23647
rect 11437 23613 11471 23647
rect 11713 23613 11747 23647
rect 12449 23613 12483 23647
rect 12725 23613 12759 23647
rect 14565 23613 14599 23647
rect 15301 23613 15335 23647
rect 16037 23613 16071 23647
rect 16129 23613 16163 23647
rect 16957 23613 16991 23647
rect 17877 23613 17911 23647
rect 18061 23613 18095 23647
rect 18613 23613 18647 23647
rect 18889 23613 18923 23647
rect 19901 23613 19935 23647
rect 20453 23613 20487 23647
rect 20637 23613 20671 23647
rect 21189 23613 21223 23647
rect 21557 23613 21591 23647
rect 22017 23613 22051 23647
rect 22753 23613 22787 23647
rect 23857 23613 23891 23647
rect 23949 23613 23983 23647
rect 25697 23613 25731 23647
rect 25973 23613 26007 23647
rect 26709 23613 26743 23647
rect 26985 23613 27019 23647
rect 29285 23613 29319 23647
rect 30021 23613 30055 23647
rect 30665 23613 30699 23647
rect 30941 23613 30975 23647
rect 33333 23613 33367 23647
rect 33793 23613 33827 23647
rect 34161 23613 34195 23647
rect 34897 23613 34931 23647
rect 36093 23613 36127 23647
rect 36369 23613 36403 23647
rect 28365 23545 28399 23579
rect 34253 23545 34287 23579
rect 4997 23477 5031 23511
rect 14749 23477 14783 23511
rect 19717 23477 19751 23511
rect 29469 23477 29503 23511
rect 35081 23477 35115 23511
rect 38393 23477 38427 23511
rect 29469 23273 29503 23307
rect 7021 23205 7055 23239
rect 15301 23205 15335 23239
rect 24961 23205 24995 23239
rect 34345 23205 34379 23239
rect 34897 23205 34931 23239
rect 39037 23205 39071 23239
rect 4905 23137 4939 23171
rect 5365 23137 5399 23171
rect 5825 23137 5859 23171
rect 6101 23137 6135 23171
rect 6285 23137 6319 23171
rect 7573 23137 7607 23171
rect 7849 23137 7883 23171
rect 8033 23137 8067 23171
rect 8493 23137 8527 23171
rect 10333 23137 10367 23171
rect 10885 23137 10919 23171
rect 11253 23137 11287 23171
rect 11713 23137 11747 23171
rect 12173 23137 12207 23171
rect 13001 23137 13035 23171
rect 14473 23137 14507 23171
rect 15761 23137 15795 23171
rect 15945 23137 15979 23171
rect 16129 23137 16163 23171
rect 16957 23137 16991 23171
rect 17141 23137 17175 23171
rect 18429 23137 18463 23171
rect 18705 23137 18739 23171
rect 19901 23137 19935 23171
rect 19993 23137 20027 23171
rect 20269 23137 20303 23171
rect 21005 23137 21039 23171
rect 21833 23137 21867 23171
rect 22937 23137 22971 23171
rect 23121 23137 23155 23171
rect 23489 23137 23523 23171
rect 24225 23137 24259 23171
rect 25789 23137 25823 23171
rect 25973 23137 26007 23171
rect 27353 23137 27387 23171
rect 28365 23137 28399 23171
rect 29193 23137 29227 23171
rect 30113 23137 30147 23171
rect 30849 23137 30883 23171
rect 32321 23137 32355 23171
rect 32505 23137 32539 23171
rect 33057 23137 33091 23171
rect 34253 23137 34287 23171
rect 34437 23137 34471 23171
rect 35357 23137 35391 23171
rect 35541 23137 35575 23171
rect 36461 23137 36495 23171
rect 37197 23137 37231 23171
rect 37749 23137 37783 23171
rect 38209 23137 38243 23171
rect 38945 23137 38979 23171
rect 1409 23069 1443 23103
rect 1685 23069 1719 23103
rect 11069 23069 11103 23103
rect 12725 23069 12759 23103
rect 13185 23069 13219 23103
rect 13645 23069 13679 23103
rect 14197 23069 14231 23103
rect 14657 23069 14691 23103
rect 18061 23069 18095 23103
rect 21925 23069 21959 23103
rect 25513 23069 25547 23103
rect 26525 23069 26559 23103
rect 27077 23069 27111 23103
rect 27537 23069 27571 23103
rect 29101 23069 29135 23103
rect 32965 23069 32999 23103
rect 36829 23069 36863 23103
rect 38485 23069 38519 23103
rect 4721 23001 4755 23035
rect 17325 23001 17359 23035
rect 18705 23001 18739 23035
rect 21833 23001 21867 23035
rect 23397 23001 23431 23035
rect 24409 23001 24443 23035
rect 31033 23001 31067 23035
rect 2973 22933 3007 22967
rect 8677 22933 8711 22967
rect 16773 22933 16807 22967
rect 30297 22933 30331 22967
rect 35633 22933 35667 22967
rect 1777 22729 1811 22763
rect 12541 22729 12575 22763
rect 20729 22729 20763 22763
rect 26525 22729 26559 22763
rect 31401 22729 31435 22763
rect 36461 22729 36495 22763
rect 38853 22729 38887 22763
rect 2513 22661 2547 22695
rect 6193 22661 6227 22695
rect 13185 22661 13219 22695
rect 18889 22661 18923 22695
rect 4261 22593 4295 22627
rect 6837 22593 6871 22627
rect 7573 22593 7607 22627
rect 8493 22593 8527 22627
rect 11713 22593 11747 22627
rect 14105 22593 14139 22627
rect 14841 22593 14875 22627
rect 15761 22593 15795 22627
rect 16497 22593 16531 22627
rect 17233 22593 17267 22627
rect 18245 22593 18279 22627
rect 21373 22593 21407 22627
rect 24225 22593 24259 22627
rect 28365 22593 28399 22627
rect 32965 22593 32999 22627
rect 37473 22593 37507 22627
rect 37749 22593 37783 22627
rect 1685 22525 1719 22559
rect 2329 22525 2363 22559
rect 3341 22525 3375 22559
rect 3525 22525 3559 22559
rect 3801 22525 3835 22559
rect 4721 22525 4755 22559
rect 5365 22525 5399 22559
rect 6009 22525 6043 22559
rect 8217 22525 8251 22559
rect 10977 22525 11011 22559
rect 12449 22525 12483 22559
rect 13185 22525 13219 22559
rect 13737 22525 13771 22559
rect 15025 22525 15059 22559
rect 15485 22525 15519 22559
rect 16773 22525 16807 22559
rect 17141 22525 17175 22559
rect 18429 22525 18463 22559
rect 18889 22525 18923 22559
rect 19809 22525 19843 22559
rect 20545 22525 20579 22559
rect 21281 22525 21315 22559
rect 21649 22525 21683 22559
rect 22293 22525 22327 22559
rect 22937 22525 22971 22559
rect 23765 22525 23799 22559
rect 24133 22525 24167 22559
rect 25145 22525 25179 22559
rect 25421 22525 25455 22559
rect 27905 22525 27939 22559
rect 28457 22525 28491 22559
rect 29469 22525 29503 22559
rect 29929 22525 29963 22559
rect 30297 22525 30331 22559
rect 31217 22525 31251 22559
rect 32505 22525 32539 22559
rect 33241 22525 33275 22559
rect 33333 22525 33367 22559
rect 33977 22525 34011 22559
rect 34897 22525 34931 22559
rect 35173 22525 35207 22559
rect 7113 22457 7147 22491
rect 7205 22457 7239 22491
rect 9873 22457 9907 22491
rect 11345 22457 11379 22491
rect 4813 22389 4847 22423
rect 5457 22389 5491 22423
rect 7021 22389 7055 22423
rect 11161 22389 11195 22423
rect 11253 22389 11287 22423
rect 19993 22389 20027 22423
rect 23029 22389 23063 22423
rect 27905 22389 27939 22423
rect 29745 22389 29779 22423
rect 8677 22185 8711 22219
rect 11437 22185 11471 22219
rect 13185 22185 13219 22219
rect 16865 22185 16899 22219
rect 18429 22185 18463 22219
rect 26709 22185 26743 22219
rect 27721 22185 27755 22219
rect 8769 22117 8803 22151
rect 11529 22117 11563 22151
rect 24777 22117 24811 22151
rect 1501 22049 1535 22083
rect 2145 22049 2179 22083
rect 2973 22049 3007 22083
rect 3525 22049 3559 22083
rect 4077 22049 4111 22083
rect 4629 22049 4663 22083
rect 5365 22049 5399 22083
rect 5825 22049 5859 22083
rect 6469 22049 6503 22083
rect 6929 22049 6963 22083
rect 7481 22049 7515 22083
rect 7757 22049 7791 22083
rect 8401 22049 8435 22083
rect 8585 22049 8619 22083
rect 9137 22049 9171 22083
rect 10517 22049 10551 22083
rect 10701 22049 10735 22083
rect 11345 22049 11379 22083
rect 11897 22049 11931 22083
rect 12357 22049 12391 22083
rect 13185 22049 13219 22083
rect 13737 22049 13771 22083
rect 14841 22049 14875 22083
rect 15301 22049 15335 22083
rect 15945 22049 15979 22083
rect 16313 22049 16347 22083
rect 17141 22049 17175 22083
rect 17601 22049 17635 22083
rect 18245 22049 18279 22083
rect 19257 22049 19291 22083
rect 19441 22049 19475 22083
rect 20177 22049 20211 22083
rect 20913 22049 20947 22083
rect 21649 22049 21683 22083
rect 22385 22049 22419 22083
rect 22753 22049 22787 22083
rect 23397 22049 23431 22083
rect 23673 22049 23707 22083
rect 6561 21981 6595 22015
rect 9689 21981 9723 22015
rect 10241 21981 10275 22015
rect 11161 21981 11195 22015
rect 13921 21981 13955 22015
rect 19533 21981 19567 22015
rect 23765 21981 23799 22015
rect 2237 21913 2271 21947
rect 12541 21913 12575 21947
rect 25421 22049 25455 22083
rect 25697 22049 25731 22083
rect 26525 22049 26559 22083
rect 27629 22049 27663 22083
rect 27905 22049 27939 22083
rect 28273 22049 28307 22083
rect 29009 22049 29043 22083
rect 29653 22049 29687 22083
rect 29929 22049 29963 22083
rect 34529 22049 34563 22083
rect 35265 22049 35299 22083
rect 35449 22049 35483 22083
rect 35817 22049 35851 22083
rect 36185 22049 36219 22083
rect 36921 22049 36955 22083
rect 37841 22049 37875 22083
rect 38301 22049 38335 22083
rect 25053 21981 25087 22015
rect 25973 21981 26007 22015
rect 31033 21981 31067 22015
rect 32137 21981 32171 22015
rect 32413 21981 32447 22015
rect 35173 21981 35207 22015
rect 38577 21981 38611 22015
rect 37841 21913 37875 21947
rect 1593 21845 1627 21879
rect 2881 21845 2915 21879
rect 4169 21845 4203 21879
rect 5365 21845 5399 21879
rect 14657 21845 14691 21879
rect 15393 21845 15427 21879
rect 20269 21845 20303 21879
rect 21097 21845 21131 21879
rect 21833 21845 21867 21879
rect 24777 21845 24811 21879
rect 29101 21845 29135 21879
rect 33701 21845 33735 21879
rect 37105 21845 37139 21879
rect 3709 21641 3743 21675
rect 8033 21641 8067 21675
rect 11529 21641 11563 21675
rect 18245 21641 18279 21675
rect 20177 21641 20211 21675
rect 25053 21641 25087 21675
rect 34161 21641 34195 21675
rect 38853 21641 38887 21675
rect 4813 21573 4847 21607
rect 7297 21573 7331 21607
rect 14289 21573 14323 21607
rect 16589 21573 16623 21607
rect 25881 21573 25915 21607
rect 9229 21505 9263 21539
rect 13185 21505 13219 21539
rect 15945 21505 15979 21539
rect 18889 21505 18923 21539
rect 19625 21505 19659 21539
rect 21925 21505 21959 21539
rect 23673 21505 23707 21539
rect 26617 21505 26651 21539
rect 27721 21505 27755 21539
rect 30297 21505 30331 21539
rect 35449 21505 35483 21539
rect 37565 21505 37599 21539
rect 1685 21437 1719 21471
rect 1777 21437 1811 21471
rect 2605 21437 2639 21471
rect 2973 21437 3007 21471
rect 3157 21437 3191 21471
rect 3617 21437 3651 21471
rect 4997 21437 5031 21471
rect 5273 21437 5307 21471
rect 5457 21437 5491 21471
rect 7113 21437 7147 21471
rect 7849 21437 7883 21471
rect 9137 21437 9171 21471
rect 9597 21437 9631 21471
rect 9873 21437 9907 21471
rect 10333 21437 10367 21471
rect 10517 21437 10551 21471
rect 11253 21437 11287 21471
rect 11345 21437 11379 21471
rect 12449 21437 12483 21471
rect 12633 21437 12667 21471
rect 12725 21437 12759 21471
rect 13829 21437 13863 21471
rect 14381 21437 14415 21471
rect 14933 21437 14967 21471
rect 15117 21437 15151 21471
rect 16313 21437 16347 21471
rect 16681 21437 16715 21471
rect 17325 21437 17359 21471
rect 18061 21437 18095 21471
rect 19073 21437 19107 21471
rect 20085 21437 20119 21471
rect 20821 21437 20855 21471
rect 21465 21437 21499 21471
rect 21649 21437 21683 21471
rect 22017 21437 22051 21471
rect 22937 21437 22971 21471
rect 23949 21437 23983 21471
rect 25881 21437 25915 21471
rect 26525 21437 26559 21471
rect 27997 21437 28031 21471
rect 28549 21437 28583 21471
rect 29285 21437 29319 21471
rect 29653 21437 29687 21471
rect 30113 21437 30147 21471
rect 30573 21437 30607 21471
rect 31217 21437 31251 21471
rect 31861 21437 31895 21471
rect 32045 21437 32079 21471
rect 32781 21437 32815 21471
rect 33241 21437 33275 21471
rect 33977 21437 34011 21471
rect 35725 21437 35759 21471
rect 35909 21437 35943 21471
rect 36369 21437 36403 21471
rect 37289 21437 37323 21471
rect 19257 21369 19291 21403
rect 28733 21369 28767 21403
rect 34897 21369 34931 21403
rect 13645 21301 13679 21335
rect 17417 21301 17451 21335
rect 19165 21301 19199 21335
rect 23029 21301 23063 21335
rect 31309 21301 31343 21335
rect 32873 21301 32907 21335
rect 36461 21301 36495 21335
rect 11253 21097 11287 21131
rect 16773 21097 16807 21131
rect 21281 21097 21315 21131
rect 23121 21097 23155 21131
rect 25605 21097 25639 21131
rect 28641 21097 28675 21131
rect 3065 21029 3099 21063
rect 5273 21029 5307 21063
rect 19625 21029 19659 21063
rect 19993 21029 20027 21063
rect 24501 21029 24535 21063
rect 24593 21029 24627 21063
rect 24961 21029 24995 21063
rect 1409 20961 1443 20995
rect 1685 20961 1719 20995
rect 4353 20961 4387 20995
rect 4629 20961 4663 20995
rect 4813 20961 4847 20995
rect 5733 20961 5767 20995
rect 6285 20961 6319 20995
rect 6745 20961 6779 20995
rect 7205 20961 7239 20995
rect 7849 20961 7883 20995
rect 8401 20961 8435 20995
rect 8861 20961 8895 20995
rect 9689 20961 9723 20995
rect 9965 20961 9999 20995
rect 11805 20961 11839 20995
rect 12541 20961 12575 20995
rect 13093 20961 13127 20995
rect 13737 20961 13771 20995
rect 14197 20961 14231 20995
rect 15853 20961 15887 20995
rect 16405 20961 16439 20995
rect 17049 20961 17083 20995
rect 17509 20961 17543 20995
rect 18521 20961 18555 20995
rect 19441 20961 19475 20995
rect 19533 20961 19567 20995
rect 21097 20961 21131 20995
rect 21833 20961 21867 20995
rect 22385 20961 22419 20995
rect 23305 20961 23339 20995
rect 23489 20961 23523 20995
rect 24409 20961 24443 20995
rect 25421 20961 25455 20995
rect 26525 20961 26559 20995
rect 27629 20961 27663 20995
rect 28181 20961 28215 20995
rect 28365 20961 28399 20995
rect 29285 20961 29319 20995
rect 29837 20961 29871 20995
rect 30297 20961 30331 20995
rect 31125 20961 31159 20995
rect 31217 20961 31251 20995
rect 31585 20961 31619 20995
rect 32413 20961 32447 20995
rect 32781 20961 32815 20995
rect 32873 20961 32907 20995
rect 33425 20961 33459 20995
rect 34345 20961 34379 20995
rect 34713 20961 34747 20995
rect 35081 20961 35115 20995
rect 36093 20961 36127 20995
rect 36829 20961 36863 20995
rect 37841 20961 37875 20995
rect 38577 20961 38611 20995
rect 5825 20893 5859 20927
rect 8033 20893 8067 20927
rect 13461 20893 13495 20927
rect 19257 20893 19291 20927
rect 22569 20893 22603 20927
rect 24225 20893 24259 20927
rect 27537 20893 27571 20927
rect 33057 20893 33091 20927
rect 34529 20893 34563 20927
rect 36921 20893 36955 20927
rect 38669 20893 38703 20927
rect 11989 20825 12023 20859
rect 18705 20825 18739 20859
rect 29377 20825 29411 20859
rect 36369 20825 36403 20859
rect 37933 20825 37967 20859
rect 8953 20757 8987 20791
rect 26617 20757 26651 20791
rect 29653 20553 29687 20587
rect 3985 20485 4019 20519
rect 9045 20485 9079 20519
rect 13277 20485 13311 20519
rect 15301 20485 15335 20519
rect 28273 20485 28307 20519
rect 6285 20417 6319 20451
rect 7113 20417 7147 20451
rect 11437 20417 11471 20451
rect 12541 20417 12575 20451
rect 14565 20417 14599 20451
rect 17509 20417 17543 20451
rect 21557 20417 21591 20451
rect 24501 20417 24535 20451
rect 26249 20417 26283 20451
rect 33609 20485 33643 20519
rect 30665 20417 30699 20451
rect 32045 20417 32079 20451
rect 34253 20417 34287 20451
rect 35725 20417 35759 20451
rect 37749 20417 37783 20451
rect 1869 20349 1903 20383
rect 2697 20349 2731 20383
rect 2881 20349 2915 20383
rect 3249 20349 3283 20383
rect 3893 20349 3927 20383
rect 4445 20349 4479 20383
rect 4721 20349 4755 20383
rect 5549 20349 5583 20383
rect 5733 20349 5767 20383
rect 5825 20349 5859 20383
rect 6837 20349 6871 20383
rect 8953 20349 8987 20383
rect 9505 20349 9539 20383
rect 9873 20349 9907 20383
rect 11713 20349 11747 20383
rect 11897 20349 11931 20383
rect 13001 20349 13035 20383
rect 13369 20349 13403 20383
rect 15025 20349 15059 20383
rect 15301 20349 15335 20383
rect 16313 20349 16347 20383
rect 16589 20349 16623 20383
rect 16957 20349 16991 20383
rect 17325 20349 17359 20383
rect 17601 20349 17635 20383
rect 21097 20349 21131 20383
rect 21281 20349 21315 20383
rect 22109 20349 22143 20383
rect 22845 20349 22879 20383
rect 23029 20349 23063 20383
rect 23673 20349 23707 20383
rect 24777 20349 24811 20383
rect 25329 20349 25363 20383
rect 25973 20349 26007 20383
rect 28457 20349 28491 20383
rect 28549 20349 28583 20383
rect 29653 20349 29687 20383
rect 29745 20349 29779 20383
rect 30389 20349 30423 20383
rect 32505 20349 32539 20383
rect 33793 20349 33827 20383
rect 34161 20349 34195 20383
rect 35265 20349 35299 20383
rect 35817 20349 35851 20383
rect 36185 20349 36219 20383
rect 36369 20349 36403 20383
rect 36737 20349 36771 20383
rect 37473 20349 37507 20383
rect 10885 20281 10919 20315
rect 18429 20281 18463 20315
rect 25513 20281 25547 20315
rect 1961 20213 1995 20247
rect 8401 20213 8435 20247
rect 16129 20213 16163 20247
rect 17785 20213 17819 20247
rect 19717 20213 19751 20247
rect 22109 20213 22143 20247
rect 23857 20213 23891 20247
rect 27353 20213 27387 20247
rect 28641 20213 28675 20247
rect 29837 20213 29871 20247
rect 32689 20213 32723 20247
rect 38853 20213 38887 20247
rect 11989 20009 12023 20043
rect 12817 20009 12851 20043
rect 17417 20009 17451 20043
rect 22293 20009 22327 20043
rect 26801 20009 26835 20043
rect 3065 19941 3099 19975
rect 34621 19941 34655 19975
rect 1409 19873 1443 19907
rect 4077 19873 4111 19907
rect 4997 19873 5031 19907
rect 5273 19873 5307 19907
rect 5549 19873 5583 19907
rect 6009 19873 6043 19907
rect 6653 19873 6687 19907
rect 7757 19873 7791 19907
rect 9137 19873 9171 19907
rect 9689 19873 9723 19907
rect 10885 19873 10919 19907
rect 12909 19873 12943 19907
rect 13369 19873 13403 19907
rect 13553 19873 13587 19907
rect 14473 19873 14507 19907
rect 15301 19873 15335 19907
rect 15485 19873 15519 19907
rect 16957 19873 16991 19907
rect 17141 19873 17175 19907
rect 17693 19873 17727 19907
rect 18061 19873 18095 19907
rect 19165 19873 19199 19907
rect 19349 19873 19383 19907
rect 19625 19873 19659 19907
rect 20269 19873 20303 19907
rect 20913 19873 20947 19907
rect 23029 19873 23063 19907
rect 24685 19873 24719 19907
rect 25145 19873 25179 19907
rect 25421 19873 25455 19907
rect 25605 19873 25639 19907
rect 26525 19873 26559 19907
rect 26709 19873 26743 19907
rect 27537 19873 27571 19907
rect 28457 19873 28491 19907
rect 28549 19873 28583 19907
rect 29009 19873 29043 19907
rect 29745 19873 29779 19907
rect 30849 19873 30883 19907
rect 32965 19873 32999 19907
rect 33333 19873 33367 19907
rect 33517 19873 33551 19907
rect 33977 19873 34011 19907
rect 35173 19873 35207 19907
rect 35357 19873 35391 19907
rect 35449 19873 35483 19907
rect 35633 19873 35667 19907
rect 35909 19873 35943 19907
rect 36921 19873 36955 19907
rect 38117 19873 38151 19907
rect 38485 19873 38519 19907
rect 38669 19873 38703 19907
rect 1685 19805 1719 19839
rect 5365 19805 5399 19839
rect 7481 19805 7515 19839
rect 10609 19805 10643 19839
rect 18981 19805 19015 19839
rect 21189 19805 21223 19839
rect 23949 19737 23983 19771
rect 24041 19737 24075 19771
rect 29101 19805 29135 19839
rect 4169 19669 4203 19703
rect 9781 19669 9815 19703
rect 14657 19669 14691 19703
rect 15577 19669 15611 19703
rect 23213 19669 23247 19703
rect 27721 19669 27755 19703
rect 28457 19669 28491 19703
rect 29837 19669 29871 19703
rect 31033 19669 31067 19703
rect 32781 19669 32815 19703
rect 37105 19669 37139 19703
rect 1593 19465 1627 19499
rect 11529 19465 11563 19499
rect 15577 19465 15611 19499
rect 31493 19465 31527 19499
rect 35081 19465 35115 19499
rect 24041 19397 24075 19431
rect 7849 19329 7883 19363
rect 13737 19329 13771 19363
rect 22569 19329 22603 19363
rect 29561 19329 29595 19363
rect 1501 19261 1535 19295
rect 2133 19261 2167 19295
rect 3157 19261 3191 19295
rect 3341 19261 3375 19295
rect 3709 19261 3743 19295
rect 4261 19261 4295 19295
rect 5457 19261 5491 19295
rect 5825 19261 5859 19295
rect 7113 19261 7147 19295
rect 7665 19261 7699 19295
rect 7757 19261 7791 19295
rect 8493 19261 8527 19295
rect 9321 19261 9355 19295
rect 9597 19261 9631 19295
rect 10977 19261 11011 19295
rect 11437 19261 11471 19295
rect 12265 19261 12299 19295
rect 12817 19261 12851 19295
rect 13185 19261 13219 19295
rect 13553 19261 13587 19295
rect 14197 19261 14231 19295
rect 14473 19261 14507 19295
rect 16313 19261 16347 19295
rect 16405 19261 16439 19295
rect 17325 19261 17359 19295
rect 17417 19261 17451 19295
rect 18061 19261 18095 19295
rect 18705 19261 18739 19295
rect 18981 19261 19015 19295
rect 20821 19261 20855 19295
rect 22661 19261 22695 19295
rect 22753 19261 22787 19295
rect 23949 19261 23983 19295
rect 24685 19261 24719 19295
rect 25145 19261 25179 19295
rect 25421 19261 25455 19295
rect 25605 19261 25639 19295
rect 26341 19261 26375 19295
rect 27077 19261 27111 19295
rect 27353 19261 27387 19295
rect 28733 19261 28767 19295
rect 29285 19261 29319 19295
rect 31677 19261 31711 19295
rect 32045 19261 32079 19295
rect 32413 19261 32447 19295
rect 33885 19261 33919 19295
rect 34069 19261 34103 19295
rect 34897 19261 34931 19295
rect 35633 19261 35667 19295
rect 36185 19261 36219 19295
rect 36921 19261 36955 19295
rect 37197 19261 37231 19295
rect 38577 19261 38611 19295
rect 6009 19193 6043 19227
rect 16865 19193 16899 19227
rect 23213 19193 23247 19227
rect 2329 19125 2363 19159
rect 4077 19125 4111 19159
rect 12081 19125 12115 19159
rect 18245 19125 18279 19159
rect 20085 19125 20119 19159
rect 26525 19125 26559 19159
rect 30665 19125 30699 19159
rect 33885 19125 33919 19159
rect 35909 19125 35943 19159
rect 4813 18921 4847 18955
rect 15577 18921 15611 18955
rect 26709 18921 26743 18955
rect 8769 18853 8803 18887
rect 10241 18853 10275 18887
rect 14013 18853 14047 18887
rect 15301 18853 15335 18887
rect 20545 18853 20579 18887
rect 21465 18853 21499 18887
rect 21649 18853 21683 18887
rect 22017 18853 22051 18887
rect 22109 18853 22143 18887
rect 36921 18853 36955 18887
rect 2605 18785 2639 18819
rect 2697 18785 2731 18819
rect 2881 18785 2915 18819
rect 3249 18785 3283 18819
rect 3525 18785 3559 18819
rect 4629 18785 4663 18819
rect 5457 18785 5491 18819
rect 5733 18785 5767 18819
rect 6101 18785 6135 18819
rect 6837 18785 6871 18819
rect 7757 18785 7791 18819
rect 8217 18785 8251 18819
rect 8677 18785 8711 18819
rect 9801 18785 9835 18819
rect 12449 18785 12483 18819
rect 13277 18785 13311 18819
rect 13829 18785 13863 18819
rect 14473 18785 14507 18819
rect 15485 18785 15519 18819
rect 16773 18785 16807 18819
rect 18429 18785 18463 18819
rect 19349 18785 19383 18819
rect 19625 18785 19659 18819
rect 20085 18785 20119 18819
rect 20913 18785 20947 18819
rect 21557 18785 21591 18819
rect 22569 18785 22603 18819
rect 22753 18785 22787 18819
rect 22937 18785 22971 18819
rect 23673 18785 23707 18819
rect 24041 18785 24075 18819
rect 25237 18785 25271 18819
rect 25605 18785 25639 18819
rect 26525 18785 26559 18819
rect 27537 18785 27571 18819
rect 27813 18785 27847 18819
rect 28457 18785 28491 18819
rect 30021 18785 30055 18819
rect 30205 18785 30239 18819
rect 30481 18785 30515 18819
rect 30665 18785 30699 18819
rect 30941 18785 30975 18819
rect 32137 18785 32171 18819
rect 32505 18785 32539 18819
rect 32965 18785 32999 18819
rect 33793 18785 33827 18819
rect 34345 18785 34379 18819
rect 34529 18785 34563 18819
rect 35081 18785 35115 18819
rect 35817 18785 35851 18819
rect 36369 18785 36403 18819
rect 36737 18785 36771 18819
rect 37197 18785 37231 18819
rect 38301 18785 38335 18819
rect 38669 18785 38703 18819
rect 5917 18717 5951 18751
rect 7849 18717 7883 18751
rect 9689 18717 9723 18751
rect 10793 18717 10827 18751
rect 11069 18717 11103 18751
rect 13001 18717 13035 18751
rect 17049 18717 17083 18751
rect 18889 18717 18923 18751
rect 19993 18717 20027 18751
rect 21281 18717 21315 18751
rect 24133 18717 24167 18751
rect 24869 18717 24903 18751
rect 29561 18717 29595 18751
rect 34621 18717 34655 18751
rect 38761 18717 38795 18751
rect 19625 18649 19659 18683
rect 23489 18649 23523 18683
rect 25513 18649 25547 18683
rect 38117 18649 38151 18683
rect 2145 18581 2179 18615
rect 14657 18581 14691 18615
rect 21097 18581 21131 18615
rect 27353 18581 27387 18615
rect 28641 18581 28675 18615
rect 32229 18581 32263 18615
rect 9229 18377 9263 18411
rect 11437 18377 11471 18411
rect 12449 18377 12483 18411
rect 19625 18377 19659 18411
rect 19993 18377 20027 18411
rect 5549 18309 5583 18343
rect 6285 18309 6319 18343
rect 4905 18241 4939 18275
rect 11805 18241 11839 18275
rect 21557 18309 21591 18343
rect 22385 18309 22419 18343
rect 23949 18309 23983 18343
rect 29469 18309 29503 18343
rect 32965 18309 32999 18343
rect 35081 18309 35115 18343
rect 15209 18241 15243 18275
rect 18061 18241 18095 18275
rect 23857 18241 23891 18275
rect 27169 18241 27203 18275
rect 33609 18241 33643 18275
rect 34253 18241 34287 18275
rect 35725 18241 35759 18275
rect 38577 18241 38611 18275
rect 2789 18173 2823 18207
rect 3525 18173 3559 18207
rect 3801 18173 3835 18207
rect 4169 18173 4203 18207
rect 5273 18173 5307 18207
rect 5641 18173 5675 18207
rect 6469 18173 6503 18207
rect 7021 18173 7055 18207
rect 7205 18173 7239 18207
rect 7573 18173 7607 18207
rect 8217 18173 8251 18207
rect 8401 18173 8435 18207
rect 8585 18173 8619 18207
rect 9229 18173 9263 18207
rect 9321 18173 9355 18207
rect 9597 18173 9631 18207
rect 11621 18173 11655 18207
rect 11713 18173 11747 18207
rect 12357 18173 12391 18207
rect 12633 18173 12667 18207
rect 13461 18173 13495 18207
rect 14289 18173 14323 18207
rect 14933 18173 14967 18207
rect 17233 18173 17267 18207
rect 18337 18173 18371 18207
rect 19809 18173 19843 18207
rect 20177 18173 20211 18207
rect 20453 18173 20487 18207
rect 22569 18173 22603 18207
rect 22845 18173 22879 18207
rect 24593 18173 24627 18207
rect 25053 18173 25087 18207
rect 25329 18173 25363 18207
rect 25513 18173 25547 18207
rect 26525 18173 26559 18207
rect 26709 18173 26743 18207
rect 27813 18173 27847 18207
rect 28365 18173 28399 18207
rect 28641 18173 28675 18207
rect 29285 18173 29319 18207
rect 29837 18173 29871 18207
rect 30297 18173 30331 18207
rect 31309 18173 31343 18207
rect 32045 18173 32079 18207
rect 33149 18173 33183 18207
rect 33517 18173 33551 18207
rect 34161 18173 34195 18207
rect 34897 18173 34931 18207
rect 36001 18173 36035 18207
rect 38209 18173 38243 18207
rect 38393 18173 38427 18207
rect 38669 18173 38703 18207
rect 4261 18105 4295 18139
rect 13277 18105 13311 18139
rect 13829 18105 13863 18139
rect 26617 18105 26651 18139
rect 32137 18105 32171 18139
rect 37381 18105 37415 18139
rect 10701 18037 10735 18071
rect 12725 18037 12759 18071
rect 14381 18037 14415 18071
rect 16313 18037 16347 18071
rect 17417 18037 17451 18071
rect 27721 18037 27755 18071
rect 31493 18037 31527 18071
rect 9781 17833 9815 17867
rect 30941 17833 30975 17867
rect 32413 17833 32447 17867
rect 33701 17833 33735 17867
rect 3157 17765 3191 17799
rect 10885 17765 10919 17799
rect 20177 17765 20211 17799
rect 30021 17765 30055 17799
rect 1501 17697 1535 17731
rect 4077 17697 4111 17731
rect 4905 17697 4939 17731
rect 5365 17697 5399 17731
rect 5733 17697 5767 17731
rect 6101 17697 6135 17731
rect 6929 17697 6963 17731
rect 7113 17697 7147 17731
rect 7665 17697 7699 17731
rect 7941 17697 7975 17731
rect 8585 17697 8619 17731
rect 9689 17697 9723 17731
rect 10425 17697 10459 17731
rect 13921 17697 13955 17731
rect 14289 17697 14323 17731
rect 15301 17697 15335 17731
rect 17601 17697 17635 17731
rect 17693 17697 17727 17731
rect 18705 17697 18739 17731
rect 19717 17697 19751 17731
rect 21833 17697 21867 17731
rect 22109 17697 22143 17731
rect 22293 17697 22327 17731
rect 22477 17697 22511 17731
rect 22661 17697 22695 17731
rect 23857 17697 23891 17731
rect 24593 17697 24627 17731
rect 25053 17697 25087 17731
rect 25329 17697 25363 17731
rect 25513 17697 25547 17731
rect 26801 17697 26835 17731
rect 27077 17697 27111 17731
rect 27537 17697 27571 17731
rect 27721 17697 27755 17731
rect 28181 17697 28215 17731
rect 29285 17697 29319 17731
rect 29745 17697 29779 17731
rect 31125 17697 31159 17731
rect 31401 17697 31435 17731
rect 32321 17697 32355 17731
rect 32689 17697 32723 17731
rect 33517 17697 33551 17731
rect 34621 17697 34655 17731
rect 34805 17697 34839 17731
rect 35357 17697 35391 17731
rect 35633 17697 35667 17731
rect 36277 17697 36311 17731
rect 36829 17697 36863 17731
rect 38301 17697 38335 17731
rect 38577 17697 38611 17731
rect 1777 17629 1811 17663
rect 8677 17629 8711 17663
rect 10333 17629 10367 17663
rect 11345 17629 11379 17663
rect 11621 17629 11655 17663
rect 13645 17629 13679 17663
rect 15577 17629 15611 17663
rect 18613 17629 18647 17663
rect 19625 17629 19659 17663
rect 21373 17629 21407 17663
rect 29101 17629 29135 17663
rect 37841 17629 37875 17663
rect 6101 17561 6135 17595
rect 14289 17561 14323 17595
rect 23949 17561 23983 17595
rect 26617 17561 26651 17595
rect 38577 17561 38611 17595
rect 4169 17493 4203 17527
rect 8033 17493 8067 17527
rect 12909 17493 12943 17527
rect 16681 17493 16715 17527
rect 17877 17493 17911 17527
rect 18889 17493 18923 17527
rect 35725 17493 35759 17527
rect 36369 17493 36403 17527
rect 6929 17289 6963 17323
rect 9229 17289 9263 17323
rect 10241 17289 10275 17323
rect 11621 17289 11655 17323
rect 16589 17289 16623 17323
rect 27445 17289 27479 17323
rect 33517 17289 33551 17323
rect 38853 17289 38887 17323
rect 15853 17221 15887 17255
rect 18245 17221 18279 17255
rect 22661 17221 22695 17255
rect 31585 17221 31619 17255
rect 3065 17153 3099 17187
rect 6193 17153 6227 17187
rect 9965 17153 9999 17187
rect 11345 17153 11379 17187
rect 13645 17153 13679 17187
rect 18889 17153 18923 17187
rect 19165 17153 19199 17187
rect 32413 17153 32447 17187
rect 36001 17153 36035 17187
rect 1685 17085 1719 17119
rect 2237 17085 2271 17119
rect 2421 17085 2455 17119
rect 3249 17085 3283 17119
rect 3433 17085 3467 17119
rect 3985 17085 4019 17119
rect 4905 17085 4939 17119
rect 5457 17085 5491 17119
rect 5549 17085 5583 17119
rect 6285 17085 6319 17119
rect 6837 17085 6871 17119
rect 7849 17085 7883 17119
rect 8125 17085 8159 17119
rect 10057 17085 10091 17119
rect 11437 17085 11471 17119
rect 12725 17085 12759 17119
rect 12909 17085 12943 17119
rect 13461 17085 13495 17119
rect 14197 17085 14231 17119
rect 14933 17085 14967 17119
rect 15393 17085 15427 17119
rect 15761 17085 15795 17119
rect 16681 17085 16715 17119
rect 17233 17085 17267 17119
rect 18061 17085 18095 17119
rect 21557 17085 21591 17119
rect 21741 17085 21775 17119
rect 22109 17085 22143 17119
rect 22477 17085 22511 17119
rect 24133 17085 24167 17119
rect 24869 17085 24903 17119
rect 26157 17085 26191 17119
rect 26249 17085 26283 17119
rect 26525 17085 26559 17119
rect 26709 17085 26743 17119
rect 27997 17085 28031 17119
rect 28089 17085 28123 17119
rect 28365 17085 28399 17119
rect 28457 17085 28491 17119
rect 29561 17085 29595 17119
rect 30021 17085 30055 17119
rect 30297 17085 30331 17119
rect 30481 17085 30515 17119
rect 31401 17085 31435 17119
rect 32137 17085 32171 17119
rect 34897 17085 34931 17119
rect 35357 17085 35391 17119
rect 35725 17085 35759 17119
rect 36553 17085 36587 17119
rect 36829 17085 36863 17119
rect 38669 17085 38703 17119
rect 25513 17017 25547 17051
rect 1685 16949 1719 16983
rect 14381 16949 14415 16983
rect 20453 16949 20487 16983
rect 24317 16949 24351 16983
rect 24961 16949 24995 16983
rect 30481 16949 30515 16983
rect 37933 16949 37967 16983
rect 3433 16745 3467 16779
rect 5457 16745 5491 16779
rect 11529 16745 11563 16779
rect 14197 16745 14231 16779
rect 18613 16745 18647 16779
rect 21281 16745 21315 16779
rect 34989 16745 35023 16779
rect 35633 16745 35667 16779
rect 37841 16745 37875 16779
rect 2789 16677 2823 16711
rect 8033 16677 8067 16711
rect 8585 16677 8619 16711
rect 32137 16677 32171 16711
rect 2597 16609 2631 16643
rect 2697 16609 2731 16643
rect 3341 16609 3375 16643
rect 4353 16609 4387 16643
rect 6193 16609 6227 16643
rect 6561 16609 6595 16643
rect 7205 16609 7239 16643
rect 7941 16609 7975 16643
rect 8125 16609 8159 16643
rect 10149 16609 10183 16643
rect 10425 16609 10459 16643
rect 15485 16609 15519 16643
rect 15577 16609 15611 16643
rect 17417 16609 17451 16643
rect 17693 16609 17727 16643
rect 18429 16609 18463 16643
rect 19165 16609 19199 16643
rect 19809 16609 19843 16643
rect 20177 16609 20211 16643
rect 21465 16609 21499 16643
rect 22017 16609 22051 16643
rect 22753 16609 22787 16643
rect 23765 16609 23799 16643
rect 24317 16609 24351 16643
rect 24869 16609 24903 16643
rect 25329 16609 25363 16643
rect 25789 16609 25823 16643
rect 25881 16609 25915 16643
rect 27077 16609 27111 16643
rect 27261 16609 27295 16643
rect 27445 16609 27479 16643
rect 28641 16609 28675 16643
rect 28825 16609 28859 16643
rect 29009 16609 29043 16643
rect 29193 16609 29227 16643
rect 29377 16609 29411 16643
rect 30205 16609 30239 16643
rect 30389 16609 30423 16643
rect 30849 16609 30883 16643
rect 32827 16609 32861 16643
rect 32965 16609 32999 16643
rect 33609 16609 33643 16643
rect 34805 16609 34839 16643
rect 35633 16609 35667 16643
rect 36277 16609 36311 16643
rect 36553 16609 36587 16643
rect 37749 16609 37783 16643
rect 38301 16609 38335 16643
rect 38577 16609 38611 16643
rect 4077 16541 4111 16575
rect 6285 16541 6319 16575
rect 12817 16541 12851 16575
rect 13093 16541 13127 16575
rect 16957 16541 16991 16575
rect 17969 16541 18003 16575
rect 19349 16541 19383 16575
rect 22109 16541 22143 16575
rect 24777 16541 24811 16575
rect 32689 16541 32723 16575
rect 22937 16473 22971 16507
rect 23673 16473 23707 16507
rect 26893 16473 26927 16507
rect 30849 16473 30883 16507
rect 2421 16405 2455 16439
rect 15761 16405 15795 16439
rect 28181 16405 28215 16439
rect 33793 16405 33827 16439
rect 2973 16201 3007 16235
rect 6193 16201 6227 16235
rect 7113 16201 7147 16235
rect 29929 16201 29963 16235
rect 36921 16201 36955 16235
rect 38853 16201 38887 16235
rect 13553 16133 13587 16167
rect 26433 16133 26467 16167
rect 3617 16065 3651 16099
rect 4629 16065 4663 16099
rect 4905 16065 4939 16099
rect 6837 16065 6871 16099
rect 8401 16065 8435 16099
rect 10517 16065 10551 16099
rect 11069 16065 11103 16099
rect 18337 16065 18371 16099
rect 21005 16065 21039 16099
rect 25789 16065 25823 16099
rect 27353 16065 27387 16099
rect 27997 16065 28031 16099
rect 30481 16065 30515 16099
rect 31171 16065 31205 16099
rect 37473 16065 37507 16099
rect 1409 15997 1443 16031
rect 1685 15997 1719 16031
rect 3709 15997 3743 16031
rect 6929 15997 6963 16031
rect 8677 15997 8711 16031
rect 10609 15997 10643 16031
rect 11529 15997 11563 16031
rect 12909 15997 12943 16031
rect 13277 15997 13311 16031
rect 13645 15997 13679 16031
rect 14565 15997 14599 16031
rect 14841 15997 14875 16031
rect 16681 15997 16715 16031
rect 18061 15997 18095 16031
rect 20545 15997 20579 16031
rect 20729 15997 20763 16031
rect 21925 15997 21959 16031
rect 22109 15997 22143 16031
rect 22293 15997 22327 16031
rect 22569 15997 22603 16031
rect 22845 15997 22879 16031
rect 24133 15997 24167 16031
rect 24409 15997 24443 16031
rect 24501 15997 24535 16031
rect 24685 15997 24719 16031
rect 24961 15997 24995 16031
rect 26157 15997 26191 16031
rect 26433 15997 26467 16031
rect 27721 15997 27755 16031
rect 28089 15997 28123 16031
rect 29745 15997 29779 16031
rect 31033 15997 31067 16031
rect 31309 15997 31343 16031
rect 31953 15997 31987 16031
rect 32873 15997 32907 16031
rect 33425 15997 33459 16031
rect 33701 15997 33735 16031
rect 35817 15997 35851 16031
rect 36001 15997 36035 16031
rect 36185 15997 36219 16031
rect 36829 15997 36863 16031
rect 37749 15997 37783 16031
rect 4169 15929 4203 15963
rect 10057 15929 10091 15963
rect 21465 15929 21499 15963
rect 23673 15929 23707 15963
rect 35357 15929 35391 15963
rect 11621 15861 11655 15895
rect 15945 15861 15979 15895
rect 16865 15861 16899 15895
rect 19441 15861 19475 15895
rect 32137 15861 32171 15895
rect 32965 15861 32999 15895
rect 5457 15657 5491 15691
rect 14105 15657 14139 15691
rect 21097 15657 21131 15691
rect 26617 15657 26651 15691
rect 29285 15657 29319 15691
rect 31125 15657 31159 15691
rect 37841 15657 37875 15691
rect 39037 15657 39071 15691
rect 2973 15589 3007 15623
rect 2513 15521 2547 15555
rect 3893 15521 3927 15555
rect 6469 15521 6503 15555
rect 8585 15521 8619 15555
rect 9689 15521 9723 15555
rect 10425 15521 10459 15555
rect 10885 15521 10919 15555
rect 11069 15521 11103 15555
rect 11713 15521 11747 15555
rect 12265 15521 12299 15555
rect 12725 15521 12759 15555
rect 13001 15521 13035 15555
rect 16037 15521 16071 15555
rect 16405 15521 16439 15555
rect 16589 15521 16623 15555
rect 17325 15521 17359 15555
rect 17509 15521 17543 15555
rect 17969 15521 18003 15555
rect 18705 15521 18739 15555
rect 21005 15521 21039 15555
rect 22109 15521 22143 15555
rect 22293 15521 22327 15555
rect 22569 15521 22603 15555
rect 22661 15521 22695 15555
rect 23029 15521 23063 15555
rect 24133 15521 24167 15555
rect 24225 15521 24259 15555
rect 24501 15521 24535 15555
rect 24593 15521 24627 15555
rect 24961 15521 24995 15555
rect 25513 15521 25547 15555
rect 26525 15521 26559 15555
rect 27169 15521 27203 15555
rect 27905 15521 27939 15555
rect 29009 15521 29043 15555
rect 29653 15521 29687 15555
rect 29837 15521 29871 15555
rect 30205 15521 30239 15555
rect 30941 15521 30975 15555
rect 32597 15521 32631 15555
rect 32689 15521 32723 15555
rect 33057 15521 33091 15555
rect 33793 15521 33827 15555
rect 35817 15521 35851 15555
rect 36185 15521 36219 15555
rect 36461 15521 36495 15555
rect 36829 15521 36863 15555
rect 37749 15521 37783 15555
rect 38209 15521 38243 15555
rect 38945 15521 38979 15555
rect 2421 15453 2455 15487
rect 4077 15453 4111 15487
rect 4353 15453 4387 15487
rect 6745 15453 6779 15487
rect 8125 15453 8159 15487
rect 10517 15453 10551 15487
rect 15669 15453 15703 15487
rect 17693 15453 17727 15487
rect 18981 15453 19015 15487
rect 21649 15453 21683 15487
rect 23581 15453 23615 15487
rect 27997 15453 28031 15487
rect 33517 15453 33551 15487
rect 36093 15453 36127 15487
rect 3709 15385 3743 15419
rect 27445 15385 27479 15419
rect 8769 15317 8803 15351
rect 9781 15317 9815 15351
rect 20269 15317 20303 15351
rect 25697 15317 25731 15351
rect 35081 15317 35115 15351
rect 2789 15113 2823 15147
rect 5641 15113 5675 15147
rect 21281 15113 21315 15147
rect 38761 15113 38795 15147
rect 8493 15045 8527 15079
rect 13369 15045 13403 15079
rect 25053 15045 25087 15079
rect 28457 15045 28491 15079
rect 33149 15045 33183 15079
rect 1685 14977 1719 15011
rect 7573 14977 7607 15011
rect 13829 14977 13863 15011
rect 16405 14977 16439 15011
rect 18981 14977 19015 15011
rect 36185 14977 36219 15011
rect 38485 14977 38519 15011
rect 1409 14909 1443 14943
rect 4077 14909 4111 14943
rect 4353 14909 4387 14943
rect 7297 14909 7331 14943
rect 7481 14909 7515 14943
rect 8585 14909 8619 14943
rect 9045 14909 9079 14943
rect 9229 14909 9263 14943
rect 9597 14909 9631 14943
rect 10333 14909 10367 14943
rect 10793 14909 10827 14943
rect 11529 14909 11563 14943
rect 12449 14909 12483 14943
rect 13553 14909 13587 14943
rect 13645 14909 13679 14943
rect 14289 14909 14323 14943
rect 14657 14909 14691 14943
rect 15853 14909 15887 14943
rect 16497 14909 16531 14943
rect 16865 14909 16899 14943
rect 18061 14909 18095 14943
rect 18889 14909 18923 14943
rect 19349 14909 19383 14943
rect 19809 14909 19843 14943
rect 19993 14909 20027 14943
rect 20729 14909 20763 14943
rect 21189 14909 21223 14943
rect 21833 14909 21867 14943
rect 22293 14909 22327 14943
rect 23673 14909 23707 14943
rect 24025 14909 24059 14943
rect 24869 14909 24903 14943
rect 25605 14909 25639 14943
rect 26341 14909 26375 14943
rect 26617 14909 26651 14943
rect 27629 14909 27663 14943
rect 28089 14909 28123 14943
rect 28457 14909 28491 14943
rect 29745 14909 29779 14943
rect 29929 14909 29963 14943
rect 30297 14909 30331 14943
rect 32321 14909 32355 14943
rect 32873 14909 32907 14943
rect 33149 14909 33183 14943
rect 34069 14909 34103 14943
rect 35265 14909 35299 14943
rect 35725 14909 35759 14943
rect 36277 14909 36311 14943
rect 36461 14909 36495 14943
rect 36921 14909 36955 14943
rect 37749 14909 37783 14943
rect 38577 14909 38611 14943
rect 22569 14841 22603 14875
rect 23857 14841 23891 14875
rect 24409 14841 24443 14875
rect 31033 14841 31067 14875
rect 31309 14841 31343 14875
rect 31401 14841 31435 14875
rect 31769 14841 31803 14875
rect 10977 14773 11011 14807
rect 11713 14773 11747 14807
rect 12633 14773 12667 14807
rect 18245 14773 18279 14807
rect 23949 14773 23983 14807
rect 25697 14773 25731 14807
rect 29561 14773 29595 14807
rect 31217 14773 31251 14807
rect 34253 14773 34287 14807
rect 37933 14773 37967 14807
rect 2053 14569 2087 14603
rect 11621 14569 11655 14603
rect 16681 14569 16715 14603
rect 20085 14569 20119 14603
rect 23949 14569 23983 14603
rect 24041 14569 24075 14603
rect 26617 14569 26651 14603
rect 28273 14569 28307 14603
rect 30573 14569 30607 14603
rect 37105 14569 37139 14603
rect 4813 14501 4847 14535
rect 24133 14501 24167 14535
rect 30021 14501 30055 14535
rect 38117 14501 38151 14535
rect 38485 14501 38519 14535
rect 2237 14433 2271 14467
rect 2513 14433 2547 14467
rect 3249 14433 3283 14467
rect 4353 14433 4387 14467
rect 4629 14433 4663 14467
rect 8401 14433 8435 14467
rect 8585 14433 8619 14467
rect 10241 14433 10275 14467
rect 10517 14433 10551 14467
rect 13461 14433 13495 14467
rect 13829 14433 13863 14467
rect 14473 14433 14507 14467
rect 15577 14433 15611 14467
rect 19889 14433 19923 14467
rect 23029 14433 23063 14467
rect 23765 14433 23799 14467
rect 25421 14433 25455 14467
rect 25605 14433 25639 14467
rect 25789 14433 25823 14467
rect 26709 14433 26743 14467
rect 27077 14433 27111 14467
rect 28089 14433 28123 14467
rect 29285 14433 29319 14467
rect 29837 14433 29871 14467
rect 30481 14433 30515 14467
rect 30941 14433 30975 14467
rect 32597 14433 32631 14467
rect 32965 14433 32999 14467
rect 34069 14433 34103 14467
rect 34253 14433 34287 14467
rect 34437 14433 34471 14467
rect 34621 14433 34655 14467
rect 34897 14433 34931 14467
rect 37933 14433 37967 14467
rect 38025 14433 38059 14467
rect 38945 14433 38979 14467
rect 5917 14365 5951 14399
rect 6193 14365 6227 14399
rect 8677 14365 8711 14399
rect 13093 14365 13127 14399
rect 15301 14365 15335 14399
rect 17785 14365 17819 14399
rect 18061 14365 18095 14399
rect 20913 14365 20947 14399
rect 21189 14365 21223 14399
rect 24501 14365 24535 14399
rect 27537 14365 27571 14399
rect 29101 14365 29135 14399
rect 33057 14365 33091 14399
rect 33609 14365 33643 14399
rect 35541 14365 35575 14399
rect 35817 14365 35851 14399
rect 37749 14365 37783 14399
rect 13737 14297 13771 14331
rect 25237 14297 25271 14331
rect 32413 14297 32447 14331
rect 3433 14229 3467 14263
rect 7481 14229 7515 14263
rect 14657 14229 14691 14263
rect 19349 14229 19383 14263
rect 22293 14229 22327 14263
rect 23213 14229 23247 14263
rect 39037 14229 39071 14263
rect 14749 14025 14783 14059
rect 25053 14025 25087 14059
rect 28641 14025 28675 14059
rect 29285 14025 29319 14059
rect 34437 14025 34471 14059
rect 3801 13957 3835 13991
rect 8309 13957 8343 13991
rect 16497 13957 16531 13991
rect 18337 13957 18371 13991
rect 1593 13889 1627 13923
rect 1869 13889 1903 13923
rect 4629 13889 4663 13923
rect 5273 13889 5307 13923
rect 17325 13889 17359 13923
rect 21189 13889 21223 13923
rect 23949 13889 23983 13923
rect 26065 13889 26099 13923
rect 29285 13889 29319 13923
rect 29837 13889 29871 13923
rect 33149 13889 33183 13923
rect 35449 13889 35483 13923
rect 36185 13889 36219 13923
rect 37013 13889 37047 13923
rect 3985 13821 4019 13855
rect 4169 13821 4203 13855
rect 4537 13821 4571 13855
rect 5365 13821 5399 13855
rect 5825 13821 5859 13855
rect 7205 13821 7239 13855
rect 7389 13821 7423 13855
rect 7573 13821 7607 13855
rect 8217 13821 8251 13855
rect 8677 13821 8711 13855
rect 9229 13821 9263 13855
rect 9597 13821 9631 13855
rect 10149 13821 10183 13855
rect 11161 13821 11195 13855
rect 11529 13821 11563 13855
rect 11897 13821 11931 13855
rect 12541 13821 12575 13855
rect 12817 13821 12851 13855
rect 14197 13821 14231 13855
rect 14657 13821 14691 13855
rect 15301 13821 15335 13855
rect 15669 13821 15703 13855
rect 16497 13821 16531 13855
rect 16865 13821 16899 13855
rect 18429 13821 18463 13855
rect 18705 13821 18739 13855
rect 19257 13821 19291 13855
rect 19625 13821 19659 13855
rect 20085 13821 20119 13855
rect 20821 13821 20855 13855
rect 21281 13821 21315 13855
rect 21649 13821 21683 13855
rect 21925 13821 21959 13855
rect 22293 13821 22327 13855
rect 23673 13821 23707 13855
rect 25789 13821 25823 13855
rect 28457 13821 28491 13855
rect 29653 13821 29687 13855
rect 29929 13821 29963 13855
rect 30573 13821 30607 13855
rect 30757 13821 30791 13855
rect 31401 13821 31435 13855
rect 31861 13821 31895 13855
rect 32505 13821 32539 13855
rect 33057 13821 33091 13855
rect 33517 13821 33551 13855
rect 33793 13821 33827 13855
rect 34621 13821 34655 13855
rect 35633 13821 35667 13855
rect 36645 13821 36679 13855
rect 37381 13821 37415 13855
rect 37565 13821 37599 13855
rect 37933 13821 37967 13855
rect 38301 13821 38335 13855
rect 35725 13753 35759 13787
rect 35817 13753 35851 13787
rect 2973 13685 3007 13719
rect 27169 13685 27203 13719
rect 31953 13685 31987 13719
rect 7205 13481 7239 13515
rect 16681 13481 16715 13515
rect 18245 13481 18279 13515
rect 19809 13481 19843 13515
rect 21465 13481 21499 13515
rect 24409 13481 24443 13515
rect 28549 13481 28583 13515
rect 33701 13481 33735 13515
rect 36645 13481 36679 13515
rect 3249 13413 3283 13447
rect 25605 13413 25639 13447
rect 36829 13413 36863 13447
rect 1777 13345 1811 13379
rect 2789 13345 2823 13379
rect 4261 13345 4295 13379
rect 7113 13345 7147 13379
rect 7665 13345 7699 13379
rect 8309 13345 8343 13379
rect 8861 13345 8895 13379
rect 9873 13345 9907 13379
rect 10241 13345 10275 13379
rect 11529 13345 11563 13379
rect 11805 13345 11839 13379
rect 11989 13345 12023 13379
rect 12909 13345 12943 13379
rect 13645 13345 13679 13379
rect 14105 13345 14139 13379
rect 15301 13345 15335 13379
rect 16221 13345 16255 13379
rect 16773 13345 16807 13379
rect 17141 13345 17175 13379
rect 18153 13345 18187 13379
rect 18705 13345 18739 13379
rect 19717 13345 19751 13379
rect 21373 13345 21407 13379
rect 22017 13345 22051 13379
rect 22569 13345 22603 13379
rect 23213 13345 23247 13379
rect 24317 13345 24351 13379
rect 24869 13345 24903 13379
rect 25513 13345 25547 13379
rect 26525 13345 26559 13379
rect 27445 13345 27479 13379
rect 29469 13345 29503 13379
rect 29653 13345 29687 13379
rect 30389 13345 30423 13379
rect 30573 13345 30607 13379
rect 30941 13345 30975 13379
rect 31309 13345 31343 13379
rect 32689 13345 32723 13379
rect 33057 13345 33091 13379
rect 33885 13345 33919 13379
rect 34805 13345 34839 13379
rect 34989 13345 35023 13379
rect 35449 13345 35483 13379
rect 35725 13345 35759 13379
rect 36737 13345 36771 13379
rect 37749 13345 37783 13379
rect 38117 13345 38151 13379
rect 38577 13345 38611 13379
rect 1685 13277 1719 13311
rect 2697 13277 2731 13311
rect 4997 13277 5031 13311
rect 5273 13277 5307 13311
rect 12265 13277 12299 13311
rect 17601 13277 17635 13311
rect 18981 13277 19015 13311
rect 22753 13277 22787 13311
rect 27169 13277 27203 13311
rect 30021 13277 30055 13311
rect 32229 13277 32263 13311
rect 34069 13277 34103 13311
rect 34437 13277 34471 13311
rect 36461 13277 36495 13311
rect 37197 13277 37231 13311
rect 4445 13209 4479 13243
rect 15485 13209 15519 13243
rect 29285 13209 29319 13243
rect 32965 13209 32999 13243
rect 38577 13209 38611 13243
rect 1961 13141 1995 13175
rect 6561 13141 6595 13175
rect 8401 13141 8435 13175
rect 9781 13141 9815 13175
rect 13001 13141 13035 13175
rect 14289 13141 14323 13175
rect 16037 13141 16071 13175
rect 23305 13141 23339 13175
rect 26617 13141 26651 13175
rect 2789 12937 2823 12971
rect 5089 12937 5123 12971
rect 5917 12937 5951 12971
rect 16865 12937 16899 12971
rect 18337 12937 18371 12971
rect 32965 12937 32999 12971
rect 36369 12937 36403 12971
rect 37197 12937 37231 12971
rect 9229 12869 9263 12903
rect 14381 12869 14415 12903
rect 25881 12869 25915 12903
rect 27537 12869 27571 12903
rect 31493 12869 31527 12903
rect 38761 12869 38795 12903
rect 1685 12801 1719 12835
rect 5641 12801 5675 12835
rect 6929 12801 6963 12835
rect 11897 12801 11931 12835
rect 19349 12801 19383 12835
rect 23949 12801 23983 12835
rect 28089 12801 28123 12835
rect 29285 12801 29319 12835
rect 30849 12801 30883 12835
rect 33241 12801 33275 12835
rect 36921 12801 36955 12835
rect 1409 12733 1443 12767
rect 3525 12733 3559 12767
rect 3801 12733 3835 12767
rect 5733 12733 5767 12767
rect 6837 12733 6871 12767
rect 7665 12733 7699 12767
rect 7941 12733 7975 12767
rect 8217 12733 8251 12767
rect 9137 12733 9171 12767
rect 9873 12733 9907 12767
rect 10977 12733 11011 12767
rect 11253 12733 11287 12767
rect 11437 12733 11471 12767
rect 12449 12733 12483 12767
rect 12909 12733 12943 12767
rect 13093 12733 13127 12767
rect 13277 12733 13311 12767
rect 14473 12733 14507 12767
rect 14749 12733 14783 12767
rect 15117 12733 15151 12767
rect 15669 12733 15703 12767
rect 16221 12733 16255 12767
rect 16681 12733 16715 12767
rect 18889 12733 18923 12767
rect 18981 12733 19015 12767
rect 19257 12733 19291 12767
rect 19993 12733 20027 12767
rect 20453 12733 20487 12767
rect 21281 12733 21315 12767
rect 21557 12733 21591 12767
rect 23673 12733 23707 12767
rect 25789 12733 25823 12767
rect 26433 12733 26467 12767
rect 27261 12733 27295 12767
rect 27997 12733 28031 12767
rect 29469 12733 29503 12767
rect 31125 12733 31159 12767
rect 31493 12733 31527 12767
rect 32229 12733 32263 12767
rect 33149 12733 33183 12767
rect 33425 12733 33459 12767
rect 35265 12733 35299 12767
rect 35449 12733 35483 12767
rect 35725 12733 35759 12767
rect 36277 12733 36311 12767
rect 37013 12733 37047 12767
rect 37933 12733 37967 12767
rect 38301 12733 38335 12767
rect 38853 12733 38887 12767
rect 8677 12665 8711 12699
rect 29653 12665 29687 12699
rect 30021 12665 30055 12699
rect 33609 12665 33643 12699
rect 33977 12665 34011 12699
rect 19993 12597 20027 12631
rect 22661 12597 22695 12631
rect 25053 12597 25087 12631
rect 26525 12597 26559 12631
rect 29561 12597 29595 12631
rect 32413 12597 32447 12631
rect 33517 12597 33551 12631
rect 17877 12393 17911 12427
rect 18613 12393 18647 12427
rect 23765 12393 23799 12427
rect 26617 12393 26651 12427
rect 28733 12393 28767 12427
rect 29469 12393 29503 12427
rect 32137 12393 32171 12427
rect 33149 12393 33183 12427
rect 3525 12325 3559 12359
rect 8585 12325 8619 12359
rect 19165 12325 19199 12359
rect 25237 12325 25271 12359
rect 2053 12257 2087 12291
rect 2789 12257 2823 12291
rect 3341 12257 3375 12291
rect 7389 12257 7423 12291
rect 7941 12257 7975 12291
rect 8125 12257 8159 12291
rect 10149 12257 10183 12291
rect 10333 12257 10367 12291
rect 10517 12257 10551 12291
rect 11805 12257 11839 12291
rect 11989 12257 12023 12291
rect 12173 12257 12207 12291
rect 15301 12257 15335 12291
rect 15853 12257 15887 12291
rect 16037 12257 16071 12291
rect 16681 12257 16715 12291
rect 17233 12257 17267 12291
rect 17693 12257 17727 12291
rect 18429 12257 18463 12291
rect 19809 12257 19843 12291
rect 20177 12257 20211 12291
rect 20361 12257 20395 12291
rect 21281 12257 21315 12291
rect 21925 12257 21959 12291
rect 22293 12257 22327 12291
rect 22661 12257 22695 12291
rect 23213 12257 23247 12291
rect 23673 12257 23707 12291
rect 24685 12257 24719 12291
rect 24777 12257 24811 12291
rect 25697 12257 25731 12291
rect 26525 12257 26559 12291
rect 27169 12257 27203 12291
rect 27813 12257 27847 12291
rect 28549 12257 28583 12291
rect 29285 12257 29319 12291
rect 30205 12257 30239 12291
rect 30665 12257 30699 12291
rect 31033 12257 31067 12291
rect 5181 12189 5215 12223
rect 5457 12189 5491 12223
rect 13093 12189 13127 12223
rect 13369 12189 13403 12223
rect 15393 12189 15427 12223
rect 19901 12189 19935 12223
rect 25789 12189 25823 12223
rect 31401 12189 31435 12223
rect 36277 12325 36311 12359
rect 36645 12325 36679 12359
rect 32229 12257 32263 12291
rect 32965 12257 32999 12291
rect 34161 12257 34195 12291
rect 34621 12257 34655 12291
rect 36093 12257 36127 12291
rect 36185 12257 36219 12291
rect 38117 12257 38151 12291
rect 38577 12257 38611 12291
rect 33885 12189 33919 12223
rect 35909 12189 35943 12223
rect 38761 12189 38795 12223
rect 9965 12121 9999 12155
rect 11621 12121 11655 12155
rect 21557 12121 21591 12155
rect 27997 12121 28031 12155
rect 30757 12121 30791 12155
rect 32137 12121 32171 12155
rect 34621 12121 34655 12155
rect 38025 12121 38059 12155
rect 2237 12053 2271 12087
rect 6745 12053 6779 12087
rect 14473 12053 14507 12087
rect 27261 12053 27295 12087
rect 30021 12053 30055 12087
rect 32413 12053 32447 12087
rect 4629 11849 4663 11883
rect 6193 11849 6227 11883
rect 7205 11849 7239 11883
rect 19809 11849 19843 11883
rect 21465 11849 21499 11883
rect 23765 11849 23799 11883
rect 27537 11849 27571 11883
rect 30389 11849 30423 11883
rect 38945 11849 38979 11883
rect 12725 11781 12759 11815
rect 14657 11781 14691 11815
rect 29745 11781 29779 11815
rect 32505 11781 32539 11815
rect 3065 11713 3099 11747
rect 8953 11713 8987 11747
rect 10517 11713 10551 11747
rect 11437 11713 11471 11747
rect 15577 11713 15611 11747
rect 19257 11713 19291 11747
rect 20269 11713 20303 11747
rect 24409 11713 24443 11747
rect 25605 11713 25639 11747
rect 26433 11713 26467 11747
rect 31217 11713 31251 11747
rect 3341 11645 3375 11679
rect 6101 11645 6135 11679
rect 7113 11645 7147 11679
rect 8033 11645 8067 11679
rect 8217 11645 8251 11679
rect 8493 11645 8527 11679
rect 9597 11645 9631 11679
rect 9873 11645 9907 11679
rect 10149 11645 10183 11679
rect 11345 11645 11379 11679
rect 11713 11645 11747 11679
rect 12909 11645 12943 11679
rect 13093 11645 13127 11679
rect 13277 11645 13311 11679
rect 13921 11645 13955 11679
rect 14749 11645 14783 11679
rect 15117 11645 15151 11679
rect 16221 11645 16255 11679
rect 16589 11645 16623 11679
rect 17141 11645 17175 11679
rect 18521 11645 18555 11679
rect 19073 11645 19107 11679
rect 20361 11645 20395 11679
rect 20729 11645 20763 11679
rect 20913 11645 20947 11679
rect 21373 11645 21407 11679
rect 22569 11645 22603 11679
rect 23673 11645 23707 11679
rect 24501 11645 24535 11679
rect 24961 11645 24995 11679
rect 25053 11645 25087 11679
rect 26157 11645 26191 11679
rect 28549 11645 28583 11679
rect 29653 11645 29687 11679
rect 30297 11645 30331 11679
rect 30941 11645 30975 11679
rect 33609 11645 33643 11679
rect 33793 11645 33827 11679
rect 33977 11645 34011 11679
rect 35357 11645 35391 11679
rect 35541 11645 35575 11679
rect 35909 11645 35943 11679
rect 36001 11645 36035 11679
rect 36829 11645 36863 11679
rect 37013 11645 37047 11679
rect 37381 11645 37415 11679
rect 37565 11645 37599 11679
rect 37749 11645 37783 11679
rect 38761 11645 38795 11679
rect 17325 11577 17359 11611
rect 33149 11577 33183 11611
rect 38301 11577 38335 11611
rect 14013 11509 14047 11543
rect 22753 11509 22787 11543
rect 28641 11509 28675 11543
rect 35173 11509 35207 11543
rect 18705 11305 18739 11339
rect 31493 11305 31527 11339
rect 32229 11305 32263 11339
rect 12633 11237 12667 11271
rect 20361 11237 20395 11271
rect 30665 11237 30699 11271
rect 36185 11237 36219 11271
rect 36369 11237 36403 11271
rect 36553 11237 36587 11271
rect 36921 11237 36955 11271
rect 38853 11237 38887 11271
rect 2789 11169 2823 11203
rect 3249 11169 3283 11203
rect 4629 11169 4663 11203
rect 5365 11169 5399 11203
rect 5917 11169 5951 11203
rect 6285 11169 6319 11203
rect 6653 11169 6687 11203
rect 6929 11169 6963 11203
rect 7665 11169 7699 11203
rect 8033 11169 8067 11203
rect 8401 11169 8435 11203
rect 9781 11169 9815 11203
rect 10057 11169 10091 11203
rect 10425 11169 10459 11203
rect 10885 11169 10919 11203
rect 11621 11169 11655 11203
rect 12081 11169 12115 11203
rect 12357 11169 12391 11203
rect 13553 11169 13587 11203
rect 13921 11169 13955 11203
rect 14565 11169 14599 11203
rect 14657 11169 14691 11203
rect 15301 11169 15335 11203
rect 16221 11169 16255 11203
rect 18521 11169 18555 11203
rect 18981 11169 19015 11203
rect 19901 11169 19935 11203
rect 20177 11169 20211 11203
rect 21557 11169 21591 11203
rect 21971 11169 22005 11203
rect 22845 11169 22879 11203
rect 22937 11169 22971 11203
rect 23305 11169 23339 11203
rect 24777 11169 24811 11203
rect 25329 11169 25363 11203
rect 25513 11169 25547 11203
rect 26617 11169 26651 11203
rect 29377 11169 29411 11203
rect 29929 11169 29963 11203
rect 31309 11169 31343 11203
rect 32229 11169 32263 11203
rect 32321 11169 32355 11203
rect 33057 11169 33091 11203
rect 33333 11169 33367 11203
rect 33517 11169 33551 11203
rect 34253 11169 34287 11203
rect 34805 11169 34839 11203
rect 35081 11169 35115 11203
rect 35725 11169 35759 11203
rect 36461 11169 36495 11203
rect 38117 11169 38151 11203
rect 38577 11169 38611 11203
rect 3341 11101 3375 11135
rect 5457 11101 5491 11135
rect 14013 11101 14047 11135
rect 16497 11101 16531 11135
rect 21833 11101 21867 11135
rect 23765 11101 23799 11135
rect 24685 11101 24719 11135
rect 25881 11101 25915 11135
rect 26893 11101 26927 11135
rect 34713 11101 34747 11135
rect 37841 11101 37875 11135
rect 10977 11033 11011 11067
rect 13369 11033 13403 11067
rect 15485 11033 15519 11067
rect 28181 11033 28215 11067
rect 32229 11033 32263 11067
rect 32413 11033 32447 11067
rect 4445 10965 4479 10999
rect 17601 10965 17635 10999
rect 2513 10761 2547 10795
rect 4353 10761 4387 10795
rect 7021 10761 7055 10795
rect 9045 10761 9079 10795
rect 29101 10761 29135 10795
rect 13277 10693 13311 10727
rect 21097 10693 21131 10727
rect 31401 10693 31435 10727
rect 2237 10625 2271 10659
rect 8033 10625 8067 10659
rect 11529 10625 11563 10659
rect 14013 10625 14047 10659
rect 17141 10625 17175 10659
rect 18889 10625 18923 10659
rect 21557 10625 21591 10659
rect 24685 10625 24719 10659
rect 29101 10625 29135 10659
rect 29285 10625 29319 10659
rect 36093 10625 36127 10659
rect 37749 10625 37783 10659
rect 38853 10625 38887 10659
rect 2329 10557 2363 10591
rect 3433 10557 3467 10591
rect 4261 10557 4295 10591
rect 6837 10557 6871 10591
rect 7665 10557 7699 10591
rect 8401 10557 8435 10591
rect 8861 10557 8895 10591
rect 9873 10557 9907 10591
rect 10057 10557 10091 10591
rect 11437 10557 11471 10591
rect 11713 10557 11747 10591
rect 12449 10557 12483 10591
rect 13001 10557 13035 10591
rect 13369 10557 13403 10591
rect 14473 10557 14507 10591
rect 14657 10557 14691 10591
rect 14841 10557 14875 10591
rect 15485 10557 15519 10591
rect 16497 10557 16531 10591
rect 16957 10557 16991 10591
rect 17325 10557 17359 10591
rect 18061 10557 18095 10591
rect 19533 10557 19567 10591
rect 19625 10557 19659 10591
rect 19901 10557 19935 10591
rect 20085 10557 20119 10591
rect 21649 10557 21683 10591
rect 22017 10557 22051 10591
rect 22109 10557 22143 10591
rect 22661 10557 22695 10591
rect 23673 10557 23707 10591
rect 24961 10557 24995 10591
rect 27077 10557 27111 10591
rect 27169 10557 27203 10591
rect 27537 10557 27571 10591
rect 27629 10557 27663 10591
rect 29469 10557 29503 10591
rect 30021 10557 30055 10591
rect 30205 10557 30239 10591
rect 31309 10557 31343 10591
rect 31677 10557 31711 10591
rect 32137 10557 32171 10591
rect 32873 10557 32907 10591
rect 33241 10557 33275 10591
rect 33517 10557 33551 10591
rect 34437 10557 34471 10591
rect 35173 10557 35207 10591
rect 36461 10557 36495 10591
rect 36737 10557 36771 10591
rect 37473 10557 37507 10591
rect 10333 10489 10367 10523
rect 23765 10489 23799 10523
rect 28181 10489 28215 10523
rect 37013 10489 37047 10523
rect 3249 10421 3283 10455
rect 15669 10421 15703 10455
rect 18245 10421 18279 10455
rect 22845 10421 22879 10455
rect 26249 10421 26283 10455
rect 30481 10421 30515 10455
rect 32781 10421 32815 10455
rect 34253 10421 34287 10455
rect 35357 10421 35391 10455
rect 5641 10217 5675 10251
rect 13369 10217 13403 10251
rect 24133 10217 24167 10251
rect 27629 10217 27663 10251
rect 30573 10217 30607 10251
rect 32229 10217 32263 10251
rect 34805 10217 34839 10251
rect 37105 10217 37139 10251
rect 37841 10217 37875 10251
rect 11069 10149 11103 10183
rect 12817 10149 12851 10183
rect 15301 10149 15335 10183
rect 1685 10081 1719 10115
rect 4077 10081 4111 10115
rect 6193 10081 6227 10115
rect 7573 10081 7607 10115
rect 8309 10081 8343 10115
rect 8867 10081 8901 10115
rect 10517 10081 10551 10115
rect 10793 10081 10827 10115
rect 12357 10081 12391 10115
rect 12541 10081 12575 10115
rect 13461 10081 13495 10115
rect 13921 10081 13955 10115
rect 15945 10081 15979 10115
rect 16313 10081 16347 10115
rect 17141 10081 17175 10115
rect 17417 10081 17451 10115
rect 17969 10081 18003 10115
rect 18981 10081 19015 10115
rect 19349 10081 19383 10115
rect 19901 10081 19935 10115
rect 21557 10081 21591 10115
rect 21925 10081 21959 10115
rect 25237 10081 25271 10115
rect 25697 10081 25731 10115
rect 26525 10081 26559 10115
rect 27537 10081 27571 10115
rect 28457 10081 28491 10115
rect 30573 10081 30607 10115
rect 31033 10081 31067 10115
rect 31309 10081 31343 10115
rect 32321 10081 32355 10115
rect 32689 10081 32723 10115
rect 33701 10081 33735 10115
rect 34805 10081 34839 10115
rect 34897 10081 34931 10115
rect 35633 10081 35667 10115
rect 35817 10081 35851 10115
rect 36093 10081 36127 10115
rect 36921 10081 36955 10115
rect 38025 10081 38059 10115
rect 38209 10081 38243 10115
rect 38945 10081 38979 10115
rect 1409 10013 1443 10047
rect 2789 10013 2823 10047
rect 4353 10013 4387 10047
rect 7941 10013 7975 10047
rect 10057 10013 10091 10047
rect 14289 10013 14323 10047
rect 15853 10013 15887 10047
rect 16405 10013 16439 10047
rect 16957 10013 16991 10047
rect 21465 10013 21499 10047
rect 22017 10013 22051 10047
rect 22753 10013 22787 10047
rect 23029 10013 23063 10047
rect 24961 10013 24995 10047
rect 28181 10013 28215 10047
rect 32965 10013 32999 10047
rect 21005 9945 21039 9979
rect 25697 9945 25731 9979
rect 26709 9945 26743 9979
rect 33885 9945 33919 9979
rect 35357 10013 35391 10047
rect 39037 9945 39071 9979
rect 6377 9877 6411 9911
rect 9045 9877 9079 9911
rect 16957 9877 16991 9911
rect 17141 9877 17175 9911
rect 18797 9877 18831 9911
rect 20085 9877 20119 9911
rect 29745 9877 29779 9911
rect 34805 9877 34839 9911
rect 19993 9673 20027 9707
rect 38301 9673 38335 9707
rect 10241 9605 10275 9639
rect 12817 9605 12851 9639
rect 13645 9605 13679 9639
rect 18521 9605 18555 9639
rect 25145 9605 25179 9639
rect 26065 9605 26099 9639
rect 30665 9605 30699 9639
rect 4261 9537 4295 9571
rect 9229 9537 9263 9571
rect 16589 9537 16623 9571
rect 17325 9537 17359 9571
rect 19257 9537 19291 9571
rect 21189 9537 21223 9571
rect 21741 9537 21775 9571
rect 26893 9537 26927 9571
rect 29561 9537 29595 9571
rect 35817 9537 35851 9571
rect 36921 9537 36955 9571
rect 2329 9469 2363 9503
rect 2789 9469 2823 9503
rect 3617 9469 3651 9503
rect 3893 9469 3927 9503
rect 4353 9469 4387 9503
rect 4813 9469 4847 9503
rect 5365 9469 5399 9503
rect 5825 9469 5859 9503
rect 7021 9469 7055 9503
rect 7297 9469 7331 9503
rect 8677 9469 8711 9503
rect 9137 9469 9171 9503
rect 9965 9469 9999 9503
rect 10701 9469 10735 9503
rect 10793 9469 10827 9503
rect 11529 9469 11563 9503
rect 12633 9469 12667 9503
rect 13553 9469 13587 9503
rect 14105 9469 14139 9503
rect 14381 9469 14415 9503
rect 15393 9469 15427 9503
rect 15577 9469 15611 9503
rect 15761 9469 15795 9503
rect 16773 9469 16807 9503
rect 17233 9469 17267 9503
rect 18429 9469 18463 9503
rect 18797 9469 18831 9503
rect 19809 9469 19843 9503
rect 21281 9469 21315 9503
rect 21649 9469 21683 9503
rect 22293 9469 22327 9503
rect 22845 9469 22879 9503
rect 24041 9469 24075 9503
rect 24225 9469 24259 9503
rect 24685 9469 24719 9503
rect 24777 9469 24811 9503
rect 25881 9469 25915 9503
rect 27077 9469 27111 9503
rect 27537 9469 27571 9503
rect 27629 9469 27663 9503
rect 29101 9469 29135 9503
rect 29285 9469 29319 9503
rect 31401 9469 31435 9503
rect 32045 9469 32079 9503
rect 32229 9469 32263 9503
rect 33425 9469 33459 9503
rect 33977 9469 34011 9503
rect 34069 9469 34103 9503
rect 35357 9469 35391 9503
rect 35725 9469 35759 9503
rect 37197 9469 37231 9503
rect 14933 9401 14967 9435
rect 20637 9401 20671 9435
rect 28181 9401 28215 9435
rect 34897 9401 34931 9435
rect 2329 9333 2363 9367
rect 5917 9333 5951 9367
rect 11713 9333 11747 9367
rect 22385 9333 22419 9367
rect 28917 9333 28951 9367
rect 31493 9333 31527 9367
rect 33333 9333 33367 9367
rect 2973 9129 3007 9163
rect 13461 9129 13495 9163
rect 18337 9129 18371 9163
rect 27445 9129 27479 9163
rect 30205 9129 30239 9163
rect 36369 9129 36403 9163
rect 37841 9129 37875 9163
rect 19165 9061 19199 9095
rect 24133 9061 24167 9095
rect 26617 9061 26651 9095
rect 1685 8993 1719 9027
rect 3893 8993 3927 9027
rect 4445 8993 4479 9027
rect 4905 8993 4939 9027
rect 5457 8993 5491 9027
rect 5825 8993 5859 9027
rect 6101 8993 6135 9027
rect 7205 8993 7239 9027
rect 7757 8993 7791 9027
rect 8125 8993 8159 9027
rect 8585 8993 8619 9027
rect 9045 8993 9079 9027
rect 10701 8993 10735 9027
rect 11069 8993 11103 9027
rect 11713 8993 11747 9027
rect 12357 8993 12391 9027
rect 12725 8993 12759 9027
rect 13369 8993 13403 9027
rect 13921 8993 13955 9027
rect 15945 8993 15979 9027
rect 16313 8993 16347 9027
rect 17233 8993 17267 9027
rect 19809 8993 19843 9027
rect 19901 8993 19935 9027
rect 20177 8993 20211 9027
rect 21833 8993 21867 9027
rect 22201 8993 22235 9027
rect 23213 8993 23247 9027
rect 23581 8993 23615 9027
rect 23857 8993 23891 9027
rect 24777 8993 24811 9027
rect 25237 8993 25271 9027
rect 25329 8993 25363 9027
rect 26525 8993 26559 9027
rect 27353 8993 27387 9027
rect 28273 8993 28307 9027
rect 30113 8993 30147 9027
rect 30757 8993 30791 9027
rect 32137 8993 32171 9027
rect 33149 8993 33183 9027
rect 35265 8993 35299 9027
rect 37749 8993 37783 9027
rect 38485 8993 38519 9027
rect 38577 8993 38611 9027
rect 1409 8925 1443 8959
rect 4813 8925 4847 8959
rect 7297 8925 7331 8959
rect 11161 8925 11195 8959
rect 12265 8925 12299 8959
rect 12817 8925 12851 8959
rect 14381 8925 14415 8959
rect 15853 8925 15887 8959
rect 16405 8925 16439 8959
rect 16957 8925 16991 8959
rect 20269 8925 20303 8959
rect 21373 8925 21407 8959
rect 24685 8925 24719 8959
rect 27997 8925 28031 8959
rect 32873 8925 32907 8959
rect 34989 8925 35023 8959
rect 10517 8857 10551 8891
rect 22109 8857 22143 8891
rect 25697 8857 25731 8891
rect 30941 8857 30975 8891
rect 3709 8789 3743 8823
rect 15393 8789 15427 8823
rect 29377 8789 29411 8823
rect 32321 8789 32355 8823
rect 34437 8789 34471 8823
rect 4077 8585 4111 8619
rect 6193 8585 6227 8619
rect 11805 8585 11839 8619
rect 24133 8585 24167 8619
rect 26249 8585 26283 8619
rect 30849 8585 30883 8619
rect 38485 8585 38519 8619
rect 11253 8517 11287 8551
rect 13093 8517 13127 8551
rect 31677 8517 31711 8551
rect 33241 8517 33275 8551
rect 2789 8449 2823 8483
rect 4905 8449 4939 8483
rect 7205 8449 7239 8483
rect 13553 8449 13587 8483
rect 14105 8449 14139 8483
rect 16037 8449 16071 8483
rect 16589 8449 16623 8483
rect 18429 8449 18463 8483
rect 20085 8449 20119 8483
rect 21465 8449 21499 8483
rect 22201 8449 22235 8483
rect 24685 8449 24719 8483
rect 24961 8449 24995 8483
rect 26801 8449 26835 8483
rect 28457 8449 28491 8483
rect 1409 8381 1443 8415
rect 1685 8381 1719 8415
rect 3985 8381 4019 8415
rect 4629 8381 4663 8415
rect 7113 8381 7147 8415
rect 7757 8381 7791 8415
rect 8125 8381 8159 8415
rect 8309 8381 8343 8415
rect 9045 8381 9079 8415
rect 10057 8381 10091 8415
rect 10609 8381 10643 8415
rect 11437 8381 11471 8415
rect 11713 8381 11747 8415
rect 13645 8381 13679 8415
rect 14013 8381 14047 8415
rect 16129 8381 16163 8415
rect 16497 8381 16531 8415
rect 17325 8381 17359 8415
rect 17417 8381 17451 8415
rect 18061 8381 18095 8415
rect 18613 8381 18647 8415
rect 19533 8381 19567 8415
rect 19993 8381 20027 8415
rect 21005 8381 21039 8415
rect 21281 8381 21315 8415
rect 21925 8381 21959 8415
rect 22477 8381 22511 8415
rect 22661 8381 22695 8415
rect 23949 8381 23983 8415
rect 27077 8381 27111 8415
rect 29285 8381 29319 8415
rect 29561 8381 29595 8415
rect 31401 8381 31435 8415
rect 32045 8381 32079 8415
rect 32229 8381 32263 8415
rect 33425 8381 33459 8415
rect 33793 8381 33827 8415
rect 33885 8381 33919 8415
rect 34897 8381 34931 8415
rect 36553 8381 36587 8415
rect 37289 8381 37323 8415
rect 38393 8381 38427 8415
rect 15485 8313 15519 8347
rect 10333 8245 10367 8279
rect 35081 8245 35115 8279
rect 8677 8041 8711 8075
rect 16681 8041 16715 8075
rect 22477 8041 22511 8075
rect 25145 8041 25179 8075
rect 25881 8041 25915 8075
rect 27721 8041 27755 8075
rect 29377 8041 29411 8075
rect 31309 8041 31343 8075
rect 35817 8041 35851 8075
rect 14473 7973 14507 8007
rect 16037 7973 16071 8007
rect 28457 7973 28491 8007
rect 33793 7973 33827 8007
rect 4077 7905 4111 7939
rect 4537 7905 4571 7939
rect 4813 7905 4847 7939
rect 5457 7905 5491 7939
rect 6009 7905 6043 7939
rect 6469 7905 6503 7939
rect 6745 7905 6779 7939
rect 8125 7905 8159 7939
rect 8585 7905 8619 7939
rect 9689 7905 9723 7939
rect 11989 7905 12023 7939
rect 12449 7905 12483 7939
rect 13737 7905 13771 7939
rect 14197 7905 14231 7939
rect 15485 7905 15519 7939
rect 15761 7905 15795 7939
rect 16865 7905 16899 7939
rect 16957 7905 16991 7939
rect 17325 7905 17359 7939
rect 17693 7905 17727 7939
rect 18797 7905 18831 7939
rect 19625 7905 19659 7939
rect 19993 7905 20027 7939
rect 21373 7905 21407 7939
rect 23305 7905 23339 7939
rect 23949 7905 23983 7939
rect 24317 7905 24351 7939
rect 24961 7905 24995 7939
rect 25697 7905 25731 7939
rect 26709 7905 26743 7939
rect 27169 7905 27203 7939
rect 27261 7905 27295 7939
rect 28365 7905 28399 7939
rect 29285 7905 29319 7939
rect 32137 7905 32171 7939
rect 35081 7905 35115 7939
rect 35725 7905 35759 7939
rect 1409 7837 1443 7871
rect 1685 7837 1719 7871
rect 9965 7837 9999 7871
rect 12633 7837 12667 7871
rect 13553 7837 13587 7871
rect 19165 7837 19199 7871
rect 21097 7837 21131 7871
rect 26617 7837 26651 7871
rect 29929 7837 29963 7871
rect 30205 7837 30239 7871
rect 32413 7837 32447 7871
rect 34253 7837 34287 7871
rect 34805 7837 34839 7871
rect 35265 7837 35299 7871
rect 4169 7769 4203 7803
rect 11897 7769 11931 7803
rect 19901 7769 19935 7803
rect 23397 7769 23431 7803
rect 2973 7701 3007 7735
rect 11253 7701 11287 7735
rect 17049 7701 17083 7735
rect 18613 7701 18647 7735
rect 7021 7497 7055 7531
rect 8585 7497 8619 7531
rect 12817 7497 12851 7531
rect 15485 7497 15519 7531
rect 17141 7497 17175 7531
rect 28457 7497 28491 7531
rect 5549 7429 5583 7463
rect 7849 7429 7883 7463
rect 14197 7429 14231 7463
rect 22385 7429 22419 7463
rect 23765 7429 23799 7463
rect 3525 7361 3559 7395
rect 4905 7361 4939 7395
rect 9965 7361 9999 7395
rect 14933 7361 14967 7395
rect 18981 7361 19015 7395
rect 19257 7361 19291 7395
rect 25421 7361 25455 7395
rect 29285 7361 29319 7395
rect 30297 7361 30331 7395
rect 31585 7361 31619 7395
rect 35357 7361 35391 7395
rect 36737 7361 36771 7395
rect 37381 7361 37415 7395
rect 37657 7361 37691 7395
rect 2329 7293 2363 7327
rect 2513 7293 2547 7327
rect 3249 7293 3283 7327
rect 5365 7293 5399 7327
rect 6837 7293 6871 7327
rect 7757 7293 7791 7327
rect 8401 7293 8435 7327
rect 9137 7293 9171 7327
rect 9781 7293 9815 7327
rect 9873 7293 9907 7327
rect 10517 7293 10551 7327
rect 10793 7293 10827 7327
rect 11529 7293 11563 7327
rect 13001 7293 13035 7327
rect 14013 7293 14047 7327
rect 14473 7293 14507 7327
rect 15669 7293 15703 7327
rect 15761 7293 15795 7327
rect 16037 7293 16071 7327
rect 18245 7293 18279 7327
rect 21281 7293 21315 7327
rect 21557 7293 21591 7327
rect 21925 7293 21959 7327
rect 22477 7293 22511 7327
rect 23857 7293 23891 7327
rect 24041 7293 24075 7327
rect 24409 7293 24443 7327
rect 25329 7293 25363 7327
rect 25789 7293 25823 7327
rect 26341 7293 26375 7327
rect 27537 7293 27571 7327
rect 28273 7293 28307 7327
rect 29837 7293 29871 7327
rect 30113 7293 30147 7327
rect 31861 7293 31895 7327
rect 32045 7293 32079 7327
rect 33057 7293 33091 7327
rect 33333 7293 33367 7327
rect 33517 7293 33551 7327
rect 35081 7293 35115 7327
rect 11621 7225 11655 7259
rect 31033 7225 31067 7259
rect 32505 7225 32539 7259
rect 2145 7157 2179 7191
rect 18429 7157 18463 7191
rect 20361 7157 20395 7191
rect 21097 7157 21131 7191
rect 27721 7157 27755 7191
rect 38761 7157 38795 7191
rect 8677 6953 8711 6987
rect 22569 6953 22603 6987
rect 16865 6885 16899 6919
rect 18429 6885 18463 6919
rect 29009 6885 29043 6919
rect 2329 6817 2363 6851
rect 4261 6817 4295 6851
rect 4905 6817 4939 6851
rect 5549 6817 5583 6851
rect 5641 6817 5675 6851
rect 6285 6817 6319 6851
rect 6561 6817 6595 6851
rect 10609 6817 10643 6851
rect 11069 6817 11103 6851
rect 11805 6817 11839 6851
rect 13461 6817 13495 6851
rect 13921 6817 13955 6851
rect 14565 6817 14599 6851
rect 16313 6817 16347 6851
rect 16681 6817 16715 6851
rect 17601 6817 17635 6851
rect 17693 6817 17727 6851
rect 18061 6817 18095 6851
rect 19165 6817 19199 6851
rect 19533 6817 19567 6851
rect 20085 6817 20119 6851
rect 20913 6817 20947 6851
rect 21557 6817 21591 6851
rect 21925 6817 21959 6851
rect 22753 6817 22787 6851
rect 23121 6817 23155 6851
rect 23489 6817 23523 6851
rect 23857 6817 23891 6851
rect 24777 6817 24811 6851
rect 25145 6817 25179 6851
rect 25513 6817 25547 6851
rect 26525 6817 26559 6851
rect 28365 6817 28399 6851
rect 29837 6817 29871 6851
rect 30573 6817 30607 6851
rect 31125 6817 31159 6851
rect 31401 6817 31435 6851
rect 32137 6817 32171 6851
rect 33701 6817 33735 6851
rect 35817 6817 35851 6851
rect 2237 6749 2271 6783
rect 7297 6749 7331 6783
rect 7573 6749 7607 6783
rect 10425 6749 10459 6783
rect 11161 6749 11195 6783
rect 12081 6749 12115 6783
rect 15945 6749 15979 6783
rect 19993 6749 20027 6783
rect 21465 6749 21499 6783
rect 24961 6749 24995 6783
rect 27537 6749 27571 6783
rect 28089 6749 28123 6783
rect 28549 6749 28583 6783
rect 29561 6749 29595 6783
rect 30021 6749 30055 6783
rect 31585 6749 31619 6783
rect 33425 6749 33459 6783
rect 35541 6749 35575 6783
rect 4997 6681 5031 6715
rect 14657 6681 14691 6715
rect 22937 6681 22971 6715
rect 2513 6613 2547 6647
rect 4353 6613 4387 6647
rect 14013 6613 14047 6647
rect 26709 6613 26743 6647
rect 32321 6613 32355 6647
rect 34805 6613 34839 6647
rect 36921 6613 36955 6647
rect 9873 6409 9907 6443
rect 20913 6409 20947 6443
rect 26065 6409 26099 6443
rect 28181 6409 28215 6443
rect 29469 6409 29503 6443
rect 10609 6341 10643 6375
rect 12725 6341 12759 6375
rect 23765 6341 23799 6375
rect 4353 6273 4387 6307
rect 7481 6273 7515 6307
rect 15761 6273 15795 6307
rect 22477 6273 22511 6307
rect 31033 6273 31067 6307
rect 31493 6273 31527 6307
rect 32229 6273 32263 6307
rect 32781 6273 32815 6307
rect 36277 6273 36311 6307
rect 3893 6205 3927 6239
rect 4261 6205 4295 6239
rect 4721 6205 4755 6239
rect 5089 6205 5123 6239
rect 5641 6205 5675 6239
rect 6101 6205 6135 6239
rect 7113 6205 7147 6239
rect 7757 6205 7791 6239
rect 8125 6205 8159 6239
rect 8309 6205 8343 6239
rect 9045 6205 9079 6239
rect 9689 6205 9723 6239
rect 10425 6205 10459 6239
rect 11161 6205 11195 6239
rect 11253 6205 11287 6239
rect 12817 6205 12851 6239
rect 13277 6205 13311 6239
rect 13369 6205 13403 6239
rect 14013 6205 14047 6239
rect 14289 6205 14323 6239
rect 15301 6205 15335 6239
rect 15577 6205 15611 6239
rect 16589 6205 16623 6239
rect 16773 6205 16807 6239
rect 17325 6205 17359 6239
rect 18613 6205 18647 6239
rect 19257 6205 19291 6239
rect 19533 6205 19567 6239
rect 19809 6205 19843 6239
rect 21833 6205 21867 6239
rect 22201 6205 22235 6239
rect 22569 6205 22603 6239
rect 23949 6205 23983 6239
rect 24041 6205 24075 6239
rect 24685 6205 24719 6239
rect 25881 6205 25915 6239
rect 26617 6205 26651 6239
rect 26893 6205 26927 6239
rect 29285 6205 29319 6239
rect 31309 6205 31343 6239
rect 33057 6205 33091 6239
rect 33241 6205 33275 6239
rect 33701 6205 33735 6239
rect 34897 6205 34931 6239
rect 35173 6205 35207 6239
rect 37013 6205 37047 6239
rect 37565 6205 37599 6239
rect 37841 6205 37875 6239
rect 38025 6205 38059 6239
rect 6193 6137 6227 6171
rect 11713 6137 11747 6171
rect 17509 6137 17543 6171
rect 30481 6137 30515 6171
rect 33793 6137 33827 6171
rect 18429 6069 18463 6103
rect 19073 6069 19107 6103
rect 12817 5865 12851 5899
rect 14289 5865 14323 5899
rect 19073 5865 19107 5899
rect 21005 5865 21039 5899
rect 23213 5865 23247 5899
rect 28733 5865 28767 5899
rect 31493 5865 31527 5899
rect 6745 5797 6779 5831
rect 27077 5797 27111 5831
rect 35173 5797 35207 5831
rect 4353 5729 4387 5763
rect 6285 5729 6319 5763
rect 7205 5729 7239 5763
rect 7849 5729 7883 5763
rect 8125 5729 8159 5763
rect 8585 5729 8619 5763
rect 9137 5729 9171 5763
rect 9689 5729 9723 5763
rect 10333 5729 10367 5763
rect 10977 5729 11011 5763
rect 11345 5729 11379 5763
rect 11529 5729 11563 5763
rect 12265 5729 12299 5763
rect 12909 5729 12943 5763
rect 13369 5729 13403 5763
rect 13553 5729 13587 5763
rect 14473 5729 14507 5763
rect 15117 5729 15151 5763
rect 15301 5729 15335 5763
rect 15945 5729 15979 5763
rect 16037 5729 16071 5763
rect 16497 5729 16531 5763
rect 17233 5729 17267 5763
rect 17969 5729 18003 5763
rect 20913 5729 20947 5763
rect 21741 5729 21775 5763
rect 22109 5729 22143 5763
rect 23949 5729 23983 5763
rect 24961 5729 24995 5763
rect 25145 5729 25179 5763
rect 25789 5729 25823 5763
rect 27629 5729 27663 5763
rect 27905 5729 27939 5763
rect 28549 5729 28583 5763
rect 29929 5729 29963 5763
rect 30205 5729 30239 5763
rect 30389 5729 30423 5763
rect 31309 5729 31343 5763
rect 32689 5729 32723 5763
rect 32965 5729 32999 5763
rect 34529 5729 34563 5763
rect 34713 5729 34747 5763
rect 35725 5729 35759 5763
rect 36001 5729 36035 5763
rect 4077 5661 4111 5695
rect 6193 5661 6227 5695
rect 10517 5661 10551 5695
rect 17693 5661 17727 5695
rect 21833 5661 21867 5695
rect 28089 5661 28123 5695
rect 29377 5661 29411 5695
rect 32137 5661 32171 5695
rect 33149 5661 33183 5695
rect 33701 5661 33735 5695
rect 34253 5661 34287 5695
rect 36185 5661 36219 5695
rect 5641 5593 5675 5627
rect 7297 5593 7331 5627
rect 15393 5593 15427 5627
rect 24869 5593 24903 5627
rect 9781 5525 9815 5559
rect 14933 5525 14967 5559
rect 21557 5525 21591 5559
rect 24041 5525 24075 5559
rect 6009 5321 6043 5355
rect 8585 5321 8619 5355
rect 11621 5321 11655 5355
rect 18153 5321 18187 5355
rect 26433 5321 26467 5355
rect 33149 5321 33183 5355
rect 36645 5321 36679 5355
rect 4629 5185 4663 5219
rect 4905 5185 4939 5219
rect 7297 5185 7331 5219
rect 9229 5185 9263 5219
rect 12725 5185 12759 5219
rect 16221 5185 16255 5219
rect 19441 5185 19475 5219
rect 20177 5185 20211 5219
rect 22017 5185 22051 5219
rect 28181 5185 28215 5219
rect 28641 5185 28675 5219
rect 31585 5185 31619 5219
rect 35081 5185 35115 5219
rect 3341 5117 3375 5151
rect 3893 5117 3927 5151
rect 7021 5117 7055 5151
rect 9137 5117 9171 5151
rect 9689 5117 9723 5151
rect 10149 5117 10183 5151
rect 10333 5117 10367 5151
rect 11069 5117 11103 5151
rect 11529 5117 11563 5151
rect 12817 5117 12851 5151
rect 13277 5117 13311 5151
rect 13645 5117 13679 5151
rect 14013 5117 14047 5151
rect 14565 5117 14599 5151
rect 15301 5117 15335 5151
rect 15761 5117 15795 5151
rect 16037 5117 16071 5151
rect 16681 5117 16715 5151
rect 16957 5117 16991 5151
rect 17877 5117 17911 5151
rect 18061 5117 18095 5151
rect 18705 5117 18739 5151
rect 19165 5117 19199 5151
rect 19901 5117 19935 5151
rect 22109 5117 22143 5151
rect 24041 5117 24075 5151
rect 24869 5117 24903 5151
rect 25145 5117 25179 5151
rect 28457 5117 28491 5151
rect 29285 5117 29319 5151
rect 29561 5117 29595 5151
rect 31861 5117 31895 5151
rect 33977 5117 34011 5151
rect 35633 5117 35667 5151
rect 35909 5117 35943 5151
rect 36093 5117 36127 5151
rect 36553 5117 36587 5151
rect 4077 5049 4111 5083
rect 21557 5049 21591 5083
rect 22569 5049 22603 5083
rect 27629 5049 27663 5083
rect 17693 4981 17727 5015
rect 24225 4981 24259 5015
rect 30665 4981 30699 5015
rect 34161 4981 34195 5015
rect 5273 4777 5307 4811
rect 7205 4777 7239 4811
rect 8125 4777 8159 4811
rect 11621 4777 11655 4811
rect 20177 4777 20211 4811
rect 24317 4777 24351 4811
rect 25421 4777 25455 4811
rect 36645 4777 36679 4811
rect 29193 4709 29227 4743
rect 32137 4709 32171 4743
rect 5089 4641 5123 4675
rect 8309 4641 8343 4675
rect 8677 4641 8711 4675
rect 8953 4641 8987 4675
rect 10517 4641 10551 4675
rect 12633 4641 12667 4675
rect 14013 4641 14047 4675
rect 14473 4641 14507 4675
rect 15577 4641 15611 4675
rect 16037 4641 16071 4675
rect 16313 4641 16347 4675
rect 16865 4641 16899 4675
rect 17233 4641 17267 4675
rect 18245 4641 18279 4675
rect 19625 4641 19659 4675
rect 20085 4641 20119 4675
rect 21281 4641 21315 4675
rect 21741 4641 21775 4675
rect 22937 4641 22971 4675
rect 25329 4641 25363 4675
rect 27629 4641 27663 4675
rect 27905 4641 27939 4675
rect 29745 4641 29779 4675
rect 30021 4641 30055 4675
rect 32689 4641 32723 4675
rect 32965 4641 32999 4675
rect 34299 4641 34333 4675
rect 34437 4641 34471 4675
rect 5825 4573 5859 4607
rect 6101 4573 6135 4607
rect 9137 4573 9171 4607
rect 10241 4573 10275 4607
rect 12357 4573 12391 4607
rect 16497 4573 16531 4607
rect 17969 4573 18003 4607
rect 21097 4573 21131 4607
rect 23213 4573 23247 4607
rect 27077 4573 27111 4607
rect 28089 4573 28123 4607
rect 30205 4573 30239 4607
rect 32827 4573 32861 4607
rect 33609 4573 33643 4607
rect 34161 4573 34195 4607
rect 35081 4573 35115 4607
rect 35357 4573 35391 4607
rect 14565 4505 14599 4539
rect 21741 4505 21775 4539
rect 29469 4165 29503 4199
rect 3709 4097 3743 4131
rect 3985 4097 4019 4131
rect 8776 4097 8810 4131
rect 9039 4097 9073 4131
rect 14749 4097 14783 4131
rect 16129 4097 16163 4131
rect 17509 4097 17543 4131
rect 20269 4097 20303 4131
rect 21649 4097 21683 4131
rect 22661 4097 22695 4131
rect 30941 4097 30975 4131
rect 34897 4097 34931 4131
rect 35587 4097 35621 4131
rect 6009 4029 6043 4063
rect 7113 4029 7147 4063
rect 7389 4029 7423 4063
rect 8033 4029 8067 4063
rect 10425 4029 10459 4063
rect 11345 4029 11379 4063
rect 11529 4029 11563 4063
rect 13277 4029 13311 4063
rect 13461 4029 13495 4063
rect 14473 4029 14507 4063
rect 16773 4029 16807 4063
rect 17233 4029 17267 4063
rect 18613 4029 18647 4063
rect 19073 4029 19107 4063
rect 19993 4029 20027 4063
rect 22109 4029 22143 4063
rect 22201 4029 22235 4063
rect 25605 4029 25639 4063
rect 25881 4029 25915 4063
rect 26065 4029 26099 4063
rect 26525 4029 26559 4063
rect 26801 4029 26835 4063
rect 29285 4029 29319 4063
rect 31217 4029 31251 4063
rect 31401 4029 31435 4063
rect 32413 4029 32447 4063
rect 32689 4029 32723 4063
rect 32873 4029 32907 4063
rect 33885 4029 33919 4063
rect 34023 4029 34057 4063
rect 34161 4029 34195 4063
rect 35449 4029 35483 4063
rect 35725 4029 35759 4063
rect 11805 3961 11839 3995
rect 13737 3961 13771 3995
rect 19349 3961 19383 3995
rect 25053 3961 25087 3995
rect 30389 3961 30423 3995
rect 31861 3961 31895 3995
rect 33333 3961 33367 3995
rect 5273 3893 5307 3927
rect 6193 3893 6227 3927
rect 6929 3893 6963 3927
rect 8217 3893 8251 3927
rect 27905 3893 27939 3927
rect 7205 3689 7239 3723
rect 9781 3689 9815 3723
rect 30481 3689 30515 3723
rect 34989 3689 35023 3723
rect 10977 3621 11011 3655
rect 24961 3621 24995 3655
rect 27445 3621 27479 3655
rect 32137 3621 32171 3655
rect 5273 3553 5307 3587
rect 6377 3553 6411 3587
rect 7113 3553 7147 3587
rect 7849 3553 7883 3587
rect 8677 3553 8711 3587
rect 9965 3553 9999 3587
rect 10149 3553 10183 3587
rect 10885 3553 10919 3587
rect 11897 3553 11931 3587
rect 13737 3553 13771 3587
rect 14197 3553 14231 3587
rect 15945 3553 15979 3587
rect 16221 3553 16255 3587
rect 18061 3553 18095 3587
rect 21373 3553 21407 3587
rect 22569 3553 22603 3587
rect 22845 3553 22879 3587
rect 25513 3553 25547 3587
rect 25789 3553 25823 3587
rect 27997 3553 28031 3587
rect 28273 3553 28307 3587
rect 28457 3553 28491 3587
rect 29193 3553 29227 3587
rect 32965 3553 32999 3587
rect 33885 3553 33919 3587
rect 35725 3553 35759 3587
rect 5181 3485 5215 3519
rect 5733 3485 5767 3519
rect 7941 3485 7975 3519
rect 11621 3485 11655 3519
rect 14289 3485 14323 3519
rect 18337 3485 18371 3519
rect 21281 3485 21315 3519
rect 21833 3485 21867 3519
rect 25973 3485 26007 3519
rect 28917 3485 28951 3519
rect 32689 3485 32723 3519
rect 33149 3485 33183 3519
rect 33609 3485 33643 3519
rect 8861 3417 8895 3451
rect 6561 3349 6595 3383
rect 13185 3349 13219 3383
rect 17509 3349 17543 3383
rect 19625 3349 19659 3383
rect 24133 3349 24167 3383
rect 35909 3349 35943 3383
rect 10885 3145 10919 3179
rect 12725 3145 12759 3179
rect 28457 3145 28491 3179
rect 31401 3145 31435 3179
rect 33701 3145 33735 3179
rect 1869 3009 1903 3043
rect 6285 3009 6319 3043
rect 7481 3009 7515 3043
rect 9597 3009 9631 3043
rect 13553 3009 13587 3043
rect 13829 3009 13863 3043
rect 15669 3009 15703 3043
rect 16221 3009 16255 3043
rect 19809 3009 19843 3043
rect 21189 3009 21223 3043
rect 32413 3009 32447 3043
rect 34897 3009 34931 3043
rect 35449 3009 35483 3043
rect 35909 3009 35943 3043
rect 2145 2941 2179 2975
rect 5825 2941 5859 2975
rect 6101 2941 6135 2975
rect 7205 2941 7239 2975
rect 9321 2941 9355 2975
rect 12449 2941 12483 2975
rect 12541 2941 12575 2975
rect 15761 2941 15795 2975
rect 16681 2941 16715 2975
rect 16773 2941 16807 2975
rect 18153 2941 18187 2975
rect 18613 2941 18647 2975
rect 19533 2941 19567 2975
rect 21649 2941 21683 2975
rect 21741 2941 21775 2975
rect 23673 2941 23707 2975
rect 23765 2941 23799 2975
rect 24961 2941 24995 2975
rect 25237 2941 25271 2975
rect 27077 2941 27111 2975
rect 27353 2941 27387 2975
rect 30021 2941 30055 2975
rect 30297 2941 30331 2975
rect 32137 2941 32171 2975
rect 35725 2941 35759 2975
rect 17233 2873 17267 2907
rect 18889 2873 18923 2907
rect 22201 2873 22235 2907
rect 24225 2873 24259 2907
rect 3249 2805 3283 2839
rect 8769 2805 8803 2839
rect 15117 2805 15151 2839
rect 26525 2805 26559 2839
rect 9137 2601 9171 2635
rect 18429 2601 18463 2635
rect 28457 2601 28491 2635
rect 14933 2533 14967 2567
rect 20637 2533 20671 2567
rect 32597 2533 32631 2567
rect 4077 2465 4111 2499
rect 4353 2465 4387 2499
rect 6929 2465 6963 2499
rect 9045 2465 9079 2499
rect 10425 2465 10459 2499
rect 10701 2465 10735 2499
rect 13553 2465 13587 2499
rect 15853 2465 15887 2499
rect 18337 2465 18371 2499
rect 19257 2465 19291 2499
rect 22109 2465 22143 2499
rect 24041 2465 24075 2499
rect 24317 2465 24351 2499
rect 26893 2465 26927 2499
rect 29009 2465 29043 2499
rect 30297 2465 30331 2499
rect 30573 2465 30607 2499
rect 33425 2465 33459 2499
rect 7205 2397 7239 2431
rect 13277 2397 13311 2431
rect 15577 2397 15611 2431
rect 18981 2397 19015 2431
rect 21833 2397 21867 2431
rect 27169 2397 27203 2431
rect 29745 2397 29779 2431
rect 30757 2397 30791 2431
rect 33149 2397 33183 2431
rect 33609 2397 33643 2431
rect 8493 2329 8527 2363
rect 5457 2261 5491 2295
rect 11989 2261 12023 2295
rect 17141 2261 17175 2295
rect 23397 2261 23431 2295
rect 25605 2261 25639 2295
rect 38485 2261 38519 2295
<< metal1 >>
rect 1104 38650 39836 38672
rect 1104 38598 19606 38650
rect 19658 38598 19670 38650
rect 19722 38598 19734 38650
rect 19786 38598 19798 38650
rect 19850 38598 39836 38650
rect 1104 38576 39836 38598
rect 7558 38496 7564 38548
rect 7616 38536 7622 38548
rect 8297 38539 8355 38545
rect 8297 38536 8309 38539
rect 7616 38508 8309 38536
rect 7616 38496 7622 38508
rect 8297 38505 8309 38508
rect 8343 38505 8355 38539
rect 8297 38499 8355 38505
rect 19242 38496 19248 38548
rect 19300 38536 19306 38548
rect 29822 38536 29828 38548
rect 19300 38508 26188 38536
rect 29783 38508 29828 38536
rect 19300 38496 19306 38508
rect 9674 38468 9680 38480
rect 7852 38440 9680 38468
rect 1302 38360 1308 38412
rect 1360 38400 1366 38412
rect 7852 38400 7880 38440
rect 9674 38428 9680 38440
rect 9732 38428 9738 38480
rect 26160 38468 26188 38508
rect 29822 38496 29828 38508
rect 29880 38496 29886 38548
rect 26160 38440 30236 38468
rect 9030 38400 9036 38412
rect 1360 38372 7880 38400
rect 8991 38372 9036 38400
rect 1360 38360 1366 38372
rect 9030 38360 9036 38372
rect 9088 38360 9094 38412
rect 10689 38403 10747 38409
rect 10689 38369 10701 38403
rect 10735 38400 10747 38403
rect 10962 38400 10968 38412
rect 10735 38372 10968 38400
rect 10735 38369 10747 38372
rect 10689 38363 10747 38369
rect 10962 38360 10968 38372
rect 11020 38360 11026 38412
rect 11330 38400 11336 38412
rect 11291 38372 11336 38400
rect 11330 38360 11336 38372
rect 11388 38360 11394 38412
rect 11422 38360 11428 38412
rect 11480 38400 11486 38412
rect 12621 38403 12679 38409
rect 12621 38400 12633 38403
rect 11480 38372 12633 38400
rect 11480 38360 11486 38372
rect 12621 38369 12633 38372
rect 12667 38400 12679 38403
rect 13722 38400 13728 38412
rect 12667 38372 13728 38400
rect 12667 38369 12679 38372
rect 12621 38363 12679 38369
rect 13722 38360 13728 38372
rect 13780 38360 13786 38412
rect 30208 38409 30236 38440
rect 30009 38403 30067 38409
rect 30009 38369 30021 38403
rect 30055 38369 30067 38403
rect 30009 38363 30067 38369
rect 30193 38403 30251 38409
rect 30193 38369 30205 38403
rect 30239 38369 30251 38403
rect 30193 38363 30251 38369
rect 6086 38292 6092 38344
rect 6144 38332 6150 38344
rect 6917 38335 6975 38341
rect 6917 38332 6929 38335
rect 6144 38304 6929 38332
rect 6144 38292 6150 38304
rect 6917 38301 6929 38304
rect 6963 38301 6975 38335
rect 6917 38295 6975 38301
rect 7193 38335 7251 38341
rect 7193 38301 7205 38335
rect 7239 38332 7251 38335
rect 7926 38332 7932 38344
rect 7239 38304 7932 38332
rect 7239 38301 7251 38304
rect 7193 38295 7251 38301
rect 7926 38292 7932 38304
rect 7984 38292 7990 38344
rect 30024 38332 30052 38363
rect 30466 38332 30472 38344
rect 30024 38304 30472 38332
rect 30466 38292 30472 38304
rect 30524 38292 30530 38344
rect 25498 38224 25504 38276
rect 25556 38264 25562 38276
rect 30650 38264 30656 38276
rect 25556 38236 30656 38264
rect 25556 38224 25562 38236
rect 30650 38224 30656 38236
rect 30708 38224 30714 38276
rect 8110 38156 8116 38208
rect 8168 38196 8174 38208
rect 9125 38199 9183 38205
rect 9125 38196 9137 38199
rect 8168 38168 9137 38196
rect 8168 38156 8174 38168
rect 9125 38165 9137 38168
rect 9171 38165 9183 38199
rect 10778 38196 10784 38208
rect 10739 38168 10784 38196
rect 9125 38159 9183 38165
rect 10778 38156 10784 38168
rect 10836 38156 10842 38208
rect 11054 38156 11060 38208
rect 11112 38196 11118 38208
rect 11425 38199 11483 38205
rect 11425 38196 11437 38199
rect 11112 38168 11437 38196
rect 11112 38156 11118 38168
rect 11425 38165 11437 38168
rect 11471 38165 11483 38199
rect 12710 38196 12716 38208
rect 12671 38168 12716 38196
rect 11425 38159 11483 38165
rect 12710 38156 12716 38168
rect 12768 38156 12774 38208
rect 26786 38156 26792 38208
rect 26844 38196 26850 38208
rect 32950 38196 32956 38208
rect 26844 38168 32956 38196
rect 26844 38156 26850 38168
rect 32950 38156 32956 38168
rect 33008 38156 33014 38208
rect 1104 38106 39836 38128
rect 1104 38054 4246 38106
rect 4298 38054 4310 38106
rect 4362 38054 4374 38106
rect 4426 38054 4438 38106
rect 4490 38054 34966 38106
rect 35018 38054 35030 38106
rect 35082 38054 35094 38106
rect 35146 38054 35158 38106
rect 35210 38054 39836 38106
rect 1104 38032 39836 38054
rect 6181 37995 6239 38001
rect 6181 37961 6193 37995
rect 6227 37992 6239 37995
rect 9766 37992 9772 38004
rect 6227 37964 9772 37992
rect 6227 37961 6239 37964
rect 6181 37955 6239 37961
rect 9766 37952 9772 37964
rect 9824 37952 9830 38004
rect 13998 37992 14004 38004
rect 13959 37964 14004 37992
rect 13998 37952 14004 37964
rect 14056 37952 14062 38004
rect 20809 37995 20867 38001
rect 20809 37961 20821 37995
rect 20855 37992 20867 37995
rect 26786 37992 26792 38004
rect 20855 37964 26792 37992
rect 20855 37961 20867 37964
rect 20809 37955 20867 37961
rect 26786 37952 26792 37964
rect 26844 37952 26850 38004
rect 36449 37995 36507 38001
rect 36449 37961 36461 37995
rect 36495 37992 36507 37995
rect 37182 37992 37188 38004
rect 36495 37964 37188 37992
rect 36495 37961 36507 37964
rect 36449 37955 36507 37961
rect 37182 37952 37188 37964
rect 37240 37952 37246 38004
rect 29825 37927 29883 37933
rect 29825 37893 29837 37927
rect 29871 37893 29883 37927
rect 29825 37887 29883 37893
rect 3326 37816 3332 37868
rect 3384 37856 3390 37868
rect 8110 37856 8116 37868
rect 3384 37828 7972 37856
rect 8071 37828 8116 37856
rect 3384 37816 3390 37828
rect 4617 37791 4675 37797
rect 4617 37757 4629 37791
rect 4663 37757 4675 37791
rect 4617 37751 4675 37757
rect 4893 37791 4951 37797
rect 4893 37757 4905 37791
rect 4939 37788 4951 37791
rect 5166 37788 5172 37800
rect 4939 37760 5172 37788
rect 4939 37757 4951 37760
rect 4893 37751 4951 37757
rect 4632 37652 4660 37751
rect 5166 37748 5172 37760
rect 5224 37748 5230 37800
rect 6825 37791 6883 37797
rect 6825 37757 6837 37791
rect 6871 37788 6883 37791
rect 7466 37788 7472 37800
rect 6871 37760 7472 37788
rect 6871 37757 6883 37760
rect 6825 37751 6883 37757
rect 7466 37748 7472 37760
rect 7524 37748 7530 37800
rect 7742 37748 7748 37800
rect 7800 37788 7806 37800
rect 7837 37791 7895 37797
rect 7837 37788 7849 37791
rect 7800 37760 7849 37788
rect 7800 37748 7806 37760
rect 7837 37757 7849 37760
rect 7883 37757 7895 37791
rect 7944 37788 7972 37828
rect 8110 37816 8116 37828
rect 8168 37816 8174 37868
rect 8202 37816 8208 37868
rect 8260 37856 8266 37868
rect 10045 37859 10103 37865
rect 10045 37856 10057 37859
rect 8260 37828 10057 37856
rect 8260 37816 8266 37828
rect 10045 37825 10057 37828
rect 10091 37825 10103 37859
rect 10045 37819 10103 37825
rect 14553 37859 14611 37865
rect 14553 37825 14565 37859
rect 14599 37856 14611 37859
rect 15286 37856 15292 37868
rect 14599 37828 15292 37856
rect 14599 37825 14611 37828
rect 14553 37819 14611 37825
rect 15286 37816 15292 37828
rect 15344 37816 15350 37868
rect 17218 37816 17224 37868
rect 17276 37856 17282 37868
rect 25498 37856 25504 37868
rect 17276 37828 25504 37856
rect 17276 37816 17282 37828
rect 25498 37816 25504 37828
rect 25556 37816 25562 37868
rect 25593 37859 25651 37865
rect 25593 37825 25605 37859
rect 25639 37856 25651 37859
rect 26329 37859 26387 37865
rect 26329 37856 26341 37859
rect 25639 37828 26341 37856
rect 25639 37825 25651 37828
rect 25593 37819 25651 37825
rect 26329 37825 26341 37828
rect 26375 37825 26387 37859
rect 26329 37819 26387 37825
rect 26694 37816 26700 37868
rect 26752 37856 26758 37868
rect 29840 37856 29868 37887
rect 26752 37828 29868 37856
rect 26752 37816 26758 37828
rect 34606 37816 34612 37868
rect 34664 37856 34670 37868
rect 35161 37859 35219 37865
rect 35161 37856 35173 37859
rect 34664 37828 35173 37856
rect 34664 37816 34670 37828
rect 35161 37825 35173 37828
rect 35207 37825 35219 37859
rect 35161 37819 35219 37825
rect 9493 37791 9551 37797
rect 9493 37788 9505 37791
rect 7944 37760 9505 37788
rect 7837 37751 7895 37757
rect 9493 37757 9505 37760
rect 9539 37788 9551 37791
rect 9674 37788 9680 37800
rect 9539 37760 9680 37788
rect 9539 37757 9551 37760
rect 9493 37751 9551 37757
rect 9674 37748 9680 37760
rect 9732 37788 9738 37800
rect 9953 37791 10011 37797
rect 9953 37788 9965 37791
rect 9732 37760 9965 37788
rect 9732 37748 9738 37760
rect 9953 37757 9965 37760
rect 9999 37757 10011 37791
rect 9953 37751 10011 37757
rect 10597 37791 10655 37797
rect 10597 37757 10609 37791
rect 10643 37757 10655 37791
rect 10962 37788 10968 37800
rect 10923 37760 10968 37788
rect 10597 37751 10655 37757
rect 6086 37652 6092 37664
rect 4632 37624 6092 37652
rect 6086 37612 6092 37624
rect 6144 37612 6150 37664
rect 6914 37652 6920 37664
rect 6875 37624 6920 37652
rect 6914 37612 6920 37624
rect 6972 37612 6978 37664
rect 10612 37652 10640 37751
rect 10962 37748 10968 37760
rect 11020 37748 11026 37800
rect 11422 37788 11428 37800
rect 11383 37760 11428 37788
rect 11422 37748 11428 37760
rect 11480 37748 11486 37800
rect 12434 37748 12440 37800
rect 12492 37788 12498 37800
rect 12713 37791 12771 37797
rect 12492 37760 12537 37788
rect 12492 37748 12498 37760
rect 12713 37757 12725 37791
rect 12759 37788 12771 37791
rect 13538 37788 13544 37800
rect 12759 37760 13544 37788
rect 12759 37757 12771 37760
rect 12713 37751 12771 37757
rect 13538 37748 13544 37760
rect 13596 37748 13602 37800
rect 14829 37791 14887 37797
rect 14829 37757 14841 37791
rect 14875 37788 14887 37791
rect 15838 37788 15844 37800
rect 14875 37760 15844 37788
rect 14875 37757 14887 37760
rect 14829 37751 14887 37757
rect 15838 37748 15844 37760
rect 15896 37748 15902 37800
rect 17954 37748 17960 37800
rect 18012 37788 18018 37800
rect 19245 37791 19303 37797
rect 19245 37788 19257 37791
rect 18012 37760 19257 37788
rect 18012 37748 18018 37760
rect 19245 37757 19257 37760
rect 19291 37757 19303 37791
rect 19521 37791 19579 37797
rect 19521 37788 19533 37791
rect 19245 37751 19303 37757
rect 19352 37760 19533 37788
rect 13998 37652 14004 37664
rect 10612 37624 14004 37652
rect 13998 37612 14004 37624
rect 14056 37652 14062 37664
rect 15933 37655 15991 37661
rect 15933 37652 15945 37655
rect 14056 37624 15945 37652
rect 14056 37612 14062 37624
rect 15933 37621 15945 37624
rect 15979 37621 15991 37655
rect 15933 37615 15991 37621
rect 18782 37612 18788 37664
rect 18840 37652 18846 37664
rect 19061 37655 19119 37661
rect 19061 37652 19073 37655
rect 18840 37624 19073 37652
rect 18840 37612 18846 37624
rect 19061 37621 19073 37624
rect 19107 37652 19119 37655
rect 19352 37652 19380 37760
rect 19521 37757 19533 37760
rect 19567 37757 19579 37791
rect 21450 37788 21456 37800
rect 21411 37760 21456 37788
rect 19521 37751 19579 37757
rect 21450 37748 21456 37760
rect 21508 37748 21514 37800
rect 21729 37791 21787 37797
rect 21729 37757 21741 37791
rect 21775 37788 21787 37791
rect 21818 37788 21824 37800
rect 21775 37760 21824 37788
rect 21775 37757 21787 37760
rect 21729 37751 21787 37757
rect 21818 37748 21824 37760
rect 21876 37748 21882 37800
rect 23937 37791 23995 37797
rect 23937 37757 23949 37791
rect 23983 37757 23995 37791
rect 24210 37788 24216 37800
rect 24171 37760 24216 37788
rect 23937 37751 23995 37757
rect 23109 37723 23167 37729
rect 23109 37689 23121 37723
rect 23155 37720 23167 37723
rect 23290 37720 23296 37732
rect 23155 37692 23296 37720
rect 23155 37689 23167 37692
rect 23109 37683 23167 37689
rect 23290 37680 23296 37692
rect 23348 37680 23354 37732
rect 19107 37624 19380 37652
rect 19107 37621 19119 37624
rect 19061 37615 19119 37621
rect 21450 37612 21456 37664
rect 21508 37652 21514 37664
rect 23014 37652 23020 37664
rect 21508 37624 23020 37652
rect 21508 37612 21514 37624
rect 23014 37612 23020 37624
rect 23072 37652 23078 37664
rect 23952 37652 23980 37751
rect 24210 37748 24216 37760
rect 24268 37748 24274 37800
rect 26053 37791 26111 37797
rect 26053 37788 26065 37791
rect 25700 37760 26065 37788
rect 24578 37652 24584 37664
rect 23072 37624 24584 37652
rect 23072 37612 23078 37624
rect 24578 37612 24584 37624
rect 24636 37652 24642 37664
rect 25700 37652 25728 37760
rect 26053 37757 26065 37760
rect 26099 37788 26111 37791
rect 26418 37788 26424 37800
rect 26099 37760 26424 37788
rect 26099 37757 26111 37760
rect 26053 37751 26111 37757
rect 26418 37748 26424 37760
rect 26476 37748 26482 37800
rect 29822 37788 29828 37800
rect 29783 37760 29828 37788
rect 29822 37748 29828 37760
rect 29880 37748 29886 37800
rect 30466 37788 30472 37800
rect 30379 37760 30472 37788
rect 30466 37748 30472 37760
rect 30524 37748 30530 37800
rect 30745 37791 30803 37797
rect 30745 37757 30757 37791
rect 30791 37788 30803 37791
rect 31478 37788 31484 37800
rect 30791 37760 31484 37788
rect 30791 37757 30803 37760
rect 30745 37751 30803 37757
rect 31478 37748 31484 37760
rect 31536 37748 31542 37800
rect 33594 37748 33600 37800
rect 33652 37788 33658 37800
rect 34885 37791 34943 37797
rect 34885 37788 34897 37791
rect 33652 37760 34897 37788
rect 33652 37748 33658 37760
rect 34885 37757 34897 37760
rect 34931 37757 34943 37791
rect 34885 37751 34943 37757
rect 30484 37720 30512 37748
rect 31018 37720 31024 37732
rect 30484 37692 31024 37720
rect 31018 37680 31024 37692
rect 31076 37680 31082 37732
rect 24636 37624 25728 37652
rect 24636 37612 24642 37624
rect 26786 37612 26792 37664
rect 26844 37652 26850 37664
rect 27433 37655 27491 37661
rect 27433 37652 27445 37655
rect 26844 37624 27445 37652
rect 26844 37612 26850 37624
rect 27433 37621 27445 37624
rect 27479 37621 27491 37655
rect 27433 37615 27491 37621
rect 1104 37562 39836 37584
rect 1104 37510 19606 37562
rect 19658 37510 19670 37562
rect 19722 37510 19734 37562
rect 19786 37510 19798 37562
rect 19850 37510 39836 37562
rect 1104 37488 39836 37510
rect 1673 37451 1731 37457
rect 1673 37417 1685 37451
rect 1719 37448 1731 37451
rect 17218 37448 17224 37460
rect 1719 37420 17224 37448
rect 1719 37417 1731 37420
rect 1673 37411 1731 37417
rect 1780 37321 1808 37420
rect 17218 37408 17224 37420
rect 17276 37408 17282 37460
rect 17954 37448 17960 37460
rect 17328 37420 17960 37448
rect 5534 37380 5540 37392
rect 5000 37352 5540 37380
rect 1765 37315 1823 37321
rect 1765 37281 1777 37315
rect 1811 37281 1823 37315
rect 1765 37275 1823 37281
rect 1854 37272 1860 37324
rect 1912 37312 1918 37324
rect 5000 37321 5028 37352
rect 5534 37340 5540 37352
rect 5592 37340 5598 37392
rect 9030 37380 9036 37392
rect 8312 37352 8524 37380
rect 8991 37352 9036 37380
rect 4985 37315 5043 37321
rect 1912 37284 1992 37312
rect 1912 37272 1918 37284
rect 1964 37185 1992 37284
rect 4985 37281 4997 37315
rect 5031 37281 5043 37315
rect 4985 37275 5043 37281
rect 5077 37315 5135 37321
rect 5077 37281 5089 37315
rect 5123 37312 5135 37315
rect 5905 37315 5963 37321
rect 5905 37312 5917 37315
rect 5123 37284 5917 37312
rect 5123 37281 5135 37284
rect 5077 37275 5135 37281
rect 5905 37281 5917 37284
rect 5951 37281 5963 37315
rect 8202 37312 8208 37324
rect 8163 37284 8208 37312
rect 5905 37275 5963 37281
rect 8202 37272 8208 37284
rect 8260 37272 8266 37324
rect 8312 37321 8340 37352
rect 8297 37315 8355 37321
rect 8297 37281 8309 37315
rect 8343 37281 8355 37315
rect 8297 37275 8355 37281
rect 8496 37256 8524 37352
rect 9030 37340 9036 37352
rect 9088 37340 9094 37392
rect 13998 37380 14004 37392
rect 13372 37352 14004 37380
rect 8662 37312 8668 37324
rect 8623 37284 8668 37312
rect 8662 37272 8668 37284
rect 8720 37272 8726 37324
rect 9674 37312 9680 37324
rect 9635 37284 9680 37312
rect 9674 37272 9680 37284
rect 9732 37272 9738 37324
rect 11054 37312 11060 37324
rect 11015 37284 11060 37312
rect 11054 37272 11060 37284
rect 11112 37272 11118 37324
rect 13372 37321 13400 37352
rect 13998 37340 14004 37352
rect 14056 37340 14062 37392
rect 13357 37315 13415 37321
rect 13357 37281 13369 37315
rect 13403 37281 13415 37315
rect 13722 37312 13728 37324
rect 13683 37284 13728 37312
rect 13357 37275 13415 37281
rect 13722 37272 13728 37284
rect 13780 37272 13786 37324
rect 14090 37312 14096 37324
rect 14051 37284 14096 37312
rect 14090 37272 14096 37284
rect 14148 37272 14154 37324
rect 14366 37312 14372 37324
rect 14327 37284 14372 37312
rect 14366 37272 14372 37284
rect 14424 37272 14430 37324
rect 15289 37315 15347 37321
rect 15289 37312 15301 37315
rect 14476 37284 15301 37312
rect 5629 37247 5687 37253
rect 5629 37213 5641 37247
rect 5675 37244 5687 37247
rect 6086 37244 6092 37256
rect 5675 37216 6092 37244
rect 5675 37213 5687 37216
rect 5629 37207 5687 37213
rect 6086 37204 6092 37216
rect 6144 37204 6150 37256
rect 8478 37244 8484 37256
rect 8391 37216 8484 37244
rect 8478 37204 8484 37216
rect 8536 37244 8542 37256
rect 9214 37244 9220 37256
rect 8536 37216 9220 37244
rect 8536 37204 8542 37216
rect 9214 37204 9220 37216
rect 9272 37204 9278 37256
rect 9858 37204 9864 37256
rect 9916 37244 9922 37256
rect 10781 37247 10839 37253
rect 10781 37244 10793 37247
rect 9916 37216 10793 37244
rect 9916 37204 9922 37216
rect 10781 37213 10793 37216
rect 10827 37244 10839 37247
rect 12434 37244 12440 37256
rect 10827 37216 12440 37244
rect 10827 37213 10839 37216
rect 10781 37207 10839 37213
rect 12434 37204 12440 37216
rect 12492 37204 12498 37256
rect 13906 37204 13912 37256
rect 13964 37244 13970 37256
rect 14476 37244 14504 37284
rect 15289 37281 15301 37284
rect 15335 37281 15347 37315
rect 15289 37275 15347 37281
rect 15746 37272 15752 37324
rect 15804 37312 15810 37324
rect 15933 37315 15991 37321
rect 15933 37312 15945 37315
rect 15804 37284 15945 37312
rect 15804 37272 15810 37284
rect 15933 37281 15945 37284
rect 15979 37281 15991 37315
rect 15933 37275 15991 37281
rect 16022 37272 16028 37324
rect 16080 37312 16086 37324
rect 17221 37315 17279 37321
rect 17221 37312 17233 37315
rect 16080 37284 16125 37312
rect 16500 37284 17233 37312
rect 16080 37272 16086 37284
rect 13964 37216 14504 37244
rect 13964 37204 13970 37216
rect 15378 37204 15384 37256
rect 15436 37244 15442 37256
rect 16500 37244 16528 37284
rect 17221 37281 17233 37284
rect 17267 37312 17279 37315
rect 17328 37312 17356 37420
rect 17954 37408 17960 37420
rect 18012 37408 18018 37460
rect 21818 37408 21824 37460
rect 21876 37448 21882 37460
rect 22281 37451 22339 37457
rect 22281 37448 22293 37451
rect 21876 37420 22293 37448
rect 21876 37408 21882 37420
rect 22281 37417 22293 37420
rect 22327 37417 22339 37451
rect 22281 37411 22339 37417
rect 23124 37420 23980 37448
rect 17494 37312 17500 37324
rect 17267 37284 17356 37312
rect 17455 37284 17500 37312
rect 17267 37281 17279 37284
rect 17221 37275 17279 37281
rect 17494 37272 17500 37284
rect 17552 37272 17558 37324
rect 18877 37315 18935 37321
rect 18877 37281 18889 37315
rect 18923 37312 18935 37315
rect 23124 37312 23152 37420
rect 23952 37380 23980 37420
rect 24210 37408 24216 37460
rect 24268 37448 24274 37460
rect 24397 37451 24455 37457
rect 24397 37448 24409 37451
rect 24268 37420 24409 37448
rect 24268 37408 24274 37420
rect 24397 37417 24409 37420
rect 24443 37417 24455 37451
rect 25314 37448 25320 37460
rect 25275 37420 25320 37448
rect 24397 37411 24455 37417
rect 25314 37408 25320 37420
rect 25372 37408 25378 37460
rect 28718 37448 28724 37460
rect 25424 37420 28724 37448
rect 25424 37380 25452 37420
rect 28718 37408 28724 37420
rect 28776 37408 28782 37460
rect 23952 37352 25452 37380
rect 35253 37383 35311 37389
rect 35253 37349 35265 37383
rect 35299 37380 35311 37383
rect 39390 37380 39396 37392
rect 35299 37352 39396 37380
rect 35299 37349 35311 37352
rect 35253 37343 35311 37349
rect 39390 37340 39396 37352
rect 39448 37340 39454 37392
rect 23290 37312 23296 37324
rect 18923 37284 23152 37312
rect 23251 37284 23296 37312
rect 18923 37281 18935 37284
rect 18877 37275 18935 37281
rect 23290 37272 23296 37284
rect 23348 37272 23354 37324
rect 25498 37312 25504 37324
rect 25459 37284 25504 37312
rect 25498 37272 25504 37284
rect 25556 37272 25562 37324
rect 25777 37315 25835 37321
rect 25777 37281 25789 37315
rect 25823 37312 25835 37315
rect 26234 37312 26240 37324
rect 25823 37284 26240 37312
rect 25823 37281 25835 37284
rect 25777 37275 25835 37281
rect 26234 37272 26240 37284
rect 26292 37272 26298 37324
rect 26418 37272 26424 37324
rect 26476 37312 26482 37324
rect 26513 37315 26571 37321
rect 26513 37312 26525 37315
rect 26476 37284 26525 37312
rect 26476 37272 26482 37284
rect 26513 37281 26525 37284
rect 26559 37281 26571 37315
rect 26786 37312 26792 37324
rect 26747 37284 26792 37312
rect 26513 37275 26571 37281
rect 15436 37216 16528 37244
rect 15436 37204 15442 37216
rect 20162 37204 20168 37256
rect 20220 37244 20226 37256
rect 20901 37247 20959 37253
rect 20901 37244 20913 37247
rect 20220 37216 20913 37244
rect 20220 37204 20226 37216
rect 20901 37213 20913 37216
rect 20947 37213 20959 37247
rect 21174 37244 21180 37256
rect 21135 37216 21180 37244
rect 20901 37207 20959 37213
rect 21174 37204 21180 37216
rect 21232 37204 21238 37256
rect 23014 37244 23020 37256
rect 22975 37216 23020 37244
rect 23014 37204 23020 37216
rect 23072 37204 23078 37256
rect 26528 37244 26556 37275
rect 26786 37272 26792 37284
rect 26844 37272 26850 37324
rect 28629 37315 28687 37321
rect 28629 37281 28641 37315
rect 28675 37281 28687 37315
rect 28629 37275 28687 37281
rect 33505 37315 33563 37321
rect 33505 37281 33517 37315
rect 33551 37312 33563 37315
rect 33873 37315 33931 37321
rect 33873 37312 33885 37315
rect 33551 37284 33885 37312
rect 33551 37281 33563 37284
rect 33505 37275 33563 37281
rect 33873 37281 33885 37284
rect 33919 37312 33931 37315
rect 33962 37312 33968 37324
rect 33919 37284 33968 37312
rect 33919 37281 33931 37284
rect 33873 37275 33931 37281
rect 28644 37244 28672 37275
rect 33962 37272 33968 37284
rect 34020 37272 34026 37324
rect 28902 37244 28908 37256
rect 26528 37216 28672 37244
rect 28863 37216 28908 37244
rect 28902 37204 28908 37216
rect 28960 37204 28966 37256
rect 33594 37244 33600 37256
rect 33555 37216 33600 37244
rect 33594 37204 33600 37216
rect 33652 37204 33658 37256
rect 1949 37179 2007 37185
rect 1949 37145 1961 37179
rect 1995 37145 2007 37179
rect 1949 37139 2007 37145
rect 11882 37136 11888 37188
rect 11940 37176 11946 37188
rect 12345 37179 12403 37185
rect 12345 37176 12357 37179
rect 11940 37148 12357 37176
rect 11940 37136 11946 37148
rect 12345 37145 12357 37148
rect 12391 37176 12403 37179
rect 14366 37176 14372 37188
rect 12391 37148 14372 37176
rect 12391 37145 12403 37148
rect 12345 37139 12403 37145
rect 14366 37136 14372 37148
rect 14424 37136 14430 37188
rect 7190 37108 7196 37120
rect 7151 37080 7196 37108
rect 7190 37068 7196 37080
rect 7248 37068 7254 37120
rect 9674 37068 9680 37120
rect 9732 37108 9738 37120
rect 9769 37111 9827 37117
rect 9769 37108 9781 37111
rect 9732 37080 9781 37108
rect 9732 37068 9738 37080
rect 9769 37077 9781 37080
rect 9815 37077 9827 37111
rect 13170 37108 13176 37120
rect 13131 37080 13176 37108
rect 9769 37071 9827 37077
rect 13170 37068 13176 37080
rect 13228 37068 13234 37120
rect 13722 37068 13728 37120
rect 13780 37108 13786 37120
rect 15010 37108 15016 37120
rect 13780 37080 15016 37108
rect 13780 37068 13786 37080
rect 15010 37068 15016 37080
rect 15068 37068 15074 37120
rect 15194 37068 15200 37120
rect 15252 37108 15258 37120
rect 15381 37111 15439 37117
rect 15381 37108 15393 37111
rect 15252 37080 15393 37108
rect 15252 37068 15258 37080
rect 15381 37077 15393 37080
rect 15427 37077 15439 37111
rect 15381 37071 15439 37077
rect 27706 37068 27712 37120
rect 27764 37108 27770 37120
rect 27893 37111 27951 37117
rect 27893 37108 27905 37111
rect 27764 37080 27905 37108
rect 27764 37068 27770 37080
rect 27893 37077 27905 37080
rect 27939 37077 27951 37111
rect 30006 37108 30012 37120
rect 29967 37080 30012 37108
rect 27893 37071 27951 37077
rect 30006 37068 30012 37080
rect 30064 37068 30070 37120
rect 1104 37018 39836 37040
rect 1104 36966 4246 37018
rect 4298 36966 4310 37018
rect 4362 36966 4374 37018
rect 4426 36966 4438 37018
rect 4490 36966 34966 37018
rect 35018 36966 35030 37018
rect 35082 36966 35094 37018
rect 35146 36966 35158 37018
rect 35210 36966 39836 37018
rect 1104 36944 39836 36966
rect 8662 36904 8668 36916
rect 8623 36876 8668 36904
rect 8662 36864 8668 36876
rect 8720 36864 8726 36916
rect 14366 36904 14372 36916
rect 8956 36876 14372 36904
rect 5626 36796 5632 36848
rect 5684 36836 5690 36848
rect 8956 36836 8984 36876
rect 14366 36864 14372 36876
rect 14424 36864 14430 36916
rect 15838 36904 15844 36916
rect 15799 36876 15844 36904
rect 15838 36864 15844 36876
rect 15896 36864 15902 36916
rect 20346 36864 20352 36916
rect 20404 36904 20410 36916
rect 20404 36876 31616 36904
rect 20404 36864 20410 36876
rect 5684 36808 8984 36836
rect 5684 36796 5690 36808
rect 9214 36796 9220 36848
rect 9272 36836 9278 36848
rect 9272 36808 10180 36836
rect 9272 36796 9278 36808
rect 5534 36768 5540 36780
rect 5495 36740 5540 36768
rect 5534 36728 5540 36740
rect 5592 36728 5598 36780
rect 8478 36768 8484 36780
rect 5736 36740 8484 36768
rect 5736 36709 5764 36740
rect 8478 36728 8484 36740
rect 8536 36728 8542 36780
rect 9674 36768 9680 36780
rect 8864 36740 9680 36768
rect 5353 36703 5411 36709
rect 5353 36669 5365 36703
rect 5399 36669 5411 36703
rect 5353 36663 5411 36669
rect 5721 36703 5779 36709
rect 5721 36669 5733 36703
rect 5767 36669 5779 36703
rect 5721 36663 5779 36669
rect 6089 36703 6147 36709
rect 6089 36669 6101 36703
rect 6135 36700 6147 36703
rect 6914 36700 6920 36712
rect 6135 36672 6920 36700
rect 6135 36669 6147 36672
rect 6089 36663 6147 36669
rect 5368 36632 5396 36663
rect 6914 36660 6920 36672
rect 6972 36660 6978 36712
rect 7190 36700 7196 36712
rect 7151 36672 7196 36700
rect 7190 36660 7196 36672
rect 7248 36660 7254 36712
rect 7929 36703 7987 36709
rect 7929 36669 7941 36703
rect 7975 36700 7987 36703
rect 8570 36700 8576 36712
rect 7975 36672 8576 36700
rect 7975 36669 7987 36672
rect 7929 36663 7987 36669
rect 8570 36660 8576 36672
rect 8628 36660 8634 36712
rect 8864 36709 8892 36740
rect 9674 36728 9680 36740
rect 9732 36728 9738 36780
rect 8849 36703 8907 36709
rect 8849 36669 8861 36703
rect 8895 36669 8907 36703
rect 8849 36663 8907 36669
rect 9309 36703 9367 36709
rect 9309 36669 9321 36703
rect 9355 36669 9367 36703
rect 10042 36700 10048 36712
rect 10003 36672 10048 36700
rect 9309 36663 9367 36669
rect 5810 36632 5816 36644
rect 5368 36604 5816 36632
rect 5810 36592 5816 36604
rect 5868 36592 5874 36644
rect 8110 36632 8116 36644
rect 7392 36604 8116 36632
rect 7392 36573 7420 36604
rect 8110 36592 8116 36604
rect 8168 36592 8174 36644
rect 9324 36632 9352 36663
rect 10042 36660 10048 36672
rect 10100 36660 10106 36712
rect 10152 36709 10180 36808
rect 22462 36796 22468 36848
rect 22520 36836 22526 36848
rect 24210 36836 24216 36848
rect 22520 36808 24216 36836
rect 22520 36796 22526 36808
rect 24210 36796 24216 36808
rect 24268 36796 24274 36848
rect 24578 36836 24584 36848
rect 24539 36808 24584 36836
rect 24578 36796 24584 36808
rect 24636 36796 24642 36848
rect 31478 36836 31484 36848
rect 31439 36808 31484 36836
rect 31478 36796 31484 36808
rect 31536 36796 31542 36848
rect 31588 36836 31616 36876
rect 33686 36836 33692 36848
rect 31588 36808 33692 36836
rect 33686 36796 33692 36808
rect 33744 36796 33750 36848
rect 10965 36771 11023 36777
rect 10965 36737 10977 36771
rect 11011 36768 11023 36771
rect 11330 36768 11336 36780
rect 11011 36740 11336 36768
rect 11011 36737 11023 36740
rect 10965 36731 11023 36737
rect 11330 36728 11336 36740
rect 11388 36728 11394 36780
rect 15194 36768 15200 36780
rect 14200 36740 15200 36768
rect 10137 36703 10195 36709
rect 10137 36669 10149 36703
rect 10183 36669 10195 36703
rect 10778 36700 10784 36712
rect 10739 36672 10784 36700
rect 10137 36663 10195 36669
rect 10778 36660 10784 36672
rect 10836 36660 10842 36712
rect 11701 36703 11759 36709
rect 11701 36669 11713 36703
rect 11747 36700 11759 36703
rect 11882 36700 11888 36712
rect 11747 36672 11888 36700
rect 11747 36669 11759 36672
rect 11701 36663 11759 36669
rect 11882 36660 11888 36672
rect 11940 36660 11946 36712
rect 12713 36703 12771 36709
rect 12713 36669 12725 36703
rect 12759 36700 12771 36703
rect 13722 36700 13728 36712
rect 12759 36672 13728 36700
rect 12759 36669 12771 36672
rect 12713 36663 12771 36669
rect 13722 36660 13728 36672
rect 13780 36660 13786 36712
rect 13998 36700 14004 36712
rect 13959 36672 14004 36700
rect 13998 36660 14004 36672
rect 14056 36660 14062 36712
rect 14200 36709 14228 36740
rect 15194 36728 15200 36740
rect 15252 36728 15258 36780
rect 17954 36728 17960 36780
rect 18012 36768 18018 36780
rect 18049 36771 18107 36777
rect 18049 36768 18061 36771
rect 18012 36740 18061 36768
rect 18012 36728 18018 36740
rect 18049 36737 18061 36740
rect 18095 36768 18107 36771
rect 20162 36768 20168 36780
rect 18095 36740 20168 36768
rect 18095 36737 18107 36740
rect 18049 36731 18107 36737
rect 20162 36728 20168 36740
rect 20220 36728 20226 36780
rect 24486 36768 24492 36780
rect 20272 36740 24492 36768
rect 14185 36703 14243 36709
rect 14185 36669 14197 36703
rect 14231 36669 14243 36703
rect 14185 36663 14243 36669
rect 14274 36660 14280 36712
rect 14332 36700 14338 36712
rect 14458 36700 14464 36712
rect 14332 36672 14377 36700
rect 14419 36672 14464 36700
rect 14332 36660 14338 36672
rect 14458 36660 14464 36672
rect 14516 36660 14522 36712
rect 14829 36703 14887 36709
rect 14829 36669 14841 36703
rect 14875 36700 14887 36703
rect 15010 36700 15016 36712
rect 14875 36672 15016 36700
rect 14875 36669 14887 36672
rect 14829 36663 14887 36669
rect 15010 36660 15016 36672
rect 15068 36660 15074 36712
rect 15381 36703 15439 36709
rect 15381 36669 15393 36703
rect 15427 36669 15439 36703
rect 15657 36703 15715 36709
rect 15657 36700 15669 36703
rect 15381 36663 15439 36669
rect 15488 36672 15669 36700
rect 13170 36632 13176 36644
rect 9324 36604 13176 36632
rect 13170 36592 13176 36604
rect 13228 36592 13234 36644
rect 13449 36635 13507 36641
rect 13449 36601 13461 36635
rect 13495 36632 13507 36635
rect 15396 36632 15424 36663
rect 13495 36604 15424 36632
rect 13495 36601 13507 36604
rect 13449 36595 13507 36601
rect 7377 36567 7435 36573
rect 7377 36533 7389 36567
rect 7423 36533 7435 36567
rect 8018 36564 8024 36576
rect 7979 36536 8024 36564
rect 7377 36527 7435 36533
rect 8018 36524 8024 36536
rect 8076 36524 8082 36576
rect 11790 36564 11796 36576
rect 11751 36536 11796 36564
rect 11790 36524 11796 36536
rect 11848 36524 11854 36576
rect 12894 36564 12900 36576
rect 12855 36536 12900 36564
rect 12894 36524 12900 36536
rect 12952 36524 12958 36576
rect 13188 36564 13216 36592
rect 15488 36564 15516 36672
rect 15657 36669 15669 36672
rect 15703 36669 15715 36703
rect 15657 36663 15715 36669
rect 18138 36660 18144 36712
rect 18196 36700 18202 36712
rect 18325 36703 18383 36709
rect 18325 36700 18337 36703
rect 18196 36672 18337 36700
rect 18196 36660 18202 36672
rect 18325 36669 18337 36672
rect 18371 36669 18383 36703
rect 18325 36663 18383 36669
rect 15565 36635 15623 36641
rect 15565 36601 15577 36635
rect 15611 36632 15623 36635
rect 15930 36632 15936 36644
rect 15611 36604 15936 36632
rect 15611 36601 15623 36604
rect 15565 36595 15623 36601
rect 15930 36592 15936 36604
rect 15988 36592 15994 36644
rect 19705 36635 19763 36641
rect 19705 36601 19717 36635
rect 19751 36632 19763 36635
rect 20070 36632 20076 36644
rect 19751 36604 20076 36632
rect 19751 36601 19763 36604
rect 19705 36595 19763 36601
rect 20070 36592 20076 36604
rect 20128 36592 20134 36644
rect 13188 36536 15516 36564
rect 15746 36524 15752 36576
rect 15804 36564 15810 36576
rect 20272 36564 20300 36740
rect 24486 36728 24492 36740
rect 24544 36728 24550 36780
rect 25498 36728 25504 36780
rect 25556 36768 25562 36780
rect 25961 36771 26019 36777
rect 25961 36768 25973 36771
rect 25556 36740 25973 36768
rect 25556 36728 25562 36740
rect 25961 36737 25973 36740
rect 26007 36737 26019 36771
rect 25961 36731 26019 36737
rect 26418 36728 26424 36780
rect 26476 36768 26482 36780
rect 27065 36771 27123 36777
rect 27065 36768 27077 36771
rect 26476 36740 27077 36768
rect 26476 36728 26482 36740
rect 27065 36737 27077 36740
rect 27111 36737 27123 36771
rect 27065 36731 27123 36737
rect 27341 36771 27399 36777
rect 27341 36737 27353 36771
rect 27387 36768 27399 36771
rect 27706 36768 27712 36780
rect 27387 36740 27712 36768
rect 27387 36737 27399 36740
rect 27341 36731 27399 36737
rect 20438 36700 20444 36712
rect 20399 36672 20444 36700
rect 20438 36660 20444 36672
rect 20496 36660 20502 36712
rect 20530 36660 20536 36712
rect 20588 36700 20594 36712
rect 22462 36700 22468 36712
rect 20588 36672 21128 36700
rect 22423 36672 22468 36700
rect 20588 36660 20594 36672
rect 21100 36632 21128 36672
rect 22462 36660 22468 36672
rect 22520 36660 22526 36712
rect 22830 36700 22836 36712
rect 22791 36672 22836 36700
rect 22830 36660 22836 36672
rect 22888 36660 22894 36712
rect 24670 36660 24676 36712
rect 24728 36700 24734 36712
rect 24765 36703 24823 36709
rect 24765 36700 24777 36703
rect 24728 36672 24777 36700
rect 24728 36660 24734 36672
rect 24765 36669 24777 36672
rect 24811 36669 24823 36703
rect 25314 36700 25320 36712
rect 25275 36672 25320 36700
rect 24765 36663 24823 36669
rect 25314 36660 25320 36672
rect 25372 36660 25378 36712
rect 25869 36703 25927 36709
rect 25869 36669 25881 36703
rect 25915 36700 25927 36703
rect 26602 36700 26608 36712
rect 25915 36672 26608 36700
rect 25915 36669 25927 36672
rect 25869 36663 25927 36669
rect 26602 36660 26608 36672
rect 26660 36660 26666 36712
rect 27080 36700 27108 36731
rect 27706 36728 27712 36740
rect 27764 36728 27770 36780
rect 28721 36771 28779 36777
rect 28721 36737 28733 36771
rect 28767 36768 28779 36771
rect 28902 36768 28908 36780
rect 28767 36740 28908 36768
rect 28767 36737 28779 36740
rect 28721 36731 28779 36737
rect 28902 36728 28908 36740
rect 28960 36728 28966 36780
rect 29549 36771 29607 36777
rect 29549 36737 29561 36771
rect 29595 36768 29607 36771
rect 30006 36768 30012 36780
rect 29595 36740 30012 36768
rect 29595 36737 29607 36740
rect 29549 36731 29607 36737
rect 30006 36728 30012 36740
rect 30064 36728 30070 36780
rect 35250 36768 35256 36780
rect 30116 36740 35256 36768
rect 29273 36703 29331 36709
rect 29273 36700 29285 36703
rect 27080 36672 29285 36700
rect 29273 36669 29285 36672
rect 29319 36669 29331 36703
rect 30116 36700 30144 36740
rect 35250 36728 35256 36740
rect 35308 36728 35314 36780
rect 31386 36700 31392 36712
rect 29273 36663 29331 36669
rect 29380 36672 30144 36700
rect 31347 36672 31392 36700
rect 21100 36604 26924 36632
rect 15804 36536 20300 36564
rect 15804 36524 15810 36536
rect 20898 36524 20904 36576
rect 20956 36564 20962 36576
rect 21174 36564 21180 36576
rect 20956 36536 21180 36564
rect 20956 36524 20962 36536
rect 21174 36524 21180 36536
rect 21232 36564 21238 36576
rect 21545 36567 21603 36573
rect 21545 36564 21557 36567
rect 21232 36536 21557 36564
rect 21232 36524 21238 36536
rect 21545 36533 21557 36536
rect 21591 36533 21603 36567
rect 22370 36564 22376 36576
rect 22331 36536 22376 36564
rect 21545 36527 21603 36533
rect 22370 36524 22376 36536
rect 22428 36524 22434 36576
rect 25222 36564 25228 36576
rect 25183 36536 25228 36564
rect 25222 36524 25228 36536
rect 25280 36524 25286 36576
rect 26896 36564 26924 36604
rect 29380 36564 29408 36672
rect 31386 36660 31392 36672
rect 31444 36660 31450 36712
rect 26896 36536 29408 36564
rect 30006 36524 30012 36576
rect 30064 36564 30070 36576
rect 30653 36567 30711 36573
rect 30653 36564 30665 36567
rect 30064 36536 30665 36564
rect 30064 36524 30070 36536
rect 30653 36533 30665 36536
rect 30699 36533 30711 36567
rect 30653 36527 30711 36533
rect 1104 36474 39836 36496
rect 1104 36422 19606 36474
rect 19658 36422 19670 36474
rect 19722 36422 19734 36474
rect 19786 36422 19798 36474
rect 19850 36422 39836 36474
rect 1104 36400 39836 36422
rect 7466 36360 7472 36372
rect 7427 36332 7472 36360
rect 7466 36320 7472 36332
rect 7524 36360 7530 36372
rect 7834 36360 7840 36372
rect 7524 36332 7840 36360
rect 7524 36320 7530 36332
rect 7834 36320 7840 36332
rect 7892 36320 7898 36372
rect 12894 36360 12900 36372
rect 11716 36332 12900 36360
rect 5718 36292 5724 36304
rect 4816 36264 5724 36292
rect 4816 36233 4844 36264
rect 5718 36252 5724 36264
rect 5776 36252 5782 36304
rect 7190 36252 7196 36304
rect 7248 36292 7254 36304
rect 11716 36292 11744 36332
rect 12894 36320 12900 36332
rect 12952 36320 12958 36372
rect 25498 36360 25504 36372
rect 25459 36332 25504 36360
rect 25498 36320 25504 36332
rect 25556 36320 25562 36372
rect 12710 36292 12716 36304
rect 7248 36264 8156 36292
rect 7248 36252 7254 36264
rect 4801 36227 4859 36233
rect 4801 36193 4813 36227
rect 4847 36193 4859 36227
rect 4801 36187 4859 36193
rect 5353 36227 5411 36233
rect 5353 36193 5365 36227
rect 5399 36224 5411 36227
rect 5534 36224 5540 36236
rect 5399 36196 5540 36224
rect 5399 36193 5411 36196
rect 5353 36187 5411 36193
rect 5534 36184 5540 36196
rect 5592 36224 5598 36236
rect 6730 36224 6736 36236
rect 5592 36196 6736 36224
rect 5592 36184 5598 36196
rect 6730 36184 6736 36196
rect 6788 36184 6794 36236
rect 7374 36224 7380 36236
rect 7335 36196 7380 36224
rect 7374 36184 7380 36196
rect 7432 36184 7438 36236
rect 8128 36233 8156 36264
rect 9968 36264 10824 36292
rect 8113 36227 8171 36233
rect 8113 36193 8125 36227
rect 8159 36193 8171 36227
rect 8113 36187 8171 36193
rect 8570 36184 8576 36236
rect 8628 36224 8634 36236
rect 8849 36227 8907 36233
rect 8849 36224 8861 36227
rect 8628 36196 8861 36224
rect 8628 36184 8634 36196
rect 8849 36193 8861 36196
rect 8895 36224 8907 36227
rect 9398 36224 9404 36236
rect 8895 36196 9404 36224
rect 8895 36193 8907 36196
rect 8849 36187 8907 36193
rect 9398 36184 9404 36196
rect 9456 36184 9462 36236
rect 9968 36233 9996 36264
rect 10796 36236 10824 36264
rect 11624 36264 11744 36292
rect 12360 36264 12716 36292
rect 9953 36227 10011 36233
rect 9953 36193 9965 36227
rect 9999 36193 10011 36227
rect 10318 36224 10324 36236
rect 10279 36196 10324 36224
rect 9953 36187 10011 36193
rect 10318 36184 10324 36196
rect 10376 36184 10382 36236
rect 10689 36227 10747 36233
rect 10689 36193 10701 36227
rect 10735 36193 10747 36227
rect 10689 36187 10747 36193
rect 5445 36159 5503 36165
rect 5445 36125 5457 36159
rect 5491 36125 5503 36159
rect 7466 36156 7472 36168
rect 7379 36128 7472 36156
rect 5445 36119 5503 36125
rect 4893 36091 4951 36097
rect 4893 36057 4905 36091
rect 4939 36088 4951 36091
rect 4982 36088 4988 36100
rect 4939 36060 4988 36088
rect 4939 36057 4951 36060
rect 4893 36051 4951 36057
rect 4982 36048 4988 36060
rect 5040 36048 5046 36100
rect 5350 36048 5356 36100
rect 5408 36088 5414 36100
rect 5460 36088 5488 36119
rect 7466 36116 7472 36128
rect 7524 36156 7530 36168
rect 8205 36159 8263 36165
rect 8205 36156 8217 36159
rect 7524 36128 8217 36156
rect 7524 36116 7530 36128
rect 8205 36125 8217 36128
rect 8251 36125 8263 36159
rect 10704 36156 10732 36187
rect 10778 36184 10784 36236
rect 10836 36224 10842 36236
rect 11624 36233 11652 36264
rect 11609 36227 11667 36233
rect 11609 36224 11621 36227
rect 10836 36196 11621 36224
rect 10836 36184 10842 36196
rect 11609 36193 11621 36196
rect 11655 36193 11667 36227
rect 11790 36224 11796 36236
rect 11751 36196 11796 36224
rect 11609 36187 11667 36193
rect 11790 36184 11796 36196
rect 11848 36184 11854 36236
rect 12360 36233 12388 36264
rect 12710 36252 12716 36264
rect 12768 36252 12774 36304
rect 14090 36252 14096 36304
rect 14148 36292 14154 36304
rect 14185 36295 14243 36301
rect 14185 36292 14197 36295
rect 14148 36264 14197 36292
rect 14148 36252 14154 36264
rect 14185 36261 14197 36264
rect 14231 36261 14243 36295
rect 14185 36255 14243 36261
rect 20349 36295 20407 36301
rect 20349 36261 20361 36295
rect 20395 36292 20407 36295
rect 20438 36292 20444 36304
rect 20395 36264 20444 36292
rect 20395 36261 20407 36264
rect 20349 36255 20407 36261
rect 20438 36252 20444 36264
rect 20496 36252 20502 36304
rect 12345 36227 12403 36233
rect 12345 36193 12357 36227
rect 12391 36193 12403 36227
rect 12526 36224 12532 36236
rect 12487 36196 12532 36224
rect 12345 36187 12403 36193
rect 12526 36184 12532 36196
rect 12584 36184 12590 36236
rect 13722 36224 13728 36236
rect 13635 36196 13728 36224
rect 13722 36184 13728 36196
rect 13780 36184 13786 36236
rect 13906 36224 13912 36236
rect 13867 36196 13912 36224
rect 13906 36184 13912 36196
rect 13964 36184 13970 36236
rect 14274 36184 14280 36236
rect 14332 36224 14338 36236
rect 15289 36227 15347 36233
rect 15289 36224 15301 36227
rect 14332 36196 15301 36224
rect 14332 36184 14338 36196
rect 15289 36193 15301 36196
rect 15335 36193 15347 36227
rect 15289 36187 15347 36193
rect 17954 36184 17960 36236
rect 18012 36224 18018 36236
rect 18690 36224 18696 36236
rect 18012 36196 18696 36224
rect 18012 36184 18018 36196
rect 18690 36184 18696 36196
rect 18748 36184 18754 36236
rect 20898 36224 20904 36236
rect 20859 36196 20904 36224
rect 20898 36184 20904 36196
rect 20956 36184 20962 36236
rect 22646 36224 22652 36236
rect 22607 36196 22652 36224
rect 22646 36184 22652 36196
rect 22704 36184 22710 36236
rect 23106 36224 23112 36236
rect 23067 36196 23112 36224
rect 23106 36184 23112 36196
rect 23164 36184 23170 36236
rect 30006 36224 30012 36236
rect 29967 36196 30012 36224
rect 30006 36184 30012 36196
rect 30064 36184 30070 36236
rect 32122 36224 32128 36236
rect 32035 36196 32128 36224
rect 32122 36184 32128 36196
rect 32180 36224 32186 36236
rect 33594 36224 33600 36236
rect 32180 36196 33600 36224
rect 32180 36184 32186 36196
rect 33594 36184 33600 36196
rect 33652 36224 33658 36236
rect 34241 36227 34299 36233
rect 34241 36224 34253 36227
rect 33652 36196 34253 36224
rect 33652 36184 33658 36196
rect 34241 36193 34253 36196
rect 34287 36193 34299 36227
rect 34241 36187 34299 36193
rect 11238 36156 11244 36168
rect 10704 36128 11244 36156
rect 8205 36119 8263 36125
rect 11238 36116 11244 36128
rect 11296 36156 11302 36168
rect 11808 36156 11836 36184
rect 11296 36128 11836 36156
rect 13740 36156 13768 36184
rect 15381 36159 15439 36165
rect 15381 36156 15393 36159
rect 13740 36128 15393 36156
rect 11296 36116 11302 36128
rect 15381 36125 15393 36128
rect 15427 36125 15439 36159
rect 15381 36119 15439 36125
rect 16393 36159 16451 36165
rect 16393 36125 16405 36159
rect 16439 36125 16451 36159
rect 16666 36156 16672 36168
rect 16627 36128 16672 36156
rect 16393 36119 16451 36125
rect 5408 36060 5488 36088
rect 5408 36048 5414 36060
rect 10042 36048 10048 36100
rect 10100 36088 10106 36100
rect 10597 36091 10655 36097
rect 10597 36088 10609 36091
rect 10100 36060 10609 36088
rect 10100 36048 10106 36060
rect 10597 36057 10609 36060
rect 10643 36057 10655 36091
rect 10597 36051 10655 36057
rect 12713 36091 12771 36097
rect 12713 36057 12725 36091
rect 12759 36088 12771 36091
rect 13814 36088 13820 36100
rect 12759 36060 13820 36088
rect 12759 36057 12771 36060
rect 12713 36051 12771 36057
rect 13814 36048 13820 36060
rect 13872 36048 13878 36100
rect 15286 36048 15292 36100
rect 15344 36088 15350 36100
rect 16408 36088 16436 36119
rect 16666 36116 16672 36128
rect 16724 36116 16730 36168
rect 18969 36159 19027 36165
rect 18969 36125 18981 36159
rect 19015 36156 19027 36159
rect 20070 36156 20076 36168
rect 19015 36128 20076 36156
rect 19015 36125 19027 36128
rect 18969 36119 19027 36125
rect 20070 36116 20076 36128
rect 20128 36116 20134 36168
rect 24118 36156 24124 36168
rect 24079 36128 24124 36156
rect 24118 36116 24124 36128
rect 24176 36116 24182 36168
rect 24394 36156 24400 36168
rect 24355 36128 24400 36156
rect 24394 36116 24400 36128
rect 24452 36116 24458 36168
rect 26326 36116 26332 36168
rect 26384 36156 26390 36168
rect 27341 36159 27399 36165
rect 27341 36156 27353 36159
rect 26384 36128 27353 36156
rect 26384 36116 26390 36128
rect 27341 36125 27353 36128
rect 27387 36125 27399 36159
rect 27341 36119 27399 36125
rect 27617 36159 27675 36165
rect 27617 36125 27629 36159
rect 27663 36156 27675 36159
rect 29638 36156 29644 36168
rect 27663 36128 29644 36156
rect 27663 36125 27675 36128
rect 27617 36119 27675 36125
rect 29638 36116 29644 36128
rect 29696 36116 29702 36168
rect 29730 36116 29736 36168
rect 29788 36156 29794 36168
rect 32398 36156 32404 36168
rect 29788 36128 29833 36156
rect 32359 36128 32404 36156
rect 29788 36116 29794 36128
rect 32398 36116 32404 36128
rect 32456 36116 32462 36168
rect 34514 36156 34520 36168
rect 34475 36128 34520 36156
rect 34514 36116 34520 36128
rect 34572 36116 34578 36168
rect 15344 36060 16436 36088
rect 15344 36048 15350 36060
rect 22830 36048 22836 36100
rect 22888 36088 22894 36100
rect 23017 36091 23075 36097
rect 23017 36088 23029 36091
rect 22888 36060 23029 36088
rect 22888 36048 22894 36060
rect 23017 36057 23029 36060
rect 23063 36057 23075 36091
rect 23017 36051 23075 36057
rect 9030 36020 9036 36032
rect 8991 35992 9036 36020
rect 9030 35980 9036 35992
rect 9088 35980 9094 36032
rect 17957 36023 18015 36029
rect 17957 35989 17969 36023
rect 18003 36020 18015 36023
rect 18138 36020 18144 36032
rect 18003 35992 18144 36020
rect 18003 35989 18015 35992
rect 17957 35983 18015 35989
rect 18138 35980 18144 35992
rect 18196 35980 18202 36032
rect 18230 35980 18236 36032
rect 18288 36020 18294 36032
rect 20806 36020 20812 36032
rect 18288 35992 20812 36020
rect 18288 35980 18294 35992
rect 20806 35980 20812 35992
rect 20864 35980 20870 36032
rect 20990 36020 20996 36032
rect 20951 35992 20996 36020
rect 20990 35980 20996 35992
rect 21048 35980 21054 36032
rect 27338 35980 27344 36032
rect 27396 36020 27402 36032
rect 28721 36023 28779 36029
rect 28721 36020 28733 36023
rect 27396 35992 28733 36020
rect 27396 35980 27402 35992
rect 28721 35989 28733 35992
rect 28767 35989 28779 36023
rect 31110 36020 31116 36032
rect 31071 35992 31116 36020
rect 28721 35983 28779 35989
rect 31110 35980 31116 35992
rect 31168 35980 31174 36032
rect 33502 36020 33508 36032
rect 33463 35992 33508 36020
rect 33502 35980 33508 35992
rect 33560 35980 33566 36032
rect 35618 36020 35624 36032
rect 35579 35992 35624 36020
rect 35618 35980 35624 35992
rect 35676 35980 35682 36032
rect 1104 35930 39836 35952
rect 1104 35878 4246 35930
rect 4298 35878 4310 35930
rect 4362 35878 4374 35930
rect 4426 35878 4438 35930
rect 4490 35878 34966 35930
rect 35018 35878 35030 35930
rect 35082 35878 35094 35930
rect 35146 35878 35158 35930
rect 35210 35878 39836 35930
rect 1104 35856 39836 35878
rect 7929 35819 7987 35825
rect 7929 35816 7941 35819
rect 1688 35788 7941 35816
rect 1688 35612 1716 35788
rect 7929 35785 7941 35788
rect 7975 35785 7987 35819
rect 9398 35816 9404 35828
rect 9359 35788 9404 35816
rect 7929 35779 7987 35785
rect 9398 35776 9404 35788
rect 9456 35776 9462 35828
rect 12253 35819 12311 35825
rect 12253 35785 12265 35819
rect 12299 35816 12311 35819
rect 15746 35816 15752 35828
rect 12299 35788 15752 35816
rect 12299 35785 12311 35788
rect 12253 35779 12311 35785
rect 15746 35776 15752 35788
rect 15804 35776 15810 35828
rect 16666 35816 16672 35828
rect 16627 35788 16672 35816
rect 16666 35776 16672 35788
rect 16724 35776 16730 35828
rect 18046 35776 18052 35828
rect 18104 35816 18110 35828
rect 18325 35819 18383 35825
rect 18325 35816 18337 35819
rect 18104 35788 18337 35816
rect 18104 35776 18110 35788
rect 18325 35785 18337 35788
rect 18371 35785 18383 35819
rect 18325 35779 18383 35785
rect 18690 35776 18696 35828
rect 18748 35816 18754 35828
rect 19061 35819 19119 35825
rect 19061 35816 19073 35819
rect 18748 35788 19073 35816
rect 18748 35776 18754 35788
rect 19061 35785 19073 35788
rect 19107 35785 19119 35819
rect 19061 35779 19119 35785
rect 20809 35819 20867 35825
rect 20809 35785 20821 35819
rect 20855 35816 20867 35819
rect 22462 35816 22468 35828
rect 20855 35788 22468 35816
rect 20855 35785 20867 35788
rect 20809 35779 20867 35785
rect 22462 35776 22468 35788
rect 22520 35776 22526 35828
rect 22646 35816 22652 35828
rect 22607 35788 22652 35816
rect 22646 35776 22652 35788
rect 22704 35776 22710 35828
rect 26436 35788 29408 35816
rect 5810 35748 5816 35760
rect 5771 35720 5816 35748
rect 5810 35708 5816 35720
rect 5868 35708 5874 35760
rect 10962 35708 10968 35760
rect 11020 35748 11026 35760
rect 11057 35751 11115 35757
rect 11057 35748 11069 35751
rect 11020 35720 11069 35748
rect 11020 35708 11026 35720
rect 11057 35717 11069 35720
rect 11103 35717 11115 35751
rect 13906 35748 13912 35760
rect 11057 35711 11115 35717
rect 12452 35720 13912 35748
rect 5169 35683 5227 35689
rect 5169 35649 5181 35683
rect 5215 35680 5227 35683
rect 5534 35680 5540 35692
rect 5215 35652 5540 35680
rect 5215 35649 5227 35652
rect 5169 35643 5227 35649
rect 5534 35640 5540 35652
rect 5592 35640 5598 35692
rect 7466 35680 7472 35692
rect 5920 35652 7472 35680
rect 1765 35615 1823 35621
rect 1765 35612 1777 35615
rect 1688 35584 1777 35612
rect 1765 35581 1777 35584
rect 1811 35581 1823 35615
rect 3786 35612 3792 35624
rect 3747 35584 3792 35612
rect 1765 35575 1823 35581
rect 3786 35572 3792 35584
rect 3844 35572 3850 35624
rect 4154 35572 4160 35624
rect 4212 35612 4218 35624
rect 5350 35612 5356 35624
rect 4212 35584 5356 35612
rect 4212 35572 4218 35584
rect 5350 35572 5356 35584
rect 5408 35572 5414 35624
rect 5920 35621 5948 35652
rect 7466 35640 7472 35652
rect 7524 35640 7530 35692
rect 7742 35640 7748 35692
rect 7800 35680 7806 35692
rect 8021 35683 8079 35689
rect 8021 35680 8033 35683
rect 7800 35652 8033 35680
rect 7800 35640 7806 35652
rect 8021 35649 8033 35652
rect 8067 35680 8079 35683
rect 9858 35680 9864 35692
rect 8067 35652 9864 35680
rect 8067 35649 8079 35652
rect 8021 35643 8079 35649
rect 9858 35640 9864 35652
rect 9916 35640 9922 35692
rect 11238 35680 11244 35692
rect 11199 35652 11244 35680
rect 11238 35640 11244 35652
rect 11296 35640 11302 35692
rect 12452 35680 12480 35720
rect 13906 35708 13912 35720
rect 13964 35708 13970 35760
rect 22480 35748 22508 35776
rect 24394 35748 24400 35760
rect 22480 35720 23980 35748
rect 24355 35720 24400 35748
rect 11624 35652 12480 35680
rect 11624 35624 11652 35652
rect 12526 35640 12532 35692
rect 12584 35680 12590 35692
rect 13265 35683 13323 35689
rect 13265 35680 13277 35683
rect 12584 35652 13277 35680
rect 12584 35640 12590 35652
rect 13265 35649 13277 35652
rect 13311 35649 13323 35683
rect 13265 35643 13323 35649
rect 14277 35683 14335 35689
rect 14277 35649 14289 35683
rect 14323 35680 14335 35683
rect 14918 35680 14924 35692
rect 14323 35652 14924 35680
rect 14323 35649 14335 35652
rect 14277 35643 14335 35649
rect 14918 35640 14924 35652
rect 14976 35680 14982 35692
rect 15565 35683 15623 35689
rect 14976 35652 15516 35680
rect 14976 35640 14982 35652
rect 5905 35615 5963 35621
rect 5905 35581 5917 35615
rect 5951 35581 5963 35615
rect 6822 35612 6828 35624
rect 6783 35584 6828 35612
rect 5905 35575 5963 35581
rect 6822 35572 6828 35584
rect 6880 35572 6886 35624
rect 8294 35612 8300 35624
rect 8255 35584 8300 35612
rect 8294 35572 8300 35584
rect 8352 35572 8358 35624
rect 10597 35615 10655 35621
rect 10597 35581 10609 35615
rect 10643 35612 10655 35615
rect 10778 35612 10784 35624
rect 10643 35584 10784 35612
rect 10643 35581 10655 35584
rect 10597 35575 10655 35581
rect 10778 35572 10784 35584
rect 10836 35572 10842 35624
rect 11149 35615 11207 35621
rect 11149 35581 11161 35615
rect 11195 35612 11207 35615
rect 11606 35612 11612 35624
rect 11195 35584 11612 35612
rect 11195 35581 11207 35584
rect 11149 35575 11207 35581
rect 11606 35572 11612 35584
rect 11664 35572 11670 35624
rect 12434 35572 12440 35624
rect 12492 35612 12498 35624
rect 12492 35584 12537 35612
rect 12492 35572 12498 35584
rect 12894 35572 12900 35624
rect 12952 35612 12958 35624
rect 12989 35615 13047 35621
rect 12989 35612 13001 35615
rect 12952 35584 13001 35612
rect 12952 35572 12958 35584
rect 12989 35581 13001 35584
rect 13035 35581 13047 35615
rect 12989 35575 13047 35581
rect 14366 35572 14372 35624
rect 14424 35612 14430 35624
rect 15286 35612 15292 35624
rect 14424 35584 14469 35612
rect 15247 35584 15292 35612
rect 14424 35572 14430 35584
rect 15286 35572 15292 35584
rect 15344 35572 15350 35624
rect 15488 35612 15516 35652
rect 15565 35649 15577 35683
rect 15611 35680 15623 35683
rect 16022 35680 16028 35692
rect 15611 35652 16028 35680
rect 15611 35649 15623 35652
rect 15565 35643 15623 35649
rect 16022 35640 16028 35652
rect 16080 35640 16086 35692
rect 20438 35680 20444 35692
rect 19996 35652 20444 35680
rect 18049 35615 18107 35621
rect 18049 35612 18061 35615
rect 15488 35584 18061 35612
rect 18049 35581 18061 35584
rect 18095 35581 18107 35615
rect 18049 35575 18107 35581
rect 18141 35615 18199 35621
rect 18141 35581 18153 35615
rect 18187 35581 18199 35615
rect 19242 35612 19248 35624
rect 19203 35584 19248 35612
rect 18141 35575 18199 35581
rect 14826 35544 14832 35556
rect 14787 35516 14832 35544
rect 14826 35504 14832 35516
rect 14884 35504 14890 35556
rect 18156 35544 18184 35575
rect 19242 35572 19248 35584
rect 19300 35572 19306 35624
rect 19996 35621 20024 35652
rect 20438 35640 20444 35652
rect 20496 35640 20502 35692
rect 21269 35683 21327 35689
rect 21269 35649 21281 35683
rect 21315 35680 21327 35683
rect 21450 35680 21456 35692
rect 21315 35652 21456 35680
rect 21315 35649 21327 35652
rect 21269 35643 21327 35649
rect 21450 35640 21456 35652
rect 21508 35640 21514 35692
rect 21545 35683 21603 35689
rect 21545 35649 21557 35683
rect 21591 35680 21603 35683
rect 22370 35680 22376 35692
rect 21591 35652 22376 35680
rect 21591 35649 21603 35652
rect 21545 35643 21603 35649
rect 22370 35640 22376 35652
rect 22428 35640 22434 35692
rect 23952 35624 23980 35720
rect 24394 35708 24400 35720
rect 24452 35708 24458 35760
rect 25130 35708 25136 35760
rect 25188 35748 25194 35760
rect 25188 35720 25452 35748
rect 25188 35708 25194 35720
rect 24581 35683 24639 35689
rect 24581 35649 24593 35683
rect 24627 35680 24639 35683
rect 24762 35680 24768 35692
rect 24627 35652 24768 35680
rect 24627 35649 24639 35652
rect 24581 35643 24639 35649
rect 24762 35640 24768 35652
rect 24820 35680 24826 35692
rect 25424 35680 25452 35720
rect 26436 35680 26464 35788
rect 27157 35751 27215 35757
rect 27157 35717 27169 35751
rect 27203 35717 27215 35751
rect 27157 35711 27215 35717
rect 24820 35652 25360 35680
rect 25424 35652 26464 35680
rect 27172 35680 27200 35711
rect 27706 35708 27712 35760
rect 27764 35748 27770 35760
rect 29273 35751 29331 35757
rect 29273 35748 29285 35751
rect 27764 35720 29285 35748
rect 27764 35708 27770 35720
rect 29273 35717 29285 35720
rect 29319 35717 29331 35751
rect 29380 35748 29408 35788
rect 29638 35776 29644 35828
rect 29696 35816 29702 35828
rect 29733 35819 29791 35825
rect 29733 35816 29745 35819
rect 29696 35788 29745 35816
rect 29696 35776 29702 35788
rect 29733 35785 29745 35788
rect 29779 35785 29791 35819
rect 32398 35816 32404 35828
rect 32359 35788 32404 35816
rect 29733 35779 29791 35785
rect 32398 35776 32404 35788
rect 32456 35776 32462 35828
rect 33226 35816 33232 35828
rect 33187 35788 33232 35816
rect 33226 35776 33232 35788
rect 33284 35776 33290 35828
rect 30834 35748 30840 35760
rect 29380 35720 30840 35748
rect 29273 35711 29331 35717
rect 30834 35708 30840 35720
rect 30892 35708 30898 35760
rect 31110 35680 31116 35692
rect 27172 35652 29592 35680
rect 31071 35652 31116 35680
rect 24820 35640 24826 35652
rect 19981 35615 20039 35621
rect 19981 35581 19993 35615
rect 20027 35581 20039 35615
rect 19981 35575 20039 35581
rect 20070 35572 20076 35624
rect 20128 35612 20134 35624
rect 20165 35615 20223 35621
rect 20165 35612 20177 35615
rect 20128 35584 20177 35612
rect 20128 35572 20134 35584
rect 20165 35581 20177 35584
rect 20211 35581 20223 35615
rect 20165 35575 20223 35581
rect 20533 35615 20591 35621
rect 20533 35581 20545 35615
rect 20579 35612 20591 35615
rect 20990 35612 20996 35624
rect 20579 35584 20996 35612
rect 20579 35581 20591 35584
rect 20533 35575 20591 35581
rect 20990 35572 20996 35584
rect 21048 35572 21054 35624
rect 23934 35612 23940 35624
rect 21376 35584 23796 35612
rect 23895 35584 23940 35612
rect 21376 35544 21404 35584
rect 18156 35516 21404 35544
rect 23768 35544 23796 35584
rect 23934 35572 23940 35584
rect 23992 35572 23998 35624
rect 24489 35615 24547 35621
rect 24489 35581 24501 35615
rect 24535 35612 24547 35615
rect 25222 35612 25228 35624
rect 24535 35584 25228 35612
rect 24535 35581 24547 35584
rect 24489 35575 24547 35581
rect 25222 35572 25228 35584
rect 25280 35572 25286 35624
rect 25130 35544 25136 35556
rect 23768 35516 25136 35544
rect 25130 35504 25136 35516
rect 25188 35504 25194 35556
rect 25332 35544 25360 35652
rect 25498 35612 25504 35624
rect 25459 35584 25504 35612
rect 25498 35572 25504 35584
rect 25556 35572 25562 35624
rect 26145 35615 26203 35621
rect 26145 35581 26157 35615
rect 26191 35612 26203 35615
rect 26234 35612 26240 35624
rect 26191 35584 26240 35612
rect 26191 35581 26203 35584
rect 26145 35575 26203 35581
rect 26234 35572 26240 35584
rect 26292 35572 26298 35624
rect 26329 35615 26387 35621
rect 26329 35581 26341 35615
rect 26375 35612 26387 35615
rect 26786 35612 26792 35624
rect 26375 35584 26792 35612
rect 26375 35581 26387 35584
rect 26329 35575 26387 35581
rect 26786 35572 26792 35584
rect 26844 35612 26850 35624
rect 27338 35612 27344 35624
rect 26844 35584 27344 35612
rect 26844 35572 26850 35584
rect 27338 35572 27344 35584
rect 27396 35572 27402 35624
rect 27525 35615 27583 35621
rect 27525 35581 27537 35615
rect 27571 35581 27583 35615
rect 27525 35575 27583 35581
rect 26421 35547 26479 35553
rect 26421 35544 26433 35547
rect 25332 35516 26433 35544
rect 26421 35513 26433 35516
rect 26467 35513 26479 35547
rect 26421 35507 26479 35513
rect 27062 35504 27068 35556
rect 27120 35544 27126 35556
rect 27540 35544 27568 35575
rect 27614 35572 27620 35624
rect 27672 35612 27678 35624
rect 29564 35621 29592 35652
rect 31110 35640 31116 35652
rect 31168 35640 31174 35692
rect 27709 35615 27767 35621
rect 27709 35612 27721 35615
rect 27672 35584 27721 35612
rect 27672 35572 27678 35584
rect 27709 35581 27721 35584
rect 27755 35581 27767 35615
rect 27709 35575 27767 35581
rect 29549 35615 29607 35621
rect 29549 35581 29561 35615
rect 29595 35581 29607 35615
rect 29549 35575 29607 35581
rect 29730 35572 29736 35624
rect 29788 35612 29794 35624
rect 30837 35615 30895 35621
rect 30837 35612 30849 35615
rect 29788 35584 30849 35612
rect 29788 35572 29794 35584
rect 30837 35581 30849 35584
rect 30883 35612 30895 35615
rect 32122 35612 32128 35624
rect 30883 35584 32128 35612
rect 30883 35581 30895 35584
rect 30837 35575 30895 35581
rect 32122 35572 32128 35584
rect 32180 35572 32186 35624
rect 32953 35615 33011 35621
rect 32953 35581 32965 35615
rect 32999 35581 33011 35615
rect 32953 35575 33011 35581
rect 27120 35516 27568 35544
rect 29457 35547 29515 35553
rect 27120 35504 27126 35516
rect 29457 35513 29469 35547
rect 29503 35513 29515 35547
rect 29457 35507 29515 35513
rect 1949 35479 2007 35485
rect 1949 35445 1961 35479
rect 1995 35476 2007 35479
rect 2866 35476 2872 35488
rect 1995 35448 2872 35476
rect 1995 35445 2007 35448
rect 1949 35439 2007 35445
rect 2866 35436 2872 35448
rect 2924 35436 2930 35488
rect 3973 35479 4031 35485
rect 3973 35445 3985 35479
rect 4019 35476 4031 35479
rect 4154 35476 4160 35488
rect 4019 35448 4160 35476
rect 4019 35445 4031 35448
rect 3973 35439 4031 35445
rect 4154 35436 4160 35448
rect 4212 35436 4218 35488
rect 6730 35436 6736 35488
rect 6788 35476 6794 35488
rect 7009 35479 7067 35485
rect 7009 35476 7021 35479
rect 6788 35448 7021 35476
rect 6788 35436 6794 35448
rect 7009 35445 7021 35448
rect 7055 35445 7067 35479
rect 7009 35439 7067 35445
rect 7929 35479 7987 35485
rect 7929 35445 7941 35479
rect 7975 35476 7987 35479
rect 12253 35479 12311 35485
rect 12253 35476 12265 35479
rect 7975 35448 12265 35476
rect 7975 35445 7987 35448
rect 7929 35439 7987 35445
rect 12253 35445 12265 35448
rect 12299 35445 12311 35479
rect 12253 35439 12311 35445
rect 12529 35479 12587 35485
rect 12529 35445 12541 35479
rect 12575 35476 12587 35479
rect 13078 35476 13084 35488
rect 12575 35448 13084 35476
rect 12575 35445 12587 35448
rect 12529 35439 12587 35445
rect 13078 35436 13084 35448
rect 13136 35436 13142 35488
rect 24118 35436 24124 35488
rect 24176 35476 24182 35488
rect 26326 35476 26332 35488
rect 24176 35448 26332 35476
rect 24176 35436 24182 35448
rect 26326 35436 26332 35448
rect 26384 35436 26390 35488
rect 26602 35436 26608 35488
rect 26660 35476 26666 35488
rect 29472 35476 29500 35507
rect 26660 35448 29500 35476
rect 26660 35436 26666 35448
rect 30742 35436 30748 35488
rect 30800 35476 30806 35488
rect 31570 35476 31576 35488
rect 30800 35448 31576 35476
rect 30800 35436 30806 35448
rect 31570 35436 31576 35448
rect 31628 35476 31634 35488
rect 32968 35476 32996 35575
rect 33042 35572 33048 35624
rect 33100 35612 33106 35624
rect 33100 35584 33145 35612
rect 33100 35572 33106 35584
rect 31628 35448 32996 35476
rect 31628 35436 31634 35448
rect 1104 35386 39836 35408
rect 1104 35334 19606 35386
rect 19658 35334 19670 35386
rect 19722 35334 19734 35386
rect 19786 35334 19798 35386
rect 19850 35334 39836 35386
rect 1104 35312 39836 35334
rect 11793 35275 11851 35281
rect 11793 35272 11805 35275
rect 10428 35244 11805 35272
rect 6365 35207 6423 35213
rect 6365 35173 6377 35207
rect 6411 35204 6423 35207
rect 6638 35204 6644 35216
rect 6411 35176 6644 35204
rect 6411 35173 6423 35176
rect 6365 35167 6423 35173
rect 6638 35164 6644 35176
rect 6696 35204 6702 35216
rect 6696 35176 8984 35204
rect 6696 35164 6702 35176
rect 1946 35096 1952 35148
rect 2004 35136 2010 35148
rect 4065 35139 4123 35145
rect 4065 35136 4077 35139
rect 2004 35108 4077 35136
rect 2004 35096 2010 35108
rect 4065 35105 4077 35108
rect 4111 35136 4123 35139
rect 4154 35136 4160 35148
rect 4111 35108 4160 35136
rect 4111 35105 4123 35108
rect 4065 35099 4123 35105
rect 4154 35096 4160 35108
rect 4212 35096 4218 35148
rect 4982 35136 4988 35148
rect 4943 35108 4988 35136
rect 4982 35096 4988 35108
rect 5040 35096 5046 35148
rect 6822 35096 6828 35148
rect 6880 35136 6886 35148
rect 7285 35139 7343 35145
rect 7285 35136 7297 35139
rect 6880 35108 7297 35136
rect 6880 35096 6886 35108
rect 7285 35105 7297 35108
rect 7331 35105 7343 35139
rect 7466 35136 7472 35148
rect 7427 35108 7472 35136
rect 7285 35099 7343 35105
rect 1397 35071 1455 35077
rect 1397 35037 1409 35071
rect 1443 35037 1455 35071
rect 1397 35031 1455 35037
rect 1673 35071 1731 35077
rect 1673 35037 1685 35071
rect 1719 35068 1731 35071
rect 2130 35068 2136 35080
rect 1719 35040 2136 35068
rect 1719 35037 1731 35040
rect 1673 35031 1731 35037
rect 1412 34932 1440 35031
rect 2130 35028 2136 35040
rect 2188 35028 2194 35080
rect 2682 35028 2688 35080
rect 2740 35068 2746 35080
rect 4709 35071 4767 35077
rect 4709 35068 4721 35071
rect 2740 35040 4721 35068
rect 2740 35028 2746 35040
rect 4709 35037 4721 35040
rect 4755 35068 4767 35071
rect 6086 35068 6092 35080
rect 4755 35040 6092 35068
rect 4755 35037 4767 35040
rect 4709 35031 4767 35037
rect 6086 35028 6092 35040
rect 6144 35028 6150 35080
rect 7300 35068 7328 35099
rect 7466 35096 7472 35108
rect 7524 35096 7530 35148
rect 8018 35136 8024 35148
rect 7979 35108 8024 35136
rect 8018 35096 8024 35108
rect 8076 35096 8082 35148
rect 8202 35136 8208 35148
rect 8163 35108 8208 35136
rect 8202 35096 8208 35108
rect 8260 35096 8266 35148
rect 8956 35145 8984 35176
rect 8941 35139 8999 35145
rect 8941 35105 8953 35139
rect 8987 35105 8999 35139
rect 8941 35099 8999 35105
rect 10318 35096 10324 35148
rect 10376 35136 10382 35148
rect 10428 35145 10456 35244
rect 11793 35241 11805 35244
rect 11839 35272 11851 35275
rect 12526 35272 12532 35284
rect 11839 35244 12532 35272
rect 11839 35241 11851 35244
rect 11793 35235 11851 35241
rect 12526 35232 12532 35244
rect 12584 35232 12590 35284
rect 24670 35232 24676 35284
rect 24728 35272 24734 35284
rect 35986 35272 35992 35284
rect 24728 35244 26372 35272
rect 24728 35232 24734 35244
rect 11149 35207 11207 35213
rect 11149 35173 11161 35207
rect 11195 35204 11207 35207
rect 12434 35204 12440 35216
rect 11195 35176 12440 35204
rect 11195 35173 11207 35176
rect 11149 35167 11207 35173
rect 12434 35164 12440 35176
rect 12492 35164 12498 35216
rect 23845 35207 23903 35213
rect 23216 35176 23520 35204
rect 10413 35139 10471 35145
rect 10413 35136 10425 35139
rect 10376 35108 10425 35136
rect 10376 35096 10382 35108
rect 10413 35105 10425 35108
rect 10459 35105 10471 35139
rect 10413 35099 10471 35105
rect 10873 35139 10931 35145
rect 10873 35105 10885 35139
rect 10919 35105 10931 35139
rect 11606 35136 11612 35148
rect 11567 35108 11612 35136
rect 10873 35099 10931 35105
rect 9033 35071 9091 35077
rect 9033 35068 9045 35071
rect 7300 35040 9045 35068
rect 9033 35037 9045 35040
rect 9079 35037 9091 35071
rect 9033 35031 9091 35037
rect 10229 35071 10287 35077
rect 10229 35037 10241 35071
rect 10275 35068 10287 35071
rect 10778 35068 10784 35080
rect 10275 35040 10784 35068
rect 10275 35037 10287 35040
rect 10229 35031 10287 35037
rect 10778 35028 10784 35040
rect 10836 35028 10842 35080
rect 2700 35000 2728 35028
rect 2332 34972 2728 35000
rect 2332 34932 2360 34972
rect 7374 34960 7380 35012
rect 7432 35000 7438 35012
rect 8202 35000 8208 35012
rect 7432 34972 8208 35000
rect 7432 34960 7438 34972
rect 8202 34960 8208 34972
rect 8260 34960 8266 35012
rect 8389 35003 8447 35009
rect 8389 34969 8401 35003
rect 8435 35000 8447 35003
rect 8478 35000 8484 35012
rect 8435 34972 8484 35000
rect 8435 34969 8447 34972
rect 8389 34963 8447 34969
rect 8478 34960 8484 34972
rect 8536 35000 8542 35012
rect 9582 35000 9588 35012
rect 8536 34972 9588 35000
rect 8536 34960 8542 34972
rect 9582 34960 9588 34972
rect 9640 34960 9646 35012
rect 10888 35000 10916 35099
rect 11606 35096 11612 35108
rect 11664 35096 11670 35148
rect 13078 35136 13084 35148
rect 13039 35108 13084 35136
rect 13078 35096 13084 35108
rect 13136 35096 13142 35148
rect 14826 35096 14832 35148
rect 14884 35136 14890 35148
rect 15565 35139 15623 35145
rect 15565 35136 15577 35139
rect 14884 35108 15577 35136
rect 14884 35096 14890 35108
rect 15565 35105 15577 35108
rect 15611 35105 15623 35139
rect 18046 35136 18052 35148
rect 18007 35108 18052 35136
rect 15565 35099 15623 35105
rect 18046 35096 18052 35108
rect 18104 35096 18110 35148
rect 22373 35139 22431 35145
rect 22373 35105 22385 35139
rect 22419 35105 22431 35139
rect 22373 35099 22431 35105
rect 22557 35139 22615 35145
rect 22557 35105 22569 35139
rect 22603 35136 22615 35139
rect 22646 35136 22652 35148
rect 22603 35108 22652 35136
rect 22603 35105 22615 35108
rect 22557 35099 22615 35105
rect 12805 35071 12863 35077
rect 12805 35037 12817 35071
rect 12851 35068 12863 35071
rect 13170 35068 13176 35080
rect 12851 35040 13176 35068
rect 12851 35037 12863 35040
rect 12805 35031 12863 35037
rect 13170 35028 13176 35040
rect 13228 35028 13234 35080
rect 15289 35071 15347 35077
rect 15289 35037 15301 35071
rect 15335 35068 15347 35071
rect 15746 35068 15752 35080
rect 15335 35040 15752 35068
rect 15335 35037 15347 35040
rect 15289 35031 15347 35037
rect 15746 35028 15752 35040
rect 15804 35068 15810 35080
rect 17773 35071 17831 35077
rect 17773 35068 17785 35071
rect 15804 35040 17785 35068
rect 15804 35028 15810 35040
rect 17773 35037 17785 35040
rect 17819 35037 17831 35071
rect 17773 35031 17831 35037
rect 20898 35028 20904 35080
rect 20956 35068 20962 35080
rect 21545 35071 21603 35077
rect 21545 35068 21557 35071
rect 20956 35040 21557 35068
rect 20956 35028 20962 35040
rect 21545 35037 21557 35040
rect 21591 35037 21603 35071
rect 21545 35031 21603 35037
rect 22094 35028 22100 35080
rect 22152 35068 22158 35080
rect 22152 35040 22197 35068
rect 22152 35028 22158 35040
rect 10796 34972 10916 35000
rect 1412 34904 2360 34932
rect 2774 34892 2780 34944
rect 2832 34932 2838 34944
rect 4157 34935 4215 34941
rect 2832 34904 2877 34932
rect 2832 34892 2838 34904
rect 4157 34901 4169 34935
rect 4203 34932 4215 34935
rect 5626 34932 5632 34944
rect 4203 34904 5632 34932
rect 4203 34901 4215 34904
rect 4157 34895 4215 34901
rect 5626 34892 5632 34904
rect 5684 34892 5690 34944
rect 5902 34892 5908 34944
rect 5960 34932 5966 34944
rect 9766 34932 9772 34944
rect 5960 34904 9772 34932
rect 5960 34892 5966 34904
rect 9766 34892 9772 34904
rect 9824 34932 9830 34944
rect 10796 34932 10824 34972
rect 22278 34960 22284 35012
rect 22336 35000 22342 35012
rect 22388 35000 22416 35099
rect 22646 35096 22652 35108
rect 22704 35096 22710 35148
rect 23106 35136 23112 35148
rect 23019 35108 23112 35136
rect 23106 35096 23112 35108
rect 23164 35096 23170 35148
rect 23216 35145 23244 35176
rect 23201 35139 23259 35145
rect 23201 35105 23213 35139
rect 23247 35105 23259 35139
rect 23382 35136 23388 35148
rect 23343 35108 23388 35136
rect 23201 35099 23259 35105
rect 23382 35096 23388 35108
rect 23440 35096 23446 35148
rect 23492 35136 23520 35176
rect 23845 35173 23857 35207
rect 23891 35204 23903 35207
rect 23891 35176 25544 35204
rect 23891 35173 23903 35176
rect 23845 35167 23903 35173
rect 23934 35136 23940 35148
rect 23492 35108 23940 35136
rect 23934 35096 23940 35108
rect 23992 35136 23998 35148
rect 24305 35139 24363 35145
rect 24305 35136 24317 35139
rect 23992 35108 24317 35136
rect 23992 35096 23998 35108
rect 24305 35105 24317 35108
rect 24351 35105 24363 35139
rect 24762 35136 24768 35148
rect 24723 35108 24768 35136
rect 24305 35099 24363 35105
rect 24762 35096 24768 35108
rect 24820 35096 24826 35148
rect 25516 35145 25544 35176
rect 26344 35145 26372 35244
rect 26436 35244 35992 35272
rect 25501 35139 25559 35145
rect 24872 35108 25452 35136
rect 23124 35068 23152 35096
rect 24780 35068 24808 35096
rect 23124 35040 24808 35068
rect 24872 35000 24900 35108
rect 25041 35071 25099 35077
rect 25041 35037 25053 35071
rect 25087 35037 25099 35071
rect 25424 35068 25452 35108
rect 25501 35105 25513 35139
rect 25547 35105 25559 35139
rect 25501 35099 25559 35105
rect 26329 35139 26387 35145
rect 26329 35105 26341 35139
rect 26375 35105 26387 35139
rect 26329 35099 26387 35105
rect 26436 35068 26464 35244
rect 35986 35232 35992 35244
rect 36044 35232 36050 35284
rect 30650 35164 30656 35216
rect 30708 35204 30714 35216
rect 34425 35207 34483 35213
rect 30708 35176 30880 35204
rect 30708 35164 30714 35176
rect 26786 35136 26792 35148
rect 26747 35108 26792 35136
rect 26786 35096 26792 35108
rect 26844 35096 26850 35148
rect 27062 35136 27068 35148
rect 27023 35108 27068 35136
rect 27062 35096 27068 35108
rect 27120 35096 27126 35148
rect 27246 35136 27252 35148
rect 27207 35108 27252 35136
rect 27246 35096 27252 35108
rect 27304 35136 27310 35148
rect 27522 35136 27528 35148
rect 27304 35108 27528 35136
rect 27304 35096 27310 35108
rect 27522 35096 27528 35108
rect 27580 35096 27586 35148
rect 29730 35136 29736 35148
rect 28644 35108 29736 35136
rect 26602 35068 26608 35080
rect 25424 35040 26464 35068
rect 26563 35040 26608 35068
rect 25041 35031 25099 35037
rect 22336 34972 24900 35000
rect 25056 35000 25084 35031
rect 26602 35028 26608 35040
rect 26660 35028 26666 35080
rect 28644 35077 28672 35108
rect 29730 35096 29736 35108
rect 29788 35096 29794 35148
rect 30742 35136 30748 35148
rect 30703 35108 30748 35136
rect 30742 35096 30748 35108
rect 30800 35096 30806 35148
rect 30852 35145 30880 35176
rect 34425 35173 34437 35207
rect 34471 35204 34483 35207
rect 34514 35204 34520 35216
rect 34471 35176 34520 35204
rect 34471 35173 34483 35176
rect 34425 35167 34483 35173
rect 34514 35164 34520 35176
rect 34572 35164 34578 35216
rect 30837 35139 30895 35145
rect 30837 35105 30849 35139
rect 30883 35136 30895 35139
rect 32030 35136 32036 35148
rect 30883 35108 32036 35136
rect 30883 35105 30895 35108
rect 30837 35099 30895 35105
rect 32030 35096 32036 35108
rect 32088 35096 32094 35148
rect 32122 35096 32128 35148
rect 32180 35136 32186 35148
rect 32769 35139 32827 35145
rect 32769 35136 32781 35139
rect 32180 35108 32781 35136
rect 32180 35096 32186 35108
rect 32769 35105 32781 35108
rect 32815 35105 32827 35139
rect 32769 35099 32827 35105
rect 33045 35139 33103 35145
rect 33045 35105 33057 35139
rect 33091 35136 33103 35139
rect 33502 35136 33508 35148
rect 33091 35108 33508 35136
rect 33091 35105 33103 35108
rect 33045 35099 33103 35105
rect 33502 35096 33508 35108
rect 33560 35096 33566 35148
rect 28629 35071 28687 35077
rect 28629 35037 28641 35071
rect 28675 35037 28687 35071
rect 28629 35031 28687 35037
rect 28905 35071 28963 35077
rect 28905 35037 28917 35071
rect 28951 35068 28963 35071
rect 31294 35068 31300 35080
rect 28951 35040 30328 35068
rect 31255 35040 31300 35068
rect 28951 35037 28963 35040
rect 28905 35031 28963 35037
rect 27706 35000 27712 35012
rect 25056 34972 27712 35000
rect 22336 34960 22342 34972
rect 27706 34960 27712 34972
rect 27764 34960 27770 35012
rect 9824 34904 10824 34932
rect 9824 34892 9830 34904
rect 13998 34892 14004 34944
rect 14056 34932 14062 34944
rect 14185 34935 14243 34941
rect 14185 34932 14197 34935
rect 14056 34904 14197 34932
rect 14056 34892 14062 34904
rect 14185 34901 14197 34904
rect 14231 34932 14243 34935
rect 14274 34932 14280 34944
rect 14231 34904 14280 34932
rect 14231 34901 14243 34904
rect 14185 34895 14243 34901
rect 14274 34892 14280 34904
rect 14332 34892 14338 34944
rect 16853 34935 16911 34941
rect 16853 34901 16865 34935
rect 16899 34932 16911 34935
rect 17034 34932 17040 34944
rect 16899 34904 17040 34932
rect 16899 34901 16911 34904
rect 16853 34895 16911 34901
rect 17034 34892 17040 34904
rect 17092 34892 17098 34944
rect 18966 34892 18972 34944
rect 19024 34932 19030 34944
rect 19153 34935 19211 34941
rect 19153 34932 19165 34935
rect 19024 34904 19165 34932
rect 19024 34892 19030 34904
rect 19153 34901 19165 34904
rect 19199 34901 19211 34935
rect 19153 34895 19211 34901
rect 24486 34892 24492 34944
rect 24544 34932 24550 34944
rect 25593 34935 25651 34941
rect 25593 34932 25605 34935
rect 24544 34904 25605 34932
rect 24544 34892 24550 34904
rect 25593 34901 25605 34904
rect 25639 34901 25651 34935
rect 25593 34895 25651 34901
rect 26145 34935 26203 34941
rect 26145 34901 26157 34935
rect 26191 34932 26203 34935
rect 26326 34932 26332 34944
rect 26191 34904 26332 34932
rect 26191 34901 26203 34904
rect 26145 34895 26203 34901
rect 26326 34892 26332 34904
rect 26384 34932 26390 34944
rect 28644 34932 28672 35031
rect 26384 34904 28672 34932
rect 26384 34892 26390 34904
rect 29546 34892 29552 34944
rect 29604 34932 29610 34944
rect 30009 34935 30067 34941
rect 30009 34932 30021 34935
rect 29604 34904 30021 34932
rect 29604 34892 29610 34904
rect 30009 34901 30021 34904
rect 30055 34901 30067 34935
rect 30300 34932 30328 35040
rect 31294 35028 31300 35040
rect 31352 35028 31358 35080
rect 35618 34932 35624 34944
rect 30300 34904 35624 34932
rect 30009 34895 30067 34901
rect 35618 34892 35624 34904
rect 35676 34892 35682 34944
rect 1104 34842 39836 34864
rect 1104 34790 4246 34842
rect 4298 34790 4310 34842
rect 4362 34790 4374 34842
rect 4426 34790 4438 34842
rect 4490 34790 34966 34842
rect 35018 34790 35030 34842
rect 35082 34790 35094 34842
rect 35146 34790 35158 34842
rect 35210 34790 39836 34842
rect 1104 34768 39836 34790
rect 2130 34728 2136 34740
rect 2091 34700 2136 34728
rect 2130 34688 2136 34700
rect 2188 34688 2194 34740
rect 3786 34688 3792 34740
rect 3844 34728 3850 34740
rect 3844 34700 7052 34728
rect 3844 34688 3850 34700
rect 5718 34620 5724 34672
rect 5776 34660 5782 34672
rect 5813 34663 5871 34669
rect 5813 34660 5825 34663
rect 5776 34632 5825 34660
rect 5776 34620 5782 34632
rect 5813 34629 5825 34632
rect 5859 34629 5871 34663
rect 5813 34623 5871 34629
rect 2682 34552 2688 34604
rect 2740 34592 2746 34604
rect 2869 34595 2927 34601
rect 2869 34592 2881 34595
rect 2740 34564 2881 34592
rect 2740 34552 2746 34564
rect 2869 34561 2881 34564
rect 2915 34561 2927 34595
rect 2869 34555 2927 34561
rect 5169 34595 5227 34601
rect 5169 34561 5181 34595
rect 5215 34592 5227 34595
rect 5215 34564 6776 34592
rect 5215 34561 5227 34564
rect 5169 34555 5227 34561
rect 6748 34536 6776 34564
rect 1762 34524 1768 34536
rect 1723 34496 1768 34524
rect 1762 34484 1768 34496
rect 1820 34484 1826 34536
rect 1946 34524 1952 34536
rect 1907 34496 1952 34524
rect 1946 34484 1952 34496
rect 2004 34484 2010 34536
rect 3145 34527 3203 34533
rect 3145 34493 3157 34527
rect 3191 34524 3203 34527
rect 4154 34524 4160 34536
rect 3191 34496 4160 34524
rect 3191 34493 3203 34496
rect 3145 34487 3203 34493
rect 4154 34484 4160 34496
rect 4212 34484 4218 34536
rect 5350 34524 5356 34536
rect 5311 34496 5356 34524
rect 5350 34484 5356 34496
rect 5408 34484 5414 34536
rect 5902 34524 5908 34536
rect 5863 34496 5908 34524
rect 5902 34484 5908 34496
rect 5960 34484 5966 34536
rect 6730 34484 6736 34536
rect 6788 34524 6794 34536
rect 6917 34527 6975 34533
rect 6917 34524 6929 34527
rect 6788 34496 6929 34524
rect 6788 34484 6794 34496
rect 6917 34493 6929 34496
rect 6963 34493 6975 34527
rect 7024 34524 7052 34700
rect 8110 34688 8116 34740
rect 8168 34728 8174 34740
rect 11425 34731 11483 34737
rect 8168 34700 9076 34728
rect 8168 34688 8174 34700
rect 8754 34660 8760 34672
rect 8312 34632 8760 34660
rect 8312 34592 8340 34632
rect 8754 34620 8760 34632
rect 8812 34620 8818 34672
rect 9048 34601 9076 34700
rect 11425 34697 11437 34731
rect 11471 34728 11483 34731
rect 11606 34728 11612 34740
rect 11471 34700 11612 34728
rect 11471 34697 11483 34700
rect 11425 34691 11483 34697
rect 11606 34688 11612 34700
rect 11664 34688 11670 34740
rect 15010 34728 15016 34740
rect 12452 34700 15016 34728
rect 12452 34669 12480 34700
rect 15010 34688 15016 34700
rect 15068 34728 15074 34740
rect 16209 34731 16267 34737
rect 16209 34728 16221 34731
rect 15068 34700 16221 34728
rect 15068 34688 15074 34700
rect 16209 34697 16221 34700
rect 16255 34697 16267 34731
rect 17218 34728 17224 34740
rect 17179 34700 17224 34728
rect 16209 34691 16267 34697
rect 17218 34688 17224 34700
rect 17276 34688 17282 34740
rect 22094 34688 22100 34740
rect 22152 34728 22158 34740
rect 23293 34731 23351 34737
rect 22152 34700 22197 34728
rect 22152 34688 22158 34700
rect 23293 34697 23305 34731
rect 23339 34728 23351 34731
rect 24670 34728 24676 34740
rect 23339 34700 24676 34728
rect 23339 34697 23351 34700
rect 23293 34691 23351 34697
rect 24670 34688 24676 34700
rect 24728 34688 24734 34740
rect 32030 34688 32036 34740
rect 32088 34728 32094 34740
rect 32953 34731 33011 34737
rect 32088 34700 32352 34728
rect 32088 34688 32094 34700
rect 12437 34663 12495 34669
rect 12437 34629 12449 34663
rect 12483 34629 12495 34663
rect 12437 34623 12495 34629
rect 23382 34620 23388 34672
rect 23440 34660 23446 34672
rect 32324 34660 32352 34700
rect 32953 34697 32965 34731
rect 32999 34728 33011 34731
rect 33042 34728 33048 34740
rect 32999 34700 33048 34728
rect 32999 34697 33011 34700
rect 32953 34691 33011 34697
rect 33042 34688 33048 34700
rect 33100 34688 33106 34740
rect 36170 34660 36176 34672
rect 23440 34632 24256 34660
rect 32324 34632 36176 34660
rect 23440 34620 23446 34632
rect 8220 34564 8340 34592
rect 9033 34595 9091 34601
rect 7374 34524 7380 34536
rect 7024 34496 7380 34524
rect 6917 34487 6975 34493
rect 7374 34484 7380 34496
rect 7432 34484 7438 34536
rect 8220 34533 8248 34564
rect 9033 34561 9045 34595
rect 9079 34561 9091 34595
rect 9033 34555 9091 34561
rect 9582 34552 9588 34604
rect 9640 34592 9646 34604
rect 12805 34595 12863 34601
rect 9640 34564 10824 34592
rect 9640 34552 9646 34564
rect 8205 34527 8263 34533
rect 8205 34493 8217 34527
rect 8251 34493 8263 34527
rect 8938 34524 8944 34536
rect 8205 34487 8263 34493
rect 8312 34496 8944 34524
rect 1857 34459 1915 34465
rect 1857 34425 1869 34459
rect 1903 34425 1915 34459
rect 1857 34419 1915 34425
rect 4525 34459 4583 34465
rect 4525 34425 4537 34459
rect 4571 34456 4583 34459
rect 4706 34456 4712 34468
rect 4571 34428 4712 34456
rect 4571 34425 4583 34428
rect 4525 34419 4583 34425
rect 1872 34388 1900 34419
rect 4706 34416 4712 34428
rect 4764 34416 4770 34468
rect 7653 34459 7711 34465
rect 7653 34425 7665 34459
rect 7699 34456 7711 34459
rect 8312 34456 8340 34496
rect 8938 34484 8944 34496
rect 8996 34484 9002 34536
rect 9953 34527 10011 34533
rect 9953 34524 9965 34527
rect 9140 34496 9965 34524
rect 7699 34428 8340 34456
rect 7699 34425 7711 34428
rect 7653 34419 7711 34425
rect 8386 34416 8392 34468
rect 8444 34456 8450 34468
rect 9140 34456 9168 34496
rect 9953 34493 9965 34496
rect 9999 34493 10011 34527
rect 10226 34524 10232 34536
rect 10187 34496 10232 34524
rect 9953 34487 10011 34493
rect 10226 34484 10232 34496
rect 10284 34484 10290 34536
rect 10796 34533 10824 34564
rect 12805 34561 12817 34595
rect 12851 34592 12863 34595
rect 13906 34592 13912 34604
rect 12851 34564 13912 34592
rect 12851 34561 12863 34564
rect 12805 34555 12863 34561
rect 13906 34552 13912 34564
rect 13964 34552 13970 34604
rect 14829 34595 14887 34601
rect 14829 34561 14841 34595
rect 14875 34592 14887 34595
rect 15286 34592 15292 34604
rect 14875 34564 15292 34592
rect 14875 34561 14887 34564
rect 14829 34555 14887 34561
rect 15286 34552 15292 34564
rect 15344 34552 15350 34604
rect 16945 34595 17003 34601
rect 16945 34561 16957 34595
rect 16991 34592 17003 34595
rect 18877 34595 18935 34601
rect 18877 34592 18889 34595
rect 16991 34564 18889 34592
rect 16991 34561 17003 34564
rect 16945 34555 17003 34561
rect 18877 34561 18889 34564
rect 18923 34592 18935 34595
rect 20346 34592 20352 34604
rect 18923 34564 20352 34592
rect 18923 34561 18935 34564
rect 18877 34555 18935 34561
rect 20346 34552 20352 34564
rect 20404 34552 20410 34604
rect 21634 34552 21640 34604
rect 21692 34592 21698 34604
rect 24228 34592 24256 34632
rect 36170 34620 36176 34632
rect 36228 34620 36234 34672
rect 24486 34592 24492 34604
rect 21692 34564 23520 34592
rect 24228 34564 24348 34592
rect 24447 34564 24492 34592
rect 21692 34552 21698 34564
rect 10689 34527 10747 34533
rect 10689 34493 10701 34527
rect 10735 34493 10747 34527
rect 10689 34487 10747 34493
rect 10781 34527 10839 34533
rect 10781 34493 10793 34527
rect 10827 34493 10839 34527
rect 10781 34487 10839 34493
rect 8444 34428 9168 34456
rect 8444 34416 8450 34428
rect 5718 34388 5724 34400
rect 1872 34360 5724 34388
rect 5718 34348 5724 34360
rect 5776 34348 5782 34400
rect 8297 34391 8355 34397
rect 8297 34357 8309 34391
rect 8343 34388 8355 34391
rect 8846 34388 8852 34400
rect 8343 34360 8852 34388
rect 8343 34357 8355 34360
rect 8297 34351 8355 34357
rect 8846 34348 8852 34360
rect 8904 34348 8910 34400
rect 9769 34391 9827 34397
rect 9769 34357 9781 34391
rect 9815 34388 9827 34391
rect 9858 34388 9864 34400
rect 9815 34360 9864 34388
rect 9815 34357 9827 34360
rect 9769 34351 9827 34357
rect 9858 34348 9864 34360
rect 9916 34348 9922 34400
rect 10502 34348 10508 34400
rect 10560 34388 10566 34400
rect 10704 34388 10732 34487
rect 11054 34484 11060 34536
rect 11112 34524 11118 34536
rect 11333 34527 11391 34533
rect 11333 34524 11345 34527
rect 11112 34496 11345 34524
rect 11112 34484 11118 34496
rect 11333 34493 11345 34496
rect 11379 34493 11391 34527
rect 11333 34487 11391 34493
rect 12618 34484 12624 34536
rect 12676 34524 12682 34536
rect 12897 34527 12955 34533
rect 12897 34524 12909 34527
rect 12676 34496 12909 34524
rect 12676 34484 12682 34496
rect 12897 34493 12909 34496
rect 12943 34493 12955 34527
rect 13357 34527 13415 34533
rect 13357 34524 13369 34527
rect 12897 34487 12955 34493
rect 13004 34496 13369 34524
rect 11514 34416 11520 34468
rect 11572 34456 11578 34468
rect 13004 34456 13032 34496
rect 13357 34493 13369 34496
rect 13403 34493 13415 34527
rect 13357 34487 13415 34493
rect 13817 34527 13875 34533
rect 13817 34493 13829 34527
rect 13863 34524 13875 34527
rect 13998 34524 14004 34536
rect 13863 34496 14004 34524
rect 13863 34493 13875 34496
rect 13817 34487 13875 34493
rect 13998 34484 14004 34496
rect 14056 34484 14062 34536
rect 14369 34527 14427 34533
rect 14369 34493 14381 34527
rect 14415 34524 14427 34527
rect 14458 34524 14464 34536
rect 14415 34496 14464 34524
rect 14415 34493 14427 34496
rect 14369 34487 14427 34493
rect 14458 34484 14464 34496
rect 14516 34484 14522 34536
rect 15102 34524 15108 34536
rect 15063 34496 15108 34524
rect 15102 34484 15108 34496
rect 15160 34484 15166 34536
rect 17034 34484 17040 34536
rect 17092 34524 17098 34536
rect 17092 34496 17137 34524
rect 17092 34484 17098 34496
rect 18966 34484 18972 34536
rect 19024 34524 19030 34536
rect 19886 34524 19892 34536
rect 19024 34496 19069 34524
rect 19847 34496 19892 34524
rect 19024 34484 19030 34496
rect 19886 34484 19892 34496
rect 19944 34484 19950 34536
rect 20162 34524 20168 34536
rect 20123 34496 20168 34524
rect 20162 34484 20168 34496
rect 20220 34484 20226 34536
rect 22278 34524 22284 34536
rect 22239 34496 22284 34524
rect 22278 34484 22284 34496
rect 22336 34484 22342 34536
rect 22738 34524 22744 34536
rect 22699 34496 22744 34524
rect 22738 34484 22744 34496
rect 22796 34484 22802 34536
rect 23492 34533 23520 34564
rect 23477 34527 23535 34533
rect 23477 34493 23489 34527
rect 23523 34493 23535 34527
rect 23477 34487 23535 34493
rect 24118 34484 24124 34536
rect 24176 34524 24182 34536
rect 24213 34527 24271 34533
rect 24213 34524 24225 34527
rect 24176 34496 24225 34524
rect 24176 34484 24182 34496
rect 24213 34493 24225 34496
rect 24259 34493 24271 34527
rect 24320 34524 24348 34564
rect 24486 34552 24492 34564
rect 24544 34552 24550 34604
rect 25593 34595 25651 34601
rect 25593 34561 25605 34595
rect 25639 34592 25651 34595
rect 27246 34592 27252 34604
rect 25639 34564 27252 34592
rect 25639 34561 25651 34564
rect 25593 34555 25651 34561
rect 25608 34524 25636 34555
rect 27246 34552 27252 34564
rect 27304 34552 27310 34604
rect 29546 34592 29552 34604
rect 29507 34564 29552 34592
rect 29546 34552 29552 34564
rect 29604 34552 29610 34604
rect 31294 34552 31300 34604
rect 31352 34592 31358 34604
rect 31665 34595 31723 34601
rect 31665 34592 31677 34595
rect 31352 34564 31677 34592
rect 31352 34552 31358 34564
rect 31665 34561 31677 34564
rect 31711 34561 31723 34595
rect 34882 34592 34888 34604
rect 34843 34564 34888 34592
rect 31665 34555 31723 34561
rect 34882 34552 34888 34564
rect 34940 34552 34946 34604
rect 24320 34496 25636 34524
rect 24213 34487 24271 34493
rect 26326 34484 26332 34536
rect 26384 34524 26390 34536
rect 26789 34527 26847 34533
rect 26789 34524 26801 34527
rect 26384 34496 26801 34524
rect 26384 34484 26390 34496
rect 26789 34493 26801 34496
rect 26835 34493 26847 34527
rect 26789 34487 26847 34493
rect 27065 34527 27123 34533
rect 27065 34493 27077 34527
rect 27111 34524 27123 34527
rect 28166 34524 28172 34536
rect 27111 34496 28172 34524
rect 27111 34493 27123 34496
rect 27065 34487 27123 34493
rect 28166 34484 28172 34496
rect 28224 34484 28230 34536
rect 29273 34527 29331 34533
rect 29273 34493 29285 34527
rect 29319 34524 29331 34527
rect 29362 34524 29368 34536
rect 29319 34496 29368 34524
rect 29319 34493 29331 34496
rect 29273 34487 29331 34493
rect 29362 34484 29368 34496
rect 29420 34484 29426 34536
rect 31389 34527 31447 34533
rect 31389 34524 31401 34527
rect 31220 34496 31401 34524
rect 19426 34456 19432 34468
rect 11572 34428 13032 34456
rect 19387 34428 19432 34456
rect 11572 34416 11578 34428
rect 19426 34416 19432 34428
rect 19484 34416 19490 34468
rect 21545 34459 21603 34465
rect 21545 34425 21557 34459
rect 21591 34456 21603 34459
rect 21818 34456 21824 34468
rect 21591 34428 21824 34456
rect 21591 34425 21603 34428
rect 21545 34419 21603 34425
rect 21818 34416 21824 34428
rect 21876 34416 21882 34468
rect 12618 34388 12624 34400
rect 10560 34360 12624 34388
rect 10560 34348 10566 34360
rect 12618 34348 12624 34360
rect 12676 34348 12682 34400
rect 28350 34388 28356 34400
rect 28311 34360 28356 34388
rect 28350 34348 28356 34360
rect 28408 34348 28414 34400
rect 30650 34388 30656 34400
rect 30611 34360 30656 34388
rect 30650 34348 30656 34360
rect 30708 34348 30714 34400
rect 31220 34388 31248 34496
rect 31389 34493 31401 34496
rect 31435 34493 31447 34527
rect 33689 34527 33747 34533
rect 33689 34524 33701 34527
rect 31389 34487 31447 34493
rect 31496 34496 33701 34524
rect 31294 34416 31300 34468
rect 31352 34456 31358 34468
rect 31496 34456 31524 34496
rect 33689 34493 33701 34496
rect 33735 34493 33747 34527
rect 33689 34487 33747 34493
rect 33778 34484 33784 34536
rect 33836 34524 33842 34536
rect 34241 34527 34299 34533
rect 33836 34496 33881 34524
rect 33836 34484 33842 34496
rect 34241 34493 34253 34527
rect 34287 34524 34299 34527
rect 34790 34524 34796 34536
rect 34287 34496 34796 34524
rect 34287 34493 34299 34496
rect 34241 34487 34299 34493
rect 34790 34484 34796 34496
rect 34848 34484 34854 34536
rect 34974 34524 34980 34536
rect 34935 34496 34980 34524
rect 34974 34484 34980 34496
rect 35032 34484 35038 34536
rect 31352 34428 31524 34456
rect 31352 34416 31358 34428
rect 35250 34416 35256 34468
rect 35308 34456 35314 34468
rect 35437 34459 35495 34465
rect 35437 34456 35449 34459
rect 35308 34428 35449 34456
rect 35308 34416 35314 34428
rect 35437 34425 35449 34428
rect 35483 34425 35495 34459
rect 35437 34419 35495 34425
rect 32490 34388 32496 34400
rect 31220 34360 32496 34388
rect 32490 34348 32496 34360
rect 32548 34348 32554 34400
rect 1104 34298 39836 34320
rect 1104 34246 19606 34298
rect 19658 34246 19670 34298
rect 19722 34246 19734 34298
rect 19786 34246 19798 34298
rect 19850 34246 39836 34298
rect 1104 34224 39836 34246
rect 8294 34184 8300 34196
rect 8255 34156 8300 34184
rect 8294 34144 8300 34156
rect 8352 34144 8358 34196
rect 10045 34187 10103 34193
rect 10045 34153 10057 34187
rect 10091 34184 10103 34187
rect 11054 34184 11060 34196
rect 10091 34156 11060 34184
rect 10091 34153 10103 34156
rect 10045 34147 10103 34153
rect 11054 34144 11060 34156
rect 11112 34144 11118 34196
rect 14185 34187 14243 34193
rect 14185 34153 14197 34187
rect 14231 34184 14243 34187
rect 15102 34184 15108 34196
rect 14231 34156 15108 34184
rect 14231 34153 14243 34156
rect 14185 34147 14243 34153
rect 15102 34144 15108 34156
rect 15160 34144 15166 34196
rect 27246 34144 27252 34196
rect 27304 34184 27310 34196
rect 27304 34156 29040 34184
rect 27304 34144 27310 34156
rect 1762 34076 1768 34128
rect 1820 34116 1826 34128
rect 2041 34119 2099 34125
rect 2041 34116 2053 34119
rect 1820 34088 2053 34116
rect 1820 34076 1826 34088
rect 2041 34085 2053 34088
rect 2087 34085 2099 34119
rect 2774 34116 2780 34128
rect 2041 34079 2099 34085
rect 2608 34088 2780 34116
rect 2608 34057 2636 34088
rect 2774 34076 2780 34088
rect 2832 34076 2838 34128
rect 3050 34116 3056 34128
rect 2884 34088 3056 34116
rect 2884 34057 2912 34088
rect 3050 34076 3056 34088
rect 3108 34076 3114 34128
rect 4065 34119 4123 34125
rect 4065 34085 4077 34119
rect 4111 34116 4123 34119
rect 4154 34116 4160 34128
rect 4111 34088 4160 34116
rect 4111 34085 4123 34088
rect 4065 34079 4123 34085
rect 4154 34076 4160 34088
rect 4212 34076 4218 34128
rect 5626 34076 5632 34128
rect 5684 34116 5690 34128
rect 8110 34116 8116 34128
rect 5684 34088 6592 34116
rect 5684 34076 5690 34088
rect 2593 34051 2651 34057
rect 2593 34017 2605 34051
rect 2639 34017 2651 34051
rect 2593 34011 2651 34017
rect 2685 34051 2743 34057
rect 2685 34017 2697 34051
rect 2731 34048 2743 34051
rect 2869 34051 2927 34057
rect 2731 34020 2820 34048
rect 2731 34017 2743 34020
rect 2685 34011 2743 34017
rect 2792 33980 2820 34020
rect 2869 34017 2881 34051
rect 2915 34017 2927 34051
rect 3142 34048 3148 34060
rect 3103 34020 3148 34048
rect 2869 34011 2927 34017
rect 3142 34008 3148 34020
rect 3200 34008 3206 34060
rect 3326 34048 3332 34060
rect 3287 34020 3332 34048
rect 3326 34008 3332 34020
rect 3384 34008 3390 34060
rect 3694 34008 3700 34060
rect 3752 34048 3758 34060
rect 6564 34057 6592 34088
rect 7024 34088 8116 34116
rect 4893 34051 4951 34057
rect 4893 34048 4905 34051
rect 3752 34020 4905 34048
rect 3752 34008 3758 34020
rect 4893 34017 4905 34020
rect 4939 34017 4951 34051
rect 4893 34011 4951 34017
rect 5813 34051 5871 34057
rect 5813 34017 5825 34051
rect 5859 34048 5871 34051
rect 6457 34051 6515 34057
rect 5859 34020 6408 34048
rect 5859 34017 5871 34020
rect 5813 34011 5871 34017
rect 2958 33980 2964 33992
rect 2792 33952 2964 33980
rect 2958 33940 2964 33952
rect 3016 33940 3022 33992
rect 4614 33980 4620 33992
rect 4575 33952 4620 33980
rect 4614 33940 4620 33952
rect 4672 33940 4678 33992
rect 5074 33980 5080 33992
rect 5035 33952 5080 33980
rect 5074 33940 5080 33952
rect 5132 33940 5138 33992
rect 5902 33980 5908 33992
rect 5863 33952 5908 33980
rect 5902 33940 5908 33952
rect 5960 33940 5966 33992
rect 5629 33915 5687 33921
rect 5629 33881 5641 33915
rect 5675 33912 5687 33915
rect 6086 33912 6092 33924
rect 5675 33884 6092 33912
rect 5675 33881 5687 33884
rect 5629 33875 5687 33881
rect 6086 33872 6092 33884
rect 6144 33872 6150 33924
rect 6380 33912 6408 34020
rect 6457 34017 6469 34051
rect 6503 34017 6515 34051
rect 6457 34011 6515 34017
rect 6549 34051 6607 34057
rect 6549 34017 6561 34051
rect 6595 34017 6607 34051
rect 6549 34011 6607 34017
rect 6472 33980 6500 34011
rect 6638 34008 6644 34060
rect 6696 34048 6702 34060
rect 6733 34051 6791 34057
rect 6733 34048 6745 34051
rect 6696 34020 6745 34048
rect 6696 34008 6702 34020
rect 6733 34017 6745 34020
rect 6779 34017 6791 34051
rect 6733 34011 6791 34017
rect 6914 34008 6920 34060
rect 6972 34048 6978 34060
rect 7024 34057 7052 34088
rect 8110 34076 8116 34088
rect 8168 34076 8174 34128
rect 8570 34076 8576 34128
rect 8628 34116 8634 34128
rect 9030 34116 9036 34128
rect 8628 34088 9036 34116
rect 8628 34076 8634 34088
rect 9030 34076 9036 34088
rect 9088 34116 9094 34128
rect 9582 34116 9588 34128
rect 9088 34088 9588 34116
rect 9088 34076 9094 34088
rect 9582 34076 9588 34088
rect 9640 34116 9646 34128
rect 9953 34119 10011 34125
rect 9953 34116 9965 34119
rect 9640 34088 9965 34116
rect 9640 34076 9646 34088
rect 9953 34085 9965 34088
rect 9999 34085 10011 34119
rect 9953 34079 10011 34085
rect 10137 34119 10195 34125
rect 10137 34085 10149 34119
rect 10183 34116 10195 34119
rect 10226 34116 10232 34128
rect 10183 34088 10232 34116
rect 10183 34085 10195 34088
rect 10137 34079 10195 34085
rect 10226 34076 10232 34088
rect 10284 34116 10290 34128
rect 10962 34116 10968 34128
rect 10284 34088 10968 34116
rect 10284 34076 10290 34088
rect 10962 34076 10968 34088
rect 11020 34076 11026 34128
rect 12618 34116 12624 34128
rect 12579 34088 12624 34116
rect 12618 34076 12624 34088
rect 12676 34076 12682 34128
rect 27062 34116 27068 34128
rect 26804 34088 27068 34116
rect 7009 34051 7067 34057
rect 7009 34048 7021 34051
rect 6972 34020 7021 34048
rect 6972 34008 6978 34020
rect 7009 34017 7021 34020
rect 7055 34017 7067 34051
rect 7190 34048 7196 34060
rect 7151 34020 7196 34048
rect 7009 34011 7067 34017
rect 7190 34008 7196 34020
rect 7248 34008 7254 34060
rect 8202 34048 8208 34060
rect 8163 34020 8208 34048
rect 8202 34008 8208 34020
rect 8260 34008 8266 34060
rect 8478 34048 8484 34060
rect 8439 34020 8484 34048
rect 8478 34008 8484 34020
rect 8536 34008 8542 34060
rect 8846 34048 8852 34060
rect 8807 34020 8852 34048
rect 8846 34008 8852 34020
rect 8904 34008 8910 34060
rect 10505 34051 10563 34057
rect 10505 34017 10517 34051
rect 10551 34048 10563 34051
rect 11514 34048 11520 34060
rect 10551 34020 11520 34048
rect 10551 34017 10563 34020
rect 10505 34011 10563 34017
rect 11514 34008 11520 34020
rect 11572 34008 11578 34060
rect 13354 34048 13360 34060
rect 13315 34020 13360 34048
rect 13354 34008 13360 34020
rect 13412 34008 13418 34060
rect 13906 34048 13912 34060
rect 13867 34020 13912 34048
rect 13906 34008 13912 34020
rect 13964 34008 13970 34060
rect 16853 34051 16911 34057
rect 16853 34017 16865 34051
rect 16899 34048 16911 34051
rect 17218 34048 17224 34060
rect 16899 34020 17224 34048
rect 16899 34017 16911 34020
rect 16853 34011 16911 34017
rect 17218 34008 17224 34020
rect 17276 34008 17282 34060
rect 18969 34051 19027 34057
rect 18969 34017 18981 34051
rect 19015 34048 19027 34051
rect 19426 34048 19432 34060
rect 19015 34020 19432 34048
rect 19015 34017 19027 34020
rect 18969 34011 19027 34017
rect 19426 34008 19432 34020
rect 19484 34008 19490 34060
rect 20990 34008 20996 34060
rect 21048 34048 21054 34060
rect 21913 34051 21971 34057
rect 21913 34048 21925 34051
rect 21048 34020 21925 34048
rect 21048 34008 21054 34020
rect 21913 34017 21925 34020
rect 21959 34017 21971 34051
rect 24210 34048 24216 34060
rect 24171 34020 24216 34048
rect 21913 34011 21971 34017
rect 24210 34008 24216 34020
rect 24268 34008 24274 34060
rect 25222 34048 25228 34060
rect 25183 34020 25228 34048
rect 25222 34008 25228 34020
rect 25280 34008 25286 34060
rect 26804 34057 26832 34088
rect 27062 34076 27068 34088
rect 27120 34116 27126 34128
rect 28350 34116 28356 34128
rect 27120 34088 28356 34116
rect 27120 34076 27126 34088
rect 28350 34076 28356 34088
rect 28408 34116 28414 34128
rect 28905 34119 28963 34125
rect 28905 34116 28917 34119
rect 28408 34088 28917 34116
rect 28408 34076 28414 34088
rect 28905 34085 28917 34088
rect 28951 34085 28963 34119
rect 28905 34079 28963 34085
rect 26789 34051 26847 34057
rect 26789 34017 26801 34051
rect 26835 34017 26847 34051
rect 27246 34048 27252 34060
rect 27207 34020 27252 34048
rect 26789 34011 26847 34017
rect 27246 34008 27252 34020
rect 27304 34008 27310 34060
rect 27706 34048 27712 34060
rect 27667 34020 27712 34048
rect 27706 34008 27712 34020
rect 27764 34008 27770 34060
rect 27893 34051 27951 34057
rect 27893 34017 27905 34051
rect 27939 34017 27951 34051
rect 27893 34011 27951 34017
rect 27985 34051 28043 34057
rect 27985 34017 27997 34051
rect 28031 34017 28043 34051
rect 29012 34048 29040 34156
rect 31386 34144 31392 34196
rect 31444 34184 31450 34196
rect 31481 34187 31539 34193
rect 31481 34184 31493 34187
rect 31444 34156 31493 34184
rect 31444 34144 31450 34156
rect 31481 34153 31493 34156
rect 31527 34153 31539 34187
rect 34882 34184 34888 34196
rect 31481 34147 31539 34153
rect 32140 34156 34888 34184
rect 29089 34051 29147 34057
rect 29089 34048 29101 34051
rect 29012 34020 29101 34048
rect 27985 34011 28043 34017
rect 29089 34017 29101 34020
rect 29135 34017 29147 34051
rect 29089 34011 29147 34017
rect 7098 33980 7104 33992
rect 6472 33952 7104 33980
rect 7098 33940 7104 33952
rect 7156 33940 7162 33992
rect 7834 33940 7840 33992
rect 7892 33980 7898 33992
rect 9769 33983 9827 33989
rect 9769 33980 9781 33983
rect 7892 33952 9781 33980
rect 7892 33940 7898 33952
rect 9769 33949 9781 33952
rect 9815 33980 9827 33983
rect 10594 33980 10600 33992
rect 9815 33952 10600 33980
rect 9815 33949 9827 33952
rect 9769 33943 9827 33949
rect 10594 33940 10600 33952
rect 10652 33940 10658 33992
rect 10965 33983 11023 33989
rect 10965 33949 10977 33983
rect 11011 33949 11023 33983
rect 11238 33980 11244 33992
rect 11199 33952 11244 33980
rect 10965 33943 11023 33949
rect 8386 33912 8392 33924
rect 6380 33884 8392 33912
rect 8386 33872 8392 33884
rect 8444 33872 8450 33924
rect 9858 33872 9864 33924
rect 9916 33912 9922 33924
rect 10042 33912 10048 33924
rect 9916 33884 10048 33912
rect 9916 33872 9922 33884
rect 10042 33872 10048 33884
rect 10100 33912 10106 33924
rect 10980 33912 11008 33943
rect 11238 33940 11244 33952
rect 11296 33940 11302 33992
rect 13814 33980 13820 33992
rect 13775 33952 13820 33980
rect 13814 33940 13820 33952
rect 13872 33940 13878 33992
rect 15930 33940 15936 33992
rect 15988 33980 15994 33992
rect 16577 33983 16635 33989
rect 16577 33980 16589 33983
rect 15988 33952 16589 33980
rect 15988 33940 15994 33952
rect 16577 33949 16589 33952
rect 16623 33980 16635 33983
rect 18693 33983 18751 33989
rect 18693 33980 18705 33983
rect 16623 33952 18705 33980
rect 16623 33949 16635 33952
rect 16577 33943 16635 33949
rect 18693 33949 18705 33952
rect 18739 33949 18751 33983
rect 18693 33943 18751 33949
rect 19886 33940 19892 33992
rect 19944 33980 19950 33992
rect 22005 33983 22063 33989
rect 22005 33980 22017 33983
rect 19944 33952 22017 33980
rect 19944 33940 19950 33952
rect 22005 33949 22017 33952
rect 22051 33949 22063 33983
rect 22278 33980 22284 33992
rect 22239 33952 22284 33980
rect 22005 33943 22063 33949
rect 22278 33940 22284 33952
rect 22336 33940 22342 33992
rect 24118 33980 24124 33992
rect 24079 33952 24124 33980
rect 24118 33940 24124 33952
rect 24176 33940 24182 33992
rect 25130 33980 25136 33992
rect 25091 33952 25136 33980
rect 25130 33940 25136 33952
rect 25188 33940 25194 33992
rect 27908 33980 27936 34011
rect 26620 33952 27936 33980
rect 28000 33980 28028 34011
rect 29365 33983 29423 33989
rect 29365 33980 29377 33983
rect 28000 33952 29377 33980
rect 10100 33884 11008 33912
rect 10100 33872 10106 33884
rect 5718 33804 5724 33856
rect 5776 33844 5782 33856
rect 8294 33844 8300 33856
rect 5776 33816 8300 33844
rect 5776 33804 5782 33816
rect 8294 33804 8300 33816
rect 8352 33804 8358 33856
rect 10980 33844 11008 33884
rect 26234 33872 26240 33924
rect 26292 33912 26298 33924
rect 26620 33921 26648 33952
rect 29365 33949 29377 33952
rect 29411 33949 29423 33983
rect 29365 33943 29423 33949
rect 29454 33940 29460 33992
rect 29512 33980 29518 33992
rect 29917 33983 29975 33989
rect 29917 33980 29929 33983
rect 29512 33952 29929 33980
rect 29512 33940 29518 33952
rect 29917 33949 29929 33952
rect 29963 33949 29975 33983
rect 29917 33943 29975 33949
rect 30193 33983 30251 33989
rect 30193 33949 30205 33983
rect 30239 33980 30251 33983
rect 30239 33952 30972 33980
rect 30239 33949 30251 33952
rect 30193 33943 30251 33949
rect 26605 33915 26663 33921
rect 26605 33912 26617 33915
rect 26292 33884 26617 33912
rect 26292 33872 26298 33884
rect 26605 33881 26617 33884
rect 26651 33881 26663 33915
rect 30944 33912 30972 33952
rect 31570 33940 31576 33992
rect 31628 33980 31634 33992
rect 32140 33989 32168 34156
rect 34882 34144 34888 34156
rect 34940 34184 34946 34196
rect 34940 34156 35480 34184
rect 34940 34144 34946 34156
rect 34974 34116 34980 34128
rect 34935 34088 34980 34116
rect 34974 34076 34980 34088
rect 35032 34076 35038 34128
rect 32217 34051 32275 34057
rect 32217 34017 32229 34051
rect 32263 34048 32275 34051
rect 32306 34048 32312 34060
rect 32263 34020 32312 34048
rect 32263 34017 32275 34020
rect 32217 34011 32275 34017
rect 32306 34008 32312 34020
rect 32364 34008 32370 34060
rect 32490 34008 32496 34060
rect 32548 34048 32554 34060
rect 33321 34051 33379 34057
rect 33321 34048 33333 34051
rect 32548 34020 33333 34048
rect 32548 34008 32554 34020
rect 33321 34017 33333 34020
rect 33367 34048 33379 34051
rect 34514 34048 34520 34060
rect 33367 34020 34520 34048
rect 33367 34017 33379 34020
rect 33321 34011 33379 34017
rect 34514 34008 34520 34020
rect 34572 34008 34578 34060
rect 35452 34057 35480 34156
rect 35437 34051 35495 34057
rect 35437 34017 35449 34051
rect 35483 34017 35495 34051
rect 35437 34011 35495 34017
rect 35529 34051 35587 34057
rect 35529 34017 35541 34051
rect 35575 34048 35587 34051
rect 36078 34048 36084 34060
rect 35575 34020 36084 34048
rect 35575 34017 35587 34020
rect 35529 34011 35587 34017
rect 36078 34008 36084 34020
rect 36136 34008 36142 34060
rect 32125 33983 32183 33989
rect 32125 33980 32137 33983
rect 31628 33952 32137 33980
rect 31628 33940 31634 33952
rect 32125 33949 32137 33952
rect 32171 33949 32183 33983
rect 32125 33943 32183 33949
rect 32677 33983 32735 33989
rect 32677 33949 32689 33983
rect 32723 33949 32735 33983
rect 32677 33943 32735 33949
rect 33597 33983 33655 33989
rect 33597 33949 33609 33983
rect 33643 33980 33655 33983
rect 33643 33952 34284 33980
rect 33643 33949 33655 33952
rect 33597 33943 33655 33949
rect 32692 33912 32720 33943
rect 30944 33884 32720 33912
rect 26605 33875 26663 33881
rect 13170 33844 13176 33856
rect 10980 33816 13176 33844
rect 13170 33804 13176 33816
rect 13228 33804 13234 33856
rect 18141 33847 18199 33853
rect 18141 33813 18153 33847
rect 18187 33844 18199 33847
rect 18414 33844 18420 33856
rect 18187 33816 18420 33844
rect 18187 33813 18199 33816
rect 18141 33807 18199 33813
rect 18414 33804 18420 33816
rect 18472 33804 18478 33856
rect 20254 33844 20260 33856
rect 20215 33816 20260 33844
rect 20254 33804 20260 33816
rect 20312 33804 20318 33856
rect 21634 33804 21640 33856
rect 21692 33844 21698 33856
rect 21729 33847 21787 33853
rect 21729 33844 21741 33847
rect 21692 33816 21741 33844
rect 21692 33804 21698 33816
rect 21729 33813 21741 33816
rect 21775 33813 21787 33847
rect 23566 33844 23572 33856
rect 23527 33816 23572 33844
rect 21729 33807 21787 33813
rect 23566 33804 23572 33816
rect 23624 33804 23630 33856
rect 24394 33844 24400 33856
rect 24355 33816 24400 33844
rect 24394 33804 24400 33816
rect 24452 33804 24458 33856
rect 24854 33804 24860 33856
rect 24912 33844 24918 33856
rect 25409 33847 25467 33853
rect 25409 33844 25421 33847
rect 24912 33816 25421 33844
rect 24912 33804 24918 33816
rect 25409 33813 25421 33816
rect 25455 33813 25467 33847
rect 28166 33844 28172 33856
rect 28127 33816 28172 33844
rect 25409 33807 25467 33813
rect 28166 33804 28172 33816
rect 28224 33804 28230 33856
rect 34256 33844 34284 33952
rect 35713 33847 35771 33853
rect 35713 33844 35725 33847
rect 34256 33816 35725 33844
rect 35713 33813 35725 33816
rect 35759 33813 35771 33847
rect 35713 33807 35771 33813
rect 1104 33754 39836 33776
rect 1104 33702 4246 33754
rect 4298 33702 4310 33754
rect 4362 33702 4374 33754
rect 4426 33702 4438 33754
rect 4490 33702 34966 33754
rect 35018 33702 35030 33754
rect 35082 33702 35094 33754
rect 35146 33702 35158 33754
rect 35210 33702 39836 33754
rect 1104 33680 39836 33702
rect 3142 33600 3148 33652
rect 3200 33640 3206 33652
rect 4893 33643 4951 33649
rect 4893 33640 4905 33643
rect 3200 33612 4905 33640
rect 3200 33600 3206 33612
rect 4893 33609 4905 33612
rect 4939 33640 4951 33643
rect 5074 33640 5080 33652
rect 4939 33612 5080 33640
rect 4939 33609 4951 33612
rect 4893 33603 4951 33609
rect 5074 33600 5080 33612
rect 5132 33600 5138 33652
rect 7190 33600 7196 33652
rect 7248 33640 7254 33652
rect 8570 33640 8576 33652
rect 7248 33612 8576 33640
rect 7248 33600 7254 33612
rect 8570 33600 8576 33612
rect 8628 33600 8634 33652
rect 9217 33643 9275 33649
rect 9217 33609 9229 33643
rect 9263 33640 9275 33643
rect 11238 33640 11244 33652
rect 9263 33612 11244 33640
rect 9263 33609 9275 33612
rect 9217 33603 9275 33609
rect 11238 33600 11244 33612
rect 11296 33600 11302 33652
rect 19981 33643 20039 33649
rect 19981 33609 19993 33643
rect 20027 33640 20039 33643
rect 20162 33640 20168 33652
rect 20027 33612 20168 33640
rect 20027 33609 20039 33612
rect 19981 33603 20039 33609
rect 20162 33600 20168 33612
rect 20220 33600 20226 33652
rect 23845 33643 23903 33649
rect 23845 33640 23857 33643
rect 21744 33612 23857 33640
rect 5552 33544 7880 33572
rect 3786 33504 3792 33516
rect 3747 33476 3792 33504
rect 3786 33464 3792 33476
rect 3844 33464 3850 33516
rect 5552 33513 5580 33544
rect 5537 33507 5595 33513
rect 5537 33473 5549 33507
rect 5583 33473 5595 33507
rect 6730 33504 6736 33516
rect 5537 33467 5595 33473
rect 5736 33476 6736 33504
rect 2774 33396 2780 33448
rect 2832 33436 2838 33448
rect 3326 33436 3332 33448
rect 2832 33408 2877 33436
rect 3287 33408 3332 33436
rect 2832 33396 2838 33408
rect 3326 33396 3332 33408
rect 3384 33396 3390 33448
rect 3694 33436 3700 33448
rect 3655 33408 3700 33436
rect 3694 33396 3700 33408
rect 3752 33396 3758 33448
rect 4249 33439 4307 33445
rect 4249 33405 4261 33439
rect 4295 33436 4307 33439
rect 4706 33436 4712 33448
rect 4295 33408 4712 33436
rect 4295 33405 4307 33408
rect 4249 33399 4307 33405
rect 4706 33396 4712 33408
rect 4764 33396 4770 33448
rect 5736 33445 5764 33476
rect 6730 33464 6736 33476
rect 6788 33464 6794 33516
rect 6914 33504 6920 33516
rect 6875 33476 6920 33504
rect 6914 33464 6920 33476
rect 6972 33464 6978 33516
rect 5721 33439 5779 33445
rect 5721 33405 5733 33439
rect 5767 33405 5779 33439
rect 7098 33436 7104 33448
rect 5721 33399 5779 33405
rect 5920 33408 7104 33436
rect 5920 33377 5948 33408
rect 7098 33396 7104 33408
rect 7156 33396 7162 33448
rect 7852 33445 7880 33544
rect 8202 33532 8208 33584
rect 8260 33572 8266 33584
rect 13354 33572 13360 33584
rect 8260 33544 13360 33572
rect 8260 33532 8266 33544
rect 13354 33532 13360 33544
rect 13412 33532 13418 33584
rect 21634 33572 21640 33584
rect 19444 33544 21640 33572
rect 8757 33507 8815 33513
rect 8757 33473 8769 33507
rect 8803 33504 8815 33507
rect 9953 33507 10011 33513
rect 9953 33504 9965 33507
rect 8803 33476 9965 33504
rect 8803 33473 8815 33476
rect 8757 33467 8815 33473
rect 9953 33473 9965 33476
rect 9999 33473 10011 33507
rect 9953 33467 10011 33473
rect 14829 33507 14887 33513
rect 14829 33473 14841 33507
rect 14875 33504 14887 33507
rect 16206 33504 16212 33516
rect 14875 33476 16212 33504
rect 14875 33473 14887 33476
rect 14829 33467 14887 33473
rect 16206 33464 16212 33476
rect 16264 33464 16270 33516
rect 7469 33439 7527 33445
rect 7469 33405 7481 33439
rect 7515 33405 7527 33439
rect 7469 33399 7527 33405
rect 7837 33439 7895 33445
rect 7837 33405 7849 33439
rect 7883 33405 7895 33439
rect 8110 33436 8116 33448
rect 8071 33408 8116 33436
rect 7837 33399 7895 33405
rect 5905 33371 5963 33377
rect 5905 33337 5917 33371
rect 5951 33337 5963 33371
rect 5905 33331 5963 33337
rect 6273 33371 6331 33377
rect 6273 33337 6285 33371
rect 6319 33368 6331 33371
rect 7374 33368 7380 33380
rect 6319 33340 7380 33368
rect 6319 33337 6331 33340
rect 6273 33331 6331 33337
rect 7374 33328 7380 33340
rect 7432 33328 7438 33380
rect 5813 33303 5871 33309
rect 5813 33269 5825 33303
rect 5859 33300 5871 33303
rect 7190 33300 7196 33312
rect 5859 33272 7196 33300
rect 5859 33269 5871 33272
rect 5813 33263 5871 33269
rect 7190 33260 7196 33272
rect 7248 33260 7254 33312
rect 7484 33300 7512 33399
rect 7852 33368 7880 33399
rect 8110 33396 8116 33408
rect 8168 33396 8174 33448
rect 8294 33396 8300 33448
rect 8352 33436 8358 33448
rect 8941 33439 8999 33445
rect 8941 33436 8953 33439
rect 8352 33408 8953 33436
rect 8352 33396 8358 33408
rect 8941 33405 8953 33408
rect 8987 33405 8999 33439
rect 8941 33399 8999 33405
rect 9033 33439 9091 33445
rect 9033 33405 9045 33439
rect 9079 33436 9091 33439
rect 10318 33436 10324 33448
rect 9079 33408 10324 33436
rect 9079 33405 9091 33408
rect 9033 33399 9091 33405
rect 10318 33396 10324 33408
rect 10376 33396 10382 33448
rect 10502 33436 10508 33448
rect 10463 33408 10508 33436
rect 10502 33396 10508 33408
rect 10560 33396 10566 33448
rect 10594 33396 10600 33448
rect 10652 33436 10658 33448
rect 10781 33439 10839 33445
rect 10652 33408 10697 33436
rect 10652 33396 10658 33408
rect 10781 33405 10793 33439
rect 10827 33405 10839 33439
rect 11054 33436 11060 33448
rect 11015 33408 11060 33436
rect 10781 33399 10839 33405
rect 8846 33368 8852 33380
rect 7852 33340 8852 33368
rect 8846 33328 8852 33340
rect 8904 33328 8910 33380
rect 9582 33328 9588 33380
rect 9640 33368 9646 33380
rect 10796 33368 10824 33399
rect 11054 33396 11060 33408
rect 11112 33396 11118 33448
rect 11241 33439 11299 33445
rect 11241 33405 11253 33439
rect 11287 33405 11299 33439
rect 13630 33436 13636 33448
rect 13591 33408 13636 33436
rect 11241 33399 11299 33405
rect 9640 33340 10824 33368
rect 9640 33328 9646 33340
rect 10962 33328 10968 33380
rect 11020 33368 11026 33380
rect 11256 33368 11284 33399
rect 13630 33396 13636 33408
rect 13688 33396 13694 33448
rect 13906 33436 13912 33448
rect 13867 33408 13912 33436
rect 13906 33396 13912 33408
rect 13964 33396 13970 33448
rect 13998 33396 14004 33448
rect 14056 33436 14062 33448
rect 14093 33439 14151 33445
rect 14093 33436 14105 33439
rect 14056 33408 14105 33436
rect 14056 33396 14062 33408
rect 14093 33405 14105 33408
rect 14139 33405 14151 33439
rect 15102 33436 15108 33448
rect 15063 33408 15108 33436
rect 14093 33399 14151 33405
rect 15102 33396 15108 33408
rect 15160 33396 15166 33448
rect 16574 33396 16580 33448
rect 16632 33436 16638 33448
rect 19444 33445 19472 33544
rect 21634 33532 21640 33544
rect 21692 33532 21698 33584
rect 19705 33507 19763 33513
rect 19705 33473 19717 33507
rect 19751 33504 19763 33507
rect 20346 33504 20352 33516
rect 19751 33476 20352 33504
rect 19751 33473 19763 33476
rect 19705 33467 19763 33473
rect 20346 33464 20352 33476
rect 20404 33464 20410 33516
rect 20717 33507 20775 33513
rect 20717 33473 20729 33507
rect 20763 33504 20775 33507
rect 21082 33504 21088 33516
rect 20763 33476 21088 33504
rect 20763 33473 20775 33476
rect 20717 33467 20775 33473
rect 21082 33464 21088 33476
rect 21140 33504 21146 33516
rect 21744 33513 21772 33612
rect 23845 33609 23857 33612
rect 23891 33640 23903 33643
rect 24118 33640 24124 33652
rect 23891 33612 24124 33640
rect 23891 33609 23903 33612
rect 23845 33603 23903 33609
rect 24118 33600 24124 33612
rect 24176 33600 24182 33652
rect 24486 33600 24492 33652
rect 24544 33640 24550 33652
rect 29546 33640 29552 33652
rect 24544 33612 29552 33640
rect 24544 33600 24550 33612
rect 29546 33600 29552 33612
rect 29604 33640 29610 33652
rect 31570 33640 31576 33652
rect 29604 33612 30880 33640
rect 31531 33612 31576 33640
rect 29604 33600 29610 33612
rect 21729 33507 21787 33513
rect 21729 33504 21741 33507
rect 21140 33476 21741 33504
rect 21140 33464 21146 33476
rect 21729 33473 21741 33476
rect 21775 33473 21787 33507
rect 22278 33504 22284 33516
rect 22239 33476 22284 33504
rect 21729 33467 21787 33473
rect 22278 33464 22284 33476
rect 22336 33464 22342 33516
rect 23198 33464 23204 33516
rect 23256 33504 23262 33516
rect 24581 33507 24639 33513
rect 24581 33504 24593 33507
rect 23256 33476 24593 33504
rect 23256 33464 23262 33476
rect 24581 33473 24593 33476
rect 24627 33473 24639 33507
rect 24854 33504 24860 33516
rect 24815 33476 24860 33504
rect 24581 33467 24639 33473
rect 17037 33439 17095 33445
rect 17037 33436 17049 33439
rect 16632 33408 17049 33436
rect 16632 33396 16638 33408
rect 17037 33405 17049 33408
rect 17083 33405 17095 33439
rect 17037 33399 17095 33405
rect 19429 33439 19487 33445
rect 19429 33405 19441 33439
rect 19475 33405 19487 33439
rect 19429 33399 19487 33405
rect 19797 33439 19855 33445
rect 19797 33405 19809 33439
rect 19843 33436 19855 33439
rect 20530 33436 20536 33448
rect 19843 33408 20536 33436
rect 19843 33405 19855 33408
rect 19797 33399 19855 33405
rect 20530 33396 20536 33408
rect 20588 33396 20594 33448
rect 20806 33436 20812 33448
rect 20767 33408 20812 33436
rect 20806 33396 20812 33408
rect 20864 33396 20870 33448
rect 21818 33396 21824 33448
rect 21876 33436 21882 33448
rect 23661 33439 23719 33445
rect 21876 33408 21921 33436
rect 21876 33396 21882 33408
rect 23661 33405 23673 33439
rect 23707 33436 23719 33439
rect 24486 33436 24492 33448
rect 23707 33408 24492 33436
rect 23707 33405 23719 33408
rect 23661 33399 23719 33405
rect 24486 33396 24492 33408
rect 24544 33396 24550 33448
rect 24596 33436 24624 33467
rect 24854 33464 24860 33476
rect 24912 33464 24918 33516
rect 27154 33504 27160 33516
rect 26712 33476 27160 33504
rect 26712 33445 26740 33476
rect 27154 33464 27160 33476
rect 27212 33504 27218 33516
rect 29273 33507 29331 33513
rect 29273 33504 29285 33507
rect 27212 33476 29285 33504
rect 27212 33464 27218 33476
rect 29273 33473 29285 33476
rect 29319 33504 29331 33507
rect 29454 33504 29460 33516
rect 29319 33476 29460 33504
rect 29319 33473 29331 33476
rect 29273 33467 29331 33473
rect 29454 33464 29460 33476
rect 29512 33464 29518 33516
rect 29549 33507 29607 33513
rect 29549 33473 29561 33507
rect 29595 33504 29607 33507
rect 30650 33504 30656 33516
rect 29595 33476 30656 33504
rect 29595 33473 29607 33476
rect 29549 33467 29607 33473
rect 30650 33464 30656 33476
rect 30708 33464 30714 33516
rect 26697 33439 26755 33445
rect 26697 33436 26709 33439
rect 24596 33408 26709 33436
rect 26697 33405 26709 33408
rect 26743 33405 26755 33439
rect 26697 33399 26755 33405
rect 26973 33439 27031 33445
rect 26973 33405 26985 33439
rect 27019 33436 27031 33439
rect 27614 33436 27620 33448
rect 27019 33408 27620 33436
rect 27019 33405 27031 33408
rect 26973 33399 27031 33405
rect 27614 33396 27620 33408
rect 27672 33396 27678 33448
rect 30852 33436 30880 33612
rect 31570 33600 31576 33612
rect 31628 33600 31634 33652
rect 33689 33643 33747 33649
rect 33689 33609 33701 33643
rect 33735 33640 33747 33643
rect 33778 33640 33784 33652
rect 33735 33612 33784 33640
rect 33735 33609 33747 33612
rect 33689 33603 33747 33609
rect 33778 33600 33784 33612
rect 33836 33600 33842 33652
rect 32309 33507 32367 33513
rect 32309 33473 32321 33507
rect 32355 33504 32367 33507
rect 32490 33504 32496 33516
rect 32355 33476 32496 33504
rect 32355 33473 32367 33476
rect 32309 33467 32367 33473
rect 32490 33464 32496 33476
rect 32548 33464 32554 33516
rect 32585 33507 32643 33513
rect 32585 33473 32597 33507
rect 32631 33504 32643 33507
rect 33226 33504 33232 33516
rect 32631 33476 33232 33504
rect 32631 33473 32643 33476
rect 32585 33467 32643 33473
rect 33226 33464 33232 33476
rect 33284 33464 33290 33516
rect 35161 33507 35219 33513
rect 35161 33473 35173 33507
rect 35207 33504 35219 33507
rect 35250 33504 35256 33516
rect 35207 33476 35256 33504
rect 35207 33473 35219 33476
rect 35161 33467 35219 33473
rect 35250 33464 35256 33476
rect 35308 33464 35314 33516
rect 31389 33439 31447 33445
rect 31389 33436 31401 33439
rect 30852 33408 31401 33436
rect 31389 33405 31401 33408
rect 31435 33405 31447 33439
rect 31389 33399 31447 33405
rect 34514 33396 34520 33448
rect 34572 33436 34578 33448
rect 34885 33439 34943 33445
rect 34885 33436 34897 33439
rect 34572 33408 34897 33436
rect 34572 33396 34578 33408
rect 34885 33405 34897 33408
rect 34931 33405 34943 33439
rect 34885 33399 34943 33405
rect 11020 33340 11284 33368
rect 13081 33371 13139 33377
rect 11020 33328 11026 33340
rect 13081 33337 13093 33371
rect 13127 33368 13139 33371
rect 13446 33368 13452 33380
rect 13127 33340 13452 33368
rect 13127 33337 13139 33340
rect 13081 33331 13139 33337
rect 13446 33328 13452 33340
rect 13504 33328 13510 33380
rect 21174 33328 21180 33380
rect 21232 33368 21238 33380
rect 21269 33371 21327 33377
rect 21269 33368 21281 33371
rect 21232 33340 21281 33368
rect 21232 33328 21238 33340
rect 21269 33337 21281 33340
rect 21315 33337 21327 33371
rect 21269 33331 21327 33337
rect 36541 33371 36599 33377
rect 36541 33337 36553 33371
rect 36587 33368 36599 33371
rect 36998 33368 37004 33380
rect 36587 33340 37004 33368
rect 36587 33337 36599 33340
rect 36541 33331 36599 33337
rect 36998 33328 37004 33340
rect 37056 33328 37062 33380
rect 8754 33300 8760 33312
rect 7484 33272 8760 33300
rect 8754 33260 8760 33272
rect 8812 33260 8818 33312
rect 15838 33260 15844 33312
rect 15896 33300 15902 33312
rect 16209 33303 16267 33309
rect 16209 33300 16221 33303
rect 15896 33272 16221 33300
rect 15896 33260 15902 33272
rect 16209 33269 16221 33272
rect 16255 33269 16267 33303
rect 17126 33300 17132 33312
rect 17087 33272 17132 33300
rect 16209 33263 16267 33269
rect 17126 33260 17132 33272
rect 17184 33260 17190 33312
rect 17954 33260 17960 33312
rect 18012 33300 18018 33312
rect 19242 33300 19248 33312
rect 18012 33272 19248 33300
rect 18012 33260 18018 33272
rect 19242 33260 19248 33272
rect 19300 33260 19306 33312
rect 23750 33260 23756 33312
rect 23808 33300 23814 33312
rect 25961 33303 26019 33309
rect 25961 33300 25973 33303
rect 23808 33272 25973 33300
rect 23808 33260 23814 33272
rect 25961 33269 25973 33272
rect 26007 33269 26019 33303
rect 25961 33263 26019 33269
rect 27890 33260 27896 33312
rect 27948 33300 27954 33312
rect 28077 33303 28135 33309
rect 28077 33300 28089 33303
rect 27948 33272 28089 33300
rect 27948 33260 27954 33272
rect 28077 33269 28089 33272
rect 28123 33269 28135 33303
rect 28077 33263 28135 33269
rect 30837 33303 30895 33309
rect 30837 33269 30849 33303
rect 30883 33300 30895 33303
rect 31478 33300 31484 33312
rect 30883 33272 31484 33300
rect 30883 33269 30895 33272
rect 30837 33263 30895 33269
rect 31478 33260 31484 33272
rect 31536 33260 31542 33312
rect 1104 33210 39836 33232
rect 1104 33158 19606 33210
rect 19658 33158 19670 33210
rect 19722 33158 19734 33210
rect 19786 33158 19798 33210
rect 19850 33158 39836 33210
rect 1104 33136 39836 33158
rect 5994 33096 6000 33108
rect 4356 33068 6000 33096
rect 3053 33031 3111 33037
rect 3053 32997 3065 33031
rect 3099 33028 3111 33031
rect 3326 33028 3332 33040
rect 3099 33000 3332 33028
rect 3099 32997 3111 33000
rect 3053 32991 3111 32997
rect 3326 32988 3332 33000
rect 3384 32988 3390 33040
rect 1397 32963 1455 32969
rect 1397 32929 1409 32963
rect 1443 32960 1455 32963
rect 2682 32960 2688 32972
rect 1443 32932 2688 32960
rect 1443 32929 1455 32932
rect 1397 32923 1455 32929
rect 2682 32920 2688 32932
rect 2740 32920 2746 32972
rect 4356 32969 4384 33068
rect 5994 33056 6000 33068
rect 6052 33056 6058 33108
rect 8386 33056 8392 33108
rect 8444 33096 8450 33108
rect 9309 33099 9367 33105
rect 9309 33096 9321 33099
rect 8444 33068 9321 33096
rect 8444 33056 8450 33068
rect 9309 33065 9321 33068
rect 9355 33065 9367 33099
rect 9309 33059 9367 33065
rect 10962 33056 10968 33108
rect 11020 33096 11026 33108
rect 14737 33099 14795 33105
rect 11020 33068 11468 33096
rect 11020 33056 11026 33068
rect 4433 33031 4491 33037
rect 4433 32997 4445 33031
rect 4479 33028 4491 33031
rect 4614 33028 4620 33040
rect 4479 33000 4620 33028
rect 4479 32997 4491 33000
rect 4433 32991 4491 32997
rect 4614 32988 4620 33000
rect 4672 32988 4678 33040
rect 5074 32988 5080 33040
rect 5132 33028 5138 33040
rect 5132 33000 5764 33028
rect 5132 32988 5138 33000
rect 4341 32963 4399 32969
rect 4341 32929 4353 32963
rect 4387 32929 4399 32963
rect 4706 32960 4712 32972
rect 4667 32932 4712 32960
rect 4341 32923 4399 32929
rect 4706 32920 4712 32932
rect 4764 32920 4770 32972
rect 4982 32960 4988 32972
rect 4943 32932 4988 32960
rect 4982 32920 4988 32932
rect 5040 32920 5046 32972
rect 5736 32969 5764 33000
rect 8938 32988 8944 33040
rect 8996 33028 9002 33040
rect 11149 33031 11207 33037
rect 11149 33028 11161 33031
rect 8996 33000 11161 33028
rect 8996 32988 9002 33000
rect 11149 32997 11161 33000
rect 11195 32997 11207 33031
rect 11440 33028 11468 33068
rect 14737 33065 14749 33099
rect 14783 33096 14795 33099
rect 15102 33096 15108 33108
rect 14783 33068 15108 33096
rect 14783 33065 14795 33068
rect 14737 33059 14795 33065
rect 15102 33056 15108 33068
rect 15160 33056 15166 33108
rect 16666 33096 16672 33108
rect 15212 33068 16672 33096
rect 11509 33031 11567 33037
rect 11509 33028 11521 33031
rect 11440 33000 11521 33028
rect 11149 32991 11207 32997
rect 11509 32997 11521 33000
rect 11555 32997 11567 33031
rect 11509 32991 11567 32997
rect 13354 32988 13360 33040
rect 13412 33028 13418 33040
rect 15212 33028 15240 33068
rect 16666 33056 16672 33068
rect 16724 33056 16730 33108
rect 24765 33099 24823 33105
rect 24765 33065 24777 33099
rect 24811 33096 24823 33099
rect 25222 33096 25228 33108
rect 24811 33068 25228 33096
rect 24811 33065 24823 33068
rect 24765 33059 24823 33065
rect 25222 33056 25228 33068
rect 25280 33056 25286 33108
rect 30469 33099 30527 33105
rect 30469 33065 30481 33099
rect 30515 33096 30527 33099
rect 31294 33096 31300 33108
rect 30515 33068 31300 33096
rect 30515 33065 30527 33068
rect 30469 33059 30527 33065
rect 16574 33028 16580 33040
rect 13412 33000 15240 33028
rect 15764 33000 16580 33028
rect 13412 32988 13418 33000
rect 5353 32963 5411 32969
rect 5353 32929 5365 32963
rect 5399 32929 5411 32963
rect 5353 32923 5411 32929
rect 5721 32963 5779 32969
rect 5721 32929 5733 32963
rect 5767 32929 5779 32963
rect 8570 32960 8576 32972
rect 8531 32932 8576 32960
rect 5721 32923 5779 32929
rect 1670 32892 1676 32904
rect 1631 32864 1676 32892
rect 1670 32852 1676 32864
rect 1728 32852 1734 32904
rect 4062 32852 4068 32904
rect 4120 32892 4126 32904
rect 5368 32892 5396 32923
rect 8570 32920 8576 32932
rect 8628 32920 8634 32972
rect 9122 32920 9128 32972
rect 9180 32960 9186 32972
rect 9493 32963 9551 32969
rect 9493 32960 9505 32963
rect 9180 32932 9505 32960
rect 9180 32920 9186 32932
rect 9493 32929 9505 32932
rect 9539 32929 9551 32963
rect 9493 32923 9551 32929
rect 10505 32963 10563 32969
rect 10505 32929 10517 32963
rect 10551 32960 10563 32963
rect 11330 32960 11336 32972
rect 10551 32932 11192 32960
rect 11291 32932 11336 32960
rect 10551 32929 10563 32932
rect 10505 32923 10563 32929
rect 4120 32864 5396 32892
rect 4120 32852 4126 32864
rect 6086 32852 6092 32904
rect 6144 32892 6150 32904
rect 6454 32892 6460 32904
rect 6144 32864 6460 32892
rect 6144 32852 6150 32864
rect 6454 32852 6460 32864
rect 6512 32852 6518 32904
rect 6730 32892 6736 32904
rect 6691 32864 6736 32892
rect 6730 32852 6736 32864
rect 6788 32852 6794 32904
rect 9674 32892 9680 32904
rect 9635 32864 9680 32892
rect 9674 32852 9680 32864
rect 9732 32852 9738 32904
rect 10226 32892 10232 32904
rect 10187 32864 10232 32892
rect 10226 32852 10232 32864
rect 10284 32852 10290 32904
rect 10689 32895 10747 32901
rect 10689 32861 10701 32895
rect 10735 32892 10747 32895
rect 11054 32892 11060 32904
rect 10735 32864 11060 32892
rect 10735 32861 10747 32864
rect 10689 32855 10747 32861
rect 11054 32852 11060 32864
rect 11112 32852 11118 32904
rect 11164 32892 11192 32932
rect 11330 32920 11336 32932
rect 11388 32920 11394 32972
rect 11422 32920 11428 32972
rect 11480 32960 11486 32972
rect 13924 32969 13952 33000
rect 13909 32963 13967 32969
rect 11480 32932 11525 32960
rect 11480 32920 11486 32932
rect 13909 32929 13921 32963
rect 13955 32929 13967 32963
rect 14458 32960 14464 32972
rect 14419 32932 14464 32960
rect 13909 32923 13967 32929
rect 14458 32920 14464 32932
rect 14516 32920 14522 32972
rect 15654 32960 15660 32972
rect 15615 32932 15660 32960
rect 15654 32920 15660 32932
rect 15712 32920 15718 32972
rect 15764 32969 15792 33000
rect 16574 32988 16580 33000
rect 16632 32988 16638 33040
rect 30484 33028 30512 33059
rect 31294 33056 31300 33068
rect 31352 33056 31358 33108
rect 29472 33000 30512 33028
rect 15749 32963 15807 32969
rect 15749 32929 15761 32963
rect 15795 32929 15807 32963
rect 16114 32960 16120 32972
rect 16075 32932 16120 32960
rect 15749 32923 15807 32929
rect 16114 32920 16120 32932
rect 16172 32920 16178 32972
rect 16206 32920 16212 32972
rect 16264 32960 16270 32972
rect 16853 32963 16911 32969
rect 16264 32932 16620 32960
rect 16264 32920 16270 32932
rect 11885 32895 11943 32901
rect 11885 32892 11897 32895
rect 11164 32864 11897 32892
rect 11885 32861 11897 32864
rect 11931 32861 11943 32895
rect 11885 32855 11943 32861
rect 14553 32895 14611 32901
rect 14553 32861 14565 32895
rect 14599 32892 14611 32895
rect 16390 32892 16396 32904
rect 14599 32864 16396 32892
rect 14599 32861 14611 32864
rect 14553 32855 14611 32861
rect 16390 32852 16396 32864
rect 16448 32852 16454 32904
rect 16592 32901 16620 32932
rect 16853 32929 16865 32963
rect 16899 32960 16911 32963
rect 17126 32960 17132 32972
rect 16899 32932 17132 32960
rect 16899 32929 16911 32932
rect 16853 32923 16911 32929
rect 17126 32920 17132 32932
rect 17184 32920 17190 32972
rect 19886 32920 19892 32972
rect 19944 32960 19950 32972
rect 20438 32960 20444 32972
rect 19944 32932 20444 32960
rect 19944 32920 19950 32932
rect 20438 32920 20444 32932
rect 20496 32960 20502 32972
rect 20901 32963 20959 32969
rect 20901 32960 20913 32963
rect 20496 32932 20913 32960
rect 20496 32920 20502 32932
rect 20901 32929 20913 32932
rect 20947 32929 20959 32963
rect 21174 32960 21180 32972
rect 21135 32932 21180 32960
rect 20901 32923 20959 32929
rect 16577 32895 16635 32901
rect 16577 32861 16589 32895
rect 16623 32861 16635 32895
rect 16577 32855 16635 32861
rect 18322 32852 18328 32904
rect 18380 32892 18386 32904
rect 18693 32895 18751 32901
rect 18693 32892 18705 32895
rect 18380 32864 18705 32892
rect 18380 32852 18386 32864
rect 18693 32861 18705 32864
rect 18739 32861 18751 32895
rect 18966 32892 18972 32904
rect 18927 32864 18972 32892
rect 18693 32855 18751 32861
rect 18966 32852 18972 32864
rect 19024 32852 19030 32904
rect 20916 32892 20944 32923
rect 21174 32920 21180 32932
rect 21232 32920 21238 32972
rect 22557 32963 22615 32969
rect 22557 32929 22569 32963
rect 22603 32960 22615 32963
rect 23477 32963 23535 32969
rect 22603 32932 23428 32960
rect 22603 32929 22615 32932
rect 22557 32923 22615 32929
rect 23198 32892 23204 32904
rect 20916 32864 23204 32892
rect 23198 32852 23204 32864
rect 23256 32852 23262 32904
rect 23400 32892 23428 32932
rect 23477 32929 23489 32963
rect 23523 32960 23535 32963
rect 24394 32960 24400 32972
rect 23523 32932 24400 32960
rect 23523 32929 23535 32932
rect 23477 32923 23535 32929
rect 24394 32920 24400 32932
rect 24452 32920 24458 32972
rect 25409 32963 25467 32969
rect 25409 32960 25421 32963
rect 24504 32932 25421 32960
rect 24504 32892 24532 32932
rect 25409 32929 25421 32932
rect 25455 32929 25467 32963
rect 28813 32963 28871 32969
rect 25409 32923 25467 32929
rect 27080 32932 28580 32960
rect 23400 32864 24532 32892
rect 25130 32852 25136 32904
rect 25188 32892 25194 32904
rect 25317 32895 25375 32901
rect 25317 32892 25329 32895
rect 25188 32864 25329 32892
rect 25188 32852 25194 32864
rect 25317 32861 25329 32864
rect 25363 32892 25375 32895
rect 27080 32892 27108 32932
rect 25363 32864 27108 32892
rect 25363 32861 25375 32864
rect 25317 32855 25375 32861
rect 27154 32852 27160 32904
rect 27212 32892 27218 32904
rect 27430 32892 27436 32904
rect 27212 32864 27257 32892
rect 27391 32864 27436 32892
rect 27212 32852 27218 32864
rect 27430 32852 27436 32864
rect 27488 32852 27494 32904
rect 28552 32892 28580 32932
rect 28813 32929 28825 32963
rect 28859 32960 28871 32963
rect 29365 32963 29423 32969
rect 29365 32960 29377 32963
rect 28859 32932 29377 32960
rect 28859 32929 28871 32932
rect 28813 32923 28871 32929
rect 29365 32929 29377 32932
rect 29411 32929 29423 32963
rect 29365 32923 29423 32929
rect 29270 32892 29276 32904
rect 28552 32864 29276 32892
rect 29270 32852 29276 32864
rect 29328 32892 29334 32904
rect 29472 32892 29500 33000
rect 29546 32920 29552 32972
rect 29604 32960 29610 32972
rect 30285 32963 30343 32969
rect 30285 32960 30297 32963
rect 29604 32932 30297 32960
rect 29604 32920 29610 32932
rect 30285 32929 30297 32932
rect 30331 32929 30343 32963
rect 30285 32923 30343 32929
rect 30374 32920 30380 32972
rect 30432 32960 30438 32972
rect 32125 32963 32183 32969
rect 32125 32960 32137 32963
rect 30432 32932 32137 32960
rect 30432 32920 30438 32932
rect 32125 32929 32137 32932
rect 32171 32929 32183 32963
rect 32858 32960 32864 32972
rect 32819 32932 32864 32960
rect 32125 32923 32183 32929
rect 32858 32920 32864 32932
rect 32916 32920 32922 32972
rect 33689 32963 33747 32969
rect 33689 32929 33701 32963
rect 33735 32960 33747 32963
rect 33778 32960 33784 32972
rect 33735 32932 33784 32960
rect 33735 32929 33747 32932
rect 33689 32923 33747 32929
rect 33778 32920 33784 32932
rect 33836 32920 33842 32972
rect 33870 32920 33876 32972
rect 33928 32960 33934 32972
rect 33928 32932 33973 32960
rect 33928 32920 33934 32932
rect 34790 32920 34796 32972
rect 34848 32960 34854 32972
rect 34977 32963 35035 32969
rect 34977 32960 34989 32963
rect 34848 32932 34989 32960
rect 34848 32920 34854 32932
rect 34977 32929 34989 32932
rect 35023 32929 35035 32963
rect 34977 32923 35035 32929
rect 38841 32963 38899 32969
rect 38841 32929 38853 32963
rect 38887 32960 38899 32963
rect 39114 32960 39120 32972
rect 38887 32932 39120 32960
rect 38887 32929 38899 32932
rect 38841 32923 38899 32929
rect 39114 32920 39120 32932
rect 39172 32920 39178 32972
rect 29328 32864 29500 32892
rect 29328 32852 29334 32864
rect 32766 32852 32772 32904
rect 32824 32892 32830 32904
rect 32953 32895 33011 32901
rect 32953 32892 32965 32895
rect 32824 32864 32965 32892
rect 32824 32852 32830 32864
rect 32953 32861 32965 32864
rect 32999 32861 33011 32895
rect 32953 32855 33011 32861
rect 34514 32852 34520 32904
rect 34572 32892 34578 32904
rect 34701 32895 34759 32901
rect 34701 32892 34713 32895
rect 34572 32864 34713 32892
rect 34572 32852 34578 32864
rect 34701 32861 34713 32864
rect 34747 32861 34759 32895
rect 34701 32855 34759 32861
rect 8110 32784 8116 32836
rect 8168 32824 8174 32836
rect 11330 32824 11336 32836
rect 8168 32796 11336 32824
rect 8168 32784 8174 32796
rect 11330 32784 11336 32796
rect 11388 32784 11394 32836
rect 32398 32824 32404 32836
rect 32359 32796 32404 32824
rect 32398 32784 32404 32796
rect 32456 32784 32462 32836
rect 7098 32716 7104 32768
rect 7156 32756 7162 32768
rect 8021 32759 8079 32765
rect 8021 32756 8033 32759
rect 7156 32728 8033 32756
rect 7156 32716 7162 32728
rect 8021 32725 8033 32728
rect 8067 32756 8079 32759
rect 8202 32756 8208 32768
rect 8067 32728 8208 32756
rect 8067 32725 8079 32728
rect 8021 32719 8079 32725
rect 8202 32716 8208 32728
rect 8260 32716 8266 32768
rect 8754 32756 8760 32768
rect 8667 32728 8760 32756
rect 8754 32716 8760 32728
rect 8812 32756 8818 32768
rect 9582 32756 9588 32768
rect 8812 32728 9588 32756
rect 8812 32716 8818 32728
rect 9582 32716 9588 32728
rect 9640 32716 9646 32768
rect 17862 32716 17868 32768
rect 17920 32756 17926 32768
rect 17957 32759 18015 32765
rect 17957 32756 17969 32759
rect 17920 32728 17969 32756
rect 17920 32716 17926 32728
rect 17957 32725 17969 32728
rect 18003 32725 18015 32759
rect 17957 32719 18015 32725
rect 19150 32716 19156 32768
rect 19208 32756 19214 32768
rect 20073 32759 20131 32765
rect 20073 32756 20085 32759
rect 19208 32728 20085 32756
rect 19208 32716 19214 32728
rect 20073 32725 20085 32728
rect 20119 32725 20131 32759
rect 25590 32756 25596 32768
rect 25551 32728 25596 32756
rect 20073 32719 20131 32725
rect 25590 32716 25596 32728
rect 25648 32716 25654 32768
rect 27614 32716 27620 32768
rect 27672 32756 27678 32768
rect 29549 32759 29607 32765
rect 29549 32756 29561 32759
rect 27672 32728 29561 32756
rect 27672 32716 27678 32728
rect 29549 32725 29561 32728
rect 29595 32725 29607 32759
rect 29549 32719 29607 32725
rect 33226 32716 33232 32768
rect 33284 32756 33290 32768
rect 33965 32759 34023 32765
rect 33965 32756 33977 32759
rect 33284 32728 33977 32756
rect 33284 32716 33290 32728
rect 33965 32725 33977 32728
rect 34011 32725 34023 32759
rect 36262 32756 36268 32768
rect 36223 32728 36268 32756
rect 33965 32719 34023 32725
rect 36262 32716 36268 32728
rect 36320 32716 36326 32768
rect 38194 32716 38200 32768
rect 38252 32756 38258 32768
rect 38933 32759 38991 32765
rect 38933 32756 38945 32759
rect 38252 32728 38945 32756
rect 38252 32716 38258 32728
rect 38933 32725 38945 32728
rect 38979 32725 38991 32759
rect 38933 32719 38991 32725
rect 1104 32666 39836 32688
rect 1104 32614 4246 32666
rect 4298 32614 4310 32666
rect 4362 32614 4374 32666
rect 4426 32614 4438 32666
rect 4490 32614 34966 32666
rect 35018 32614 35030 32666
rect 35082 32614 35094 32666
rect 35146 32614 35158 32666
rect 35210 32614 39836 32666
rect 1104 32592 39836 32614
rect 5537 32555 5595 32561
rect 5537 32521 5549 32555
rect 5583 32552 5595 32555
rect 5902 32552 5908 32564
rect 5583 32524 5908 32552
rect 5583 32521 5595 32524
rect 5537 32515 5595 32521
rect 5902 32512 5908 32524
rect 5960 32512 5966 32564
rect 15654 32512 15660 32564
rect 15712 32552 15718 32564
rect 15749 32555 15807 32561
rect 15749 32552 15761 32555
rect 15712 32524 15761 32552
rect 15712 32512 15718 32524
rect 15749 32521 15761 32524
rect 15795 32521 15807 32555
rect 15749 32515 15807 32521
rect 16206 32512 16212 32564
rect 16264 32552 16270 32564
rect 17681 32555 17739 32561
rect 17681 32552 17693 32555
rect 16264 32524 17693 32552
rect 16264 32512 16270 32524
rect 17681 32521 17693 32524
rect 17727 32552 17739 32555
rect 18322 32552 18328 32564
rect 17727 32524 18328 32552
rect 17727 32521 17739 32524
rect 17681 32515 17739 32521
rect 18322 32512 18328 32524
rect 18380 32512 18386 32564
rect 22646 32512 22652 32564
rect 22704 32552 22710 32564
rect 22833 32555 22891 32561
rect 22833 32552 22845 32555
rect 22704 32524 22845 32552
rect 22704 32512 22710 32524
rect 22833 32521 22845 32524
rect 22879 32521 22891 32555
rect 22833 32515 22891 32521
rect 27430 32512 27436 32564
rect 27488 32552 27494 32564
rect 29549 32555 29607 32561
rect 29549 32552 29561 32555
rect 27488 32524 29561 32552
rect 27488 32512 27494 32524
rect 29549 32521 29561 32524
rect 29595 32521 29607 32555
rect 29549 32515 29607 32521
rect 3050 32484 3056 32496
rect 2056 32456 3056 32484
rect 2056 32348 2084 32456
rect 3050 32444 3056 32456
rect 3108 32444 3114 32496
rect 3234 32484 3240 32496
rect 3195 32456 3240 32484
rect 3234 32444 3240 32456
rect 3292 32444 3298 32496
rect 4154 32444 4160 32496
rect 4212 32484 4218 32496
rect 4614 32484 4620 32496
rect 4212 32456 4620 32484
rect 4212 32444 4218 32456
rect 4614 32444 4620 32456
rect 4672 32484 4678 32496
rect 4982 32484 4988 32496
rect 4672 32456 4988 32484
rect 4672 32444 4678 32456
rect 4982 32444 4988 32456
rect 5040 32444 5046 32496
rect 7193 32487 7251 32493
rect 7193 32453 7205 32487
rect 7239 32484 7251 32487
rect 10962 32484 10968 32496
rect 7239 32456 10968 32484
rect 7239 32453 7251 32456
rect 7193 32447 7251 32453
rect 10962 32444 10968 32456
rect 11020 32484 11026 32496
rect 18966 32484 18972 32496
rect 11020 32456 11192 32484
rect 18927 32456 18972 32484
rect 11020 32444 11026 32456
rect 2958 32416 2964 32428
rect 2240 32388 2964 32416
rect 2133 32351 2191 32357
rect 2133 32348 2145 32351
rect 2056 32320 2145 32348
rect 2133 32317 2145 32320
rect 2179 32317 2191 32351
rect 2133 32311 2191 32317
rect 1949 32283 2007 32289
rect 1949 32249 1961 32283
rect 1995 32280 2007 32283
rect 2240 32280 2268 32388
rect 2958 32376 2964 32388
rect 3016 32376 3022 32428
rect 3068 32416 3096 32444
rect 4062 32416 4068 32428
rect 3068 32388 4068 32416
rect 4062 32376 4068 32388
rect 4120 32416 4126 32428
rect 6273 32419 6331 32425
rect 4120 32388 4476 32416
rect 4120 32376 4126 32388
rect 3326 32348 3332 32360
rect 2332 32320 3332 32348
rect 2332 32289 2360 32320
rect 3326 32308 3332 32320
rect 3384 32308 3390 32360
rect 3881 32351 3939 32357
rect 3881 32317 3893 32351
rect 3927 32317 3939 32351
rect 4154 32348 4160 32360
rect 4115 32320 4160 32348
rect 3881 32311 3939 32317
rect 1995 32252 2268 32280
rect 2317 32283 2375 32289
rect 1995 32249 2007 32252
rect 1949 32243 2007 32249
rect 2317 32249 2329 32283
rect 2363 32249 2375 32283
rect 2317 32243 2375 32249
rect 2685 32283 2743 32289
rect 2685 32249 2697 32283
rect 2731 32280 2743 32283
rect 3050 32280 3056 32292
rect 2731 32252 3056 32280
rect 2731 32249 2743 32252
rect 2685 32243 2743 32249
rect 3050 32240 3056 32252
rect 3108 32240 3114 32292
rect 3896 32280 3924 32311
rect 4154 32308 4160 32320
rect 4212 32308 4218 32360
rect 4448 32357 4476 32388
rect 6273 32385 6285 32419
rect 6319 32416 6331 32419
rect 6730 32416 6736 32428
rect 6319 32388 6736 32416
rect 6319 32385 6331 32388
rect 6273 32379 6331 32385
rect 6730 32376 6736 32388
rect 6788 32376 6794 32428
rect 7374 32376 7380 32428
rect 7432 32416 7438 32428
rect 9953 32419 10011 32425
rect 7432 32388 8616 32416
rect 7432 32376 7438 32388
rect 4433 32351 4491 32357
rect 4433 32317 4445 32351
rect 4479 32317 4491 32351
rect 5074 32348 5080 32360
rect 5035 32320 5080 32348
rect 4433 32311 4491 32317
rect 5074 32308 5080 32320
rect 5132 32308 5138 32360
rect 5718 32348 5724 32360
rect 5679 32320 5724 32348
rect 5718 32308 5724 32320
rect 5776 32308 5782 32360
rect 5813 32351 5871 32357
rect 5813 32317 5825 32351
rect 5859 32348 5871 32351
rect 6914 32348 6920 32360
rect 5859 32320 6920 32348
rect 5859 32317 5871 32320
rect 5813 32311 5871 32317
rect 6914 32308 6920 32320
rect 6972 32308 6978 32360
rect 7101 32351 7159 32357
rect 7101 32317 7113 32351
rect 7147 32348 7159 32351
rect 8294 32348 8300 32360
rect 7147 32320 8156 32348
rect 8255 32320 8300 32348
rect 7147 32317 7159 32320
rect 7101 32311 7159 32317
rect 4706 32280 4712 32292
rect 3896 32252 4712 32280
rect 4706 32240 4712 32252
rect 4764 32240 4770 32292
rect 5736 32280 5764 32308
rect 6546 32280 6552 32292
rect 5736 32252 6552 32280
rect 6546 32240 6552 32252
rect 6604 32240 6610 32292
rect 7282 32240 7288 32292
rect 7340 32280 7346 32292
rect 7745 32283 7803 32289
rect 7745 32280 7757 32283
rect 7340 32252 7757 32280
rect 7340 32240 7346 32252
rect 7745 32249 7757 32252
rect 7791 32249 7803 32283
rect 8128 32280 8156 32320
rect 8294 32308 8300 32320
rect 8352 32308 8358 32360
rect 8588 32357 8616 32388
rect 9953 32385 9965 32419
rect 9999 32416 10011 32419
rect 10226 32416 10232 32428
rect 9999 32388 10232 32416
rect 9999 32385 10011 32388
rect 9953 32379 10011 32385
rect 10226 32376 10232 32388
rect 10284 32376 10290 32428
rect 8573 32351 8631 32357
rect 8573 32317 8585 32351
rect 8619 32317 8631 32351
rect 8754 32348 8760 32360
rect 8715 32320 8760 32348
rect 8573 32311 8631 32317
rect 8754 32308 8760 32320
rect 8812 32308 8818 32360
rect 9858 32348 9864 32360
rect 9819 32320 9864 32348
rect 9858 32308 9864 32320
rect 9916 32308 9922 32360
rect 10321 32351 10379 32357
rect 10321 32317 10333 32351
rect 10367 32317 10379 32351
rect 10594 32348 10600 32360
rect 10555 32320 10600 32348
rect 10321 32311 10379 32317
rect 9490 32280 9496 32292
rect 8128 32252 9496 32280
rect 7745 32243 7803 32249
rect 9490 32240 9496 32252
rect 9548 32240 9554 32292
rect 9582 32240 9588 32292
rect 9640 32280 9646 32292
rect 10336 32280 10364 32311
rect 10594 32308 10600 32320
rect 10652 32308 10658 32360
rect 11054 32348 11060 32360
rect 11015 32320 11060 32348
rect 11054 32308 11060 32320
rect 11112 32308 11118 32360
rect 11164 32348 11192 32456
rect 18966 32444 18972 32456
rect 19024 32444 19030 32496
rect 28074 32484 28080 32496
rect 28035 32456 28080 32484
rect 28074 32444 28080 32456
rect 28132 32444 28138 32496
rect 32858 32444 32864 32496
rect 32916 32484 32922 32496
rect 34057 32487 34115 32493
rect 34057 32484 34069 32487
rect 32916 32456 34069 32484
rect 32916 32444 32922 32456
rect 34057 32453 34069 32456
rect 34103 32453 34115 32487
rect 34057 32447 34115 32453
rect 13170 32416 13176 32428
rect 13131 32388 13176 32416
rect 13170 32376 13176 32388
rect 13228 32376 13234 32428
rect 13446 32416 13452 32428
rect 13407 32388 13452 32416
rect 13446 32376 13452 32388
rect 13504 32376 13510 32428
rect 14550 32376 14556 32428
rect 14608 32416 14614 32428
rect 14608 32388 16436 32416
rect 14608 32376 14614 32388
rect 11241 32351 11299 32357
rect 11241 32348 11253 32351
rect 11164 32320 11253 32348
rect 11241 32317 11253 32320
rect 11287 32317 11299 32351
rect 11241 32311 11299 32317
rect 15102 32308 15108 32360
rect 15160 32348 15166 32360
rect 15657 32351 15715 32357
rect 15657 32348 15669 32351
rect 15160 32320 15669 32348
rect 15160 32308 15166 32320
rect 15657 32317 15669 32320
rect 15703 32317 15715 32351
rect 15657 32311 15715 32317
rect 15838 32308 15844 32360
rect 15896 32348 15902 32360
rect 16408 32357 16436 32388
rect 16666 32376 16672 32428
rect 16724 32416 16730 32428
rect 20438 32416 20444 32428
rect 16724 32388 18092 32416
rect 20399 32388 20444 32416
rect 16724 32376 16730 32388
rect 16025 32351 16083 32357
rect 16025 32348 16037 32351
rect 15896 32320 16037 32348
rect 15896 32308 15902 32320
rect 16025 32317 16037 32320
rect 16071 32317 16083 32351
rect 16025 32311 16083 32317
rect 16393 32351 16451 32357
rect 16393 32317 16405 32351
rect 16439 32317 16451 32351
rect 16393 32311 16451 32317
rect 17129 32351 17187 32357
rect 17129 32317 17141 32351
rect 17175 32348 17187 32351
rect 17494 32348 17500 32360
rect 17175 32320 17500 32348
rect 17175 32317 17187 32320
rect 17129 32311 17187 32317
rect 11422 32280 11428 32292
rect 9640 32252 11428 32280
rect 9640 32240 9646 32252
rect 11422 32240 11428 32252
rect 11480 32240 11486 32292
rect 14826 32280 14832 32292
rect 14787 32252 14832 32280
rect 14826 32240 14832 32252
rect 14884 32240 14890 32292
rect 16408 32280 16436 32311
rect 17494 32308 17500 32320
rect 17552 32308 17558 32360
rect 17865 32351 17923 32357
rect 17865 32317 17877 32351
rect 17911 32348 17923 32351
rect 17954 32348 17960 32360
rect 17911 32320 17960 32348
rect 17911 32317 17923 32320
rect 17865 32311 17923 32317
rect 17954 32308 17960 32320
rect 18012 32308 18018 32360
rect 18064 32357 18092 32388
rect 20438 32376 20444 32388
rect 20496 32376 20502 32428
rect 21082 32376 21088 32428
rect 21140 32416 21146 32428
rect 22557 32419 22615 32425
rect 22557 32416 22569 32419
rect 21140 32388 22569 32416
rect 21140 32376 21146 32388
rect 22557 32385 22569 32388
rect 22603 32385 22615 32419
rect 22557 32379 22615 32385
rect 23198 32376 23204 32428
rect 23256 32416 23262 32428
rect 23661 32419 23719 32425
rect 23661 32416 23673 32419
rect 23256 32388 23673 32416
rect 23256 32376 23262 32388
rect 23661 32385 23673 32388
rect 23707 32385 23719 32419
rect 23661 32379 23719 32385
rect 23937 32419 23995 32425
rect 23937 32385 23949 32419
rect 23983 32416 23995 32419
rect 25590 32416 25596 32428
rect 23983 32388 25596 32416
rect 23983 32385 23995 32388
rect 23937 32379 23995 32385
rect 18049 32351 18107 32357
rect 18049 32317 18061 32351
rect 18095 32317 18107 32351
rect 18506 32348 18512 32360
rect 18467 32320 18512 32348
rect 18049 32311 18107 32317
rect 18506 32308 18512 32320
rect 18564 32308 18570 32360
rect 18874 32348 18880 32360
rect 18835 32320 18880 32348
rect 18874 32308 18880 32320
rect 18932 32308 18938 32360
rect 20714 32348 20720 32360
rect 20675 32320 20720 32348
rect 20714 32308 20720 32320
rect 20772 32308 20778 32360
rect 22097 32351 22155 32357
rect 22097 32317 22109 32351
rect 22143 32348 22155 32351
rect 22649 32351 22707 32357
rect 22649 32348 22661 32351
rect 22143 32320 22661 32348
rect 22143 32317 22155 32320
rect 22097 32311 22155 32317
rect 22649 32317 22661 32320
rect 22695 32317 22707 32351
rect 23676 32348 23704 32379
rect 25590 32376 25596 32388
rect 25648 32376 25654 32428
rect 29270 32416 29276 32428
rect 29231 32388 29276 32416
rect 29270 32376 29276 32388
rect 29328 32376 29334 32428
rect 33321 32419 33379 32425
rect 33321 32385 33333 32419
rect 33367 32416 33379 32419
rect 33870 32416 33876 32428
rect 33367 32388 33876 32416
rect 33367 32385 33379 32388
rect 33321 32379 33379 32385
rect 33870 32376 33876 32388
rect 33928 32376 33934 32428
rect 25774 32348 25780 32360
rect 23676 32320 25780 32348
rect 22649 32311 22707 32317
rect 25774 32308 25780 32320
rect 25832 32308 25838 32360
rect 26050 32348 26056 32360
rect 26011 32320 26056 32348
rect 26050 32308 26056 32320
rect 26108 32308 26114 32360
rect 28261 32351 28319 32357
rect 28261 32317 28273 32351
rect 28307 32348 28319 32351
rect 28626 32348 28632 32360
rect 28307 32320 28632 32348
rect 28307 32317 28319 32320
rect 28261 32311 28319 32317
rect 28626 32308 28632 32320
rect 28684 32308 28690 32360
rect 28721 32351 28779 32357
rect 28721 32317 28733 32351
rect 28767 32348 28779 32351
rect 28810 32348 28816 32360
rect 28767 32320 28816 32348
rect 28767 32317 28779 32320
rect 28721 32311 28779 32317
rect 28810 32308 28816 32320
rect 28868 32308 28874 32360
rect 29365 32351 29423 32357
rect 29365 32317 29377 32351
rect 29411 32348 29423 32351
rect 30190 32348 30196 32360
rect 29411 32320 30196 32348
rect 29411 32317 29423 32320
rect 29365 32311 29423 32317
rect 30190 32308 30196 32320
rect 30248 32308 30254 32360
rect 30561 32351 30619 32357
rect 30561 32317 30573 32351
rect 30607 32317 30619 32351
rect 30834 32348 30840 32360
rect 30795 32320 30840 32348
rect 30561 32311 30619 32317
rect 17770 32280 17776 32292
rect 16408 32252 17776 32280
rect 17770 32240 17776 32252
rect 17828 32240 17834 32292
rect 2225 32215 2283 32221
rect 2225 32181 2237 32215
rect 2271 32212 2283 32215
rect 3142 32212 3148 32224
rect 2271 32184 3148 32212
rect 2271 32181 2283 32184
rect 2225 32175 2283 32181
rect 3142 32172 3148 32184
rect 3200 32172 3206 32224
rect 16206 32172 16212 32224
rect 16264 32212 16270 32224
rect 18506 32212 18512 32224
rect 16264 32184 18512 32212
rect 16264 32172 16270 32184
rect 18506 32172 18512 32184
rect 18564 32172 18570 32224
rect 24394 32172 24400 32224
rect 24452 32212 24458 32224
rect 25041 32215 25099 32221
rect 25041 32212 25053 32215
rect 24452 32184 25053 32212
rect 24452 32172 24458 32184
rect 25041 32181 25053 32184
rect 25087 32181 25099 32215
rect 27154 32212 27160 32224
rect 27115 32184 27160 32212
rect 25041 32175 25099 32181
rect 27154 32172 27160 32184
rect 27212 32172 27218 32224
rect 30576 32212 30604 32311
rect 30834 32308 30840 32320
rect 30892 32308 30898 32360
rect 32950 32348 32956 32360
rect 32911 32320 32956 32348
rect 32950 32308 32956 32320
rect 33008 32308 33014 32360
rect 33597 32351 33655 32357
rect 33597 32348 33609 32351
rect 33336 32320 33609 32348
rect 33336 32292 33364 32320
rect 33597 32317 33609 32320
rect 33643 32317 33655 32351
rect 33597 32311 33655 32317
rect 34149 32351 34207 32357
rect 34149 32317 34161 32351
rect 34195 32348 34207 32351
rect 34790 32348 34796 32360
rect 34195 32320 34796 32348
rect 34195 32317 34207 32320
rect 34149 32311 34207 32317
rect 34790 32308 34796 32320
rect 34848 32308 34854 32360
rect 35437 32351 35495 32357
rect 35437 32317 35449 32351
rect 35483 32348 35495 32351
rect 36078 32348 36084 32360
rect 35483 32320 36084 32348
rect 35483 32317 35495 32320
rect 35437 32311 35495 32317
rect 36078 32308 36084 32320
rect 36136 32308 36142 32360
rect 36262 32348 36268 32360
rect 36223 32320 36268 32348
rect 36262 32308 36268 32320
rect 36320 32308 36326 32360
rect 38654 32348 38660 32360
rect 38615 32320 38660 32348
rect 38654 32308 38660 32320
rect 38712 32308 38718 32360
rect 32214 32280 32220 32292
rect 32175 32252 32220 32280
rect 32214 32240 32220 32252
rect 32272 32240 32278 32292
rect 33318 32240 33324 32292
rect 33376 32240 33382 32292
rect 35253 32283 35311 32289
rect 35253 32249 35265 32283
rect 35299 32249 35311 32283
rect 35802 32280 35808 32292
rect 35763 32252 35808 32280
rect 35253 32243 35311 32249
rect 32122 32212 32128 32224
rect 30576 32184 32128 32212
rect 32122 32172 32128 32184
rect 32180 32212 32186 32224
rect 32769 32215 32827 32221
rect 32769 32212 32781 32215
rect 32180 32184 32781 32212
rect 32180 32172 32186 32184
rect 32769 32181 32781 32184
rect 32815 32212 32827 32215
rect 34514 32212 34520 32224
rect 32815 32184 34520 32212
rect 32815 32181 32827 32184
rect 32769 32175 32827 32181
rect 34514 32172 34520 32184
rect 34572 32172 34578 32224
rect 35268 32212 35296 32243
rect 35802 32240 35808 32252
rect 35860 32240 35866 32292
rect 36170 32212 36176 32224
rect 35268 32184 36176 32212
rect 36170 32172 36176 32184
rect 36228 32172 36234 32224
rect 36357 32215 36415 32221
rect 36357 32181 36369 32215
rect 36403 32212 36415 32215
rect 36538 32212 36544 32224
rect 36403 32184 36544 32212
rect 36403 32181 36415 32184
rect 36357 32175 36415 32181
rect 36538 32172 36544 32184
rect 36596 32172 36602 32224
rect 38746 32212 38752 32224
rect 38707 32184 38752 32212
rect 38746 32172 38752 32184
rect 38804 32172 38810 32224
rect 1104 32122 39836 32144
rect 1104 32070 19606 32122
rect 19658 32070 19670 32122
rect 19722 32070 19734 32122
rect 19786 32070 19798 32122
rect 19850 32070 39836 32122
rect 1104 32048 39836 32070
rect 1670 31968 1676 32020
rect 1728 32008 1734 32020
rect 2317 32011 2375 32017
rect 2317 32008 2329 32011
rect 1728 31980 2329 32008
rect 1728 31968 1734 31980
rect 2317 31977 2329 31980
rect 2363 31977 2375 32011
rect 2317 31971 2375 31977
rect 4062 31968 4068 32020
rect 4120 32008 4126 32020
rect 4249 32011 4307 32017
rect 4249 32008 4261 32011
rect 4120 31980 4261 32008
rect 4120 31968 4126 31980
rect 4249 31977 4261 31980
rect 4295 31977 4307 32011
rect 10594 32008 10600 32020
rect 4249 31971 4307 31977
rect 8864 31980 10600 32008
rect 7190 31940 7196 31952
rect 5552 31912 7196 31940
rect 2498 31872 2504 31884
rect 2459 31844 2504 31872
rect 2498 31832 2504 31844
rect 2556 31832 2562 31884
rect 3050 31872 3056 31884
rect 3011 31844 3056 31872
rect 3050 31832 3056 31844
rect 3108 31832 3114 31884
rect 3234 31872 3240 31884
rect 3195 31844 3240 31872
rect 3234 31832 3240 31844
rect 3292 31832 3298 31884
rect 4062 31872 4068 31884
rect 4023 31844 4068 31872
rect 4062 31832 4068 31844
rect 4120 31832 4126 31884
rect 5552 31881 5580 31912
rect 7190 31900 7196 31912
rect 7248 31900 7254 31952
rect 8754 31940 8760 31952
rect 7852 31912 8760 31940
rect 5537 31875 5595 31881
rect 5537 31841 5549 31875
rect 5583 31841 5595 31875
rect 5537 31835 5595 31841
rect 6641 31875 6699 31881
rect 6641 31841 6653 31875
rect 6687 31841 6699 31875
rect 6641 31835 6699 31841
rect 7101 31875 7159 31881
rect 7101 31841 7113 31875
rect 7147 31872 7159 31875
rect 7282 31872 7288 31884
rect 7147 31844 7288 31872
rect 7147 31841 7159 31844
rect 7101 31835 7159 31841
rect 6656 31804 6684 31835
rect 7282 31832 7288 31844
rect 7340 31832 7346 31884
rect 7852 31881 7880 31912
rect 8754 31900 8760 31912
rect 8812 31900 8818 31952
rect 7837 31875 7895 31881
rect 7837 31841 7849 31875
rect 7883 31841 7895 31875
rect 8202 31872 8208 31884
rect 8163 31844 8208 31872
rect 7837 31835 7895 31841
rect 8202 31832 8208 31844
rect 8260 31832 8266 31884
rect 8573 31875 8631 31881
rect 8573 31841 8585 31875
rect 8619 31872 8631 31875
rect 8864 31872 8892 31980
rect 10594 31968 10600 31980
rect 10652 31968 10658 32020
rect 11054 31968 11060 32020
rect 11112 32008 11118 32020
rect 11241 32011 11299 32017
rect 11241 32008 11253 32011
rect 11112 31980 11253 32008
rect 11112 31968 11118 31980
rect 11241 31977 11253 31980
rect 11287 31977 11299 32011
rect 11241 31971 11299 31977
rect 13081 32011 13139 32017
rect 13081 31977 13093 32011
rect 13127 32008 13139 32011
rect 13630 32008 13636 32020
rect 13127 31980 13636 32008
rect 13127 31977 13139 31980
rect 13081 31971 13139 31977
rect 13630 31968 13636 31980
rect 13688 31968 13694 32020
rect 14458 31968 14464 32020
rect 14516 32008 14522 32020
rect 15381 32011 15439 32017
rect 15381 32008 15393 32011
rect 14516 31980 15393 32008
rect 14516 31968 14522 31980
rect 15381 31977 15393 31980
rect 15427 31977 15439 32011
rect 15381 31971 15439 31977
rect 17696 31980 18828 32008
rect 13906 31940 13912 31952
rect 13740 31912 13912 31940
rect 8619 31844 8892 31872
rect 9033 31875 9091 31881
rect 8619 31841 8631 31844
rect 8573 31835 8631 31841
rect 9033 31841 9045 31875
rect 9079 31872 9091 31875
rect 9582 31872 9588 31884
rect 9079 31844 9588 31872
rect 9079 31841 9091 31844
rect 9033 31835 9091 31841
rect 9582 31832 9588 31844
rect 9640 31832 9646 31884
rect 9674 31832 9680 31884
rect 9732 31872 9738 31884
rect 10137 31875 10195 31881
rect 10137 31872 10149 31875
rect 9732 31844 10149 31872
rect 9732 31832 9738 31844
rect 10137 31841 10149 31844
rect 10183 31841 10195 31875
rect 10137 31835 10195 31841
rect 11977 31875 12035 31881
rect 11977 31841 11989 31875
rect 12023 31872 12035 31875
rect 12250 31872 12256 31884
rect 12023 31844 12256 31872
rect 12023 31841 12035 31844
rect 11977 31835 12035 31841
rect 12250 31832 12256 31844
rect 12308 31832 12314 31884
rect 12986 31872 12992 31884
rect 12947 31844 12992 31872
rect 12986 31832 12992 31844
rect 13044 31832 13050 31884
rect 13630 31832 13636 31884
rect 13688 31872 13694 31884
rect 13740 31881 13768 31912
rect 13906 31900 13912 31912
rect 13964 31940 13970 31952
rect 13964 31912 16068 31940
rect 13964 31900 13970 31912
rect 13725 31875 13783 31881
rect 13725 31872 13737 31875
rect 13688 31844 13737 31872
rect 13688 31832 13694 31844
rect 13725 31841 13737 31844
rect 13771 31841 13783 31875
rect 13998 31872 14004 31884
rect 13959 31844 14004 31872
rect 13725 31835 13783 31841
rect 13998 31832 14004 31844
rect 14056 31832 14062 31884
rect 14553 31875 14611 31881
rect 14553 31841 14565 31875
rect 14599 31872 14611 31875
rect 15194 31872 15200 31884
rect 14599 31844 15200 31872
rect 14599 31841 14611 31844
rect 14553 31835 14611 31841
rect 15194 31832 15200 31844
rect 15252 31832 15258 31884
rect 15473 31875 15531 31881
rect 15473 31841 15485 31875
rect 15519 31872 15531 31875
rect 15838 31872 15844 31884
rect 15519 31844 15844 31872
rect 15519 31841 15531 31844
rect 15473 31835 15531 31841
rect 15838 31832 15844 31844
rect 15896 31832 15902 31884
rect 16040 31881 16068 31912
rect 16114 31900 16120 31952
rect 16172 31940 16178 31952
rect 16853 31943 16911 31949
rect 16853 31940 16865 31943
rect 16172 31912 16865 31940
rect 16172 31900 16178 31912
rect 16853 31909 16865 31912
rect 16899 31909 16911 31943
rect 16853 31903 16911 31909
rect 16025 31875 16083 31881
rect 16025 31841 16037 31875
rect 16071 31872 16083 31875
rect 16206 31872 16212 31884
rect 16071 31844 16212 31872
rect 16071 31841 16083 31844
rect 16025 31835 16083 31841
rect 16206 31832 16212 31844
rect 16264 31832 16270 31884
rect 16390 31832 16396 31884
rect 16448 31872 16454 31884
rect 17696 31881 17724 31980
rect 18509 31943 18567 31949
rect 18509 31940 18521 31943
rect 17972 31912 18521 31940
rect 17681 31875 17739 31881
rect 17681 31872 17693 31875
rect 16448 31844 17693 31872
rect 16448 31832 16454 31844
rect 17681 31841 17693 31844
rect 17727 31841 17739 31875
rect 17862 31872 17868 31884
rect 17823 31844 17868 31872
rect 17681 31835 17739 31841
rect 17862 31832 17868 31844
rect 17920 31832 17926 31884
rect 7653 31807 7711 31813
rect 7653 31804 7665 31807
rect 6656 31776 7665 31804
rect 7653 31773 7665 31776
rect 7699 31773 7711 31807
rect 7653 31767 7711 31773
rect 9861 31807 9919 31813
rect 9861 31773 9873 31807
rect 9907 31804 9919 31807
rect 10042 31804 10048 31816
rect 9907 31776 10048 31804
rect 9907 31773 9919 31776
rect 9861 31767 9919 31773
rect 10042 31764 10048 31776
rect 10100 31764 10106 31816
rect 11330 31764 11336 31816
rect 11388 31804 11394 31816
rect 12069 31807 12127 31813
rect 12069 31804 12081 31807
rect 11388 31776 12081 31804
rect 11388 31764 11394 31776
rect 12069 31773 12081 31776
rect 12115 31773 12127 31807
rect 14016 31804 14044 31832
rect 15102 31804 15108 31816
rect 14016 31776 15108 31804
rect 12069 31767 12127 31773
rect 15102 31764 15108 31776
rect 15160 31804 15166 31816
rect 16117 31807 16175 31813
rect 16117 31804 16129 31807
rect 15160 31776 16129 31804
rect 15160 31764 15166 31776
rect 16117 31773 16129 31776
rect 16163 31773 16175 31807
rect 16117 31767 16175 31773
rect 17218 31764 17224 31816
rect 17276 31804 17282 31816
rect 17405 31807 17463 31813
rect 17405 31804 17417 31807
rect 17276 31776 17417 31804
rect 17276 31764 17282 31776
rect 17405 31773 17417 31776
rect 17451 31773 17463 31807
rect 17405 31767 17463 31773
rect 17494 31764 17500 31816
rect 17552 31804 17558 31816
rect 17880 31804 17908 31832
rect 17552 31776 17908 31804
rect 17552 31764 17558 31776
rect 5994 31696 6000 31748
rect 6052 31736 6058 31748
rect 6052 31708 9904 31736
rect 6052 31696 6058 31708
rect 9876 31680 9904 31708
rect 15838 31696 15844 31748
rect 15896 31736 15902 31748
rect 17972 31736 18000 31912
rect 18509 31909 18521 31912
rect 18555 31909 18567 31943
rect 18509 31903 18567 31909
rect 18693 31943 18751 31949
rect 18693 31909 18705 31943
rect 18739 31909 18751 31943
rect 18800 31940 18828 31980
rect 18874 31968 18880 32020
rect 18932 32008 18938 32020
rect 19613 32011 19671 32017
rect 19613 32008 19625 32011
rect 18932 31980 19625 32008
rect 18932 31968 18938 31980
rect 19613 31977 19625 31980
rect 19659 31977 19671 32011
rect 19613 31971 19671 31977
rect 25774 31968 25780 32020
rect 25832 32008 25838 32020
rect 26881 32011 26939 32017
rect 26881 32008 26893 32011
rect 25832 31980 26893 32008
rect 25832 31968 25838 31980
rect 26881 31977 26893 31980
rect 26927 32008 26939 32011
rect 27246 32008 27252 32020
rect 26927 31980 27252 32008
rect 26927 31977 26939 31980
rect 26881 31971 26939 31977
rect 27246 31968 27252 31980
rect 27304 31968 27310 32020
rect 31113 32011 31171 32017
rect 31113 31977 31125 32011
rect 31159 31977 31171 32011
rect 31113 31971 31171 31977
rect 19061 31943 19119 31949
rect 19061 31940 19073 31943
rect 18800 31912 19073 31940
rect 18693 31903 18751 31909
rect 19061 31909 19073 31912
rect 19107 31909 19119 31943
rect 27338 31940 27344 31952
rect 19061 31903 19119 31909
rect 25148 31912 27344 31940
rect 18598 31872 18604 31884
rect 18559 31844 18604 31872
rect 18598 31832 18604 31844
rect 18656 31832 18662 31884
rect 18708 31872 18736 31903
rect 19150 31872 19156 31884
rect 18708 31844 19156 31872
rect 19150 31832 19156 31844
rect 19208 31872 19214 31884
rect 19521 31875 19579 31881
rect 19521 31872 19533 31875
rect 19208 31844 19533 31872
rect 19208 31832 19214 31844
rect 19521 31841 19533 31844
rect 19567 31841 19579 31875
rect 19521 31835 19579 31841
rect 19981 31875 20039 31881
rect 19981 31841 19993 31875
rect 20027 31841 20039 31875
rect 19981 31835 20039 31841
rect 20993 31875 21051 31881
rect 20993 31841 21005 31875
rect 21039 31872 21051 31875
rect 21450 31872 21456 31884
rect 21039 31844 21456 31872
rect 21039 31841 21051 31844
rect 20993 31835 21051 31841
rect 18322 31804 18328 31816
rect 18235 31776 18328 31804
rect 18322 31764 18328 31776
rect 18380 31804 18386 31816
rect 18380 31776 18405 31804
rect 18380 31764 18386 31776
rect 15896 31708 18000 31736
rect 18340 31736 18368 31764
rect 19996 31736 20024 31835
rect 21450 31832 21456 31844
rect 21508 31872 21514 31884
rect 21545 31875 21603 31881
rect 21545 31872 21557 31875
rect 21508 31844 21557 31872
rect 21508 31832 21514 31844
rect 21545 31841 21557 31844
rect 21591 31841 21603 31875
rect 22646 31872 22652 31884
rect 22607 31844 22652 31872
rect 21545 31835 21603 31841
rect 22646 31832 22652 31844
rect 22704 31832 22710 31884
rect 25148 31881 25176 31912
rect 27338 31900 27344 31912
rect 27396 31900 27402 31952
rect 31128 31940 31156 31971
rect 33686 31968 33692 32020
rect 33744 32008 33750 32020
rect 33744 31980 37872 32008
rect 33744 31968 33750 31980
rect 30300 31912 31156 31940
rect 33781 31943 33839 31949
rect 30300 31884 30328 31912
rect 33781 31909 33793 31943
rect 33827 31940 33839 31943
rect 33870 31940 33876 31952
rect 33827 31912 33876 31940
rect 33827 31909 33839 31912
rect 33781 31903 33839 31909
rect 33870 31900 33876 31912
rect 33928 31900 33934 31952
rect 36170 31900 36176 31952
rect 36228 31940 36234 31952
rect 37090 31940 37096 31952
rect 36228 31912 37096 31940
rect 36228 31900 36234 31912
rect 37090 31900 37096 31912
rect 37148 31940 37154 31952
rect 37148 31912 37780 31940
rect 37148 31900 37154 31912
rect 25133 31875 25191 31881
rect 25133 31841 25145 31875
rect 25179 31841 25191 31875
rect 25685 31875 25743 31881
rect 25685 31872 25697 31875
rect 25133 31835 25191 31841
rect 25240 31844 25697 31872
rect 20901 31807 20959 31813
rect 20901 31773 20913 31807
rect 20947 31804 20959 31807
rect 21082 31804 21088 31816
rect 20947 31776 21088 31804
rect 20947 31773 20959 31776
rect 20901 31767 20959 31773
rect 21082 31764 21088 31776
rect 21140 31764 21146 31816
rect 22373 31807 22431 31813
rect 22373 31773 22385 31807
rect 22419 31773 22431 31807
rect 22373 31767 22431 31773
rect 18340 31708 20024 31736
rect 15896 31696 15902 31708
rect 20438 31696 20444 31748
rect 20496 31736 20502 31748
rect 22388 31736 22416 31767
rect 23474 31764 23480 31816
rect 23532 31804 23538 31816
rect 24394 31804 24400 31816
rect 23532 31776 24400 31804
rect 23532 31764 23538 31776
rect 24394 31764 24400 31776
rect 24452 31764 24458 31816
rect 24670 31764 24676 31816
rect 24728 31804 24734 31816
rect 25240 31804 25268 31844
rect 25685 31841 25697 31844
rect 25731 31841 25743 31875
rect 25685 31835 25743 31841
rect 27065 31875 27123 31881
rect 27065 31841 27077 31875
rect 27111 31841 27123 31875
rect 27065 31835 27123 31841
rect 24728 31776 25268 31804
rect 25501 31807 25559 31813
rect 24728 31764 24734 31776
rect 25501 31773 25513 31807
rect 25547 31804 25559 31807
rect 26050 31804 26056 31816
rect 25547 31776 26056 31804
rect 25547 31773 25559 31776
rect 25501 31767 25559 31773
rect 26050 31764 26056 31776
rect 26108 31764 26114 31816
rect 20496 31708 22416 31736
rect 20496 31696 20502 31708
rect 5626 31668 5632 31680
rect 5587 31640 5632 31668
rect 5626 31628 5632 31640
rect 5684 31628 5690 31680
rect 6086 31628 6092 31680
rect 6144 31668 6150 31680
rect 6457 31671 6515 31677
rect 6457 31668 6469 31671
rect 6144 31640 6469 31668
rect 6144 31628 6150 31640
rect 6457 31637 6469 31640
rect 6503 31637 6515 31671
rect 6457 31631 6515 31637
rect 9858 31628 9864 31680
rect 9916 31628 9922 31680
rect 14642 31668 14648 31680
rect 14603 31640 14648 31668
rect 14642 31628 14648 31640
rect 14700 31628 14706 31680
rect 20714 31628 20720 31680
rect 20772 31668 20778 31680
rect 21177 31671 21235 31677
rect 21177 31668 21189 31671
rect 20772 31640 21189 31668
rect 20772 31628 20778 31640
rect 21177 31637 21189 31640
rect 21223 31637 21235 31671
rect 21177 31631 21235 31637
rect 23937 31671 23995 31677
rect 23937 31637 23949 31671
rect 23983 31668 23995 31671
rect 24026 31668 24032 31680
rect 23983 31640 24032 31668
rect 23983 31637 23995 31640
rect 23937 31631 23995 31637
rect 24026 31628 24032 31640
rect 24084 31628 24090 31680
rect 27080 31668 27108 31835
rect 27154 31832 27160 31884
rect 27212 31872 27218 31884
rect 29365 31875 29423 31881
rect 29365 31872 29377 31875
rect 27212 31844 29377 31872
rect 27212 31832 27218 31844
rect 29365 31841 29377 31844
rect 29411 31841 29423 31875
rect 29365 31835 29423 31841
rect 29917 31875 29975 31881
rect 29917 31841 29929 31875
rect 29963 31872 29975 31875
rect 30006 31872 30012 31884
rect 29963 31844 30012 31872
rect 29963 31841 29975 31844
rect 29917 31835 29975 31841
rect 30006 31832 30012 31844
rect 30064 31832 30070 31884
rect 30282 31872 30288 31884
rect 30195 31844 30288 31872
rect 30282 31832 30288 31844
rect 30340 31832 30346 31884
rect 30929 31875 30987 31881
rect 30929 31872 30941 31875
rect 30392 31844 30941 31872
rect 27246 31804 27252 31816
rect 27207 31776 27252 31804
rect 27246 31764 27252 31776
rect 27304 31764 27310 31816
rect 27525 31807 27583 31813
rect 27525 31773 27537 31807
rect 27571 31804 27583 31807
rect 27614 31804 27620 31816
rect 27571 31776 27620 31804
rect 27571 31773 27583 31776
rect 27525 31767 27583 31773
rect 27614 31764 27620 31776
rect 27672 31764 27678 31816
rect 28905 31807 28963 31813
rect 28905 31773 28917 31807
rect 28951 31804 28963 31807
rect 29454 31804 29460 31816
rect 28951 31776 29460 31804
rect 28951 31773 28963 31776
rect 28905 31767 28963 31773
rect 29454 31764 29460 31776
rect 29512 31764 29518 31816
rect 29546 31764 29552 31816
rect 29604 31804 29610 31816
rect 30392 31804 30420 31844
rect 30929 31841 30941 31844
rect 30975 31841 30987 31875
rect 32122 31872 32128 31884
rect 32083 31844 32128 31872
rect 30929 31835 30987 31841
rect 32122 31832 32128 31844
rect 32180 31832 32186 31884
rect 32398 31872 32404 31884
rect 32359 31844 32404 31872
rect 32398 31832 32404 31844
rect 32456 31832 32462 31884
rect 34514 31872 34520 31884
rect 34427 31844 34520 31872
rect 34514 31832 34520 31844
rect 34572 31872 34578 31884
rect 36630 31872 36636 31884
rect 34572 31844 34928 31872
rect 36591 31844 36636 31872
rect 34572 31832 34578 31844
rect 29604 31776 30420 31804
rect 29604 31764 29610 31776
rect 34698 31764 34704 31816
rect 34756 31804 34762 31816
rect 34793 31807 34851 31813
rect 34793 31804 34805 31807
rect 34756 31776 34805 31804
rect 34756 31764 34762 31776
rect 34793 31773 34805 31776
rect 34839 31773 34851 31807
rect 34900 31804 34928 31844
rect 36630 31832 36636 31844
rect 36688 31832 36694 31884
rect 37752 31881 37780 31912
rect 37737 31875 37795 31881
rect 37737 31841 37749 31875
rect 37783 31841 37795 31875
rect 37844 31872 37872 31980
rect 38749 31875 38807 31881
rect 38749 31872 38761 31875
rect 37844 31844 38761 31872
rect 37737 31835 37795 31841
rect 38749 31841 38761 31844
rect 38795 31841 38807 31875
rect 38749 31835 38807 31841
rect 36814 31804 36820 31816
rect 34900 31776 36820 31804
rect 34793 31767 34851 31773
rect 36814 31764 36820 31776
rect 36872 31764 36878 31816
rect 30285 31739 30343 31745
rect 30285 31705 30297 31739
rect 30331 31736 30343 31739
rect 30466 31736 30472 31748
rect 30331 31708 30472 31736
rect 30331 31705 30343 31708
rect 30285 31699 30343 31705
rect 30466 31696 30472 31708
rect 30524 31696 30530 31748
rect 28442 31668 28448 31680
rect 27080 31640 28448 31668
rect 28442 31628 28448 31640
rect 28500 31628 28506 31680
rect 36078 31668 36084 31680
rect 36039 31640 36084 31668
rect 36078 31628 36084 31640
rect 36136 31628 36142 31680
rect 36722 31668 36728 31680
rect 36683 31640 36728 31668
rect 36722 31628 36728 31640
rect 36780 31628 36786 31680
rect 37921 31671 37979 31677
rect 37921 31637 37933 31671
rect 37967 31668 37979 31671
rect 38010 31668 38016 31680
rect 37967 31640 38016 31668
rect 37967 31637 37979 31640
rect 37921 31631 37979 31637
rect 38010 31628 38016 31640
rect 38068 31628 38074 31680
rect 38930 31668 38936 31680
rect 38891 31640 38936 31668
rect 38930 31628 38936 31640
rect 38988 31628 38994 31680
rect 1104 31578 39836 31600
rect 1104 31526 4246 31578
rect 4298 31526 4310 31578
rect 4362 31526 4374 31578
rect 4426 31526 4438 31578
rect 4490 31526 34966 31578
rect 35018 31526 35030 31578
rect 35082 31526 35094 31578
rect 35146 31526 35158 31578
rect 35210 31526 39836 31578
rect 1104 31504 39836 31526
rect 2866 31424 2872 31476
rect 2924 31464 2930 31476
rect 2961 31467 3019 31473
rect 2961 31464 2973 31467
rect 2924 31436 2973 31464
rect 2924 31424 2930 31436
rect 2961 31433 2973 31436
rect 3007 31464 3019 31467
rect 4062 31464 4068 31476
rect 3007 31436 4068 31464
rect 3007 31433 3019 31436
rect 2961 31427 3019 31433
rect 4062 31424 4068 31436
rect 4120 31424 4126 31476
rect 9490 31464 9496 31476
rect 9451 31436 9496 31464
rect 9490 31424 9496 31436
rect 9548 31424 9554 31476
rect 15102 31424 15108 31476
rect 15160 31464 15166 31476
rect 17405 31467 17463 31473
rect 17405 31464 17417 31467
rect 15160 31436 17417 31464
rect 15160 31424 15166 31436
rect 17405 31433 17417 31436
rect 17451 31433 17463 31467
rect 17405 31427 17463 31433
rect 18325 31467 18383 31473
rect 18325 31433 18337 31467
rect 18371 31464 18383 31467
rect 18506 31464 18512 31476
rect 18371 31436 18512 31464
rect 18371 31433 18383 31436
rect 18325 31427 18383 31433
rect 18506 31424 18512 31436
rect 18564 31424 18570 31476
rect 27338 31464 27344 31476
rect 27299 31436 27344 31464
rect 27338 31424 27344 31436
rect 27396 31424 27402 31476
rect 31128 31436 33180 31464
rect 9858 31356 9864 31408
rect 9916 31396 9922 31408
rect 12437 31399 12495 31405
rect 12437 31396 12449 31399
rect 9916 31368 12449 31396
rect 9916 31356 9922 31368
rect 12437 31365 12449 31368
rect 12483 31365 12495 31399
rect 12437 31359 12495 31365
rect 12529 31399 12587 31405
rect 12529 31365 12541 31399
rect 12575 31365 12587 31399
rect 12529 31359 12587 31365
rect 20533 31399 20591 31405
rect 20533 31365 20545 31399
rect 20579 31365 20591 31399
rect 20533 31359 20591 31365
rect 22465 31399 22523 31405
rect 22465 31365 22477 31399
rect 22511 31396 22523 31399
rect 23474 31396 23480 31408
rect 22511 31368 23480 31396
rect 22511 31365 22523 31368
rect 22465 31359 22523 31365
rect 1397 31331 1455 31337
rect 1397 31297 1409 31331
rect 1443 31328 1455 31331
rect 2682 31328 2688 31340
rect 1443 31300 2688 31328
rect 1443 31297 1455 31300
rect 1397 31291 1455 31297
rect 2682 31288 2688 31300
rect 2740 31288 2746 31340
rect 4614 31328 4620 31340
rect 4264 31300 4620 31328
rect 1670 31260 1676 31272
rect 1631 31232 1676 31260
rect 1670 31220 1676 31232
rect 1728 31220 1734 31272
rect 3697 31263 3755 31269
rect 3697 31229 3709 31263
rect 3743 31260 3755 31263
rect 3970 31260 3976 31272
rect 3743 31232 3976 31260
rect 3743 31229 3755 31232
rect 3697 31223 3755 31229
rect 3970 31220 3976 31232
rect 4028 31220 4034 31272
rect 4264 31269 4292 31300
rect 4614 31288 4620 31300
rect 4672 31288 4678 31340
rect 6181 31331 6239 31337
rect 6181 31297 6193 31331
rect 6227 31328 6239 31331
rect 7561 31331 7619 31337
rect 7561 31328 7573 31331
rect 6227 31300 7573 31328
rect 6227 31297 6239 31300
rect 6181 31291 6239 31297
rect 7561 31297 7573 31300
rect 7607 31297 7619 31331
rect 7561 31291 7619 31297
rect 8202 31288 8208 31340
rect 8260 31328 8266 31340
rect 11425 31331 11483 31337
rect 8260 31300 9996 31328
rect 8260 31288 8266 31300
rect 4249 31263 4307 31269
rect 4249 31229 4261 31263
rect 4295 31229 4307 31263
rect 4249 31223 4307 31229
rect 4525 31263 4583 31269
rect 4525 31229 4537 31263
rect 4571 31260 4583 31263
rect 4706 31260 4712 31272
rect 4571 31232 4712 31260
rect 4571 31229 4583 31232
rect 4525 31223 4583 31229
rect 4706 31220 4712 31232
rect 4764 31260 4770 31272
rect 4890 31260 4896 31272
rect 4764 31232 4896 31260
rect 4764 31220 4770 31232
rect 4890 31220 4896 31232
rect 4948 31220 4954 31272
rect 5445 31263 5503 31269
rect 5445 31229 5457 31263
rect 5491 31229 5503 31263
rect 6086 31260 6092 31272
rect 6047 31232 6092 31260
rect 5445 31223 5503 31229
rect 5460 31192 5488 31223
rect 6086 31220 6092 31232
rect 6144 31220 6150 31272
rect 6454 31220 6460 31272
rect 6512 31260 6518 31272
rect 7285 31263 7343 31269
rect 7285 31260 7297 31263
rect 6512 31232 7297 31260
rect 6512 31220 6518 31232
rect 7285 31229 7297 31232
rect 7331 31229 7343 31263
rect 7285 31223 7343 31229
rect 8754 31220 8760 31272
rect 8812 31260 8818 31272
rect 9968 31269 9996 31300
rect 11425 31297 11437 31331
rect 11471 31328 11483 31331
rect 12544 31328 12572 31359
rect 11471 31300 12572 31328
rect 16025 31331 16083 31337
rect 11471 31297 11483 31300
rect 11425 31291 11483 31297
rect 16025 31297 16037 31331
rect 16071 31328 16083 31331
rect 18322 31328 18328 31340
rect 16071 31300 18328 31328
rect 16071 31297 16083 31300
rect 16025 31291 16083 31297
rect 18322 31288 18328 31300
rect 18380 31288 18386 31340
rect 19426 31288 19432 31340
rect 19484 31328 19490 31340
rect 19797 31331 19855 31337
rect 19797 31328 19809 31331
rect 19484 31300 19809 31328
rect 19484 31288 19490 31300
rect 19797 31297 19809 31300
rect 19843 31328 19855 31331
rect 20548 31328 20576 31359
rect 23474 31356 23480 31368
rect 23532 31356 23538 31408
rect 23566 31356 23572 31408
rect 23624 31396 23630 31408
rect 23937 31399 23995 31405
rect 23937 31396 23949 31399
rect 23624 31368 23949 31396
rect 23624 31356 23630 31368
rect 23937 31365 23949 31368
rect 23983 31396 23995 31399
rect 24210 31396 24216 31408
rect 23983 31368 24216 31396
rect 23983 31365 23995 31368
rect 23937 31359 23995 31365
rect 24210 31356 24216 31368
rect 24268 31356 24274 31408
rect 27706 31356 27712 31408
rect 27764 31396 27770 31408
rect 29365 31399 29423 31405
rect 29365 31396 29377 31399
rect 27764 31368 29377 31396
rect 27764 31356 27770 31368
rect 29365 31365 29377 31368
rect 29411 31365 29423 31399
rect 29365 31359 29423 31365
rect 30745 31399 30803 31405
rect 30745 31365 30757 31399
rect 30791 31396 30803 31399
rect 30834 31396 30840 31408
rect 30791 31368 30840 31396
rect 30791 31365 30803 31368
rect 30745 31359 30803 31365
rect 30834 31356 30840 31368
rect 30892 31356 30898 31408
rect 24305 31331 24363 31337
rect 24305 31328 24317 31331
rect 19843 31300 20576 31328
rect 22388 31300 24317 31328
rect 19843 31297 19855 31300
rect 19797 31291 19855 31297
rect 8941 31263 8999 31269
rect 8941 31260 8953 31263
rect 8812 31232 8953 31260
rect 8812 31220 8818 31232
rect 8941 31229 8953 31232
rect 8987 31260 8999 31263
rect 9401 31263 9459 31269
rect 9401 31260 9413 31263
rect 8987 31232 9413 31260
rect 8987 31229 8999 31232
rect 8941 31223 8999 31229
rect 9401 31229 9413 31232
rect 9447 31229 9459 31263
rect 9401 31223 9459 31229
rect 9953 31263 10011 31269
rect 9953 31229 9965 31263
rect 9999 31229 10011 31263
rect 9953 31223 10011 31229
rect 11701 31263 11759 31269
rect 11701 31229 11713 31263
rect 11747 31229 11759 31263
rect 11701 31223 11759 31229
rect 11885 31263 11943 31269
rect 11885 31229 11897 31263
rect 11931 31260 11943 31263
rect 12894 31260 12900 31272
rect 11931 31232 12900 31260
rect 11931 31229 11943 31232
rect 11885 31223 11943 31229
rect 7374 31192 7380 31204
rect 5460 31164 7380 31192
rect 7374 31152 7380 31164
rect 7432 31152 7438 31204
rect 10870 31192 10876 31204
rect 10831 31164 10876 31192
rect 10870 31152 10876 31164
rect 10928 31152 10934 31204
rect 3234 31084 3240 31136
rect 3292 31124 3298 31136
rect 3605 31127 3663 31133
rect 3605 31124 3617 31127
rect 3292 31096 3617 31124
rect 3292 31084 3298 31096
rect 3605 31093 3617 31096
rect 3651 31093 3663 31127
rect 3605 31087 3663 31093
rect 5537 31127 5595 31133
rect 5537 31093 5549 31127
rect 5583 31124 5595 31127
rect 5810 31124 5816 31136
rect 5583 31096 5816 31124
rect 5583 31093 5595 31096
rect 5537 31087 5595 31093
rect 5810 31084 5816 31096
rect 5868 31084 5874 31136
rect 11716 31124 11744 31223
rect 12894 31220 12900 31232
rect 12952 31220 12958 31272
rect 13630 31260 13636 31272
rect 13591 31232 13636 31260
rect 13630 31220 13636 31232
rect 13688 31220 13694 31272
rect 13909 31263 13967 31269
rect 13909 31229 13921 31263
rect 13955 31260 13967 31263
rect 13998 31260 14004 31272
rect 13955 31232 14004 31260
rect 13955 31229 13967 31232
rect 13909 31223 13967 31229
rect 13998 31220 14004 31232
rect 14056 31220 14062 31272
rect 14369 31263 14427 31269
rect 14369 31229 14381 31263
rect 14415 31260 14427 31263
rect 14642 31260 14648 31272
rect 14415 31232 14648 31260
rect 14415 31229 14427 31232
rect 14369 31223 14427 31229
rect 14642 31220 14648 31232
rect 14700 31220 14706 31272
rect 15105 31263 15163 31269
rect 15105 31229 15117 31263
rect 15151 31229 15163 31263
rect 15105 31223 15163 31229
rect 15197 31263 15255 31269
rect 15197 31229 15209 31263
rect 15243 31260 15255 31263
rect 15378 31260 15384 31272
rect 15243 31232 15384 31260
rect 15243 31229 15255 31232
rect 15197 31223 15255 31229
rect 15120 31192 15148 31223
rect 15378 31220 15384 31232
rect 15436 31220 15442 31272
rect 15562 31260 15568 31272
rect 15523 31232 15568 31260
rect 15562 31220 15568 31232
rect 15620 31220 15626 31272
rect 15654 31220 15660 31272
rect 15712 31260 15718 31272
rect 16209 31263 16267 31269
rect 16209 31260 16221 31263
rect 15712 31232 16221 31260
rect 15712 31220 15718 31232
rect 16209 31229 16221 31232
rect 16255 31260 16267 31263
rect 17221 31263 17279 31269
rect 17221 31260 17233 31263
rect 16255 31232 17233 31260
rect 16255 31229 16267 31232
rect 16209 31223 16267 31229
rect 17221 31229 17233 31232
rect 17267 31260 17279 31263
rect 17267 31232 17448 31260
rect 17267 31229 17279 31232
rect 17221 31223 17279 31229
rect 15286 31192 15292 31204
rect 15120 31164 15292 31192
rect 15286 31152 15292 31164
rect 15344 31152 15350 31204
rect 16393 31195 16451 31201
rect 16393 31192 16405 31195
rect 15396 31164 16405 31192
rect 13354 31124 13360 31136
rect 11716 31096 13360 31124
rect 13354 31084 13360 31096
rect 13412 31084 13418 31136
rect 14642 31084 14648 31136
rect 14700 31124 14706 31136
rect 15396 31124 15424 31164
rect 16393 31161 16405 31164
rect 16439 31161 16451 31195
rect 16393 31155 16451 31161
rect 16761 31195 16819 31201
rect 16761 31161 16773 31195
rect 16807 31192 16819 31195
rect 17310 31192 17316 31204
rect 16807 31164 17316 31192
rect 16807 31161 16819 31164
rect 16761 31155 16819 31161
rect 17310 31152 17316 31164
rect 17368 31152 17374 31204
rect 17420 31192 17448 31232
rect 17770 31220 17776 31272
rect 17828 31260 17834 31272
rect 18141 31263 18199 31269
rect 18141 31260 18153 31263
rect 17828 31232 18153 31260
rect 17828 31220 17834 31232
rect 18141 31229 18153 31232
rect 18187 31229 18199 31263
rect 19150 31260 19156 31272
rect 19111 31232 19156 31260
rect 18141 31223 18199 31229
rect 19150 31220 19156 31232
rect 19208 31220 19214 31272
rect 19705 31263 19763 31269
rect 19705 31229 19717 31263
rect 19751 31260 19763 31263
rect 19886 31260 19892 31272
rect 19751 31232 19892 31260
rect 19751 31229 19763 31232
rect 19705 31223 19763 31229
rect 19886 31220 19892 31232
rect 19944 31220 19950 31272
rect 20438 31260 20444 31272
rect 20399 31232 20444 31260
rect 20438 31220 20444 31232
rect 20496 31220 20502 31272
rect 21177 31263 21235 31269
rect 21177 31229 21189 31263
rect 21223 31229 21235 31263
rect 21634 31260 21640 31272
rect 21595 31232 21640 31260
rect 21177 31223 21235 31229
rect 18598 31192 18604 31204
rect 17420 31164 18604 31192
rect 18598 31152 18604 31164
rect 18656 31152 18662 31204
rect 21192 31192 21220 31223
rect 21634 31220 21640 31232
rect 21692 31220 21698 31272
rect 22388 31269 22416 31300
rect 24305 31297 24317 31300
rect 24351 31297 24363 31331
rect 24305 31291 24363 31297
rect 26804 31300 28028 31328
rect 22373 31263 22431 31269
rect 22373 31229 22385 31263
rect 22419 31229 22431 31263
rect 22373 31223 22431 31229
rect 22649 31263 22707 31269
rect 22649 31229 22661 31263
rect 22695 31260 22707 31263
rect 23566 31260 23572 31272
rect 22695 31232 23572 31260
rect 22695 31229 22707 31232
rect 22649 31223 22707 31229
rect 23566 31220 23572 31232
rect 23624 31220 23630 31272
rect 23845 31263 23903 31269
rect 23845 31229 23857 31263
rect 23891 31229 23903 31263
rect 23845 31223 23903 31229
rect 22554 31192 22560 31204
rect 21192 31164 22560 31192
rect 22554 31152 22560 31164
rect 22612 31152 22618 31204
rect 23860 31192 23888 31223
rect 24026 31220 24032 31272
rect 24084 31260 24090 31272
rect 24121 31263 24179 31269
rect 24121 31260 24133 31263
rect 24084 31232 24133 31260
rect 24084 31220 24090 31232
rect 24121 31229 24133 31232
rect 24167 31229 24179 31263
rect 26234 31260 26240 31272
rect 26195 31232 26240 31260
rect 24121 31223 24179 31229
rect 26234 31220 26240 31232
rect 26292 31220 26298 31272
rect 26418 31260 26424 31272
rect 26379 31232 26424 31260
rect 26418 31220 26424 31232
rect 26476 31220 26482 31272
rect 26804 31269 26832 31300
rect 26789 31263 26847 31269
rect 26789 31229 26801 31263
rect 26835 31229 26847 31263
rect 26789 31223 26847 31229
rect 27154 31220 27160 31272
rect 27212 31260 27218 31272
rect 28000 31269 28028 31300
rect 27249 31263 27307 31269
rect 27249 31260 27261 31263
rect 27212 31232 27261 31260
rect 27212 31220 27218 31232
rect 27249 31229 27261 31232
rect 27295 31229 27307 31263
rect 27249 31223 27307 31229
rect 27985 31263 28043 31269
rect 27985 31229 27997 31263
rect 28031 31229 28043 31263
rect 27985 31223 28043 31229
rect 28629 31263 28687 31269
rect 28629 31229 28641 31263
rect 28675 31260 28687 31263
rect 28994 31260 29000 31272
rect 28675 31232 29000 31260
rect 28675 31229 28687 31232
rect 28629 31223 28687 31229
rect 27890 31192 27896 31204
rect 23860 31164 27896 31192
rect 27890 31152 27896 31164
rect 27948 31152 27954 31204
rect 28000 31192 28028 31223
rect 28994 31220 29000 31232
rect 29052 31220 29058 31272
rect 29454 31260 29460 31272
rect 29415 31232 29460 31260
rect 29454 31220 29460 31232
rect 29512 31220 29518 31272
rect 29825 31263 29883 31269
rect 29825 31229 29837 31263
rect 29871 31229 29883 31263
rect 30466 31260 30472 31272
rect 30427 31232 30472 31260
rect 29825 31223 29883 31229
rect 28534 31192 28540 31204
rect 28000 31164 28540 31192
rect 28534 31152 28540 31164
rect 28592 31192 28598 31204
rect 28810 31192 28816 31204
rect 28592 31164 28816 31192
rect 28592 31152 28598 31164
rect 28810 31152 28816 31164
rect 28868 31192 28874 31204
rect 29840 31192 29868 31223
rect 30466 31220 30472 31232
rect 30524 31220 30530 31272
rect 31128 31269 31156 31436
rect 33152 31405 33180 31436
rect 34790 31424 34796 31476
rect 34848 31464 34854 31476
rect 36725 31467 36783 31473
rect 36725 31464 36737 31467
rect 34848 31436 36737 31464
rect 34848 31424 34854 31436
rect 36725 31433 36737 31436
rect 36771 31433 36783 31467
rect 36725 31427 36783 31433
rect 33137 31399 33195 31405
rect 33137 31365 33149 31399
rect 33183 31365 33195 31399
rect 33137 31359 33195 31365
rect 34882 31356 34888 31408
rect 34940 31396 34946 31408
rect 35713 31399 35771 31405
rect 35713 31396 35725 31399
rect 34940 31368 35725 31396
rect 34940 31356 34946 31368
rect 35713 31365 35725 31368
rect 35759 31365 35771 31399
rect 35713 31359 35771 31365
rect 33318 31328 33324 31340
rect 33060 31300 33324 31328
rect 31113 31263 31171 31269
rect 31113 31229 31125 31263
rect 31159 31229 31171 31263
rect 31113 31223 31171 31229
rect 31481 31263 31539 31269
rect 31481 31229 31493 31263
rect 31527 31260 31539 31263
rect 31570 31260 31576 31272
rect 31527 31232 31576 31260
rect 31527 31229 31539 31232
rect 31481 31223 31539 31229
rect 31570 31220 31576 31232
rect 31628 31220 31634 31272
rect 32214 31220 32220 31272
rect 32272 31260 32278 31272
rect 32401 31263 32459 31269
rect 32401 31260 32413 31263
rect 32272 31232 32413 31260
rect 32272 31220 32278 31232
rect 32401 31229 32413 31232
rect 32447 31229 32459 31263
rect 32401 31223 32459 31229
rect 32769 31263 32827 31269
rect 32769 31229 32781 31263
rect 32815 31260 32827 31263
rect 33060 31260 33088 31300
rect 33318 31288 33324 31300
rect 33376 31288 33382 31340
rect 32815 31232 33088 31260
rect 33137 31263 33195 31269
rect 32815 31229 32827 31232
rect 32769 31223 32827 31229
rect 33137 31229 33149 31263
rect 33183 31260 33195 31263
rect 33226 31260 33232 31272
rect 33183 31232 33232 31260
rect 33183 31229 33195 31232
rect 33137 31223 33195 31229
rect 28868 31164 29868 31192
rect 32416 31192 32444 31223
rect 33226 31220 33232 31232
rect 33284 31220 33290 31272
rect 33965 31263 34023 31269
rect 33965 31260 33977 31263
rect 33336 31232 33977 31260
rect 33336 31192 33364 31232
rect 33965 31229 33977 31232
rect 34011 31229 34023 31263
rect 33965 31223 34023 31229
rect 34790 31220 34796 31272
rect 34848 31260 34854 31272
rect 34885 31263 34943 31269
rect 34885 31260 34897 31263
rect 34848 31232 34897 31260
rect 34848 31220 34854 31232
rect 34885 31229 34897 31232
rect 34931 31229 34943 31263
rect 34885 31223 34943 31229
rect 35253 31263 35311 31269
rect 35253 31229 35265 31263
rect 35299 31229 35311 31263
rect 35802 31260 35808 31272
rect 35763 31232 35808 31260
rect 35253 31223 35311 31229
rect 32416 31164 33364 31192
rect 28868 31152 28874 31164
rect 33594 31152 33600 31204
rect 33652 31192 33658 31204
rect 33778 31192 33784 31204
rect 33652 31164 33784 31192
rect 33652 31152 33658 31164
rect 33778 31152 33784 31164
rect 33836 31192 33842 31204
rect 35268 31192 35296 31223
rect 35802 31220 35808 31232
rect 35860 31220 35866 31272
rect 36078 31220 36084 31272
rect 36136 31260 36142 31272
rect 36633 31263 36691 31269
rect 36633 31260 36645 31263
rect 36136 31232 36645 31260
rect 36136 31220 36142 31232
rect 36633 31229 36645 31232
rect 36679 31229 36691 31263
rect 36633 31223 36691 31229
rect 36814 31220 36820 31272
rect 36872 31260 36878 31272
rect 37461 31263 37519 31269
rect 37461 31260 37473 31263
rect 36872 31232 37473 31260
rect 36872 31220 36878 31232
rect 37461 31229 37473 31232
rect 37507 31229 37519 31263
rect 37734 31260 37740 31272
rect 37695 31232 37740 31260
rect 37461 31223 37519 31229
rect 37734 31220 37740 31232
rect 37792 31220 37798 31272
rect 33836 31164 35296 31192
rect 33836 31152 33842 31164
rect 35894 31152 35900 31204
rect 35952 31192 35958 31204
rect 36449 31195 36507 31201
rect 36449 31192 36461 31195
rect 35952 31164 36461 31192
rect 35952 31152 35958 31164
rect 36449 31161 36461 31164
rect 36495 31161 36507 31195
rect 36449 31155 36507 31161
rect 14700 31096 15424 31124
rect 16301 31127 16359 31133
rect 14700 31084 14706 31096
rect 16301 31093 16313 31127
rect 16347 31124 16359 31127
rect 18046 31124 18052 31136
rect 16347 31096 18052 31124
rect 16347 31093 16359 31096
rect 16301 31087 16359 31093
rect 18046 31084 18052 31096
rect 18104 31084 18110 31136
rect 18322 31084 18328 31136
rect 18380 31124 18386 31136
rect 18969 31127 19027 31133
rect 18969 31124 18981 31127
rect 18380 31096 18981 31124
rect 18380 31084 18386 31096
rect 18969 31093 18981 31096
rect 19015 31093 19027 31127
rect 18969 31087 19027 31093
rect 21542 31084 21548 31136
rect 21600 31124 21606 31136
rect 21729 31127 21787 31133
rect 21729 31124 21741 31127
rect 21600 31096 21741 31124
rect 21600 31084 21606 31096
rect 21729 31093 21741 31096
rect 21775 31093 21787 31127
rect 21729 31087 21787 31093
rect 22370 31084 22376 31136
rect 22428 31124 22434 31136
rect 22833 31127 22891 31133
rect 22833 31124 22845 31127
rect 22428 31096 22845 31124
rect 22428 31084 22434 31096
rect 22833 31093 22845 31096
rect 22879 31093 22891 31127
rect 28442 31124 28448 31136
rect 28355 31096 28448 31124
rect 22833 31087 22891 31093
rect 28442 31084 28448 31096
rect 28500 31124 28506 31136
rect 28902 31124 28908 31136
rect 28500 31096 28908 31124
rect 28500 31084 28506 31096
rect 28902 31084 28908 31096
rect 28960 31084 28966 31136
rect 33042 31084 33048 31136
rect 33100 31124 33106 31136
rect 34057 31127 34115 31133
rect 34057 31124 34069 31127
rect 33100 31096 34069 31124
rect 33100 31084 33106 31096
rect 34057 31093 34069 31096
rect 34103 31093 34115 31127
rect 34057 31087 34115 31093
rect 38654 31084 38660 31136
rect 38712 31124 38718 31136
rect 38841 31127 38899 31133
rect 38841 31124 38853 31127
rect 38712 31096 38853 31124
rect 38712 31084 38718 31096
rect 38841 31093 38853 31096
rect 38887 31093 38899 31127
rect 38841 31087 38899 31093
rect 1104 31034 39836 31056
rect 1104 30982 19606 31034
rect 19658 30982 19670 31034
rect 19722 30982 19734 31034
rect 19786 30982 19798 31034
rect 19850 30982 39836 31034
rect 1104 30960 39836 30982
rect 1670 30880 1676 30932
rect 1728 30920 1734 30932
rect 2501 30923 2559 30929
rect 2501 30920 2513 30923
rect 1728 30892 2513 30920
rect 1728 30880 1734 30892
rect 2501 30889 2513 30892
rect 2547 30889 2559 30923
rect 2501 30883 2559 30889
rect 17770 30880 17776 30932
rect 17828 30920 17834 30932
rect 18601 30923 18659 30929
rect 18601 30920 18613 30923
rect 17828 30892 18613 30920
rect 17828 30880 17834 30892
rect 18601 30889 18613 30892
rect 18647 30889 18659 30923
rect 18601 30883 18659 30889
rect 34241 30923 34299 30929
rect 34241 30889 34253 30923
rect 34287 30920 34299 30923
rect 34698 30920 34704 30932
rect 34287 30892 34704 30920
rect 34287 30889 34299 30892
rect 34241 30883 34299 30889
rect 34698 30880 34704 30892
rect 34756 30880 34762 30932
rect 2866 30852 2872 30864
rect 1780 30824 2872 30852
rect 1780 30793 1808 30824
rect 2866 30812 2872 30824
rect 2924 30812 2930 30864
rect 7190 30852 7196 30864
rect 7151 30824 7196 30852
rect 7190 30812 7196 30824
rect 7248 30812 7254 30864
rect 17494 30852 17500 30864
rect 17144 30824 17500 30852
rect 17144 30796 17172 30824
rect 17494 30812 17500 30824
rect 17552 30812 17558 30864
rect 30009 30855 30067 30861
rect 30009 30821 30021 30855
rect 30055 30852 30067 30855
rect 30374 30852 30380 30864
rect 30055 30824 30380 30852
rect 30055 30821 30067 30824
rect 30009 30815 30067 30821
rect 30374 30812 30380 30824
rect 30432 30812 30438 30864
rect 33318 30852 33324 30864
rect 32692 30824 33324 30852
rect 1765 30787 1823 30793
rect 1765 30753 1777 30787
rect 1811 30753 1823 30787
rect 2682 30784 2688 30796
rect 2643 30756 2688 30784
rect 1765 30747 1823 30753
rect 2682 30744 2688 30756
rect 2740 30744 2746 30796
rect 3234 30784 3240 30796
rect 3195 30756 3240 30784
rect 3234 30744 3240 30756
rect 3292 30744 3298 30796
rect 3421 30787 3479 30793
rect 3421 30753 3433 30787
rect 3467 30784 3479 30787
rect 3694 30784 3700 30796
rect 3467 30756 3700 30784
rect 3467 30753 3479 30756
rect 3421 30747 3479 30753
rect 3694 30744 3700 30756
rect 3752 30744 3758 30796
rect 4062 30784 4068 30796
rect 4023 30756 4068 30784
rect 4062 30744 4068 30756
rect 4120 30744 4126 30796
rect 5353 30787 5411 30793
rect 5353 30753 5365 30787
rect 5399 30784 5411 30787
rect 5626 30784 5632 30796
rect 5399 30756 5632 30784
rect 5399 30753 5411 30756
rect 5353 30747 5411 30753
rect 5626 30744 5632 30756
rect 5684 30744 5690 30796
rect 7650 30784 7656 30796
rect 7611 30756 7656 30784
rect 7650 30744 7656 30756
rect 7708 30744 7714 30796
rect 7834 30784 7840 30796
rect 7795 30756 7840 30784
rect 7834 30744 7840 30756
rect 7892 30744 7898 30796
rect 8021 30787 8079 30793
rect 8021 30753 8033 30787
rect 8067 30753 8079 30787
rect 8021 30747 8079 30753
rect 5074 30716 5080 30728
rect 5035 30688 5080 30716
rect 5074 30676 5080 30688
rect 5132 30676 5138 30728
rect 6733 30719 6791 30725
rect 6733 30685 6745 30719
rect 6779 30716 6791 30719
rect 7006 30716 7012 30728
rect 6779 30688 7012 30716
rect 6779 30685 6791 30688
rect 6733 30679 6791 30685
rect 7006 30676 7012 30688
rect 7064 30716 7070 30728
rect 8036 30716 8064 30747
rect 8386 30744 8392 30796
rect 8444 30784 8450 30796
rect 8665 30787 8723 30793
rect 8665 30784 8677 30787
rect 8444 30756 8677 30784
rect 8444 30744 8450 30756
rect 8665 30753 8677 30756
rect 8711 30784 8723 30787
rect 9677 30787 9735 30793
rect 9677 30784 9689 30787
rect 8711 30756 9689 30784
rect 8711 30753 8723 30756
rect 8665 30747 8723 30753
rect 9677 30753 9689 30756
rect 9723 30753 9735 30787
rect 10410 30784 10416 30796
rect 10371 30756 10416 30784
rect 9677 30747 9735 30753
rect 10410 30744 10416 30756
rect 10468 30744 10474 30796
rect 10870 30744 10876 30796
rect 10928 30784 10934 30796
rect 11977 30787 12035 30793
rect 11977 30784 11989 30787
rect 10928 30756 11989 30784
rect 10928 30744 10934 30756
rect 11977 30753 11989 30756
rect 12023 30753 12035 30787
rect 11977 30747 12035 30753
rect 13357 30787 13415 30793
rect 13357 30753 13369 30787
rect 13403 30784 13415 30787
rect 14093 30787 14151 30793
rect 14093 30784 14105 30787
rect 13403 30756 14105 30784
rect 13403 30753 13415 30756
rect 13357 30747 13415 30753
rect 14093 30753 14105 30756
rect 14139 30784 14151 30787
rect 14274 30784 14280 30796
rect 14139 30756 14280 30784
rect 14139 30753 14151 30756
rect 14093 30747 14151 30753
rect 14274 30744 14280 30756
rect 14332 30744 14338 30796
rect 14553 30787 14611 30793
rect 14553 30753 14565 30787
rect 14599 30753 14611 30787
rect 14553 30747 14611 30753
rect 7064 30688 8064 30716
rect 7064 30676 7070 30688
rect 11146 30676 11152 30728
rect 11204 30716 11210 30728
rect 11701 30719 11759 30725
rect 11701 30716 11713 30719
rect 11204 30688 11713 30716
rect 11204 30676 11210 30688
rect 11701 30685 11713 30688
rect 11747 30685 11759 30719
rect 14182 30716 14188 30728
rect 14143 30688 14188 30716
rect 11701 30679 11759 30685
rect 14182 30676 14188 30688
rect 14240 30676 14246 30728
rect 14568 30716 14596 30747
rect 14826 30744 14832 30796
rect 14884 30784 14890 30796
rect 15289 30787 15347 30793
rect 15289 30784 15301 30787
rect 14884 30756 15301 30784
rect 14884 30744 14890 30756
rect 15289 30753 15301 30756
rect 15335 30753 15347 30787
rect 15289 30747 15347 30753
rect 15838 30744 15844 30796
rect 15896 30784 15902 30796
rect 16206 30784 16212 30796
rect 15896 30756 16212 30784
rect 15896 30744 15902 30756
rect 16206 30744 16212 30756
rect 16264 30744 16270 30796
rect 16945 30787 17003 30793
rect 16945 30753 16957 30787
rect 16991 30784 17003 30787
rect 17126 30784 17132 30796
rect 16991 30756 17132 30784
rect 16991 30753 17003 30756
rect 16945 30747 17003 30753
rect 17126 30744 17132 30756
rect 17184 30744 17190 30796
rect 17310 30744 17316 30796
rect 17368 30784 17374 30796
rect 17405 30787 17463 30793
rect 17405 30784 17417 30787
rect 17368 30756 17417 30784
rect 17368 30744 17374 30756
rect 17405 30753 17417 30756
rect 17451 30753 17463 30787
rect 17405 30747 17463 30753
rect 17954 30744 17960 30796
rect 18012 30784 18018 30796
rect 18509 30787 18567 30793
rect 18509 30784 18521 30787
rect 18012 30756 18521 30784
rect 18012 30744 18018 30756
rect 18509 30753 18521 30756
rect 18555 30753 18567 30787
rect 19150 30784 19156 30796
rect 19111 30756 19156 30784
rect 18509 30747 18567 30753
rect 19150 30744 19156 30756
rect 19208 30744 19214 30796
rect 19426 30784 19432 30796
rect 19387 30756 19432 30784
rect 19426 30744 19432 30756
rect 19484 30744 19490 30796
rect 19886 30784 19892 30796
rect 19847 30756 19892 30784
rect 19886 30744 19892 30756
rect 19944 30744 19950 30796
rect 21542 30784 21548 30796
rect 21503 30756 21548 30784
rect 21542 30744 21548 30756
rect 21600 30744 21606 30796
rect 23658 30784 23664 30796
rect 23619 30756 23664 30784
rect 23658 30744 23664 30756
rect 23716 30744 23722 30796
rect 23937 30787 23995 30793
rect 23937 30784 23949 30787
rect 23768 30756 23949 30784
rect 15470 30716 15476 30728
rect 14568 30688 15476 30716
rect 15470 30676 15476 30688
rect 15528 30676 15534 30728
rect 18230 30676 18236 30728
rect 18288 30716 18294 30728
rect 21269 30719 21327 30725
rect 21269 30716 21281 30719
rect 18288 30688 21281 30716
rect 18288 30676 18294 30688
rect 21269 30685 21281 30688
rect 21315 30685 21327 30719
rect 21269 30679 21327 30685
rect 23014 30676 23020 30728
rect 23072 30716 23078 30728
rect 23768 30716 23796 30756
rect 23937 30753 23949 30756
rect 23983 30753 23995 30787
rect 24210 30784 24216 30796
rect 24171 30756 24216 30784
rect 23937 30747 23995 30753
rect 24210 30744 24216 30756
rect 24268 30744 24274 30796
rect 24578 30784 24584 30796
rect 24539 30756 24584 30784
rect 24578 30744 24584 30756
rect 24636 30744 24642 30796
rect 25314 30784 25320 30796
rect 25275 30756 25320 30784
rect 25314 30744 25320 30756
rect 25372 30744 25378 30796
rect 27157 30787 27215 30793
rect 27157 30784 27169 30787
rect 25424 30756 27169 30784
rect 23072 30688 23796 30716
rect 23845 30719 23903 30725
rect 23072 30676 23078 30688
rect 23845 30685 23857 30719
rect 23891 30716 23903 30719
rect 25424 30716 25452 30756
rect 27157 30753 27169 30756
rect 27203 30753 27215 30787
rect 27706 30784 27712 30796
rect 27667 30756 27712 30784
rect 27157 30747 27215 30753
rect 27706 30744 27712 30756
rect 27764 30744 27770 30796
rect 28166 30744 28172 30796
rect 28224 30784 28230 30796
rect 28813 30787 28871 30793
rect 28813 30784 28825 30787
rect 28224 30756 28825 30784
rect 28224 30744 28230 30756
rect 28813 30753 28825 30756
rect 28859 30753 28871 30787
rect 28813 30747 28871 30753
rect 29457 30787 29515 30793
rect 29457 30753 29469 30787
rect 29503 30753 29515 30787
rect 29457 30747 29515 30753
rect 29825 30787 29883 30793
rect 29825 30753 29837 30787
rect 29871 30784 29883 30787
rect 30282 30784 30288 30796
rect 29871 30756 30288 30784
rect 29871 30753 29883 30756
rect 29825 30747 29883 30753
rect 26878 30716 26884 30728
rect 23891 30688 25452 30716
rect 26839 30688 26884 30716
rect 23891 30685 23903 30688
rect 23845 30679 23903 30685
rect 26878 30676 26884 30688
rect 26936 30676 26942 30728
rect 26970 30676 26976 30728
rect 27028 30716 27034 30728
rect 28997 30719 29055 30725
rect 28997 30716 29009 30719
rect 27028 30688 29009 30716
rect 27028 30676 27034 30688
rect 28997 30685 29009 30688
rect 29043 30685 29055 30719
rect 29472 30716 29500 30747
rect 30282 30744 30288 30756
rect 30340 30744 30346 30796
rect 30558 30784 30564 30796
rect 30519 30756 30564 30784
rect 30558 30744 30564 30756
rect 30616 30744 30622 30796
rect 32692 30793 32720 30824
rect 33318 30812 33324 30824
rect 33376 30852 33382 30864
rect 33376 30824 36216 30852
rect 33376 30812 33382 30824
rect 31205 30787 31263 30793
rect 31205 30753 31217 30787
rect 31251 30784 31263 30787
rect 32677 30787 32735 30793
rect 31251 30756 32352 30784
rect 31251 30753 31263 30756
rect 31205 30747 31263 30753
rect 30006 30716 30012 30728
rect 29472 30688 30012 30716
rect 28997 30679 29055 30685
rect 30006 30676 30012 30688
rect 30064 30676 30070 30728
rect 31297 30719 31355 30725
rect 31297 30685 31309 30719
rect 31343 30685 31355 30719
rect 32214 30716 32220 30728
rect 32175 30688 32220 30716
rect 31297 30679 31355 30685
rect 7098 30608 7104 30660
rect 7156 30648 7162 30660
rect 7156 30620 11744 30648
rect 7156 30608 7162 30620
rect 11716 30592 11744 30620
rect 15194 30608 15200 30660
rect 15252 30648 15258 30660
rect 16301 30651 16359 30657
rect 16301 30648 16313 30651
rect 15252 30620 16313 30648
rect 15252 30608 15258 30620
rect 16301 30617 16313 30620
rect 16347 30617 16359 30651
rect 27614 30648 27620 30660
rect 27575 30620 27620 30648
rect 16301 30611 16359 30617
rect 27614 30608 27620 30620
rect 27672 30608 27678 30660
rect 30745 30651 30803 30657
rect 30745 30617 30757 30651
rect 30791 30648 30803 30651
rect 31110 30648 31116 30660
rect 30791 30620 31116 30648
rect 30791 30617 30803 30620
rect 30745 30611 30803 30617
rect 31110 30608 31116 30620
rect 31168 30608 31174 30660
rect 31312 30648 31340 30679
rect 32214 30676 32220 30688
rect 32272 30676 32278 30728
rect 32324 30716 32352 30756
rect 32677 30753 32689 30787
rect 32723 30753 32735 30787
rect 33042 30784 33048 30796
rect 33003 30756 33048 30784
rect 32677 30747 32735 30753
rect 33042 30744 33048 30756
rect 33100 30744 33106 30796
rect 33134 30744 33140 30796
rect 33192 30784 33198 30796
rect 34149 30787 34207 30793
rect 34149 30784 34161 30787
rect 33192 30756 34161 30784
rect 33192 30744 33198 30756
rect 34149 30753 34161 30756
rect 34195 30753 34207 30787
rect 34882 30784 34888 30796
rect 34843 30756 34888 30784
rect 34149 30747 34207 30753
rect 34882 30744 34888 30756
rect 34940 30744 34946 30796
rect 32953 30719 33011 30725
rect 32953 30716 32965 30719
rect 32324 30688 32965 30716
rect 32953 30685 32965 30688
rect 32999 30685 33011 30719
rect 32953 30679 33011 30685
rect 34238 30676 34244 30728
rect 34296 30716 34302 30728
rect 34977 30719 35035 30725
rect 34977 30716 34989 30719
rect 34296 30688 34989 30716
rect 34296 30676 34302 30688
rect 34977 30685 34989 30688
rect 35023 30685 35035 30719
rect 36078 30716 36084 30728
rect 36039 30688 36084 30716
rect 34977 30679 35035 30685
rect 36078 30676 36084 30688
rect 36136 30676 36142 30728
rect 36188 30716 36216 30824
rect 36633 30787 36691 30793
rect 36633 30753 36645 30787
rect 36679 30784 36691 30787
rect 36722 30784 36728 30796
rect 36679 30756 36728 30784
rect 36679 30753 36691 30756
rect 36633 30747 36691 30753
rect 36722 30744 36728 30756
rect 36780 30744 36786 30796
rect 36909 30787 36967 30793
rect 36909 30753 36921 30787
rect 36955 30784 36967 30787
rect 37458 30784 37464 30796
rect 36955 30756 37464 30784
rect 36955 30753 36967 30756
rect 36909 30747 36967 30753
rect 37458 30744 37464 30756
rect 37516 30784 37522 30796
rect 37737 30787 37795 30793
rect 37737 30784 37749 30787
rect 37516 30756 37749 30784
rect 37516 30744 37522 30756
rect 37737 30753 37749 30756
rect 37783 30753 37795 30787
rect 37737 30747 37795 30753
rect 37918 30744 37924 30796
rect 37976 30784 37982 30796
rect 38105 30787 38163 30793
rect 38105 30784 38117 30787
rect 37976 30756 38117 30784
rect 37976 30744 37982 30756
rect 38105 30753 38117 30756
rect 38151 30753 38163 30787
rect 38105 30747 38163 30753
rect 38473 30787 38531 30793
rect 38473 30753 38485 30787
rect 38519 30753 38531 30787
rect 38473 30747 38531 30753
rect 37093 30719 37151 30725
rect 37093 30716 37105 30719
rect 36188 30688 37105 30716
rect 37093 30685 37105 30688
rect 37139 30716 37151 30719
rect 38010 30716 38016 30728
rect 37139 30688 38016 30716
rect 37139 30685 37151 30688
rect 37093 30679 37151 30685
rect 38010 30676 38016 30688
rect 38068 30716 38074 30728
rect 38488 30716 38516 30747
rect 38838 30716 38844 30728
rect 38068 30688 38516 30716
rect 38799 30688 38844 30716
rect 38068 30676 38074 30688
rect 38838 30676 38844 30688
rect 38896 30676 38902 30728
rect 31312 30620 31432 30648
rect 1857 30583 1915 30589
rect 1857 30549 1869 30583
rect 1903 30580 1915 30583
rect 2774 30580 2780 30592
rect 1903 30552 2780 30580
rect 1903 30549 1915 30552
rect 1857 30543 1915 30549
rect 2774 30540 2780 30552
rect 2832 30540 2838 30592
rect 4249 30583 4307 30589
rect 4249 30549 4261 30583
rect 4295 30580 4307 30583
rect 4706 30580 4712 30592
rect 4295 30552 4712 30580
rect 4295 30549 4307 30552
rect 4249 30543 4307 30549
rect 4706 30540 4712 30552
rect 4764 30540 4770 30592
rect 8849 30583 8907 30589
rect 8849 30549 8861 30583
rect 8895 30580 8907 30583
rect 8938 30580 8944 30592
rect 8895 30552 8944 30580
rect 8895 30549 8907 30552
rect 8849 30543 8907 30549
rect 8938 30540 8944 30552
rect 8996 30580 9002 30592
rect 9214 30580 9220 30592
rect 8996 30552 9220 30580
rect 8996 30540 9002 30552
rect 9214 30540 9220 30552
rect 9272 30540 9278 30592
rect 9858 30580 9864 30592
rect 9819 30552 9864 30580
rect 9858 30540 9864 30552
rect 9916 30540 9922 30592
rect 10134 30540 10140 30592
rect 10192 30580 10198 30592
rect 10594 30580 10600 30592
rect 10192 30552 10600 30580
rect 10192 30540 10198 30552
rect 10594 30540 10600 30552
rect 10652 30540 10658 30592
rect 11698 30540 11704 30592
rect 11756 30540 11762 30592
rect 15473 30583 15531 30589
rect 15473 30549 15485 30583
rect 15519 30580 15531 30583
rect 15654 30580 15660 30592
rect 15519 30552 15660 30580
rect 15519 30549 15531 30552
rect 15473 30543 15531 30549
rect 15654 30540 15660 30552
rect 15712 30540 15718 30592
rect 16114 30540 16120 30592
rect 16172 30580 16178 30592
rect 17589 30583 17647 30589
rect 17589 30580 17601 30583
rect 16172 30552 17601 30580
rect 16172 30540 16178 30552
rect 17589 30549 17601 30552
rect 17635 30549 17647 30583
rect 22646 30580 22652 30592
rect 22607 30552 22652 30580
rect 17589 30543 17647 30549
rect 22646 30540 22652 30552
rect 22704 30540 22710 30592
rect 25409 30583 25467 30589
rect 25409 30549 25421 30583
rect 25455 30580 25467 30583
rect 25590 30580 25596 30592
rect 25455 30552 25596 30580
rect 25455 30549 25467 30552
rect 25409 30543 25467 30549
rect 25590 30540 25596 30552
rect 25648 30540 25654 30592
rect 28629 30583 28687 30589
rect 28629 30549 28641 30583
rect 28675 30580 28687 30583
rect 28994 30580 29000 30592
rect 28675 30552 29000 30580
rect 28675 30549 28687 30552
rect 28629 30543 28687 30549
rect 28994 30540 29000 30552
rect 29052 30580 29058 30592
rect 29270 30580 29276 30592
rect 29052 30552 29276 30580
rect 29052 30540 29058 30552
rect 29270 30540 29276 30552
rect 29328 30540 29334 30592
rect 31404 30580 31432 30620
rect 31570 30580 31576 30592
rect 31404 30552 31576 30580
rect 31570 30540 31576 30552
rect 31628 30580 31634 30592
rect 32766 30580 32772 30592
rect 31628 30552 32772 30580
rect 31628 30540 31634 30552
rect 32766 30540 32772 30552
rect 32824 30580 32830 30592
rect 34238 30580 34244 30592
rect 32824 30552 34244 30580
rect 32824 30540 32830 30552
rect 34238 30540 34244 30552
rect 34296 30540 34302 30592
rect 1104 30490 39836 30512
rect 1104 30438 4246 30490
rect 4298 30438 4310 30490
rect 4362 30438 4374 30490
rect 4426 30438 4438 30490
rect 4490 30438 34966 30490
rect 35018 30438 35030 30490
rect 35082 30438 35094 30490
rect 35146 30438 35158 30490
rect 35210 30438 39836 30490
rect 1104 30416 39836 30438
rect 9858 30336 9864 30388
rect 9916 30376 9922 30388
rect 10226 30376 10232 30388
rect 9916 30348 10232 30376
rect 9916 30336 9922 30348
rect 10226 30336 10232 30348
rect 10284 30336 10290 30388
rect 10410 30336 10416 30388
rect 10468 30376 10474 30388
rect 10962 30376 10968 30388
rect 10468 30348 10968 30376
rect 10468 30336 10474 30348
rect 10962 30336 10968 30348
rect 11020 30376 11026 30388
rect 11020 30348 11652 30376
rect 11020 30336 11026 30348
rect 3694 30308 3700 30320
rect 3655 30280 3700 30308
rect 3694 30268 3700 30280
rect 3752 30268 3758 30320
rect 7650 30308 7656 30320
rect 7611 30280 7656 30308
rect 7650 30268 7656 30280
rect 7708 30268 7714 30320
rect 9950 30268 9956 30320
rect 10008 30308 10014 30320
rect 10321 30311 10379 30317
rect 10321 30308 10333 30311
rect 10008 30280 10333 30308
rect 10008 30268 10014 30280
rect 10321 30277 10333 30280
rect 10367 30277 10379 30311
rect 10321 30271 10379 30277
rect 10594 30268 10600 30320
rect 10652 30308 10658 30320
rect 10652 30280 11560 30308
rect 10652 30268 10658 30280
rect 3160 30212 4568 30240
rect 1673 30175 1731 30181
rect 1673 30141 1685 30175
rect 1719 30141 1731 30175
rect 1673 30135 1731 30141
rect 1765 30175 1823 30181
rect 1765 30141 1777 30175
rect 1811 30172 1823 30175
rect 2406 30172 2412 30184
rect 1811 30144 2412 30172
rect 1811 30141 1823 30144
rect 1765 30135 1823 30141
rect 1688 30036 1716 30135
rect 2406 30132 2412 30144
rect 2464 30132 2470 30184
rect 2774 30132 2780 30184
rect 2832 30172 2838 30184
rect 2832 30144 2877 30172
rect 2832 30132 2838 30144
rect 3050 30132 3056 30184
rect 3108 30172 3114 30184
rect 3160 30181 3188 30212
rect 4540 30184 4568 30212
rect 4614 30200 4620 30252
rect 4672 30240 4678 30252
rect 4801 30243 4859 30249
rect 4801 30240 4813 30243
rect 4672 30212 4813 30240
rect 4672 30200 4678 30212
rect 4801 30209 4813 30212
rect 4847 30209 4859 30243
rect 4801 30203 4859 30209
rect 6273 30243 6331 30249
rect 6273 30209 6285 30243
rect 6319 30240 6331 30243
rect 7834 30240 7840 30252
rect 6319 30212 7840 30240
rect 6319 30209 6331 30212
rect 6273 30203 6331 30209
rect 3145 30175 3203 30181
rect 3145 30172 3157 30175
rect 3108 30144 3157 30172
rect 3108 30132 3114 30144
rect 3145 30141 3157 30144
rect 3191 30141 3203 30175
rect 3145 30135 3203 30141
rect 3234 30132 3240 30184
rect 3292 30172 3298 30184
rect 3513 30175 3571 30181
rect 3513 30172 3525 30175
rect 3292 30144 3525 30172
rect 3292 30132 3298 30144
rect 3513 30141 3525 30144
rect 3559 30172 3571 30175
rect 4062 30172 4068 30184
rect 3559 30144 4068 30172
rect 3559 30141 3571 30144
rect 3513 30135 3571 30141
rect 4062 30132 4068 30144
rect 4120 30132 4126 30184
rect 4522 30172 4528 30184
rect 4483 30144 4528 30172
rect 4522 30132 4528 30144
rect 4580 30132 4586 30184
rect 4706 30172 4712 30184
rect 4619 30144 4712 30172
rect 4706 30132 4712 30144
rect 4764 30172 4770 30184
rect 5810 30172 5816 30184
rect 4764 30144 5488 30172
rect 5771 30144 5816 30172
rect 4764 30132 4770 30144
rect 5460 30116 5488 30144
rect 5810 30132 5816 30144
rect 5868 30132 5874 30184
rect 5997 30175 6055 30181
rect 5997 30141 6009 30175
rect 6043 30141 6055 30175
rect 7006 30172 7012 30184
rect 6967 30144 7012 30172
rect 5997 30135 6055 30141
rect 5442 30064 5448 30116
rect 5500 30104 5506 30116
rect 6012 30104 6040 30135
rect 7006 30132 7012 30144
rect 7064 30132 7070 30184
rect 7208 30181 7236 30212
rect 7834 30200 7840 30212
rect 7892 30200 7898 30252
rect 8294 30240 8300 30252
rect 8207 30212 8300 30240
rect 7193 30175 7251 30181
rect 7193 30141 7205 30175
rect 7239 30141 7251 30175
rect 7193 30135 7251 30141
rect 7745 30175 7803 30181
rect 7745 30141 7757 30175
rect 7791 30172 7803 30175
rect 8220 30172 8248 30212
rect 8294 30200 8300 30212
rect 8352 30240 8358 30252
rect 8478 30240 8484 30252
rect 8352 30212 8484 30240
rect 8352 30200 8358 30212
rect 8478 30200 8484 30212
rect 8536 30240 8542 30252
rect 9582 30240 9588 30252
rect 8536 30212 9588 30240
rect 8536 30200 8542 30212
rect 9582 30200 9588 30212
rect 9640 30200 9646 30252
rect 9677 30243 9735 30249
rect 9677 30209 9689 30243
rect 9723 30240 9735 30243
rect 9723 30212 11376 30240
rect 9723 30209 9735 30212
rect 9677 30203 9735 30209
rect 11348 30184 11376 30212
rect 8386 30172 8392 30184
rect 7791 30144 8248 30172
rect 8347 30144 8392 30172
rect 7791 30141 7803 30144
rect 7745 30135 7803 30141
rect 8386 30132 8392 30144
rect 8444 30132 8450 30184
rect 9306 30172 9312 30184
rect 9267 30144 9312 30172
rect 9306 30132 9312 30144
rect 9364 30132 9370 30184
rect 10045 30175 10103 30181
rect 10045 30141 10057 30175
rect 10091 30172 10103 30175
rect 10134 30172 10140 30184
rect 10091 30144 10140 30172
rect 10091 30141 10103 30144
rect 10045 30135 10103 30141
rect 10134 30132 10140 30144
rect 10192 30132 10198 30184
rect 10226 30132 10232 30184
rect 10284 30172 10290 30184
rect 10321 30175 10379 30181
rect 10321 30172 10333 30175
rect 10284 30144 10333 30172
rect 10284 30132 10290 30144
rect 10321 30141 10333 30144
rect 10367 30141 10379 30175
rect 11330 30172 11336 30184
rect 11291 30144 11336 30172
rect 10321 30135 10379 30141
rect 11330 30132 11336 30144
rect 11388 30132 11394 30184
rect 11532 30181 11560 30280
rect 11624 30240 11652 30348
rect 11698 30336 11704 30388
rect 11756 30376 11762 30388
rect 12986 30376 12992 30388
rect 11756 30348 12992 30376
rect 11756 30336 11762 30348
rect 12986 30336 12992 30348
rect 13044 30336 13050 30388
rect 19334 30336 19340 30388
rect 19392 30376 19398 30388
rect 19613 30379 19671 30385
rect 19613 30376 19625 30379
rect 19392 30348 19625 30376
rect 19392 30336 19398 30348
rect 19613 30345 19625 30348
rect 19659 30376 19671 30379
rect 20438 30376 20444 30388
rect 19659 30348 20444 30376
rect 19659 30345 19671 30348
rect 19613 30339 19671 30345
rect 20438 30336 20444 30348
rect 20496 30336 20502 30388
rect 26234 30336 26240 30388
rect 26292 30376 26298 30388
rect 26513 30379 26571 30385
rect 26513 30376 26525 30379
rect 26292 30348 26525 30376
rect 26292 30336 26298 30348
rect 26513 30345 26525 30348
rect 26559 30376 26571 30379
rect 26970 30376 26976 30388
rect 26559 30348 26976 30376
rect 26559 30345 26571 30348
rect 26513 30339 26571 30345
rect 26970 30336 26976 30348
rect 27028 30336 27034 30388
rect 32030 30376 32036 30388
rect 30852 30348 32036 30376
rect 12434 30268 12440 30320
rect 12492 30308 12498 30320
rect 12529 30311 12587 30317
rect 12529 30308 12541 30311
rect 12492 30280 12541 30308
rect 12492 30268 12498 30280
rect 12529 30277 12541 30280
rect 12575 30277 12587 30311
rect 12529 30271 12587 30277
rect 17405 30311 17463 30317
rect 17405 30277 17417 30311
rect 17451 30308 17463 30311
rect 17954 30308 17960 30320
rect 17451 30280 17960 30308
rect 17451 30277 17463 30280
rect 17405 30271 17463 30277
rect 17954 30268 17960 30280
rect 18012 30268 18018 30320
rect 18046 30268 18052 30320
rect 18104 30268 18110 30320
rect 13725 30243 13783 30249
rect 13725 30240 13737 30243
rect 11624 30212 13737 30240
rect 13725 30209 13737 30212
rect 13771 30209 13783 30243
rect 13725 30203 13783 30209
rect 14826 30200 14832 30252
rect 14884 30240 14890 30252
rect 15562 30240 15568 30252
rect 14884 30212 14964 30240
rect 15523 30212 15568 30240
rect 14884 30200 14890 30212
rect 11517 30175 11575 30181
rect 11517 30141 11529 30175
rect 11563 30141 11575 30175
rect 12526 30172 12532 30184
rect 12487 30144 12532 30172
rect 11517 30135 11575 30141
rect 12526 30132 12532 30144
rect 12584 30132 12590 30184
rect 12989 30175 13047 30181
rect 12989 30141 13001 30175
rect 13035 30141 13047 30175
rect 13906 30172 13912 30184
rect 13867 30144 13912 30172
rect 12989 30135 13047 30141
rect 5500 30076 6040 30104
rect 5500 30064 5506 30076
rect 8294 30064 8300 30116
rect 8352 30104 8358 30116
rect 13004 30104 13032 30135
rect 13906 30132 13912 30144
rect 13964 30132 13970 30184
rect 14277 30175 14335 30181
rect 14277 30141 14289 30175
rect 14323 30141 14335 30175
rect 14458 30172 14464 30184
rect 14419 30144 14464 30172
rect 14277 30135 14335 30141
rect 8352 30076 13032 30104
rect 14292 30104 14320 30135
rect 14458 30132 14464 30144
rect 14516 30132 14522 30184
rect 14936 30181 14964 30212
rect 15562 30200 15568 30212
rect 15620 30200 15626 30252
rect 17218 30240 17224 30252
rect 16132 30212 17224 30240
rect 14921 30175 14979 30181
rect 14921 30141 14933 30175
rect 14967 30141 14979 30175
rect 14921 30135 14979 30141
rect 15838 30132 15844 30184
rect 15896 30172 15902 30184
rect 16132 30181 16160 30212
rect 17218 30200 17224 30212
rect 17276 30200 17282 30252
rect 18064 30240 18092 30268
rect 19242 30240 19248 30252
rect 17328 30212 19248 30240
rect 16117 30175 16175 30181
rect 16117 30172 16129 30175
rect 15896 30144 16129 30172
rect 15896 30132 15902 30144
rect 16117 30141 16129 30144
rect 16163 30141 16175 30175
rect 16390 30172 16396 30184
rect 16351 30144 16396 30172
rect 16117 30135 16175 30141
rect 16390 30132 16396 30144
rect 16448 30132 16454 30184
rect 16577 30175 16635 30181
rect 16577 30141 16589 30175
rect 16623 30172 16635 30175
rect 16758 30172 16764 30184
rect 16623 30144 16764 30172
rect 16623 30141 16635 30144
rect 16577 30135 16635 30141
rect 16758 30132 16764 30144
rect 16816 30132 16822 30184
rect 14642 30104 14648 30116
rect 14292 30076 14648 30104
rect 8352 30064 8358 30076
rect 14642 30064 14648 30076
rect 14700 30064 14706 30116
rect 17236 30104 17264 30200
rect 17328 30181 17356 30212
rect 19242 30200 19248 30212
rect 19300 30200 19306 30252
rect 19886 30200 19892 30252
rect 19944 30240 19950 30252
rect 19944 30212 21036 30240
rect 19944 30200 19950 30212
rect 17313 30175 17371 30181
rect 17313 30141 17325 30175
rect 17359 30141 17371 30175
rect 17313 30135 17371 30141
rect 17862 30132 17868 30184
rect 17920 30172 17926 30184
rect 18049 30175 18107 30181
rect 18049 30172 18061 30175
rect 17920 30144 18061 30172
rect 17920 30132 17926 30144
rect 18049 30141 18061 30144
rect 18095 30141 18107 30175
rect 18322 30172 18328 30184
rect 18283 30144 18328 30172
rect 18049 30135 18107 30141
rect 18322 30132 18328 30144
rect 18380 30132 18386 30184
rect 20162 30172 20168 30184
rect 20123 30144 20168 30172
rect 20162 30132 20168 30144
rect 20220 30132 20226 30184
rect 21008 30181 21036 30212
rect 21634 30200 21640 30252
rect 21692 30240 21698 30252
rect 21729 30243 21787 30249
rect 21729 30240 21741 30243
rect 21692 30212 21741 30240
rect 21692 30200 21698 30212
rect 21729 30209 21741 30212
rect 21775 30209 21787 30243
rect 21729 30203 21787 30209
rect 24949 30243 25007 30249
rect 24949 30209 24961 30243
rect 24995 30240 25007 30243
rect 26050 30240 26056 30252
rect 24995 30212 26056 30240
rect 24995 30209 25007 30212
rect 24949 30203 25007 30209
rect 26050 30200 26056 30212
rect 26108 30240 26114 30252
rect 27065 30243 27123 30249
rect 27065 30240 27077 30243
rect 26108 30212 27077 30240
rect 26108 30200 26114 30212
rect 27065 30209 27077 30212
rect 27111 30209 27123 30243
rect 29454 30240 29460 30252
rect 29415 30212 29460 30240
rect 27065 30203 27123 30209
rect 29454 30200 29460 30212
rect 29512 30200 29518 30252
rect 30852 30249 30880 30348
rect 32030 30336 32036 30348
rect 32088 30336 32094 30388
rect 32214 30376 32220 30388
rect 32175 30348 32220 30376
rect 32214 30336 32220 30348
rect 32272 30336 32278 30388
rect 37458 30376 37464 30388
rect 37419 30348 37464 30376
rect 37458 30336 37464 30348
rect 37516 30336 37522 30388
rect 35894 30268 35900 30320
rect 35952 30268 35958 30320
rect 37734 30268 37740 30320
rect 37792 30308 37798 30320
rect 38105 30311 38163 30317
rect 38105 30308 38117 30311
rect 37792 30280 38117 30308
rect 37792 30268 37798 30280
rect 38105 30277 38117 30280
rect 38151 30277 38163 30311
rect 38105 30271 38163 30277
rect 30837 30243 30895 30249
rect 30837 30209 30849 30243
rect 30883 30209 30895 30243
rect 31110 30240 31116 30252
rect 31071 30212 31116 30240
rect 30837 30203 30895 30209
rect 31110 30200 31116 30212
rect 31168 30200 31174 30252
rect 34238 30240 34244 30252
rect 34199 30212 34244 30240
rect 34238 30200 34244 30212
rect 34296 30200 34302 30252
rect 35912 30240 35940 30268
rect 34900 30212 35940 30240
rect 20625 30175 20683 30181
rect 20625 30141 20637 30175
rect 20671 30141 20683 30175
rect 20625 30135 20683 30141
rect 20993 30175 21051 30181
rect 20993 30141 21005 30175
rect 21039 30141 21051 30175
rect 20993 30135 21051 30141
rect 17236 30076 18092 30104
rect 3142 30036 3148 30048
rect 1688 30008 3148 30036
rect 3142 29996 3148 30008
rect 3200 29996 3206 30048
rect 8573 30039 8631 30045
rect 8573 30005 8585 30039
rect 8619 30036 8631 30039
rect 8754 30036 8760 30048
rect 8619 30008 8760 30036
rect 8619 30005 8631 30008
rect 8573 29999 8631 30005
rect 8754 29996 8760 30008
rect 8812 29996 8818 30048
rect 9122 30036 9128 30048
rect 9083 30008 9128 30036
rect 9122 29996 9128 30008
rect 9180 29996 9186 30048
rect 9214 29996 9220 30048
rect 9272 30036 9278 30048
rect 11149 30039 11207 30045
rect 11149 30036 11161 30039
rect 9272 30008 11161 30036
rect 9272 29996 9278 30008
rect 11149 30005 11161 30008
rect 11195 30005 11207 30039
rect 11149 29999 11207 30005
rect 13814 29996 13820 30048
rect 13872 30036 13878 30048
rect 17954 30036 17960 30048
rect 13872 30008 17960 30036
rect 13872 29996 13878 30008
rect 17954 29996 17960 30008
rect 18012 29996 18018 30048
rect 18064 30036 18092 30076
rect 19150 30064 19156 30116
rect 19208 30104 19214 30116
rect 20640 30104 20668 30135
rect 22002 30132 22008 30184
rect 22060 30172 22066 30184
rect 22189 30175 22247 30181
rect 22189 30172 22201 30175
rect 22060 30144 22201 30172
rect 22060 30132 22066 30144
rect 22189 30141 22201 30144
rect 22235 30141 22247 30175
rect 22189 30135 22247 30141
rect 22373 30175 22431 30181
rect 22373 30141 22385 30175
rect 22419 30141 22431 30175
rect 22373 30135 22431 30141
rect 22557 30175 22615 30181
rect 22557 30141 22569 30175
rect 22603 30172 22615 30175
rect 22646 30172 22652 30184
rect 22603 30144 22652 30172
rect 22603 30141 22615 30144
rect 22557 30135 22615 30141
rect 21266 30104 21272 30116
rect 19208 30076 20668 30104
rect 21179 30076 21272 30104
rect 19208 30064 19214 30076
rect 21266 30064 21272 30076
rect 21324 30104 21330 30116
rect 22388 30104 22416 30135
rect 22646 30132 22652 30144
rect 22704 30172 22710 30184
rect 23198 30172 23204 30184
rect 22704 30144 23204 30172
rect 22704 30132 22710 30144
rect 23198 30132 23204 30144
rect 23256 30132 23262 30184
rect 23934 30172 23940 30184
rect 23895 30144 23940 30172
rect 23934 30132 23940 30144
rect 23992 30132 23998 30184
rect 24121 30175 24179 30181
rect 24121 30141 24133 30175
rect 24167 30141 24179 30175
rect 25222 30172 25228 30184
rect 25183 30144 25228 30172
rect 24121 30135 24179 30141
rect 21324 30076 22416 30104
rect 21324 30064 21330 30076
rect 23290 30064 23296 30116
rect 23348 30104 23354 30116
rect 24136 30104 24164 30135
rect 25222 30132 25228 30144
rect 25280 30132 25286 30184
rect 27338 30172 27344 30184
rect 27299 30144 27344 30172
rect 27338 30132 27344 30144
rect 27396 30132 27402 30184
rect 29825 30175 29883 30181
rect 29825 30141 29837 30175
rect 29871 30172 29883 30175
rect 30006 30172 30012 30184
rect 29871 30144 30012 30172
rect 29871 30141 29883 30144
rect 29825 30135 29883 30141
rect 30006 30132 30012 30144
rect 30064 30132 30070 30184
rect 30193 30175 30251 30181
rect 30193 30141 30205 30175
rect 30239 30172 30251 30175
rect 30282 30172 30288 30184
rect 30239 30144 30288 30172
rect 30239 30141 30251 30144
rect 30193 30135 30251 30141
rect 30282 30132 30288 30144
rect 30340 30132 30346 30184
rect 30377 30175 30435 30181
rect 30377 30141 30389 30175
rect 30423 30172 30435 30175
rect 33134 30172 33140 30184
rect 30423 30144 33140 30172
rect 30423 30141 30435 30144
rect 30377 30135 30435 30141
rect 33134 30132 33140 30144
rect 33192 30132 33198 30184
rect 34900 30181 34928 30212
rect 36078 30200 36084 30252
rect 36136 30240 36142 30252
rect 36173 30243 36231 30249
rect 36173 30240 36185 30243
rect 36136 30212 36185 30240
rect 36136 30200 36142 30212
rect 36173 30209 36185 30212
rect 36219 30209 36231 30243
rect 38838 30240 38844 30252
rect 38799 30212 38844 30240
rect 36173 30203 36231 30209
rect 38838 30200 38844 30212
rect 38896 30200 38902 30252
rect 33229 30175 33287 30181
rect 33229 30141 33241 30175
rect 33275 30141 33287 30175
rect 33229 30135 33287 30141
rect 33965 30175 34023 30181
rect 33965 30141 33977 30175
rect 34011 30141 34023 30175
rect 33965 30135 34023 30141
rect 34885 30175 34943 30181
rect 34885 30141 34897 30175
rect 34931 30141 34943 30175
rect 34885 30135 34943 30141
rect 35069 30175 35127 30181
rect 35069 30141 35081 30175
rect 35115 30172 35127 30175
rect 35250 30172 35256 30184
rect 35115 30144 35256 30172
rect 35115 30141 35127 30144
rect 35069 30135 35127 30141
rect 28718 30104 28724 30116
rect 23348 30076 24164 30104
rect 28679 30076 28724 30104
rect 23348 30064 23354 30076
rect 28718 30064 28724 30076
rect 28776 30064 28782 30116
rect 32490 30064 32496 30116
rect 32548 30104 32554 30116
rect 33244 30104 33272 30135
rect 32548 30076 33272 30104
rect 33980 30104 34008 30135
rect 35250 30132 35256 30144
rect 35308 30132 35314 30184
rect 35897 30175 35955 30181
rect 35897 30141 35909 30175
rect 35943 30172 35955 30175
rect 36814 30172 36820 30184
rect 35943 30144 36820 30172
rect 35943 30141 35955 30144
rect 35897 30135 35955 30141
rect 36814 30132 36820 30144
rect 36872 30132 36878 30184
rect 38102 30172 38108 30184
rect 38063 30144 38108 30172
rect 38102 30132 38108 30144
rect 38160 30132 38166 30184
rect 38746 30172 38752 30184
rect 38707 30144 38752 30172
rect 38746 30132 38752 30144
rect 38804 30132 38810 30184
rect 34698 30104 34704 30116
rect 33980 30076 34704 30104
rect 32548 30064 32554 30076
rect 34698 30064 34704 30076
rect 34756 30064 34762 30116
rect 35437 30107 35495 30113
rect 35437 30073 35449 30107
rect 35483 30104 35495 30107
rect 35710 30104 35716 30116
rect 35483 30076 35716 30104
rect 35483 30073 35495 30076
rect 35437 30067 35495 30073
rect 35710 30064 35716 30076
rect 35768 30064 35774 30116
rect 21726 30036 21732 30048
rect 18064 30008 21732 30036
rect 21726 29996 21732 30008
rect 21784 29996 21790 30048
rect 23658 29996 23664 30048
rect 23716 30036 23722 30048
rect 23753 30039 23811 30045
rect 23753 30036 23765 30039
rect 23716 30008 23765 30036
rect 23716 29996 23722 30008
rect 23753 30005 23765 30008
rect 23799 30005 23811 30039
rect 23753 29999 23811 30005
rect 33321 30039 33379 30045
rect 33321 30005 33333 30039
rect 33367 30036 33379 30039
rect 33870 30036 33876 30048
rect 33367 30008 33876 30036
rect 33367 30005 33379 30008
rect 33321 29999 33379 30005
rect 33870 29996 33876 30008
rect 33928 29996 33934 30048
rect 1104 29946 39836 29968
rect 1104 29894 19606 29946
rect 19658 29894 19670 29946
rect 19722 29894 19734 29946
rect 19786 29894 19798 29946
rect 19850 29894 39836 29946
rect 1104 29872 39836 29894
rect 5534 29792 5540 29844
rect 5592 29832 5598 29844
rect 6546 29832 6552 29844
rect 5592 29804 6552 29832
rect 5592 29792 5598 29804
rect 6546 29792 6552 29804
rect 6604 29832 6610 29844
rect 6604 29804 7696 29832
rect 6604 29792 6610 29804
rect 4522 29724 4528 29776
rect 4580 29764 4586 29776
rect 7668 29764 7696 29804
rect 9306 29792 9312 29844
rect 9364 29832 9370 29844
rect 13630 29832 13636 29844
rect 9364 29804 13636 29832
rect 9364 29792 9370 29804
rect 13630 29792 13636 29804
rect 13688 29792 13694 29844
rect 13998 29792 14004 29844
rect 14056 29832 14062 29844
rect 16298 29832 16304 29844
rect 14056 29804 16304 29832
rect 14056 29792 14062 29804
rect 16298 29792 16304 29804
rect 16356 29792 16362 29844
rect 17129 29835 17187 29841
rect 17129 29801 17141 29835
rect 17175 29832 17187 29835
rect 25225 29835 25283 29841
rect 17175 29804 19196 29832
rect 17175 29801 17187 29804
rect 17129 29795 17187 29801
rect 9582 29764 9588 29776
rect 4580 29736 7604 29764
rect 7668 29736 9588 29764
rect 4580 29724 4586 29736
rect 4065 29699 4123 29705
rect 4065 29665 4077 29699
rect 4111 29665 4123 29699
rect 4614 29696 4620 29708
rect 4575 29668 4620 29696
rect 4065 29659 4123 29665
rect 1394 29628 1400 29640
rect 1355 29600 1400 29628
rect 1394 29588 1400 29600
rect 1452 29588 1458 29640
rect 1673 29631 1731 29637
rect 1673 29597 1685 29631
rect 1719 29628 1731 29631
rect 1854 29628 1860 29640
rect 1719 29600 1860 29628
rect 1719 29597 1731 29600
rect 1673 29591 1731 29597
rect 1854 29588 1860 29600
rect 1912 29588 1918 29640
rect 2961 29495 3019 29501
rect 2961 29461 2973 29495
rect 3007 29492 3019 29495
rect 3142 29492 3148 29504
rect 3007 29464 3148 29492
rect 3007 29461 3019 29464
rect 2961 29455 3019 29461
rect 3142 29452 3148 29464
rect 3200 29452 3206 29504
rect 3970 29452 3976 29504
rect 4028 29492 4034 29504
rect 4080 29492 4108 29659
rect 4614 29656 4620 29668
rect 4672 29656 4678 29708
rect 5442 29656 5448 29708
rect 5500 29696 5506 29708
rect 5997 29699 6055 29705
rect 5997 29696 6009 29699
rect 5500 29668 6009 29696
rect 5500 29656 5506 29668
rect 5997 29665 6009 29668
rect 6043 29665 6055 29699
rect 5997 29659 6055 29665
rect 6549 29699 6607 29705
rect 6549 29665 6561 29699
rect 6595 29665 6607 29699
rect 6549 29659 6607 29665
rect 4890 29628 4896 29640
rect 4851 29600 4896 29628
rect 4890 29588 4896 29600
rect 4948 29588 4954 29640
rect 5810 29628 5816 29640
rect 5771 29600 5816 29628
rect 5810 29588 5816 29600
rect 5868 29588 5874 29640
rect 4341 29563 4399 29569
rect 4341 29529 4353 29563
rect 4387 29560 4399 29563
rect 4798 29560 4804 29572
rect 4387 29532 4804 29560
rect 4387 29529 4399 29532
rect 4341 29523 4399 29529
rect 4798 29520 4804 29532
rect 4856 29520 4862 29572
rect 5626 29520 5632 29572
rect 5684 29560 5690 29572
rect 6457 29563 6515 29569
rect 6457 29560 6469 29563
rect 5684 29532 6469 29560
rect 5684 29520 5690 29532
rect 6457 29529 6469 29532
rect 6503 29529 6515 29563
rect 6564 29560 6592 29659
rect 7006 29656 7012 29708
rect 7064 29696 7070 29708
rect 7576 29705 7604 29736
rect 9582 29724 9588 29736
rect 9640 29724 9646 29776
rect 9766 29724 9772 29776
rect 9824 29764 9830 29776
rect 13906 29764 13912 29776
rect 9824 29736 9904 29764
rect 9824 29724 9830 29736
rect 7193 29699 7251 29705
rect 7193 29696 7205 29699
rect 7064 29668 7205 29696
rect 7064 29656 7070 29668
rect 7193 29665 7205 29668
rect 7239 29665 7251 29699
rect 7193 29659 7251 29665
rect 7561 29699 7619 29705
rect 7561 29665 7573 29699
rect 7607 29665 7619 29699
rect 7561 29659 7619 29665
rect 7745 29699 7803 29705
rect 7745 29665 7757 29699
rect 7791 29665 7803 29699
rect 7745 29659 7803 29665
rect 7374 29588 7380 29640
rect 7432 29628 7438 29640
rect 7760 29628 7788 29659
rect 8110 29656 8116 29708
rect 8168 29696 8174 29708
rect 8389 29699 8447 29705
rect 8389 29696 8401 29699
rect 8168 29668 8401 29696
rect 8168 29656 8174 29668
rect 8389 29665 8401 29668
rect 8435 29665 8447 29699
rect 9876 29696 9904 29736
rect 12636 29736 13912 29764
rect 12636 29705 12664 29736
rect 13906 29724 13912 29736
rect 13964 29724 13970 29776
rect 15470 29724 15476 29776
rect 15528 29764 15534 29776
rect 16758 29764 16764 29776
rect 15528 29736 16764 29764
rect 15528 29724 15534 29736
rect 10045 29699 10103 29705
rect 10045 29696 10057 29699
rect 9876 29668 10057 29696
rect 8389 29659 8447 29665
rect 10045 29665 10057 29668
rect 10091 29665 10103 29699
rect 10045 29659 10103 29665
rect 12621 29699 12679 29705
rect 12621 29665 12633 29699
rect 12667 29665 12679 29699
rect 12621 29659 12679 29665
rect 12713 29699 12771 29705
rect 12713 29665 12725 29699
rect 12759 29665 12771 29699
rect 13354 29696 13360 29708
rect 13267 29668 13360 29696
rect 12713 29659 12771 29665
rect 7432 29600 7788 29628
rect 9769 29631 9827 29637
rect 7432 29588 7438 29600
rect 9769 29597 9781 29631
rect 9815 29628 9827 29631
rect 11146 29628 11152 29640
rect 9815 29600 11152 29628
rect 9815 29597 9827 29600
rect 9769 29591 9827 29597
rect 11146 29588 11152 29600
rect 11204 29588 11210 29640
rect 12526 29628 12532 29640
rect 12487 29600 12532 29628
rect 12526 29588 12532 29600
rect 12584 29588 12590 29640
rect 9674 29560 9680 29572
rect 6564 29532 9680 29560
rect 6457 29523 6515 29529
rect 9674 29520 9680 29532
rect 9732 29520 9738 29572
rect 11333 29563 11391 29569
rect 11333 29529 11345 29563
rect 11379 29560 11391 29563
rect 12250 29560 12256 29572
rect 11379 29532 12256 29560
rect 11379 29529 11391 29532
rect 11333 29523 11391 29529
rect 12250 29520 12256 29532
rect 12308 29560 12314 29572
rect 12728 29560 12756 29659
rect 13354 29656 13360 29668
rect 13412 29656 13418 29708
rect 13817 29699 13875 29705
rect 13817 29665 13829 29699
rect 13863 29696 13875 29699
rect 14090 29696 14096 29708
rect 13863 29668 14096 29696
rect 13863 29665 13875 29668
rect 13817 29659 13875 29665
rect 14090 29656 14096 29668
rect 14148 29656 14154 29708
rect 14274 29696 14280 29708
rect 14235 29668 14280 29696
rect 14274 29656 14280 29668
rect 14332 29656 14338 29708
rect 15194 29656 15200 29708
rect 15252 29696 15258 29708
rect 15289 29699 15347 29705
rect 15289 29696 15301 29699
rect 15252 29668 15301 29696
rect 15252 29656 15258 29668
rect 15289 29665 15301 29668
rect 15335 29696 15347 29699
rect 15838 29696 15844 29708
rect 15335 29668 15844 29696
rect 15335 29665 15347 29668
rect 15289 29659 15347 29665
rect 15838 29656 15844 29668
rect 15896 29656 15902 29708
rect 15948 29705 15976 29736
rect 16758 29724 16764 29736
rect 16816 29724 16822 29776
rect 15933 29699 15991 29705
rect 15933 29665 15945 29699
rect 15979 29665 15991 29699
rect 16114 29696 16120 29708
rect 16075 29668 16120 29696
rect 15933 29659 15991 29665
rect 16114 29656 16120 29668
rect 16172 29656 16178 29708
rect 16298 29656 16304 29708
rect 16356 29696 16362 29708
rect 17037 29699 17095 29705
rect 17037 29696 17049 29699
rect 16356 29668 17049 29696
rect 16356 29656 16362 29668
rect 17037 29665 17049 29668
rect 17083 29665 17095 29699
rect 17037 29659 17095 29665
rect 17773 29699 17831 29705
rect 17773 29665 17785 29699
rect 17819 29696 17831 29699
rect 19058 29696 19064 29708
rect 17819 29668 19064 29696
rect 17819 29665 17831 29668
rect 17773 29659 17831 29665
rect 19058 29656 19064 29668
rect 19116 29656 19122 29708
rect 19168 29696 19196 29804
rect 25225 29801 25237 29835
rect 25271 29832 25283 29835
rect 25314 29832 25320 29844
rect 25271 29804 25320 29832
rect 25271 29801 25283 29804
rect 25225 29795 25283 29801
rect 25314 29792 25320 29804
rect 25372 29792 25378 29844
rect 25406 29792 25412 29844
rect 25464 29832 25470 29844
rect 31021 29835 31079 29841
rect 25464 29804 28488 29832
rect 25464 29792 25470 29804
rect 22002 29764 22008 29776
rect 21963 29736 22008 29764
rect 22002 29724 22008 29736
rect 22060 29724 22066 29776
rect 24578 29764 24584 29776
rect 24228 29736 24584 29764
rect 24228 29708 24256 29736
rect 24578 29724 24584 29736
rect 24636 29764 24642 29776
rect 24636 29736 25452 29764
rect 24636 29724 24642 29736
rect 19429 29699 19487 29705
rect 19429 29696 19441 29699
rect 19168 29668 19441 29696
rect 19429 29665 19441 29668
rect 19475 29665 19487 29699
rect 19429 29659 19487 29665
rect 19978 29656 19984 29708
rect 20036 29696 20042 29708
rect 20165 29699 20223 29705
rect 20165 29696 20177 29699
rect 20036 29668 20177 29696
rect 20036 29656 20042 29668
rect 20165 29665 20177 29668
rect 20211 29665 20223 29699
rect 21266 29696 21272 29708
rect 21227 29668 21272 29696
rect 20165 29659 20223 29665
rect 21266 29656 21272 29668
rect 21324 29656 21330 29708
rect 21726 29696 21732 29708
rect 21687 29668 21732 29696
rect 21726 29656 21732 29668
rect 21784 29656 21790 29708
rect 23293 29699 23351 29705
rect 23293 29665 23305 29699
rect 23339 29665 23351 29699
rect 23293 29659 23351 29665
rect 13372 29628 13400 29656
rect 16132 29628 16160 29656
rect 13372 29600 16160 29628
rect 18049 29631 18107 29637
rect 18049 29597 18061 29631
rect 18095 29628 18107 29631
rect 18785 29631 18843 29637
rect 18785 29628 18797 29631
rect 18095 29600 18797 29628
rect 18095 29597 18107 29600
rect 18049 29591 18107 29597
rect 18785 29597 18797 29600
rect 18831 29628 18843 29631
rect 19334 29628 19340 29640
rect 18831 29600 19340 29628
rect 18831 29597 18843 29600
rect 18785 29591 18843 29597
rect 19334 29588 19340 29600
rect 19392 29588 19398 29640
rect 21085 29631 21143 29637
rect 21085 29597 21097 29631
rect 21131 29628 21143 29631
rect 22646 29628 22652 29640
rect 21131 29600 22652 29628
rect 21131 29597 21143 29600
rect 21085 29591 21143 29597
rect 22646 29588 22652 29600
rect 22704 29588 22710 29640
rect 12308 29532 12756 29560
rect 12308 29520 12314 29532
rect 12894 29520 12900 29572
rect 12952 29560 12958 29572
rect 14461 29563 14519 29569
rect 14461 29560 14473 29563
rect 12952 29532 14473 29560
rect 12952 29520 12958 29532
rect 14461 29529 14473 29532
rect 14507 29560 14519 29563
rect 15194 29560 15200 29572
rect 14507 29532 15200 29560
rect 14507 29529 14519 29532
rect 14461 29523 14519 29529
rect 15194 29520 15200 29532
rect 15252 29520 15258 29572
rect 15286 29520 15292 29572
rect 15344 29560 15350 29572
rect 15381 29563 15439 29569
rect 15381 29560 15393 29563
rect 15344 29532 15393 29560
rect 15344 29520 15350 29532
rect 15381 29529 15393 29532
rect 15427 29529 15439 29563
rect 15381 29523 15439 29529
rect 17310 29520 17316 29572
rect 17368 29560 17374 29572
rect 19429 29563 19487 29569
rect 19429 29560 19441 29563
rect 17368 29532 19441 29560
rect 17368 29520 17374 29532
rect 19429 29529 19441 29532
rect 19475 29529 19487 29563
rect 23308 29560 23336 29659
rect 23382 29656 23388 29708
rect 23440 29696 23446 29708
rect 23569 29699 23627 29705
rect 23569 29696 23581 29699
rect 23440 29668 23581 29696
rect 23440 29656 23446 29668
rect 23569 29665 23581 29668
rect 23615 29665 23627 29699
rect 24026 29696 24032 29708
rect 23987 29668 24032 29696
rect 23569 29659 23627 29665
rect 24026 29656 24032 29668
rect 24084 29656 24090 29708
rect 24210 29696 24216 29708
rect 24171 29668 24216 29696
rect 24210 29656 24216 29668
rect 24268 29656 24274 29708
rect 25225 29699 25283 29705
rect 25225 29665 25237 29699
rect 25271 29696 25283 29699
rect 25314 29696 25320 29708
rect 25271 29668 25320 29696
rect 25271 29665 25283 29668
rect 25225 29659 25283 29665
rect 25314 29656 25320 29668
rect 25372 29656 25378 29708
rect 25424 29705 25452 29736
rect 27338 29724 27344 29776
rect 27396 29764 27402 29776
rect 27985 29767 28043 29773
rect 27985 29764 27997 29767
rect 27396 29736 27997 29764
rect 27396 29724 27402 29736
rect 27985 29733 27997 29736
rect 28031 29733 28043 29767
rect 27985 29727 28043 29733
rect 25409 29699 25467 29705
rect 25409 29665 25421 29699
rect 25455 29665 25467 29699
rect 27249 29699 27307 29705
rect 27249 29696 27261 29699
rect 25409 29659 25467 29665
rect 25516 29668 27261 29696
rect 23477 29631 23535 29637
rect 23477 29597 23489 29631
rect 23523 29628 23535 29631
rect 25516 29628 25544 29668
rect 27249 29665 27261 29668
rect 27295 29665 27307 29699
rect 27249 29659 27307 29665
rect 27801 29699 27859 29705
rect 27801 29665 27813 29699
rect 27847 29696 27859 29699
rect 28074 29696 28080 29708
rect 27847 29668 28080 29696
rect 27847 29665 27859 29668
rect 27801 29659 27859 29665
rect 28074 29656 28080 29668
rect 28132 29656 28138 29708
rect 28460 29705 28488 29804
rect 31021 29801 31033 29835
rect 31067 29832 31079 29835
rect 32950 29832 32956 29844
rect 31067 29804 32956 29832
rect 31067 29801 31079 29804
rect 31021 29795 31079 29801
rect 32950 29792 32956 29804
rect 33008 29792 33014 29844
rect 34790 29792 34796 29844
rect 34848 29832 34854 29844
rect 34977 29835 35035 29841
rect 34977 29832 34989 29835
rect 34848 29804 34989 29832
rect 34848 29792 34854 29804
rect 34977 29801 34989 29804
rect 35023 29801 35035 29835
rect 34977 29795 35035 29801
rect 35897 29835 35955 29841
rect 35897 29801 35909 29835
rect 35943 29832 35955 29835
rect 38470 29832 38476 29844
rect 35943 29804 38476 29832
rect 35943 29801 35955 29804
rect 35897 29795 35955 29801
rect 38470 29792 38476 29804
rect 38528 29792 38534 29844
rect 29270 29724 29276 29776
rect 29328 29764 29334 29776
rect 30558 29764 30564 29776
rect 29328 29736 30420 29764
rect 30519 29736 30564 29764
rect 29328 29724 29334 29736
rect 28445 29699 28503 29705
rect 28445 29665 28457 29699
rect 28491 29665 28503 29699
rect 28445 29659 28503 29665
rect 29362 29656 29368 29708
rect 29420 29696 29426 29708
rect 29457 29699 29515 29705
rect 29457 29696 29469 29699
rect 29420 29668 29469 29696
rect 29420 29656 29426 29668
rect 29457 29665 29469 29668
rect 29503 29665 29515 29699
rect 30006 29696 30012 29708
rect 29967 29668 30012 29696
rect 29457 29659 29515 29665
rect 30006 29656 30012 29668
rect 30064 29656 30070 29708
rect 30282 29696 30288 29708
rect 30243 29668 30288 29696
rect 30282 29656 30288 29668
rect 30340 29656 30346 29708
rect 30392 29696 30420 29736
rect 30558 29724 30564 29736
rect 30616 29724 30622 29776
rect 32214 29724 32220 29776
rect 32272 29764 32278 29776
rect 37458 29764 37464 29776
rect 32272 29736 32720 29764
rect 32272 29724 32278 29736
rect 31205 29699 31263 29705
rect 31205 29696 31217 29699
rect 30392 29668 31217 29696
rect 31205 29665 31217 29668
rect 31251 29665 31263 29699
rect 31205 29659 31263 29665
rect 31297 29699 31355 29705
rect 31297 29665 31309 29699
rect 31343 29665 31355 29699
rect 31297 29659 31355 29665
rect 32493 29699 32551 29705
rect 32493 29665 32505 29699
rect 32539 29696 32551 29699
rect 32582 29696 32588 29708
rect 32539 29668 32588 29696
rect 32539 29665 32551 29668
rect 32493 29659 32551 29665
rect 23523 29600 25544 29628
rect 23523 29597 23535 29600
rect 23477 29591 23535 29597
rect 26878 29588 26884 29640
rect 26936 29628 26942 29640
rect 27065 29631 27123 29637
rect 27065 29628 27077 29631
rect 26936 29600 27077 29628
rect 26936 29588 26942 29600
rect 27065 29597 27077 29600
rect 27111 29597 27123 29631
rect 27065 29591 27123 29597
rect 23658 29560 23664 29572
rect 23308 29532 23664 29560
rect 19429 29523 19487 29529
rect 23658 29520 23664 29532
rect 23716 29520 23722 29572
rect 27080 29560 27108 29591
rect 30374 29588 30380 29640
rect 30432 29628 30438 29640
rect 31312 29628 31340 29659
rect 32582 29656 32588 29668
rect 32640 29656 32646 29708
rect 32692 29705 32720 29736
rect 36740 29736 37464 29764
rect 32677 29699 32735 29705
rect 32677 29665 32689 29699
rect 32723 29665 32735 29699
rect 33870 29696 33876 29708
rect 33831 29668 33876 29696
rect 32677 29659 32735 29665
rect 33870 29656 33876 29668
rect 33928 29656 33934 29708
rect 36740 29705 36768 29736
rect 37458 29724 37464 29736
rect 37516 29724 37522 29776
rect 35805 29699 35863 29705
rect 35805 29665 35817 29699
rect 35851 29665 35863 29699
rect 35805 29659 35863 29665
rect 36725 29699 36783 29705
rect 36725 29665 36737 29699
rect 36771 29665 36783 29699
rect 36725 29659 36783 29665
rect 30432 29600 31340 29628
rect 33045 29631 33103 29637
rect 30432 29588 30438 29600
rect 33045 29597 33057 29631
rect 33091 29628 33103 29631
rect 33226 29628 33232 29640
rect 33091 29600 33232 29628
rect 33091 29597 33103 29600
rect 33045 29591 33103 29597
rect 33226 29588 33232 29600
rect 33284 29588 33290 29640
rect 33597 29631 33655 29637
rect 33597 29597 33609 29631
rect 33643 29628 33655 29631
rect 34514 29628 34520 29640
rect 33643 29600 34520 29628
rect 33643 29597 33655 29600
rect 33597 29591 33655 29597
rect 34514 29588 34520 29600
rect 34572 29588 34578 29640
rect 35820 29628 35848 29659
rect 36814 29656 36820 29708
rect 36872 29696 36878 29708
rect 37001 29699 37059 29705
rect 37001 29696 37013 29699
rect 36872 29668 37013 29696
rect 36872 29656 36878 29668
rect 37001 29665 37013 29668
rect 37047 29665 37059 29699
rect 37001 29659 37059 29665
rect 37921 29699 37979 29705
rect 37921 29665 37933 29699
rect 37967 29665 37979 29699
rect 38102 29696 38108 29708
rect 38063 29668 38108 29696
rect 37921 29659 37979 29665
rect 35820 29600 36584 29628
rect 27246 29560 27252 29572
rect 27080 29532 27252 29560
rect 27246 29520 27252 29532
rect 27304 29520 27310 29572
rect 31481 29563 31539 29569
rect 31481 29529 31493 29563
rect 31527 29560 31539 29563
rect 31570 29560 31576 29572
rect 31527 29532 31576 29560
rect 31527 29529 31539 29532
rect 31481 29523 31539 29529
rect 31570 29520 31576 29532
rect 31628 29520 31634 29572
rect 36556 29504 36584 29600
rect 37936 29560 37964 29659
rect 38102 29656 38108 29668
rect 38160 29656 38166 29708
rect 38289 29699 38347 29705
rect 38289 29665 38301 29699
rect 38335 29665 38347 29699
rect 38933 29699 38991 29705
rect 38933 29696 38945 29699
rect 38289 29659 38347 29665
rect 38764 29668 38945 29696
rect 38010 29588 38016 29640
rect 38068 29628 38074 29640
rect 38304 29628 38332 29659
rect 38068 29600 38332 29628
rect 38068 29588 38074 29600
rect 38764 29572 38792 29668
rect 38933 29665 38945 29668
rect 38979 29665 38991 29699
rect 38933 29659 38991 29665
rect 38746 29560 38752 29572
rect 37936 29532 38752 29560
rect 38746 29520 38752 29532
rect 38804 29520 38810 29572
rect 7742 29492 7748 29504
rect 4028 29464 7748 29492
rect 4028 29452 4034 29464
rect 7742 29452 7748 29464
rect 7800 29452 7806 29504
rect 8386 29452 8392 29504
rect 8444 29492 8450 29504
rect 8573 29495 8631 29501
rect 8573 29492 8585 29495
rect 8444 29464 8585 29492
rect 8444 29452 8450 29464
rect 8573 29461 8585 29464
rect 8619 29492 8631 29495
rect 10778 29492 10784 29504
rect 8619 29464 10784 29492
rect 8619 29461 8631 29464
rect 8573 29455 8631 29461
rect 10778 29452 10784 29464
rect 10836 29452 10842 29504
rect 10870 29452 10876 29504
rect 10928 29492 10934 29504
rect 13998 29492 14004 29504
rect 10928 29464 14004 29492
rect 10928 29452 10934 29464
rect 13998 29452 14004 29464
rect 14056 29452 14062 29504
rect 19150 29452 19156 29504
rect 19208 29492 19214 29504
rect 20257 29495 20315 29501
rect 20257 29492 20269 29495
rect 19208 29464 20269 29492
rect 19208 29452 19214 29464
rect 20257 29461 20269 29464
rect 20303 29461 20315 29495
rect 28626 29492 28632 29504
rect 28587 29464 28632 29492
rect 20257 29455 20315 29461
rect 28626 29452 28632 29464
rect 28684 29452 28690 29504
rect 36538 29492 36544 29504
rect 36499 29464 36544 29492
rect 36538 29452 36544 29464
rect 36596 29452 36602 29504
rect 39022 29492 39028 29504
rect 38983 29464 39028 29492
rect 39022 29452 39028 29464
rect 39080 29452 39086 29504
rect 1104 29402 39836 29424
rect 1104 29350 4246 29402
rect 4298 29350 4310 29402
rect 4362 29350 4374 29402
rect 4426 29350 4438 29402
rect 4490 29350 34966 29402
rect 35018 29350 35030 29402
rect 35082 29350 35094 29402
rect 35146 29350 35158 29402
rect 35210 29350 39836 29402
rect 1104 29328 39836 29350
rect 1854 29288 1860 29300
rect 1815 29260 1860 29288
rect 1854 29248 1860 29260
rect 1912 29248 1918 29300
rect 5074 29248 5080 29300
rect 5132 29288 5138 29300
rect 5721 29291 5779 29297
rect 5721 29288 5733 29291
rect 5132 29260 5733 29288
rect 5132 29248 5138 29260
rect 5721 29257 5733 29260
rect 5767 29257 5779 29291
rect 5721 29251 5779 29257
rect 6181 29291 6239 29297
rect 6181 29257 6193 29291
rect 6227 29288 6239 29291
rect 8478 29288 8484 29300
rect 6227 29260 8484 29288
rect 6227 29257 6239 29260
rect 6181 29251 6239 29257
rect 8478 29248 8484 29260
rect 8536 29248 8542 29300
rect 13814 29288 13820 29300
rect 8680 29260 13820 29288
rect 2958 29180 2964 29232
rect 3016 29220 3022 29232
rect 3145 29223 3203 29229
rect 3145 29220 3157 29223
rect 3016 29192 3157 29220
rect 3016 29180 3022 29192
rect 3145 29189 3157 29192
rect 3191 29189 3203 29223
rect 7006 29220 7012 29232
rect 3145 29183 3203 29189
rect 6012 29192 7012 29220
rect 4893 29155 4951 29161
rect 4893 29152 4905 29155
rect 1780 29124 4905 29152
rect 1780 29093 1808 29124
rect 4893 29121 4905 29124
rect 4939 29121 4951 29155
rect 4893 29115 4951 29121
rect 1765 29087 1823 29093
rect 1765 29053 1777 29087
rect 1811 29053 1823 29087
rect 2406 29084 2412 29096
rect 2367 29056 2412 29084
rect 1765 29047 1823 29053
rect 2406 29044 2412 29056
rect 2464 29044 2470 29096
rect 3050 29084 3056 29096
rect 3011 29056 3056 29084
rect 3050 29044 3056 29056
rect 3108 29044 3114 29096
rect 3234 29084 3240 29096
rect 3195 29056 3240 29084
rect 3234 29044 3240 29056
rect 3292 29044 3298 29096
rect 4154 29084 4160 29096
rect 4115 29056 4160 29084
rect 4154 29044 4160 29056
rect 4212 29044 4218 29096
rect 4525 29087 4583 29093
rect 4525 29053 4537 29087
rect 4571 29084 4583 29087
rect 4614 29084 4620 29096
rect 4571 29056 4620 29084
rect 4571 29053 4583 29056
rect 4525 29047 4583 29053
rect 4614 29044 4620 29056
rect 4672 29044 4678 29096
rect 4798 29084 4804 29096
rect 4759 29056 4804 29084
rect 4798 29044 4804 29056
rect 4856 29044 4862 29096
rect 6012 29093 6040 29192
rect 7006 29180 7012 29192
rect 7064 29180 7070 29232
rect 8386 29220 8392 29232
rect 7208 29192 8392 29220
rect 7208 29152 7236 29192
rect 8386 29180 8392 29192
rect 8444 29180 8450 29232
rect 8110 29152 8116 29164
rect 6840 29124 7236 29152
rect 7484 29124 8116 29152
rect 6840 29093 6868 29124
rect 5905 29087 5963 29093
rect 5905 29053 5917 29087
rect 5951 29053 5963 29087
rect 5905 29047 5963 29053
rect 5997 29087 6055 29093
rect 5997 29053 6009 29087
rect 6043 29053 6055 29087
rect 5997 29047 6055 29053
rect 6831 29087 6889 29093
rect 6831 29053 6843 29087
rect 6877 29053 6889 29087
rect 6831 29047 6889 29053
rect 4172 29016 4200 29044
rect 4890 29016 4896 29028
rect 4172 28988 4896 29016
rect 4890 28976 4896 28988
rect 4948 28976 4954 29028
rect 5920 29016 5948 29047
rect 7006 29044 7012 29096
rect 7064 29084 7070 29096
rect 7484 29084 7512 29124
rect 8110 29112 8116 29124
rect 8168 29112 8174 29164
rect 8294 29152 8300 29164
rect 8255 29124 8300 29152
rect 8294 29112 8300 29124
rect 8352 29112 8358 29164
rect 7064 29056 7512 29084
rect 7064 29044 7070 29056
rect 7558 29044 7564 29096
rect 7616 29084 7622 29096
rect 8680 29084 8708 29260
rect 13814 29248 13820 29260
rect 13872 29248 13878 29300
rect 13906 29248 13912 29300
rect 13964 29288 13970 29300
rect 14645 29291 14703 29297
rect 14645 29288 14657 29291
rect 13964 29260 14657 29288
rect 13964 29248 13970 29260
rect 14645 29257 14657 29260
rect 14691 29257 14703 29291
rect 16114 29288 16120 29300
rect 14645 29251 14703 29257
rect 14752 29260 16120 29288
rect 9766 29180 9772 29232
rect 9824 29220 9830 29232
rect 9861 29223 9919 29229
rect 9861 29220 9873 29223
rect 9824 29192 9873 29220
rect 9824 29180 9830 29192
rect 9861 29189 9873 29192
rect 9907 29189 9919 29223
rect 10870 29220 10876 29232
rect 9861 29183 9919 29189
rect 10152 29192 10876 29220
rect 10152 29152 10180 29192
rect 10870 29180 10876 29192
rect 10928 29180 10934 29232
rect 11330 29180 11336 29232
rect 11388 29180 11394 29232
rect 13630 29180 13636 29232
rect 13688 29220 13694 29232
rect 14752 29220 14780 29260
rect 16114 29248 16120 29260
rect 16172 29248 16178 29300
rect 16666 29248 16672 29300
rect 16724 29288 16730 29300
rect 16761 29291 16819 29297
rect 16761 29288 16773 29291
rect 16724 29260 16773 29288
rect 16724 29248 16730 29260
rect 16761 29257 16773 29260
rect 16807 29257 16819 29291
rect 16761 29251 16819 29257
rect 17405 29291 17463 29297
rect 17405 29257 17417 29291
rect 17451 29288 17463 29291
rect 18322 29288 18328 29300
rect 17451 29260 18328 29288
rect 17451 29257 17463 29260
rect 17405 29251 17463 29257
rect 13688 29192 14780 29220
rect 13688 29180 13694 29192
rect 11348 29152 11376 29180
rect 14090 29152 14096 29164
rect 8956 29124 10180 29152
rect 10520 29124 11376 29152
rect 11440 29124 14096 29152
rect 8846 29084 8852 29096
rect 7616 29056 8708 29084
rect 8807 29056 8852 29084
rect 7616 29044 7622 29056
rect 8846 29044 8852 29056
rect 8904 29044 8910 29096
rect 6914 29016 6920 29028
rect 5920 28988 6920 29016
rect 6914 28976 6920 28988
rect 6972 28976 6978 29028
rect 8864 29016 8892 29044
rect 7668 28988 8892 29016
rect 7009 28951 7067 28957
rect 7009 28917 7021 28951
rect 7055 28948 7067 28951
rect 7668 28948 7696 28988
rect 7055 28920 7696 28948
rect 7055 28917 7067 28920
rect 7009 28911 7067 28917
rect 7742 28908 7748 28960
rect 7800 28948 7806 28960
rect 8956 28948 8984 29124
rect 9125 29087 9183 29093
rect 9125 29053 9137 29087
rect 9171 29084 9183 29087
rect 9214 29084 9220 29096
rect 9171 29056 9220 29084
rect 9171 29053 9183 29056
rect 9125 29047 9183 29053
rect 9214 29044 9220 29056
rect 9272 29044 9278 29096
rect 9309 29087 9367 29093
rect 9309 29053 9321 29087
rect 9355 29053 9367 29087
rect 9950 29084 9956 29096
rect 9911 29056 9956 29084
rect 9309 29047 9367 29053
rect 9324 29016 9352 29047
rect 9950 29044 9956 29056
rect 10008 29044 10014 29096
rect 10520 29093 10548 29124
rect 10505 29087 10563 29093
rect 10505 29053 10517 29087
rect 10551 29053 10563 29087
rect 10505 29047 10563 29053
rect 10594 29044 10600 29096
rect 10652 29084 10658 29096
rect 10652 29056 10697 29084
rect 10652 29044 10658 29056
rect 10778 29044 10784 29096
rect 10836 29084 10842 29096
rect 11333 29087 11391 29093
rect 11333 29084 11345 29087
rect 10836 29056 11345 29084
rect 10836 29044 10842 29056
rect 11333 29053 11345 29056
rect 11379 29053 11391 29087
rect 11333 29047 11391 29053
rect 10410 29016 10416 29028
rect 9324 28988 10416 29016
rect 10410 28976 10416 28988
rect 10468 29016 10474 29028
rect 11440 29016 11468 29124
rect 14090 29112 14096 29124
rect 14148 29112 14154 29164
rect 14458 29112 14464 29164
rect 14516 29152 14522 29164
rect 15381 29155 15439 29161
rect 15381 29152 15393 29155
rect 14516 29124 15393 29152
rect 14516 29112 14522 29124
rect 15381 29121 15393 29124
rect 15427 29121 15439 29155
rect 15381 29115 15439 29121
rect 16117 29155 16175 29161
rect 16117 29121 16129 29155
rect 16163 29152 16175 29155
rect 16390 29152 16396 29164
rect 16163 29124 16396 29152
rect 16163 29121 16175 29124
rect 16117 29115 16175 29121
rect 16390 29112 16396 29124
rect 16448 29112 16454 29164
rect 16776 29152 16804 29251
rect 18322 29248 18328 29260
rect 18380 29248 18386 29300
rect 20990 29288 20996 29300
rect 19260 29260 20996 29288
rect 16776 29124 18092 29152
rect 12437 29087 12495 29093
rect 12437 29053 12449 29087
rect 12483 29053 12495 29087
rect 12710 29084 12716 29096
rect 12671 29056 12716 29084
rect 12437 29047 12495 29053
rect 10468 28988 11468 29016
rect 10468 28976 10474 28988
rect 7800 28920 8984 28948
rect 7800 28908 7806 28920
rect 9582 28908 9588 28960
rect 9640 28948 9646 28960
rect 11517 28951 11575 28957
rect 11517 28948 11529 28951
rect 9640 28920 11529 28948
rect 9640 28908 9646 28920
rect 11517 28917 11529 28920
rect 11563 28917 11575 28951
rect 11517 28911 11575 28917
rect 11698 28908 11704 28960
rect 11756 28948 11762 28960
rect 12452 28948 12480 29047
rect 12710 29044 12716 29056
rect 12768 29044 12774 29096
rect 14182 29044 14188 29096
rect 14240 29084 14246 29096
rect 14553 29087 14611 29093
rect 14553 29084 14565 29087
rect 14240 29056 14565 29084
rect 14240 29044 14246 29056
rect 14553 29053 14565 29056
rect 14599 29053 14611 29087
rect 14553 29047 14611 29053
rect 14642 29044 14648 29096
rect 14700 29084 14706 29096
rect 14700 29056 15792 29084
rect 14700 29044 14706 29056
rect 14090 29016 14096 29028
rect 14051 28988 14096 29016
rect 14090 28976 14096 28988
rect 14148 28976 14154 29028
rect 15654 29016 15660 29028
rect 15615 28988 15660 29016
rect 15654 28976 15660 28988
rect 15712 28976 15718 29028
rect 15764 29025 15792 29056
rect 16298 29044 16304 29096
rect 16356 29084 16362 29096
rect 16577 29087 16635 29093
rect 16577 29084 16589 29087
rect 16356 29056 16589 29084
rect 16356 29044 16362 29056
rect 16577 29053 16589 29056
rect 16623 29053 16635 29087
rect 17310 29084 17316 29096
rect 17271 29056 17316 29084
rect 16577 29047 16635 29053
rect 17310 29044 17316 29056
rect 17368 29044 17374 29096
rect 18064 29093 18092 29124
rect 18049 29087 18107 29093
rect 18049 29053 18061 29087
rect 18095 29053 18107 29087
rect 18049 29047 18107 29053
rect 18877 29087 18935 29093
rect 18877 29053 18889 29087
rect 18923 29084 18935 29087
rect 18966 29084 18972 29096
rect 18923 29056 18972 29084
rect 18923 29053 18935 29056
rect 18877 29047 18935 29053
rect 18966 29044 18972 29056
rect 19024 29044 19030 29096
rect 19058 29044 19064 29096
rect 19116 29084 19122 29096
rect 19116 29056 19161 29084
rect 19116 29044 19122 29056
rect 15749 29019 15807 29025
rect 15749 28985 15761 29019
rect 15795 28985 15807 29019
rect 15749 28979 15807 28985
rect 15838 28976 15844 29028
rect 15896 28976 15902 29028
rect 16114 28976 16120 29028
rect 16172 29016 16178 29028
rect 19260 29016 19288 29260
rect 20990 29248 20996 29260
rect 21048 29248 21054 29300
rect 21358 29248 21364 29300
rect 21416 29288 21422 29300
rect 29733 29291 29791 29297
rect 21416 29260 24256 29288
rect 21416 29248 21422 29260
rect 20162 29180 20168 29232
rect 20220 29220 20226 29232
rect 21729 29223 21787 29229
rect 20220 29192 21220 29220
rect 20220 29180 20226 29192
rect 20073 29155 20131 29161
rect 20073 29121 20085 29155
rect 20119 29152 20131 29155
rect 21082 29152 21088 29164
rect 20119 29124 21088 29152
rect 20119 29121 20131 29124
rect 20073 29115 20131 29121
rect 21082 29112 21088 29124
rect 21140 29112 21146 29164
rect 21192 29152 21220 29192
rect 21729 29189 21741 29223
rect 21775 29220 21787 29223
rect 22830 29220 22836 29232
rect 21775 29192 22836 29220
rect 21775 29189 21787 29192
rect 21729 29183 21787 29189
rect 22830 29180 22836 29192
rect 22888 29180 22894 29232
rect 22281 29155 22339 29161
rect 22281 29152 22293 29155
rect 21192 29124 22293 29152
rect 22281 29121 22293 29124
rect 22327 29121 22339 29155
rect 22281 29115 22339 29121
rect 24121 29155 24179 29161
rect 24121 29121 24133 29155
rect 24167 29121 24179 29155
rect 24121 29115 24179 29121
rect 20438 29084 20444 29096
rect 20399 29056 20444 29084
rect 20438 29044 20444 29056
rect 20496 29044 20502 29096
rect 20717 29087 20775 29093
rect 20717 29053 20729 29087
rect 20763 29053 20775 29087
rect 21542 29084 21548 29096
rect 21503 29056 21548 29084
rect 20717 29047 20775 29053
rect 16172 28988 19288 29016
rect 16172 28976 16178 28988
rect 19426 28976 19432 29028
rect 19484 29016 19490 29028
rect 20732 29016 20760 29047
rect 21542 29044 21548 29056
rect 21600 29044 21606 29096
rect 22094 29044 22100 29096
rect 22152 29084 22158 29096
rect 23658 29084 23664 29096
rect 22152 29056 22197 29084
rect 23619 29056 23664 29084
rect 22152 29044 22158 29056
rect 23658 29044 23664 29056
rect 23716 29044 23722 29096
rect 19484 28988 20760 29016
rect 20993 29019 21051 29025
rect 19484 28976 19490 28988
rect 20993 28985 21005 29019
rect 21039 29016 21051 29019
rect 23014 29016 23020 29028
rect 21039 28988 23020 29016
rect 21039 28985 21051 28988
rect 20993 28979 21051 28985
rect 23014 28976 23020 28988
rect 23072 28976 23078 29028
rect 24136 29016 24164 29115
rect 24228 29093 24256 29260
rect 29733 29257 29745 29291
rect 29779 29288 29791 29291
rect 30742 29288 30748 29300
rect 29779 29260 30748 29288
rect 29779 29257 29791 29260
rect 29733 29251 29791 29257
rect 30742 29248 30748 29260
rect 30800 29248 30806 29300
rect 32508 29260 34652 29288
rect 25222 29180 25228 29232
rect 25280 29220 25286 29232
rect 26421 29223 26479 29229
rect 26421 29220 26433 29223
rect 25280 29192 26433 29220
rect 25280 29180 25286 29192
rect 26421 29189 26433 29192
rect 26467 29189 26479 29223
rect 26421 29183 26479 29189
rect 24578 29112 24584 29164
rect 24636 29152 24642 29164
rect 28074 29152 28080 29164
rect 24636 29124 26004 29152
rect 28035 29124 28080 29152
rect 24636 29112 24642 29124
rect 24213 29087 24271 29093
rect 24213 29053 24225 29087
rect 24259 29053 24271 29087
rect 24213 29047 24271 29053
rect 24394 29044 24400 29096
rect 24452 29084 24458 29096
rect 24489 29087 24547 29093
rect 24489 29084 24501 29087
rect 24452 29056 24501 29084
rect 24452 29044 24458 29056
rect 24489 29053 24501 29056
rect 24535 29053 24547 29087
rect 24489 29047 24547 29053
rect 24762 29044 24768 29096
rect 24820 29084 24826 29096
rect 24857 29087 24915 29093
rect 24857 29084 24869 29087
rect 24820 29056 24869 29084
rect 24820 29044 24826 29056
rect 24857 29053 24869 29056
rect 24903 29053 24915 29087
rect 25590 29084 25596 29096
rect 25551 29056 25596 29084
rect 24857 29047 24915 29053
rect 25590 29044 25596 29056
rect 25648 29044 25654 29096
rect 25976 29093 26004 29124
rect 28074 29112 28080 29124
rect 28132 29112 28138 29164
rect 30285 29155 30343 29161
rect 30285 29121 30297 29155
rect 30331 29152 30343 29155
rect 31570 29152 31576 29164
rect 30331 29124 31576 29152
rect 30331 29121 30343 29124
rect 30285 29115 30343 29121
rect 31570 29112 31576 29124
rect 31628 29112 31634 29164
rect 25961 29087 26019 29093
rect 25961 29053 25973 29087
rect 26007 29053 26019 29087
rect 26418 29084 26424 29096
rect 26379 29056 26424 29084
rect 25961 29047 26019 29053
rect 26418 29044 26424 29056
rect 26476 29044 26482 29096
rect 27246 29084 27252 29096
rect 27207 29056 27252 29084
rect 27246 29044 27252 29056
rect 27304 29044 27310 29096
rect 27525 29087 27583 29093
rect 27525 29053 27537 29087
rect 27571 29053 27583 29087
rect 27525 29047 27583 29053
rect 27985 29087 28043 29093
rect 27985 29053 27997 29087
rect 28031 29053 28043 29087
rect 28902 29084 28908 29096
rect 28863 29056 28908 29084
rect 27985 29047 28043 29053
rect 27540 29016 27568 29047
rect 24136 28988 27568 29016
rect 28000 29016 28028 29047
rect 28902 29044 28908 29056
rect 28960 29044 28966 29096
rect 29546 29084 29552 29096
rect 29507 29056 29552 29084
rect 29546 29044 29552 29056
rect 29604 29044 29610 29096
rect 30561 29087 30619 29093
rect 30561 29053 30573 29087
rect 30607 29084 30619 29087
rect 31294 29084 31300 29096
rect 30607 29056 31300 29084
rect 30607 29053 30619 29056
rect 30561 29047 30619 29053
rect 31294 29044 31300 29056
rect 31352 29044 31358 29096
rect 31941 29087 31999 29093
rect 31941 29053 31953 29087
rect 31987 29084 31999 29087
rect 32306 29084 32312 29096
rect 31987 29056 32312 29084
rect 31987 29053 31999 29056
rect 31941 29047 31999 29053
rect 32306 29044 32312 29056
rect 32364 29084 32370 29096
rect 32401 29087 32459 29093
rect 32401 29084 32413 29087
rect 32364 29056 32413 29084
rect 32364 29044 32370 29056
rect 32401 29053 32413 29056
rect 32447 29053 32459 29087
rect 32508 29084 32536 29260
rect 33134 29180 33140 29232
rect 33192 29220 33198 29232
rect 33229 29223 33287 29229
rect 33229 29220 33241 29223
rect 33192 29192 33241 29220
rect 33192 29180 33198 29192
rect 33229 29189 33241 29192
rect 33275 29189 33287 29223
rect 33229 29183 33287 29189
rect 32582 29112 32588 29164
rect 32640 29152 32646 29164
rect 34624 29152 34652 29260
rect 34698 29180 34704 29232
rect 34756 29220 34762 29232
rect 35713 29223 35771 29229
rect 35713 29220 35725 29223
rect 34756 29192 35725 29220
rect 34756 29180 34762 29192
rect 35713 29189 35725 29192
rect 35759 29189 35771 29223
rect 35713 29183 35771 29189
rect 36633 29223 36691 29229
rect 36633 29189 36645 29223
rect 36679 29220 36691 29223
rect 37090 29220 37096 29232
rect 36679 29192 37096 29220
rect 36679 29189 36691 29192
rect 36633 29183 36691 29189
rect 36648 29152 36676 29183
rect 37090 29180 37096 29192
rect 37148 29220 37154 29232
rect 37148 29192 38148 29220
rect 37148 29180 37154 29192
rect 38010 29152 38016 29164
rect 32640 29124 34008 29152
rect 34624 29124 36676 29152
rect 37971 29124 38016 29152
rect 32640 29112 32646 29124
rect 32769 29087 32827 29093
rect 32769 29084 32781 29087
rect 32508 29056 32781 29084
rect 32401 29047 32459 29053
rect 32769 29053 32781 29056
rect 32815 29053 32827 29087
rect 33226 29084 33232 29096
rect 33187 29056 33232 29084
rect 32769 29047 32827 29053
rect 33226 29044 33232 29056
rect 33284 29044 33290 29096
rect 33980 29093 34008 29124
rect 33965 29087 34023 29093
rect 33965 29053 33977 29087
rect 34011 29084 34023 29087
rect 34011 29056 34284 29084
rect 34011 29053 34023 29056
rect 33965 29047 34023 29053
rect 29270 29016 29276 29028
rect 28000 28988 29276 29016
rect 29270 28976 29276 28988
rect 29328 28976 29334 29028
rect 34256 29016 34284 29056
rect 34790 29044 34796 29096
rect 34848 29084 34854 29096
rect 35268 29093 35296 29124
rect 38010 29112 38016 29124
rect 38068 29112 38074 29164
rect 34885 29087 34943 29093
rect 34885 29084 34897 29087
rect 34848 29056 34897 29084
rect 34848 29044 34854 29056
rect 34885 29053 34897 29056
rect 34931 29053 34943 29087
rect 34885 29047 34943 29053
rect 35253 29087 35311 29093
rect 35253 29053 35265 29087
rect 35299 29053 35311 29087
rect 35710 29084 35716 29096
rect 35671 29056 35716 29084
rect 35253 29047 35311 29053
rect 35710 29044 35716 29056
rect 35768 29044 35774 29096
rect 36449 29087 36507 29093
rect 36449 29053 36461 29087
rect 36495 29084 36507 29087
rect 36814 29084 36820 29096
rect 36495 29056 36820 29084
rect 36495 29053 36507 29056
rect 36449 29047 36507 29053
rect 36814 29044 36820 29056
rect 36872 29044 36878 29096
rect 37458 29084 37464 29096
rect 37419 29056 37464 29084
rect 37458 29044 37464 29056
rect 37516 29044 37522 29096
rect 37918 29084 37924 29096
rect 37879 29056 37924 29084
rect 37918 29044 37924 29056
rect 37976 29044 37982 29096
rect 38120 29093 38148 29192
rect 38105 29087 38163 29093
rect 38105 29053 38117 29087
rect 38151 29053 38163 29087
rect 38654 29084 38660 29096
rect 38615 29056 38660 29084
rect 38105 29047 38163 29053
rect 38654 29044 38660 29056
rect 38712 29044 38718 29096
rect 35894 29016 35900 29028
rect 34256 28988 35900 29016
rect 35894 28976 35900 28988
rect 35952 28976 35958 29028
rect 15286 28948 15292 28960
rect 11756 28920 15292 28948
rect 11756 28908 11762 28920
rect 15286 28908 15292 28920
rect 15344 28908 15350 28960
rect 15565 28951 15623 28957
rect 15565 28917 15577 28951
rect 15611 28948 15623 28951
rect 15856 28948 15884 28976
rect 15611 28920 15884 28948
rect 18325 28951 18383 28957
rect 15611 28917 15623 28920
rect 15565 28911 15623 28917
rect 18325 28917 18337 28951
rect 18371 28948 18383 28951
rect 18506 28948 18512 28960
rect 18371 28920 18512 28948
rect 18371 28917 18383 28920
rect 18325 28911 18383 28917
rect 18506 28908 18512 28920
rect 18564 28908 18570 28960
rect 18782 28908 18788 28960
rect 18840 28948 18846 28960
rect 18874 28948 18880 28960
rect 18840 28920 18880 28948
rect 18840 28908 18846 28920
rect 18874 28908 18880 28920
rect 18932 28908 18938 28960
rect 20162 28908 20168 28960
rect 20220 28948 20226 28960
rect 20622 28948 20628 28960
rect 20220 28920 20628 28948
rect 20220 28908 20226 28920
rect 20622 28908 20628 28920
rect 20680 28908 20686 28960
rect 27706 28908 27712 28960
rect 27764 28948 27770 28960
rect 28721 28951 28779 28957
rect 28721 28948 28733 28951
rect 27764 28920 28733 28948
rect 27764 28908 27770 28920
rect 28721 28917 28733 28920
rect 28767 28917 28779 28951
rect 28721 28911 28779 28917
rect 33594 28908 33600 28960
rect 33652 28948 33658 28960
rect 34149 28951 34207 28957
rect 34149 28948 34161 28951
rect 33652 28920 34161 28948
rect 33652 28908 33658 28920
rect 34149 28917 34161 28920
rect 34195 28917 34207 28951
rect 34149 28911 34207 28917
rect 36446 28908 36452 28960
rect 36504 28948 36510 28960
rect 36722 28948 36728 28960
rect 36504 28920 36728 28948
rect 36504 28908 36510 28920
rect 36722 28908 36728 28920
rect 36780 28908 36786 28960
rect 1104 28858 39836 28880
rect 1104 28806 19606 28858
rect 19658 28806 19670 28858
rect 19722 28806 19734 28858
rect 19786 28806 19798 28858
rect 19850 28806 39836 28858
rect 1104 28784 39836 28806
rect 3329 28747 3387 28753
rect 3329 28713 3341 28747
rect 3375 28744 3387 28747
rect 4154 28744 4160 28756
rect 3375 28716 4160 28744
rect 3375 28713 3387 28716
rect 3329 28707 3387 28713
rect 4154 28704 4160 28716
rect 4212 28704 4218 28756
rect 6914 28704 6920 28756
rect 6972 28744 6978 28756
rect 7653 28747 7711 28753
rect 7653 28744 7665 28747
rect 6972 28716 7665 28744
rect 6972 28704 6978 28716
rect 7653 28713 7665 28716
rect 7699 28744 7711 28747
rect 13449 28747 13507 28753
rect 7699 28716 11560 28744
rect 7699 28713 7711 28716
rect 7653 28707 7711 28713
rect 2133 28679 2191 28685
rect 2133 28645 2145 28679
rect 2179 28676 2191 28679
rect 4249 28679 4307 28685
rect 4249 28676 4261 28679
rect 2179 28648 4261 28676
rect 2179 28645 2191 28648
rect 2133 28639 2191 28645
rect 4249 28645 4261 28648
rect 4295 28676 4307 28679
rect 5534 28676 5540 28688
rect 4295 28648 5540 28676
rect 4295 28645 4307 28648
rect 4249 28639 4307 28645
rect 5534 28636 5540 28648
rect 5592 28636 5598 28688
rect 7101 28679 7159 28685
rect 7101 28645 7113 28679
rect 7147 28676 7159 28679
rect 7374 28676 7380 28688
rect 7147 28648 7380 28676
rect 7147 28645 7159 28648
rect 7101 28639 7159 28645
rect 7374 28636 7380 28648
rect 7432 28636 7438 28688
rect 9122 28676 9128 28688
rect 7852 28648 9128 28676
rect 2225 28611 2283 28617
rect 2225 28577 2237 28611
rect 2271 28608 2283 28611
rect 2314 28608 2320 28620
rect 2271 28580 2320 28608
rect 2271 28577 2283 28580
rect 2225 28571 2283 28577
rect 2314 28568 2320 28580
rect 2372 28568 2378 28620
rect 3142 28608 3148 28620
rect 3103 28580 3148 28608
rect 3142 28568 3148 28580
rect 3200 28568 3206 28620
rect 4157 28611 4215 28617
rect 4157 28577 4169 28611
rect 4203 28577 4215 28611
rect 4157 28571 4215 28577
rect 4341 28611 4399 28617
rect 4341 28577 4353 28611
rect 4387 28608 4399 28611
rect 5350 28608 5356 28620
rect 4387 28580 5356 28608
rect 4387 28577 4399 28580
rect 4341 28571 4399 28577
rect 4172 28540 4200 28571
rect 5350 28568 5356 28580
rect 5408 28568 5414 28620
rect 7852 28617 7880 28648
rect 9122 28636 9128 28648
rect 9180 28636 9186 28688
rect 11330 28676 11336 28688
rect 9784 28648 11336 28676
rect 9784 28617 9812 28648
rect 11330 28636 11336 28648
rect 11388 28636 11394 28688
rect 7837 28611 7895 28617
rect 7837 28577 7849 28611
rect 7883 28577 7895 28611
rect 7837 28571 7895 28577
rect 8573 28611 8631 28617
rect 8573 28577 8585 28611
rect 8619 28577 8631 28611
rect 8573 28571 8631 28577
rect 8941 28611 8999 28617
rect 8941 28577 8953 28611
rect 8987 28608 8999 28611
rect 9769 28611 9827 28617
rect 9769 28608 9781 28611
rect 8987 28580 9781 28608
rect 8987 28577 8999 28580
rect 8941 28571 8999 28577
rect 9769 28577 9781 28580
rect 9815 28577 9827 28611
rect 10134 28608 10140 28620
rect 10047 28580 10140 28608
rect 9769 28571 9827 28577
rect 4706 28540 4712 28552
rect 4172 28512 4712 28540
rect 4706 28500 4712 28512
rect 4764 28500 4770 28552
rect 5074 28500 5080 28552
rect 5132 28540 5138 28552
rect 5445 28543 5503 28549
rect 5445 28540 5457 28543
rect 5132 28512 5457 28540
rect 5132 28500 5138 28512
rect 5445 28509 5457 28512
rect 5491 28509 5503 28543
rect 5718 28540 5724 28552
rect 5679 28512 5724 28540
rect 5445 28503 5503 28509
rect 5718 28500 5724 28512
rect 5776 28500 5782 28552
rect 8202 28540 8208 28552
rect 8163 28512 8208 28540
rect 8202 28500 8208 28512
rect 8260 28500 8266 28552
rect 8588 28472 8616 28571
rect 10134 28568 10140 28580
rect 10192 28608 10198 28620
rect 10594 28608 10600 28620
rect 10192 28580 10600 28608
rect 10192 28568 10198 28580
rect 10594 28568 10600 28580
rect 10652 28568 10658 28620
rect 10781 28611 10839 28617
rect 10781 28577 10793 28611
rect 10827 28608 10839 28611
rect 10870 28608 10876 28620
rect 10827 28580 10876 28608
rect 10827 28577 10839 28580
rect 10781 28571 10839 28577
rect 10870 28568 10876 28580
rect 10928 28568 10934 28620
rect 11532 28617 11560 28716
rect 13449 28713 13461 28747
rect 13495 28713 13507 28747
rect 13449 28707 13507 28713
rect 13464 28676 13492 28707
rect 15562 28704 15568 28756
rect 15620 28744 15626 28756
rect 23477 28747 23535 28753
rect 15620 28716 21680 28744
rect 15620 28704 15626 28716
rect 11992 28648 12664 28676
rect 11992 28617 12020 28648
rect 11517 28611 11575 28617
rect 11517 28577 11529 28611
rect 11563 28577 11575 28611
rect 11517 28571 11575 28577
rect 11977 28611 12035 28617
rect 11977 28577 11989 28611
rect 12023 28577 12035 28611
rect 11977 28571 12035 28577
rect 12345 28611 12403 28617
rect 12345 28577 12357 28611
rect 12391 28577 12403 28611
rect 12345 28571 12403 28577
rect 9122 28540 9128 28552
rect 9083 28512 9128 28540
rect 9122 28500 9128 28512
rect 9180 28500 9186 28552
rect 10152 28472 10180 28568
rect 12360 28540 12388 28571
rect 12636 28540 12664 28648
rect 12728 28648 13492 28676
rect 12728 28617 12756 28648
rect 20070 28636 20076 28688
rect 20128 28676 20134 28688
rect 20346 28676 20352 28688
rect 20128 28648 20352 28676
rect 20128 28636 20134 28648
rect 20346 28636 20352 28648
rect 20404 28636 20410 28688
rect 12713 28611 12771 28617
rect 12713 28577 12725 28611
rect 12759 28577 12771 28611
rect 12713 28571 12771 28577
rect 13541 28611 13599 28617
rect 13541 28577 13553 28611
rect 13587 28608 13599 28611
rect 13630 28608 13636 28620
rect 13587 28580 13636 28608
rect 13587 28577 13599 28580
rect 13541 28571 13599 28577
rect 13630 28568 13636 28580
rect 13688 28568 13694 28620
rect 13909 28611 13967 28617
rect 13909 28577 13921 28611
rect 13955 28577 13967 28611
rect 13909 28571 13967 28577
rect 13924 28540 13952 28571
rect 14090 28568 14096 28620
rect 14148 28608 14154 28620
rect 14185 28611 14243 28617
rect 14185 28608 14197 28611
rect 14148 28580 14197 28608
rect 14148 28568 14154 28580
rect 14185 28577 14197 28580
rect 14231 28577 14243 28611
rect 15286 28608 15292 28620
rect 15199 28580 15292 28608
rect 14185 28571 14243 28577
rect 15286 28568 15292 28580
rect 15344 28608 15350 28620
rect 17589 28611 17647 28617
rect 15344 28580 15792 28608
rect 15344 28568 15350 28580
rect 15764 28552 15792 28580
rect 17589 28577 17601 28611
rect 17635 28608 17647 28611
rect 18046 28608 18052 28620
rect 17635 28580 18052 28608
rect 17635 28577 17647 28580
rect 17589 28571 17647 28577
rect 18046 28568 18052 28580
rect 18104 28568 18110 28620
rect 18506 28608 18512 28620
rect 18467 28580 18512 28608
rect 18506 28568 18512 28580
rect 18564 28568 18570 28620
rect 20990 28568 20996 28620
rect 21048 28608 21054 28620
rect 21361 28611 21419 28617
rect 21361 28608 21373 28611
rect 21048 28580 21373 28608
rect 21048 28568 21054 28580
rect 21361 28577 21373 28580
rect 21407 28608 21419 28611
rect 21542 28608 21548 28620
rect 21407 28580 21548 28608
rect 21407 28577 21419 28580
rect 21361 28571 21419 28577
rect 21542 28568 21548 28580
rect 21600 28568 21606 28620
rect 21652 28608 21680 28716
rect 23477 28713 23489 28747
rect 23523 28744 23535 28747
rect 24210 28744 24216 28756
rect 23523 28716 24216 28744
rect 23523 28713 23535 28716
rect 23477 28707 23535 28713
rect 24210 28704 24216 28716
rect 24268 28744 24274 28756
rect 24762 28744 24768 28756
rect 24268 28716 24768 28744
rect 24268 28704 24274 28716
rect 24762 28704 24768 28716
rect 24820 28704 24826 28756
rect 25869 28747 25927 28753
rect 25869 28713 25881 28747
rect 25915 28744 25927 28747
rect 27246 28744 27252 28756
rect 25915 28716 27252 28744
rect 25915 28713 25927 28716
rect 25869 28707 25927 28713
rect 27246 28704 27252 28716
rect 27304 28704 27310 28756
rect 30282 28704 30288 28756
rect 30340 28744 30346 28756
rect 35618 28744 35624 28756
rect 30340 28716 30788 28744
rect 30340 28704 30346 28716
rect 21913 28611 21971 28617
rect 21913 28608 21925 28611
rect 21652 28580 21925 28608
rect 21913 28577 21925 28580
rect 21959 28608 21971 28611
rect 22094 28608 22100 28620
rect 21959 28580 22100 28608
rect 21959 28577 21971 28580
rect 21913 28571 21971 28577
rect 22094 28568 22100 28580
rect 22152 28568 22158 28620
rect 23290 28608 23296 28620
rect 23251 28580 23296 28608
rect 23290 28568 23296 28580
rect 23348 28568 23354 28620
rect 23842 28568 23848 28620
rect 23900 28608 23906 28620
rect 24029 28611 24087 28617
rect 24029 28608 24041 28611
rect 23900 28580 24041 28608
rect 23900 28568 23906 28580
rect 24029 28577 24041 28580
rect 24075 28577 24087 28611
rect 24394 28608 24400 28620
rect 24355 28580 24400 28608
rect 24029 28571 24087 28577
rect 24394 28568 24400 28580
rect 24452 28568 24458 28620
rect 24762 28608 24768 28620
rect 24723 28580 24768 28608
rect 24762 28568 24768 28580
rect 24820 28568 24826 28620
rect 25406 28568 25412 28620
rect 25464 28608 25470 28620
rect 25685 28611 25743 28617
rect 25685 28608 25697 28611
rect 25464 28580 25697 28608
rect 25464 28568 25470 28580
rect 25685 28577 25697 28580
rect 25731 28577 25743 28611
rect 25685 28571 25743 28577
rect 26789 28611 26847 28617
rect 26789 28577 26801 28611
rect 26835 28577 26847 28611
rect 27246 28608 27252 28620
rect 27207 28580 27252 28608
rect 26789 28571 26847 28577
rect 13998 28540 14004 28552
rect 12360 28512 12572 28540
rect 12636 28512 14004 28540
rect 8588 28444 10180 28472
rect 10873 28475 10931 28481
rect 10873 28441 10885 28475
rect 10919 28472 10931 28475
rect 11238 28472 11244 28484
rect 10919 28444 11244 28472
rect 10919 28441 10931 28444
rect 10873 28435 10931 28441
rect 11238 28432 11244 28444
rect 11296 28472 11302 28484
rect 11606 28472 11612 28484
rect 11296 28444 11612 28472
rect 11296 28432 11302 28444
rect 11606 28432 11612 28444
rect 11664 28432 11670 28484
rect 12544 28472 12572 28512
rect 13998 28500 14004 28512
rect 14056 28500 14062 28552
rect 15470 28500 15476 28552
rect 15528 28540 15534 28552
rect 15565 28543 15623 28549
rect 15565 28540 15577 28543
rect 15528 28512 15577 28540
rect 15528 28500 15534 28512
rect 15565 28509 15577 28512
rect 15611 28509 15623 28543
rect 15565 28503 15623 28509
rect 15746 28500 15752 28552
rect 15804 28500 15810 28552
rect 17954 28500 17960 28552
rect 18012 28540 18018 28552
rect 18230 28540 18236 28552
rect 18012 28512 18236 28540
rect 18012 28500 18018 28512
rect 18230 28500 18236 28512
rect 18288 28500 18294 28552
rect 19242 28500 19248 28552
rect 19300 28540 19306 28552
rect 22189 28543 22247 28549
rect 22189 28540 22201 28543
rect 19300 28512 22201 28540
rect 19300 28500 19306 28512
rect 22189 28509 22201 28512
rect 22235 28509 22247 28543
rect 24670 28540 24676 28552
rect 24631 28512 24676 28540
rect 22189 28503 22247 28509
rect 24670 28500 24676 28512
rect 24728 28500 24734 28552
rect 12618 28472 12624 28484
rect 12544 28444 12624 28472
rect 12618 28432 12624 28444
rect 12676 28432 12682 28484
rect 12713 28475 12771 28481
rect 12713 28441 12725 28475
rect 12759 28441 12771 28475
rect 12713 28435 12771 28441
rect 21637 28475 21695 28481
rect 21637 28441 21649 28475
rect 21683 28472 21695 28475
rect 22278 28472 22284 28484
rect 21683 28444 22284 28472
rect 21683 28441 21695 28444
rect 21637 28435 21695 28441
rect 1946 28404 1952 28416
rect 1907 28376 1952 28404
rect 1946 28364 1952 28376
rect 2004 28364 2010 28416
rect 2406 28404 2412 28416
rect 2367 28376 2412 28404
rect 2406 28364 2412 28376
rect 2464 28364 2470 28416
rect 4525 28407 4583 28413
rect 4525 28373 4537 28407
rect 4571 28404 4583 28407
rect 4614 28404 4620 28416
rect 4571 28376 4620 28404
rect 4571 28373 4583 28376
rect 4525 28367 4583 28373
rect 4614 28364 4620 28376
rect 4672 28364 4678 28416
rect 11146 28364 11152 28416
rect 11204 28404 11210 28416
rect 11333 28407 11391 28413
rect 11333 28404 11345 28407
rect 11204 28376 11345 28404
rect 11204 28364 11210 28376
rect 11333 28373 11345 28376
rect 11379 28404 11391 28407
rect 11698 28404 11704 28416
rect 11379 28376 11704 28404
rect 11379 28373 11391 28376
rect 11333 28367 11391 28373
rect 11698 28364 11704 28376
rect 11756 28364 11762 28416
rect 12728 28404 12756 28435
rect 22278 28432 22284 28444
rect 22336 28432 22342 28484
rect 23750 28432 23756 28484
rect 23808 28472 23814 28484
rect 25424 28472 25452 28568
rect 26804 28540 26832 28571
rect 27246 28568 27252 28580
rect 27304 28568 27310 28620
rect 28074 28608 28080 28620
rect 28035 28580 28080 28608
rect 28074 28568 28080 28580
rect 28132 28568 28138 28620
rect 28718 28568 28724 28620
rect 28776 28608 28782 28620
rect 29917 28611 29975 28617
rect 29917 28608 29929 28611
rect 28776 28580 29929 28608
rect 28776 28568 28782 28580
rect 29917 28577 29929 28580
rect 29963 28577 29975 28611
rect 30374 28608 30380 28620
rect 30335 28580 30380 28608
rect 29917 28571 29975 28577
rect 30374 28568 30380 28580
rect 30432 28568 30438 28620
rect 30760 28617 30788 28716
rect 32876 28716 35624 28744
rect 31021 28679 31079 28685
rect 31021 28645 31033 28679
rect 31067 28676 31079 28679
rect 32490 28676 32496 28688
rect 31067 28648 32496 28676
rect 31067 28645 31079 28648
rect 31021 28639 31079 28645
rect 32490 28636 32496 28648
rect 32548 28636 32554 28688
rect 30745 28611 30803 28617
rect 30745 28577 30757 28611
rect 30791 28577 30803 28611
rect 30745 28571 30803 28577
rect 32309 28611 32367 28617
rect 32309 28577 32321 28611
rect 32355 28608 32367 28611
rect 32876 28608 32904 28716
rect 35618 28704 35624 28716
rect 35676 28704 35682 28756
rect 35250 28676 35256 28688
rect 35211 28648 35256 28676
rect 35250 28636 35256 28648
rect 35308 28636 35314 28688
rect 36630 28636 36636 28688
rect 36688 28676 36694 28688
rect 36817 28679 36875 28685
rect 36817 28676 36829 28679
rect 36688 28648 36829 28676
rect 36688 28636 36694 28648
rect 36817 28645 36829 28648
rect 36863 28645 36875 28679
rect 36817 28639 36875 28645
rect 32355 28580 32904 28608
rect 32953 28611 33011 28617
rect 32355 28577 32367 28580
rect 32309 28571 32367 28577
rect 32953 28577 32965 28611
rect 32999 28608 33011 28611
rect 35710 28608 35716 28620
rect 32999 28580 35572 28608
rect 35671 28580 35716 28608
rect 32999 28577 33011 28580
rect 32953 28571 33011 28577
rect 27614 28540 27620 28552
rect 26804 28512 27620 28540
rect 27614 28500 27620 28512
rect 27672 28500 27678 28552
rect 27706 28500 27712 28552
rect 27764 28540 27770 28552
rect 27801 28543 27859 28549
rect 27801 28540 27813 28543
rect 27764 28512 27813 28540
rect 27764 28500 27770 28512
rect 27801 28509 27813 28512
rect 27847 28509 27859 28543
rect 27801 28503 27859 28509
rect 32766 28500 32772 28552
rect 32824 28540 32830 28552
rect 33597 28543 33655 28549
rect 33597 28540 33609 28543
rect 32824 28512 33609 28540
rect 32824 28500 32830 28512
rect 33597 28509 33609 28512
rect 33643 28509 33655 28543
rect 33870 28540 33876 28552
rect 33831 28512 33876 28540
rect 33597 28503 33655 28509
rect 33870 28500 33876 28512
rect 33928 28500 33934 28552
rect 35544 28540 35572 28580
rect 35710 28568 35716 28580
rect 35768 28568 35774 28620
rect 36354 28608 36360 28620
rect 36315 28580 36360 28608
rect 36354 28568 36360 28580
rect 36412 28568 36418 28620
rect 36538 28608 36544 28620
rect 36499 28580 36544 28608
rect 36538 28568 36544 28580
rect 36596 28568 36602 28620
rect 38286 28608 38292 28620
rect 38247 28580 38292 28608
rect 38286 28568 38292 28580
rect 38344 28568 38350 28620
rect 38470 28608 38476 28620
rect 38431 28580 38476 28608
rect 38470 28568 38476 28580
rect 38528 28568 38534 28620
rect 38657 28611 38715 28617
rect 38657 28577 38669 28611
rect 38703 28608 38715 28611
rect 38838 28608 38844 28620
rect 38703 28580 38844 28608
rect 38703 28577 38715 28580
rect 38657 28571 38715 28577
rect 38838 28568 38844 28580
rect 38896 28568 38902 28620
rect 37829 28543 37887 28549
rect 37829 28540 37841 28543
rect 35544 28512 37841 28540
rect 37829 28509 37841 28512
rect 37875 28509 37887 28543
rect 37829 28503 37887 28509
rect 23808 28444 25452 28472
rect 32401 28475 32459 28481
rect 23808 28432 23814 28444
rect 32401 28441 32413 28475
rect 32447 28472 32459 28475
rect 33502 28472 33508 28484
rect 32447 28444 33508 28472
rect 32447 28441 32459 28444
rect 32401 28435 32459 28441
rect 33502 28432 33508 28444
rect 33560 28432 33566 28484
rect 16574 28404 16580 28416
rect 12728 28376 16580 28404
rect 16574 28364 16580 28376
rect 16632 28364 16638 28416
rect 16669 28407 16727 28413
rect 16669 28373 16681 28407
rect 16715 28404 16727 28407
rect 16758 28404 16764 28416
rect 16715 28376 16764 28404
rect 16715 28373 16727 28376
rect 16669 28367 16727 28373
rect 16758 28364 16764 28376
rect 16816 28364 16822 28416
rect 17681 28407 17739 28413
rect 17681 28373 17693 28407
rect 17727 28404 17739 28407
rect 19242 28404 19248 28416
rect 17727 28376 19248 28404
rect 17727 28373 17739 28376
rect 17681 28367 17739 28373
rect 19242 28364 19248 28376
rect 19300 28364 19306 28416
rect 19797 28407 19855 28413
rect 19797 28373 19809 28407
rect 19843 28404 19855 28407
rect 19978 28404 19984 28416
rect 19843 28376 19984 28404
rect 19843 28373 19855 28376
rect 19797 28367 19855 28373
rect 19978 28364 19984 28376
rect 20036 28364 20042 28416
rect 26602 28404 26608 28416
rect 26563 28376 26608 28404
rect 26602 28364 26608 28376
rect 26660 28364 26666 28416
rect 29365 28407 29423 28413
rect 29365 28373 29377 28407
rect 29411 28404 29423 28407
rect 29638 28404 29644 28416
rect 29411 28376 29644 28404
rect 29411 28373 29423 28376
rect 29365 28367 29423 28373
rect 29638 28364 29644 28376
rect 29696 28364 29702 28416
rect 33045 28407 33103 28413
rect 33045 28373 33057 28407
rect 33091 28404 33103 28407
rect 34238 28404 34244 28416
rect 33091 28376 34244 28404
rect 33091 28373 33103 28376
rect 33045 28367 33103 28373
rect 34238 28364 34244 28376
rect 34296 28364 34302 28416
rect 1104 28314 39836 28336
rect 1104 28262 4246 28314
rect 4298 28262 4310 28314
rect 4362 28262 4374 28314
rect 4426 28262 4438 28314
rect 4490 28262 34966 28314
rect 35018 28262 35030 28314
rect 35082 28262 35094 28314
rect 35146 28262 35158 28314
rect 35210 28262 39836 28314
rect 1104 28240 39836 28262
rect 9953 28203 10011 28209
rect 9953 28200 9965 28203
rect 4540 28172 9965 28200
rect 4062 28132 4068 28144
rect 2608 28104 4068 28132
rect 1949 27999 2007 28005
rect 1949 27965 1961 27999
rect 1995 27996 2007 27999
rect 2314 27996 2320 28008
rect 1995 27968 2320 27996
rect 1995 27965 2007 27968
rect 1949 27959 2007 27965
rect 2314 27956 2320 27968
rect 2372 27956 2378 28008
rect 2608 28005 2636 28104
rect 4062 28092 4068 28104
rect 4120 28092 4126 28144
rect 3234 28064 3240 28076
rect 3195 28036 3240 28064
rect 3234 28024 3240 28036
rect 3292 28024 3298 28076
rect 2593 27999 2651 28005
rect 2593 27965 2605 27999
rect 2639 27965 2651 27999
rect 2958 27996 2964 28008
rect 2919 27968 2964 27996
rect 2593 27959 2651 27965
rect 2958 27956 2964 27968
rect 3016 27956 3022 28008
rect 3326 27996 3332 28008
rect 3287 27968 3332 27996
rect 3326 27956 3332 27968
rect 3384 27956 3390 28008
rect 4065 27999 4123 28005
rect 4065 27965 4077 27999
rect 4111 27996 4123 27999
rect 4430 27996 4436 28008
rect 4111 27968 4436 27996
rect 4111 27965 4123 27968
rect 4065 27959 4123 27965
rect 4430 27956 4436 27968
rect 4488 27956 4494 28008
rect 4540 28005 4568 28172
rect 9953 28169 9965 28172
rect 9999 28169 10011 28203
rect 15470 28200 15476 28212
rect 15431 28172 15476 28200
rect 9953 28163 10011 28169
rect 15470 28160 15476 28172
rect 15528 28160 15534 28212
rect 16114 28200 16120 28212
rect 16075 28172 16120 28200
rect 16114 28160 16120 28172
rect 16172 28160 16178 28212
rect 16574 28160 16580 28212
rect 16632 28200 16638 28212
rect 24762 28200 24768 28212
rect 16632 28172 24768 28200
rect 16632 28160 16638 28172
rect 24762 28160 24768 28172
rect 24820 28160 24826 28212
rect 31754 28160 31760 28212
rect 31812 28200 31818 28212
rect 32766 28200 32772 28212
rect 31812 28172 32772 28200
rect 31812 28160 31818 28172
rect 32766 28160 32772 28172
rect 32824 28160 32830 28212
rect 35069 28203 35127 28209
rect 35069 28169 35081 28203
rect 35115 28200 35127 28203
rect 35802 28200 35808 28212
rect 35115 28172 35808 28200
rect 35115 28169 35127 28172
rect 35069 28163 35127 28169
rect 35802 28160 35808 28172
rect 35860 28160 35866 28212
rect 36814 28160 36820 28212
rect 36872 28200 36878 28212
rect 37369 28203 37427 28209
rect 37369 28200 37381 28203
rect 36872 28172 37381 28200
rect 36872 28160 36878 28172
rect 37369 28169 37381 28172
rect 37415 28169 37427 28203
rect 37369 28163 37427 28169
rect 5445 28135 5503 28141
rect 5445 28101 5457 28135
rect 5491 28132 5503 28135
rect 5718 28132 5724 28144
rect 5491 28104 5724 28132
rect 5491 28101 5503 28104
rect 5445 28095 5503 28101
rect 5718 28092 5724 28104
rect 5776 28092 5782 28144
rect 7009 28135 7067 28141
rect 7009 28101 7021 28135
rect 7055 28132 7067 28135
rect 7098 28132 7104 28144
rect 7055 28104 7104 28132
rect 7055 28101 7067 28104
rect 7009 28095 7067 28101
rect 7098 28092 7104 28104
rect 7156 28092 7162 28144
rect 11146 28132 11152 28144
rect 9600 28104 11152 28132
rect 4617 28067 4675 28073
rect 4617 28033 4629 28067
rect 4663 28064 4675 28067
rect 8021 28067 8079 28073
rect 8021 28064 8033 28067
rect 4663 28036 8033 28064
rect 4663 28033 4675 28036
rect 4617 28027 4675 28033
rect 8021 28033 8033 28036
rect 8067 28033 8079 28067
rect 9600 28064 9628 28104
rect 11146 28092 11152 28104
rect 11204 28092 11210 28144
rect 11330 28092 11336 28144
rect 11388 28132 11394 28144
rect 11388 28104 11652 28132
rect 11388 28092 11394 28104
rect 8021 28027 8079 28033
rect 9048 28036 9628 28064
rect 4525 27999 4583 28005
rect 4525 27965 4537 27999
rect 4571 27965 4583 27999
rect 4525 27959 4583 27965
rect 5353 27999 5411 28005
rect 5353 27965 5365 27999
rect 5399 27996 5411 27999
rect 5626 27996 5632 28008
rect 5399 27968 5632 27996
rect 5399 27965 5411 27968
rect 5353 27959 5411 27965
rect 5626 27956 5632 27968
rect 5684 27956 5690 28008
rect 5810 27996 5816 28008
rect 5771 27968 5816 27996
rect 5810 27956 5816 27968
rect 5868 27956 5874 28008
rect 5997 27999 6055 28005
rect 5997 27965 6009 27999
rect 6043 27965 6055 27999
rect 6822 27996 6828 28008
rect 6783 27968 6828 27996
rect 5997 27959 6055 27965
rect 5442 27888 5448 27940
rect 5500 27928 5506 27940
rect 6012 27928 6040 27959
rect 6822 27956 6828 27968
rect 6880 27956 6886 28008
rect 7745 27999 7803 28005
rect 7745 27965 7757 27999
rect 7791 27996 7803 27999
rect 9048 27996 9076 28036
rect 9674 28024 9680 28076
rect 9732 28064 9738 28076
rect 11624 28064 11652 28104
rect 12158 28092 12164 28144
rect 12216 28132 12222 28144
rect 16666 28132 16672 28144
rect 12216 28104 15332 28132
rect 16627 28104 16672 28132
rect 12216 28092 12222 28104
rect 14277 28067 14335 28073
rect 14277 28064 14289 28067
rect 9732 28036 11560 28064
rect 11624 28036 14289 28064
rect 9732 28024 9738 28036
rect 7791 27968 9076 27996
rect 7791 27965 7803 27968
rect 7745 27959 7803 27965
rect 9122 27956 9128 28008
rect 9180 27996 9186 28008
rect 11532 28005 11560 28036
rect 14277 28033 14289 28036
rect 14323 28033 14335 28067
rect 15304 28064 15332 28104
rect 16666 28092 16672 28104
rect 16724 28092 16730 28144
rect 18230 28092 18236 28144
rect 18288 28132 18294 28144
rect 18288 28104 19380 28132
rect 18288 28092 18294 28104
rect 19352 28073 19380 28104
rect 20530 28092 20536 28144
rect 20588 28132 20594 28144
rect 20717 28135 20775 28141
rect 20717 28132 20729 28135
rect 20588 28104 20729 28132
rect 20588 28092 20594 28104
rect 20717 28101 20729 28104
rect 20763 28101 20775 28135
rect 20717 28095 20775 28101
rect 22281 28135 22339 28141
rect 22281 28101 22293 28135
rect 22327 28132 22339 28135
rect 24578 28132 24584 28144
rect 22327 28104 24584 28132
rect 22327 28101 22339 28104
rect 22281 28095 22339 28101
rect 24578 28092 24584 28104
rect 24636 28092 24642 28144
rect 27798 28092 27804 28144
rect 27856 28132 27862 28144
rect 28077 28135 28135 28141
rect 28077 28132 28089 28135
rect 27856 28104 28089 28132
rect 27856 28092 27862 28104
rect 28077 28101 28089 28104
rect 28123 28101 28135 28135
rect 28077 28095 28135 28101
rect 30561 28135 30619 28141
rect 30561 28101 30573 28135
rect 30607 28132 30619 28135
rect 33042 28132 33048 28144
rect 30607 28104 33048 28132
rect 30607 28101 30619 28104
rect 30561 28095 30619 28101
rect 33042 28092 33048 28104
rect 33100 28092 33106 28144
rect 18509 28067 18567 28073
rect 15304 28036 18184 28064
rect 14277 28027 14335 28033
rect 9861 27999 9919 28005
rect 9861 27996 9873 27999
rect 9180 27968 9873 27996
rect 9180 27956 9186 27968
rect 9861 27965 9873 27968
rect 9907 27965 9919 27999
rect 9861 27959 9919 27965
rect 10229 27999 10287 28005
rect 10229 27965 10241 27999
rect 10275 27965 10287 27999
rect 10229 27959 10287 27965
rect 10873 27999 10931 28005
rect 10873 27965 10885 27999
rect 10919 27996 10931 27999
rect 11517 27999 11575 28005
rect 10919 27968 11468 27996
rect 10919 27965 10931 27968
rect 10873 27959 10931 27965
rect 5500 27900 6040 27928
rect 5500 27888 5506 27900
rect 8938 27888 8944 27940
rect 8996 27928 9002 27940
rect 10244 27928 10272 27959
rect 8996 27900 10272 27928
rect 11440 27928 11468 27968
rect 11517 27965 11529 27999
rect 11563 27965 11575 27999
rect 11517 27959 11575 27965
rect 11606 27956 11612 28008
rect 11664 27996 11670 28008
rect 12437 27999 12495 28005
rect 12437 27996 12449 27999
rect 11664 27968 12449 27996
rect 11664 27956 11670 27968
rect 12437 27965 12449 27968
rect 12483 27965 12495 27999
rect 13630 27996 13636 28008
rect 13543 27968 13636 27996
rect 12437 27959 12495 27965
rect 13630 27956 13636 27968
rect 13688 27956 13694 28008
rect 13998 27996 14004 28008
rect 13959 27968 14004 27996
rect 13998 27956 14004 27968
rect 14056 27956 14062 28008
rect 15378 27996 15384 28008
rect 15339 27968 15384 27996
rect 15378 27956 15384 27968
rect 15436 27956 15442 28008
rect 16298 27996 16304 28008
rect 16259 27968 16304 27996
rect 16298 27956 16304 27968
rect 16356 27956 16362 28008
rect 16390 27956 16396 28008
rect 16448 27996 16454 28008
rect 17034 27996 17040 28008
rect 16448 27968 16493 27996
rect 16995 27968 17040 27996
rect 16448 27956 16454 27968
rect 17034 27956 17040 27968
rect 17092 27956 17098 28008
rect 17218 27996 17224 28008
rect 17179 27968 17224 27996
rect 17218 27956 17224 27968
rect 17276 27956 17282 28008
rect 18156 28005 18184 28036
rect 18509 28033 18521 28067
rect 18555 28064 18567 28067
rect 19337 28067 19395 28073
rect 18555 28036 19288 28064
rect 18555 28033 18567 28036
rect 18509 28027 18567 28033
rect 18141 27999 18199 28005
rect 18141 27965 18153 27999
rect 18187 27965 18199 27999
rect 18141 27959 18199 27965
rect 18877 27999 18935 28005
rect 18877 27965 18889 27999
rect 18923 27965 18935 27999
rect 18877 27959 18935 27965
rect 12529 27931 12587 27937
rect 12529 27928 12541 27931
rect 11440 27900 12541 27928
rect 8996 27888 9002 27900
rect 12529 27897 12541 27900
rect 12575 27897 12587 27931
rect 13648 27928 13676 27956
rect 15562 27928 15568 27940
rect 13648 27900 15568 27928
rect 12529 27891 12587 27897
rect 15562 27888 15568 27900
rect 15620 27888 15626 27940
rect 2041 27863 2099 27869
rect 2041 27829 2053 27863
rect 2087 27860 2099 27863
rect 3878 27860 3884 27872
rect 2087 27832 3884 27860
rect 2087 27829 2099 27832
rect 2041 27823 2099 27829
rect 3878 27820 3884 27832
rect 3936 27820 3942 27872
rect 9306 27860 9312 27872
rect 9267 27832 9312 27860
rect 9306 27820 9312 27832
rect 9364 27820 9370 27872
rect 11606 27860 11612 27872
rect 11567 27832 11612 27860
rect 11606 27820 11612 27832
rect 11664 27820 11670 27872
rect 13541 27863 13599 27869
rect 13541 27829 13553 27863
rect 13587 27860 13599 27863
rect 14550 27860 14556 27872
rect 13587 27832 14556 27860
rect 13587 27829 13599 27832
rect 13541 27823 13599 27829
rect 14550 27820 14556 27832
rect 14608 27820 14614 27872
rect 18892 27860 18920 27959
rect 19260 27928 19288 28036
rect 19337 28033 19349 28067
rect 19383 28033 19395 28067
rect 22830 28064 22836 28076
rect 22791 28036 22836 28064
rect 19337 28027 19395 28033
rect 22830 28024 22836 28036
rect 22888 28024 22894 28076
rect 24210 28024 24216 28076
rect 24268 28064 24274 28076
rect 25869 28067 25927 28073
rect 24268 28036 24900 28064
rect 24268 28024 24274 28036
rect 19613 27999 19671 28005
rect 19613 27965 19625 27999
rect 19659 27996 19671 27999
rect 20346 27996 20352 28008
rect 19659 27968 20352 27996
rect 19659 27965 19671 27968
rect 19613 27959 19671 27965
rect 20346 27956 20352 27968
rect 20404 27956 20410 28008
rect 22005 27999 22063 28005
rect 22005 27965 22017 27999
rect 22051 27965 22063 27999
rect 22554 27996 22560 28008
rect 22515 27968 22560 27996
rect 22005 27959 22063 27965
rect 19426 27928 19432 27940
rect 19260 27900 19432 27928
rect 19426 27888 19432 27900
rect 19484 27888 19490 27940
rect 20990 27928 20996 27940
rect 20640 27900 20996 27928
rect 20640 27860 20668 27900
rect 20990 27888 20996 27900
rect 21048 27888 21054 27940
rect 22020 27928 22048 27959
rect 22554 27956 22560 27968
rect 22612 27956 22618 28008
rect 23750 27996 23756 28008
rect 23711 27968 23756 27996
rect 23750 27956 23756 27968
rect 23808 27956 23814 28008
rect 24305 27999 24363 28005
rect 24305 27965 24317 27999
rect 24351 27965 24363 27999
rect 24578 27996 24584 28008
rect 24539 27968 24584 27996
rect 24305 27959 24363 27965
rect 24026 27928 24032 27940
rect 22020 27900 24032 27928
rect 24026 27888 24032 27900
rect 24084 27888 24090 27940
rect 24320 27928 24348 27959
rect 24578 27956 24584 27968
rect 24636 27956 24642 28008
rect 24872 28005 24900 28036
rect 25869 28033 25881 28067
rect 25915 28064 25927 28067
rect 26050 28064 26056 28076
rect 25915 28036 26056 28064
rect 25915 28033 25927 28036
rect 25869 28027 25927 28033
rect 26050 28024 26056 28036
rect 26108 28024 26114 28076
rect 27246 28024 27252 28076
rect 27304 28064 27310 28076
rect 33134 28064 33140 28076
rect 27304 28036 28580 28064
rect 27304 28024 27310 28036
rect 24857 27999 24915 28005
rect 24857 27965 24869 27999
rect 24903 27965 24915 27999
rect 24857 27959 24915 27965
rect 26145 27999 26203 28005
rect 26145 27965 26157 27999
rect 26191 27996 26203 27999
rect 26234 27996 26240 28008
rect 26191 27968 26240 27996
rect 26191 27965 26203 27968
rect 26145 27959 26203 27965
rect 26234 27956 26240 27968
rect 26292 27956 26298 28008
rect 28552 28005 28580 28036
rect 31956 28036 33140 28064
rect 28261 27999 28319 28005
rect 28261 27965 28273 27999
rect 28307 27965 28319 27999
rect 28261 27959 28319 27965
rect 28537 27999 28595 28005
rect 28537 27965 28549 27999
rect 28583 27965 28595 27999
rect 29638 27996 29644 28008
rect 29599 27968 29644 27996
rect 28537 27959 28595 27965
rect 24670 27928 24676 27940
rect 24320 27900 24676 27928
rect 24670 27888 24676 27900
rect 24728 27888 24734 27940
rect 27525 27931 27583 27937
rect 27525 27897 27537 27931
rect 27571 27928 27583 27931
rect 27614 27928 27620 27940
rect 27571 27900 27620 27928
rect 27571 27897 27583 27900
rect 27525 27891 27583 27897
rect 27614 27888 27620 27900
rect 27672 27888 27678 27940
rect 28276 27928 28304 27959
rect 29638 27956 29644 27968
rect 29696 27956 29702 28008
rect 30193 27999 30251 28005
rect 30193 27965 30205 27999
rect 30239 27996 30251 27999
rect 30374 27996 30380 28008
rect 30239 27968 30380 27996
rect 30239 27965 30251 27968
rect 30193 27959 30251 27965
rect 30374 27956 30380 27968
rect 30432 27956 30438 28008
rect 30561 27999 30619 28005
rect 30561 27965 30573 27999
rect 30607 27996 30619 27999
rect 30742 27996 30748 28008
rect 30607 27968 30748 27996
rect 30607 27965 30619 27968
rect 30561 27959 30619 27965
rect 30742 27956 30748 27968
rect 30800 27956 30806 28008
rect 30926 27956 30932 28008
rect 30984 27996 30990 28008
rect 31956 28005 31984 28036
rect 33134 28024 33140 28036
rect 33192 28024 33198 28076
rect 35342 28064 35348 28076
rect 34992 28036 35348 28064
rect 31205 27999 31263 28005
rect 31205 27996 31217 27999
rect 30984 27968 31217 27996
rect 30984 27956 30990 27968
rect 31205 27965 31217 27968
rect 31251 27965 31263 27999
rect 31205 27959 31263 27965
rect 31941 27999 31999 28005
rect 31941 27965 31953 27999
rect 31987 27965 31999 27999
rect 31941 27959 31999 27965
rect 32217 27999 32275 28005
rect 32217 27965 32229 27999
rect 32263 27965 32275 27999
rect 32950 27996 32956 28008
rect 32911 27968 32956 27996
rect 32217 27959 32275 27965
rect 29362 27928 29368 27940
rect 28276 27900 29368 27928
rect 29362 27888 29368 27900
rect 29420 27888 29426 27940
rect 32232 27928 32260 27959
rect 32950 27956 32956 27968
rect 33008 27956 33014 28008
rect 33226 27996 33232 28008
rect 33187 27968 33232 27996
rect 33226 27956 33232 27968
rect 33284 27956 33290 28008
rect 33594 27996 33600 28008
rect 33555 27968 33600 27996
rect 33594 27956 33600 27968
rect 33652 27956 33658 28008
rect 34149 27999 34207 28005
rect 34149 27965 34161 27999
rect 34195 27996 34207 27999
rect 34514 27996 34520 28008
rect 34195 27968 34520 27996
rect 34195 27965 34207 27968
rect 34149 27959 34207 27965
rect 34514 27956 34520 27968
rect 34572 27956 34578 28008
rect 34992 28005 35020 28036
rect 35342 28024 35348 28036
rect 35400 28064 35406 28076
rect 36832 28064 36860 28160
rect 38286 28092 38292 28144
rect 38344 28132 38350 28144
rect 38749 28135 38807 28141
rect 38749 28132 38761 28135
rect 38344 28104 38761 28132
rect 38344 28092 38350 28104
rect 38749 28101 38761 28104
rect 38795 28101 38807 28135
rect 38749 28095 38807 28101
rect 35400 28036 36860 28064
rect 35400 28024 35406 28036
rect 37918 28024 37924 28076
rect 37976 28064 37982 28076
rect 38105 28067 38163 28073
rect 38105 28064 38117 28067
rect 37976 28036 38117 28064
rect 37976 28024 37982 28036
rect 38105 28033 38117 28036
rect 38151 28064 38163 28067
rect 38838 28064 38844 28076
rect 38151 28036 38844 28064
rect 38151 28033 38163 28036
rect 38105 28027 38163 28033
rect 38838 28024 38844 28036
rect 38896 28024 38902 28076
rect 34977 27999 35035 28005
rect 34977 27965 34989 27999
rect 35023 27965 35035 27999
rect 34977 27959 35035 27965
rect 35526 27956 35532 28008
rect 35584 27996 35590 28008
rect 35805 27999 35863 28005
rect 35805 27996 35817 27999
rect 35584 27968 35817 27996
rect 35584 27956 35590 27968
rect 35805 27965 35817 27968
rect 35851 27965 35863 27999
rect 35805 27959 35863 27965
rect 36081 27999 36139 28005
rect 36081 27965 36093 27999
rect 36127 27996 36139 27999
rect 37090 27996 37096 28008
rect 36127 27968 37096 27996
rect 36127 27965 36139 27968
rect 36081 27959 36139 27965
rect 37090 27956 37096 27968
rect 37148 27956 37154 28008
rect 38470 27996 38476 28008
rect 38431 27968 38476 27996
rect 38470 27956 38476 27968
rect 38528 27956 38534 28008
rect 38746 27996 38752 28008
rect 38707 27968 38752 27996
rect 38746 27956 38752 27968
rect 38804 27956 38810 28008
rect 34054 27928 34060 27940
rect 32232 27900 34060 27928
rect 34054 27888 34060 27900
rect 34112 27888 34118 27940
rect 34330 27928 34336 27940
rect 34291 27900 34336 27928
rect 34330 27888 34336 27900
rect 34388 27888 34394 27940
rect 18892 27832 20668 27860
rect 23937 27863 23995 27869
rect 23937 27829 23949 27863
rect 23983 27860 23995 27863
rect 24394 27860 24400 27872
rect 23983 27832 24400 27860
rect 23983 27829 23995 27832
rect 23937 27823 23995 27829
rect 24394 27820 24400 27832
rect 24452 27820 24458 27872
rect 31294 27860 31300 27872
rect 31255 27832 31300 27860
rect 31294 27820 31300 27832
rect 31352 27820 31358 27872
rect 1104 27770 39836 27792
rect 1104 27718 19606 27770
rect 19658 27718 19670 27770
rect 19722 27718 19734 27770
rect 19786 27718 19798 27770
rect 19850 27718 39836 27770
rect 1104 27696 39836 27718
rect 2958 27656 2964 27668
rect 2919 27628 2964 27656
rect 2958 27616 2964 27628
rect 3016 27616 3022 27668
rect 7098 27656 7104 27668
rect 3068 27628 7104 27656
rect 2682 27548 2688 27600
rect 2740 27588 2746 27600
rect 3068 27588 3096 27628
rect 7098 27616 7104 27628
rect 7156 27616 7162 27668
rect 8202 27616 8208 27668
rect 8260 27656 8266 27668
rect 17589 27659 17647 27665
rect 17589 27656 17601 27659
rect 8260 27628 10272 27656
rect 8260 27616 8266 27628
rect 2740 27560 3096 27588
rect 2740 27548 2746 27560
rect 1394 27520 1400 27532
rect 1355 27492 1400 27520
rect 1394 27480 1400 27492
rect 1452 27480 1458 27532
rect 1673 27523 1731 27529
rect 1673 27489 1685 27523
rect 1719 27520 1731 27523
rect 2406 27520 2412 27532
rect 1719 27492 2412 27520
rect 1719 27489 1731 27492
rect 1673 27483 1731 27489
rect 2406 27480 2412 27492
rect 2464 27480 2470 27532
rect 4341 27523 4399 27529
rect 4341 27489 4353 27523
rect 4387 27520 4399 27523
rect 4614 27520 4620 27532
rect 4387 27492 4620 27520
rect 4387 27489 4399 27492
rect 4341 27483 4399 27489
rect 4614 27480 4620 27492
rect 4672 27480 4678 27532
rect 6181 27523 6239 27529
rect 6181 27489 6193 27523
rect 6227 27489 6239 27523
rect 6181 27483 6239 27489
rect 7009 27523 7067 27529
rect 7009 27489 7021 27523
rect 7055 27520 7067 27523
rect 7558 27520 7564 27532
rect 7055 27492 7564 27520
rect 7055 27489 7067 27492
rect 7009 27483 7067 27489
rect 1412 27452 1440 27480
rect 2774 27452 2780 27464
rect 1412 27424 2780 27452
rect 2774 27412 2780 27424
rect 2832 27452 2838 27464
rect 4065 27455 4123 27461
rect 4065 27452 4077 27455
rect 2832 27424 4077 27452
rect 2832 27412 2838 27424
rect 4065 27421 4077 27424
rect 4111 27452 4123 27455
rect 5074 27452 5080 27464
rect 4111 27424 5080 27452
rect 4111 27421 4123 27424
rect 4065 27415 4123 27421
rect 5074 27412 5080 27424
rect 5132 27412 5138 27464
rect 6196 27452 6224 27483
rect 7558 27480 7564 27492
rect 7616 27520 7622 27532
rect 7653 27523 7711 27529
rect 7653 27520 7665 27523
rect 7616 27492 7665 27520
rect 7616 27480 7622 27492
rect 7653 27489 7665 27492
rect 7699 27489 7711 27523
rect 8662 27520 8668 27532
rect 8623 27492 8668 27520
rect 7653 27483 7711 27489
rect 8662 27480 8668 27492
rect 8720 27480 8726 27532
rect 9122 27520 9128 27532
rect 9083 27492 9128 27520
rect 9122 27480 9128 27492
rect 9180 27480 9186 27532
rect 10137 27523 10195 27529
rect 10137 27489 10149 27523
rect 10183 27489 10195 27523
rect 10137 27483 10195 27489
rect 6822 27452 6828 27464
rect 6196 27424 6828 27452
rect 6822 27412 6828 27424
rect 6880 27452 6886 27464
rect 7374 27452 7380 27464
rect 6880 27424 7380 27452
rect 6880 27412 6886 27424
rect 7374 27412 7380 27424
rect 7432 27452 7438 27464
rect 8757 27455 8815 27461
rect 7432 27424 7880 27452
rect 7432 27412 7438 27424
rect 7852 27393 7880 27424
rect 8757 27421 8769 27455
rect 8803 27452 8815 27455
rect 9674 27452 9680 27464
rect 8803 27424 9680 27452
rect 8803 27421 8815 27424
rect 8757 27415 8815 27421
rect 9674 27412 9680 27424
rect 9732 27412 9738 27464
rect 7837 27387 7895 27393
rect 7837 27353 7849 27387
rect 7883 27353 7895 27387
rect 10152 27384 10180 27483
rect 10244 27461 10272 27628
rect 15580 27628 17601 27656
rect 13998 27588 14004 27600
rect 13924 27560 14004 27588
rect 10410 27520 10416 27532
rect 10371 27492 10416 27520
rect 10410 27480 10416 27492
rect 10468 27480 10474 27532
rect 11057 27523 11115 27529
rect 11057 27489 11069 27523
rect 11103 27520 11115 27523
rect 11146 27520 11152 27532
rect 11103 27492 11152 27520
rect 11103 27489 11115 27492
rect 11057 27483 11115 27489
rect 11146 27480 11152 27492
rect 11204 27480 11210 27532
rect 11333 27523 11391 27529
rect 11333 27489 11345 27523
rect 11379 27520 11391 27523
rect 11606 27520 11612 27532
rect 11379 27492 11612 27520
rect 11379 27489 11391 27492
rect 11333 27483 11391 27489
rect 11606 27480 11612 27492
rect 11664 27480 11670 27532
rect 13357 27523 13415 27529
rect 13357 27489 13369 27523
rect 13403 27520 13415 27523
rect 13630 27520 13636 27532
rect 13403 27492 13636 27520
rect 13403 27489 13415 27492
rect 13357 27483 13415 27489
rect 13630 27480 13636 27492
rect 13688 27480 13694 27532
rect 13924 27529 13952 27560
rect 13998 27548 14004 27560
rect 14056 27548 14062 27600
rect 15580 27529 15608 27628
rect 17589 27625 17601 27628
rect 17635 27656 17647 27659
rect 18322 27656 18328 27668
rect 17635 27628 18328 27656
rect 17635 27625 17647 27628
rect 17589 27619 17647 27625
rect 18322 27616 18328 27628
rect 18380 27616 18386 27668
rect 19058 27656 19064 27668
rect 19019 27628 19064 27656
rect 19058 27616 19064 27628
rect 19116 27616 19122 27668
rect 20073 27659 20131 27665
rect 20073 27625 20085 27659
rect 20119 27656 20131 27659
rect 20622 27656 20628 27668
rect 20119 27628 20628 27656
rect 20119 27625 20131 27628
rect 20073 27619 20131 27625
rect 20622 27616 20628 27628
rect 20680 27616 20686 27668
rect 20990 27616 20996 27668
rect 21048 27656 21054 27668
rect 21085 27659 21143 27665
rect 21085 27656 21097 27659
rect 21048 27628 21097 27656
rect 21048 27616 21054 27628
rect 21085 27625 21097 27628
rect 21131 27656 21143 27659
rect 24670 27656 24676 27668
rect 21131 27628 24676 27656
rect 21131 27625 21143 27628
rect 21085 27619 21143 27625
rect 24670 27616 24676 27628
rect 24728 27616 24734 27668
rect 33870 27656 33876 27668
rect 33831 27628 33876 27656
rect 33870 27616 33876 27628
rect 33928 27616 33934 27668
rect 34514 27616 34520 27668
rect 34572 27656 34578 27668
rect 35621 27659 35679 27665
rect 35621 27656 35633 27659
rect 34572 27628 35633 27656
rect 34572 27616 34578 27628
rect 35621 27625 35633 27628
rect 35667 27625 35679 27659
rect 35621 27619 35679 27625
rect 36541 27659 36599 27665
rect 36541 27625 36553 27659
rect 36587 27656 36599 27659
rect 36630 27656 36636 27668
rect 36587 27628 36636 27656
rect 36587 27625 36599 27628
rect 36541 27619 36599 27625
rect 36630 27616 36636 27628
rect 36688 27616 36694 27668
rect 18138 27548 18144 27600
rect 18196 27588 18202 27600
rect 23842 27588 23848 27600
rect 18196 27560 23704 27588
rect 23803 27560 23848 27588
rect 18196 27548 18202 27560
rect 13909 27523 13967 27529
rect 13909 27489 13921 27523
rect 13955 27489 13967 27523
rect 13909 27483 13967 27489
rect 15565 27523 15623 27529
rect 15565 27489 15577 27523
rect 15611 27489 15623 27523
rect 15565 27483 15623 27489
rect 15657 27523 15715 27529
rect 15657 27489 15669 27523
rect 15703 27520 15715 27523
rect 16114 27520 16120 27532
rect 15703 27492 16120 27520
rect 15703 27489 15715 27492
rect 15657 27483 15715 27489
rect 16114 27480 16120 27492
rect 16172 27520 16178 27532
rect 17218 27520 17224 27532
rect 16172 27492 17224 27520
rect 16172 27480 16178 27492
rect 17218 27480 17224 27492
rect 17276 27480 17282 27532
rect 19061 27523 19119 27529
rect 19061 27489 19073 27523
rect 19107 27520 19119 27523
rect 19150 27520 19156 27532
rect 19107 27492 19156 27520
rect 19107 27489 19119 27492
rect 19061 27483 19119 27489
rect 19150 27480 19156 27492
rect 19208 27480 19214 27532
rect 19245 27523 19303 27529
rect 19245 27489 19257 27523
rect 19291 27489 19303 27523
rect 19245 27483 19303 27489
rect 10229 27455 10287 27461
rect 10229 27421 10241 27455
rect 10275 27452 10287 27455
rect 10870 27452 10876 27464
rect 10275 27424 10876 27452
rect 10275 27421 10287 27424
rect 10229 27415 10287 27421
rect 10870 27412 10876 27424
rect 10928 27412 10934 27464
rect 11422 27412 11428 27464
rect 11480 27452 11486 27464
rect 12713 27455 12771 27461
rect 12713 27452 12725 27455
rect 11480 27424 12725 27452
rect 11480 27412 11486 27424
rect 12713 27421 12725 27424
rect 12759 27452 12771 27455
rect 14001 27455 14059 27461
rect 14001 27452 14013 27455
rect 12759 27424 14013 27452
rect 12759 27421 12771 27424
rect 12713 27415 12771 27421
rect 14001 27421 14013 27424
rect 14047 27421 14059 27455
rect 14001 27415 14059 27421
rect 15746 27412 15752 27464
rect 15804 27452 15810 27464
rect 16209 27455 16267 27461
rect 16209 27452 16221 27455
rect 15804 27424 16221 27452
rect 15804 27412 15810 27424
rect 16209 27421 16221 27424
rect 16255 27421 16267 27455
rect 16209 27415 16267 27421
rect 16390 27412 16396 27464
rect 16448 27452 16454 27464
rect 16485 27455 16543 27461
rect 16485 27452 16497 27455
rect 16448 27424 16497 27452
rect 16448 27412 16454 27424
rect 16485 27421 16497 27424
rect 16531 27421 16543 27455
rect 19260 27452 19288 27483
rect 19334 27480 19340 27532
rect 19392 27520 19398 27532
rect 19981 27523 20039 27529
rect 19981 27520 19993 27523
rect 19392 27492 19993 27520
rect 19392 27480 19398 27492
rect 19981 27489 19993 27492
rect 20027 27489 20039 27523
rect 19981 27483 20039 27489
rect 20901 27523 20959 27529
rect 20901 27489 20913 27523
rect 20947 27520 20959 27523
rect 21634 27520 21640 27532
rect 20947 27492 21640 27520
rect 20947 27489 20959 27492
rect 20901 27483 20959 27489
rect 21634 27480 21640 27492
rect 21692 27480 21698 27532
rect 22097 27523 22155 27529
rect 22097 27489 22109 27523
rect 22143 27489 22155 27523
rect 22278 27520 22284 27532
rect 22239 27492 22284 27520
rect 22097 27483 22155 27489
rect 19886 27452 19892 27464
rect 19260 27424 19892 27452
rect 16485 27415 16543 27421
rect 19886 27412 19892 27424
rect 19944 27412 19950 27464
rect 22112 27452 22140 27483
rect 22278 27480 22284 27492
rect 22336 27480 22342 27532
rect 22462 27520 22468 27532
rect 22423 27492 22468 27520
rect 22462 27480 22468 27492
rect 22520 27480 22526 27532
rect 23109 27523 23167 27529
rect 23109 27489 23121 27523
rect 23155 27520 23167 27523
rect 23155 27492 23612 27520
rect 23155 27489 23167 27492
rect 23109 27483 23167 27489
rect 23014 27452 23020 27464
rect 22112 27424 23020 27452
rect 23014 27412 23020 27424
rect 23072 27412 23078 27464
rect 23198 27412 23204 27464
rect 23256 27452 23262 27464
rect 23477 27455 23535 27461
rect 23477 27452 23489 27455
rect 23256 27424 23489 27452
rect 23256 27412 23262 27424
rect 23477 27421 23489 27424
rect 23523 27421 23535 27455
rect 23477 27415 23535 27421
rect 13449 27387 13507 27393
rect 10152 27356 10272 27384
rect 7837 27347 7895 27353
rect 4062 27276 4068 27328
rect 4120 27316 4126 27328
rect 5629 27319 5687 27325
rect 5629 27316 5641 27319
rect 4120 27288 5641 27316
rect 4120 27276 4126 27288
rect 5629 27285 5641 27288
rect 5675 27285 5687 27319
rect 5629 27279 5687 27285
rect 5994 27276 6000 27328
rect 6052 27316 6058 27328
rect 6365 27319 6423 27325
rect 6365 27316 6377 27319
rect 6052 27288 6377 27316
rect 6052 27276 6058 27288
rect 6365 27285 6377 27288
rect 6411 27316 6423 27319
rect 6454 27316 6460 27328
rect 6411 27288 6460 27316
rect 6411 27285 6423 27288
rect 6365 27279 6423 27285
rect 6454 27276 6460 27288
rect 6512 27276 6518 27328
rect 7101 27319 7159 27325
rect 7101 27285 7113 27319
rect 7147 27316 7159 27319
rect 8110 27316 8116 27328
rect 7147 27288 8116 27316
rect 7147 27285 7159 27288
rect 7101 27279 7159 27285
rect 8110 27276 8116 27288
rect 8168 27316 8174 27328
rect 8386 27316 8392 27328
rect 8168 27288 8392 27316
rect 8168 27276 8174 27288
rect 8386 27276 8392 27288
rect 8444 27276 8450 27328
rect 10244 27316 10272 27356
rect 13449 27353 13461 27387
rect 13495 27384 13507 27387
rect 13906 27384 13912 27396
rect 13495 27356 13912 27384
rect 13495 27353 13507 27356
rect 13449 27347 13507 27353
rect 13906 27344 13912 27356
rect 13964 27344 13970 27396
rect 21913 27387 21971 27393
rect 21913 27353 21925 27387
rect 21959 27384 21971 27387
rect 22922 27384 22928 27396
rect 21959 27356 22928 27384
rect 21959 27353 21971 27356
rect 21913 27347 21971 27353
rect 22922 27344 22928 27356
rect 22980 27344 22986 27396
rect 12250 27316 12256 27328
rect 10244 27288 12256 27316
rect 12250 27276 12256 27288
rect 12308 27276 12314 27328
rect 22830 27276 22836 27328
rect 22888 27316 22894 27328
rect 23247 27319 23305 27325
rect 23247 27316 23259 27319
rect 22888 27288 23259 27316
rect 22888 27276 22894 27288
rect 23247 27285 23259 27288
rect 23293 27285 23305 27319
rect 23247 27279 23305 27285
rect 23385 27319 23443 27325
rect 23385 27285 23397 27319
rect 23431 27316 23443 27319
rect 23474 27316 23480 27328
rect 23431 27288 23480 27316
rect 23431 27285 23443 27288
rect 23385 27279 23443 27285
rect 23474 27276 23480 27288
rect 23532 27276 23538 27328
rect 23584 27316 23612 27492
rect 23676 27452 23704 27560
rect 23842 27548 23848 27560
rect 23900 27548 23906 27600
rect 24026 27548 24032 27600
rect 24084 27588 24090 27600
rect 24578 27588 24584 27600
rect 24084 27560 24584 27588
rect 24084 27548 24090 27560
rect 24578 27548 24584 27560
rect 24636 27548 24642 27600
rect 29362 27588 29368 27600
rect 29323 27560 29368 27588
rect 29362 27548 29368 27560
rect 29420 27548 29426 27600
rect 30926 27588 30932 27600
rect 30887 27560 30932 27588
rect 30926 27548 30932 27560
rect 30984 27548 30990 27600
rect 33226 27588 33232 27600
rect 32324 27560 33232 27588
rect 24394 27520 24400 27532
rect 24355 27492 24400 27520
rect 24394 27480 24400 27492
rect 24452 27480 24458 27532
rect 24486 27480 24492 27532
rect 24544 27520 24550 27532
rect 24765 27523 24823 27529
rect 24765 27520 24777 27523
rect 24544 27492 24777 27520
rect 24544 27480 24550 27492
rect 24765 27489 24777 27492
rect 24811 27489 24823 27523
rect 24765 27483 24823 27489
rect 25133 27523 25191 27529
rect 25133 27489 25145 27523
rect 25179 27489 25191 27523
rect 26602 27520 26608 27532
rect 26563 27492 26608 27520
rect 25133 27483 25191 27489
rect 25148 27452 25176 27483
rect 26602 27480 26608 27492
rect 26660 27480 26666 27532
rect 27065 27523 27123 27529
rect 27065 27489 27077 27523
rect 27111 27489 27123 27523
rect 27065 27483 27123 27489
rect 23676 27424 25176 27452
rect 25593 27455 25651 27461
rect 25593 27421 25605 27455
rect 25639 27452 25651 27455
rect 27080 27452 27108 27483
rect 27614 27480 27620 27532
rect 27672 27520 27678 27532
rect 29825 27523 29883 27529
rect 29825 27520 29837 27523
rect 27672 27492 29837 27520
rect 27672 27480 27678 27492
rect 29825 27489 29837 27492
rect 29871 27489 29883 27523
rect 29825 27483 29883 27489
rect 30285 27523 30343 27529
rect 30285 27489 30297 27523
rect 30331 27489 30343 27523
rect 30742 27520 30748 27532
rect 30703 27492 30748 27520
rect 30285 27483 30343 27489
rect 27706 27452 27712 27464
rect 25639 27424 27108 27452
rect 27667 27424 27712 27452
rect 25639 27421 25651 27424
rect 25593 27415 25651 27421
rect 27706 27412 27712 27424
rect 27764 27412 27770 27464
rect 27982 27452 27988 27464
rect 27943 27424 27988 27452
rect 27982 27412 27988 27424
rect 28040 27412 28046 27464
rect 30300 27452 30328 27483
rect 30742 27480 30748 27492
rect 30800 27480 30806 27532
rect 31386 27520 31392 27532
rect 31347 27492 31392 27520
rect 31386 27480 31392 27492
rect 31444 27480 31450 27532
rect 32324 27529 32352 27560
rect 33226 27548 33232 27560
rect 33284 27548 33290 27600
rect 35250 27548 35256 27600
rect 35308 27588 35314 27600
rect 36722 27588 36728 27600
rect 35308 27560 35572 27588
rect 36683 27560 36728 27588
rect 35308 27548 35314 27560
rect 32309 27523 32367 27529
rect 32309 27489 32321 27523
rect 32355 27489 32367 27523
rect 32490 27520 32496 27532
rect 32451 27492 32496 27520
rect 32309 27483 32367 27489
rect 32490 27480 32496 27492
rect 32548 27480 32554 27532
rect 32953 27523 33011 27529
rect 32953 27489 32965 27523
rect 32999 27489 33011 27523
rect 32953 27483 33011 27489
rect 30374 27452 30380 27464
rect 30287 27424 30380 27452
rect 30374 27412 30380 27424
rect 30432 27452 30438 27464
rect 31662 27452 31668 27464
rect 30432 27424 31668 27452
rect 30432 27412 30438 27424
rect 31662 27412 31668 27424
rect 31720 27412 31726 27464
rect 32968 27452 32996 27483
rect 33042 27480 33048 27532
rect 33100 27520 33106 27532
rect 33781 27523 33839 27529
rect 33781 27520 33793 27523
rect 33100 27492 33793 27520
rect 33100 27480 33106 27492
rect 33781 27489 33793 27492
rect 33827 27489 33839 27523
rect 34330 27520 34336 27532
rect 34291 27492 34336 27520
rect 33781 27483 33839 27489
rect 34330 27480 34336 27492
rect 34388 27480 34394 27532
rect 35342 27520 35348 27532
rect 35303 27492 35348 27520
rect 35342 27480 35348 27492
rect 35400 27480 35406 27532
rect 35544 27529 35572 27560
rect 36722 27548 36728 27560
rect 36780 27548 36786 27600
rect 37090 27588 37096 27600
rect 37051 27560 37096 27588
rect 37090 27548 37096 27560
rect 37148 27548 37154 27600
rect 35529 27523 35587 27529
rect 35529 27489 35541 27523
rect 35575 27489 35587 27523
rect 36633 27523 36691 27529
rect 36633 27520 36645 27523
rect 35529 27483 35587 27489
rect 35636 27492 36645 27520
rect 33594 27452 33600 27464
rect 32968 27424 33600 27452
rect 33594 27412 33600 27424
rect 33652 27412 33658 27464
rect 34054 27412 34060 27464
rect 34112 27452 34118 27464
rect 34609 27455 34667 27461
rect 34609 27452 34621 27455
rect 34112 27424 34621 27452
rect 34112 27412 34118 27424
rect 34609 27421 34621 27424
rect 34655 27421 34667 27455
rect 34609 27415 34667 27421
rect 26234 27344 26240 27396
rect 26292 27384 26298 27396
rect 26605 27387 26663 27393
rect 26605 27384 26617 27387
rect 26292 27356 26617 27384
rect 26292 27344 26298 27356
rect 26605 27353 26617 27356
rect 26651 27353 26663 27387
rect 26605 27347 26663 27353
rect 31481 27387 31539 27393
rect 31481 27353 31493 27387
rect 31527 27384 31539 27387
rect 31527 27356 33456 27384
rect 31527 27353 31539 27356
rect 31481 27347 31539 27353
rect 23842 27316 23848 27328
rect 23584 27288 23848 27316
rect 23842 27276 23848 27288
rect 23900 27276 23906 27328
rect 32214 27316 32220 27328
rect 32175 27288 32220 27316
rect 32214 27276 32220 27288
rect 32272 27276 32278 27328
rect 33428 27316 33456 27356
rect 33502 27344 33508 27396
rect 33560 27384 33566 27396
rect 35636 27384 35664 27492
rect 36633 27489 36645 27492
rect 36679 27520 36691 27523
rect 37737 27523 37795 27529
rect 37737 27520 37749 27523
rect 36679 27492 37749 27520
rect 36679 27489 36691 27492
rect 36633 27483 36691 27489
rect 37737 27489 37749 27492
rect 37783 27489 37795 27523
rect 37737 27483 37795 27489
rect 37918 27480 37924 27532
rect 37976 27520 37982 27532
rect 38289 27523 38347 27529
rect 38289 27520 38301 27523
rect 37976 27492 38301 27520
rect 37976 27480 37982 27492
rect 38289 27489 38301 27492
rect 38335 27489 38347 27523
rect 38289 27483 38347 27489
rect 38933 27523 38991 27529
rect 38933 27489 38945 27523
rect 38979 27489 38991 27523
rect 38933 27483 38991 27489
rect 36357 27455 36415 27461
rect 36357 27421 36369 27455
rect 36403 27452 36415 27455
rect 36446 27452 36452 27464
rect 36403 27424 36452 27452
rect 36403 27421 36415 27424
rect 36357 27415 36415 27421
rect 36446 27412 36452 27424
rect 36504 27412 36510 27464
rect 37182 27412 37188 27464
rect 37240 27452 37246 27464
rect 38948 27452 38976 27483
rect 37240 27424 38976 27452
rect 37240 27412 37246 27424
rect 39025 27387 39083 27393
rect 39025 27384 39037 27387
rect 33560 27356 35664 27384
rect 36740 27356 39037 27384
rect 33560 27344 33566 27356
rect 35710 27316 35716 27328
rect 33428 27288 35716 27316
rect 35710 27276 35716 27288
rect 35768 27276 35774 27328
rect 35802 27276 35808 27328
rect 35860 27316 35866 27328
rect 36740 27316 36768 27356
rect 39025 27353 39037 27356
rect 39071 27353 39083 27387
rect 39025 27347 39083 27353
rect 37826 27316 37832 27328
rect 35860 27288 36768 27316
rect 37787 27288 37832 27316
rect 35860 27276 35866 27288
rect 37826 27276 37832 27288
rect 37884 27276 37890 27328
rect 1104 27226 39836 27248
rect 1104 27174 4246 27226
rect 4298 27174 4310 27226
rect 4362 27174 4374 27226
rect 4426 27174 4438 27226
rect 4490 27174 34966 27226
rect 35018 27174 35030 27226
rect 35082 27174 35094 27226
rect 35146 27174 35158 27226
rect 35210 27174 39836 27226
rect 1104 27152 39836 27174
rect 2314 27112 2320 27124
rect 2275 27084 2320 27112
rect 2314 27072 2320 27084
rect 2372 27072 2378 27124
rect 8662 27072 8668 27124
rect 8720 27112 8726 27124
rect 9677 27115 9735 27121
rect 9677 27112 9689 27115
rect 8720 27084 9689 27112
rect 8720 27072 8726 27084
rect 9677 27081 9689 27084
rect 9723 27081 9735 27115
rect 11330 27112 11336 27124
rect 11291 27084 11336 27112
rect 9677 27075 9735 27081
rect 11330 27072 11336 27084
rect 11388 27072 11394 27124
rect 12529 27115 12587 27121
rect 12529 27081 12541 27115
rect 12575 27112 12587 27115
rect 12710 27112 12716 27124
rect 12575 27084 12716 27112
rect 12575 27081 12587 27084
rect 12529 27075 12587 27081
rect 12710 27072 12716 27084
rect 12768 27072 12774 27124
rect 14829 27115 14887 27121
rect 14829 27081 14841 27115
rect 14875 27112 14887 27115
rect 16390 27112 16396 27124
rect 14875 27084 16396 27112
rect 14875 27081 14887 27084
rect 14829 27075 14887 27081
rect 16390 27072 16396 27084
rect 16448 27072 16454 27124
rect 21082 27112 21088 27124
rect 21043 27084 21088 27112
rect 21082 27072 21088 27084
rect 21140 27072 21146 27124
rect 22922 27072 22928 27124
rect 22980 27112 22986 27124
rect 24486 27112 24492 27124
rect 22980 27084 24256 27112
rect 24447 27084 24492 27112
rect 22980 27072 22986 27084
rect 2958 27044 2964 27056
rect 2424 27016 2964 27044
rect 2424 26920 2452 27016
rect 2958 27004 2964 27016
rect 3016 27004 3022 27056
rect 4798 27004 4804 27056
rect 4856 27044 4862 27056
rect 5629 27047 5687 27053
rect 5629 27044 5641 27047
rect 4856 27016 5641 27044
rect 4856 27004 4862 27016
rect 5629 27013 5641 27016
rect 5675 27013 5687 27047
rect 5629 27007 5687 27013
rect 8481 27047 8539 27053
rect 8481 27013 8493 27047
rect 8527 27044 8539 27047
rect 8570 27044 8576 27056
rect 8527 27016 8576 27044
rect 8527 27013 8539 27016
rect 8481 27007 8539 27013
rect 8570 27004 8576 27016
rect 8628 27004 8634 27056
rect 13998 27044 14004 27056
rect 13372 27016 14004 27044
rect 3326 26976 3332 26988
rect 2884 26948 3332 26976
rect 2884 26920 2912 26948
rect 3326 26936 3332 26948
rect 3384 26936 3390 26988
rect 4433 26979 4491 26985
rect 4433 26945 4445 26979
rect 4479 26976 4491 26979
rect 4706 26976 4712 26988
rect 4479 26948 4712 26976
rect 4479 26945 4491 26948
rect 4433 26939 4491 26945
rect 4706 26936 4712 26948
rect 4764 26936 4770 26988
rect 9306 26976 9312 26988
rect 8680 26948 9312 26976
rect 2406 26908 2412 26920
rect 2319 26880 2412 26908
rect 2406 26868 2412 26880
rect 2464 26868 2470 26920
rect 2866 26908 2872 26920
rect 2779 26880 2872 26908
rect 2866 26868 2872 26880
rect 2924 26868 2930 26920
rect 3050 26908 3056 26920
rect 3011 26880 3056 26908
rect 3050 26868 3056 26880
rect 3108 26868 3114 26920
rect 3878 26908 3884 26920
rect 3839 26880 3884 26908
rect 3878 26868 3884 26880
rect 3936 26868 3942 26920
rect 4062 26908 4068 26920
rect 4023 26880 4068 26908
rect 4062 26868 4068 26880
rect 4120 26868 4126 26920
rect 4893 26911 4951 26917
rect 4893 26877 4905 26911
rect 4939 26877 4951 26911
rect 5534 26908 5540 26920
rect 5495 26880 5540 26908
rect 4893 26871 4951 26877
rect 4908 26840 4936 26871
rect 5534 26868 5540 26880
rect 5592 26868 5598 26920
rect 6273 26911 6331 26917
rect 6273 26877 6285 26911
rect 6319 26908 6331 26911
rect 6825 26911 6883 26917
rect 6825 26908 6837 26911
rect 6319 26880 6837 26908
rect 6319 26877 6331 26880
rect 6273 26871 6331 26877
rect 6825 26877 6837 26880
rect 6871 26877 6883 26911
rect 6825 26871 6883 26877
rect 7377 26911 7435 26917
rect 7377 26877 7389 26911
rect 7423 26877 7435 26911
rect 7377 26871 7435 26877
rect 7653 26911 7711 26917
rect 7653 26877 7665 26911
rect 7699 26877 7711 26911
rect 7834 26908 7840 26920
rect 7795 26880 7840 26908
rect 7653 26871 7711 26877
rect 6178 26840 6184 26852
rect 4908 26812 6184 26840
rect 6178 26800 6184 26812
rect 6236 26800 6242 26852
rect 4982 26772 4988 26784
rect 4943 26744 4988 26772
rect 4982 26732 4988 26744
rect 5040 26732 5046 26784
rect 7392 26772 7420 26871
rect 7668 26840 7696 26871
rect 7834 26868 7840 26880
rect 7892 26868 7898 26920
rect 8680 26917 8708 26948
rect 9306 26936 9312 26948
rect 9364 26976 9370 26988
rect 13372 26985 13400 27016
rect 13998 27004 14004 27016
rect 14056 27004 14062 27056
rect 14093 27047 14151 27053
rect 14093 27013 14105 27047
rect 14139 27044 14151 27047
rect 18138 27044 18144 27056
rect 14139 27016 18144 27044
rect 14139 27013 14151 27016
rect 14093 27007 14151 27013
rect 18138 27004 18144 27016
rect 18196 27004 18202 27056
rect 20438 27004 20444 27056
rect 20496 27044 20502 27056
rect 20622 27044 20628 27056
rect 20496 27016 20628 27044
rect 20496 27004 20502 27016
rect 20622 27004 20628 27016
rect 20680 27004 20686 27056
rect 24118 27044 24124 27056
rect 24079 27016 24124 27044
rect 24118 27004 24124 27016
rect 24176 27004 24182 27056
rect 24228 27044 24256 27084
rect 24486 27072 24492 27084
rect 24544 27072 24550 27124
rect 29270 27072 29276 27124
rect 29328 27112 29334 27124
rect 29365 27115 29423 27121
rect 29365 27112 29377 27115
rect 29328 27084 29377 27112
rect 29328 27072 29334 27084
rect 29365 27081 29377 27084
rect 29411 27081 29423 27115
rect 29365 27075 29423 27081
rect 30006 27072 30012 27124
rect 30064 27112 30070 27124
rect 31021 27115 31079 27121
rect 31021 27112 31033 27115
rect 30064 27084 31033 27112
rect 30064 27072 30070 27084
rect 31021 27081 31033 27084
rect 31067 27112 31079 27115
rect 32490 27112 32496 27124
rect 31067 27084 32496 27112
rect 31067 27081 31079 27084
rect 31021 27075 31079 27081
rect 32490 27072 32496 27084
rect 32548 27072 32554 27124
rect 33137 27115 33195 27121
rect 33137 27081 33149 27115
rect 33183 27112 33195 27115
rect 33226 27112 33232 27124
rect 33183 27084 33232 27112
rect 33183 27081 33195 27084
rect 33137 27075 33195 27081
rect 33226 27072 33232 27084
rect 33284 27072 33290 27124
rect 34514 27072 34520 27124
rect 34572 27112 34578 27124
rect 35802 27112 35808 27124
rect 34572 27084 35808 27112
rect 34572 27072 34578 27084
rect 35802 27072 35808 27084
rect 35860 27072 35866 27124
rect 38838 27112 38844 27124
rect 38799 27084 38844 27112
rect 38838 27072 38844 27084
rect 38896 27072 38902 27124
rect 35069 27047 35127 27053
rect 35069 27044 35081 27047
rect 24228 27016 28120 27044
rect 13357 26979 13415 26985
rect 9364 26948 11284 26976
rect 9364 26936 9370 26948
rect 9876 26917 9904 26948
rect 8665 26911 8723 26917
rect 8665 26877 8677 26911
rect 8711 26877 8723 26911
rect 8665 26871 8723 26877
rect 9125 26911 9183 26917
rect 9125 26877 9137 26911
rect 9171 26877 9183 26911
rect 9125 26871 9183 26877
rect 9861 26911 9919 26917
rect 9861 26877 9873 26911
rect 9907 26877 9919 26911
rect 9861 26871 9919 26877
rect 10229 26911 10287 26917
rect 10229 26877 10241 26911
rect 10275 26877 10287 26911
rect 10502 26908 10508 26920
rect 10463 26880 10508 26908
rect 10229 26871 10287 26877
rect 8110 26840 8116 26852
rect 7668 26812 8116 26840
rect 8110 26800 8116 26812
rect 8168 26800 8174 26852
rect 9140 26840 9168 26871
rect 10244 26840 10272 26871
rect 10502 26868 10508 26880
rect 10560 26868 10566 26920
rect 11256 26917 11284 26948
rect 13357 26945 13369 26979
rect 13403 26945 13415 26979
rect 17037 26979 17095 26985
rect 17037 26976 17049 26979
rect 13357 26939 13415 26945
rect 14752 26948 17049 26976
rect 11241 26911 11299 26917
rect 11241 26877 11253 26911
rect 11287 26877 11299 26911
rect 11241 26871 11299 26877
rect 12434 26868 12440 26920
rect 12492 26908 12498 26920
rect 13538 26908 13544 26920
rect 12492 26880 12537 26908
rect 13499 26880 13544 26908
rect 12492 26868 12498 26880
rect 13538 26868 13544 26880
rect 13596 26868 13602 26920
rect 13906 26868 13912 26920
rect 13964 26908 13970 26920
rect 14752 26917 14780 26948
rect 17037 26945 17049 26948
rect 17083 26945 17095 26979
rect 18966 26976 18972 26988
rect 18927 26948 18972 26976
rect 17037 26939 17095 26945
rect 18966 26936 18972 26948
rect 19024 26936 19030 26988
rect 20530 26976 20536 26988
rect 19536 26948 20536 26976
rect 14001 26911 14059 26917
rect 14001 26908 14013 26911
rect 13964 26880 14013 26908
rect 13964 26868 13970 26880
rect 14001 26877 14013 26880
rect 14047 26877 14059 26911
rect 14001 26871 14059 26877
rect 14737 26911 14795 26917
rect 14737 26877 14749 26911
rect 14783 26877 14795 26911
rect 14737 26871 14795 26877
rect 15381 26911 15439 26917
rect 15381 26877 15393 26911
rect 15427 26908 15439 26911
rect 15470 26908 15476 26920
rect 15427 26880 15476 26908
rect 15427 26877 15439 26880
rect 15381 26871 15439 26877
rect 15470 26868 15476 26880
rect 15528 26868 15534 26920
rect 16114 26908 16120 26920
rect 16075 26880 16120 26908
rect 16114 26868 16120 26880
rect 16172 26868 16178 26920
rect 16485 26911 16543 26917
rect 16485 26877 16497 26911
rect 16531 26908 16543 26911
rect 16531 26880 16620 26908
rect 16531 26877 16543 26880
rect 16485 26871 16543 26877
rect 11422 26840 11428 26852
rect 9140 26812 11428 26840
rect 11422 26800 11428 26812
rect 11480 26800 11486 26852
rect 13814 26800 13820 26852
rect 13872 26840 13878 26852
rect 16022 26840 16028 26852
rect 13872 26812 16028 26840
rect 13872 26800 13878 26812
rect 16022 26800 16028 26812
rect 16080 26800 16086 26852
rect 8846 26772 8852 26784
rect 7392 26744 8852 26772
rect 8846 26732 8852 26744
rect 8904 26772 8910 26784
rect 10778 26772 10784 26784
rect 8904 26744 10784 26772
rect 8904 26732 8910 26744
rect 10778 26732 10784 26744
rect 10836 26732 10842 26784
rect 15562 26772 15568 26784
rect 15523 26744 15568 26772
rect 15562 26732 15568 26744
rect 15620 26732 15626 26784
rect 16592 26772 16620 26880
rect 16666 26868 16672 26920
rect 16724 26908 16730 26920
rect 16945 26911 17003 26917
rect 16945 26908 16957 26911
rect 16724 26880 16957 26908
rect 16724 26868 16730 26880
rect 16945 26877 16957 26880
rect 16991 26877 17003 26911
rect 16945 26871 17003 26877
rect 18877 26911 18935 26917
rect 18877 26877 18889 26911
rect 18923 26877 18935 26911
rect 19058 26908 19064 26920
rect 19019 26880 19064 26908
rect 18877 26871 18935 26877
rect 18892 26840 18920 26871
rect 19058 26868 19064 26880
rect 19116 26868 19122 26920
rect 19426 26868 19432 26920
rect 19484 26908 19490 26920
rect 19536 26917 19564 26948
rect 20530 26936 20536 26948
rect 20588 26936 20594 26988
rect 24213 26979 24271 26985
rect 22112 26948 22876 26976
rect 19521 26911 19579 26917
rect 19521 26908 19533 26911
rect 19484 26880 19533 26908
rect 19484 26868 19490 26880
rect 19521 26877 19533 26880
rect 19567 26877 19579 26911
rect 20070 26908 20076 26920
rect 20031 26880 20076 26908
rect 19521 26871 19579 26877
rect 20070 26868 20076 26880
rect 20128 26868 20134 26920
rect 20438 26908 20444 26920
rect 20399 26880 20444 26908
rect 20438 26868 20444 26880
rect 20496 26868 20502 26920
rect 20806 26868 20812 26920
rect 20864 26908 20870 26920
rect 20993 26911 21051 26917
rect 20993 26908 21005 26911
rect 20864 26880 21005 26908
rect 20864 26868 20870 26880
rect 20993 26877 21005 26880
rect 21039 26877 21051 26911
rect 20993 26871 21051 26877
rect 21729 26911 21787 26917
rect 21729 26877 21741 26911
rect 21775 26908 21787 26911
rect 21910 26908 21916 26920
rect 21775 26880 21916 26908
rect 21775 26877 21787 26880
rect 21729 26871 21787 26877
rect 21910 26868 21916 26880
rect 21968 26868 21974 26920
rect 22112 26917 22140 26948
rect 22848 26920 22876 26948
rect 24213 26945 24225 26979
rect 24259 26945 24271 26979
rect 24213 26939 24271 26945
rect 27709 26979 27767 26985
rect 27709 26945 27721 26979
rect 27755 26976 27767 26979
rect 27982 26976 27988 26988
rect 27755 26948 27988 26976
rect 27755 26945 27767 26948
rect 27709 26939 27767 26945
rect 22097 26911 22155 26917
rect 22097 26877 22109 26911
rect 22143 26877 22155 26911
rect 22278 26908 22284 26920
rect 22239 26880 22284 26908
rect 22097 26871 22155 26877
rect 22278 26868 22284 26880
rect 22336 26868 22342 26920
rect 22649 26911 22707 26917
rect 22649 26877 22661 26911
rect 22695 26877 22707 26911
rect 22649 26871 22707 26877
rect 19978 26840 19984 26852
rect 18892 26812 19984 26840
rect 19978 26800 19984 26812
rect 20036 26840 20042 26852
rect 22664 26840 22692 26871
rect 22830 26868 22836 26920
rect 22888 26908 22894 26920
rect 23992 26911 24050 26917
rect 23992 26908 24004 26911
rect 22888 26880 24004 26908
rect 22888 26868 22894 26880
rect 23992 26877 24004 26880
rect 24038 26877 24050 26911
rect 23992 26871 24050 26877
rect 23842 26840 23848 26852
rect 20036 26812 22692 26840
rect 23803 26812 23848 26840
rect 20036 26800 20042 26812
rect 23842 26800 23848 26812
rect 23900 26800 23906 26852
rect 17034 26772 17040 26784
rect 16592 26744 17040 26772
rect 17034 26732 17040 26744
rect 17092 26772 17098 26784
rect 17494 26772 17500 26784
rect 17092 26744 17500 26772
rect 17092 26732 17098 26744
rect 17494 26732 17500 26744
rect 17552 26732 17558 26784
rect 18506 26732 18512 26784
rect 18564 26772 18570 26784
rect 24228 26772 24256 26939
rect 27982 26936 27988 26948
rect 28040 26936 28046 26988
rect 25590 26908 25596 26920
rect 25551 26880 25596 26908
rect 25590 26868 25596 26880
rect 25648 26868 25654 26920
rect 27525 26911 27583 26917
rect 27525 26877 27537 26911
rect 27571 26908 27583 26911
rect 27798 26908 27804 26920
rect 27571 26880 27804 26908
rect 27571 26877 27583 26880
rect 27525 26871 27583 26877
rect 27798 26868 27804 26880
rect 27856 26868 27862 26920
rect 28092 26917 28120 27016
rect 33704 27016 35081 27044
rect 28626 26936 28632 26988
rect 28684 26976 28690 26988
rect 28684 26948 29868 26976
rect 28684 26936 28690 26948
rect 28077 26911 28135 26917
rect 28077 26877 28089 26911
rect 28123 26877 28135 26911
rect 28534 26908 28540 26920
rect 28495 26880 28540 26908
rect 28077 26871 28135 26877
rect 28534 26868 28540 26880
rect 28592 26868 28598 26920
rect 29546 26908 29552 26920
rect 29507 26880 29552 26908
rect 29546 26868 29552 26880
rect 29604 26868 29610 26920
rect 29840 26917 29868 26948
rect 32306 26936 32312 26988
rect 32364 26976 32370 26988
rect 33704 26976 33732 27016
rect 35069 27013 35081 27016
rect 35115 27044 35127 27047
rect 35621 27047 35679 27053
rect 35621 27044 35633 27047
rect 35115 27016 35633 27044
rect 35115 27013 35127 27016
rect 35069 27007 35127 27013
rect 35621 27013 35633 27016
rect 35667 27013 35679 27047
rect 35621 27007 35679 27013
rect 32364 26948 33732 26976
rect 32364 26936 32370 26948
rect 34238 26936 34244 26988
rect 34296 26976 34302 26988
rect 37737 26979 37795 26985
rect 37737 26976 37749 26979
rect 34296 26948 37749 26976
rect 34296 26936 34302 26948
rect 37737 26945 37749 26948
rect 37783 26945 37795 26979
rect 37737 26939 37795 26945
rect 29825 26911 29883 26917
rect 29825 26877 29837 26911
rect 29871 26877 29883 26911
rect 30834 26908 30840 26920
rect 30795 26880 30840 26908
rect 29825 26871 29883 26877
rect 30834 26868 30840 26880
rect 30892 26868 30898 26920
rect 31570 26908 31576 26920
rect 31531 26880 31576 26908
rect 31570 26868 31576 26880
rect 31628 26868 31634 26920
rect 31846 26908 31852 26920
rect 31807 26880 31852 26908
rect 31846 26868 31852 26880
rect 31904 26868 31910 26920
rect 33686 26908 33692 26920
rect 33647 26880 33692 26908
rect 33686 26868 33692 26880
rect 33744 26868 33750 26920
rect 33873 26911 33931 26917
rect 33873 26877 33885 26911
rect 33919 26908 33931 26911
rect 34790 26908 34796 26920
rect 33919 26880 34796 26908
rect 33919 26877 33931 26880
rect 33873 26871 33931 26877
rect 34790 26868 34796 26880
rect 34848 26908 34854 26920
rect 34885 26911 34943 26917
rect 34885 26908 34897 26911
rect 34848 26880 34897 26908
rect 34848 26868 34854 26880
rect 34885 26877 34897 26880
rect 34931 26877 34943 26911
rect 34885 26871 34943 26877
rect 35621 26911 35679 26917
rect 35621 26877 35633 26911
rect 35667 26908 35679 26911
rect 35713 26911 35771 26917
rect 35713 26908 35725 26911
rect 35667 26880 35725 26908
rect 35667 26877 35679 26880
rect 35621 26871 35679 26877
rect 35713 26877 35725 26880
rect 35759 26877 35771 26911
rect 35713 26871 35771 26877
rect 36265 26911 36323 26917
rect 36265 26877 36277 26911
rect 36311 26908 36323 26911
rect 36630 26908 36636 26920
rect 36311 26880 36636 26908
rect 36311 26877 36323 26880
rect 36265 26871 36323 26877
rect 36630 26868 36636 26880
rect 36688 26868 36694 26920
rect 37458 26908 37464 26920
rect 37419 26880 37464 26908
rect 37458 26868 37464 26880
rect 37516 26868 37522 26920
rect 18564 26744 24256 26772
rect 18564 26732 18570 26744
rect 25406 26732 25412 26784
rect 25464 26772 25470 26784
rect 25685 26775 25743 26781
rect 25685 26772 25697 26775
rect 25464 26744 25697 26772
rect 25464 26732 25470 26744
rect 25685 26741 25697 26744
rect 25731 26741 25743 26775
rect 25685 26735 25743 26741
rect 28629 26775 28687 26781
rect 28629 26741 28641 26775
rect 28675 26772 28687 26775
rect 30098 26772 30104 26784
rect 28675 26744 30104 26772
rect 28675 26741 28687 26744
rect 28629 26735 28687 26741
rect 30098 26732 30104 26744
rect 30156 26732 30162 26784
rect 33502 26732 33508 26784
rect 33560 26772 33566 26784
rect 33965 26775 34023 26781
rect 33965 26772 33977 26775
rect 33560 26744 33977 26772
rect 33560 26732 33566 26744
rect 33965 26741 33977 26744
rect 34011 26741 34023 26775
rect 35802 26772 35808 26784
rect 35763 26744 35808 26772
rect 33965 26735 34023 26741
rect 35802 26732 35808 26744
rect 35860 26732 35866 26784
rect 1104 26682 39836 26704
rect 1104 26630 19606 26682
rect 19658 26630 19670 26682
rect 19722 26630 19734 26682
rect 19786 26630 19798 26682
rect 19850 26630 39836 26682
rect 1104 26608 39836 26630
rect 7742 26528 7748 26580
rect 7800 26568 7806 26580
rect 8297 26571 8355 26577
rect 8297 26568 8309 26571
rect 7800 26540 8309 26568
rect 7800 26528 7806 26540
rect 8297 26537 8309 26540
rect 8343 26537 8355 26571
rect 8297 26531 8355 26537
rect 8754 26528 8760 26580
rect 8812 26568 8818 26580
rect 9030 26568 9036 26580
rect 8812 26540 9036 26568
rect 8812 26528 8818 26540
rect 9030 26528 9036 26540
rect 9088 26568 9094 26580
rect 13814 26568 13820 26580
rect 9088 26540 13820 26568
rect 9088 26528 9094 26540
rect 13814 26528 13820 26540
rect 13872 26528 13878 26580
rect 13998 26528 14004 26580
rect 14056 26568 14062 26580
rect 14553 26571 14611 26577
rect 14553 26568 14565 26571
rect 14056 26540 14565 26568
rect 14056 26528 14062 26540
rect 14553 26537 14565 26540
rect 14599 26537 14611 26571
rect 14553 26531 14611 26537
rect 16206 26528 16212 26580
rect 16264 26528 16270 26580
rect 20438 26568 20444 26580
rect 18248 26540 20444 26568
rect 1946 26500 1952 26512
rect 1907 26472 1952 26500
rect 1946 26460 1952 26472
rect 2004 26460 2010 26512
rect 9122 26460 9128 26512
rect 9180 26500 9186 26512
rect 10413 26503 10471 26509
rect 10413 26500 10425 26503
rect 9180 26472 10425 26500
rect 9180 26460 9186 26472
rect 10413 26469 10425 26472
rect 10459 26469 10471 26503
rect 10413 26463 10471 26469
rect 12250 26460 12256 26512
rect 12308 26500 12314 26512
rect 15378 26500 15384 26512
rect 12308 26472 13676 26500
rect 12308 26460 12314 26472
rect 2406 26432 2412 26444
rect 2367 26404 2412 26432
rect 2406 26392 2412 26404
rect 2464 26392 2470 26444
rect 2777 26435 2835 26441
rect 2777 26401 2789 26435
rect 2823 26401 2835 26435
rect 2777 26395 2835 26401
rect 2792 26364 2820 26395
rect 2866 26392 2872 26444
rect 2924 26432 2930 26444
rect 2924 26404 2969 26432
rect 2924 26392 2930 26404
rect 3970 26392 3976 26444
rect 4028 26432 4034 26444
rect 4065 26435 4123 26441
rect 4065 26432 4077 26435
rect 4028 26404 4077 26432
rect 4028 26392 4034 26404
rect 4065 26401 4077 26404
rect 4111 26401 4123 26435
rect 4798 26432 4804 26444
rect 4759 26404 4804 26432
rect 4065 26395 4123 26401
rect 4798 26392 4804 26404
rect 4856 26392 4862 26444
rect 4893 26435 4951 26441
rect 4893 26401 4905 26435
rect 4939 26432 4951 26435
rect 5721 26435 5779 26441
rect 5721 26432 5733 26435
rect 4939 26404 5733 26432
rect 4939 26401 4951 26404
rect 4893 26395 4951 26401
rect 5721 26401 5733 26404
rect 5767 26401 5779 26435
rect 8202 26432 8208 26444
rect 8163 26404 8208 26432
rect 5721 26395 5779 26401
rect 8202 26392 8208 26404
rect 8260 26392 8266 26444
rect 8573 26435 8631 26441
rect 8573 26401 8585 26435
rect 8619 26432 8631 26435
rect 8662 26432 8668 26444
rect 8619 26404 8668 26432
rect 8619 26401 8631 26404
rect 8573 26395 8631 26401
rect 8662 26392 8668 26404
rect 8720 26392 8726 26444
rect 9677 26435 9735 26441
rect 9677 26401 9689 26435
rect 9723 26432 9735 26435
rect 11054 26432 11060 26444
rect 9723 26404 11060 26432
rect 9723 26401 9735 26404
rect 9677 26395 9735 26401
rect 11054 26392 11060 26404
rect 11112 26392 11118 26444
rect 11238 26432 11244 26444
rect 11199 26404 11244 26432
rect 11238 26392 11244 26404
rect 11296 26392 11302 26444
rect 11422 26432 11428 26444
rect 11383 26404 11428 26432
rect 11422 26392 11428 26404
rect 11480 26392 11486 26444
rect 11514 26392 11520 26444
rect 11572 26432 11578 26444
rect 13648 26441 13676 26472
rect 14384 26472 15384 26500
rect 14384 26441 14412 26472
rect 15378 26460 15384 26472
rect 15436 26500 15442 26512
rect 15436 26472 15884 26500
rect 15436 26460 15442 26472
rect 11885 26435 11943 26441
rect 11885 26432 11897 26435
rect 11572 26404 11897 26432
rect 11572 26392 11578 26404
rect 11885 26401 11897 26404
rect 11931 26401 11943 26435
rect 11885 26395 11943 26401
rect 12989 26435 13047 26441
rect 12989 26401 13001 26435
rect 13035 26432 13047 26435
rect 13541 26435 13599 26441
rect 13035 26404 13492 26432
rect 13035 26401 13047 26404
rect 12989 26395 13047 26401
rect 2958 26364 2964 26376
rect 2792 26336 2964 26364
rect 2958 26324 2964 26336
rect 3016 26324 3022 26376
rect 5074 26324 5080 26376
rect 5132 26364 5138 26376
rect 5445 26367 5503 26373
rect 5445 26364 5457 26367
rect 5132 26336 5457 26364
rect 5132 26324 5138 26336
rect 5445 26333 5457 26336
rect 5491 26333 5503 26367
rect 5445 26327 5503 26333
rect 7101 26367 7159 26373
rect 7101 26333 7113 26367
rect 7147 26333 7159 26367
rect 7101 26327 7159 26333
rect 4249 26231 4307 26237
rect 4249 26197 4261 26231
rect 4295 26228 4307 26231
rect 5074 26228 5080 26240
rect 4295 26200 5080 26228
rect 4295 26197 4307 26200
rect 4249 26191 4307 26197
rect 5074 26188 5080 26200
rect 5132 26188 5138 26240
rect 6822 26188 6828 26240
rect 6880 26228 6886 26240
rect 7116 26228 7144 26327
rect 10778 26324 10784 26376
rect 10836 26364 10842 26376
rect 10965 26367 11023 26373
rect 10965 26364 10977 26367
rect 10836 26336 10977 26364
rect 10836 26324 10842 26336
rect 10965 26333 10977 26336
rect 11011 26333 11023 26367
rect 10965 26327 11023 26333
rect 9766 26296 9772 26308
rect 9727 26268 9772 26296
rect 9766 26256 9772 26268
rect 9824 26256 9830 26308
rect 11974 26296 11980 26308
rect 11935 26268 11980 26296
rect 11974 26256 11980 26268
rect 12032 26256 12038 26308
rect 13081 26299 13139 26305
rect 13081 26265 13093 26299
rect 13127 26296 13139 26299
rect 13262 26296 13268 26308
rect 13127 26268 13268 26296
rect 13127 26265 13139 26268
rect 13081 26259 13139 26265
rect 13262 26256 13268 26268
rect 13320 26256 13326 26308
rect 13464 26296 13492 26404
rect 13541 26401 13553 26435
rect 13587 26401 13599 26435
rect 13541 26395 13599 26401
rect 13633 26435 13691 26441
rect 13633 26401 13645 26435
rect 13679 26401 13691 26435
rect 13633 26395 13691 26401
rect 14369 26435 14427 26441
rect 14369 26401 14381 26435
rect 14415 26401 14427 26435
rect 14369 26395 14427 26401
rect 15749 26435 15807 26441
rect 15749 26401 15761 26435
rect 15795 26401 15807 26435
rect 15856 26432 15884 26472
rect 16224 26441 16252 26528
rect 18248 26500 18276 26540
rect 20438 26528 20444 26540
rect 20496 26568 20502 26580
rect 21085 26571 21143 26577
rect 21085 26568 21097 26571
rect 20496 26540 21097 26568
rect 20496 26528 20502 26540
rect 21085 26537 21097 26540
rect 21131 26568 21143 26571
rect 21131 26540 23704 26568
rect 21131 26537 21143 26540
rect 21085 26531 21143 26537
rect 19797 26503 19855 26509
rect 19797 26500 19809 26503
rect 17052 26472 18276 26500
rect 16117 26435 16175 26441
rect 16117 26432 16129 26435
rect 15856 26404 16129 26432
rect 15749 26395 15807 26401
rect 16117 26401 16129 26404
rect 16163 26401 16175 26435
rect 16117 26395 16175 26401
rect 16209 26435 16267 26441
rect 16209 26401 16221 26435
rect 16255 26401 16267 26435
rect 16209 26395 16267 26401
rect 13556 26364 13584 26395
rect 14384 26364 14412 26395
rect 15286 26364 15292 26376
rect 13556 26336 14412 26364
rect 15247 26336 15292 26364
rect 15286 26324 15292 26336
rect 15344 26324 15350 26376
rect 15470 26296 15476 26308
rect 13464 26268 15476 26296
rect 15470 26256 15476 26268
rect 15528 26296 15534 26308
rect 15764 26296 15792 26395
rect 16942 26392 16948 26444
rect 17000 26432 17006 26444
rect 17052 26441 17080 26472
rect 17037 26435 17095 26441
rect 17037 26432 17049 26435
rect 17000 26404 17049 26432
rect 17000 26392 17006 26404
rect 17037 26401 17049 26404
rect 17083 26401 17095 26435
rect 17037 26395 17095 26401
rect 17405 26435 17463 26441
rect 17405 26401 17417 26435
rect 17451 26432 17463 26435
rect 17678 26432 17684 26444
rect 17451 26404 17684 26432
rect 17451 26401 17463 26404
rect 17405 26395 17463 26401
rect 17678 26392 17684 26404
rect 17736 26432 17742 26444
rect 18248 26441 18276 26472
rect 19168 26472 19809 26500
rect 18233 26435 18291 26441
rect 17736 26404 18184 26432
rect 17736 26392 17742 26404
rect 16022 26324 16028 26376
rect 16080 26364 16086 26376
rect 17129 26367 17187 26373
rect 16080 26336 17080 26364
rect 16080 26324 16086 26336
rect 16390 26296 16396 26308
rect 15528 26268 16396 26296
rect 15528 26256 15534 26268
rect 16390 26256 16396 26268
rect 16448 26256 16454 26308
rect 17052 26296 17080 26336
rect 17129 26333 17141 26367
rect 17175 26364 17187 26367
rect 17494 26364 17500 26376
rect 17175 26336 17500 26364
rect 17175 26333 17187 26336
rect 17129 26327 17187 26333
rect 17494 26324 17500 26336
rect 17552 26324 17558 26376
rect 18046 26364 18052 26376
rect 18007 26336 18052 26364
rect 18046 26324 18052 26336
rect 18104 26324 18110 26376
rect 18156 26364 18184 26404
rect 18233 26401 18245 26435
rect 18279 26401 18291 26435
rect 18233 26395 18291 26401
rect 18322 26392 18328 26444
rect 18380 26432 18386 26444
rect 18598 26432 18604 26444
rect 18380 26404 18604 26432
rect 18380 26392 18386 26404
rect 18598 26392 18604 26404
rect 18656 26392 18662 26444
rect 18693 26435 18751 26441
rect 18693 26401 18705 26435
rect 18739 26432 18751 26435
rect 19058 26432 19064 26444
rect 18739 26404 19064 26432
rect 18739 26401 18751 26404
rect 18693 26395 18751 26401
rect 18708 26364 18736 26395
rect 19058 26392 19064 26404
rect 19116 26392 19122 26444
rect 19168 26364 19196 26472
rect 19797 26469 19809 26472
rect 19843 26469 19855 26503
rect 20346 26500 20352 26512
rect 20307 26472 20352 26500
rect 19797 26463 19855 26469
rect 20346 26460 20352 26472
rect 20404 26460 20410 26512
rect 20806 26460 20812 26512
rect 20864 26500 20870 26512
rect 20864 26472 21864 26500
rect 20864 26460 20870 26472
rect 19886 26432 19892 26444
rect 19847 26404 19892 26432
rect 19886 26392 19892 26404
rect 19944 26392 19950 26444
rect 19978 26392 19984 26444
rect 20036 26432 20042 26444
rect 21836 26441 21864 26472
rect 20901 26435 20959 26441
rect 20901 26432 20913 26435
rect 20036 26404 20913 26432
rect 20036 26392 20042 26404
rect 20901 26401 20913 26404
rect 20947 26401 20959 26435
rect 20901 26395 20959 26401
rect 21821 26435 21879 26441
rect 21821 26401 21833 26435
rect 21867 26401 21879 26435
rect 21821 26395 21879 26401
rect 21910 26392 21916 26444
rect 21968 26432 21974 26444
rect 22557 26435 22615 26441
rect 22557 26432 22569 26435
rect 21968 26404 22569 26432
rect 21968 26392 21974 26404
rect 22557 26401 22569 26404
rect 22603 26401 22615 26435
rect 22830 26432 22836 26444
rect 22791 26404 22836 26432
rect 22557 26395 22615 26401
rect 18156 26336 18736 26364
rect 18892 26336 19196 26364
rect 18322 26296 18328 26308
rect 17052 26268 18328 26296
rect 18322 26256 18328 26268
rect 18380 26296 18386 26308
rect 18892 26296 18920 26336
rect 22094 26324 22100 26376
rect 22152 26364 22158 26376
rect 22572 26364 22600 26395
rect 22830 26392 22836 26404
rect 22888 26392 22894 26444
rect 23293 26435 23351 26441
rect 23293 26401 23305 26435
rect 23339 26432 23351 26435
rect 23474 26432 23480 26444
rect 23339 26404 23480 26432
rect 23339 26401 23351 26404
rect 23293 26395 23351 26401
rect 23474 26392 23480 26404
rect 23532 26432 23538 26444
rect 23676 26441 23704 26540
rect 24578 26528 24584 26580
rect 24636 26568 24642 26580
rect 25593 26571 25651 26577
rect 25593 26568 25605 26571
rect 24636 26540 25605 26568
rect 24636 26528 24642 26540
rect 25593 26537 25605 26540
rect 25639 26537 25651 26571
rect 26602 26568 26608 26580
rect 26563 26540 26608 26568
rect 25593 26531 25651 26537
rect 26602 26528 26608 26540
rect 26660 26528 26666 26580
rect 37642 26528 37648 26580
rect 37700 26568 37706 26580
rect 37921 26571 37979 26577
rect 37921 26568 37933 26571
rect 37700 26540 37933 26568
rect 37700 26528 37706 26540
rect 37921 26537 37933 26540
rect 37967 26537 37979 26571
rect 37921 26531 37979 26537
rect 30834 26460 30840 26512
rect 30892 26500 30898 26512
rect 30892 26472 32352 26500
rect 30892 26460 30898 26472
rect 23661 26435 23719 26441
rect 23532 26404 23612 26432
rect 23532 26392 23538 26404
rect 23584 26364 23612 26404
rect 23661 26401 23673 26435
rect 23707 26401 23719 26435
rect 24210 26432 24216 26444
rect 24171 26404 24216 26432
rect 23661 26395 23719 26401
rect 24210 26392 24216 26404
rect 24268 26392 24274 26444
rect 24946 26392 24952 26444
rect 25004 26432 25010 26444
rect 25409 26435 25467 26441
rect 25409 26432 25421 26435
rect 25004 26404 25421 26432
rect 25004 26392 25010 26404
rect 25409 26401 25421 26404
rect 25455 26401 25467 26435
rect 26510 26432 26516 26444
rect 26471 26404 26516 26432
rect 25409 26395 25467 26401
rect 26510 26392 26516 26404
rect 26568 26392 26574 26444
rect 27065 26435 27123 26441
rect 27065 26401 27077 26435
rect 27111 26432 27123 26435
rect 30101 26435 30159 26441
rect 27111 26404 28028 26432
rect 27111 26401 27123 26404
rect 27065 26395 27123 26401
rect 28000 26376 28028 26404
rect 30101 26401 30113 26435
rect 30147 26432 30159 26435
rect 30558 26432 30564 26444
rect 30147 26404 30564 26432
rect 30147 26401 30159 26404
rect 30101 26395 30159 26401
rect 30558 26392 30564 26404
rect 30616 26392 30622 26444
rect 30653 26435 30711 26441
rect 30653 26401 30665 26435
rect 30699 26432 30711 26435
rect 32122 26432 32128 26444
rect 30699 26404 32128 26432
rect 30699 26401 30711 26404
rect 30653 26395 30711 26401
rect 32122 26392 32128 26404
rect 32180 26392 32186 26444
rect 32324 26441 32352 26472
rect 32309 26435 32367 26441
rect 32309 26401 32321 26435
rect 32355 26432 32367 26435
rect 33318 26432 33324 26444
rect 32355 26404 33324 26432
rect 32355 26401 32367 26404
rect 32309 26395 32367 26401
rect 33318 26392 33324 26404
rect 33376 26392 33382 26444
rect 33502 26432 33508 26444
rect 33463 26404 33508 26432
rect 33502 26392 33508 26404
rect 33560 26392 33566 26444
rect 35526 26432 35532 26444
rect 35487 26404 35532 26432
rect 35526 26392 35532 26404
rect 35584 26392 35590 26444
rect 35802 26432 35808 26444
rect 35763 26404 35808 26432
rect 35802 26392 35808 26404
rect 35860 26392 35866 26444
rect 38010 26432 38016 26444
rect 37971 26404 38016 26432
rect 38010 26392 38016 26404
rect 38068 26392 38074 26444
rect 38381 26435 38439 26441
rect 38381 26401 38393 26435
rect 38427 26432 38439 26435
rect 39022 26432 39028 26444
rect 38427 26404 39028 26432
rect 38427 26401 38439 26404
rect 38381 26395 38439 26401
rect 39022 26392 39028 26404
rect 39080 26392 39086 26444
rect 24118 26364 24124 26376
rect 22152 26336 22197 26364
rect 22572 26336 23520 26364
rect 23584 26336 24124 26364
rect 22152 26324 22158 26336
rect 20070 26296 20076 26308
rect 18380 26268 18920 26296
rect 18984 26268 20076 26296
rect 18380 26256 18386 26268
rect 7834 26228 7840 26240
rect 6880 26200 7840 26228
rect 6880 26188 6886 26200
rect 7834 26188 7840 26200
rect 7892 26228 7898 26240
rect 11422 26228 11428 26240
rect 7892 26200 11428 26228
rect 7892 26188 7898 26200
rect 11422 26188 11428 26200
rect 11480 26188 11486 26240
rect 18598 26188 18604 26240
rect 18656 26228 18662 26240
rect 18984 26228 19012 26268
rect 20070 26256 20076 26268
rect 20128 26256 20134 26308
rect 23492 26240 23520 26336
rect 24118 26324 24124 26336
rect 24176 26364 24182 26376
rect 24394 26364 24400 26376
rect 24176 26336 24400 26364
rect 24176 26324 24182 26336
rect 24394 26324 24400 26336
rect 24452 26364 24458 26376
rect 24581 26367 24639 26373
rect 24581 26364 24593 26367
rect 24452 26336 24593 26364
rect 24452 26324 24458 26336
rect 24581 26333 24593 26336
rect 24627 26333 24639 26367
rect 24581 26327 24639 26333
rect 27801 26367 27859 26373
rect 27801 26333 27813 26367
rect 27847 26333 27859 26367
rect 27801 26327 27859 26333
rect 23566 26256 23572 26308
rect 23624 26296 23630 26308
rect 24489 26299 24547 26305
rect 24489 26296 24501 26299
rect 23624 26268 24501 26296
rect 23624 26256 23630 26268
rect 24489 26265 24501 26268
rect 24535 26265 24547 26299
rect 27706 26296 27712 26308
rect 24489 26259 24547 26265
rect 27540 26268 27712 26296
rect 18656 26200 19012 26228
rect 18656 26188 18662 26200
rect 19426 26188 19432 26240
rect 19484 26228 19490 26240
rect 19613 26231 19671 26237
rect 19613 26228 19625 26231
rect 19484 26200 19625 26228
rect 19484 26188 19490 26200
rect 19613 26197 19625 26200
rect 19659 26197 19671 26231
rect 19613 26191 19671 26197
rect 23474 26188 23480 26240
rect 23532 26228 23538 26240
rect 23842 26228 23848 26240
rect 23532 26200 23848 26228
rect 23532 26188 23538 26200
rect 23842 26188 23848 26200
rect 23900 26228 23906 26240
rect 24351 26231 24409 26237
rect 24351 26228 24363 26231
rect 23900 26200 24363 26228
rect 23900 26188 23906 26200
rect 24351 26197 24363 26200
rect 24397 26197 24409 26231
rect 24854 26228 24860 26240
rect 24815 26200 24860 26228
rect 24351 26191 24409 26197
rect 24854 26188 24860 26200
rect 24912 26188 24918 26240
rect 26142 26188 26148 26240
rect 26200 26228 26206 26240
rect 27540 26228 27568 26268
rect 27706 26256 27712 26268
rect 27764 26296 27770 26308
rect 27816 26296 27844 26327
rect 27982 26324 27988 26376
rect 28040 26324 28046 26376
rect 28077 26367 28135 26373
rect 28077 26333 28089 26367
rect 28123 26364 28135 26367
rect 29270 26364 29276 26376
rect 28123 26336 29276 26364
rect 28123 26333 28135 26336
rect 28077 26327 28135 26333
rect 29270 26324 29276 26336
rect 29328 26324 29334 26376
rect 30745 26367 30803 26373
rect 30745 26364 30757 26367
rect 30116 26336 30757 26364
rect 30116 26308 30144 26336
rect 30745 26333 30757 26336
rect 30791 26333 30803 26367
rect 31570 26364 31576 26376
rect 30745 26327 30803 26333
rect 31220 26336 31576 26364
rect 27764 26268 27844 26296
rect 27764 26256 27770 26268
rect 29638 26256 29644 26308
rect 29696 26296 29702 26308
rect 30009 26299 30067 26305
rect 30009 26296 30021 26299
rect 29696 26268 30021 26296
rect 29696 26256 29702 26268
rect 30009 26265 30021 26268
rect 30055 26265 30067 26299
rect 30009 26259 30067 26265
rect 30098 26256 30104 26308
rect 30156 26256 30162 26308
rect 29178 26228 29184 26240
rect 26200 26200 27568 26228
rect 29139 26200 29184 26228
rect 26200 26188 26206 26200
rect 29178 26188 29184 26200
rect 29236 26188 29242 26240
rect 29730 26188 29736 26240
rect 29788 26228 29794 26240
rect 31220 26228 31248 26336
rect 31570 26324 31576 26336
rect 31628 26364 31634 26376
rect 33229 26367 33287 26373
rect 33229 26364 33241 26367
rect 31628 26336 33241 26364
rect 31628 26324 31634 26336
rect 33229 26333 33241 26336
rect 33275 26364 33287 26367
rect 35544 26364 35572 26392
rect 33275 26336 35572 26364
rect 33275 26333 33287 26336
rect 33229 26327 33287 26333
rect 31662 26256 31668 26308
rect 31720 26296 31726 26308
rect 32493 26299 32551 26305
rect 32493 26296 32505 26299
rect 31720 26268 32505 26296
rect 31720 26256 31726 26268
rect 32493 26265 32505 26268
rect 32539 26265 32551 26299
rect 32493 26259 32551 26265
rect 34606 26228 34612 26240
rect 29788 26200 31248 26228
rect 34567 26200 34612 26228
rect 29788 26188 29794 26200
rect 34606 26188 34612 26200
rect 34664 26188 34670 26240
rect 36538 26188 36544 26240
rect 36596 26228 36602 26240
rect 36722 26228 36728 26240
rect 36596 26200 36728 26228
rect 36596 26188 36602 26200
rect 36722 26188 36728 26200
rect 36780 26228 36786 26240
rect 36909 26231 36967 26237
rect 36909 26228 36921 26231
rect 36780 26200 36921 26228
rect 36780 26188 36786 26200
rect 36909 26197 36921 26200
rect 36955 26197 36967 26231
rect 36909 26191 36967 26197
rect 1104 26138 39836 26160
rect 1104 26086 4246 26138
rect 4298 26086 4310 26138
rect 4362 26086 4374 26138
rect 4426 26086 4438 26138
rect 4490 26086 34966 26138
rect 35018 26086 35030 26138
rect 35082 26086 35094 26138
rect 35146 26086 35158 26138
rect 35210 26086 39836 26138
rect 1104 26064 39836 26086
rect 4157 26027 4215 26033
rect 4157 25993 4169 26027
rect 4203 26024 4215 26027
rect 4614 26024 4620 26036
rect 4203 25996 4620 26024
rect 4203 25993 4215 25996
rect 4157 25987 4215 25993
rect 4614 25984 4620 25996
rect 4672 25984 4678 26036
rect 22462 26024 22468 26036
rect 14660 25996 22468 26024
rect 10962 25956 10968 25968
rect 8956 25928 10968 25956
rect 2774 25888 2780 25900
rect 2700 25860 2780 25888
rect 2593 25823 2651 25829
rect 2593 25789 2605 25823
rect 2639 25820 2651 25823
rect 2700 25820 2728 25860
rect 2774 25848 2780 25860
rect 2832 25848 2838 25900
rect 8956 25888 8984 25928
rect 10962 25916 10968 25928
rect 11020 25916 11026 25968
rect 11054 25916 11060 25968
rect 11112 25956 11118 25968
rect 11238 25956 11244 25968
rect 11112 25928 11244 25956
rect 11112 25916 11118 25928
rect 11238 25916 11244 25928
rect 11296 25956 11302 25968
rect 14660 25965 14688 25996
rect 22462 25984 22468 25996
rect 22520 25984 22526 26036
rect 25498 25984 25504 26036
rect 25556 26024 25562 26036
rect 25593 26027 25651 26033
rect 25593 26024 25605 26027
rect 25556 25996 25605 26024
rect 25556 25984 25562 25996
rect 25593 25993 25605 25996
rect 25639 26024 25651 26027
rect 25774 26024 25780 26036
rect 25639 25996 25780 26024
rect 25639 25993 25651 25996
rect 25593 25987 25651 25993
rect 25774 25984 25780 25996
rect 25832 25984 25838 26036
rect 32122 25984 32128 26036
rect 32180 26024 32186 26036
rect 33229 26027 33287 26033
rect 33229 26024 33241 26027
rect 32180 25996 33241 26024
rect 32180 25984 32186 25996
rect 33229 25993 33241 25996
rect 33275 25993 33287 26027
rect 33229 25987 33287 25993
rect 35618 25984 35624 26036
rect 35676 26024 35682 26036
rect 36265 26027 36323 26033
rect 36265 26024 36277 26027
rect 35676 25996 36277 26024
rect 35676 25984 35682 25996
rect 36265 25993 36277 25996
rect 36311 25993 36323 26027
rect 36265 25987 36323 25993
rect 39025 26027 39083 26033
rect 39025 25993 39037 26027
rect 39071 26024 39083 26027
rect 39114 26024 39120 26036
rect 39071 25996 39120 26024
rect 39071 25993 39083 25996
rect 39025 25987 39083 25993
rect 39114 25984 39120 25996
rect 39172 25984 39178 26036
rect 11793 25959 11851 25965
rect 11793 25956 11805 25959
rect 11296 25928 11805 25956
rect 11296 25916 11302 25928
rect 11793 25925 11805 25928
rect 11839 25925 11851 25959
rect 11793 25919 11851 25925
rect 14645 25959 14703 25965
rect 14645 25925 14657 25959
rect 14691 25925 14703 25959
rect 14645 25919 14703 25925
rect 15565 25959 15623 25965
rect 15565 25925 15577 25959
rect 15611 25956 15623 25959
rect 23937 25959 23995 25965
rect 15611 25928 22416 25956
rect 15611 25925 15623 25928
rect 15565 25919 15623 25925
rect 11974 25888 11980 25900
rect 8772 25860 8984 25888
rect 10704 25860 11980 25888
rect 2639 25792 2728 25820
rect 2869 25823 2927 25829
rect 2639 25789 2651 25792
rect 2593 25783 2651 25789
rect 2869 25789 2881 25823
rect 2915 25820 2927 25823
rect 4154 25820 4160 25832
rect 2915 25792 4160 25820
rect 2915 25789 2927 25792
rect 2869 25783 2927 25789
rect 4154 25780 4160 25792
rect 4212 25780 4218 25832
rect 4614 25780 4620 25832
rect 4672 25820 4678 25832
rect 4709 25823 4767 25829
rect 4709 25820 4721 25823
rect 4672 25792 4721 25820
rect 4672 25780 4678 25792
rect 4709 25789 4721 25792
rect 4755 25789 4767 25823
rect 5718 25820 5724 25832
rect 5679 25792 5724 25820
rect 4709 25783 4767 25789
rect 5718 25780 5724 25792
rect 5776 25780 5782 25832
rect 7098 25820 7104 25832
rect 7059 25792 7104 25820
rect 7098 25780 7104 25792
rect 7156 25780 7162 25832
rect 8113 25823 8171 25829
rect 8113 25789 8125 25823
rect 8159 25820 8171 25823
rect 8202 25820 8208 25832
rect 8159 25792 8208 25820
rect 8159 25789 8171 25792
rect 8113 25783 8171 25789
rect 8202 25780 8208 25792
rect 8260 25780 8266 25832
rect 8662 25820 8668 25832
rect 8575 25792 8668 25820
rect 8662 25780 8668 25792
rect 8720 25820 8726 25832
rect 8772 25820 8800 25860
rect 8720 25792 8800 25820
rect 8849 25823 8907 25829
rect 8720 25780 8726 25792
rect 8849 25789 8861 25823
rect 8895 25789 8907 25823
rect 9398 25820 9404 25832
rect 9359 25792 9404 25820
rect 8849 25783 8907 25789
rect 7466 25712 7472 25764
rect 7524 25752 7530 25764
rect 7524 25724 8248 25752
rect 7524 25712 7530 25724
rect 4062 25644 4068 25696
rect 4120 25684 4126 25696
rect 4893 25687 4951 25693
rect 4893 25684 4905 25687
rect 4120 25656 4905 25684
rect 4120 25644 4126 25656
rect 4893 25653 4905 25656
rect 4939 25653 4951 25687
rect 4893 25647 4951 25653
rect 5810 25644 5816 25696
rect 5868 25684 5874 25696
rect 5905 25687 5963 25693
rect 5905 25684 5917 25687
rect 5868 25656 5917 25684
rect 5868 25644 5874 25656
rect 5905 25653 5917 25656
rect 5951 25653 5963 25687
rect 5905 25647 5963 25653
rect 7285 25687 7343 25693
rect 7285 25653 7297 25687
rect 7331 25684 7343 25687
rect 7650 25684 7656 25696
rect 7331 25656 7656 25684
rect 7331 25653 7343 25656
rect 7285 25647 7343 25653
rect 7650 25644 7656 25656
rect 7708 25644 7714 25696
rect 8018 25644 8024 25696
rect 8076 25684 8082 25696
rect 8113 25687 8171 25693
rect 8113 25684 8125 25687
rect 8076 25656 8125 25684
rect 8076 25644 8082 25656
rect 8113 25653 8125 25656
rect 8159 25653 8171 25687
rect 8220 25684 8248 25724
rect 8570 25712 8576 25764
rect 8628 25752 8634 25764
rect 8864 25752 8892 25783
rect 9398 25780 9404 25792
rect 9456 25780 9462 25832
rect 10704 25829 10732 25860
rect 11974 25848 11980 25860
rect 12032 25848 12038 25900
rect 12437 25891 12495 25897
rect 12437 25857 12449 25891
rect 12483 25888 12495 25891
rect 13078 25888 13084 25900
rect 12483 25860 13084 25888
rect 12483 25857 12495 25860
rect 12437 25851 12495 25857
rect 13078 25848 13084 25860
rect 13136 25848 13142 25900
rect 19334 25888 19340 25900
rect 18616 25860 19340 25888
rect 10689 25823 10747 25829
rect 10689 25789 10701 25823
rect 10735 25789 10747 25823
rect 10870 25820 10876 25832
rect 10831 25792 10876 25820
rect 10689 25783 10747 25789
rect 10870 25780 10876 25792
rect 10928 25780 10934 25832
rect 11241 25823 11299 25829
rect 11241 25789 11253 25823
rect 11287 25789 11299 25823
rect 11609 25823 11667 25829
rect 11609 25820 11621 25823
rect 11241 25783 11299 25789
rect 11348 25792 11621 25820
rect 11256 25752 11284 25783
rect 8628 25724 11284 25752
rect 8628 25712 8634 25724
rect 9493 25687 9551 25693
rect 9493 25684 9505 25687
rect 8220 25656 9505 25684
rect 8113 25647 8171 25653
rect 9493 25653 9505 25656
rect 9539 25653 9551 25687
rect 9493 25647 9551 25653
rect 10962 25644 10968 25696
rect 11020 25684 11026 25696
rect 11348 25684 11376 25792
rect 11609 25789 11621 25792
rect 11655 25789 11667 25823
rect 11609 25783 11667 25789
rect 12526 25780 12532 25832
rect 12584 25820 12590 25832
rect 12713 25823 12771 25829
rect 12713 25820 12725 25823
rect 12584 25792 12725 25820
rect 12584 25780 12590 25792
rect 12713 25789 12725 25792
rect 12759 25789 12771 25823
rect 13814 25820 13820 25832
rect 13775 25792 13820 25820
rect 12713 25783 12771 25789
rect 13814 25780 13820 25792
rect 13872 25780 13878 25832
rect 14274 25820 14280 25832
rect 14235 25792 14280 25820
rect 14274 25780 14280 25792
rect 14332 25780 14338 25832
rect 14550 25820 14556 25832
rect 14511 25792 14556 25820
rect 14550 25780 14556 25792
rect 14608 25780 14614 25832
rect 15286 25820 15292 25832
rect 15247 25792 15292 25820
rect 15286 25780 15292 25792
rect 15344 25780 15350 25832
rect 15746 25780 15752 25832
rect 15804 25820 15810 25832
rect 15841 25823 15899 25829
rect 15841 25820 15853 25823
rect 15804 25792 15853 25820
rect 15804 25780 15810 25792
rect 15841 25789 15853 25792
rect 15887 25789 15899 25823
rect 16114 25820 16120 25832
rect 16075 25792 16120 25820
rect 15841 25783 15899 25789
rect 16114 25780 16120 25792
rect 16172 25780 16178 25832
rect 16942 25820 16948 25832
rect 16903 25792 16948 25820
rect 16942 25780 16948 25792
rect 17000 25780 17006 25832
rect 17129 25823 17187 25829
rect 17129 25789 17141 25823
rect 17175 25820 17187 25823
rect 17678 25820 17684 25832
rect 17175 25792 17684 25820
rect 17175 25789 17187 25792
rect 17129 25783 17187 25789
rect 17678 25780 17684 25792
rect 17736 25780 17742 25832
rect 18616 25829 18644 25860
rect 19334 25848 19340 25860
rect 19392 25888 19398 25900
rect 19978 25888 19984 25900
rect 19392 25860 19984 25888
rect 19392 25848 19398 25860
rect 19978 25848 19984 25860
rect 20036 25848 20042 25900
rect 21358 25888 21364 25900
rect 21319 25860 21364 25888
rect 21358 25848 21364 25860
rect 21416 25848 21422 25900
rect 22094 25848 22100 25900
rect 22152 25888 22158 25900
rect 22152 25860 22197 25888
rect 22152 25848 22158 25860
rect 18601 25823 18659 25829
rect 18601 25789 18613 25823
rect 18647 25789 18659 25823
rect 18601 25783 18659 25789
rect 18690 25780 18696 25832
rect 18748 25820 18754 25832
rect 19150 25820 19156 25832
rect 18748 25792 18793 25820
rect 19111 25792 19156 25820
rect 18748 25780 18754 25792
rect 19150 25780 19156 25792
rect 19208 25820 19214 25832
rect 19610 25820 19616 25832
rect 19208 25792 19616 25820
rect 19208 25780 19214 25792
rect 19610 25780 19616 25792
rect 19668 25780 19674 25832
rect 19797 25823 19855 25829
rect 19797 25789 19809 25823
rect 19843 25820 19855 25823
rect 19886 25820 19892 25832
rect 19843 25792 19892 25820
rect 19843 25789 19855 25792
rect 19797 25783 19855 25789
rect 19886 25780 19892 25792
rect 19944 25780 19950 25832
rect 20438 25820 20444 25832
rect 20399 25792 20444 25820
rect 20438 25780 20444 25792
rect 20496 25780 20502 25832
rect 20625 25823 20683 25829
rect 20625 25789 20637 25823
rect 20671 25789 20683 25823
rect 21174 25820 21180 25832
rect 21135 25792 21180 25820
rect 20625 25783 20683 25789
rect 11422 25712 11428 25764
rect 11480 25752 11486 25764
rect 12621 25755 12679 25761
rect 12621 25752 12633 25755
rect 11480 25724 12633 25752
rect 11480 25712 11486 25724
rect 12621 25721 12633 25724
rect 12667 25721 12679 25755
rect 13170 25752 13176 25764
rect 13131 25724 13176 25752
rect 12621 25715 12679 25721
rect 13170 25712 13176 25724
rect 13228 25712 13234 25764
rect 17497 25755 17555 25761
rect 17497 25721 17509 25755
rect 17543 25752 17555 25755
rect 18046 25752 18052 25764
rect 17543 25724 18052 25752
rect 17543 25721 17555 25724
rect 17497 25715 17555 25721
rect 18046 25712 18052 25724
rect 18104 25712 18110 25764
rect 19521 25755 19579 25761
rect 19521 25721 19533 25755
rect 19567 25752 19579 25755
rect 19702 25752 19708 25764
rect 19567 25724 19708 25752
rect 19567 25721 19579 25724
rect 19521 25715 19579 25721
rect 19702 25712 19708 25724
rect 19760 25712 19766 25764
rect 19978 25712 19984 25764
rect 20036 25752 20042 25764
rect 20640 25752 20668 25783
rect 21174 25780 21180 25792
rect 21232 25780 21238 25832
rect 22388 25829 22416 25928
rect 23937 25925 23949 25959
rect 23983 25925 23995 25959
rect 31846 25956 31852 25968
rect 31807 25928 31852 25956
rect 23937 25919 23995 25925
rect 23952 25888 23980 25919
rect 31846 25916 31852 25928
rect 31904 25916 31910 25968
rect 24670 25888 24676 25900
rect 22940 25860 23980 25888
rect 24631 25860 24676 25888
rect 22940 25829 22968 25860
rect 24670 25848 24676 25860
rect 24728 25848 24734 25900
rect 25222 25848 25228 25900
rect 25280 25888 25286 25900
rect 26142 25888 26148 25900
rect 25280 25860 26148 25888
rect 25280 25848 25286 25860
rect 26142 25848 26148 25860
rect 26200 25888 26206 25900
rect 26421 25891 26479 25897
rect 26421 25888 26433 25891
rect 26200 25860 26433 25888
rect 26200 25848 26206 25860
rect 26421 25857 26433 25860
rect 26467 25857 26479 25891
rect 29638 25888 29644 25900
rect 29599 25860 29644 25888
rect 26421 25851 26479 25857
rect 29638 25848 29644 25860
rect 29696 25848 29702 25900
rect 32306 25888 32312 25900
rect 31680 25860 32312 25888
rect 22373 25823 22431 25829
rect 22373 25789 22385 25823
rect 22419 25789 22431 25823
rect 22373 25783 22431 25789
rect 22925 25823 22983 25829
rect 22925 25789 22937 25823
rect 22971 25789 22983 25823
rect 23658 25820 23664 25832
rect 23619 25792 23664 25820
rect 22925 25783 22983 25789
rect 23658 25780 23664 25792
rect 23716 25780 23722 25832
rect 24578 25820 24584 25832
rect 24539 25792 24584 25820
rect 24578 25780 24584 25792
rect 24636 25780 24642 25832
rect 25314 25780 25320 25832
rect 25372 25820 25378 25832
rect 25409 25823 25467 25829
rect 25409 25820 25421 25823
rect 25372 25792 25421 25820
rect 25372 25780 25378 25792
rect 25409 25789 25421 25792
rect 25455 25789 25467 25823
rect 26694 25820 26700 25832
rect 26655 25792 26700 25820
rect 25409 25783 25467 25789
rect 26694 25780 26700 25792
rect 26752 25780 26758 25832
rect 28537 25823 28595 25829
rect 28537 25789 28549 25823
rect 28583 25820 28595 25823
rect 29178 25820 29184 25832
rect 28583 25792 29184 25820
rect 28583 25789 28595 25792
rect 28537 25783 28595 25789
rect 29178 25780 29184 25792
rect 29236 25780 29242 25832
rect 31680 25829 31708 25860
rect 32306 25848 32312 25860
rect 32364 25848 32370 25900
rect 34885 25891 34943 25897
rect 34885 25857 34897 25891
rect 34931 25888 34943 25891
rect 35526 25888 35532 25900
rect 34931 25860 35532 25888
rect 34931 25857 34943 25860
rect 34885 25851 34943 25857
rect 35526 25848 35532 25860
rect 35584 25848 35590 25900
rect 37458 25888 37464 25900
rect 37419 25860 37464 25888
rect 37458 25848 37464 25860
rect 37516 25848 37522 25900
rect 37737 25891 37795 25897
rect 37737 25857 37749 25891
rect 37783 25888 37795 25891
rect 37826 25888 37832 25900
rect 37783 25860 37832 25888
rect 37783 25857 37795 25860
rect 37737 25851 37795 25857
rect 37826 25848 37832 25860
rect 37884 25848 37890 25900
rect 29365 25823 29423 25829
rect 29365 25789 29377 25823
rect 29411 25789 29423 25823
rect 29365 25783 29423 25789
rect 31665 25823 31723 25829
rect 31665 25789 31677 25823
rect 31711 25789 31723 25823
rect 32214 25820 32220 25832
rect 32175 25792 32220 25820
rect 31665 25783 31723 25789
rect 20036 25724 20668 25752
rect 23109 25755 23167 25761
rect 20036 25712 20042 25724
rect 23109 25721 23121 25755
rect 23155 25752 23167 25755
rect 25130 25752 25136 25764
rect 23155 25724 25136 25752
rect 23155 25721 23167 25724
rect 23109 25715 23167 25721
rect 25130 25712 25136 25724
rect 25188 25712 25194 25764
rect 28074 25752 28080 25764
rect 28035 25724 28080 25752
rect 28074 25712 28080 25724
rect 28132 25712 28138 25764
rect 11020 25656 11376 25684
rect 11020 25644 11026 25656
rect 13722 25644 13728 25696
rect 13780 25684 13786 25696
rect 22554 25684 22560 25696
rect 13780 25656 22560 25684
rect 13780 25644 13786 25656
rect 22554 25644 22560 25656
rect 22612 25644 22618 25696
rect 28626 25684 28632 25696
rect 28587 25656 28632 25684
rect 28626 25644 28632 25656
rect 28684 25644 28690 25696
rect 29380 25684 29408 25783
rect 32214 25780 32220 25792
rect 32272 25780 32278 25832
rect 32490 25820 32496 25832
rect 32451 25792 32496 25820
rect 32490 25780 32496 25792
rect 32548 25780 32554 25832
rect 33137 25823 33195 25829
rect 33137 25789 33149 25823
rect 33183 25789 33195 25823
rect 33137 25783 33195 25789
rect 33873 25823 33931 25829
rect 33873 25789 33885 25823
rect 33919 25820 33931 25823
rect 34054 25820 34060 25832
rect 33919 25792 34060 25820
rect 33919 25789 33931 25792
rect 33873 25783 33931 25789
rect 30374 25712 30380 25764
rect 30432 25752 30438 25764
rect 31021 25755 31079 25761
rect 31021 25752 31033 25755
rect 30432 25724 31033 25752
rect 30432 25712 30438 25724
rect 31021 25721 31033 25724
rect 31067 25752 31079 25755
rect 33152 25752 33180 25783
rect 34054 25780 34060 25792
rect 34112 25780 34118 25832
rect 35158 25820 35164 25832
rect 35119 25792 35164 25820
rect 35158 25780 35164 25792
rect 35216 25780 35222 25832
rect 31067 25724 33180 25752
rect 31067 25721 31079 25724
rect 31021 25715 31079 25721
rect 29638 25684 29644 25696
rect 29380 25656 29644 25684
rect 29638 25644 29644 25656
rect 29696 25644 29702 25696
rect 1104 25594 39836 25616
rect 1104 25542 19606 25594
rect 19658 25542 19670 25594
rect 19722 25542 19734 25594
rect 19786 25542 19798 25594
rect 19850 25542 39836 25594
rect 1104 25520 39836 25542
rect 2866 25440 2872 25492
rect 2924 25480 2930 25492
rect 2961 25483 3019 25489
rect 2961 25480 2973 25483
rect 2924 25452 2973 25480
rect 2924 25440 2930 25452
rect 2961 25449 2973 25452
rect 3007 25449 3019 25483
rect 4154 25480 4160 25492
rect 4115 25452 4160 25480
rect 2961 25443 3019 25449
rect 4154 25440 4160 25452
rect 4212 25440 4218 25492
rect 7006 25480 7012 25492
rect 5644 25452 7012 25480
rect 4062 25412 4068 25424
rect 2976 25384 4068 25412
rect 2976 25356 3004 25384
rect 4062 25372 4068 25384
rect 4120 25412 4126 25424
rect 4120 25384 4568 25412
rect 4120 25372 4126 25384
rect 1397 25347 1455 25353
rect 1397 25313 1409 25347
rect 1443 25344 1455 25347
rect 2774 25344 2780 25356
rect 1443 25316 2780 25344
rect 1443 25313 1455 25316
rect 1397 25307 1455 25313
rect 2774 25304 2780 25316
rect 2832 25304 2838 25356
rect 2958 25304 2964 25356
rect 3016 25304 3022 25356
rect 4540 25353 4568 25384
rect 5644 25353 5672 25452
rect 7006 25440 7012 25452
rect 7064 25480 7070 25492
rect 15381 25483 15439 25489
rect 7064 25452 7788 25480
rect 7064 25440 7070 25452
rect 7760 25421 7788 25452
rect 15381 25449 15393 25483
rect 15427 25480 15439 25483
rect 16114 25480 16120 25492
rect 15427 25452 16120 25480
rect 15427 25449 15439 25452
rect 15381 25443 15439 25449
rect 16114 25440 16120 25452
rect 16172 25440 16178 25492
rect 18693 25483 18751 25489
rect 18693 25449 18705 25483
rect 18739 25480 18751 25483
rect 19334 25480 19340 25492
rect 18739 25452 19340 25480
rect 18739 25449 18751 25452
rect 18693 25443 18751 25449
rect 19334 25440 19340 25452
rect 19392 25440 19398 25492
rect 19426 25440 19432 25492
rect 19484 25480 19490 25492
rect 19521 25483 19579 25489
rect 19521 25480 19533 25483
rect 19484 25452 19533 25480
rect 19484 25440 19490 25452
rect 19521 25449 19533 25452
rect 19567 25449 19579 25483
rect 23474 25480 23480 25492
rect 23435 25452 23480 25480
rect 19521 25443 19579 25449
rect 23474 25440 23480 25452
rect 23532 25440 23538 25492
rect 26605 25483 26663 25489
rect 26605 25449 26617 25483
rect 26651 25480 26663 25483
rect 26694 25480 26700 25492
rect 26651 25452 26700 25480
rect 26651 25449 26663 25452
rect 26605 25443 26663 25449
rect 26694 25440 26700 25452
rect 26752 25440 26758 25492
rect 28074 25440 28080 25492
rect 28132 25480 28138 25492
rect 33505 25483 33563 25489
rect 28132 25452 32720 25480
rect 28132 25440 28138 25452
rect 7745 25415 7803 25421
rect 7745 25381 7757 25415
rect 7791 25381 7803 25415
rect 8110 25412 8116 25424
rect 8071 25384 8116 25412
rect 7745 25375 7803 25381
rect 8110 25372 8116 25384
rect 8168 25372 8174 25424
rect 11146 25372 11152 25424
rect 11204 25412 11210 25424
rect 11514 25412 11520 25424
rect 11204 25384 11520 25412
rect 11204 25372 11210 25384
rect 11514 25372 11520 25384
rect 11572 25372 11578 25424
rect 11974 25372 11980 25424
rect 12032 25412 12038 25424
rect 19242 25412 19248 25424
rect 12032 25384 16160 25412
rect 19203 25384 19248 25412
rect 12032 25372 12038 25384
rect 4341 25347 4399 25353
rect 4341 25313 4353 25347
rect 4387 25313 4399 25347
rect 4341 25307 4399 25313
rect 4525 25347 4583 25353
rect 4525 25313 4537 25347
rect 4571 25313 4583 25347
rect 4525 25307 4583 25313
rect 5629 25347 5687 25353
rect 5629 25313 5641 25347
rect 5675 25313 5687 25347
rect 5810 25344 5816 25356
rect 5771 25316 5816 25344
rect 5629 25307 5687 25313
rect 1670 25276 1676 25288
rect 1631 25248 1676 25276
rect 1670 25236 1676 25248
rect 1728 25236 1734 25288
rect 4356 25276 4384 25307
rect 5810 25304 5816 25316
rect 5868 25304 5874 25356
rect 6086 25304 6092 25356
rect 6144 25344 6150 25356
rect 6822 25344 6828 25356
rect 6144 25316 6189 25344
rect 6783 25316 6828 25344
rect 6144 25304 6150 25316
rect 6822 25304 6828 25316
rect 6880 25304 6886 25356
rect 7558 25344 7564 25356
rect 7519 25316 7564 25344
rect 7558 25304 7564 25316
rect 7616 25304 7622 25356
rect 7653 25347 7711 25353
rect 7653 25313 7665 25347
rect 7699 25344 7711 25347
rect 8570 25344 8576 25356
rect 7699 25316 8340 25344
rect 8531 25316 8576 25344
rect 7699 25313 7711 25316
rect 7653 25307 7711 25313
rect 5074 25276 5080 25288
rect 4356 25248 5080 25276
rect 5074 25236 5080 25248
rect 5132 25236 5138 25288
rect 5534 25276 5540 25288
rect 5495 25248 5540 25276
rect 5534 25236 5540 25248
rect 5592 25236 5598 25288
rect 7098 25236 7104 25288
rect 7156 25276 7162 25288
rect 7377 25279 7435 25285
rect 7377 25276 7389 25279
rect 7156 25248 7389 25276
rect 7156 25236 7162 25248
rect 7377 25245 7389 25248
rect 7423 25276 7435 25279
rect 7742 25276 7748 25288
rect 7423 25248 7748 25276
rect 7423 25245 7435 25248
rect 7377 25239 7435 25245
rect 7742 25236 7748 25248
rect 7800 25236 7806 25288
rect 8312 25276 8340 25316
rect 8570 25304 8576 25316
rect 8628 25304 8634 25356
rect 9861 25347 9919 25353
rect 9861 25313 9873 25347
rect 9907 25344 9919 25347
rect 11054 25344 11060 25356
rect 9907 25316 11060 25344
rect 9907 25313 9919 25316
rect 9861 25307 9919 25313
rect 11054 25304 11060 25316
rect 11112 25304 11118 25356
rect 12802 25344 12808 25356
rect 12763 25316 12808 25344
rect 12802 25304 12808 25316
rect 12860 25304 12866 25356
rect 13262 25344 13268 25356
rect 13223 25316 13268 25344
rect 13262 25304 13268 25316
rect 13320 25304 13326 25356
rect 13541 25347 13599 25353
rect 13541 25313 13553 25347
rect 13587 25344 13599 25347
rect 13722 25344 13728 25356
rect 13587 25316 13728 25344
rect 13587 25313 13599 25316
rect 13541 25307 13599 25313
rect 13722 25304 13728 25316
rect 13780 25304 13786 25356
rect 14550 25344 14556 25356
rect 14511 25316 14556 25344
rect 14550 25304 14556 25316
rect 14608 25304 14614 25356
rect 15378 25344 15384 25356
rect 15339 25316 15384 25344
rect 15378 25304 15384 25316
rect 15436 25304 15442 25356
rect 15470 25304 15476 25356
rect 15528 25344 15534 25356
rect 16132 25353 16160 25384
rect 19242 25372 19248 25384
rect 19300 25372 19306 25424
rect 20070 25372 20076 25424
rect 20128 25412 20134 25424
rect 26510 25412 26516 25424
rect 20128 25384 22600 25412
rect 20128 25372 20134 25384
rect 15841 25347 15899 25353
rect 15841 25344 15853 25347
rect 15528 25316 15853 25344
rect 15528 25304 15534 25316
rect 15841 25313 15853 25316
rect 15887 25313 15899 25347
rect 15841 25307 15899 25313
rect 16117 25347 16175 25353
rect 16117 25313 16129 25347
rect 16163 25313 16175 25347
rect 16117 25307 16175 25313
rect 17129 25347 17187 25353
rect 17129 25313 17141 25347
rect 17175 25344 17187 25347
rect 18230 25344 18236 25356
rect 17175 25316 18236 25344
rect 17175 25313 17187 25316
rect 17129 25307 17187 25313
rect 18230 25304 18236 25316
rect 18288 25304 18294 25356
rect 19150 25304 19156 25356
rect 19208 25344 19214 25356
rect 19426 25344 19432 25356
rect 19208 25316 19432 25344
rect 19208 25304 19214 25316
rect 19426 25304 19432 25316
rect 19484 25304 19490 25356
rect 20806 25304 20812 25356
rect 20864 25344 20870 25356
rect 20901 25347 20959 25353
rect 20901 25344 20913 25347
rect 20864 25316 20913 25344
rect 20864 25304 20870 25316
rect 20901 25313 20913 25316
rect 20947 25313 20959 25347
rect 20901 25307 20959 25313
rect 21637 25347 21695 25353
rect 21637 25313 21649 25347
rect 21683 25313 21695 25347
rect 21637 25307 21695 25313
rect 8478 25276 8484 25288
rect 8312 25248 8484 25276
rect 8478 25236 8484 25248
rect 8536 25276 8542 25288
rect 8665 25279 8723 25285
rect 8665 25276 8677 25279
rect 8536 25248 8677 25276
rect 8536 25236 8542 25248
rect 8665 25245 8677 25248
rect 8711 25245 8723 25279
rect 8665 25239 8723 25245
rect 10137 25279 10195 25285
rect 10137 25245 10149 25279
rect 10183 25276 10195 25279
rect 11330 25276 11336 25288
rect 10183 25248 11336 25276
rect 10183 25245 10195 25248
rect 10137 25239 10195 25245
rect 11330 25236 11336 25248
rect 11388 25236 11394 25288
rect 12618 25276 12624 25288
rect 12579 25248 12624 25276
rect 12618 25236 12624 25248
rect 12676 25236 12682 25288
rect 17405 25279 17463 25285
rect 17405 25245 17417 25279
rect 17451 25276 17463 25279
rect 18506 25276 18512 25288
rect 17451 25248 18512 25276
rect 17451 25245 17463 25248
rect 17405 25239 17463 25245
rect 18506 25236 18512 25248
rect 18564 25236 18570 25288
rect 20438 25236 20444 25288
rect 20496 25276 20502 25288
rect 20993 25279 21051 25285
rect 20993 25276 21005 25279
rect 20496 25248 21005 25276
rect 20496 25236 20502 25248
rect 20993 25245 21005 25248
rect 21039 25245 21051 25279
rect 21652 25276 21680 25307
rect 21726 25304 21732 25356
rect 21784 25344 21790 25356
rect 22278 25344 22284 25356
rect 21784 25316 21829 25344
rect 22239 25316 22284 25344
rect 21784 25304 21790 25316
rect 22278 25304 22284 25316
rect 22336 25304 22342 25356
rect 22572 25353 22600 25384
rect 25792 25384 26516 25412
rect 22557 25347 22615 25353
rect 22557 25313 22569 25347
rect 22603 25313 22615 25347
rect 22557 25307 22615 25313
rect 23293 25347 23351 25353
rect 23293 25313 23305 25347
rect 23339 25313 23351 25347
rect 23293 25307 23351 25313
rect 24765 25347 24823 25353
rect 24765 25313 24777 25347
rect 24811 25344 24823 25347
rect 24854 25344 24860 25356
rect 24811 25316 24860 25344
rect 24811 25313 24823 25316
rect 24765 25307 24823 25313
rect 22002 25276 22008 25288
rect 21652 25248 22008 25276
rect 20993 25239 21051 25245
rect 22002 25236 22008 25248
rect 22060 25276 22066 25288
rect 23308 25276 23336 25307
rect 24854 25304 24860 25316
rect 24912 25304 24918 25356
rect 25130 25344 25136 25356
rect 25091 25316 25136 25344
rect 25130 25304 25136 25316
rect 25188 25304 25194 25356
rect 25792 25353 25820 25384
rect 26510 25372 26516 25384
rect 26568 25412 26574 25424
rect 29270 25412 29276 25424
rect 26568 25384 27384 25412
rect 29231 25384 29276 25412
rect 26568 25372 26574 25384
rect 25777 25347 25835 25353
rect 25777 25313 25789 25347
rect 25823 25313 25835 25347
rect 26602 25344 26608 25356
rect 26563 25316 26608 25344
rect 25777 25307 25835 25313
rect 26602 25304 26608 25316
rect 26660 25304 26666 25356
rect 27356 25353 27384 25384
rect 29270 25372 29276 25384
rect 29328 25372 29334 25424
rect 27065 25347 27123 25353
rect 27065 25313 27077 25347
rect 27111 25313 27123 25347
rect 27065 25307 27123 25313
rect 27341 25347 27399 25353
rect 27341 25313 27353 25347
rect 27387 25313 27399 25347
rect 27341 25307 27399 25313
rect 28629 25347 28687 25353
rect 28629 25313 28641 25347
rect 28675 25344 28687 25347
rect 28902 25344 28908 25356
rect 28675 25316 28908 25344
rect 28675 25313 28687 25316
rect 28629 25307 28687 25313
rect 22060 25248 23336 25276
rect 24949 25279 25007 25285
rect 22060 25236 22066 25248
rect 24949 25245 24961 25279
rect 24995 25276 25007 25279
rect 27080 25276 27108 25307
rect 28902 25304 28908 25316
rect 28960 25304 28966 25356
rect 29914 25344 29920 25356
rect 29875 25316 29920 25344
rect 29914 25304 29920 25316
rect 29972 25304 29978 25356
rect 30285 25347 30343 25353
rect 30285 25313 30297 25347
rect 30331 25344 30343 25347
rect 30929 25347 30987 25353
rect 30331 25316 30880 25344
rect 30331 25313 30343 25316
rect 30285 25307 30343 25313
rect 30006 25276 30012 25288
rect 24995 25248 27108 25276
rect 29967 25248 30012 25276
rect 24995 25245 25007 25248
rect 24949 25239 25007 25245
rect 30006 25236 30012 25248
rect 30064 25236 30070 25288
rect 30374 25276 30380 25288
rect 30335 25248 30380 25276
rect 30374 25236 30380 25248
rect 30432 25236 30438 25288
rect 30852 25276 30880 25316
rect 30929 25313 30941 25347
rect 30975 25344 30987 25347
rect 31018 25344 31024 25356
rect 30975 25316 31024 25344
rect 30975 25313 30987 25316
rect 30929 25307 30987 25313
rect 31018 25304 31024 25316
rect 31076 25304 31082 25356
rect 32309 25347 32367 25353
rect 32309 25313 32321 25347
rect 32355 25313 32367 25347
rect 32490 25344 32496 25356
rect 32451 25316 32496 25344
rect 32309 25307 32367 25313
rect 32324 25276 32352 25307
rect 32490 25304 32496 25316
rect 32548 25304 32554 25356
rect 32692 25353 32720 25452
rect 33505 25449 33517 25483
rect 33551 25480 33563 25483
rect 33594 25480 33600 25492
rect 33551 25452 33600 25480
rect 33551 25449 33563 25452
rect 33505 25443 33563 25449
rect 33594 25440 33600 25452
rect 33652 25480 33658 25492
rect 34054 25480 34060 25492
rect 33652 25452 34060 25480
rect 33652 25440 33658 25452
rect 34054 25440 34060 25452
rect 34112 25440 34118 25492
rect 34517 25415 34575 25421
rect 34517 25381 34529 25415
rect 34563 25412 34575 25415
rect 34606 25412 34612 25424
rect 34563 25384 34612 25412
rect 34563 25381 34575 25384
rect 34517 25375 34575 25381
rect 34606 25372 34612 25384
rect 34664 25372 34670 25424
rect 35069 25415 35127 25421
rect 35069 25381 35081 25415
rect 35115 25412 35127 25415
rect 35158 25412 35164 25424
rect 35115 25384 35164 25412
rect 35115 25381 35127 25384
rect 35069 25375 35127 25381
rect 35158 25372 35164 25384
rect 35216 25372 35222 25424
rect 38194 25412 38200 25424
rect 38155 25384 38200 25412
rect 38194 25372 38200 25384
rect 38252 25372 38258 25424
rect 32677 25347 32735 25353
rect 32677 25313 32689 25347
rect 32723 25313 32735 25347
rect 33318 25344 33324 25356
rect 33231 25316 33324 25344
rect 32677 25307 32735 25313
rect 33318 25304 33324 25316
rect 33376 25344 33382 25356
rect 34330 25344 34336 25356
rect 33376 25316 34336 25344
rect 33376 25304 33382 25316
rect 34330 25304 34336 25316
rect 34388 25304 34394 25356
rect 34701 25347 34759 25353
rect 34701 25313 34713 25347
rect 34747 25344 34759 25347
rect 34790 25344 34796 25356
rect 34747 25316 34796 25344
rect 34747 25313 34759 25316
rect 34701 25307 34759 25313
rect 34790 25304 34796 25316
rect 34848 25304 34854 25356
rect 35434 25304 35440 25356
rect 35492 25344 35498 25356
rect 35529 25347 35587 25353
rect 35529 25344 35541 25347
rect 35492 25316 35541 25344
rect 35492 25304 35498 25316
rect 35529 25313 35541 25316
rect 35575 25313 35587 25347
rect 35529 25307 35587 25313
rect 35618 25304 35624 25356
rect 35676 25344 35682 25356
rect 35989 25347 36047 25353
rect 35989 25344 36001 25347
rect 35676 25316 36001 25344
rect 35676 25304 35682 25316
rect 35989 25313 36001 25316
rect 36035 25313 36047 25347
rect 36538 25344 36544 25356
rect 36499 25316 36544 25344
rect 35989 25307 36047 25313
rect 36538 25304 36544 25316
rect 36596 25304 36602 25356
rect 36630 25304 36636 25356
rect 36688 25344 36694 25356
rect 36725 25347 36783 25353
rect 36725 25344 36737 25347
rect 36688 25316 36737 25344
rect 36688 25304 36694 25316
rect 36725 25313 36737 25316
rect 36771 25313 36783 25347
rect 36725 25307 36783 25313
rect 38286 25304 38292 25356
rect 38344 25344 38350 25356
rect 38344 25316 38389 25344
rect 38344 25304 38350 25316
rect 33410 25276 33416 25288
rect 30852 25248 33416 25276
rect 33410 25236 33416 25248
rect 33468 25236 33474 25288
rect 38746 25276 38752 25288
rect 38707 25248 38752 25276
rect 38746 25236 38752 25248
rect 38804 25236 38810 25288
rect 3970 25168 3976 25220
rect 4028 25208 4034 25220
rect 7190 25208 7196 25220
rect 4028 25180 7196 25208
rect 4028 25168 4034 25180
rect 7190 25168 7196 25180
rect 7248 25168 7254 25220
rect 8386 25168 8392 25220
rect 8444 25208 8450 25220
rect 8570 25208 8576 25220
rect 8444 25180 8576 25208
rect 8444 25168 8450 25180
rect 8570 25168 8576 25180
rect 8628 25168 8634 25220
rect 30558 25168 30564 25220
rect 30616 25208 30622 25220
rect 31110 25208 31116 25220
rect 30616 25180 31116 25208
rect 30616 25168 30622 25180
rect 31110 25168 31116 25180
rect 31168 25168 31174 25220
rect 36906 25208 36912 25220
rect 36867 25180 36912 25208
rect 36906 25168 36912 25180
rect 36964 25168 36970 25220
rect 14366 25100 14372 25152
rect 14424 25140 14430 25152
rect 14645 25143 14703 25149
rect 14645 25140 14657 25143
rect 14424 25112 14657 25140
rect 14424 25100 14430 25112
rect 14645 25109 14657 25112
rect 14691 25109 14703 25143
rect 14645 25103 14703 25109
rect 23750 25100 23756 25152
rect 23808 25140 23814 25152
rect 25314 25140 25320 25152
rect 23808 25112 25320 25140
rect 23808 25100 23814 25112
rect 25314 25100 25320 25112
rect 25372 25140 25378 25152
rect 25869 25143 25927 25149
rect 25869 25140 25881 25143
rect 25372 25112 25881 25140
rect 25372 25100 25378 25112
rect 25869 25109 25881 25112
rect 25915 25109 25927 25143
rect 25869 25103 25927 25109
rect 28721 25143 28779 25149
rect 28721 25109 28733 25143
rect 28767 25140 28779 25143
rect 28994 25140 29000 25152
rect 28767 25112 29000 25140
rect 28767 25109 28779 25112
rect 28721 25103 28779 25109
rect 28994 25100 29000 25112
rect 29052 25100 29058 25152
rect 36538 25100 36544 25152
rect 36596 25140 36602 25152
rect 38013 25143 38071 25149
rect 38013 25140 38025 25143
rect 36596 25112 38025 25140
rect 36596 25100 36602 25112
rect 38013 25109 38025 25112
rect 38059 25109 38071 25143
rect 38013 25103 38071 25109
rect 1104 25050 39836 25072
rect 1104 24998 4246 25050
rect 4298 24998 4310 25050
rect 4362 24998 4374 25050
rect 4426 24998 4438 25050
rect 4490 24998 34966 25050
rect 35018 24998 35030 25050
rect 35082 24998 35094 25050
rect 35146 24998 35158 25050
rect 35210 24998 39836 25050
rect 1104 24976 39836 24998
rect 1673 24939 1731 24945
rect 1673 24905 1685 24939
rect 1719 24936 1731 24939
rect 5629 24939 5687 24945
rect 1719 24908 5580 24936
rect 1719 24905 1731 24908
rect 1673 24899 1731 24905
rect 2774 24828 2780 24880
rect 2832 24868 2838 24880
rect 3418 24868 3424 24880
rect 2832 24840 3424 24868
rect 2832 24828 2838 24840
rect 3418 24828 3424 24840
rect 3476 24868 3482 24880
rect 5552 24868 5580 24908
rect 5629 24905 5641 24939
rect 5675 24936 5687 24939
rect 5718 24936 5724 24948
rect 5675 24908 5724 24936
rect 5675 24905 5687 24908
rect 5629 24899 5687 24905
rect 5718 24896 5724 24908
rect 5776 24896 5782 24948
rect 15197 24939 15255 24945
rect 15197 24905 15209 24939
rect 15243 24936 15255 24939
rect 15378 24936 15384 24948
rect 15243 24908 15384 24936
rect 15243 24905 15255 24908
rect 15197 24899 15255 24905
rect 8202 24868 8208 24880
rect 3476 24840 4108 24868
rect 5552 24840 8208 24868
rect 3476 24828 3482 24840
rect 2866 24760 2872 24812
rect 2924 24800 2930 24812
rect 4080 24809 4108 24840
rect 8202 24828 8208 24840
rect 8260 24828 8266 24880
rect 11514 24868 11520 24880
rect 10428 24840 11520 24868
rect 3053 24803 3111 24809
rect 3053 24800 3065 24803
rect 2924 24772 3065 24800
rect 2924 24760 2930 24772
rect 3053 24769 3065 24772
rect 3099 24769 3111 24803
rect 3053 24763 3111 24769
rect 4065 24803 4123 24809
rect 4065 24769 4077 24803
rect 4111 24769 4123 24803
rect 4065 24763 4123 24769
rect 4341 24803 4399 24809
rect 4341 24769 4353 24803
rect 4387 24800 4399 24803
rect 4982 24800 4988 24812
rect 4387 24772 4988 24800
rect 4387 24769 4399 24772
rect 4341 24763 4399 24769
rect 4982 24760 4988 24772
rect 5040 24760 5046 24812
rect 7006 24760 7012 24812
rect 7064 24800 7070 24812
rect 9858 24800 9864 24812
rect 7064 24772 8524 24800
rect 7064 24760 7070 24772
rect 1578 24732 1584 24744
rect 1539 24704 1584 24732
rect 1578 24692 1584 24704
rect 1636 24692 1642 24744
rect 2222 24732 2228 24744
rect 2183 24704 2228 24732
rect 2222 24692 2228 24704
rect 2280 24732 2286 24744
rect 2682 24732 2688 24744
rect 2280 24704 2688 24732
rect 2280 24692 2286 24704
rect 2682 24692 2688 24704
rect 2740 24692 2746 24744
rect 2958 24732 2964 24744
rect 2919 24704 2964 24732
rect 2958 24692 2964 24704
rect 3016 24692 3022 24744
rect 7101 24735 7159 24741
rect 7101 24701 7113 24735
rect 7147 24732 7159 24735
rect 7374 24732 7380 24744
rect 7147 24704 7380 24732
rect 7147 24701 7159 24704
rect 7101 24695 7159 24701
rect 7374 24692 7380 24704
rect 7432 24692 7438 24744
rect 7469 24735 7527 24741
rect 7469 24701 7481 24735
rect 7515 24732 7527 24735
rect 7558 24732 7564 24744
rect 7515 24704 7564 24732
rect 7515 24701 7527 24704
rect 7469 24695 7527 24701
rect 6270 24624 6276 24676
rect 6328 24664 6334 24676
rect 7193 24667 7251 24673
rect 7193 24664 7205 24667
rect 6328 24636 7205 24664
rect 6328 24624 6334 24636
rect 7193 24633 7205 24636
rect 7239 24633 7251 24667
rect 7193 24627 7251 24633
rect 7484 24664 7512 24695
rect 7558 24692 7564 24704
rect 7616 24692 7622 24744
rect 7650 24692 7656 24744
rect 7708 24732 7714 24744
rect 8021 24735 8079 24741
rect 8021 24732 8033 24735
rect 7708 24704 8033 24732
rect 7708 24692 7714 24704
rect 8021 24701 8033 24704
rect 8067 24732 8079 24735
rect 8110 24732 8116 24744
rect 8067 24704 8116 24732
rect 8067 24701 8079 24704
rect 8021 24695 8079 24701
rect 8110 24692 8116 24704
rect 8168 24692 8174 24744
rect 8297 24735 8355 24741
rect 8297 24701 8309 24735
rect 8343 24732 8355 24735
rect 8386 24732 8392 24744
rect 8343 24704 8392 24732
rect 8343 24701 8355 24704
rect 8297 24695 8355 24701
rect 8386 24692 8392 24704
rect 8444 24692 8450 24744
rect 8496 24741 8524 24772
rect 9508 24772 9864 24800
rect 9508 24741 9536 24772
rect 9858 24760 9864 24772
rect 9916 24760 9922 24812
rect 10428 24809 10456 24840
rect 11514 24828 11520 24840
rect 11572 24828 11578 24880
rect 13814 24868 13820 24880
rect 13775 24840 13820 24868
rect 13814 24828 13820 24840
rect 13872 24828 13878 24880
rect 10413 24803 10471 24809
rect 10413 24769 10425 24803
rect 10459 24769 10471 24803
rect 10413 24763 10471 24769
rect 11330 24760 11336 24812
rect 11388 24800 11394 24812
rect 12529 24803 12587 24809
rect 12529 24800 12541 24803
rect 11388 24772 12541 24800
rect 11388 24760 11394 24772
rect 12529 24769 12541 24772
rect 12575 24769 12587 24803
rect 15212 24800 15240 24899
rect 15378 24896 15384 24908
rect 15436 24896 15442 24948
rect 18506 24936 18512 24948
rect 18467 24908 18512 24936
rect 18506 24896 18512 24908
rect 18564 24896 18570 24948
rect 23017 24939 23075 24945
rect 23017 24905 23029 24939
rect 23063 24936 23075 24939
rect 24394 24936 24400 24948
rect 23063 24908 24400 24936
rect 23063 24905 23075 24908
rect 23017 24899 23075 24905
rect 24394 24896 24400 24908
rect 24452 24936 24458 24948
rect 25498 24936 25504 24948
rect 24452 24908 25504 24936
rect 24452 24896 24458 24908
rect 25498 24896 25504 24908
rect 25556 24896 25562 24948
rect 26510 24936 26516 24948
rect 26471 24908 26516 24936
rect 26510 24896 26516 24908
rect 26568 24896 26574 24948
rect 16117 24871 16175 24877
rect 16117 24837 16129 24871
rect 16163 24868 16175 24871
rect 16206 24868 16212 24880
rect 16163 24840 16212 24868
rect 16163 24837 16175 24840
rect 16117 24831 16175 24837
rect 16206 24828 16212 24840
rect 16264 24828 16270 24880
rect 20806 24868 20812 24880
rect 20364 24840 20812 24868
rect 16758 24800 16764 24812
rect 12529 24763 12587 24769
rect 14016 24772 15240 24800
rect 16224 24772 16528 24800
rect 16719 24772 16764 24800
rect 8481 24735 8539 24741
rect 8481 24701 8493 24735
rect 8527 24701 8539 24735
rect 8481 24695 8539 24701
rect 9493 24735 9551 24741
rect 9493 24701 9505 24735
rect 9539 24701 9551 24735
rect 9766 24732 9772 24744
rect 9727 24704 9772 24732
rect 9493 24695 9551 24701
rect 9766 24692 9772 24704
rect 9824 24692 9830 24744
rect 9950 24732 9956 24744
rect 9911 24704 9956 24732
rect 9950 24692 9956 24704
rect 10008 24692 10014 24744
rect 11054 24732 11060 24744
rect 11015 24704 11060 24732
rect 11054 24692 11060 24704
rect 11112 24692 11118 24744
rect 11241 24735 11299 24741
rect 11241 24701 11253 24735
rect 11287 24701 11299 24735
rect 11422 24732 11428 24744
rect 11383 24704 11428 24732
rect 11241 24695 11299 24701
rect 10226 24664 10232 24676
rect 7484 24636 10232 24664
rect 2317 24599 2375 24605
rect 2317 24565 2329 24599
rect 2363 24596 2375 24599
rect 2406 24596 2412 24608
rect 2363 24568 2412 24596
rect 2363 24565 2375 24568
rect 2317 24559 2375 24565
rect 2406 24556 2412 24568
rect 2464 24556 2470 24608
rect 5810 24556 5816 24608
rect 5868 24596 5874 24608
rect 7484 24596 7512 24636
rect 10226 24624 10232 24636
rect 10284 24624 10290 24676
rect 5868 24568 7512 24596
rect 5868 24556 5874 24568
rect 8110 24556 8116 24608
rect 8168 24596 8174 24608
rect 10502 24596 10508 24608
rect 8168 24568 10508 24596
rect 8168 24556 8174 24568
rect 10502 24556 10508 24568
rect 10560 24556 10566 24608
rect 11256 24596 11284 24695
rect 11422 24692 11428 24704
rect 11480 24692 11486 24744
rect 11514 24692 11520 24744
rect 11572 24732 11578 24744
rect 14016 24741 14044 24772
rect 12437 24735 12495 24741
rect 12437 24732 12449 24735
rect 11572 24704 12449 24732
rect 11572 24692 11578 24704
rect 12437 24701 12449 24704
rect 12483 24701 12495 24735
rect 12437 24695 12495 24701
rect 14001 24735 14059 24741
rect 14001 24701 14013 24735
rect 14047 24701 14059 24735
rect 14001 24695 14059 24701
rect 14185 24735 14243 24741
rect 14185 24701 14197 24735
rect 14231 24701 14243 24735
rect 14185 24695 14243 24701
rect 14369 24735 14427 24741
rect 14369 24701 14381 24735
rect 14415 24701 14427 24735
rect 14369 24695 14427 24701
rect 11882 24624 11888 24676
rect 11940 24664 11946 24676
rect 14200 24664 14228 24695
rect 11940 24636 14228 24664
rect 14384 24664 14412 24695
rect 14550 24692 14556 24744
rect 14608 24732 14614 24744
rect 15013 24735 15071 24741
rect 15013 24732 15025 24735
rect 14608 24704 15025 24732
rect 14608 24692 14614 24704
rect 15013 24701 15025 24704
rect 15059 24732 15071 24735
rect 16224 24732 16252 24772
rect 15059 24704 16252 24732
rect 16301 24735 16359 24741
rect 15059 24701 15071 24704
rect 15013 24695 15071 24701
rect 16301 24701 16313 24735
rect 16347 24732 16359 24735
rect 16390 24732 16396 24744
rect 16347 24704 16396 24732
rect 16347 24701 16359 24704
rect 16301 24695 16359 24701
rect 15470 24664 15476 24676
rect 14384 24636 15476 24664
rect 11940 24624 11946 24636
rect 15470 24624 15476 24636
rect 15528 24624 15534 24676
rect 12434 24596 12440 24608
rect 11256 24568 12440 24596
rect 12434 24556 12440 24568
rect 12492 24556 12498 24608
rect 15654 24556 15660 24608
rect 15712 24596 15718 24608
rect 16316 24596 16344 24695
rect 16390 24692 16396 24704
rect 16448 24692 16454 24744
rect 16500 24732 16528 24772
rect 16758 24760 16764 24772
rect 16816 24760 16822 24812
rect 18046 24800 18052 24812
rect 18007 24772 18052 24800
rect 18046 24760 18052 24772
rect 18104 24760 18110 24812
rect 16666 24732 16672 24744
rect 16500 24704 16672 24732
rect 16666 24692 16672 24704
rect 16724 24692 16730 24744
rect 17313 24735 17371 24741
rect 17313 24701 17325 24735
rect 17359 24701 17371 24735
rect 17313 24695 17371 24701
rect 17328 24664 17356 24695
rect 17494 24692 17500 24744
rect 17552 24732 17558 24744
rect 18325 24735 18383 24741
rect 18325 24732 18337 24735
rect 17552 24704 18337 24732
rect 17552 24692 17558 24704
rect 18325 24701 18337 24704
rect 18371 24701 18383 24735
rect 19797 24735 19855 24741
rect 19797 24732 19809 24735
rect 18325 24695 18383 24701
rect 19352 24704 19809 24732
rect 18138 24664 18144 24676
rect 17328 24636 18144 24664
rect 18138 24624 18144 24636
rect 18196 24624 18202 24676
rect 18230 24624 18236 24676
rect 18288 24664 18294 24676
rect 18288 24636 18333 24664
rect 18288 24624 18294 24636
rect 15712 24568 16344 24596
rect 17405 24599 17463 24605
rect 15712 24556 15718 24568
rect 17405 24565 17417 24599
rect 17451 24596 17463 24599
rect 19352 24596 19380 24704
rect 19797 24701 19809 24704
rect 19843 24732 19855 24735
rect 20364 24732 20392 24840
rect 20806 24828 20812 24840
rect 20864 24828 20870 24880
rect 22186 24868 22192 24880
rect 21192 24840 22192 24868
rect 20441 24803 20499 24809
rect 20441 24769 20453 24803
rect 20487 24800 20499 24803
rect 21082 24800 21088 24812
rect 20487 24772 21088 24800
rect 20487 24769 20499 24772
rect 20441 24763 20499 24769
rect 21082 24760 21088 24772
rect 21140 24760 21146 24812
rect 19843 24704 20392 24732
rect 20533 24735 20591 24741
rect 19843 24701 19855 24704
rect 19797 24695 19855 24701
rect 20533 24701 20545 24735
rect 20579 24701 20591 24735
rect 20806 24732 20812 24744
rect 20767 24704 20812 24732
rect 20533 24695 20591 24701
rect 20548 24664 20576 24695
rect 20806 24692 20812 24704
rect 20864 24692 20870 24744
rect 21192 24741 21220 24840
rect 22186 24828 22192 24840
rect 22244 24828 22250 24880
rect 29914 24828 29920 24880
rect 29972 24868 29978 24880
rect 30009 24871 30067 24877
rect 30009 24868 30021 24871
rect 29972 24840 30021 24868
rect 29972 24828 29978 24840
rect 30009 24837 30021 24840
rect 30055 24837 30067 24871
rect 30009 24831 30067 24837
rect 22281 24803 22339 24809
rect 22281 24769 22293 24803
rect 22327 24800 22339 24803
rect 23658 24800 23664 24812
rect 22327 24772 23664 24800
rect 22327 24769 22339 24772
rect 22281 24763 22339 24769
rect 23658 24760 23664 24772
rect 23716 24800 23722 24812
rect 24210 24800 24216 24812
rect 23716 24772 24216 24800
rect 23716 24760 23722 24772
rect 24210 24760 24216 24772
rect 24268 24760 24274 24812
rect 25406 24800 25412 24812
rect 25367 24772 25412 24800
rect 25406 24760 25412 24772
rect 25464 24760 25470 24812
rect 27985 24803 28043 24809
rect 27985 24769 27997 24803
rect 28031 24800 28043 24803
rect 29178 24800 29184 24812
rect 28031 24772 29184 24800
rect 28031 24769 28043 24772
rect 27985 24763 28043 24769
rect 29178 24760 29184 24772
rect 29236 24760 29242 24812
rect 31757 24803 31815 24809
rect 29472 24772 30144 24800
rect 21177 24735 21235 24741
rect 21177 24701 21189 24735
rect 21223 24701 21235 24735
rect 21177 24695 21235 24701
rect 21453 24735 21511 24741
rect 21453 24701 21465 24735
rect 21499 24701 21511 24735
rect 22186 24732 22192 24744
rect 22147 24704 22192 24732
rect 21453 24695 21511 24701
rect 20714 24664 20720 24676
rect 20548 24636 20720 24664
rect 20714 24624 20720 24636
rect 20772 24624 20778 24676
rect 17451 24568 19380 24596
rect 17451 24565 17463 24568
rect 17405 24559 17463 24565
rect 19426 24556 19432 24608
rect 19484 24596 19490 24608
rect 21468 24596 21496 24695
rect 22186 24692 22192 24704
rect 22244 24692 22250 24744
rect 22833 24735 22891 24741
rect 22833 24732 22845 24735
rect 22296 24704 22845 24732
rect 22296 24676 22324 24704
rect 22833 24701 22845 24704
rect 22879 24732 22891 24735
rect 22922 24732 22928 24744
rect 22879 24704 22928 24732
rect 22879 24701 22891 24704
rect 22833 24695 22891 24701
rect 22922 24692 22928 24704
rect 22980 24692 22986 24744
rect 23842 24692 23848 24744
rect 23900 24732 23906 24744
rect 24029 24735 24087 24741
rect 24029 24732 24041 24735
rect 23900 24704 24041 24732
rect 23900 24692 23906 24704
rect 24029 24701 24041 24704
rect 24075 24701 24087 24735
rect 25130 24732 25136 24744
rect 25091 24704 25136 24732
rect 24029 24695 24087 24701
rect 25130 24692 25136 24704
rect 25188 24692 25194 24744
rect 28258 24732 28264 24744
rect 28219 24704 28264 24732
rect 28258 24692 28264 24704
rect 28316 24692 28322 24744
rect 28445 24735 28503 24741
rect 28445 24701 28457 24735
rect 28491 24701 28503 24735
rect 28445 24695 28503 24701
rect 22278 24624 22284 24676
rect 22336 24624 22342 24676
rect 26786 24624 26792 24676
rect 26844 24664 26850 24676
rect 27433 24667 27491 24673
rect 27433 24664 27445 24667
rect 26844 24636 27445 24664
rect 26844 24624 26850 24636
rect 27433 24633 27445 24636
rect 27479 24633 27491 24667
rect 27433 24627 27491 24633
rect 27614 24624 27620 24676
rect 27672 24664 27678 24676
rect 28460 24664 28488 24695
rect 28626 24692 28632 24744
rect 28684 24732 28690 24744
rect 29472 24732 29500 24772
rect 30116 24741 30144 24772
rect 31757 24769 31769 24803
rect 31803 24800 31815 24803
rect 34606 24800 34612 24812
rect 31803 24772 34612 24800
rect 31803 24769 31815 24772
rect 31757 24763 31815 24769
rect 34606 24760 34612 24772
rect 34664 24760 34670 24812
rect 34882 24760 34888 24812
rect 34940 24800 34946 24812
rect 35434 24800 35440 24812
rect 34940 24772 35440 24800
rect 34940 24760 34946 24772
rect 35434 24760 35440 24772
rect 35492 24760 35498 24812
rect 36998 24760 37004 24812
rect 37056 24800 37062 24812
rect 37277 24803 37335 24809
rect 37277 24800 37289 24803
rect 37056 24772 37289 24800
rect 37056 24760 37062 24772
rect 37277 24769 37289 24772
rect 37323 24800 37335 24803
rect 37458 24800 37464 24812
rect 37323 24772 37464 24800
rect 37323 24769 37335 24772
rect 37277 24763 37335 24769
rect 37458 24760 37464 24772
rect 37516 24760 37522 24812
rect 38286 24760 38292 24812
rect 38344 24800 38350 24812
rect 38657 24803 38715 24809
rect 38657 24800 38669 24803
rect 38344 24772 38669 24800
rect 38344 24760 38350 24772
rect 38657 24769 38669 24772
rect 38703 24769 38715 24803
rect 38657 24763 38715 24769
rect 28684 24704 29500 24732
rect 29549 24735 29607 24741
rect 28684 24692 28690 24704
rect 29549 24701 29561 24735
rect 29595 24701 29607 24735
rect 29549 24695 29607 24701
rect 30101 24735 30159 24741
rect 30101 24701 30113 24735
rect 30147 24701 30159 24735
rect 30101 24695 30159 24701
rect 30285 24735 30343 24741
rect 30285 24701 30297 24735
rect 30331 24732 30343 24735
rect 30650 24732 30656 24744
rect 30331 24704 30656 24732
rect 30331 24701 30343 24704
rect 30285 24695 30343 24701
rect 27672 24636 28488 24664
rect 29564 24664 29592 24695
rect 30650 24692 30656 24704
rect 30708 24692 30714 24744
rect 31018 24732 31024 24744
rect 30760 24704 31024 24732
rect 29564 24636 30512 24664
rect 27672 24624 27678 24636
rect 30484 24608 30512 24636
rect 30558 24624 30564 24676
rect 30616 24664 30622 24676
rect 30760 24664 30788 24704
rect 31018 24692 31024 24704
rect 31076 24732 31082 24744
rect 31297 24735 31355 24741
rect 31297 24732 31309 24735
rect 31076 24704 31309 24732
rect 31076 24692 31082 24704
rect 31297 24701 31309 24704
rect 31343 24701 31355 24735
rect 31662 24732 31668 24744
rect 31623 24704 31668 24732
rect 31297 24695 31355 24701
rect 31662 24692 31668 24704
rect 31720 24692 31726 24744
rect 32214 24692 32220 24744
rect 32272 24732 32278 24744
rect 32309 24735 32367 24741
rect 32309 24732 32321 24735
rect 32272 24704 32321 24732
rect 32272 24692 32278 24704
rect 32309 24701 32321 24704
rect 32355 24701 32367 24735
rect 32582 24732 32588 24744
rect 32543 24704 32588 24732
rect 32309 24695 32367 24701
rect 32582 24692 32588 24704
rect 32640 24692 32646 24744
rect 35250 24692 35256 24744
rect 35308 24732 35314 24744
rect 35529 24735 35587 24741
rect 35529 24732 35541 24735
rect 35308 24704 35541 24732
rect 35308 24692 35314 24704
rect 35529 24701 35541 24704
rect 35575 24701 35587 24735
rect 35529 24695 35587 24701
rect 35710 24692 35716 24744
rect 35768 24732 35774 24744
rect 35897 24735 35955 24741
rect 35897 24732 35909 24735
rect 35768 24704 35909 24732
rect 35768 24692 35774 24704
rect 35897 24701 35909 24704
rect 35943 24701 35955 24735
rect 35897 24695 35955 24701
rect 36081 24735 36139 24741
rect 36081 24701 36093 24735
rect 36127 24701 36139 24735
rect 36081 24695 36139 24701
rect 30616 24636 30788 24664
rect 30837 24667 30895 24673
rect 30616 24624 30622 24636
rect 30837 24633 30849 24667
rect 30883 24664 30895 24667
rect 32398 24664 32404 24676
rect 30883 24636 32404 24664
rect 30883 24633 30895 24636
rect 30837 24627 30895 24633
rect 32398 24624 32404 24636
rect 32456 24624 32462 24676
rect 33318 24624 33324 24676
rect 33376 24664 33382 24676
rect 34514 24664 34520 24676
rect 33376 24636 34520 24664
rect 33376 24624 33382 24636
rect 34514 24624 34520 24636
rect 34572 24624 34578 24676
rect 34885 24667 34943 24673
rect 34885 24633 34897 24667
rect 34931 24664 34943 24667
rect 35066 24664 35072 24676
rect 34931 24636 35072 24664
rect 34931 24633 34943 24636
rect 34885 24627 34943 24633
rect 35066 24624 35072 24636
rect 35124 24624 35130 24676
rect 36096 24664 36124 24695
rect 36354 24692 36360 24744
rect 36412 24732 36418 24744
rect 36541 24735 36599 24741
rect 36541 24732 36553 24735
rect 36412 24704 36553 24732
rect 36412 24692 36418 24704
rect 36541 24701 36553 24704
rect 36587 24701 36599 24735
rect 36541 24695 36599 24701
rect 37366 24692 37372 24744
rect 37424 24732 37430 24744
rect 37553 24735 37611 24741
rect 37553 24732 37565 24735
rect 37424 24704 37565 24732
rect 37424 24692 37430 24704
rect 37553 24701 37565 24704
rect 37599 24701 37611 24735
rect 37553 24695 37611 24701
rect 36096 24636 36400 24664
rect 36372 24608 36400 24636
rect 19484 24568 21496 24596
rect 24213 24599 24271 24605
rect 19484 24556 19490 24568
rect 24213 24565 24225 24599
rect 24259 24596 24271 24599
rect 24302 24596 24308 24608
rect 24259 24568 24308 24596
rect 24259 24565 24271 24568
rect 24213 24559 24271 24565
rect 24302 24556 24308 24568
rect 24360 24556 24366 24608
rect 30466 24556 30472 24608
rect 30524 24596 30530 24608
rect 33689 24599 33747 24605
rect 33689 24596 33701 24599
rect 30524 24568 33701 24596
rect 30524 24556 30530 24568
rect 33689 24565 33701 24568
rect 33735 24565 33747 24599
rect 33689 24559 33747 24565
rect 36354 24556 36360 24608
rect 36412 24556 36418 24608
rect 36722 24596 36728 24608
rect 36683 24568 36728 24596
rect 36722 24556 36728 24568
rect 36780 24596 36786 24608
rect 37918 24596 37924 24608
rect 36780 24568 37924 24596
rect 36780 24556 36786 24568
rect 37918 24556 37924 24568
rect 37976 24556 37982 24608
rect 1104 24506 39836 24528
rect 1104 24454 19606 24506
rect 19658 24454 19670 24506
rect 19722 24454 19734 24506
rect 19786 24454 19798 24506
rect 19850 24454 39836 24506
rect 1104 24432 39836 24454
rect 15930 24392 15936 24404
rect 15891 24364 15936 24392
rect 15930 24352 15936 24364
rect 15988 24352 15994 24404
rect 20257 24395 20315 24401
rect 20257 24361 20269 24395
rect 20303 24392 20315 24395
rect 20714 24392 20720 24404
rect 20303 24364 20720 24392
rect 20303 24361 20315 24364
rect 20257 24355 20315 24361
rect 20714 24352 20720 24364
rect 20772 24392 20778 24404
rect 22002 24392 22008 24404
rect 20772 24364 22008 24392
rect 20772 24352 20778 24364
rect 22002 24352 22008 24364
rect 22060 24352 22066 24404
rect 22094 24352 22100 24404
rect 22152 24392 22158 24404
rect 22152 24364 24164 24392
rect 22152 24352 22158 24364
rect 1670 24284 1676 24336
rect 1728 24324 1734 24336
rect 1857 24327 1915 24333
rect 1857 24324 1869 24327
rect 1728 24296 1869 24324
rect 1728 24284 1734 24296
rect 1857 24293 1869 24296
rect 1903 24293 1915 24327
rect 12986 24324 12992 24336
rect 1857 24287 1915 24293
rect 8220 24296 8340 24324
rect 8220 24268 8248 24296
rect 2406 24256 2412 24268
rect 2367 24228 2412 24256
rect 2406 24216 2412 24228
rect 2464 24216 2470 24268
rect 2685 24259 2743 24265
rect 2685 24225 2697 24259
rect 2731 24256 2743 24259
rect 2774 24256 2780 24268
rect 2731 24228 2780 24256
rect 2731 24225 2743 24228
rect 2685 24219 2743 24225
rect 2774 24216 2780 24228
rect 2832 24216 2838 24268
rect 2869 24259 2927 24265
rect 2869 24225 2881 24259
rect 2915 24256 2927 24259
rect 2958 24256 2964 24268
rect 2915 24228 2964 24256
rect 2915 24225 2927 24228
rect 2869 24219 2927 24225
rect 2958 24216 2964 24228
rect 3016 24216 3022 24268
rect 3329 24259 3387 24265
rect 3329 24225 3341 24259
rect 3375 24256 3387 24259
rect 4341 24259 4399 24265
rect 3375 24228 4200 24256
rect 3375 24225 3387 24228
rect 3329 24219 3387 24225
rect 4172 24129 4200 24228
rect 4341 24225 4353 24259
rect 4387 24256 4399 24259
rect 4522 24256 4528 24268
rect 4387 24228 4528 24256
rect 4387 24225 4399 24228
rect 4341 24219 4399 24225
rect 4522 24216 4528 24228
rect 4580 24216 4586 24268
rect 4801 24259 4859 24265
rect 4801 24225 4813 24259
rect 4847 24256 4859 24259
rect 5534 24256 5540 24268
rect 4847 24228 5540 24256
rect 4847 24225 4859 24228
rect 4801 24219 4859 24225
rect 5534 24216 5540 24228
rect 5592 24216 5598 24268
rect 5905 24259 5963 24265
rect 5905 24225 5917 24259
rect 5951 24225 5963 24259
rect 6270 24256 6276 24268
rect 6231 24228 6276 24256
rect 5905 24219 5963 24225
rect 5445 24191 5503 24197
rect 5445 24157 5457 24191
rect 5491 24188 5503 24191
rect 5810 24188 5816 24200
rect 5491 24160 5816 24188
rect 5491 24157 5503 24160
rect 5445 24151 5503 24157
rect 5810 24148 5816 24160
rect 5868 24148 5874 24200
rect 4157 24123 4215 24129
rect 4157 24089 4169 24123
rect 4203 24089 4215 24123
rect 5920 24120 5948 24219
rect 6270 24216 6276 24228
rect 6328 24216 6334 24268
rect 7006 24256 7012 24268
rect 6967 24228 7012 24256
rect 7006 24216 7012 24228
rect 7064 24216 7070 24268
rect 7561 24259 7619 24265
rect 7561 24225 7573 24259
rect 7607 24225 7619 24259
rect 7742 24256 7748 24268
rect 7703 24228 7748 24256
rect 7561 24219 7619 24225
rect 6178 24188 6184 24200
rect 6139 24160 6184 24188
rect 6178 24148 6184 24160
rect 6236 24148 6242 24200
rect 7466 24120 7472 24132
rect 5920 24092 7472 24120
rect 4157 24083 4215 24089
rect 7466 24080 7472 24092
rect 7524 24080 7530 24132
rect 3421 24055 3479 24061
rect 3421 24021 3433 24055
rect 3467 24052 3479 24055
rect 3694 24052 3700 24064
rect 3467 24024 3700 24052
rect 3467 24021 3479 24024
rect 3421 24015 3479 24021
rect 3694 24012 3700 24024
rect 3752 24012 3758 24064
rect 7576 24052 7604 24219
rect 7742 24216 7748 24228
rect 7800 24216 7806 24268
rect 8202 24216 8208 24268
rect 8260 24216 8266 24268
rect 8312 24256 8340 24296
rect 8404 24296 12992 24324
rect 8404 24256 8432 24296
rect 12986 24284 12992 24296
rect 13044 24284 13050 24336
rect 16206 24284 16212 24336
rect 16264 24324 16270 24336
rect 16264 24296 16344 24324
rect 16264 24284 16270 24296
rect 8312 24228 8432 24256
rect 8478 24216 8484 24268
rect 8536 24256 8542 24268
rect 8573 24259 8631 24265
rect 8573 24256 8585 24259
rect 8536 24228 8585 24256
rect 8536 24216 8542 24228
rect 8573 24225 8585 24228
rect 8619 24225 8631 24259
rect 8573 24219 8631 24225
rect 10137 24259 10195 24265
rect 10137 24225 10149 24259
rect 10183 24225 10195 24259
rect 10318 24256 10324 24268
rect 10279 24228 10324 24256
rect 10137 24219 10195 24225
rect 8113 24191 8171 24197
rect 8113 24157 8125 24191
rect 8159 24188 8171 24191
rect 9398 24188 9404 24200
rect 8159 24160 9404 24188
rect 8159 24157 8171 24160
rect 8113 24151 8171 24157
rect 9398 24148 9404 24160
rect 9456 24148 9462 24200
rect 9858 24148 9864 24200
rect 9916 24188 9922 24200
rect 10152 24188 10180 24219
rect 10318 24216 10324 24228
rect 10376 24216 10382 24268
rect 10502 24256 10508 24268
rect 10463 24228 10508 24256
rect 10502 24216 10508 24228
rect 10560 24216 10566 24268
rect 11146 24256 11152 24268
rect 11107 24228 11152 24256
rect 11146 24216 11152 24228
rect 11204 24256 11210 24268
rect 11606 24256 11612 24268
rect 11204 24228 11612 24256
rect 11204 24216 11210 24228
rect 11606 24216 11612 24228
rect 11664 24216 11670 24268
rect 12713 24259 12771 24265
rect 12713 24225 12725 24259
rect 12759 24225 12771 24259
rect 12713 24219 12771 24225
rect 13081 24259 13139 24265
rect 13081 24225 13093 24259
rect 13127 24256 13139 24259
rect 14277 24259 14335 24265
rect 14277 24256 14289 24259
rect 13127 24228 14289 24256
rect 13127 24225 13139 24228
rect 13081 24219 13139 24225
rect 14277 24225 14289 24228
rect 14323 24256 14335 24259
rect 14366 24256 14372 24268
rect 14323 24228 14372 24256
rect 14323 24225 14335 24228
rect 14277 24219 14335 24225
rect 9916 24160 10180 24188
rect 9916 24148 9922 24160
rect 9950 24120 9956 24132
rect 9911 24092 9956 24120
rect 9950 24080 9956 24092
rect 10008 24080 10014 24132
rect 10152 24120 10180 24160
rect 10226 24148 10232 24200
rect 10284 24188 10290 24200
rect 12253 24191 12311 24197
rect 12253 24188 12265 24191
rect 10284 24160 12265 24188
rect 10284 24148 10290 24160
rect 12253 24157 12265 24160
rect 12299 24157 12311 24191
rect 12728 24188 12756 24219
rect 14366 24216 14372 24228
rect 14424 24216 14430 24268
rect 14458 24216 14464 24268
rect 14516 24256 14522 24268
rect 14553 24259 14611 24265
rect 14553 24256 14565 24259
rect 14516 24228 14565 24256
rect 14516 24216 14522 24228
rect 14553 24225 14565 24228
rect 14599 24225 14611 24259
rect 14553 24219 14611 24225
rect 15289 24259 15347 24265
rect 15289 24225 15301 24259
rect 15335 24256 15347 24259
rect 15470 24256 15476 24268
rect 15335 24228 15476 24256
rect 15335 24225 15347 24228
rect 15289 24219 15347 24225
rect 15470 24216 15476 24228
rect 15528 24216 15534 24268
rect 16022 24216 16028 24268
rect 16080 24256 16086 24268
rect 16316 24265 16344 24296
rect 17126 24284 17132 24336
rect 17184 24324 17190 24336
rect 17184 24296 18460 24324
rect 17184 24284 17190 24296
rect 16125 24259 16183 24265
rect 16125 24256 16137 24259
rect 16080 24228 16137 24256
rect 16080 24216 16086 24228
rect 16125 24225 16137 24228
rect 16171 24225 16183 24259
rect 16125 24219 16183 24225
rect 16301 24259 16359 24265
rect 16301 24225 16313 24259
rect 16347 24225 16359 24259
rect 16301 24219 16359 24225
rect 16945 24259 17003 24265
rect 16945 24225 16957 24259
rect 16991 24256 17003 24259
rect 17218 24256 17224 24268
rect 16991 24228 17224 24256
rect 16991 24225 17003 24228
rect 16945 24219 17003 24225
rect 17218 24216 17224 24228
rect 17276 24216 17282 24268
rect 18230 24256 18236 24268
rect 18191 24228 18236 24256
rect 18230 24216 18236 24228
rect 18288 24216 18294 24268
rect 18432 24265 18460 24296
rect 18506 24284 18512 24336
rect 18564 24324 18570 24336
rect 22738 24324 22744 24336
rect 18564 24296 22744 24324
rect 18564 24284 18570 24296
rect 22738 24284 22744 24296
rect 22796 24284 22802 24336
rect 23014 24324 23020 24336
rect 22975 24296 23020 24324
rect 23014 24284 23020 24296
rect 23072 24284 23078 24336
rect 18417 24259 18475 24265
rect 18417 24225 18429 24259
rect 18463 24225 18475 24259
rect 18417 24219 18475 24225
rect 18601 24259 18659 24265
rect 18601 24225 18613 24259
rect 18647 24225 18659 24259
rect 18601 24219 18659 24225
rect 19245 24259 19303 24265
rect 19245 24225 19257 24259
rect 19291 24256 19303 24259
rect 19886 24256 19892 24268
rect 19291 24228 19892 24256
rect 19291 24225 19303 24228
rect 19245 24219 19303 24225
rect 13725 24191 13783 24197
rect 12728 24160 13676 24188
rect 12253 24151 12311 24157
rect 10962 24120 10968 24132
rect 10152 24092 10968 24120
rect 10962 24080 10968 24092
rect 11020 24120 11026 24132
rect 11333 24123 11391 24129
rect 11333 24120 11345 24123
rect 11020 24092 11345 24120
rect 11020 24080 11026 24092
rect 11333 24089 11345 24092
rect 11379 24089 11391 24123
rect 11333 24083 11391 24089
rect 12618 24080 12624 24132
rect 12676 24120 12682 24132
rect 12989 24123 13047 24129
rect 12989 24120 13001 24123
rect 12676 24092 13001 24120
rect 12676 24080 12682 24092
rect 12989 24089 13001 24092
rect 13035 24089 13047 24123
rect 12989 24083 13047 24089
rect 8386 24052 8392 24064
rect 7576 24024 8392 24052
rect 8386 24012 8392 24024
rect 8444 24052 8450 24064
rect 8754 24052 8760 24064
rect 8444 24024 8760 24052
rect 8444 24012 8450 24024
rect 8754 24012 8760 24024
rect 8812 24052 8818 24064
rect 10318 24052 10324 24064
rect 8812 24024 10324 24052
rect 8812 24012 8818 24024
rect 10318 24012 10324 24024
rect 10376 24012 10382 24064
rect 13648 24052 13676 24160
rect 13725 24157 13737 24191
rect 13771 24188 13783 24191
rect 14734 24188 14740 24200
rect 13771 24160 14228 24188
rect 14695 24160 14740 24188
rect 13771 24157 13783 24160
rect 13725 24151 13783 24157
rect 14200 24120 14228 24160
rect 14734 24148 14740 24160
rect 14792 24148 14798 24200
rect 17037 24191 17095 24197
rect 17037 24188 17049 24191
rect 14844 24160 17049 24188
rect 14844 24120 14872 24160
rect 17037 24157 17049 24160
rect 17083 24157 17095 24191
rect 18616 24188 18644 24219
rect 19886 24216 19892 24228
rect 19944 24216 19950 24268
rect 20070 24256 20076 24268
rect 20031 24228 20076 24256
rect 20070 24216 20076 24228
rect 20128 24216 20134 24268
rect 21361 24259 21419 24265
rect 21361 24225 21373 24259
rect 21407 24256 21419 24259
rect 21634 24256 21640 24268
rect 21407 24228 21496 24256
rect 21595 24228 21640 24256
rect 21407 24225 21419 24228
rect 21361 24219 21419 24225
rect 21468 24188 21496 24228
rect 21634 24216 21640 24228
rect 21692 24216 21698 24268
rect 21726 24216 21732 24268
rect 21784 24256 21790 24268
rect 22281 24259 22339 24265
rect 22281 24256 22293 24259
rect 21784 24228 22293 24256
rect 21784 24216 21790 24228
rect 22281 24225 22293 24228
rect 22327 24225 22339 24259
rect 22281 24219 22339 24225
rect 23290 24216 23296 24268
rect 23348 24256 23354 24268
rect 23661 24259 23719 24265
rect 23661 24256 23673 24259
rect 23348 24228 23673 24256
rect 23348 24216 23354 24228
rect 23661 24225 23673 24228
rect 23707 24225 23719 24259
rect 23661 24219 23719 24225
rect 23750 24216 23756 24268
rect 23808 24256 23814 24268
rect 24026 24256 24032 24268
rect 23808 24228 23853 24256
rect 23987 24228 24032 24256
rect 23808 24216 23814 24228
rect 24026 24216 24032 24228
rect 24084 24216 24090 24268
rect 24136 24265 24164 24364
rect 25682 24352 25688 24404
rect 25740 24392 25746 24404
rect 27157 24395 27215 24401
rect 27157 24392 27169 24395
rect 25740 24364 27169 24392
rect 25740 24352 25746 24364
rect 27157 24361 27169 24364
rect 27203 24361 27215 24395
rect 27157 24355 27215 24361
rect 27338 24352 27344 24404
rect 27396 24392 27402 24404
rect 28534 24392 28540 24404
rect 27396 24364 28540 24392
rect 27396 24352 27402 24364
rect 28534 24352 28540 24364
rect 28592 24352 28598 24404
rect 30377 24395 30435 24401
rect 30377 24392 30389 24395
rect 29840 24364 30389 24392
rect 28629 24327 28687 24333
rect 28629 24324 28641 24327
rect 25608 24296 28641 24324
rect 24121 24259 24179 24265
rect 24121 24225 24133 24259
rect 24167 24225 24179 24259
rect 24854 24256 24860 24268
rect 24815 24228 24860 24256
rect 24121 24219 24179 24225
rect 24854 24216 24860 24228
rect 24912 24216 24918 24268
rect 25314 24216 25320 24268
rect 25372 24256 25378 24268
rect 25608 24265 25636 24296
rect 28629 24293 28641 24296
rect 28675 24293 28687 24327
rect 28629 24287 28687 24293
rect 28902 24284 28908 24336
rect 28960 24324 28966 24336
rect 28960 24296 29684 24324
rect 28960 24284 28966 24296
rect 25593 24259 25651 24265
rect 25593 24256 25605 24259
rect 25372 24228 25605 24256
rect 25372 24216 25378 24228
rect 25593 24225 25605 24228
rect 25639 24225 25651 24259
rect 25774 24256 25780 24268
rect 25735 24228 25780 24256
rect 25593 24219 25651 24225
rect 25774 24216 25780 24228
rect 25832 24216 25838 24268
rect 27338 24256 27344 24268
rect 27299 24228 27344 24256
rect 27338 24216 27344 24228
rect 27396 24216 27402 24268
rect 27614 24256 27620 24268
rect 27575 24228 27620 24256
rect 27614 24216 27620 24228
rect 27672 24216 27678 24268
rect 27893 24259 27951 24265
rect 27893 24225 27905 24259
rect 27939 24256 27951 24259
rect 29178 24256 29184 24268
rect 27939 24228 29184 24256
rect 27939 24225 27951 24228
rect 27893 24219 27951 24225
rect 29178 24216 29184 24228
rect 29236 24216 29242 24268
rect 29656 24265 29684 24296
rect 29840 24265 29868 24364
rect 30377 24361 30389 24364
rect 30423 24361 30435 24395
rect 30377 24355 30435 24361
rect 30834 24352 30840 24404
rect 30892 24392 30898 24404
rect 35894 24392 35900 24404
rect 30892 24364 35900 24392
rect 30892 24352 30898 24364
rect 35894 24352 35900 24364
rect 35952 24352 35958 24404
rect 37274 24352 37280 24404
rect 37332 24392 37338 24404
rect 37829 24395 37887 24401
rect 37829 24392 37841 24395
rect 37332 24364 37841 24392
rect 37332 24352 37338 24364
rect 37829 24361 37841 24364
rect 37875 24361 37887 24395
rect 37829 24355 37887 24361
rect 30006 24284 30012 24336
rect 30064 24324 30070 24336
rect 34882 24324 34888 24336
rect 30064 24296 34888 24324
rect 30064 24284 30070 24296
rect 29273 24259 29331 24265
rect 29273 24225 29285 24259
rect 29319 24256 29331 24259
rect 29641 24259 29699 24265
rect 29319 24228 29592 24256
rect 29319 24225 29331 24228
rect 29273 24219 29331 24225
rect 29362 24188 29368 24200
rect 17037 24151 17095 24157
rect 17788 24160 18644 24188
rect 18708 24160 21312 24188
rect 21468 24160 28212 24188
rect 29323 24160 29368 24188
rect 14200 24092 14872 24120
rect 16485 24123 16543 24129
rect 16485 24089 16497 24123
rect 16531 24089 16543 24123
rect 16485 24083 16543 24089
rect 14458 24052 14464 24064
rect 13648 24024 14464 24052
rect 14458 24012 14464 24024
rect 14516 24012 14522 24064
rect 14550 24012 14556 24064
rect 14608 24052 14614 24064
rect 15381 24055 15439 24061
rect 15381 24052 15393 24055
rect 14608 24024 15393 24052
rect 14608 24012 14614 24024
rect 15381 24021 15393 24024
rect 15427 24021 15439 24055
rect 16500 24052 16528 24083
rect 16666 24080 16672 24132
rect 16724 24120 16730 24132
rect 17788 24120 17816 24160
rect 18046 24120 18052 24132
rect 16724 24092 17816 24120
rect 18007 24092 18052 24120
rect 16724 24080 16730 24092
rect 18046 24080 18052 24092
rect 18104 24080 18110 24132
rect 18138 24080 18144 24132
rect 18196 24120 18202 24132
rect 18708 24120 18736 24160
rect 18196 24092 18736 24120
rect 18196 24080 18202 24092
rect 19334 24080 19340 24132
rect 19392 24120 19398 24132
rect 20622 24120 20628 24132
rect 19392 24092 20628 24120
rect 19392 24080 19398 24092
rect 20622 24080 20628 24092
rect 20680 24080 20686 24132
rect 21174 24120 21180 24132
rect 21135 24092 21180 24120
rect 21174 24080 21180 24092
rect 21232 24080 21238 24132
rect 21284 24120 21312 24160
rect 21634 24120 21640 24132
rect 21284 24092 21640 24120
rect 21634 24080 21640 24092
rect 21692 24080 21698 24132
rect 25133 24123 25191 24129
rect 25133 24089 25145 24123
rect 25179 24120 25191 24123
rect 25958 24120 25964 24132
rect 25179 24092 25964 24120
rect 25179 24089 25191 24092
rect 25133 24083 25191 24089
rect 25958 24080 25964 24092
rect 26016 24080 26022 24132
rect 17310 24052 17316 24064
rect 16500 24024 17316 24052
rect 15381 24015 15439 24021
rect 17310 24012 17316 24024
rect 17368 24012 17374 24064
rect 17678 24012 17684 24064
rect 17736 24052 17742 24064
rect 19429 24055 19487 24061
rect 19429 24052 19441 24055
rect 17736 24024 19441 24052
rect 17736 24012 17742 24024
rect 19429 24021 19441 24024
rect 19475 24021 19487 24055
rect 19429 24015 19487 24021
rect 22465 24055 22523 24061
rect 22465 24021 22477 24055
rect 22511 24052 22523 24055
rect 22830 24052 22836 24064
rect 22511 24024 22836 24052
rect 22511 24021 22523 24024
rect 22465 24015 22523 24021
rect 22830 24012 22836 24024
rect 22888 24052 22894 24064
rect 23198 24052 23204 24064
rect 22888 24024 23204 24052
rect 22888 24012 22894 24024
rect 23198 24012 23204 24024
rect 23256 24012 23262 24064
rect 28184 24052 28212 24160
rect 29362 24148 29368 24160
rect 29420 24148 29426 24200
rect 29564 24188 29592 24228
rect 29641 24225 29653 24259
rect 29687 24225 29699 24259
rect 29641 24219 29699 24225
rect 29825 24259 29883 24265
rect 29825 24225 29837 24259
rect 29871 24256 29883 24259
rect 30466 24256 30472 24268
rect 29871 24228 30328 24256
rect 30427 24228 30472 24256
rect 29871 24225 29883 24228
rect 29825 24219 29883 24225
rect 29914 24188 29920 24200
rect 29564 24160 29920 24188
rect 29914 24148 29920 24160
rect 29972 24148 29978 24200
rect 30300 24120 30328 24228
rect 30466 24216 30472 24228
rect 30524 24216 30530 24268
rect 30650 24216 30656 24268
rect 30708 24256 30714 24268
rect 30745 24259 30803 24265
rect 30745 24256 30757 24259
rect 30708 24228 30757 24256
rect 30708 24216 30714 24228
rect 30745 24225 30757 24228
rect 30791 24225 30803 24259
rect 32490 24256 32496 24268
rect 32451 24228 32496 24256
rect 30745 24219 30803 24225
rect 32490 24216 32496 24228
rect 32548 24216 32554 24268
rect 33045 24259 33103 24265
rect 33045 24225 33057 24259
rect 33091 24225 33103 24259
rect 33318 24256 33324 24268
rect 33279 24228 33324 24256
rect 33045 24219 33103 24225
rect 32582 24188 32588 24200
rect 32543 24160 32588 24188
rect 32582 24148 32588 24160
rect 32640 24148 32646 24200
rect 33060 24188 33088 24219
rect 33318 24216 33324 24228
rect 33376 24216 33382 24268
rect 33594 24256 33600 24268
rect 33555 24228 33600 24256
rect 33594 24216 33600 24228
rect 33652 24216 33658 24268
rect 34072 24265 34100 24296
rect 34882 24284 34888 24296
rect 34940 24284 34946 24336
rect 36078 24284 36084 24336
rect 36136 24324 36142 24336
rect 38194 24324 38200 24336
rect 36136 24296 38200 24324
rect 36136 24284 36142 24296
rect 38194 24284 38200 24296
rect 38252 24324 38258 24336
rect 38252 24296 38608 24324
rect 38252 24284 38258 24296
rect 34057 24259 34115 24265
rect 34057 24225 34069 24259
rect 34103 24225 34115 24259
rect 35066 24256 35072 24268
rect 35027 24228 35072 24256
rect 34057 24219 34115 24225
rect 35066 24216 35072 24228
rect 35124 24216 35130 24268
rect 35342 24216 35348 24268
rect 35400 24216 35406 24268
rect 35526 24216 35532 24268
rect 35584 24256 35590 24268
rect 36909 24259 36967 24265
rect 36909 24256 36921 24259
rect 35584 24228 36921 24256
rect 35584 24216 35590 24228
rect 36909 24225 36921 24228
rect 36955 24225 36967 24259
rect 36909 24219 36967 24225
rect 36998 24216 37004 24268
rect 37056 24216 37062 24268
rect 37826 24256 37832 24268
rect 37787 24228 37832 24256
rect 37826 24216 37832 24228
rect 37884 24216 37890 24268
rect 38286 24256 38292 24268
rect 38247 24228 38292 24256
rect 38286 24216 38292 24228
rect 38344 24216 38350 24268
rect 38580 24265 38608 24296
rect 38565 24259 38623 24265
rect 38565 24225 38577 24259
rect 38611 24225 38623 24259
rect 38565 24219 38623 24225
rect 34514 24188 34520 24200
rect 33060 24160 34520 24188
rect 34514 24148 34520 24160
rect 34572 24148 34578 24200
rect 34793 24191 34851 24197
rect 34793 24157 34805 24191
rect 34839 24188 34851 24191
rect 35360 24188 35388 24216
rect 37016 24188 37044 24216
rect 34839 24160 37044 24188
rect 34839 24157 34851 24160
rect 34793 24151 34851 24157
rect 33594 24120 33600 24132
rect 30300 24092 33600 24120
rect 33594 24080 33600 24092
rect 33652 24080 33658 24132
rect 34808 24120 34836 24151
rect 37001 24123 37059 24129
rect 37001 24120 37013 24123
rect 33704 24092 34836 24120
rect 35728 24092 37013 24120
rect 30834 24052 30840 24064
rect 28184 24024 30840 24052
rect 30834 24012 30840 24024
rect 30892 24012 30898 24064
rect 31018 24012 31024 24064
rect 31076 24052 31082 24064
rect 32214 24052 32220 24064
rect 31076 24024 32220 24052
rect 31076 24012 31082 24024
rect 32214 24012 32220 24024
rect 32272 24052 32278 24064
rect 33704 24052 33732 24092
rect 32272 24024 33732 24052
rect 32272 24012 32278 24024
rect 34330 24012 34336 24064
rect 34388 24052 34394 24064
rect 35728 24052 35756 24092
rect 37001 24089 37013 24092
rect 37047 24089 37059 24123
rect 37001 24083 37059 24089
rect 36354 24052 36360 24064
rect 34388 24024 35756 24052
rect 36315 24024 36360 24052
rect 34388 24012 34394 24024
rect 36354 24012 36360 24024
rect 36412 24012 36418 24064
rect 1104 23962 39836 23984
rect 1104 23910 4246 23962
rect 4298 23910 4310 23962
rect 4362 23910 4374 23962
rect 4426 23910 4438 23962
rect 4490 23910 34966 23962
rect 35018 23910 35030 23962
rect 35082 23910 35094 23962
rect 35146 23910 35158 23962
rect 35210 23910 39836 23962
rect 1104 23888 39836 23910
rect 8202 23848 8208 23860
rect 6932 23820 8208 23848
rect 5626 23780 5632 23792
rect 5587 23752 5632 23780
rect 5626 23740 5632 23752
rect 5684 23740 5690 23792
rect 2774 23672 2780 23724
rect 2832 23712 2838 23724
rect 3418 23712 3424 23724
rect 2832 23684 2877 23712
rect 3379 23684 3424 23712
rect 2832 23672 2838 23684
rect 3418 23672 3424 23684
rect 3476 23672 3482 23724
rect 3694 23712 3700 23724
rect 3655 23684 3700 23712
rect 3694 23672 3700 23684
rect 3752 23672 3758 23724
rect 6932 23721 6960 23820
rect 8202 23808 8208 23820
rect 8260 23808 8266 23860
rect 14001 23851 14059 23857
rect 14001 23848 14013 23851
rect 11900 23820 14013 23848
rect 8481 23783 8539 23789
rect 8481 23780 8493 23783
rect 7484 23752 8493 23780
rect 7484 23721 7512 23752
rect 8481 23749 8493 23752
rect 8527 23749 8539 23783
rect 11238 23780 11244 23792
rect 8481 23743 8539 23749
rect 8588 23752 11244 23780
rect 6917 23715 6975 23721
rect 6917 23681 6929 23715
rect 6963 23681 6975 23715
rect 6917 23675 6975 23681
rect 7469 23715 7527 23721
rect 7469 23681 7481 23715
rect 7515 23681 7527 23715
rect 8588 23712 8616 23752
rect 11238 23740 11244 23752
rect 11296 23740 11302 23792
rect 11422 23740 11428 23792
rect 11480 23740 11486 23792
rect 10502 23712 10508 23724
rect 7469 23675 7527 23681
rect 7852 23684 8616 23712
rect 9600 23684 10508 23712
rect 2038 23644 2044 23656
rect 1999 23616 2044 23644
rect 2038 23604 2044 23616
rect 2096 23604 2102 23656
rect 2406 23644 2412 23656
rect 2367 23616 2412 23644
rect 2406 23604 2412 23616
rect 2464 23604 2470 23656
rect 2685 23647 2743 23653
rect 2685 23613 2697 23647
rect 2731 23613 2743 23647
rect 5718 23644 5724 23656
rect 5679 23616 5724 23644
rect 2685 23607 2743 23613
rect 2700 23508 2728 23607
rect 5718 23604 5724 23616
rect 5776 23604 5782 23656
rect 6273 23647 6331 23653
rect 6273 23613 6285 23647
rect 6319 23644 6331 23647
rect 6822 23644 6828 23656
rect 6319 23616 6828 23644
rect 6319 23613 6331 23616
rect 6273 23607 6331 23613
rect 6822 23604 6828 23616
rect 6880 23604 6886 23656
rect 7745 23647 7803 23653
rect 7745 23613 7757 23647
rect 7791 23644 7803 23647
rect 7852 23644 7880 23684
rect 7791 23616 7880 23644
rect 7929 23647 7987 23653
rect 7791 23613 7803 23616
rect 7745 23607 7803 23613
rect 7929 23613 7941 23647
rect 7975 23644 7987 23647
rect 8386 23644 8392 23656
rect 7975 23616 8156 23644
rect 8347 23616 8392 23644
rect 7975 23613 7987 23616
rect 7929 23607 7987 23613
rect 4706 23508 4712 23520
rect 2700 23480 4712 23508
rect 4706 23468 4712 23480
rect 4764 23468 4770 23520
rect 4982 23508 4988 23520
rect 4943 23480 4988 23508
rect 4982 23468 4988 23480
rect 5040 23468 5046 23520
rect 8128 23508 8156 23616
rect 8386 23604 8392 23616
rect 8444 23604 8450 23656
rect 9600 23653 9628 23684
rect 10502 23672 10508 23684
rect 10560 23672 10566 23724
rect 10873 23715 10931 23721
rect 10873 23681 10885 23715
rect 10919 23712 10931 23715
rect 11440 23712 11468 23740
rect 10919 23684 11468 23712
rect 10919 23681 10931 23684
rect 10873 23675 10931 23681
rect 11790 23672 11796 23724
rect 11848 23712 11854 23724
rect 11900 23721 11928 23820
rect 14001 23817 14013 23820
rect 14047 23848 14059 23851
rect 14734 23848 14740 23860
rect 14047 23820 14740 23848
rect 14047 23817 14059 23820
rect 14001 23811 14059 23817
rect 14734 23808 14740 23820
rect 14792 23808 14798 23860
rect 15654 23808 15660 23860
rect 15712 23848 15718 23860
rect 17129 23851 17187 23857
rect 17129 23848 17141 23851
rect 15712 23820 17141 23848
rect 15712 23808 15718 23820
rect 17129 23817 17141 23820
rect 17175 23817 17187 23851
rect 17129 23811 17187 23817
rect 17310 23808 17316 23860
rect 17368 23848 17374 23860
rect 19334 23848 19340 23860
rect 17368 23820 19340 23848
rect 17368 23808 17374 23820
rect 19334 23808 19340 23820
rect 19392 23808 19398 23860
rect 22922 23848 22928 23860
rect 22883 23820 22928 23848
rect 22922 23808 22928 23820
rect 22980 23808 22986 23860
rect 23566 23808 23572 23860
rect 23624 23848 23630 23860
rect 24121 23851 24179 23857
rect 24121 23848 24133 23851
rect 23624 23820 24133 23848
rect 23624 23808 23630 23820
rect 24121 23817 24133 23820
rect 24167 23817 24179 23851
rect 24121 23811 24179 23817
rect 30101 23851 30159 23857
rect 30101 23817 30113 23851
rect 30147 23848 30159 23851
rect 35897 23851 35955 23857
rect 30147 23820 34192 23848
rect 30147 23817 30159 23820
rect 30101 23811 30159 23817
rect 15565 23783 15623 23789
rect 15565 23749 15577 23783
rect 15611 23749 15623 23783
rect 15565 23743 15623 23749
rect 17865 23783 17923 23789
rect 17865 23749 17877 23783
rect 17911 23780 17923 23783
rect 18230 23780 18236 23792
rect 17911 23752 18236 23780
rect 17911 23749 17923 23752
rect 17865 23743 17923 23749
rect 11885 23715 11943 23721
rect 11885 23712 11897 23715
rect 11848 23684 11897 23712
rect 11848 23672 11854 23684
rect 11885 23681 11897 23684
rect 11931 23681 11943 23715
rect 15580 23712 15608 23743
rect 18230 23740 18236 23752
rect 18288 23740 18294 23792
rect 18325 23783 18383 23789
rect 18325 23749 18337 23783
rect 18371 23780 18383 23783
rect 19978 23780 19984 23792
rect 18371 23752 19984 23780
rect 18371 23749 18383 23752
rect 18325 23743 18383 23749
rect 19978 23740 19984 23752
rect 20036 23740 20042 23792
rect 21634 23740 21640 23792
rect 21692 23780 21698 23792
rect 21818 23780 21824 23792
rect 21692 23752 21824 23780
rect 21692 23740 21698 23752
rect 21818 23740 21824 23752
rect 21876 23740 21882 23792
rect 25590 23740 25596 23792
rect 25648 23780 25654 23792
rect 25961 23783 26019 23789
rect 25961 23780 25973 23783
rect 25648 23752 25973 23780
rect 25648 23740 25654 23752
rect 25961 23749 25973 23752
rect 26007 23749 26019 23783
rect 25961 23743 26019 23749
rect 30650 23740 30656 23792
rect 30708 23740 30714 23792
rect 22281 23715 22339 23721
rect 15580 23684 21588 23712
rect 11885 23675 11943 23681
rect 8849 23647 8907 23653
rect 8849 23644 8861 23647
rect 8772 23616 8861 23644
rect 8202 23536 8208 23588
rect 8260 23576 8266 23588
rect 8478 23576 8484 23588
rect 8260 23548 8484 23576
rect 8260 23536 8266 23548
rect 8478 23536 8484 23548
rect 8536 23536 8542 23588
rect 8772 23508 8800 23616
rect 8849 23613 8861 23616
rect 8895 23613 8907 23647
rect 8849 23607 8907 23613
rect 9585 23647 9643 23653
rect 9585 23613 9597 23647
rect 9631 23613 9643 23647
rect 9858 23644 9864 23656
rect 9819 23616 9864 23644
rect 9585 23607 9643 23613
rect 9858 23604 9864 23616
rect 9916 23604 9922 23656
rect 10318 23644 10324 23656
rect 10279 23616 10324 23644
rect 10318 23604 10324 23616
rect 10376 23604 10382 23656
rect 10778 23604 10784 23656
rect 10836 23644 10842 23656
rect 11425 23647 11483 23653
rect 11425 23644 11437 23647
rect 10836 23616 11437 23644
rect 10836 23604 10842 23616
rect 11425 23613 11437 23616
rect 11471 23613 11483 23647
rect 11698 23644 11704 23656
rect 11659 23616 11704 23644
rect 11425 23607 11483 23613
rect 11698 23604 11704 23616
rect 11756 23604 11762 23656
rect 12437 23647 12495 23653
rect 12437 23613 12449 23647
rect 12483 23613 12495 23647
rect 12710 23644 12716 23656
rect 12671 23616 12716 23644
rect 12437 23607 12495 23613
rect 9766 23536 9772 23588
rect 9824 23576 9830 23588
rect 12452 23576 12480 23607
rect 12710 23604 12716 23616
rect 12768 23604 12774 23656
rect 14550 23644 14556 23656
rect 14511 23616 14556 23644
rect 14550 23604 14556 23616
rect 14608 23604 14614 23656
rect 15286 23644 15292 23656
rect 15247 23616 15292 23644
rect 15286 23604 15292 23616
rect 15344 23604 15350 23656
rect 16025 23647 16083 23653
rect 16025 23613 16037 23647
rect 16071 23613 16083 23647
rect 16025 23607 16083 23613
rect 9824 23548 12480 23576
rect 16040 23576 16068 23607
rect 16114 23604 16120 23656
rect 16172 23644 16178 23656
rect 16945 23647 17003 23653
rect 16172 23616 16217 23644
rect 16172 23604 16178 23616
rect 16945 23613 16957 23647
rect 16991 23644 17003 23647
rect 17865 23647 17923 23653
rect 17865 23644 17877 23647
rect 16991 23616 17877 23644
rect 16991 23613 17003 23616
rect 16945 23607 17003 23613
rect 17865 23613 17877 23616
rect 17911 23613 17923 23647
rect 18046 23644 18052 23656
rect 18007 23616 18052 23644
rect 17865 23607 17923 23613
rect 18046 23604 18052 23616
rect 18104 23604 18110 23656
rect 18601 23647 18659 23653
rect 18601 23613 18613 23647
rect 18647 23613 18659 23647
rect 18874 23644 18880 23656
rect 18835 23616 18880 23644
rect 18601 23607 18659 23613
rect 16574 23576 16580 23588
rect 16040 23548 16580 23576
rect 9824 23536 9830 23548
rect 16574 23536 16580 23548
rect 16632 23536 16638 23588
rect 17494 23536 17500 23588
rect 17552 23576 17558 23588
rect 18616 23576 18644 23607
rect 18874 23604 18880 23616
rect 18932 23604 18938 23656
rect 19889 23647 19947 23653
rect 19889 23613 19901 23647
rect 19935 23613 19947 23647
rect 19889 23607 19947 23613
rect 17552 23548 18644 23576
rect 19904 23576 19932 23607
rect 20070 23604 20076 23656
rect 20128 23644 20134 23656
rect 20441 23647 20499 23653
rect 20441 23644 20453 23647
rect 20128 23616 20453 23644
rect 20128 23604 20134 23616
rect 20441 23613 20453 23616
rect 20487 23613 20499 23647
rect 20441 23607 20499 23613
rect 20625 23647 20683 23653
rect 20625 23613 20637 23647
rect 20671 23644 20683 23647
rect 20714 23644 20720 23656
rect 20671 23616 20720 23644
rect 20671 23613 20683 23616
rect 20625 23607 20683 23613
rect 20714 23604 20720 23616
rect 20772 23604 20778 23656
rect 21082 23604 21088 23656
rect 21140 23644 21146 23656
rect 21560 23653 21588 23684
rect 22281 23681 22293 23715
rect 22327 23712 22339 23715
rect 23382 23712 23388 23724
rect 22327 23684 23388 23712
rect 22327 23681 22339 23684
rect 22281 23675 22339 23681
rect 23382 23672 23388 23684
rect 23440 23672 23446 23724
rect 25314 23712 25320 23724
rect 25275 23684 25320 23712
rect 25314 23672 25320 23684
rect 25372 23672 25378 23724
rect 30558 23712 30564 23724
rect 25516 23684 30564 23712
rect 21177 23647 21235 23653
rect 21177 23644 21189 23647
rect 21140 23616 21189 23644
rect 21140 23604 21146 23616
rect 21177 23613 21189 23616
rect 21223 23613 21235 23647
rect 21177 23607 21235 23613
rect 21545 23647 21603 23653
rect 21545 23613 21557 23647
rect 21591 23613 21603 23647
rect 21545 23607 21603 23613
rect 21634 23604 21640 23656
rect 21692 23644 21698 23656
rect 22005 23647 22063 23653
rect 22005 23644 22017 23647
rect 21692 23616 22017 23644
rect 21692 23604 21698 23616
rect 22005 23613 22017 23616
rect 22051 23613 22063 23647
rect 22005 23607 22063 23613
rect 22741 23647 22799 23653
rect 22741 23613 22753 23647
rect 22787 23644 22799 23647
rect 23014 23644 23020 23656
rect 22787 23616 23020 23644
rect 22787 23613 22799 23616
rect 22741 23607 22799 23613
rect 23014 23604 23020 23616
rect 23072 23604 23078 23656
rect 23842 23644 23848 23656
rect 23803 23616 23848 23644
rect 23842 23604 23848 23616
rect 23900 23604 23906 23656
rect 23937 23647 23995 23653
rect 23937 23613 23949 23647
rect 23983 23613 23995 23647
rect 23937 23607 23995 23613
rect 20990 23576 20996 23588
rect 19904 23548 20996 23576
rect 17552 23536 17558 23548
rect 20990 23536 20996 23548
rect 21048 23536 21054 23588
rect 23952 23576 23980 23607
rect 24854 23604 24860 23656
rect 24912 23644 24918 23656
rect 25516 23644 25544 23684
rect 30558 23672 30564 23684
rect 30616 23672 30622 23724
rect 30668 23712 30696 23740
rect 32033 23715 32091 23721
rect 32033 23712 32045 23715
rect 30668 23684 32045 23712
rect 32033 23681 32045 23684
rect 32079 23681 32091 23715
rect 32033 23675 32091 23681
rect 25682 23644 25688 23656
rect 24912 23616 25544 23644
rect 25643 23616 25688 23644
rect 24912 23604 24918 23616
rect 25682 23604 25688 23616
rect 25740 23604 25746 23656
rect 25958 23644 25964 23656
rect 25919 23616 25964 23644
rect 25958 23604 25964 23616
rect 26016 23604 26022 23656
rect 26697 23647 26755 23653
rect 26697 23613 26709 23647
rect 26743 23613 26755 23647
rect 26970 23644 26976 23656
rect 26931 23616 26976 23644
rect 26697 23607 26755 23613
rect 26510 23576 26516 23588
rect 23952 23548 26516 23576
rect 26510 23536 26516 23548
rect 26568 23536 26574 23588
rect 10318 23508 10324 23520
rect 8128 23480 10324 23508
rect 10318 23468 10324 23480
rect 10376 23468 10382 23520
rect 14458 23468 14464 23520
rect 14516 23508 14522 23520
rect 14737 23511 14795 23517
rect 14737 23508 14749 23511
rect 14516 23480 14749 23508
rect 14516 23468 14522 23480
rect 14737 23477 14749 23480
rect 14783 23477 14795 23511
rect 14737 23471 14795 23477
rect 18230 23468 18236 23520
rect 18288 23508 18294 23520
rect 19705 23511 19763 23517
rect 19705 23508 19717 23511
rect 18288 23480 19717 23508
rect 18288 23468 18294 23480
rect 19705 23477 19717 23480
rect 19751 23477 19763 23511
rect 19705 23471 19763 23477
rect 19978 23468 19984 23520
rect 20036 23508 20042 23520
rect 20162 23508 20168 23520
rect 20036 23480 20168 23508
rect 20036 23468 20042 23480
rect 20162 23468 20168 23480
rect 20220 23468 20226 23520
rect 20714 23468 20720 23520
rect 20772 23508 20778 23520
rect 21358 23508 21364 23520
rect 20772 23480 21364 23508
rect 20772 23468 20778 23480
rect 21358 23468 21364 23480
rect 21416 23508 21422 23520
rect 21726 23508 21732 23520
rect 21416 23480 21732 23508
rect 21416 23468 21422 23480
rect 21726 23468 21732 23480
rect 21784 23468 21790 23520
rect 25130 23468 25136 23520
rect 25188 23508 25194 23520
rect 26712 23508 26740 23607
rect 26970 23604 26976 23616
rect 27028 23604 27034 23656
rect 29273 23647 29331 23653
rect 29273 23613 29285 23647
rect 29319 23644 29331 23647
rect 30009 23647 30067 23653
rect 30009 23644 30021 23647
rect 29319 23616 30021 23644
rect 29319 23613 29331 23616
rect 29273 23607 29331 23613
rect 30009 23613 30021 23616
rect 30055 23644 30067 23647
rect 30466 23644 30472 23656
rect 30055 23616 30472 23644
rect 30055 23613 30067 23616
rect 30009 23607 30067 23613
rect 30466 23604 30472 23616
rect 30524 23604 30530 23656
rect 30653 23647 30711 23653
rect 30653 23613 30665 23647
rect 30699 23613 30711 23647
rect 30653 23607 30711 23613
rect 30929 23647 30987 23653
rect 30929 23613 30941 23647
rect 30975 23644 30987 23647
rect 32950 23644 32956 23656
rect 30975 23616 32956 23644
rect 30975 23613 30987 23616
rect 30929 23607 30987 23613
rect 28350 23576 28356 23588
rect 28311 23548 28356 23576
rect 28350 23536 28356 23548
rect 28408 23536 28414 23588
rect 29638 23536 29644 23588
rect 29696 23576 29702 23588
rect 30668 23576 30696 23607
rect 32950 23604 32956 23616
rect 33008 23604 33014 23656
rect 33318 23644 33324 23656
rect 33279 23616 33324 23644
rect 33318 23604 33324 23616
rect 33376 23604 33382 23656
rect 33778 23644 33784 23656
rect 33739 23616 33784 23644
rect 33778 23604 33784 23616
rect 33836 23604 33842 23656
rect 34164 23653 34192 23820
rect 35897 23817 35909 23851
rect 35943 23848 35955 23851
rect 37366 23848 37372 23860
rect 35943 23820 37372 23848
rect 35943 23817 35955 23820
rect 35897 23811 35955 23817
rect 37366 23808 37372 23820
rect 37424 23808 37430 23860
rect 34422 23740 34428 23792
rect 34480 23780 34486 23792
rect 35158 23780 35164 23792
rect 34480 23752 35164 23780
rect 34480 23740 34486 23752
rect 35158 23740 35164 23752
rect 35216 23740 35222 23792
rect 36998 23712 37004 23724
rect 36959 23684 37004 23712
rect 36998 23672 37004 23684
rect 37056 23672 37062 23724
rect 37274 23712 37280 23724
rect 37235 23684 37280 23712
rect 37274 23672 37280 23684
rect 37332 23672 37338 23724
rect 34149 23647 34207 23653
rect 34149 23613 34161 23647
rect 34195 23644 34207 23647
rect 34885 23647 34943 23653
rect 34195 23616 34376 23644
rect 34195 23613 34207 23616
rect 34149 23607 34207 23613
rect 34238 23576 34244 23588
rect 29696 23548 30696 23576
rect 34199 23548 34244 23576
rect 29696 23536 29702 23548
rect 25188 23480 26740 23508
rect 25188 23468 25194 23480
rect 27614 23468 27620 23520
rect 27672 23508 27678 23520
rect 29457 23511 29515 23517
rect 29457 23508 29469 23511
rect 27672 23480 29469 23508
rect 27672 23468 27678 23480
rect 29457 23477 29469 23480
rect 29503 23477 29515 23511
rect 30668 23508 30696 23548
rect 34238 23536 34244 23548
rect 34296 23536 34302 23588
rect 34348 23576 34376 23616
rect 34885 23613 34897 23647
rect 34931 23644 34943 23647
rect 35526 23644 35532 23656
rect 34931 23616 35532 23644
rect 34931 23613 34943 23616
rect 34885 23607 34943 23613
rect 35526 23604 35532 23616
rect 35584 23604 35590 23656
rect 36078 23644 36084 23656
rect 36039 23616 36084 23644
rect 36078 23604 36084 23616
rect 36136 23604 36142 23656
rect 36262 23604 36268 23656
rect 36320 23644 36326 23656
rect 36357 23647 36415 23653
rect 36357 23644 36369 23647
rect 36320 23616 36369 23644
rect 36320 23604 36326 23616
rect 36357 23613 36369 23616
rect 36403 23644 36415 23647
rect 36722 23644 36728 23656
rect 36403 23616 36728 23644
rect 36403 23613 36415 23616
rect 36357 23607 36415 23613
rect 36722 23604 36728 23616
rect 36780 23604 36786 23656
rect 34514 23576 34520 23588
rect 34348 23548 34520 23576
rect 34514 23536 34520 23548
rect 34572 23576 34578 23588
rect 35618 23576 35624 23588
rect 34572 23548 35624 23576
rect 34572 23536 34578 23548
rect 35618 23536 35624 23548
rect 35676 23536 35682 23588
rect 31018 23508 31024 23520
rect 30668 23480 31024 23508
rect 29457 23471 29515 23477
rect 31018 23468 31024 23480
rect 31076 23468 31082 23520
rect 31386 23468 31392 23520
rect 31444 23508 31450 23520
rect 33318 23508 33324 23520
rect 31444 23480 33324 23508
rect 31444 23468 31450 23480
rect 33318 23468 33324 23480
rect 33376 23468 33382 23520
rect 33410 23468 33416 23520
rect 33468 23508 33474 23520
rect 35069 23511 35127 23517
rect 35069 23508 35081 23511
rect 33468 23480 35081 23508
rect 33468 23468 33474 23480
rect 35069 23477 35081 23480
rect 35115 23477 35127 23511
rect 35069 23471 35127 23477
rect 35434 23468 35440 23520
rect 35492 23508 35498 23520
rect 38381 23511 38439 23517
rect 38381 23508 38393 23511
rect 35492 23480 38393 23508
rect 35492 23468 35498 23480
rect 38381 23477 38393 23480
rect 38427 23477 38439 23511
rect 38381 23471 38439 23477
rect 1104 23418 39836 23440
rect 1104 23366 19606 23418
rect 19658 23366 19670 23418
rect 19722 23366 19734 23418
rect 19786 23366 19798 23418
rect 19850 23366 39836 23418
rect 1104 23344 39836 23366
rect 5534 23264 5540 23316
rect 5592 23304 5598 23316
rect 10778 23304 10784 23316
rect 5592 23276 7052 23304
rect 5592 23264 5598 23276
rect 5994 23236 6000 23248
rect 5828 23208 6000 23236
rect 4890 23168 4896 23180
rect 4851 23140 4896 23168
rect 4890 23128 4896 23140
rect 4948 23128 4954 23180
rect 5828 23177 5856 23208
rect 5994 23196 6000 23208
rect 6052 23196 6058 23248
rect 7024 23245 7052 23276
rect 7576 23276 10784 23304
rect 7009 23239 7067 23245
rect 7009 23205 7021 23239
rect 7055 23205 7067 23239
rect 7009 23199 7067 23205
rect 5353 23171 5411 23177
rect 5353 23137 5365 23171
rect 5399 23137 5411 23171
rect 5353 23131 5411 23137
rect 5813 23171 5871 23177
rect 5813 23137 5825 23171
rect 5859 23137 5871 23171
rect 6086 23168 6092 23180
rect 6047 23140 6092 23168
rect 5813 23131 5871 23137
rect 1394 23100 1400 23112
rect 1355 23072 1400 23100
rect 1394 23060 1400 23072
rect 1452 23060 1458 23112
rect 1673 23103 1731 23109
rect 1673 23069 1685 23103
rect 1719 23100 1731 23103
rect 1762 23100 1768 23112
rect 1719 23072 1768 23100
rect 1719 23069 1731 23072
rect 1673 23063 1731 23069
rect 1762 23060 1768 23072
rect 1820 23060 1826 23112
rect 3326 23060 3332 23112
rect 3384 23100 3390 23112
rect 5368 23100 5396 23131
rect 6086 23128 6092 23140
rect 6144 23128 6150 23180
rect 6178 23128 6184 23180
rect 6236 23168 6242 23180
rect 7576 23177 7604 23276
rect 10778 23264 10784 23276
rect 10836 23264 10842 23316
rect 13998 23264 14004 23316
rect 14056 23304 14062 23316
rect 16114 23304 16120 23316
rect 14056 23276 16120 23304
rect 14056 23264 14062 23276
rect 16114 23264 16120 23276
rect 16172 23264 16178 23316
rect 20990 23264 20996 23316
rect 21048 23304 21054 23316
rect 23014 23304 23020 23316
rect 21048 23276 23020 23304
rect 21048 23264 21054 23276
rect 23014 23264 23020 23276
rect 23072 23264 23078 23316
rect 23198 23264 23204 23316
rect 23256 23304 23262 23316
rect 23256 23276 27108 23304
rect 23256 23264 23262 23276
rect 12618 23236 12624 23248
rect 8036 23208 12624 23236
rect 6273 23171 6331 23177
rect 6273 23168 6285 23171
rect 6236 23140 6285 23168
rect 6236 23128 6242 23140
rect 6273 23137 6285 23140
rect 6319 23137 6331 23171
rect 6273 23131 6331 23137
rect 7561 23171 7619 23177
rect 7561 23137 7573 23171
rect 7607 23137 7619 23171
rect 7834 23168 7840 23180
rect 7795 23140 7840 23168
rect 7561 23131 7619 23137
rect 7834 23128 7840 23140
rect 7892 23128 7898 23180
rect 8036 23177 8064 23208
rect 12618 23196 12624 23208
rect 12676 23196 12682 23248
rect 15286 23236 15292 23248
rect 15247 23208 15292 23236
rect 15286 23196 15292 23208
rect 15344 23196 15350 23248
rect 16666 23236 16672 23248
rect 16316 23208 16672 23236
rect 8021 23171 8079 23177
rect 8021 23137 8033 23171
rect 8067 23137 8079 23171
rect 8021 23131 8079 23137
rect 8481 23171 8539 23177
rect 8481 23137 8493 23171
rect 8527 23168 8539 23171
rect 10134 23168 10140 23180
rect 8527 23140 10140 23168
rect 8527 23137 8539 23140
rect 8481 23131 8539 23137
rect 7282 23100 7288 23112
rect 3384 23072 7288 23100
rect 3384 23060 3390 23072
rect 7282 23060 7288 23072
rect 7340 23060 7346 23112
rect 4706 22992 4712 23044
rect 4764 23032 4770 23044
rect 4764 23004 4809 23032
rect 4764 22992 4770 23004
rect 4982 22992 4988 23044
rect 5040 23032 5046 23044
rect 8036 23032 8064 23131
rect 10134 23128 10140 23140
rect 10192 23128 10198 23180
rect 10318 23168 10324 23180
rect 10279 23140 10324 23168
rect 10318 23128 10324 23140
rect 10376 23128 10382 23180
rect 10870 23168 10876 23180
rect 10831 23140 10876 23168
rect 10870 23128 10876 23140
rect 10928 23128 10934 23180
rect 11238 23168 11244 23180
rect 11199 23140 11244 23168
rect 11238 23128 11244 23140
rect 11296 23128 11302 23180
rect 11701 23171 11759 23177
rect 11701 23137 11713 23171
rect 11747 23168 11759 23171
rect 11790 23168 11796 23180
rect 11747 23140 11796 23168
rect 11747 23137 11759 23140
rect 11701 23131 11759 23137
rect 11790 23128 11796 23140
rect 11848 23128 11854 23180
rect 12158 23168 12164 23180
rect 12119 23140 12164 23168
rect 12158 23128 12164 23140
rect 12216 23128 12222 23180
rect 12342 23128 12348 23180
rect 12400 23168 12406 23180
rect 12989 23171 13047 23177
rect 12400 23140 12848 23168
rect 12400 23128 12406 23140
rect 11054 23100 11060 23112
rect 11015 23072 11060 23100
rect 11054 23060 11060 23072
rect 11112 23060 11118 23112
rect 12713 23103 12771 23109
rect 12713 23069 12725 23103
rect 12759 23069 12771 23103
rect 12820 23100 12848 23140
rect 12989 23137 13001 23171
rect 13035 23168 13047 23171
rect 14461 23171 14519 23177
rect 14461 23168 14473 23171
rect 13035 23140 14473 23168
rect 13035 23137 13047 23140
rect 12989 23131 13047 23137
rect 14461 23137 14473 23140
rect 14507 23168 14519 23171
rect 14550 23168 14556 23180
rect 14507 23140 14556 23168
rect 14507 23137 14519 23140
rect 14461 23131 14519 23137
rect 14550 23128 14556 23140
rect 14608 23128 14614 23180
rect 15654 23128 15660 23180
rect 15712 23168 15718 23180
rect 15749 23171 15807 23177
rect 15749 23168 15761 23171
rect 15712 23140 15761 23168
rect 15712 23128 15718 23140
rect 15749 23137 15761 23140
rect 15795 23137 15807 23171
rect 15749 23131 15807 23137
rect 15838 23128 15844 23180
rect 15896 23168 15902 23180
rect 15933 23171 15991 23177
rect 15933 23168 15945 23171
rect 15896 23140 15945 23168
rect 15896 23128 15902 23140
rect 15933 23137 15945 23140
rect 15979 23137 15991 23171
rect 15933 23131 15991 23137
rect 16117 23171 16175 23177
rect 16117 23137 16129 23171
rect 16163 23168 16175 23171
rect 16316 23168 16344 23208
rect 16666 23196 16672 23208
rect 16724 23236 16730 23248
rect 19242 23236 19248 23248
rect 16724 23208 17080 23236
rect 16724 23196 16730 23208
rect 16163 23140 16344 23168
rect 16163 23137 16175 23140
rect 16117 23131 16175 23137
rect 16390 23128 16396 23180
rect 16448 23168 16454 23180
rect 16945 23171 17003 23177
rect 16945 23168 16957 23171
rect 16448 23140 16957 23168
rect 16448 23128 16454 23140
rect 16945 23137 16957 23140
rect 16991 23137 17003 23171
rect 16945 23131 17003 23137
rect 13173 23103 13231 23109
rect 13173 23100 13185 23103
rect 12820 23072 13185 23100
rect 12713 23063 12771 23069
rect 13173 23069 13185 23072
rect 13219 23069 13231 23103
rect 13173 23063 13231 23069
rect 13633 23103 13691 23109
rect 13633 23069 13645 23103
rect 13679 23100 13691 23103
rect 13998 23100 14004 23112
rect 13679 23072 14004 23100
rect 13679 23069 13691 23072
rect 13633 23063 13691 23069
rect 5040 23004 8064 23032
rect 12728 23032 12756 23063
rect 13998 23060 14004 23072
rect 14056 23060 14062 23112
rect 14185 23103 14243 23109
rect 14185 23069 14197 23103
rect 14231 23100 14243 23103
rect 14366 23100 14372 23112
rect 14231 23072 14372 23100
rect 14231 23069 14243 23072
rect 14185 23063 14243 23069
rect 14200 23032 14228 23063
rect 14366 23060 14372 23072
rect 14424 23060 14430 23112
rect 14645 23103 14703 23109
rect 14645 23069 14657 23103
rect 14691 23069 14703 23103
rect 14645 23063 14703 23069
rect 12728 23004 14228 23032
rect 5040 22992 5046 23004
rect 2958 22964 2964 22976
rect 2919 22936 2964 22964
rect 2958 22924 2964 22936
rect 3016 22924 3022 22976
rect 3510 22924 3516 22976
rect 3568 22964 3574 22976
rect 5000 22964 5028 22992
rect 3568 22936 5028 22964
rect 3568 22924 3574 22936
rect 7098 22924 7104 22976
rect 7156 22964 7162 22976
rect 8665 22967 8723 22973
rect 8665 22964 8677 22967
rect 7156 22936 8677 22964
rect 7156 22924 7162 22936
rect 8665 22933 8677 22936
rect 8711 22933 8723 22967
rect 8665 22927 8723 22933
rect 10870 22924 10876 22976
rect 10928 22964 10934 22976
rect 14660 22964 14688 23063
rect 17052 23032 17080 23208
rect 17144 23208 19248 23236
rect 17144 23177 17172 23208
rect 19242 23196 19248 23208
rect 19300 23196 19306 23248
rect 21634 23236 21640 23248
rect 19996 23208 21640 23236
rect 17129 23171 17187 23177
rect 17129 23137 17141 23171
rect 17175 23137 17187 23171
rect 17129 23131 17187 23137
rect 18417 23171 18475 23177
rect 18417 23137 18429 23171
rect 18463 23137 18475 23171
rect 18690 23168 18696 23180
rect 18651 23140 18696 23168
rect 18417 23131 18475 23137
rect 18049 23103 18107 23109
rect 18049 23069 18061 23103
rect 18095 23100 18107 23103
rect 18322 23100 18328 23112
rect 18095 23072 18328 23100
rect 18095 23069 18107 23072
rect 18049 23063 18107 23069
rect 18322 23060 18328 23072
rect 18380 23060 18386 23112
rect 18432 23100 18460 23131
rect 18690 23128 18696 23140
rect 18748 23128 18754 23180
rect 19996 23177 20024 23208
rect 21634 23196 21640 23208
rect 21692 23196 21698 23248
rect 22002 23196 22008 23248
rect 22060 23236 22066 23248
rect 24949 23239 25007 23245
rect 22060 23208 23152 23236
rect 22060 23196 22066 23208
rect 19889 23171 19947 23177
rect 19889 23137 19901 23171
rect 19935 23137 19947 23171
rect 19889 23131 19947 23137
rect 19981 23171 20039 23177
rect 19981 23137 19993 23171
rect 20027 23137 20039 23171
rect 19981 23131 20039 23137
rect 20257 23171 20315 23177
rect 20257 23137 20269 23171
rect 20303 23168 20315 23171
rect 20990 23168 20996 23180
rect 20303 23140 20484 23168
rect 20951 23140 20996 23168
rect 20303 23137 20315 23140
rect 20257 23131 20315 23137
rect 19904 23100 19932 23131
rect 20346 23100 20352 23112
rect 18432 23072 18828 23100
rect 19904 23072 20352 23100
rect 17313 23035 17371 23041
rect 17313 23032 17325 23035
rect 17052 23004 17325 23032
rect 17313 23001 17325 23004
rect 17359 23001 17371 23035
rect 17313 22995 17371 23001
rect 17586 22992 17592 23044
rect 17644 23032 17650 23044
rect 18693 23035 18751 23041
rect 18693 23032 18705 23035
rect 17644 23004 18705 23032
rect 17644 22992 17650 23004
rect 18693 23001 18705 23004
rect 18739 23001 18751 23035
rect 18800 23032 18828 23072
rect 20346 23060 20352 23072
rect 20404 23060 20410 23112
rect 20456 23100 20484 23140
rect 20990 23128 20996 23140
rect 21048 23128 21054 23180
rect 21821 23171 21879 23177
rect 21821 23137 21833 23171
rect 21867 23168 21879 23171
rect 22112 23168 22140 23208
rect 22922 23168 22928 23180
rect 21867 23140 22140 23168
rect 22883 23140 22928 23168
rect 21867 23137 21879 23140
rect 21821 23131 21879 23137
rect 22922 23128 22928 23140
rect 22980 23128 22986 23180
rect 23124 23177 23152 23208
rect 24949 23205 24961 23239
rect 24995 23236 25007 23239
rect 26970 23236 26976 23248
rect 24995 23208 26976 23236
rect 24995 23205 25007 23208
rect 24949 23199 25007 23205
rect 26970 23196 26976 23208
rect 27028 23196 27034 23248
rect 23109 23171 23167 23177
rect 23109 23137 23121 23171
rect 23155 23137 23167 23171
rect 23109 23131 23167 23137
rect 23477 23171 23535 23177
rect 23477 23137 23489 23171
rect 23523 23168 23535 23171
rect 23658 23168 23664 23180
rect 23523 23140 23664 23168
rect 23523 23137 23535 23140
rect 23477 23131 23535 23137
rect 23658 23128 23664 23140
rect 23716 23128 23722 23180
rect 23934 23128 23940 23180
rect 23992 23168 23998 23180
rect 24213 23171 24271 23177
rect 24213 23168 24225 23171
rect 23992 23140 24225 23168
rect 23992 23128 23998 23140
rect 24213 23137 24225 23140
rect 24259 23168 24271 23171
rect 25682 23168 25688 23180
rect 24259 23140 25688 23168
rect 24259 23137 24271 23140
rect 24213 23131 24271 23137
rect 25682 23128 25688 23140
rect 25740 23128 25746 23180
rect 25777 23171 25835 23177
rect 25777 23137 25789 23171
rect 25823 23137 25835 23171
rect 25777 23131 25835 23137
rect 25961 23171 26019 23177
rect 25961 23137 25973 23171
rect 26007 23168 26019 23171
rect 26786 23168 26792 23180
rect 26007 23140 26792 23168
rect 26007 23137 26019 23140
rect 25961 23131 26019 23137
rect 21910 23100 21916 23112
rect 20456 23072 21588 23100
rect 21871 23072 21916 23100
rect 20254 23032 20260 23044
rect 18800 23004 20260 23032
rect 18693 22995 18751 23001
rect 20254 22992 20260 23004
rect 20312 22992 20318 23044
rect 21560 23032 21588 23072
rect 21910 23060 21916 23072
rect 21968 23060 21974 23112
rect 22002 23060 22008 23112
rect 22060 23100 22066 23112
rect 22060 23072 24440 23100
rect 22060 23060 22066 23072
rect 21818 23032 21824 23044
rect 21560 23004 21824 23032
rect 21818 22992 21824 23004
rect 21876 22992 21882 23044
rect 23290 22992 23296 23044
rect 23348 23032 23354 23044
rect 24412 23041 24440 23072
rect 25038 23060 25044 23112
rect 25096 23100 25102 23112
rect 25501 23103 25559 23109
rect 25501 23100 25513 23103
rect 25096 23072 25513 23100
rect 25096 23060 25102 23072
rect 25501 23069 25513 23072
rect 25547 23100 25559 23103
rect 25547 23072 25728 23100
rect 25547 23069 25559 23072
rect 25501 23063 25559 23069
rect 23385 23035 23443 23041
rect 23385 23032 23397 23035
rect 23348 23004 23397 23032
rect 23348 22992 23354 23004
rect 23385 23001 23397 23004
rect 23431 23001 23443 23035
rect 23385 22995 23443 23001
rect 24397 23035 24455 23041
rect 24397 23001 24409 23035
rect 24443 23001 24455 23035
rect 24397 22995 24455 23001
rect 10928 22936 14688 22964
rect 10928 22924 10934 22936
rect 16022 22924 16028 22976
rect 16080 22964 16086 22976
rect 16298 22964 16304 22976
rect 16080 22936 16304 22964
rect 16080 22924 16086 22936
rect 16298 22924 16304 22936
rect 16356 22964 16362 22976
rect 16761 22967 16819 22973
rect 16761 22964 16773 22967
rect 16356 22936 16773 22964
rect 16356 22924 16362 22936
rect 16761 22933 16773 22936
rect 16807 22933 16819 22967
rect 25700 22964 25728 23072
rect 25792 23032 25820 23131
rect 26786 23128 26792 23140
rect 26844 23128 26850 23180
rect 26234 23060 26240 23112
rect 26292 23100 26298 23112
rect 27080 23109 27108 23276
rect 29362 23264 29368 23316
rect 29420 23304 29426 23316
rect 29457 23307 29515 23313
rect 29457 23304 29469 23307
rect 29420 23276 29469 23304
rect 29420 23264 29426 23276
rect 29457 23273 29469 23276
rect 29503 23273 29515 23307
rect 29457 23267 29515 23273
rect 27890 23196 27896 23248
rect 27948 23236 27954 23248
rect 28534 23236 28540 23248
rect 27948 23208 28540 23236
rect 27948 23196 27954 23208
rect 27341 23171 27399 23177
rect 27341 23137 27353 23171
rect 27387 23168 27399 23171
rect 27798 23168 27804 23180
rect 27387 23140 27804 23168
rect 27387 23137 27399 23140
rect 27341 23131 27399 23137
rect 27798 23128 27804 23140
rect 27856 23168 27862 23180
rect 28258 23168 28264 23180
rect 27856 23140 28264 23168
rect 27856 23128 27862 23140
rect 28258 23128 28264 23140
rect 28316 23128 28322 23180
rect 28368 23177 28396 23208
rect 28534 23196 28540 23208
rect 28592 23196 28598 23248
rect 33778 23236 33784 23248
rect 32324 23208 33784 23236
rect 28353 23171 28411 23177
rect 28353 23137 28365 23171
rect 28399 23137 28411 23171
rect 28353 23131 28411 23137
rect 28442 23128 28448 23180
rect 28500 23168 28506 23180
rect 28902 23168 28908 23180
rect 28500 23140 28908 23168
rect 28500 23128 28506 23140
rect 28902 23128 28908 23140
rect 28960 23168 28966 23180
rect 29181 23171 29239 23177
rect 29181 23168 29193 23171
rect 28960 23140 29193 23168
rect 28960 23128 28966 23140
rect 29181 23137 29193 23140
rect 29227 23137 29239 23171
rect 29181 23131 29239 23137
rect 29914 23128 29920 23180
rect 29972 23168 29978 23180
rect 30101 23171 30159 23177
rect 30101 23168 30113 23171
rect 29972 23140 30113 23168
rect 29972 23128 29978 23140
rect 30101 23137 30113 23140
rect 30147 23137 30159 23171
rect 30101 23131 30159 23137
rect 30650 23128 30656 23180
rect 30708 23168 30714 23180
rect 30834 23168 30840 23180
rect 30708 23140 30840 23168
rect 30708 23128 30714 23140
rect 30834 23128 30840 23140
rect 30892 23128 30898 23180
rect 32324 23177 32352 23208
rect 33778 23196 33784 23208
rect 33836 23196 33842 23248
rect 34330 23236 34336 23248
rect 34291 23208 34336 23236
rect 34330 23196 34336 23208
rect 34388 23196 34394 23248
rect 34885 23239 34943 23245
rect 34885 23205 34897 23239
rect 34931 23236 34943 23239
rect 35250 23236 35256 23248
rect 34931 23208 35256 23236
rect 34931 23205 34943 23208
rect 34885 23199 34943 23205
rect 35250 23196 35256 23208
rect 35308 23196 35314 23248
rect 38654 23236 38660 23248
rect 37200 23208 38660 23236
rect 32309 23171 32367 23177
rect 32309 23137 32321 23171
rect 32355 23137 32367 23171
rect 32490 23168 32496 23180
rect 32451 23140 32496 23168
rect 32309 23131 32367 23137
rect 32490 23128 32496 23140
rect 32548 23128 32554 23180
rect 33042 23168 33048 23180
rect 33003 23140 33048 23168
rect 33042 23128 33048 23140
rect 33100 23128 33106 23180
rect 34238 23168 34244 23180
rect 34199 23140 34244 23168
rect 34238 23128 34244 23140
rect 34296 23128 34302 23180
rect 34425 23171 34483 23177
rect 34425 23137 34437 23171
rect 34471 23168 34483 23171
rect 34606 23168 34612 23180
rect 34471 23140 34612 23168
rect 34471 23137 34483 23140
rect 34425 23131 34483 23137
rect 34606 23128 34612 23140
rect 34664 23168 34670 23180
rect 35345 23171 35403 23177
rect 35345 23168 35357 23171
rect 34664 23140 35357 23168
rect 34664 23128 34670 23140
rect 35345 23137 35357 23140
rect 35391 23137 35403 23171
rect 35526 23168 35532 23180
rect 35487 23140 35532 23168
rect 35345 23131 35403 23137
rect 26513 23103 26571 23109
rect 26513 23100 26525 23103
rect 26292 23072 26525 23100
rect 26292 23060 26298 23072
rect 26513 23069 26525 23072
rect 26559 23069 26571 23103
rect 26513 23063 26571 23069
rect 27065 23103 27123 23109
rect 27065 23069 27077 23103
rect 27111 23069 27123 23103
rect 27065 23063 27123 23069
rect 27525 23103 27583 23109
rect 27525 23069 27537 23103
rect 27571 23100 27583 23103
rect 27614 23100 27620 23112
rect 27571 23072 27620 23100
rect 27571 23069 27583 23072
rect 27525 23063 27583 23069
rect 27614 23060 27620 23072
rect 27672 23060 27678 23112
rect 29086 23100 29092 23112
rect 27816 23072 28948 23100
rect 29047 23072 29092 23100
rect 27706 23032 27712 23044
rect 25792 23004 27712 23032
rect 27706 22992 27712 23004
rect 27764 22992 27770 23044
rect 27816 22964 27844 23072
rect 28920 23032 28948 23072
rect 29086 23060 29092 23072
rect 29144 23060 29150 23112
rect 29822 23060 29828 23112
rect 29880 23100 29886 23112
rect 32950 23100 32956 23112
rect 29880 23072 31064 23100
rect 32911 23072 32956 23100
rect 29880 23060 29886 23072
rect 31036 23044 31064 23072
rect 32950 23060 32956 23072
rect 33008 23060 33014 23112
rect 35360 23100 35388 23131
rect 35526 23128 35532 23140
rect 35584 23128 35590 23180
rect 36446 23168 36452 23180
rect 36407 23140 36452 23168
rect 36446 23128 36452 23140
rect 36504 23128 36510 23180
rect 37200 23177 37228 23208
rect 38654 23196 38660 23208
rect 38712 23236 38718 23248
rect 39025 23239 39083 23245
rect 39025 23236 39037 23239
rect 38712 23208 39037 23236
rect 38712 23196 38718 23208
rect 39025 23205 39037 23208
rect 39071 23205 39083 23239
rect 39025 23199 39083 23205
rect 37185 23171 37243 23177
rect 37185 23137 37197 23171
rect 37231 23137 37243 23171
rect 37185 23131 37243 23137
rect 37737 23171 37795 23177
rect 37737 23137 37749 23171
rect 37783 23137 37795 23171
rect 38194 23168 38200 23180
rect 38155 23140 38200 23168
rect 37737 23131 37795 23137
rect 35434 23100 35440 23112
rect 35360 23072 35440 23100
rect 35434 23060 35440 23072
rect 35492 23060 35498 23112
rect 36814 23100 36820 23112
rect 36775 23072 36820 23100
rect 36814 23060 36820 23072
rect 36872 23060 36878 23112
rect 29270 23032 29276 23044
rect 28920 23004 29276 23032
rect 29270 22992 29276 23004
rect 29328 22992 29334 23044
rect 29546 22992 29552 23044
rect 29604 23032 29610 23044
rect 31018 23032 31024 23044
rect 29604 23004 30420 23032
rect 30931 23004 31024 23032
rect 29604 22992 29610 23004
rect 25700 22936 27844 22964
rect 16761 22927 16819 22933
rect 29454 22924 29460 22976
rect 29512 22964 29518 22976
rect 30006 22964 30012 22976
rect 29512 22936 30012 22964
rect 29512 22924 29518 22936
rect 30006 22924 30012 22936
rect 30064 22964 30070 22976
rect 30285 22967 30343 22973
rect 30285 22964 30297 22967
rect 30064 22936 30297 22964
rect 30064 22924 30070 22936
rect 30285 22933 30297 22936
rect 30331 22933 30343 22967
rect 30392 22964 30420 23004
rect 31018 22992 31024 23004
rect 31076 22992 31082 23044
rect 31202 22992 31208 23044
rect 31260 23032 31266 23044
rect 37752 23032 37780 23131
rect 38194 23128 38200 23140
rect 38252 23128 38258 23180
rect 38378 23128 38384 23180
rect 38436 23168 38442 23180
rect 38933 23171 38991 23177
rect 38933 23168 38945 23171
rect 38436 23140 38945 23168
rect 38436 23128 38442 23140
rect 38933 23137 38945 23140
rect 38979 23137 38991 23171
rect 38933 23131 38991 23137
rect 38473 23103 38531 23109
rect 38473 23069 38485 23103
rect 38519 23100 38531 23103
rect 38838 23100 38844 23112
rect 38519 23072 38844 23100
rect 38519 23069 38531 23072
rect 38473 23063 38531 23069
rect 38838 23060 38844 23072
rect 38896 23060 38902 23112
rect 31260 23004 37780 23032
rect 31260 22992 31266 23004
rect 31478 22964 31484 22976
rect 30392 22936 31484 22964
rect 30285 22927 30343 22933
rect 31478 22924 31484 22936
rect 31536 22924 31542 22976
rect 34606 22924 34612 22976
rect 34664 22964 34670 22976
rect 35342 22964 35348 22976
rect 34664 22936 35348 22964
rect 34664 22924 34670 22936
rect 35342 22924 35348 22936
rect 35400 22924 35406 22976
rect 35621 22967 35679 22973
rect 35621 22933 35633 22967
rect 35667 22964 35679 22967
rect 35710 22964 35716 22976
rect 35667 22936 35716 22964
rect 35667 22933 35679 22936
rect 35621 22927 35679 22933
rect 35710 22924 35716 22936
rect 35768 22924 35774 22976
rect 1104 22874 39836 22896
rect 1104 22822 4246 22874
rect 4298 22822 4310 22874
rect 4362 22822 4374 22874
rect 4426 22822 4438 22874
rect 4490 22822 34966 22874
rect 35018 22822 35030 22874
rect 35082 22822 35094 22874
rect 35146 22822 35158 22874
rect 35210 22822 39836 22874
rect 1104 22800 39836 22822
rect 1762 22760 1768 22772
rect 1723 22732 1768 22760
rect 1762 22720 1768 22732
rect 1820 22720 1826 22772
rect 7282 22760 7288 22772
rect 7195 22732 7288 22760
rect 7282 22720 7288 22732
rect 7340 22760 7346 22772
rect 11882 22760 11888 22772
rect 7340 22732 11888 22760
rect 7340 22720 7346 22732
rect 11882 22720 11888 22732
rect 11940 22720 11946 22772
rect 12529 22763 12587 22769
rect 12529 22729 12541 22763
rect 12575 22760 12587 22763
rect 12710 22760 12716 22772
rect 12575 22732 12716 22760
rect 12575 22729 12587 22732
rect 12529 22723 12587 22729
rect 12710 22720 12716 22732
rect 12768 22720 12774 22772
rect 20717 22763 20775 22769
rect 20717 22729 20729 22763
rect 20763 22760 20775 22763
rect 21174 22760 21180 22772
rect 20763 22732 21180 22760
rect 20763 22729 20775 22732
rect 20717 22723 20775 22729
rect 21174 22720 21180 22732
rect 21232 22760 21238 22772
rect 26510 22760 26516 22772
rect 21232 22732 22968 22760
rect 26471 22732 26516 22760
rect 21232 22720 21238 22732
rect 2038 22652 2044 22704
rect 2096 22692 2102 22704
rect 2501 22695 2559 22701
rect 2501 22692 2513 22695
rect 2096 22664 2513 22692
rect 2096 22652 2102 22664
rect 2501 22661 2513 22664
rect 2547 22692 2559 22695
rect 3326 22692 3332 22704
rect 2547 22664 3332 22692
rect 2547 22661 2559 22664
rect 2501 22655 2559 22661
rect 3326 22652 3332 22664
rect 3384 22652 3390 22704
rect 5994 22652 6000 22704
rect 6052 22652 6058 22704
rect 6086 22652 6092 22704
rect 6144 22692 6150 22704
rect 6181 22695 6239 22701
rect 6181 22692 6193 22695
rect 6144 22664 6193 22692
rect 6144 22652 6150 22664
rect 6181 22661 6193 22664
rect 6227 22692 6239 22695
rect 7006 22692 7012 22704
rect 6227 22664 7012 22692
rect 6227 22661 6239 22664
rect 6181 22655 6239 22661
rect 7006 22652 7012 22664
rect 7064 22652 7070 22704
rect 2774 22624 2780 22636
rect 1688 22596 2780 22624
rect 1688 22565 1716 22596
rect 2774 22584 2780 22596
rect 2832 22584 2838 22636
rect 4249 22627 4307 22633
rect 4249 22593 4261 22627
rect 4295 22624 4307 22627
rect 4614 22624 4620 22636
rect 4295 22596 4620 22624
rect 4295 22593 4307 22596
rect 4249 22587 4307 22593
rect 4614 22584 4620 22596
rect 4672 22584 4678 22636
rect 6012 22624 6040 22652
rect 6822 22624 6828 22636
rect 6012 22596 6828 22624
rect 6822 22584 6828 22596
rect 6880 22584 6886 22636
rect 1673 22559 1731 22565
rect 1673 22525 1685 22559
rect 1719 22525 1731 22559
rect 1673 22519 1731 22525
rect 2317 22559 2375 22565
rect 2317 22525 2329 22559
rect 2363 22556 2375 22559
rect 2958 22556 2964 22568
rect 2363 22528 2964 22556
rect 2363 22525 2375 22528
rect 2317 22519 2375 22525
rect 2792 22500 2820 22528
rect 2958 22516 2964 22528
rect 3016 22516 3022 22568
rect 3326 22556 3332 22568
rect 3287 22528 3332 22556
rect 3326 22516 3332 22528
rect 3384 22516 3390 22568
rect 3510 22556 3516 22568
rect 3471 22528 3516 22556
rect 3510 22516 3516 22528
rect 3568 22516 3574 22568
rect 3786 22556 3792 22568
rect 3747 22528 3792 22556
rect 3786 22516 3792 22528
rect 3844 22516 3850 22568
rect 4706 22556 4712 22568
rect 4667 22528 4712 22556
rect 4706 22516 4712 22528
rect 4764 22516 4770 22568
rect 5353 22559 5411 22565
rect 5353 22525 5365 22559
rect 5399 22556 5411 22559
rect 5626 22556 5632 22568
rect 5399 22528 5632 22556
rect 5399 22525 5411 22528
rect 5353 22519 5411 22525
rect 5626 22516 5632 22528
rect 5684 22516 5690 22568
rect 5997 22559 6055 22565
rect 5997 22525 6009 22559
rect 6043 22525 6055 22559
rect 5997 22519 6055 22525
rect 2774 22448 2780 22500
rect 2832 22448 2838 22500
rect 3528 22488 3556 22516
rect 3694 22488 3700 22500
rect 3528 22460 3700 22488
rect 3694 22448 3700 22460
rect 3752 22448 3758 22500
rect 6012 22488 6040 22519
rect 6178 22516 6184 22568
rect 6236 22556 6242 22568
rect 6236 22528 7236 22556
rect 6236 22516 6242 22528
rect 7098 22488 7104 22500
rect 6012 22460 7104 22488
rect 7098 22448 7104 22460
rect 7156 22448 7162 22500
rect 7208 22497 7236 22528
rect 7193 22491 7251 22497
rect 7193 22457 7205 22491
rect 7239 22457 7251 22491
rect 7193 22451 7251 22457
rect 4801 22423 4859 22429
rect 4801 22389 4813 22423
rect 4847 22420 4859 22423
rect 5350 22420 5356 22432
rect 4847 22392 5356 22420
rect 4847 22389 4859 22392
rect 4801 22383 4859 22389
rect 5350 22380 5356 22392
rect 5408 22380 5414 22432
rect 5445 22423 5503 22429
rect 5445 22389 5457 22423
rect 5491 22420 5503 22423
rect 6178 22420 6184 22432
rect 5491 22392 6184 22420
rect 5491 22389 5503 22392
rect 5445 22383 5503 22389
rect 6178 22380 6184 22392
rect 6236 22380 6242 22432
rect 7009 22423 7067 22429
rect 7009 22389 7021 22423
rect 7055 22420 7067 22423
rect 7300 22420 7328 22720
rect 12894 22652 12900 22704
rect 12952 22692 12958 22704
rect 13173 22695 13231 22701
rect 13173 22692 13185 22695
rect 12952 22664 13185 22692
rect 12952 22652 12958 22664
rect 13173 22661 13185 22664
rect 13219 22661 13231 22695
rect 18877 22695 18935 22701
rect 18877 22692 18889 22695
rect 13173 22655 13231 22661
rect 16500 22664 18889 22692
rect 7561 22627 7619 22633
rect 7561 22593 7573 22627
rect 7607 22624 7619 22627
rect 7834 22624 7840 22636
rect 7607 22596 7840 22624
rect 7607 22593 7619 22596
rect 7561 22587 7619 22593
rect 7834 22584 7840 22596
rect 7892 22584 7898 22636
rect 8478 22624 8484 22636
rect 8439 22596 8484 22624
rect 8478 22584 8484 22596
rect 8536 22584 8542 22636
rect 10134 22584 10140 22636
rect 10192 22624 10198 22636
rect 11701 22627 11759 22633
rect 11701 22624 11713 22627
rect 10192 22596 11713 22624
rect 10192 22584 10198 22596
rect 11701 22593 11713 22596
rect 11747 22593 11759 22627
rect 11701 22587 11759 22593
rect 13906 22584 13912 22636
rect 13964 22624 13970 22636
rect 14093 22627 14151 22633
rect 14093 22624 14105 22627
rect 13964 22596 14105 22624
rect 13964 22584 13970 22596
rect 14093 22593 14105 22596
rect 14139 22624 14151 22627
rect 14458 22624 14464 22636
rect 14139 22596 14464 22624
rect 14139 22593 14151 22596
rect 14093 22587 14151 22593
rect 14458 22584 14464 22596
rect 14516 22584 14522 22636
rect 14829 22627 14887 22633
rect 14829 22593 14841 22627
rect 14875 22624 14887 22627
rect 15286 22624 15292 22636
rect 14875 22596 15292 22624
rect 14875 22593 14887 22596
rect 14829 22587 14887 22593
rect 15286 22584 15292 22596
rect 15344 22584 15350 22636
rect 15746 22624 15752 22636
rect 15707 22596 15752 22624
rect 15746 22584 15752 22596
rect 15804 22584 15810 22636
rect 16500 22633 16528 22664
rect 18877 22661 18889 22664
rect 18923 22661 18935 22695
rect 21818 22692 21824 22704
rect 18877 22655 18935 22661
rect 21192 22664 21824 22692
rect 16485 22627 16543 22633
rect 16485 22593 16497 22627
rect 16531 22593 16543 22627
rect 17218 22624 17224 22636
rect 17179 22596 17224 22624
rect 16485 22587 16543 22593
rect 17218 22584 17224 22596
rect 17276 22584 17282 22636
rect 18233 22627 18291 22633
rect 18233 22593 18245 22627
rect 18279 22624 18291 22627
rect 18322 22624 18328 22636
rect 18279 22596 18328 22624
rect 18279 22593 18291 22596
rect 18233 22587 18291 22593
rect 18322 22584 18328 22596
rect 18380 22584 18386 22636
rect 8205 22559 8263 22565
rect 8205 22525 8217 22559
rect 8251 22525 8263 22559
rect 8205 22519 8263 22525
rect 10965 22559 11023 22565
rect 10965 22525 10977 22559
rect 11011 22556 11023 22559
rect 11790 22556 11796 22568
rect 11011 22528 11796 22556
rect 11011 22525 11023 22528
rect 10965 22519 11023 22525
rect 8220 22432 8248 22519
rect 11790 22516 11796 22528
rect 11848 22516 11854 22568
rect 12434 22516 12440 22568
rect 12492 22556 12498 22568
rect 13170 22556 13176 22568
rect 12492 22528 12537 22556
rect 13131 22528 13176 22556
rect 12492 22516 12498 22528
rect 13170 22516 13176 22528
rect 13228 22516 13234 22568
rect 13722 22556 13728 22568
rect 13683 22528 13728 22556
rect 13722 22516 13728 22528
rect 13780 22516 13786 22568
rect 15013 22559 15071 22565
rect 15013 22525 15025 22559
rect 15059 22525 15071 22559
rect 15013 22519 15071 22525
rect 9861 22491 9919 22497
rect 9861 22457 9873 22491
rect 9907 22488 9919 22491
rect 11333 22491 11391 22497
rect 9907 22460 11284 22488
rect 9907 22457 9919 22460
rect 9861 22451 9919 22457
rect 11256 22432 11284 22460
rect 11333 22457 11345 22491
rect 11379 22488 11391 22491
rect 11606 22488 11612 22500
rect 11379 22460 11612 22488
rect 11379 22457 11391 22460
rect 11333 22451 11391 22457
rect 11606 22448 11612 22460
rect 11664 22448 11670 22500
rect 14366 22448 14372 22500
rect 14424 22488 14430 22500
rect 15028 22488 15056 22519
rect 15102 22516 15108 22568
rect 15160 22556 15166 22568
rect 15473 22559 15531 22565
rect 15473 22556 15485 22559
rect 15160 22528 15485 22556
rect 15160 22516 15166 22528
rect 15473 22525 15485 22528
rect 15519 22525 15531 22559
rect 16758 22556 16764 22568
rect 16719 22528 16764 22556
rect 15473 22519 15531 22525
rect 16758 22516 16764 22528
rect 16816 22516 16822 22568
rect 16850 22516 16856 22568
rect 16908 22556 16914 22568
rect 17129 22559 17187 22565
rect 17129 22556 17141 22559
rect 16908 22528 17141 22556
rect 16908 22516 16914 22528
rect 17129 22525 17141 22528
rect 17175 22525 17187 22559
rect 18414 22556 18420 22568
rect 18375 22528 18420 22556
rect 17129 22519 17187 22525
rect 18414 22516 18420 22528
rect 18472 22516 18478 22568
rect 18877 22559 18935 22565
rect 18877 22525 18889 22559
rect 18923 22525 18935 22559
rect 18877 22519 18935 22525
rect 19797 22559 19855 22565
rect 19797 22525 19809 22559
rect 19843 22525 19855 22559
rect 19797 22519 19855 22525
rect 20533 22559 20591 22565
rect 20533 22525 20545 22559
rect 20579 22556 20591 22559
rect 21082 22556 21088 22568
rect 20579 22528 21088 22556
rect 20579 22525 20591 22528
rect 20533 22519 20591 22525
rect 14424 22460 15056 22488
rect 14424 22448 14430 22460
rect 17954 22448 17960 22500
rect 18012 22488 18018 22500
rect 18690 22488 18696 22500
rect 18012 22460 18696 22488
rect 18012 22448 18018 22460
rect 18690 22448 18696 22460
rect 18748 22488 18754 22500
rect 18892 22488 18920 22519
rect 18748 22460 18920 22488
rect 19812 22488 19840 22519
rect 21082 22516 21088 22528
rect 21140 22516 21146 22568
rect 21192 22556 21220 22664
rect 21818 22652 21824 22664
rect 21876 22652 21882 22704
rect 22940 22692 22968 22732
rect 26510 22720 26516 22732
rect 26568 22720 26574 22772
rect 28718 22720 28724 22772
rect 28776 22760 28782 22772
rect 29822 22760 29828 22772
rect 28776 22732 29828 22760
rect 28776 22720 28782 22732
rect 29822 22720 29828 22732
rect 29880 22720 29886 22772
rect 30558 22720 30564 22772
rect 30616 22760 30622 22772
rect 31389 22763 31447 22769
rect 31389 22760 31401 22763
rect 30616 22732 31401 22760
rect 30616 22720 30622 22732
rect 31389 22729 31401 22732
rect 31435 22729 31447 22763
rect 31389 22723 31447 22729
rect 36262 22720 36268 22772
rect 36320 22760 36326 22772
rect 36449 22763 36507 22769
rect 36449 22760 36461 22763
rect 36320 22732 36461 22760
rect 36320 22720 36326 22732
rect 36449 22729 36461 22732
rect 36495 22760 36507 22763
rect 37182 22760 37188 22772
rect 36495 22732 37188 22760
rect 36495 22729 36507 22732
rect 36449 22723 36507 22729
rect 37182 22720 37188 22732
rect 37240 22720 37246 22772
rect 38194 22720 38200 22772
rect 38252 22760 38258 22772
rect 38841 22763 38899 22769
rect 38841 22760 38853 22763
rect 38252 22732 38853 22760
rect 38252 22720 38258 22732
rect 38841 22729 38853 22732
rect 38887 22729 38899 22763
rect 38841 22723 38899 22729
rect 22940 22664 24348 22692
rect 21358 22624 21364 22636
rect 21319 22596 21364 22624
rect 21358 22584 21364 22596
rect 21416 22584 21422 22636
rect 23934 22624 23940 22636
rect 22940 22596 23940 22624
rect 21269 22559 21327 22565
rect 21269 22556 21281 22559
rect 21192 22528 21281 22556
rect 21269 22525 21281 22528
rect 21315 22525 21327 22559
rect 21269 22519 21327 22525
rect 21450 22516 21456 22568
rect 21508 22556 21514 22568
rect 21637 22559 21695 22565
rect 21637 22556 21649 22559
rect 21508 22528 21649 22556
rect 21508 22516 21514 22528
rect 21637 22525 21649 22528
rect 21683 22525 21695 22559
rect 21637 22519 21695 22525
rect 22281 22559 22339 22565
rect 22281 22525 22293 22559
rect 22327 22556 22339 22559
rect 22830 22556 22836 22568
rect 22327 22528 22836 22556
rect 22327 22525 22339 22528
rect 22281 22519 22339 22525
rect 22830 22516 22836 22528
rect 22888 22516 22894 22568
rect 22940 22565 22968 22596
rect 23934 22584 23940 22596
rect 23992 22584 23998 22636
rect 24026 22584 24032 22636
rect 24084 22624 24090 22636
rect 24210 22624 24216 22636
rect 24084 22596 24216 22624
rect 24084 22584 24090 22596
rect 24210 22584 24216 22596
rect 24268 22584 24274 22636
rect 24320 22624 24348 22664
rect 28184 22664 28488 22692
rect 28184 22624 28212 22664
rect 28350 22624 28356 22636
rect 24320 22596 28212 22624
rect 28311 22596 28356 22624
rect 28350 22584 28356 22596
rect 28408 22584 28414 22636
rect 28460 22624 28488 22664
rect 31018 22652 31024 22704
rect 31076 22692 31082 22704
rect 34514 22692 34520 22704
rect 31076 22664 34520 22692
rect 31076 22652 31082 22664
rect 34514 22652 34520 22664
rect 34572 22652 34578 22704
rect 32953 22627 33011 22633
rect 28460 22596 31156 22624
rect 22925 22559 22983 22565
rect 22925 22525 22937 22559
rect 22971 22525 22983 22559
rect 22925 22519 22983 22525
rect 23014 22516 23020 22568
rect 23072 22556 23078 22568
rect 23750 22556 23756 22568
rect 23072 22528 23756 22556
rect 23072 22516 23078 22528
rect 23750 22516 23756 22528
rect 23808 22516 23814 22568
rect 23842 22516 23848 22568
rect 23900 22556 23906 22568
rect 24121 22559 24179 22565
rect 24121 22556 24133 22559
rect 23900 22528 24133 22556
rect 23900 22516 23906 22528
rect 24121 22525 24133 22528
rect 24167 22556 24179 22559
rect 24670 22556 24676 22568
rect 24167 22528 24676 22556
rect 24167 22525 24179 22528
rect 24121 22519 24179 22525
rect 24670 22516 24676 22528
rect 24728 22516 24734 22568
rect 25130 22556 25136 22568
rect 25091 22528 25136 22556
rect 25130 22516 25136 22528
rect 25188 22516 25194 22568
rect 25406 22556 25412 22568
rect 25367 22528 25412 22556
rect 25406 22516 25412 22528
rect 25464 22516 25470 22568
rect 25682 22516 25688 22568
rect 25740 22556 25746 22568
rect 27890 22556 27896 22568
rect 25740 22528 26096 22556
rect 27851 22528 27896 22556
rect 25740 22516 25746 22528
rect 23566 22488 23572 22500
rect 19812 22460 23572 22488
rect 18748 22448 18754 22460
rect 23566 22448 23572 22460
rect 23624 22448 23630 22500
rect 26068 22488 26096 22528
rect 27890 22516 27896 22528
rect 27948 22516 27954 22568
rect 28445 22559 28503 22565
rect 28445 22525 28457 22559
rect 28491 22556 28503 22559
rect 28626 22556 28632 22568
rect 28491 22528 28632 22556
rect 28491 22525 28503 22528
rect 28445 22519 28503 22525
rect 28626 22516 28632 22528
rect 28684 22516 28690 22568
rect 29454 22556 29460 22568
rect 29415 22528 29460 22556
rect 29454 22516 29460 22528
rect 29512 22516 29518 22568
rect 29917 22559 29975 22565
rect 29917 22556 29929 22559
rect 29564 22528 29929 22556
rect 26068 22460 28120 22488
rect 7055 22392 7328 22420
rect 7055 22389 7067 22392
rect 7009 22383 7067 22389
rect 8202 22380 8208 22432
rect 8260 22420 8266 22432
rect 9766 22420 9772 22432
rect 8260 22392 9772 22420
rect 8260 22380 8266 22392
rect 9766 22380 9772 22392
rect 9824 22380 9830 22432
rect 11146 22420 11152 22432
rect 11107 22392 11152 22420
rect 11146 22380 11152 22392
rect 11204 22380 11210 22432
rect 11238 22380 11244 22432
rect 11296 22420 11302 22432
rect 11296 22392 11341 22420
rect 11296 22380 11302 22392
rect 19150 22380 19156 22432
rect 19208 22420 19214 22432
rect 19981 22423 20039 22429
rect 19981 22420 19993 22423
rect 19208 22392 19993 22420
rect 19208 22380 19214 22392
rect 19981 22389 19993 22392
rect 20027 22389 20039 22423
rect 19981 22383 20039 22389
rect 23017 22423 23075 22429
rect 23017 22389 23029 22423
rect 23063 22420 23075 22423
rect 23658 22420 23664 22432
rect 23063 22392 23664 22420
rect 23063 22389 23075 22392
rect 23017 22383 23075 22389
rect 23658 22380 23664 22392
rect 23716 22380 23722 22432
rect 27893 22423 27951 22429
rect 27893 22389 27905 22423
rect 27939 22420 27951 22423
rect 27982 22420 27988 22432
rect 27939 22392 27988 22420
rect 27939 22389 27951 22392
rect 27893 22383 27951 22389
rect 27982 22380 27988 22392
rect 28040 22380 28046 22432
rect 28092 22420 28120 22460
rect 28994 22448 29000 22500
rect 29052 22488 29058 22500
rect 29564 22488 29592 22528
rect 29917 22525 29929 22528
rect 29963 22525 29975 22559
rect 29917 22519 29975 22525
rect 30285 22559 30343 22565
rect 30285 22525 30297 22559
rect 30331 22525 30343 22559
rect 31128 22556 31156 22596
rect 32953 22593 32965 22627
rect 32999 22624 33011 22627
rect 33686 22624 33692 22636
rect 32999 22596 33692 22624
rect 32999 22593 33011 22596
rect 32953 22587 33011 22593
rect 33686 22584 33692 22596
rect 33744 22584 33750 22636
rect 36354 22624 36360 22636
rect 33980 22596 36360 22624
rect 31202 22556 31208 22568
rect 31128 22528 31208 22556
rect 30285 22519 30343 22525
rect 29052 22460 29592 22488
rect 29052 22448 29058 22460
rect 29822 22448 29828 22500
rect 29880 22488 29886 22500
rect 30300 22488 30328 22519
rect 31202 22516 31208 22528
rect 31260 22516 31266 22568
rect 31570 22516 31576 22568
rect 31628 22556 31634 22568
rect 32493 22559 32551 22565
rect 32493 22556 32505 22559
rect 31628 22528 32505 22556
rect 31628 22516 31634 22528
rect 32493 22525 32505 22528
rect 32539 22525 32551 22559
rect 32493 22519 32551 22525
rect 33229 22559 33287 22565
rect 33229 22525 33241 22559
rect 33275 22525 33287 22559
rect 33229 22519 33287 22525
rect 29880 22460 30328 22488
rect 33244 22488 33272 22519
rect 33318 22516 33324 22568
rect 33376 22556 33382 22568
rect 33980 22565 34008 22596
rect 36354 22584 36360 22596
rect 36412 22584 36418 22636
rect 37458 22624 37464 22636
rect 37419 22596 37464 22624
rect 37458 22584 37464 22596
rect 37516 22584 37522 22636
rect 37737 22627 37795 22633
rect 37737 22593 37749 22627
rect 37783 22624 37795 22627
rect 38746 22624 38752 22636
rect 37783 22596 38752 22624
rect 37783 22593 37795 22596
rect 37737 22587 37795 22593
rect 38746 22584 38752 22596
rect 38804 22584 38810 22636
rect 33965 22559 34023 22565
rect 33376 22528 33421 22556
rect 33376 22516 33382 22528
rect 33965 22525 33977 22559
rect 34011 22525 34023 22559
rect 33965 22519 34023 22525
rect 34606 22516 34612 22568
rect 34664 22556 34670 22568
rect 34885 22559 34943 22565
rect 34885 22556 34897 22559
rect 34664 22528 34897 22556
rect 34664 22516 34670 22528
rect 34885 22525 34897 22528
rect 34931 22525 34943 22559
rect 35158 22556 35164 22568
rect 35119 22528 35164 22556
rect 34885 22519 34943 22525
rect 35158 22516 35164 22528
rect 35216 22516 35222 22568
rect 33502 22488 33508 22500
rect 33244 22460 33508 22488
rect 29880 22448 29886 22460
rect 33502 22448 33508 22460
rect 33560 22448 33566 22500
rect 29546 22420 29552 22432
rect 28092 22392 29552 22420
rect 29546 22380 29552 22392
rect 29604 22380 29610 22432
rect 29733 22423 29791 22429
rect 29733 22389 29745 22423
rect 29779 22420 29791 22423
rect 30006 22420 30012 22432
rect 29779 22392 30012 22420
rect 29779 22389 29791 22392
rect 29733 22383 29791 22389
rect 30006 22380 30012 22392
rect 30064 22380 30070 22432
rect 30926 22380 30932 22432
rect 30984 22420 30990 22432
rect 36446 22420 36452 22432
rect 30984 22392 36452 22420
rect 30984 22380 30990 22392
rect 36446 22380 36452 22392
rect 36504 22420 36510 22432
rect 38838 22420 38844 22432
rect 36504 22392 38844 22420
rect 36504 22380 36510 22392
rect 38838 22380 38844 22392
rect 38896 22380 38902 22432
rect 1104 22330 39836 22352
rect 1104 22278 19606 22330
rect 19658 22278 19670 22330
rect 19722 22278 19734 22330
rect 19786 22278 19798 22330
rect 19850 22278 39836 22330
rect 1104 22256 39836 22278
rect 4890 22176 4896 22228
rect 4948 22216 4954 22228
rect 7190 22216 7196 22228
rect 4948 22188 7196 22216
rect 4948 22176 4954 22188
rect 7190 22176 7196 22188
rect 7248 22216 7254 22228
rect 7374 22216 7380 22228
rect 7248 22188 7380 22216
rect 7248 22176 7254 22188
rect 7374 22176 7380 22188
rect 7432 22176 7438 22228
rect 8570 22216 8576 22228
rect 8496 22188 8576 22216
rect 2608 22120 2912 22148
rect 1486 22080 1492 22092
rect 1447 22052 1492 22080
rect 1486 22040 1492 22052
rect 1544 22040 1550 22092
rect 2133 22083 2191 22089
rect 2133 22049 2145 22083
rect 2179 22080 2191 22083
rect 2608 22080 2636 22120
rect 2179 22052 2636 22080
rect 2179 22049 2191 22052
rect 2133 22043 2191 22049
rect 2884 22012 2912 22120
rect 3436 22120 3832 22148
rect 2958 22040 2964 22092
rect 3016 22080 3022 22092
rect 3016 22052 3061 22080
rect 3016 22040 3022 22052
rect 3436 22012 3464 22120
rect 3513 22083 3571 22089
rect 3513 22049 3525 22083
rect 3559 22080 3571 22083
rect 3694 22080 3700 22092
rect 3559 22052 3700 22080
rect 3559 22049 3571 22052
rect 3513 22043 3571 22049
rect 3694 22040 3700 22052
rect 3752 22040 3758 22092
rect 2884 21984 3464 22012
rect 3804 22012 3832 22120
rect 4062 22080 4068 22092
rect 4023 22052 4068 22080
rect 4062 22040 4068 22052
rect 4120 22040 4126 22092
rect 4614 22080 4620 22092
rect 4575 22052 4620 22080
rect 4614 22040 4620 22052
rect 4672 22040 4678 22092
rect 5350 22080 5356 22092
rect 5311 22052 5356 22080
rect 5350 22040 5356 22052
rect 5408 22040 5414 22092
rect 5810 22080 5816 22092
rect 5771 22052 5816 22080
rect 5810 22040 5816 22052
rect 5868 22040 5874 22092
rect 6270 22040 6276 22092
rect 6328 22080 6334 22092
rect 6457 22083 6515 22089
rect 6457 22080 6469 22083
rect 6328 22052 6469 22080
rect 6328 22040 6334 22052
rect 6457 22049 6469 22052
rect 6503 22049 6515 22083
rect 6914 22080 6920 22092
rect 6875 22052 6920 22080
rect 6457 22043 6515 22049
rect 6914 22040 6920 22052
rect 6972 22080 6978 22092
rect 7098 22080 7104 22092
rect 6972 22052 7104 22080
rect 6972 22040 6978 22052
rect 7098 22040 7104 22052
rect 7156 22040 7162 22092
rect 7469 22083 7527 22089
rect 7469 22049 7481 22083
rect 7515 22049 7527 22083
rect 7742 22080 7748 22092
rect 7703 22052 7748 22080
rect 7469 22043 7527 22049
rect 4890 22012 4896 22024
rect 3804 21984 4896 22012
rect 4890 21972 4896 21984
rect 4948 22012 4954 22024
rect 6549 22015 6607 22021
rect 6549 22012 6561 22015
rect 4948 21984 6561 22012
rect 4948 21972 4954 21984
rect 6549 21981 6561 21984
rect 6595 21981 6607 22015
rect 7484 22012 7512 22043
rect 7742 22040 7748 22052
rect 7800 22040 7806 22092
rect 8110 22040 8116 22092
rect 8168 22080 8174 22092
rect 8389 22083 8447 22089
rect 8389 22080 8401 22083
rect 8168 22052 8401 22080
rect 8168 22040 8174 22052
rect 8389 22049 8401 22052
rect 8435 22049 8447 22083
rect 8389 22043 8447 22049
rect 8496 22024 8524 22188
rect 8570 22176 8576 22188
rect 8628 22176 8634 22228
rect 8665 22219 8723 22225
rect 8665 22185 8677 22219
rect 8711 22216 8723 22219
rect 8711 22188 9720 22216
rect 8711 22185 8723 22188
rect 8665 22179 8723 22185
rect 9692 22160 9720 22188
rect 11238 22176 11244 22228
rect 11296 22216 11302 22228
rect 11425 22219 11483 22225
rect 11425 22216 11437 22219
rect 11296 22188 11437 22216
rect 11296 22176 11302 22188
rect 11425 22185 11437 22188
rect 11471 22216 11483 22219
rect 12342 22216 12348 22228
rect 11471 22188 12348 22216
rect 11471 22185 11483 22188
rect 11425 22179 11483 22185
rect 12342 22176 12348 22188
rect 12400 22176 12406 22228
rect 13173 22219 13231 22225
rect 13173 22185 13185 22219
rect 13219 22216 13231 22219
rect 13538 22216 13544 22228
rect 13219 22188 13544 22216
rect 13219 22185 13231 22188
rect 13173 22179 13231 22185
rect 13538 22176 13544 22188
rect 13596 22176 13602 22228
rect 15746 22176 15752 22228
rect 15804 22216 15810 22228
rect 16850 22216 16856 22228
rect 15804 22188 16528 22216
rect 16811 22188 16856 22216
rect 15804 22176 15810 22188
rect 8754 22148 8760 22160
rect 8715 22120 8760 22148
rect 8754 22108 8760 22120
rect 8812 22108 8818 22160
rect 9674 22108 9680 22160
rect 9732 22148 9738 22160
rect 10962 22148 10968 22160
rect 9732 22120 10968 22148
rect 9732 22108 9738 22120
rect 10962 22108 10968 22120
rect 11020 22148 11026 22160
rect 11517 22151 11575 22157
rect 11517 22148 11529 22151
rect 11020 22120 11529 22148
rect 11020 22108 11026 22120
rect 11517 22117 11529 22120
rect 11563 22117 11575 22151
rect 16390 22148 16396 22160
rect 11517 22111 11575 22117
rect 15212 22120 16396 22148
rect 8573 22083 8631 22089
rect 8573 22049 8585 22083
rect 8619 22049 8631 22083
rect 8573 22043 8631 22049
rect 9125 22083 9183 22089
rect 9125 22049 9137 22083
rect 9171 22080 9183 22083
rect 10505 22083 10563 22089
rect 10505 22080 10517 22083
rect 9171 22052 10517 22080
rect 9171 22049 9183 22052
rect 9125 22043 9183 22049
rect 10505 22049 10517 22052
rect 10551 22049 10563 22083
rect 10505 22043 10563 22049
rect 10689 22083 10747 22089
rect 10689 22049 10701 22083
rect 10735 22080 10747 22083
rect 10870 22080 10876 22092
rect 10735 22052 10876 22080
rect 10735 22049 10747 22052
rect 10689 22043 10747 22049
rect 8294 22012 8300 22024
rect 7484 21984 8300 22012
rect 6549 21975 6607 21981
rect 8294 21972 8300 21984
rect 8352 21972 8358 22024
rect 8478 21972 8484 22024
rect 8536 21972 8542 22024
rect 2225 21947 2283 21953
rect 2225 21913 2237 21947
rect 2271 21944 2283 21947
rect 2406 21944 2412 21956
rect 2271 21916 2412 21944
rect 2271 21913 2283 21916
rect 2225 21907 2283 21913
rect 2406 21904 2412 21916
rect 2464 21944 2470 21956
rect 3786 21944 3792 21956
rect 2464 21916 3792 21944
rect 2464 21904 2470 21916
rect 3786 21904 3792 21916
rect 3844 21904 3850 21956
rect 8588 21944 8616 22043
rect 10870 22040 10876 22052
rect 10928 22080 10934 22092
rect 11333 22083 11391 22089
rect 11333 22080 11345 22083
rect 10928 22052 11345 22080
rect 10928 22040 10934 22052
rect 11333 22049 11345 22052
rect 11379 22049 11391 22083
rect 11333 22043 11391 22049
rect 11698 22040 11704 22092
rect 11756 22080 11762 22092
rect 11885 22083 11943 22089
rect 11885 22080 11897 22083
rect 11756 22052 11897 22080
rect 11756 22040 11762 22052
rect 11885 22049 11897 22052
rect 11931 22049 11943 22083
rect 12342 22080 12348 22092
rect 12303 22052 12348 22080
rect 11885 22043 11943 22049
rect 12342 22040 12348 22052
rect 12400 22040 12406 22092
rect 13170 22080 13176 22092
rect 13131 22052 13176 22080
rect 13170 22040 13176 22052
rect 13228 22040 13234 22092
rect 13725 22083 13783 22089
rect 13725 22049 13737 22083
rect 13771 22080 13783 22083
rect 13998 22080 14004 22092
rect 13771 22052 14004 22080
rect 13771 22049 13783 22052
rect 13725 22043 13783 22049
rect 13998 22040 14004 22052
rect 14056 22040 14062 22092
rect 14826 22080 14832 22092
rect 14787 22052 14832 22080
rect 14826 22040 14832 22052
rect 14884 22040 14890 22092
rect 9677 22015 9735 22021
rect 9677 21981 9689 22015
rect 9723 22012 9735 22015
rect 9950 22012 9956 22024
rect 9723 21984 9956 22012
rect 9723 21981 9735 21984
rect 9677 21975 9735 21981
rect 9950 21972 9956 21984
rect 10008 21972 10014 22024
rect 10226 22012 10232 22024
rect 10187 21984 10232 22012
rect 10226 21972 10232 21984
rect 10284 21972 10290 22024
rect 11054 21972 11060 22024
rect 11112 22012 11118 22024
rect 11149 22015 11207 22021
rect 11149 22012 11161 22015
rect 11112 21984 11161 22012
rect 11112 21972 11118 21984
rect 11149 21981 11161 21984
rect 11195 21981 11207 22015
rect 13906 22012 13912 22024
rect 11149 21975 11207 21981
rect 11256 21984 12572 22012
rect 13867 21984 13912 22012
rect 10318 21944 10324 21956
rect 8588 21916 10324 21944
rect 10318 21904 10324 21916
rect 10376 21944 10382 21956
rect 11256 21944 11284 21984
rect 12544 21953 12572 21984
rect 13906 21972 13912 21984
rect 13964 21972 13970 22024
rect 15212 22012 15240 22120
rect 16390 22108 16396 22120
rect 16448 22108 16454 22160
rect 16500 22148 16528 22188
rect 16850 22176 16856 22188
rect 16908 22176 16914 22228
rect 18417 22219 18475 22225
rect 18417 22185 18429 22219
rect 18463 22185 18475 22219
rect 23750 22216 23756 22228
rect 23663 22188 23756 22216
rect 18417 22179 18475 22185
rect 18432 22148 18460 22179
rect 23750 22176 23756 22188
rect 23808 22216 23814 22228
rect 26697 22219 26755 22225
rect 26697 22216 26709 22219
rect 23808 22188 26709 22216
rect 23808 22176 23814 22188
rect 26697 22185 26709 22188
rect 26743 22185 26755 22219
rect 27706 22216 27712 22228
rect 27667 22188 27712 22216
rect 26697 22179 26755 22185
rect 27706 22176 27712 22188
rect 27764 22176 27770 22228
rect 27890 22176 27896 22228
rect 27948 22216 27954 22228
rect 27948 22188 29776 22216
rect 27948 22176 27954 22188
rect 16500 22120 18460 22148
rect 21082 22108 21088 22160
rect 21140 22148 21146 22160
rect 22002 22148 22008 22160
rect 21140 22120 22008 22148
rect 21140 22108 21146 22120
rect 15289 22083 15347 22089
rect 15289 22049 15301 22083
rect 15335 22049 15347 22083
rect 15289 22043 15347 22049
rect 14660 21984 15240 22012
rect 10376 21916 11284 21944
rect 12529 21947 12587 21953
rect 10376 21904 10382 21916
rect 12529 21913 12541 21947
rect 12575 21913 12587 21947
rect 12529 21907 12587 21913
rect 1581 21879 1639 21885
rect 1581 21845 1593 21879
rect 1627 21876 1639 21879
rect 1670 21876 1676 21888
rect 1627 21848 1676 21876
rect 1627 21845 1639 21848
rect 1581 21839 1639 21845
rect 1670 21836 1676 21848
rect 1728 21836 1734 21888
rect 2866 21876 2872 21888
rect 2827 21848 2872 21876
rect 2866 21836 2872 21848
rect 2924 21836 2930 21888
rect 3050 21836 3056 21888
rect 3108 21876 3114 21888
rect 4157 21879 4215 21885
rect 4157 21876 4169 21879
rect 3108 21848 4169 21876
rect 3108 21836 3114 21848
rect 4157 21845 4169 21848
rect 4203 21845 4215 21879
rect 4157 21839 4215 21845
rect 4982 21836 4988 21888
rect 5040 21876 5046 21888
rect 5353 21879 5411 21885
rect 5353 21876 5365 21879
rect 5040 21848 5365 21876
rect 5040 21836 5046 21848
rect 5353 21845 5365 21848
rect 5399 21845 5411 21879
rect 5353 21839 5411 21845
rect 13814 21836 13820 21888
rect 13872 21876 13878 21888
rect 14660 21885 14688 21984
rect 15304 21944 15332 22043
rect 15746 22040 15752 22092
rect 15804 22080 15810 22092
rect 15933 22083 15991 22089
rect 15933 22080 15945 22083
rect 15804 22052 15945 22080
rect 15804 22040 15810 22052
rect 15933 22049 15945 22052
rect 15979 22049 15991 22083
rect 15933 22043 15991 22049
rect 16206 22040 16212 22092
rect 16264 22080 16270 22092
rect 16301 22083 16359 22089
rect 16301 22080 16313 22083
rect 16264 22052 16313 22080
rect 16264 22040 16270 22052
rect 16301 22049 16313 22052
rect 16347 22049 16359 22083
rect 17129 22083 17187 22089
rect 17129 22080 17141 22083
rect 16301 22043 16359 22049
rect 16408 22052 17141 22080
rect 16408 22024 16436 22052
rect 17129 22049 17141 22052
rect 17175 22049 17187 22083
rect 17129 22043 17187 22049
rect 17589 22083 17647 22089
rect 17589 22049 17601 22083
rect 17635 22080 17647 22083
rect 17954 22080 17960 22092
rect 17635 22052 17960 22080
rect 17635 22049 17647 22052
rect 17589 22043 17647 22049
rect 17954 22040 17960 22052
rect 18012 22040 18018 22092
rect 18233 22083 18291 22089
rect 18233 22049 18245 22083
rect 18279 22080 18291 22083
rect 19150 22080 19156 22092
rect 18279 22052 19156 22080
rect 18279 22049 18291 22052
rect 18233 22043 18291 22049
rect 19150 22040 19156 22052
rect 19208 22040 19214 22092
rect 19245 22083 19303 22089
rect 19245 22049 19257 22083
rect 19291 22080 19303 22083
rect 19334 22080 19340 22092
rect 19291 22052 19340 22080
rect 19291 22049 19303 22052
rect 19245 22043 19303 22049
rect 19334 22040 19340 22052
rect 19392 22040 19398 22092
rect 19426 22040 19432 22092
rect 19484 22080 19490 22092
rect 20165 22083 20223 22089
rect 19484 22052 19529 22080
rect 19484 22040 19490 22052
rect 20165 22049 20177 22083
rect 20211 22080 20223 22083
rect 20254 22080 20260 22092
rect 20211 22052 20260 22080
rect 20211 22049 20223 22052
rect 20165 22043 20223 22049
rect 20254 22040 20260 22052
rect 20312 22040 20318 22092
rect 20901 22083 20959 22089
rect 20901 22049 20913 22083
rect 20947 22049 20959 22083
rect 20901 22043 20959 22049
rect 16390 21972 16396 22024
rect 16448 21972 16454 22024
rect 17862 21972 17868 22024
rect 17920 22012 17926 22024
rect 19521 22015 19579 22021
rect 19521 22012 19533 22015
rect 17920 21984 19533 22012
rect 17920 21972 17926 21984
rect 19521 21981 19533 21984
rect 19567 21981 19579 22015
rect 20916 22012 20944 22043
rect 20990 22040 20996 22092
rect 21048 22080 21054 22092
rect 21542 22080 21548 22092
rect 21048 22052 21548 22080
rect 21048 22040 21054 22052
rect 21542 22040 21548 22052
rect 21600 22040 21606 22092
rect 21652 22089 21680 22120
rect 22002 22108 22008 22120
rect 22060 22108 22066 22160
rect 23768 22148 23796 22176
rect 23676 22120 23796 22148
rect 24765 22151 24823 22157
rect 21637 22083 21695 22089
rect 21637 22049 21649 22083
rect 21683 22049 21695 22083
rect 21637 22043 21695 22049
rect 21818 22040 21824 22092
rect 21876 22080 21882 22092
rect 22373 22083 22431 22089
rect 22373 22080 22385 22083
rect 21876 22052 22385 22080
rect 21876 22040 21882 22052
rect 22373 22049 22385 22052
rect 22419 22049 22431 22083
rect 22738 22080 22744 22092
rect 22699 22052 22744 22080
rect 22373 22043 22431 22049
rect 22738 22040 22744 22052
rect 22796 22040 22802 22092
rect 22830 22040 22836 22092
rect 22888 22080 22894 22092
rect 23382 22080 23388 22092
rect 22888 22052 23388 22080
rect 22888 22040 22894 22052
rect 23382 22040 23388 22052
rect 23440 22040 23446 22092
rect 23676 22089 23704 22120
rect 24765 22117 24777 22151
rect 24811 22148 24823 22151
rect 25130 22148 25136 22160
rect 24811 22120 25136 22148
rect 24811 22117 24823 22120
rect 24765 22111 24823 22117
rect 25130 22108 25136 22120
rect 25188 22108 25194 22160
rect 25498 22108 25504 22160
rect 25556 22148 25562 22160
rect 29086 22148 29092 22160
rect 25556 22120 25728 22148
rect 25556 22108 25562 22120
rect 23661 22083 23719 22089
rect 23661 22049 23673 22083
rect 23707 22049 23719 22083
rect 25222 22080 25228 22092
rect 23661 22043 23719 22049
rect 23768 22052 25228 22080
rect 22848 22012 22876 22040
rect 23768 22021 23796 22052
rect 25222 22040 25228 22052
rect 25280 22040 25286 22092
rect 25409 22083 25467 22089
rect 25409 22049 25421 22083
rect 25455 22080 25467 22083
rect 25590 22080 25596 22092
rect 25455 22052 25596 22080
rect 25455 22049 25467 22052
rect 25409 22043 25467 22049
rect 25590 22040 25596 22052
rect 25648 22040 25654 22092
rect 25700 22089 25728 22120
rect 28920 22120 29092 22148
rect 25685 22083 25743 22089
rect 25685 22049 25697 22083
rect 25731 22049 25743 22083
rect 26510 22080 26516 22092
rect 26471 22052 26516 22080
rect 25685 22043 25743 22049
rect 26510 22040 26516 22052
rect 26568 22040 26574 22092
rect 27614 22080 27620 22092
rect 27575 22052 27620 22080
rect 27614 22040 27620 22052
rect 27672 22040 27678 22092
rect 27798 22040 27804 22092
rect 27856 22080 27862 22092
rect 27893 22083 27951 22089
rect 27893 22080 27905 22083
rect 27856 22052 27905 22080
rect 27856 22040 27862 22052
rect 27893 22049 27905 22052
rect 27939 22049 27951 22083
rect 27893 22043 27951 22049
rect 28261 22083 28319 22089
rect 28261 22049 28273 22083
rect 28307 22080 28319 22083
rect 28920 22080 28948 22120
rect 29086 22108 29092 22120
rect 29144 22108 29150 22160
rect 28307 22052 28948 22080
rect 28997 22083 29055 22089
rect 28307 22049 28319 22052
rect 28261 22043 28319 22049
rect 28997 22049 29009 22083
rect 29043 22080 29055 22083
rect 29638 22080 29644 22092
rect 29043 22052 29132 22080
rect 29599 22052 29644 22080
rect 29043 22049 29055 22052
rect 28997 22043 29055 22049
rect 20916 21984 22876 22012
rect 23753 22015 23811 22021
rect 19521 21975 19579 21981
rect 23753 21981 23765 22015
rect 23799 21981 23811 22015
rect 23753 21975 23811 21981
rect 25041 22015 25099 22021
rect 25041 21981 25053 22015
rect 25087 22012 25099 22015
rect 25958 22012 25964 22024
rect 25087 21984 25820 22012
rect 25919 21984 25964 22012
rect 25087 21981 25099 21984
rect 25041 21975 25099 21981
rect 22646 21944 22652 21956
rect 15304 21916 22652 21944
rect 22646 21904 22652 21916
rect 22704 21904 22710 21956
rect 25792 21944 25820 21984
rect 25958 21972 25964 21984
rect 26016 21972 26022 22024
rect 27908 22012 27936 22043
rect 29104 22024 29132 22052
rect 29638 22040 29644 22052
rect 29696 22040 29702 22092
rect 28718 22012 28724 22024
rect 27908 21984 28724 22012
rect 28718 21972 28724 21984
rect 28776 21972 28782 22024
rect 29086 21972 29092 22024
rect 29144 21972 29150 22024
rect 29748 22012 29776 22188
rect 30190 22176 30196 22228
rect 30248 22216 30254 22228
rect 35894 22216 35900 22228
rect 30248 22188 35900 22216
rect 30248 22176 30254 22188
rect 35894 22176 35900 22188
rect 35952 22176 35958 22228
rect 33226 22108 33232 22160
rect 33284 22148 33290 22160
rect 33686 22148 33692 22160
rect 33284 22120 33692 22148
rect 33284 22108 33290 22120
rect 33686 22108 33692 22120
rect 33744 22108 33750 22160
rect 35084 22120 35572 22148
rect 35084 22092 35112 22120
rect 29917 22083 29975 22089
rect 29917 22049 29929 22083
rect 29963 22080 29975 22083
rect 30006 22080 30012 22092
rect 29963 22052 30012 22080
rect 29963 22049 29975 22052
rect 29917 22043 29975 22049
rect 30006 22040 30012 22052
rect 30064 22040 30070 22092
rect 34517 22083 34575 22089
rect 34517 22049 34529 22083
rect 34563 22080 34575 22083
rect 34563 22052 34652 22080
rect 34563 22049 34575 22052
rect 34517 22043 34575 22049
rect 34624 22024 34652 22052
rect 35066 22040 35072 22092
rect 35124 22040 35130 22092
rect 35250 22080 35256 22092
rect 35211 22052 35256 22080
rect 35250 22040 35256 22052
rect 35308 22040 35314 22092
rect 35434 22080 35440 22092
rect 35395 22052 35440 22080
rect 35434 22040 35440 22052
rect 35492 22040 35498 22092
rect 35544 22080 35572 22120
rect 36998 22108 37004 22160
rect 37056 22148 37062 22160
rect 37056 22120 38332 22148
rect 37056 22108 37062 22120
rect 35805 22083 35863 22089
rect 35805 22080 35817 22083
rect 35544 22052 35817 22080
rect 35805 22049 35817 22052
rect 35851 22049 35863 22083
rect 36173 22083 36231 22089
rect 36173 22080 36185 22083
rect 35805 22043 35863 22049
rect 35912 22052 36185 22080
rect 31021 22015 31079 22021
rect 31021 22012 31033 22015
rect 29748 21984 31033 22012
rect 31021 21981 31033 21984
rect 31067 21981 31079 22015
rect 32122 22012 32128 22024
rect 32083 21984 32128 22012
rect 31021 21975 31079 21981
rect 32122 21972 32128 21984
rect 32180 21972 32186 22024
rect 32398 22012 32404 22024
rect 32359 21984 32404 22012
rect 32398 21972 32404 21984
rect 32456 21972 32462 22024
rect 34606 21972 34612 22024
rect 34664 21972 34670 22024
rect 35158 22012 35164 22024
rect 35119 21984 35164 22012
rect 35158 21972 35164 21984
rect 35216 21972 35222 22024
rect 26234 21944 26240 21956
rect 25792 21916 26240 21944
rect 26234 21904 26240 21916
rect 26292 21904 26298 21956
rect 33502 21904 33508 21956
rect 33560 21944 33566 21956
rect 34882 21944 34888 21956
rect 33560 21916 34888 21944
rect 33560 21904 33566 21916
rect 34882 21904 34888 21916
rect 34940 21904 34946 21956
rect 14645 21879 14703 21885
rect 14645 21876 14657 21879
rect 13872 21848 14657 21876
rect 13872 21836 13878 21848
rect 14645 21845 14657 21848
rect 14691 21845 14703 21879
rect 15378 21876 15384 21888
rect 15339 21848 15384 21876
rect 14645 21839 14703 21845
rect 15378 21836 15384 21848
rect 15436 21836 15442 21888
rect 19426 21836 19432 21888
rect 19484 21876 19490 21888
rect 20257 21879 20315 21885
rect 20257 21876 20269 21879
rect 19484 21848 20269 21876
rect 19484 21836 19490 21848
rect 20257 21845 20269 21848
rect 20303 21876 20315 21879
rect 20530 21876 20536 21888
rect 20303 21848 20536 21876
rect 20303 21845 20315 21848
rect 20257 21839 20315 21845
rect 20530 21836 20536 21848
rect 20588 21836 20594 21888
rect 21085 21879 21143 21885
rect 21085 21845 21097 21879
rect 21131 21876 21143 21879
rect 21358 21876 21364 21888
rect 21131 21848 21364 21876
rect 21131 21845 21143 21848
rect 21085 21839 21143 21845
rect 21358 21836 21364 21848
rect 21416 21876 21422 21888
rect 21542 21876 21548 21888
rect 21416 21848 21548 21876
rect 21416 21836 21422 21848
rect 21542 21836 21548 21848
rect 21600 21836 21606 21888
rect 21821 21879 21879 21885
rect 21821 21845 21833 21879
rect 21867 21876 21879 21879
rect 22922 21876 22928 21888
rect 21867 21848 22928 21876
rect 21867 21845 21879 21848
rect 21821 21839 21879 21845
rect 22922 21836 22928 21848
rect 22980 21836 22986 21888
rect 24765 21879 24823 21885
rect 24765 21845 24777 21879
rect 24811 21876 24823 21879
rect 24854 21876 24860 21888
rect 24811 21848 24860 21876
rect 24811 21845 24823 21848
rect 24765 21839 24823 21845
rect 24854 21836 24860 21848
rect 24912 21836 24918 21888
rect 29086 21876 29092 21888
rect 29047 21848 29092 21876
rect 29086 21836 29092 21848
rect 29144 21836 29150 21888
rect 33686 21876 33692 21888
rect 33647 21848 33692 21876
rect 33686 21836 33692 21848
rect 33744 21836 33750 21888
rect 34790 21836 34796 21888
rect 34848 21876 34854 21888
rect 35912 21876 35940 22052
rect 36173 22049 36185 22052
rect 36219 22080 36231 22083
rect 36909 22083 36967 22089
rect 36909 22080 36921 22083
rect 36219 22052 36921 22080
rect 36219 22049 36231 22052
rect 36173 22043 36231 22049
rect 36909 22049 36921 22052
rect 36955 22049 36967 22083
rect 36909 22043 36967 22049
rect 37826 22040 37832 22092
rect 37884 22080 37890 22092
rect 38304 22089 38332 22120
rect 38289 22083 38347 22089
rect 37884 22052 37929 22080
rect 37884 22040 37890 22052
rect 38289 22049 38301 22083
rect 38335 22049 38347 22083
rect 38289 22043 38347 22049
rect 38565 22015 38623 22021
rect 38565 21981 38577 22015
rect 38611 21981 38623 22015
rect 38565 21975 38623 21981
rect 36814 21904 36820 21956
rect 36872 21944 36878 21956
rect 36872 21916 37228 21944
rect 36872 21904 36878 21916
rect 34848 21848 35940 21876
rect 34848 21836 34854 21848
rect 36446 21836 36452 21888
rect 36504 21876 36510 21888
rect 37093 21879 37151 21885
rect 37093 21876 37105 21879
rect 36504 21848 37105 21876
rect 36504 21836 36510 21848
rect 37093 21845 37105 21848
rect 37139 21845 37151 21879
rect 37200 21876 37228 21916
rect 37550 21904 37556 21956
rect 37608 21944 37614 21956
rect 37829 21947 37887 21953
rect 37829 21944 37841 21947
rect 37608 21916 37841 21944
rect 37608 21904 37614 21916
rect 37829 21913 37841 21916
rect 37875 21913 37887 21947
rect 37829 21907 37887 21913
rect 38580 21876 38608 21975
rect 37200 21848 38608 21876
rect 37093 21839 37151 21845
rect 1104 21786 39836 21808
rect 1104 21734 4246 21786
rect 4298 21734 4310 21786
rect 4362 21734 4374 21786
rect 4426 21734 4438 21786
rect 4490 21734 34966 21786
rect 35018 21734 35030 21786
rect 35082 21734 35094 21786
rect 35146 21734 35158 21786
rect 35210 21734 39836 21786
rect 1104 21712 39836 21734
rect 3697 21675 3755 21681
rect 3697 21641 3709 21675
rect 3743 21672 3755 21675
rect 4062 21672 4068 21684
rect 3743 21644 4068 21672
rect 3743 21641 3755 21644
rect 3697 21635 3755 21641
rect 4062 21632 4068 21644
rect 4120 21632 4126 21684
rect 6822 21632 6828 21684
rect 6880 21672 6886 21684
rect 8021 21675 8079 21681
rect 8021 21672 8033 21675
rect 6880 21644 8033 21672
rect 6880 21632 6886 21644
rect 8021 21641 8033 21644
rect 8067 21672 8079 21675
rect 9858 21672 9864 21684
rect 8067 21644 9864 21672
rect 8067 21641 8079 21644
rect 8021 21635 8079 21641
rect 9858 21632 9864 21644
rect 9916 21672 9922 21684
rect 11054 21672 11060 21684
rect 9916 21644 11060 21672
rect 9916 21632 9922 21644
rect 11054 21632 11060 21644
rect 11112 21632 11118 21684
rect 11514 21672 11520 21684
rect 11475 21644 11520 21672
rect 11514 21632 11520 21644
rect 11572 21632 11578 21684
rect 15470 21632 15476 21684
rect 15528 21672 15534 21684
rect 18233 21675 18291 21681
rect 18233 21672 18245 21675
rect 15528 21644 18245 21672
rect 15528 21632 15534 21644
rect 18233 21641 18245 21644
rect 18279 21641 18291 21675
rect 18233 21635 18291 21641
rect 19334 21632 19340 21684
rect 19392 21672 19398 21684
rect 20070 21672 20076 21684
rect 19392 21644 20076 21672
rect 19392 21632 19398 21644
rect 20070 21632 20076 21644
rect 20128 21672 20134 21684
rect 20165 21675 20223 21681
rect 20165 21672 20177 21675
rect 20128 21644 20177 21672
rect 20128 21632 20134 21644
rect 20165 21641 20177 21644
rect 20211 21641 20223 21675
rect 20165 21635 20223 21641
rect 20824 21644 23336 21672
rect 1486 21564 1492 21616
rect 1544 21604 1550 21616
rect 4801 21607 4859 21613
rect 4801 21604 4813 21607
rect 1544 21576 4813 21604
rect 1544 21564 1550 21576
rect 4801 21573 4813 21576
rect 4847 21573 4859 21607
rect 4801 21567 4859 21573
rect 7285 21607 7343 21613
rect 7285 21573 7297 21607
rect 7331 21604 7343 21607
rect 8386 21604 8392 21616
rect 7331 21576 8392 21604
rect 7331 21573 7343 21576
rect 7285 21567 7343 21573
rect 8386 21564 8392 21576
rect 8444 21564 8450 21616
rect 9674 21564 9680 21616
rect 9732 21604 9738 21616
rect 14274 21604 14280 21616
rect 9732 21576 10548 21604
rect 14235 21576 14280 21604
rect 9732 21564 9738 21576
rect 2866 21536 2872 21548
rect 1688 21508 2872 21536
rect 1688 21477 1716 21508
rect 2866 21496 2872 21508
rect 2924 21496 2930 21548
rect 8938 21536 8944 21548
rect 5276 21508 8944 21536
rect 1673 21471 1731 21477
rect 1673 21437 1685 21471
rect 1719 21437 1731 21471
rect 1673 21431 1731 21437
rect 1765 21471 1823 21477
rect 1765 21437 1777 21471
rect 1811 21468 1823 21471
rect 2590 21468 2596 21480
rect 1811 21440 2596 21468
rect 1811 21437 1823 21440
rect 1765 21431 1823 21437
rect 2590 21428 2596 21440
rect 2648 21428 2654 21480
rect 2958 21468 2964 21480
rect 2919 21440 2964 21468
rect 2958 21428 2964 21440
rect 3016 21428 3022 21480
rect 3145 21471 3203 21477
rect 3145 21437 3157 21471
rect 3191 21437 3203 21471
rect 3145 21431 3203 21437
rect 3160 21400 3188 21431
rect 3234 21428 3240 21480
rect 3292 21468 3298 21480
rect 3605 21471 3663 21477
rect 3605 21468 3617 21471
rect 3292 21440 3617 21468
rect 3292 21428 3298 21440
rect 3605 21437 3617 21440
rect 3651 21437 3663 21471
rect 4982 21468 4988 21480
rect 4943 21440 4988 21468
rect 3605 21431 3663 21437
rect 4982 21428 4988 21440
rect 5040 21428 5046 21480
rect 5276 21477 5304 21508
rect 8938 21496 8944 21508
rect 8996 21496 9002 21548
rect 9217 21539 9275 21545
rect 9217 21505 9229 21539
rect 9263 21536 9275 21539
rect 10226 21536 10232 21548
rect 9263 21508 10232 21536
rect 9263 21505 9275 21508
rect 9217 21499 9275 21505
rect 10226 21496 10232 21508
rect 10284 21496 10290 21548
rect 5261 21471 5319 21477
rect 5261 21437 5273 21471
rect 5307 21437 5319 21471
rect 5442 21468 5448 21480
rect 5403 21440 5448 21468
rect 5261 21431 5319 21437
rect 5442 21428 5448 21440
rect 5500 21428 5506 21480
rect 7101 21471 7159 21477
rect 7101 21437 7113 21471
rect 7147 21468 7159 21471
rect 7190 21468 7196 21480
rect 7147 21440 7196 21468
rect 7147 21437 7159 21440
rect 7101 21431 7159 21437
rect 7190 21428 7196 21440
rect 7248 21428 7254 21480
rect 7837 21471 7895 21477
rect 7837 21437 7849 21471
rect 7883 21468 7895 21471
rect 8018 21468 8024 21480
rect 7883 21440 8024 21468
rect 7883 21437 7895 21440
rect 7837 21431 7895 21437
rect 8018 21428 8024 21440
rect 8076 21428 8082 21480
rect 8386 21428 8392 21480
rect 8444 21468 8450 21480
rect 9125 21471 9183 21477
rect 9125 21468 9137 21471
rect 8444 21440 9137 21468
rect 8444 21428 8450 21440
rect 9125 21437 9137 21440
rect 9171 21437 9183 21471
rect 9125 21431 9183 21437
rect 9585 21471 9643 21477
rect 9585 21437 9597 21471
rect 9631 21437 9643 21471
rect 9858 21468 9864 21480
rect 9819 21440 9864 21468
rect 9585 21431 9643 21437
rect 3786 21400 3792 21412
rect 3160 21372 3792 21400
rect 3786 21360 3792 21372
rect 3844 21400 3850 21412
rect 4798 21400 4804 21412
rect 3844 21372 4804 21400
rect 3844 21360 3850 21372
rect 4798 21360 4804 21372
rect 4856 21360 4862 21412
rect 9140 21400 9168 21431
rect 9214 21400 9220 21412
rect 9140 21372 9220 21400
rect 9214 21360 9220 21372
rect 9272 21360 9278 21412
rect 9600 21400 9628 21431
rect 9858 21428 9864 21440
rect 9916 21428 9922 21480
rect 10318 21468 10324 21480
rect 10279 21440 10324 21468
rect 10318 21428 10324 21440
rect 10376 21428 10382 21480
rect 10520 21477 10548 21576
rect 14274 21564 14280 21576
rect 14332 21564 14338 21616
rect 12526 21496 12532 21548
rect 12584 21536 12590 21548
rect 13170 21536 13176 21548
rect 12584 21508 12756 21536
rect 13131 21508 13176 21536
rect 12584 21496 12590 21508
rect 10505 21471 10563 21477
rect 10505 21437 10517 21471
rect 10551 21437 10563 21471
rect 11238 21468 11244 21480
rect 11199 21440 11244 21468
rect 10505 21431 10563 21437
rect 11238 21428 11244 21440
rect 11296 21428 11302 21480
rect 11333 21471 11391 21477
rect 11333 21437 11345 21471
rect 11379 21437 11391 21471
rect 11333 21431 11391 21437
rect 12437 21471 12495 21477
rect 12437 21437 12449 21471
rect 12483 21437 12495 21471
rect 12618 21468 12624 21480
rect 12579 21440 12624 21468
rect 12437 21431 12495 21437
rect 10870 21400 10876 21412
rect 9600 21372 10876 21400
rect 10870 21360 10876 21372
rect 10928 21360 10934 21412
rect 10962 21360 10968 21412
rect 11020 21400 11026 21412
rect 11348 21400 11376 21431
rect 11020 21372 11376 21400
rect 12452 21400 12480 21431
rect 12618 21428 12624 21440
rect 12676 21428 12682 21480
rect 12728 21477 12756 21508
rect 13170 21496 13176 21508
rect 13228 21496 13234 21548
rect 15488 21536 15516 21632
rect 16574 21604 16580 21616
rect 16535 21576 16580 21604
rect 16574 21564 16580 21576
rect 16632 21564 16638 21616
rect 20714 21604 20720 21616
rect 17880 21576 20720 21604
rect 14384 21508 15516 21536
rect 15933 21539 15991 21545
rect 12713 21471 12771 21477
rect 12713 21437 12725 21471
rect 12759 21437 12771 21471
rect 13814 21468 13820 21480
rect 13775 21440 13820 21468
rect 12713 21431 12771 21437
rect 13814 21428 13820 21440
rect 13872 21428 13878 21480
rect 14384 21477 14412 21508
rect 15933 21505 15945 21539
rect 15979 21536 15991 21539
rect 17586 21536 17592 21548
rect 15979 21508 17592 21536
rect 15979 21505 15991 21508
rect 15933 21499 15991 21505
rect 17586 21496 17592 21508
rect 17644 21496 17650 21548
rect 14369 21471 14427 21477
rect 14369 21437 14381 21471
rect 14415 21437 14427 21471
rect 14369 21431 14427 21437
rect 14921 21471 14979 21477
rect 14921 21437 14933 21471
rect 14967 21437 14979 21471
rect 14921 21431 14979 21437
rect 15105 21471 15163 21477
rect 15105 21437 15117 21471
rect 15151 21468 15163 21471
rect 15562 21468 15568 21480
rect 15151 21440 15568 21468
rect 15151 21437 15163 21440
rect 15105 21431 15163 21437
rect 13078 21400 13084 21412
rect 12452 21372 13084 21400
rect 11020 21360 11026 21372
rect 13078 21360 13084 21372
rect 13136 21360 13142 21412
rect 14936 21400 14964 21431
rect 15562 21428 15568 21440
rect 15620 21428 15626 21480
rect 16301 21471 16359 21477
rect 16301 21437 16313 21471
rect 16347 21468 16359 21471
rect 16574 21468 16580 21480
rect 16347 21440 16580 21468
rect 16347 21437 16359 21440
rect 16301 21431 16359 21437
rect 16574 21428 16580 21440
rect 16632 21428 16638 21480
rect 16669 21471 16727 21477
rect 16669 21437 16681 21471
rect 16715 21468 16727 21471
rect 16758 21468 16764 21480
rect 16715 21440 16764 21468
rect 16715 21437 16727 21440
rect 16669 21431 16727 21437
rect 16758 21428 16764 21440
rect 16816 21428 16822 21480
rect 17313 21471 17371 21477
rect 17313 21437 17325 21471
rect 17359 21468 17371 21471
rect 17880 21468 17908 21576
rect 20714 21564 20720 21576
rect 20772 21564 20778 21616
rect 18877 21539 18935 21545
rect 18877 21505 18889 21539
rect 18923 21536 18935 21539
rect 19150 21536 19156 21548
rect 18923 21508 19156 21536
rect 18923 21505 18935 21508
rect 18877 21499 18935 21505
rect 19150 21496 19156 21508
rect 19208 21496 19214 21548
rect 19242 21496 19248 21548
rect 19300 21536 19306 21548
rect 19613 21539 19671 21545
rect 19613 21536 19625 21539
rect 19300 21508 19625 21536
rect 19300 21496 19306 21508
rect 19613 21505 19625 21508
rect 19659 21505 19671 21539
rect 19613 21499 19671 21505
rect 18046 21468 18052 21480
rect 17359 21440 17908 21468
rect 18007 21440 18052 21468
rect 17359 21437 17371 21440
rect 17313 21431 17371 21437
rect 18046 21428 18052 21440
rect 18104 21428 18110 21480
rect 19061 21471 19119 21477
rect 19061 21437 19073 21471
rect 19107 21468 19119 21471
rect 19426 21468 19432 21480
rect 19107 21440 19432 21468
rect 19107 21437 19119 21440
rect 19061 21431 19119 21437
rect 19426 21428 19432 21440
rect 19484 21428 19490 21480
rect 20073 21471 20131 21477
rect 20073 21437 20085 21471
rect 20119 21437 20131 21471
rect 20073 21431 20131 21437
rect 15838 21400 15844 21412
rect 14936 21372 15844 21400
rect 15838 21360 15844 21372
rect 15896 21360 15902 21412
rect 19242 21400 19248 21412
rect 19155 21372 19248 21400
rect 19242 21360 19248 21372
rect 19300 21400 19306 21412
rect 19886 21400 19892 21412
rect 19300 21372 19892 21400
rect 19300 21360 19306 21372
rect 19886 21360 19892 21372
rect 19944 21400 19950 21412
rect 20088 21400 20116 21431
rect 20162 21428 20168 21480
rect 20220 21468 20226 21480
rect 20824 21477 20852 21644
rect 21726 21564 21732 21616
rect 21784 21604 21790 21616
rect 22002 21604 22008 21616
rect 21784 21576 22008 21604
rect 21784 21564 21790 21576
rect 22002 21564 22008 21576
rect 22060 21564 22066 21616
rect 23308 21604 23336 21644
rect 23382 21632 23388 21684
rect 23440 21672 23446 21684
rect 25041 21675 25099 21681
rect 25041 21672 25053 21675
rect 23440 21644 25053 21672
rect 23440 21632 23446 21644
rect 25041 21641 25053 21644
rect 25087 21641 25099 21675
rect 25041 21635 25099 21641
rect 25222 21632 25228 21684
rect 25280 21672 25286 21684
rect 28994 21672 29000 21684
rect 25280 21644 29000 21672
rect 25280 21632 25286 21644
rect 28994 21632 29000 21644
rect 29052 21632 29058 21684
rect 29086 21632 29092 21684
rect 29144 21672 29150 21684
rect 33778 21672 33784 21684
rect 29144 21644 33784 21672
rect 29144 21632 29150 21644
rect 33778 21632 33784 21644
rect 33836 21632 33842 21684
rect 34149 21675 34207 21681
rect 34149 21641 34161 21675
rect 34195 21672 34207 21675
rect 34790 21672 34796 21684
rect 34195 21644 34796 21672
rect 34195 21641 34207 21644
rect 34149 21635 34207 21641
rect 34790 21632 34796 21644
rect 34848 21632 34854 21684
rect 38838 21672 38844 21684
rect 38799 21644 38844 21672
rect 38838 21632 38844 21644
rect 38896 21632 38902 21684
rect 23566 21604 23572 21616
rect 23308 21576 23572 21604
rect 23566 21564 23572 21576
rect 23624 21564 23630 21616
rect 25406 21564 25412 21616
rect 25464 21604 25470 21616
rect 25869 21607 25927 21613
rect 25869 21604 25881 21607
rect 25464 21576 25881 21604
rect 25464 21564 25470 21576
rect 25869 21573 25881 21576
rect 25915 21573 25927 21607
rect 25869 21567 25927 21573
rect 28626 21564 28632 21616
rect 28684 21604 28690 21616
rect 28684 21576 29684 21604
rect 28684 21564 28690 21576
rect 21266 21496 21272 21548
rect 21324 21536 21330 21548
rect 21910 21536 21916 21548
rect 21324 21508 21772 21536
rect 21871 21508 21916 21536
rect 21324 21496 21330 21508
rect 20809 21471 20867 21477
rect 20809 21468 20821 21471
rect 20220 21440 20821 21468
rect 20220 21428 20226 21440
rect 20809 21437 20821 21440
rect 20855 21437 20867 21471
rect 21450 21468 21456 21480
rect 21411 21440 21456 21468
rect 20809 21431 20867 21437
rect 21450 21428 21456 21440
rect 21508 21428 21514 21480
rect 21542 21428 21548 21480
rect 21600 21468 21606 21480
rect 21637 21471 21695 21477
rect 21637 21468 21649 21471
rect 21600 21440 21649 21468
rect 21600 21428 21606 21440
rect 21637 21437 21649 21440
rect 21683 21437 21695 21471
rect 21744 21468 21772 21508
rect 21910 21496 21916 21508
rect 21968 21496 21974 21548
rect 23474 21536 23480 21548
rect 22020 21508 23480 21536
rect 22020 21477 22048 21508
rect 23474 21496 23480 21508
rect 23532 21496 23538 21548
rect 23661 21539 23719 21545
rect 23661 21505 23673 21539
rect 23707 21536 23719 21539
rect 24854 21536 24860 21548
rect 23707 21508 24860 21536
rect 23707 21505 23719 21508
rect 23661 21499 23719 21505
rect 24854 21496 24860 21508
rect 24912 21496 24918 21548
rect 25958 21496 25964 21548
rect 26016 21536 26022 21548
rect 26605 21539 26663 21545
rect 26605 21536 26617 21539
rect 26016 21508 26617 21536
rect 26016 21496 26022 21508
rect 26605 21505 26617 21508
rect 26651 21505 26663 21539
rect 27706 21536 27712 21548
rect 27667 21508 27712 21536
rect 26605 21499 26663 21505
rect 27706 21496 27712 21508
rect 27764 21496 27770 21548
rect 22005 21471 22063 21477
rect 22005 21468 22017 21471
rect 21744 21440 22017 21468
rect 21637 21431 21695 21437
rect 22005 21437 22017 21440
rect 22051 21437 22063 21471
rect 22005 21431 22063 21437
rect 22925 21471 22983 21477
rect 22925 21437 22937 21471
rect 22971 21468 22983 21471
rect 23382 21468 23388 21480
rect 22971 21440 23388 21468
rect 22971 21437 22983 21440
rect 22925 21431 22983 21437
rect 23382 21428 23388 21440
rect 23440 21428 23446 21480
rect 23934 21468 23940 21480
rect 23895 21440 23940 21468
rect 23934 21428 23940 21440
rect 23992 21428 23998 21480
rect 25869 21471 25927 21477
rect 25869 21437 25881 21471
rect 25915 21437 25927 21471
rect 26510 21468 26516 21480
rect 26471 21440 26516 21468
rect 25869 21431 25927 21437
rect 23198 21400 23204 21412
rect 19944 21372 23204 21400
rect 19944 21360 19950 21372
rect 23198 21360 23204 21372
rect 23256 21360 23262 21412
rect 12250 21292 12256 21344
rect 12308 21332 12314 21344
rect 13633 21335 13691 21341
rect 13633 21332 13645 21335
rect 12308 21304 13645 21332
rect 12308 21292 12314 21304
rect 13633 21301 13645 21304
rect 13679 21301 13691 21335
rect 13633 21295 13691 21301
rect 17126 21292 17132 21344
rect 17184 21332 17190 21344
rect 17405 21335 17463 21341
rect 17405 21332 17417 21335
rect 17184 21304 17417 21332
rect 17184 21292 17190 21304
rect 17405 21301 17417 21304
rect 17451 21301 17463 21335
rect 17405 21295 17463 21301
rect 19153 21335 19211 21341
rect 19153 21301 19165 21335
rect 19199 21332 19211 21335
rect 19334 21332 19340 21344
rect 19199 21304 19340 21332
rect 19199 21301 19211 21304
rect 19153 21295 19211 21301
rect 19334 21292 19340 21304
rect 19392 21292 19398 21344
rect 19426 21292 19432 21344
rect 19484 21332 19490 21344
rect 22922 21332 22928 21344
rect 19484 21304 22928 21332
rect 19484 21292 19490 21304
rect 22922 21292 22928 21304
rect 22980 21292 22986 21344
rect 23017 21335 23075 21341
rect 23017 21301 23029 21335
rect 23063 21332 23075 21335
rect 24670 21332 24676 21344
rect 23063 21304 24676 21332
rect 23063 21301 23075 21304
rect 23017 21295 23075 21301
rect 24670 21292 24676 21304
rect 24728 21292 24734 21344
rect 25884 21332 25912 21431
rect 26510 21428 26516 21440
rect 26568 21428 26574 21480
rect 27982 21468 27988 21480
rect 27943 21440 27988 21468
rect 27982 21428 27988 21440
rect 28040 21428 28046 21480
rect 28537 21471 28595 21477
rect 28537 21437 28549 21471
rect 28583 21468 28595 21471
rect 28626 21468 28632 21480
rect 28583 21440 28632 21468
rect 28583 21437 28595 21440
rect 28537 21431 28595 21437
rect 28626 21428 28632 21440
rect 28684 21428 28690 21480
rect 29178 21428 29184 21480
rect 29236 21468 29242 21480
rect 29656 21477 29684 21576
rect 30282 21536 30288 21548
rect 30243 21508 30288 21536
rect 30282 21496 30288 21508
rect 30340 21496 30346 21548
rect 35437 21539 35495 21545
rect 35437 21536 35449 21539
rect 31864 21508 35449 21536
rect 31864 21480 31892 21508
rect 35437 21505 35449 21508
rect 35483 21536 35495 21539
rect 36630 21536 36636 21548
rect 35483 21508 36636 21536
rect 35483 21505 35495 21508
rect 35437 21499 35495 21505
rect 36630 21496 36636 21508
rect 36688 21496 36694 21548
rect 37550 21536 37556 21548
rect 37511 21508 37556 21536
rect 37550 21496 37556 21508
rect 37608 21496 37614 21548
rect 29273 21471 29331 21477
rect 29273 21468 29285 21471
rect 29236 21440 29285 21468
rect 29236 21428 29242 21440
rect 29273 21437 29285 21440
rect 29319 21437 29331 21471
rect 29273 21431 29331 21437
rect 29641 21471 29699 21477
rect 29641 21437 29653 21471
rect 29687 21437 29699 21471
rect 30098 21468 30104 21480
rect 30059 21440 30104 21468
rect 29641 21431 29699 21437
rect 30098 21428 30104 21440
rect 30156 21428 30162 21480
rect 30558 21468 30564 21480
rect 30519 21440 30564 21468
rect 30558 21428 30564 21440
rect 30616 21428 30622 21480
rect 31110 21428 31116 21480
rect 31168 21468 31174 21480
rect 31205 21471 31263 21477
rect 31205 21468 31217 21471
rect 31168 21440 31217 21468
rect 31168 21428 31174 21440
rect 31205 21437 31217 21440
rect 31251 21437 31263 21471
rect 31846 21468 31852 21480
rect 31759 21440 31852 21468
rect 31205 21431 31263 21437
rect 31846 21428 31852 21440
rect 31904 21428 31910 21480
rect 32030 21468 32036 21480
rect 31991 21440 32036 21468
rect 32030 21428 32036 21440
rect 32088 21428 32094 21480
rect 32306 21428 32312 21480
rect 32364 21468 32370 21480
rect 32769 21471 32827 21477
rect 32769 21468 32781 21471
rect 32364 21440 32781 21468
rect 32364 21428 32370 21440
rect 32769 21437 32781 21440
rect 32815 21437 32827 21471
rect 33226 21468 33232 21480
rect 33187 21440 33232 21468
rect 32769 21431 32827 21437
rect 33226 21428 33232 21440
rect 33284 21428 33290 21480
rect 33965 21471 34023 21477
rect 33965 21437 33977 21471
rect 34011 21437 34023 21471
rect 35710 21468 35716 21480
rect 35671 21440 35716 21468
rect 33965 21431 34023 21437
rect 28721 21403 28779 21409
rect 28721 21369 28733 21403
rect 28767 21400 28779 21403
rect 29822 21400 29828 21412
rect 28767 21372 29828 21400
rect 28767 21369 28779 21372
rect 28721 21363 28779 21369
rect 29822 21360 29828 21372
rect 29880 21360 29886 21412
rect 30006 21360 30012 21412
rect 30064 21400 30070 21412
rect 33980 21400 34008 21431
rect 35710 21428 35716 21440
rect 35768 21428 35774 21480
rect 35802 21428 35808 21480
rect 35860 21468 35866 21480
rect 35897 21471 35955 21477
rect 35897 21468 35909 21471
rect 35860 21440 35909 21468
rect 35860 21428 35866 21440
rect 35897 21437 35909 21440
rect 35943 21437 35955 21471
rect 35897 21431 35955 21437
rect 36078 21428 36084 21480
rect 36136 21468 36142 21480
rect 36354 21468 36360 21480
rect 36136 21440 36360 21468
rect 36136 21428 36142 21440
rect 36354 21428 36360 21440
rect 36412 21428 36418 21480
rect 37274 21468 37280 21480
rect 37235 21440 37280 21468
rect 37274 21428 37280 21440
rect 37332 21428 37338 21480
rect 30064 21372 34008 21400
rect 34885 21403 34943 21409
rect 30064 21360 30070 21372
rect 34885 21369 34897 21403
rect 34931 21400 34943 21403
rect 35250 21400 35256 21412
rect 34931 21372 35256 21400
rect 34931 21369 34943 21372
rect 34885 21363 34943 21369
rect 35250 21360 35256 21372
rect 35308 21360 35314 21412
rect 29270 21332 29276 21344
rect 25884 21304 29276 21332
rect 29270 21292 29276 21304
rect 29328 21292 29334 21344
rect 31294 21332 31300 21344
rect 31255 21304 31300 21332
rect 31294 21292 31300 21304
rect 31352 21292 31358 21344
rect 32398 21292 32404 21344
rect 32456 21332 32462 21344
rect 32861 21335 32919 21341
rect 32861 21332 32873 21335
rect 32456 21304 32873 21332
rect 32456 21292 32462 21304
rect 32861 21301 32873 21304
rect 32907 21301 32919 21335
rect 32861 21295 32919 21301
rect 34330 21292 34336 21344
rect 34388 21332 34394 21344
rect 36449 21335 36507 21341
rect 36449 21332 36461 21335
rect 34388 21304 36461 21332
rect 34388 21292 34394 21304
rect 36449 21301 36461 21304
rect 36495 21301 36507 21335
rect 36449 21295 36507 21301
rect 1104 21242 39836 21264
rect 1104 21190 19606 21242
rect 19658 21190 19670 21242
rect 19722 21190 19734 21242
rect 19786 21190 19798 21242
rect 19850 21190 39836 21242
rect 1104 21168 39836 21190
rect 11146 21088 11152 21140
rect 11204 21128 11210 21140
rect 11241 21131 11299 21137
rect 11241 21128 11253 21131
rect 11204 21100 11253 21128
rect 11204 21088 11210 21100
rect 11241 21097 11253 21100
rect 11287 21097 11299 21131
rect 11241 21091 11299 21097
rect 2958 21020 2964 21072
rect 3016 21060 3022 21072
rect 3053 21063 3111 21069
rect 3053 21060 3065 21063
rect 3016 21032 3065 21060
rect 3016 21020 3022 21032
rect 3053 21029 3065 21032
rect 3099 21060 3111 21063
rect 4706 21060 4712 21072
rect 3099 21032 4712 21060
rect 3099 21029 3111 21032
rect 3053 21023 3111 21029
rect 1394 20992 1400 21004
rect 1355 20964 1400 20992
rect 1394 20952 1400 20964
rect 1452 20952 1458 21004
rect 1670 20992 1676 21004
rect 1631 20964 1676 20992
rect 1670 20952 1676 20964
rect 1728 20952 1734 21004
rect 2590 20952 2596 21004
rect 2648 20992 2654 21004
rect 4632 21001 4660 21032
rect 4706 21020 4712 21032
rect 4764 21020 4770 21072
rect 5261 21063 5319 21069
rect 5261 21029 5273 21063
rect 5307 21060 5319 21063
rect 5442 21060 5448 21072
rect 5307 21032 5448 21060
rect 5307 21029 5319 21032
rect 5261 21023 5319 21029
rect 5442 21020 5448 21032
rect 5500 21020 5506 21072
rect 8018 21060 8024 21072
rect 7208 21032 8024 21060
rect 4341 20995 4399 21001
rect 4341 20992 4353 20995
rect 2648 20964 4353 20992
rect 2648 20952 2654 20964
rect 4341 20961 4353 20964
rect 4387 20961 4399 20995
rect 4341 20955 4399 20961
rect 4617 20995 4675 21001
rect 4617 20961 4629 20995
rect 4663 20961 4675 20995
rect 4798 20992 4804 21004
rect 4759 20964 4804 20992
rect 4617 20955 4675 20961
rect 4356 20924 4384 20955
rect 4798 20952 4804 20964
rect 4856 20952 4862 21004
rect 5721 20995 5779 21001
rect 5721 20961 5733 20995
rect 5767 20961 5779 20995
rect 6270 20992 6276 21004
rect 6231 20964 6276 20992
rect 5721 20955 5779 20961
rect 5736 20924 5764 20955
rect 6270 20952 6276 20964
rect 6328 20952 6334 21004
rect 6733 20995 6791 21001
rect 6733 20961 6745 20995
rect 6779 20992 6791 20995
rect 6914 20992 6920 21004
rect 6779 20964 6920 20992
rect 6779 20961 6791 20964
rect 6733 20955 6791 20961
rect 6914 20952 6920 20964
rect 6972 20952 6978 21004
rect 7208 21001 7236 21032
rect 8018 21020 8024 21032
rect 8076 21020 8082 21072
rect 7193 20995 7251 21001
rect 7193 20961 7205 20995
rect 7239 20961 7251 20995
rect 7834 20992 7840 21004
rect 7795 20964 7840 20992
rect 7193 20955 7251 20961
rect 7834 20952 7840 20964
rect 7892 20952 7898 21004
rect 8386 20992 8392 21004
rect 8347 20964 8392 20992
rect 8386 20952 8392 20964
rect 8444 20952 8450 21004
rect 8849 20995 8907 21001
rect 8849 20961 8861 20995
rect 8895 20961 8907 20995
rect 8849 20955 8907 20961
rect 9677 20995 9735 21001
rect 9677 20961 9689 20995
rect 9723 20992 9735 20995
rect 9766 20992 9772 21004
rect 9723 20964 9772 20992
rect 9723 20961 9735 20964
rect 9677 20955 9735 20961
rect 4356 20896 5764 20924
rect 5810 20884 5816 20936
rect 5868 20924 5874 20936
rect 8021 20927 8079 20933
rect 5868 20896 5913 20924
rect 5868 20884 5874 20896
rect 8021 20893 8033 20927
rect 8067 20924 8079 20927
rect 8864 20924 8892 20955
rect 9766 20952 9772 20964
rect 9824 20952 9830 21004
rect 9950 20992 9956 21004
rect 9911 20964 9956 20992
rect 9950 20952 9956 20964
rect 10008 20952 10014 21004
rect 11256 20992 11284 21091
rect 12526 21088 12532 21140
rect 12584 21128 12590 21140
rect 16758 21128 16764 21140
rect 12584 21100 13676 21128
rect 16719 21100 16764 21128
rect 12584 21088 12590 21100
rect 13648 21060 13676 21100
rect 16758 21088 16764 21100
rect 16816 21088 16822 21140
rect 18046 21088 18052 21140
rect 18104 21128 18110 21140
rect 21269 21131 21327 21137
rect 18104 21100 20024 21128
rect 18104 21088 18110 21100
rect 15746 21060 15752 21072
rect 13648 21032 15752 21060
rect 15746 21020 15752 21032
rect 15804 21060 15810 21072
rect 16942 21060 16948 21072
rect 15804 21032 15884 21060
rect 15804 21020 15810 21032
rect 11793 20995 11851 21001
rect 11793 20992 11805 20995
rect 11256 20964 11805 20992
rect 11793 20961 11805 20964
rect 11839 20961 11851 20995
rect 11793 20955 11851 20961
rect 12526 20952 12532 21004
rect 12584 20992 12590 21004
rect 13078 20992 13084 21004
rect 12584 20964 12629 20992
rect 13039 20964 13084 20992
rect 12584 20952 12590 20964
rect 13078 20952 13084 20964
rect 13136 20952 13142 21004
rect 13725 20995 13783 21001
rect 13725 20992 13737 20995
rect 13188 20964 13737 20992
rect 13188 20924 13216 20964
rect 13725 20961 13737 20964
rect 13771 20961 13783 20995
rect 13725 20955 13783 20961
rect 14185 20995 14243 21001
rect 14185 20961 14197 20995
rect 14231 20992 14243 20995
rect 14642 20992 14648 21004
rect 14231 20964 14648 20992
rect 14231 20961 14243 20964
rect 14185 20955 14243 20961
rect 14642 20952 14648 20964
rect 14700 20952 14706 21004
rect 15856 21001 15884 21032
rect 16408 21032 16948 21060
rect 16408 21001 16436 21032
rect 16942 21020 16948 21032
rect 17000 21060 17006 21072
rect 17000 21032 17908 21060
rect 17000 21020 17006 21032
rect 17880 21004 17908 21032
rect 19334 21020 19340 21072
rect 19392 21060 19398 21072
rect 19613 21063 19671 21069
rect 19392 21032 19564 21060
rect 19392 21020 19398 21032
rect 15841 20995 15899 21001
rect 15841 20961 15853 20995
rect 15887 20961 15899 20995
rect 15841 20955 15899 20961
rect 16393 20995 16451 21001
rect 16393 20961 16405 20995
rect 16439 20961 16451 20995
rect 16393 20955 16451 20961
rect 16758 20952 16764 21004
rect 16816 20992 16822 21004
rect 17037 20995 17095 21001
rect 17037 20992 17049 20995
rect 16816 20964 17049 20992
rect 16816 20952 16822 20964
rect 17037 20961 17049 20964
rect 17083 20961 17095 20995
rect 17037 20955 17095 20961
rect 17497 20995 17555 21001
rect 17497 20961 17509 20995
rect 17543 20961 17555 20995
rect 17497 20955 17555 20961
rect 8067 20896 8892 20924
rect 8956 20896 13216 20924
rect 13449 20927 13507 20933
rect 8067 20893 8079 20896
rect 8021 20887 8079 20893
rect 5350 20816 5356 20868
rect 5408 20856 5414 20868
rect 8956 20856 8984 20896
rect 13449 20893 13461 20927
rect 13495 20924 13507 20927
rect 15102 20924 15108 20936
rect 13495 20896 15108 20924
rect 13495 20893 13507 20896
rect 13449 20887 13507 20893
rect 15102 20884 15108 20896
rect 15160 20884 15166 20936
rect 17512 20924 17540 20955
rect 17862 20952 17868 21004
rect 17920 20992 17926 21004
rect 19536 21001 19564 21032
rect 19613 21029 19625 21063
rect 19659 21060 19671 21063
rect 19886 21060 19892 21072
rect 19659 21032 19892 21060
rect 19659 21029 19671 21032
rect 19613 21023 19671 21029
rect 19886 21020 19892 21032
rect 19944 21020 19950 21072
rect 19996 21069 20024 21100
rect 21269 21097 21281 21131
rect 21315 21128 21327 21131
rect 21450 21128 21456 21140
rect 21315 21100 21456 21128
rect 21315 21097 21327 21100
rect 21269 21091 21327 21097
rect 21450 21088 21456 21100
rect 21508 21088 21514 21140
rect 22094 21128 22100 21140
rect 21652 21100 22100 21128
rect 19981 21063 20039 21069
rect 19981 21029 19993 21063
rect 20027 21029 20039 21063
rect 19981 21023 20039 21029
rect 18509 20995 18567 21001
rect 18509 20992 18521 20995
rect 17920 20964 18521 20992
rect 17920 20952 17926 20964
rect 18509 20961 18521 20964
rect 18555 20961 18567 20995
rect 18509 20955 18567 20961
rect 19429 20995 19487 21001
rect 19429 20961 19441 20995
rect 19475 20961 19487 20995
rect 19429 20955 19487 20961
rect 19521 20995 19579 21001
rect 19521 20961 19533 20995
rect 19567 20992 19579 20995
rect 20162 20992 20168 21004
rect 19567 20964 20168 20992
rect 19567 20961 19579 20964
rect 19521 20955 19579 20961
rect 17954 20924 17960 20936
rect 17512 20896 17960 20924
rect 17954 20884 17960 20896
rect 18012 20884 18018 20936
rect 19150 20884 19156 20936
rect 19208 20924 19214 20936
rect 19245 20927 19303 20933
rect 19245 20924 19257 20927
rect 19208 20896 19257 20924
rect 19208 20884 19214 20896
rect 19245 20893 19257 20896
rect 19291 20893 19303 20927
rect 19444 20924 19472 20955
rect 20162 20952 20168 20964
rect 20220 20952 20226 21004
rect 21082 20992 21088 21004
rect 21043 20964 21088 20992
rect 21082 20952 21088 20964
rect 21140 20952 21146 21004
rect 20254 20924 20260 20936
rect 19444 20896 20260 20924
rect 19245 20887 19303 20893
rect 20254 20884 20260 20896
rect 20312 20924 20318 20936
rect 21542 20924 21548 20936
rect 20312 20896 21548 20924
rect 20312 20884 20318 20896
rect 21542 20884 21548 20896
rect 21600 20884 21606 20936
rect 5408 20828 8984 20856
rect 5408 20816 5414 20828
rect 10870 20816 10876 20868
rect 10928 20856 10934 20868
rect 11977 20859 12035 20865
rect 11977 20856 11989 20859
rect 10928 20828 11989 20856
rect 10928 20816 10934 20828
rect 11977 20825 11989 20828
rect 12023 20825 12035 20859
rect 11977 20819 12035 20825
rect 18693 20859 18751 20865
rect 18693 20825 18705 20859
rect 18739 20856 18751 20859
rect 21652 20856 21680 21100
rect 22094 21088 22100 21100
rect 22152 21088 22158 21140
rect 22922 21088 22928 21140
rect 22980 21128 22986 21140
rect 23106 21128 23112 21140
rect 22980 21100 23112 21128
rect 22980 21088 22986 21100
rect 23106 21088 23112 21100
rect 23164 21088 23170 21140
rect 23198 21088 23204 21140
rect 23256 21128 23262 21140
rect 23256 21100 25084 21128
rect 23256 21088 23262 21100
rect 22204 21032 23520 21060
rect 21818 20992 21824 21004
rect 21779 20964 21824 20992
rect 21818 20952 21824 20964
rect 21876 20992 21882 21004
rect 22204 20992 22232 21032
rect 21876 20964 22232 20992
rect 21876 20952 21882 20964
rect 22278 20952 22284 21004
rect 22336 20992 22342 21004
rect 22373 20995 22431 21001
rect 22373 20992 22385 20995
rect 22336 20964 22385 20992
rect 22336 20952 22342 20964
rect 22373 20961 22385 20964
rect 22419 20992 22431 20995
rect 22830 20992 22836 21004
rect 22419 20964 22836 20992
rect 22419 20961 22431 20964
rect 22373 20955 22431 20961
rect 22830 20952 22836 20964
rect 22888 20952 22894 21004
rect 23492 21001 23520 21032
rect 23566 21020 23572 21072
rect 23624 21060 23630 21072
rect 24118 21060 24124 21072
rect 23624 21032 24124 21060
rect 23624 21020 23630 21032
rect 24118 21020 24124 21032
rect 24176 21060 24182 21072
rect 24596 21069 24624 21100
rect 24489 21063 24547 21069
rect 24489 21060 24501 21063
rect 24176 21032 24501 21060
rect 24176 21020 24182 21032
rect 24489 21029 24501 21032
rect 24535 21029 24547 21063
rect 24489 21023 24547 21029
rect 24581 21063 24639 21069
rect 24581 21029 24593 21063
rect 24627 21029 24639 21063
rect 24946 21060 24952 21072
rect 24907 21032 24952 21060
rect 24581 21023 24639 21029
rect 24946 21020 24952 21032
rect 25004 21020 25010 21072
rect 25056 21060 25084 21100
rect 25130 21088 25136 21140
rect 25188 21128 25194 21140
rect 25593 21131 25651 21137
rect 25593 21128 25605 21131
rect 25188 21100 25605 21128
rect 25188 21088 25194 21100
rect 25593 21097 25605 21100
rect 25639 21097 25651 21131
rect 28626 21128 28632 21140
rect 28587 21100 28632 21128
rect 25593 21091 25651 21097
rect 28626 21088 28632 21100
rect 28684 21088 28690 21140
rect 35710 21088 35716 21140
rect 35768 21128 35774 21140
rect 36446 21128 36452 21140
rect 35768 21100 36452 21128
rect 35768 21088 35774 21100
rect 36446 21088 36452 21100
rect 36504 21088 36510 21140
rect 29086 21060 29092 21072
rect 25056 21032 29092 21060
rect 29086 21020 29092 21032
rect 29144 21020 29150 21072
rect 32030 21060 32036 21072
rect 31220 21032 32036 21060
rect 23293 20995 23351 21001
rect 23293 20961 23305 20995
rect 23339 20992 23351 20995
rect 23477 20995 23535 21001
rect 23339 20964 23428 20992
rect 23339 20961 23351 20964
rect 23293 20955 23351 20961
rect 22554 20924 22560 20936
rect 22515 20896 22560 20924
rect 22554 20884 22560 20896
rect 22612 20884 22618 20936
rect 18739 20828 21680 20856
rect 18739 20825 18751 20828
rect 18693 20819 18751 20825
rect 7466 20748 7472 20800
rect 7524 20788 7530 20800
rect 8202 20788 8208 20800
rect 7524 20760 8208 20788
rect 7524 20748 7530 20760
rect 8202 20748 8208 20760
rect 8260 20748 8266 20800
rect 8938 20788 8944 20800
rect 8899 20760 8944 20788
rect 8938 20748 8944 20760
rect 8996 20748 9002 20800
rect 13078 20748 13084 20800
rect 13136 20788 13142 20800
rect 16206 20788 16212 20800
rect 13136 20760 16212 20788
rect 13136 20748 13142 20760
rect 16206 20748 16212 20760
rect 16264 20788 16270 20800
rect 18708 20788 18736 20819
rect 22002 20816 22008 20868
rect 22060 20856 22066 20868
rect 23400 20856 23428 20964
rect 23477 20961 23489 20995
rect 23523 20961 23535 20995
rect 24394 20992 24400 21004
rect 24355 20964 24400 20992
rect 23477 20955 23535 20961
rect 24394 20952 24400 20964
rect 24452 20952 24458 21004
rect 24670 20952 24676 21004
rect 24728 20992 24734 21004
rect 25409 20995 25467 21001
rect 25409 20992 25421 20995
rect 24728 20964 25421 20992
rect 24728 20952 24734 20964
rect 25409 20961 25421 20964
rect 25455 20961 25467 20995
rect 25409 20955 25467 20961
rect 26513 20995 26571 21001
rect 26513 20961 26525 20995
rect 26559 20961 26571 20995
rect 27614 20992 27620 21004
rect 27575 20964 27620 20992
rect 26513 20955 26571 20961
rect 24210 20924 24216 20936
rect 24171 20896 24216 20924
rect 24210 20884 24216 20896
rect 24268 20884 24274 20936
rect 26528 20856 26556 20955
rect 27614 20952 27620 20964
rect 27672 20952 27678 21004
rect 27706 20952 27712 21004
rect 27764 20992 27770 21004
rect 28169 20995 28227 21001
rect 28169 20992 28181 20995
rect 27764 20964 28181 20992
rect 27764 20952 27770 20964
rect 28169 20961 28181 20964
rect 28215 20961 28227 20995
rect 28350 20992 28356 21004
rect 28311 20964 28356 20992
rect 28169 20955 28227 20961
rect 28350 20952 28356 20964
rect 28408 20952 28414 21004
rect 29270 20992 29276 21004
rect 29231 20964 29276 20992
rect 29270 20952 29276 20964
rect 29328 20952 29334 21004
rect 29822 20992 29828 21004
rect 29783 20964 29828 20992
rect 29822 20952 29828 20964
rect 29880 20952 29886 21004
rect 30282 20992 30288 21004
rect 30243 20964 30288 20992
rect 30282 20952 30288 20964
rect 30340 20952 30346 21004
rect 31220 21001 31248 21032
rect 32030 21020 32036 21032
rect 32088 21020 32094 21072
rect 33502 21060 33508 21072
rect 32324 21032 33508 21060
rect 31113 20995 31171 21001
rect 31113 20961 31125 20995
rect 31159 20961 31171 20995
rect 31113 20955 31171 20961
rect 31205 20995 31263 21001
rect 31205 20961 31217 20995
rect 31251 20961 31263 20995
rect 31205 20955 31263 20961
rect 31573 20995 31631 21001
rect 31573 20961 31585 20995
rect 31619 20992 31631 20995
rect 32324 20992 32352 21032
rect 31619 20964 32352 20992
rect 32401 20995 32459 21001
rect 31619 20961 31631 20964
rect 31573 20955 31631 20961
rect 32401 20961 32413 20995
rect 32447 20992 32459 20995
rect 32674 20992 32680 21004
rect 32447 20964 32680 20992
rect 32447 20961 32459 20964
rect 32401 20955 32459 20961
rect 27525 20927 27583 20933
rect 27525 20893 27537 20927
rect 27571 20893 27583 20927
rect 31128 20924 31156 20955
rect 32674 20952 32680 20964
rect 32732 20952 32738 21004
rect 32784 21001 32812 21032
rect 33502 21020 33508 21032
rect 33560 21020 33566 21072
rect 33778 21020 33784 21072
rect 33836 21060 33842 21072
rect 38654 21060 38660 21072
rect 33836 21032 35112 21060
rect 33836 21020 33842 21032
rect 32769 20995 32827 21001
rect 32769 20961 32781 20995
rect 32815 20961 32827 20995
rect 32769 20955 32827 20961
rect 32858 20952 32864 21004
rect 32916 20992 32922 21004
rect 33410 20992 33416 21004
rect 32916 20964 32961 20992
rect 33371 20964 33416 20992
rect 32916 20952 32922 20964
rect 33410 20952 33416 20964
rect 33468 20952 33474 21004
rect 34330 20992 34336 21004
rect 34291 20964 34336 20992
rect 34330 20952 34336 20964
rect 34388 20952 34394 21004
rect 34701 20995 34759 21001
rect 34701 20961 34713 20995
rect 34747 20992 34759 20995
rect 34974 20992 34980 21004
rect 34747 20964 34980 20992
rect 34747 20961 34759 20964
rect 34701 20955 34759 20961
rect 34974 20952 34980 20964
rect 35032 20952 35038 21004
rect 35084 21001 35112 21032
rect 36832 21032 38660 21060
rect 35069 20995 35127 21001
rect 35069 20961 35081 20995
rect 35115 20961 35127 20995
rect 35069 20955 35127 20961
rect 33042 20924 33048 20936
rect 31128 20896 31616 20924
rect 33003 20896 33048 20924
rect 27525 20887 27583 20893
rect 22060 20828 26556 20856
rect 22060 20816 22066 20828
rect 16264 20760 18736 20788
rect 16264 20748 16270 20760
rect 19886 20748 19892 20800
rect 19944 20788 19950 20800
rect 20070 20788 20076 20800
rect 19944 20760 20076 20788
rect 19944 20748 19950 20760
rect 20070 20748 20076 20760
rect 20128 20748 20134 20800
rect 21450 20748 21456 20800
rect 21508 20788 21514 20800
rect 22738 20788 22744 20800
rect 21508 20760 22744 20788
rect 21508 20748 21514 20760
rect 22738 20748 22744 20760
rect 22796 20748 22802 20800
rect 22830 20748 22836 20800
rect 22888 20788 22894 20800
rect 26605 20791 26663 20797
rect 26605 20788 26617 20791
rect 22888 20760 26617 20788
rect 22888 20748 22894 20760
rect 26605 20757 26617 20760
rect 26651 20757 26663 20791
rect 27540 20788 27568 20887
rect 31588 20868 31616 20896
rect 33042 20884 33048 20896
rect 33100 20884 33106 20936
rect 34514 20924 34520 20936
rect 34475 20896 34520 20924
rect 34514 20884 34520 20896
rect 34572 20884 34578 20936
rect 35084 20924 35112 20955
rect 35342 20952 35348 21004
rect 35400 20992 35406 21004
rect 36832 21001 36860 21032
rect 38654 21020 38660 21032
rect 38712 21020 38718 21072
rect 36081 20995 36139 21001
rect 36081 20992 36093 20995
rect 35400 20964 36093 20992
rect 35400 20952 35406 20964
rect 36081 20961 36093 20964
rect 36127 20961 36139 20995
rect 36081 20955 36139 20961
rect 36817 20995 36875 21001
rect 36817 20961 36829 20995
rect 36863 20961 36875 20995
rect 37826 20992 37832 21004
rect 37787 20964 37832 20992
rect 36817 20955 36875 20961
rect 37826 20952 37832 20964
rect 37884 20952 37890 21004
rect 38562 20992 38568 21004
rect 38523 20964 38568 20992
rect 38562 20952 38568 20964
rect 38620 20952 38626 21004
rect 35434 20924 35440 20936
rect 35084 20896 35440 20924
rect 35434 20884 35440 20896
rect 35492 20884 35498 20936
rect 35894 20884 35900 20936
rect 35952 20924 35958 20936
rect 36909 20927 36967 20933
rect 36909 20924 36921 20927
rect 35952 20896 36921 20924
rect 35952 20884 35958 20896
rect 36909 20893 36921 20896
rect 36955 20893 36967 20927
rect 36909 20887 36967 20893
rect 38470 20884 38476 20936
rect 38528 20924 38534 20936
rect 38657 20927 38715 20933
rect 38657 20924 38669 20927
rect 38528 20896 38669 20924
rect 38528 20884 38534 20896
rect 38657 20893 38669 20896
rect 38703 20893 38715 20927
rect 38657 20887 38715 20893
rect 27614 20816 27620 20868
rect 27672 20856 27678 20868
rect 29365 20859 29423 20865
rect 29365 20856 29377 20859
rect 27672 20828 29377 20856
rect 27672 20816 27678 20828
rect 29365 20825 29377 20828
rect 29411 20825 29423 20859
rect 29365 20819 29423 20825
rect 31570 20816 31576 20868
rect 31628 20816 31634 20868
rect 36357 20859 36415 20865
rect 36357 20825 36369 20859
rect 36403 20856 36415 20859
rect 37182 20856 37188 20868
rect 36403 20828 37188 20856
rect 36403 20825 36415 20828
rect 36357 20819 36415 20825
rect 37182 20816 37188 20828
rect 37240 20816 37246 20868
rect 37734 20816 37740 20868
rect 37792 20856 37798 20868
rect 37921 20859 37979 20865
rect 37921 20856 37933 20859
rect 37792 20828 37933 20856
rect 37792 20816 37798 20828
rect 37921 20825 37933 20828
rect 37967 20825 37979 20859
rect 37921 20819 37979 20825
rect 38102 20788 38108 20800
rect 27540 20760 38108 20788
rect 26605 20751 26663 20757
rect 38102 20748 38108 20760
rect 38160 20748 38166 20800
rect 1104 20698 39836 20720
rect 1104 20646 4246 20698
rect 4298 20646 4310 20698
rect 4362 20646 4374 20698
rect 4426 20646 4438 20698
rect 4490 20646 34966 20698
rect 35018 20646 35030 20698
rect 35082 20646 35094 20698
rect 35146 20646 35158 20698
rect 35210 20646 39836 20698
rect 1104 20624 39836 20646
rect 6454 20584 6460 20596
rect 3896 20556 6460 20584
rect 2958 20448 2964 20460
rect 2700 20420 2964 20448
rect 2700 20389 2728 20420
rect 2958 20408 2964 20420
rect 3016 20408 3022 20460
rect 1857 20383 1915 20389
rect 1857 20349 1869 20383
rect 1903 20349 1915 20383
rect 1857 20343 1915 20349
rect 2685 20383 2743 20389
rect 2685 20349 2697 20383
rect 2731 20349 2743 20383
rect 2685 20343 2743 20349
rect 1872 20312 1900 20343
rect 2774 20340 2780 20392
rect 2832 20380 2838 20392
rect 2869 20383 2927 20389
rect 2869 20380 2881 20383
rect 2832 20352 2881 20380
rect 2832 20340 2838 20352
rect 2869 20349 2881 20352
rect 2915 20349 2927 20383
rect 3234 20380 3240 20392
rect 3195 20352 3240 20380
rect 2869 20343 2927 20349
rect 3234 20340 3240 20352
rect 3292 20340 3298 20392
rect 3896 20389 3924 20556
rect 6454 20544 6460 20556
rect 6512 20584 6518 20596
rect 6512 20556 7788 20584
rect 6512 20544 6518 20556
rect 3973 20519 4031 20525
rect 3973 20485 3985 20519
rect 4019 20516 4031 20519
rect 4614 20516 4620 20528
rect 4019 20488 4620 20516
rect 4019 20485 4031 20488
rect 3973 20479 4031 20485
rect 4614 20476 4620 20488
rect 4672 20476 4678 20528
rect 6822 20516 6828 20528
rect 5736 20488 6828 20516
rect 5442 20448 5448 20460
rect 4448 20420 5448 20448
rect 4448 20389 4476 20420
rect 5442 20408 5448 20420
rect 5500 20408 5506 20460
rect 3881 20383 3939 20389
rect 3881 20349 3893 20383
rect 3927 20349 3939 20383
rect 3881 20343 3939 20349
rect 4433 20383 4491 20389
rect 4433 20349 4445 20383
rect 4479 20349 4491 20383
rect 4433 20343 4491 20349
rect 4709 20383 4767 20389
rect 4709 20349 4721 20383
rect 4755 20380 4767 20383
rect 4755 20352 4844 20380
rect 4755 20349 4767 20352
rect 4709 20343 4767 20349
rect 3252 20312 3280 20340
rect 1872 20284 3280 20312
rect 1949 20247 2007 20253
rect 1949 20213 1961 20247
rect 1995 20244 2007 20247
rect 4816 20244 4844 20352
rect 5350 20340 5356 20392
rect 5408 20380 5414 20392
rect 5736 20389 5764 20488
rect 6822 20476 6828 20488
rect 6880 20476 6886 20528
rect 6273 20451 6331 20457
rect 6273 20417 6285 20451
rect 6319 20448 6331 20451
rect 7101 20451 7159 20457
rect 7101 20448 7113 20451
rect 6319 20420 7113 20448
rect 6319 20417 6331 20420
rect 6273 20411 6331 20417
rect 7101 20417 7113 20420
rect 7147 20417 7159 20451
rect 7101 20411 7159 20417
rect 5537 20383 5595 20389
rect 5537 20380 5549 20383
rect 5408 20352 5549 20380
rect 5408 20340 5414 20352
rect 5537 20349 5549 20352
rect 5583 20349 5595 20383
rect 5537 20343 5595 20349
rect 5721 20383 5779 20389
rect 5721 20349 5733 20383
rect 5767 20349 5779 20383
rect 5721 20343 5779 20349
rect 5813 20383 5871 20389
rect 5813 20349 5825 20383
rect 5859 20380 5871 20383
rect 5902 20380 5908 20392
rect 5859 20352 5908 20380
rect 5859 20349 5871 20352
rect 5813 20343 5871 20349
rect 5902 20340 5908 20352
rect 5960 20340 5966 20392
rect 6822 20380 6828 20392
rect 6783 20352 6828 20380
rect 6822 20340 6828 20352
rect 6880 20340 6886 20392
rect 7760 20380 7788 20556
rect 8110 20544 8116 20596
rect 8168 20584 8174 20596
rect 16390 20584 16396 20596
rect 8168 20556 16396 20584
rect 8168 20544 8174 20556
rect 16390 20544 16396 20556
rect 16448 20544 16454 20596
rect 20254 20544 20260 20596
rect 20312 20584 20318 20596
rect 20312 20556 22416 20584
rect 20312 20544 20318 20556
rect 8386 20476 8392 20528
rect 8444 20516 8450 20528
rect 9033 20519 9091 20525
rect 9033 20516 9045 20519
rect 8444 20488 9045 20516
rect 8444 20476 8450 20488
rect 9033 20485 9045 20488
rect 9079 20485 9091 20519
rect 9033 20479 9091 20485
rect 11440 20488 12848 20516
rect 8018 20408 8024 20460
rect 8076 20448 8082 20460
rect 11440 20457 11468 20488
rect 11425 20451 11483 20457
rect 8076 20420 9536 20448
rect 8076 20408 8082 20420
rect 9508 20389 9536 20420
rect 11425 20417 11437 20451
rect 11471 20417 11483 20451
rect 12529 20451 12587 20457
rect 12529 20448 12541 20451
rect 11425 20411 11483 20417
rect 11532 20420 12541 20448
rect 8941 20383 8999 20389
rect 8941 20380 8953 20383
rect 7760 20352 8953 20380
rect 8941 20349 8953 20352
rect 8987 20349 8999 20383
rect 8941 20343 8999 20349
rect 9493 20383 9551 20389
rect 9493 20349 9505 20383
rect 9539 20349 9551 20383
rect 9858 20380 9864 20392
rect 9819 20352 9864 20380
rect 9493 20343 9551 20349
rect 9858 20340 9864 20352
rect 9916 20340 9922 20392
rect 11330 20340 11336 20392
rect 11388 20380 11394 20392
rect 11532 20380 11560 20420
rect 12529 20417 12541 20420
rect 12575 20417 12587 20451
rect 12820 20448 12848 20488
rect 12894 20476 12900 20528
rect 12952 20516 12958 20528
rect 13265 20519 13323 20525
rect 13265 20516 13277 20519
rect 12952 20488 13277 20516
rect 12952 20476 12958 20488
rect 13265 20485 13277 20488
rect 13311 20485 13323 20519
rect 15286 20516 15292 20528
rect 15247 20488 15292 20516
rect 13265 20479 13323 20485
rect 15286 20476 15292 20488
rect 15344 20476 15350 20528
rect 18230 20516 18236 20528
rect 16960 20488 18236 20516
rect 12820 20420 13032 20448
rect 12529 20411 12587 20417
rect 13004 20392 13032 20420
rect 13078 20408 13084 20460
rect 13136 20448 13142 20460
rect 14553 20451 14611 20457
rect 14553 20448 14565 20451
rect 13136 20420 14565 20448
rect 13136 20408 13142 20420
rect 14553 20417 14565 20420
rect 14599 20417 14611 20451
rect 14553 20411 14611 20417
rect 14734 20408 14740 20460
rect 14792 20448 14798 20460
rect 14918 20448 14924 20460
rect 14792 20420 14924 20448
rect 14792 20408 14798 20420
rect 14918 20408 14924 20420
rect 14976 20408 14982 20460
rect 15102 20408 15108 20460
rect 15160 20448 15166 20460
rect 15160 20420 15332 20448
rect 15160 20408 15166 20420
rect 11698 20380 11704 20392
rect 11388 20352 11560 20380
rect 11659 20352 11704 20380
rect 11388 20340 11394 20352
rect 11698 20340 11704 20352
rect 11756 20340 11762 20392
rect 11885 20383 11943 20389
rect 11885 20349 11897 20383
rect 11931 20380 11943 20383
rect 12710 20380 12716 20392
rect 11931 20352 12716 20380
rect 11931 20349 11943 20352
rect 11885 20343 11943 20349
rect 12710 20340 12716 20352
rect 12768 20340 12774 20392
rect 12986 20380 12992 20392
rect 12947 20352 12992 20380
rect 12986 20340 12992 20352
rect 13044 20340 13050 20392
rect 13357 20383 13415 20389
rect 13357 20349 13369 20383
rect 13403 20380 13415 20383
rect 13906 20380 13912 20392
rect 13403 20352 13912 20380
rect 13403 20349 13415 20352
rect 13357 20343 13415 20349
rect 13906 20340 13912 20352
rect 13964 20340 13970 20392
rect 15013 20383 15071 20389
rect 15013 20349 15025 20383
rect 15059 20380 15071 20383
rect 15194 20380 15200 20392
rect 15059 20352 15200 20380
rect 15059 20349 15071 20352
rect 15013 20343 15071 20349
rect 15194 20340 15200 20352
rect 15252 20340 15258 20392
rect 15304 20389 15332 20420
rect 15289 20383 15347 20389
rect 15289 20349 15301 20383
rect 15335 20349 15347 20383
rect 16298 20380 16304 20392
rect 16259 20352 16304 20380
rect 15289 20343 15347 20349
rect 16298 20340 16304 20352
rect 16356 20340 16362 20392
rect 16577 20383 16635 20389
rect 16577 20349 16589 20383
rect 16623 20380 16635 20383
rect 16666 20380 16672 20392
rect 16623 20352 16672 20380
rect 16623 20349 16635 20352
rect 16577 20343 16635 20349
rect 16666 20340 16672 20352
rect 16724 20340 16730 20392
rect 16960 20389 16988 20488
rect 18230 20476 18236 20488
rect 18288 20476 18294 20528
rect 21082 20516 21088 20528
rect 20995 20488 21088 20516
rect 21082 20476 21088 20488
rect 21140 20516 21146 20528
rect 22002 20516 22008 20528
rect 21140 20488 22008 20516
rect 21140 20476 21146 20488
rect 22002 20476 22008 20488
rect 22060 20476 22066 20528
rect 17494 20448 17500 20460
rect 17455 20420 17500 20448
rect 17494 20408 17500 20420
rect 17552 20408 17558 20460
rect 16945 20383 17003 20389
rect 16945 20349 16957 20383
rect 16991 20349 17003 20383
rect 16945 20343 17003 20349
rect 17313 20383 17371 20389
rect 17313 20349 17325 20383
rect 17359 20380 17371 20383
rect 17402 20380 17408 20392
rect 17359 20352 17408 20380
rect 17359 20349 17371 20352
rect 17313 20343 17371 20349
rect 17402 20340 17408 20352
rect 17460 20340 17466 20392
rect 17589 20383 17647 20389
rect 17589 20349 17601 20383
rect 17635 20380 17647 20383
rect 17770 20380 17776 20392
rect 17635 20352 17776 20380
rect 17635 20349 17647 20352
rect 17589 20343 17647 20349
rect 17770 20340 17776 20352
rect 17828 20340 17834 20392
rect 21100 20389 21128 20476
rect 21542 20448 21548 20460
rect 21455 20420 21548 20448
rect 21542 20408 21548 20420
rect 21600 20448 21606 20460
rect 22388 20448 22416 20556
rect 25590 20544 25596 20596
rect 25648 20584 25654 20596
rect 26694 20584 26700 20596
rect 25648 20556 26700 20584
rect 25648 20544 25654 20556
rect 26694 20544 26700 20556
rect 26752 20544 26758 20596
rect 29641 20587 29699 20593
rect 29641 20553 29653 20587
rect 29687 20584 29699 20587
rect 31110 20584 31116 20596
rect 29687 20556 31116 20584
rect 29687 20553 29699 20556
rect 29641 20547 29699 20553
rect 31110 20544 31116 20556
rect 31168 20584 31174 20596
rect 31168 20556 32076 20584
rect 31168 20544 31174 20556
rect 28166 20476 28172 20528
rect 28224 20516 28230 20528
rect 28261 20519 28319 20525
rect 28261 20516 28273 20519
rect 28224 20488 28273 20516
rect 28224 20476 28230 20488
rect 28261 20485 28273 20488
rect 28307 20485 28319 20519
rect 28261 20479 28319 20485
rect 22554 20448 22560 20460
rect 21600 20420 22324 20448
rect 22388 20420 22560 20448
rect 21600 20408 21606 20420
rect 21085 20383 21143 20389
rect 21085 20349 21097 20383
rect 21131 20349 21143 20383
rect 21266 20380 21272 20392
rect 21227 20352 21272 20380
rect 21085 20343 21143 20349
rect 21266 20340 21272 20352
rect 21324 20340 21330 20392
rect 21358 20340 21364 20392
rect 21416 20380 21422 20392
rect 22097 20383 22155 20389
rect 22097 20380 22109 20383
rect 21416 20352 22109 20380
rect 21416 20340 21422 20352
rect 22097 20349 22109 20352
rect 22143 20349 22155 20383
rect 22097 20343 22155 20349
rect 10873 20315 10931 20321
rect 7760 20284 8524 20312
rect 7760 20244 7788 20284
rect 8386 20244 8392 20256
rect 1995 20216 7788 20244
rect 8347 20216 8392 20244
rect 1995 20213 2007 20216
rect 1949 20207 2007 20213
rect 8386 20204 8392 20216
rect 8444 20204 8450 20256
rect 8496 20244 8524 20284
rect 10873 20281 10885 20315
rect 10919 20312 10931 20315
rect 13538 20312 13544 20324
rect 10919 20284 13544 20312
rect 10919 20281 10931 20284
rect 10873 20275 10931 20281
rect 13538 20272 13544 20284
rect 13596 20272 13602 20324
rect 18414 20312 18420 20324
rect 18375 20284 18420 20312
rect 18414 20272 18420 20284
rect 18472 20272 18478 20324
rect 22296 20312 22324 20420
rect 22554 20408 22560 20420
rect 22612 20448 22618 20460
rect 24489 20451 24547 20457
rect 24489 20448 24501 20451
rect 22612 20420 24501 20448
rect 22612 20408 22618 20420
rect 24489 20417 24501 20420
rect 24535 20417 24547 20451
rect 26237 20451 26295 20457
rect 24489 20411 24547 20417
rect 25332 20420 26096 20448
rect 22830 20380 22836 20392
rect 22791 20352 22836 20380
rect 22830 20340 22836 20352
rect 22888 20340 22894 20392
rect 22922 20340 22928 20392
rect 22980 20380 22986 20392
rect 23017 20383 23075 20389
rect 23017 20380 23029 20383
rect 22980 20352 23029 20380
rect 22980 20340 22986 20352
rect 23017 20349 23029 20352
rect 23063 20349 23075 20383
rect 23017 20343 23075 20349
rect 23474 20340 23480 20392
rect 23532 20380 23538 20392
rect 23661 20383 23719 20389
rect 23661 20380 23673 20383
rect 23532 20352 23673 20380
rect 23532 20340 23538 20352
rect 23661 20349 23673 20352
rect 23707 20349 23719 20383
rect 23661 20343 23719 20349
rect 24394 20340 24400 20392
rect 24452 20380 24458 20392
rect 25332 20389 25360 20420
rect 24765 20383 24823 20389
rect 24765 20380 24777 20383
rect 24452 20352 24777 20380
rect 24452 20340 24458 20352
rect 24765 20349 24777 20352
rect 24811 20349 24823 20383
rect 24765 20343 24823 20349
rect 25317 20383 25375 20389
rect 25317 20349 25329 20383
rect 25363 20349 25375 20383
rect 25958 20380 25964 20392
rect 25919 20352 25964 20380
rect 25317 20343 25375 20349
rect 25958 20340 25964 20352
rect 26016 20340 26022 20392
rect 26068 20380 26096 20420
rect 26237 20417 26249 20451
rect 26283 20448 26295 20451
rect 27614 20448 27620 20460
rect 26283 20420 27620 20448
rect 26283 20417 26295 20420
rect 26237 20411 26295 20417
rect 27614 20408 27620 20420
rect 27672 20408 27678 20460
rect 28276 20448 28304 20479
rect 30653 20451 30711 20457
rect 28276 20420 30604 20448
rect 27522 20380 27528 20392
rect 26068 20352 27528 20380
rect 27522 20340 27528 20352
rect 27580 20340 27586 20392
rect 28442 20380 28448 20392
rect 28403 20352 28448 20380
rect 28442 20340 28448 20352
rect 28500 20340 28506 20392
rect 28534 20340 28540 20392
rect 28592 20380 28598 20392
rect 29641 20383 29699 20389
rect 28592 20352 28637 20380
rect 28592 20340 28598 20352
rect 29641 20349 29653 20383
rect 29687 20380 29699 20383
rect 29733 20383 29791 20389
rect 29733 20380 29745 20383
rect 29687 20352 29745 20380
rect 29687 20349 29699 20352
rect 29641 20343 29699 20349
rect 29733 20349 29745 20352
rect 29779 20349 29791 20383
rect 29733 20343 29791 20349
rect 30282 20340 30288 20392
rect 30340 20380 30346 20392
rect 30377 20383 30435 20389
rect 30377 20380 30389 20383
rect 30340 20352 30389 20380
rect 30340 20340 30346 20352
rect 30377 20349 30389 20352
rect 30423 20349 30435 20383
rect 30576 20380 30604 20420
rect 30653 20417 30665 20451
rect 30699 20448 30711 20451
rect 31294 20448 31300 20460
rect 30699 20420 31300 20448
rect 30699 20417 30711 20420
rect 30653 20411 30711 20417
rect 31294 20408 31300 20420
rect 31352 20408 31358 20460
rect 32048 20457 32076 20556
rect 33042 20544 33048 20596
rect 33100 20584 33106 20596
rect 33100 20556 36308 20584
rect 33100 20544 33106 20556
rect 33597 20519 33655 20525
rect 33597 20485 33609 20519
rect 33643 20516 33655 20519
rect 35342 20516 35348 20528
rect 33643 20488 35348 20516
rect 33643 20485 33655 20488
rect 33597 20479 33655 20485
rect 35342 20476 35348 20488
rect 35400 20476 35406 20528
rect 36280 20516 36308 20556
rect 36280 20488 36400 20516
rect 32033 20451 32091 20457
rect 32033 20417 32045 20451
rect 32079 20448 32091 20451
rect 34241 20451 34299 20457
rect 32079 20420 32536 20448
rect 32079 20417 32091 20420
rect 32033 20411 32091 20417
rect 32508 20389 32536 20420
rect 34241 20417 34253 20451
rect 34287 20448 34299 20451
rect 34514 20448 34520 20460
rect 34287 20420 34520 20448
rect 34287 20417 34299 20420
rect 34241 20411 34299 20417
rect 34514 20408 34520 20420
rect 34572 20408 34578 20460
rect 35713 20451 35771 20457
rect 35713 20417 35725 20451
rect 35759 20448 35771 20451
rect 35894 20448 35900 20460
rect 35759 20420 35900 20448
rect 35759 20417 35771 20420
rect 35713 20411 35771 20417
rect 35894 20408 35900 20420
rect 35952 20408 35958 20460
rect 32493 20383 32551 20389
rect 30576 20352 31340 20380
rect 30377 20343 30435 20349
rect 24412 20312 24440 20340
rect 25498 20312 25504 20324
rect 22296 20284 24440 20312
rect 25459 20284 25504 20312
rect 25498 20272 25504 20284
rect 25556 20272 25562 20324
rect 31312 20312 31340 20352
rect 32493 20349 32505 20383
rect 32539 20349 32551 20383
rect 32493 20343 32551 20349
rect 33781 20383 33839 20389
rect 33781 20349 33793 20383
rect 33827 20380 33839 20383
rect 34054 20380 34060 20392
rect 33827 20352 34060 20380
rect 33827 20349 33839 20352
rect 33781 20343 33839 20349
rect 34054 20340 34060 20352
rect 34112 20340 34118 20392
rect 34149 20383 34207 20389
rect 34149 20349 34161 20383
rect 34195 20380 34207 20383
rect 35250 20380 35256 20392
rect 34195 20352 35256 20380
rect 34195 20349 34207 20352
rect 34149 20343 34207 20349
rect 35250 20340 35256 20352
rect 35308 20340 35314 20392
rect 35805 20383 35863 20389
rect 35805 20349 35817 20383
rect 35851 20380 35863 20383
rect 36078 20380 36084 20392
rect 35851 20352 36084 20380
rect 35851 20349 35863 20352
rect 35805 20343 35863 20349
rect 36078 20340 36084 20352
rect 36136 20340 36142 20392
rect 36173 20383 36231 20389
rect 36173 20349 36185 20383
rect 36219 20380 36231 20383
rect 36262 20380 36268 20392
rect 36219 20352 36268 20380
rect 36219 20349 36231 20352
rect 36173 20343 36231 20349
rect 36262 20340 36268 20352
rect 36320 20340 36326 20392
rect 36372 20389 36400 20488
rect 37734 20448 37740 20460
rect 37695 20420 37740 20448
rect 37734 20408 37740 20420
rect 37792 20408 37798 20460
rect 36357 20383 36415 20389
rect 36357 20349 36369 20383
rect 36403 20349 36415 20383
rect 36357 20343 36415 20349
rect 36725 20383 36783 20389
rect 36725 20349 36737 20383
rect 36771 20349 36783 20383
rect 36725 20343 36783 20349
rect 31312 20284 33824 20312
rect 33796 20256 33824 20284
rect 34514 20272 34520 20324
rect 34572 20312 34578 20324
rect 36740 20312 36768 20343
rect 37274 20340 37280 20392
rect 37332 20380 37338 20392
rect 37461 20383 37519 20389
rect 37461 20380 37473 20383
rect 37332 20352 37473 20380
rect 37332 20340 37338 20352
rect 37461 20349 37473 20352
rect 37507 20349 37519 20383
rect 37461 20343 37519 20349
rect 34572 20284 36768 20312
rect 34572 20272 34578 20284
rect 13814 20244 13820 20256
rect 8496 20216 13820 20244
rect 13814 20204 13820 20216
rect 13872 20204 13878 20256
rect 16114 20244 16120 20256
rect 16075 20216 16120 20244
rect 16114 20204 16120 20216
rect 16172 20204 16178 20256
rect 16206 20204 16212 20256
rect 16264 20244 16270 20256
rect 17773 20247 17831 20253
rect 17773 20244 17785 20247
rect 16264 20216 17785 20244
rect 16264 20204 16270 20216
rect 17773 20213 17785 20216
rect 17819 20213 17831 20247
rect 17773 20207 17831 20213
rect 19426 20204 19432 20256
rect 19484 20244 19490 20256
rect 19705 20247 19763 20253
rect 19705 20244 19717 20247
rect 19484 20216 19717 20244
rect 19484 20204 19490 20216
rect 19705 20213 19717 20216
rect 19751 20213 19763 20247
rect 19705 20207 19763 20213
rect 22097 20247 22155 20253
rect 22097 20213 22109 20247
rect 22143 20244 22155 20247
rect 22186 20244 22192 20256
rect 22143 20216 22192 20244
rect 22143 20213 22155 20216
rect 22097 20207 22155 20213
rect 22186 20204 22192 20216
rect 22244 20204 22250 20256
rect 23842 20204 23848 20256
rect 23900 20244 23906 20256
rect 23900 20216 23945 20244
rect 23900 20204 23906 20216
rect 24302 20204 24308 20256
rect 24360 20244 24366 20256
rect 25130 20244 25136 20256
rect 24360 20216 25136 20244
rect 24360 20204 24366 20216
rect 25130 20204 25136 20216
rect 25188 20204 25194 20256
rect 26326 20204 26332 20256
rect 26384 20244 26390 20256
rect 27341 20247 27399 20253
rect 27341 20244 27353 20247
rect 26384 20216 27353 20244
rect 26384 20204 26390 20216
rect 27341 20213 27353 20216
rect 27387 20213 27399 20247
rect 27341 20207 27399 20213
rect 28629 20247 28687 20253
rect 28629 20213 28641 20247
rect 28675 20244 28687 20247
rect 29730 20244 29736 20256
rect 28675 20216 29736 20244
rect 28675 20213 28687 20216
rect 28629 20207 28687 20213
rect 29730 20204 29736 20216
rect 29788 20204 29794 20256
rect 29825 20247 29883 20253
rect 29825 20213 29837 20247
rect 29871 20244 29883 20247
rect 32490 20244 32496 20256
rect 29871 20216 32496 20244
rect 29871 20213 29883 20216
rect 29825 20207 29883 20213
rect 32490 20204 32496 20216
rect 32548 20204 32554 20256
rect 32674 20244 32680 20256
rect 32587 20216 32680 20244
rect 32674 20204 32680 20216
rect 32732 20244 32738 20256
rect 33042 20244 33048 20256
rect 32732 20216 33048 20244
rect 32732 20204 32738 20216
rect 33042 20204 33048 20216
rect 33100 20204 33106 20256
rect 33778 20204 33784 20256
rect 33836 20204 33842 20256
rect 38102 20204 38108 20256
rect 38160 20244 38166 20256
rect 38841 20247 38899 20253
rect 38841 20244 38853 20247
rect 38160 20216 38853 20244
rect 38160 20204 38166 20216
rect 38841 20213 38853 20216
rect 38887 20213 38899 20247
rect 38841 20207 38899 20213
rect 1104 20154 39836 20176
rect 1104 20102 19606 20154
rect 19658 20102 19670 20154
rect 19722 20102 19734 20154
rect 19786 20102 19798 20154
rect 19850 20102 39836 20154
rect 1104 20080 39836 20102
rect 11330 20040 11336 20052
rect 5000 20012 11336 20040
rect 3053 19975 3111 19981
rect 3053 19941 3065 19975
rect 3099 19972 3111 19975
rect 3234 19972 3240 19984
rect 3099 19944 3240 19972
rect 3099 19941 3111 19944
rect 3053 19935 3111 19941
rect 3234 19932 3240 19944
rect 3292 19932 3298 19984
rect 1394 19904 1400 19916
rect 1355 19876 1400 19904
rect 1394 19864 1400 19876
rect 1452 19864 1458 19916
rect 3878 19864 3884 19916
rect 3936 19904 3942 19916
rect 5000 19913 5028 20012
rect 11330 20000 11336 20012
rect 11388 20000 11394 20052
rect 11698 20000 11704 20052
rect 11756 20040 11762 20052
rect 11977 20043 12035 20049
rect 11977 20040 11989 20043
rect 11756 20012 11989 20040
rect 11756 20000 11762 20012
rect 11977 20009 11989 20012
rect 12023 20009 12035 20043
rect 12802 20040 12808 20052
rect 12763 20012 12808 20040
rect 11977 20003 12035 20009
rect 12802 20000 12808 20012
rect 12860 20000 12866 20052
rect 12986 20000 12992 20052
rect 13044 20040 13050 20052
rect 13354 20040 13360 20052
rect 13044 20012 13360 20040
rect 13044 20000 13050 20012
rect 13354 20000 13360 20012
rect 13412 20040 13418 20052
rect 16206 20040 16212 20052
rect 13412 20012 16212 20040
rect 13412 20000 13418 20012
rect 16206 20000 16212 20012
rect 16264 20000 16270 20052
rect 17402 20040 17408 20052
rect 17363 20012 17408 20040
rect 17402 20000 17408 20012
rect 17460 20000 17466 20052
rect 17494 20000 17500 20052
rect 17552 20040 17558 20052
rect 19150 20040 19156 20052
rect 17552 20012 19156 20040
rect 17552 20000 17558 20012
rect 19150 20000 19156 20012
rect 19208 20040 19214 20052
rect 19208 20012 19472 20040
rect 19208 20000 19214 20012
rect 5810 19972 5816 19984
rect 5276 19944 5816 19972
rect 5276 19913 5304 19944
rect 5810 19932 5816 19944
rect 5868 19932 5874 19984
rect 19242 19972 19248 19984
rect 15396 19944 17080 19972
rect 4065 19907 4123 19913
rect 4065 19904 4077 19907
rect 3936 19876 4077 19904
rect 3936 19864 3942 19876
rect 4065 19873 4077 19876
rect 4111 19873 4123 19907
rect 4065 19867 4123 19873
rect 4985 19907 5043 19913
rect 4985 19873 4997 19907
rect 5031 19873 5043 19907
rect 4985 19867 5043 19873
rect 5261 19907 5319 19913
rect 5261 19873 5273 19907
rect 5307 19873 5319 19907
rect 5534 19904 5540 19916
rect 5495 19876 5540 19904
rect 5261 19867 5319 19873
rect 5534 19864 5540 19876
rect 5592 19864 5598 19916
rect 5626 19864 5632 19916
rect 5684 19904 5690 19916
rect 5997 19907 6055 19913
rect 5997 19904 6009 19907
rect 5684 19876 6009 19904
rect 5684 19864 5690 19876
rect 5997 19873 6009 19876
rect 6043 19873 6055 19907
rect 5997 19867 6055 19873
rect 6641 19907 6699 19913
rect 6641 19873 6653 19907
rect 6687 19904 6699 19907
rect 6687 19876 6776 19904
rect 6687 19873 6699 19876
rect 6641 19867 6699 19873
rect 1670 19836 1676 19848
rect 1631 19808 1676 19836
rect 1670 19796 1676 19808
rect 1728 19796 1734 19848
rect 5350 19836 5356 19848
rect 5311 19808 5356 19836
rect 5350 19796 5356 19808
rect 5408 19796 5414 19848
rect 3418 19660 3424 19712
rect 3476 19700 3482 19712
rect 4157 19703 4215 19709
rect 4157 19700 4169 19703
rect 3476 19672 4169 19700
rect 3476 19660 3482 19672
rect 4157 19669 4169 19672
rect 4203 19700 4215 19703
rect 6748 19700 6776 19876
rect 6914 19864 6920 19916
rect 6972 19904 6978 19916
rect 7745 19907 7803 19913
rect 6972 19876 7604 19904
rect 6972 19864 6978 19876
rect 6822 19796 6828 19848
rect 6880 19836 6886 19848
rect 7466 19836 7472 19848
rect 6880 19808 7472 19836
rect 6880 19796 6886 19808
rect 7466 19796 7472 19808
rect 7524 19796 7530 19848
rect 7576 19836 7604 19876
rect 7745 19873 7757 19907
rect 7791 19904 7803 19907
rect 8938 19904 8944 19916
rect 7791 19876 8944 19904
rect 7791 19873 7803 19876
rect 7745 19867 7803 19873
rect 8938 19864 8944 19876
rect 8996 19864 9002 19916
rect 9122 19904 9128 19916
rect 9035 19876 9128 19904
rect 9122 19864 9128 19876
rect 9180 19904 9186 19916
rect 9677 19907 9735 19913
rect 9677 19904 9689 19907
rect 9180 19876 9689 19904
rect 9180 19864 9186 19876
rect 9677 19873 9689 19876
rect 9723 19873 9735 19907
rect 9677 19867 9735 19873
rect 10873 19907 10931 19913
rect 10873 19873 10885 19907
rect 10919 19904 10931 19907
rect 11514 19904 11520 19916
rect 10919 19876 11520 19904
rect 10919 19873 10931 19876
rect 10873 19867 10931 19873
rect 11514 19864 11520 19876
rect 11572 19864 11578 19916
rect 12894 19904 12900 19916
rect 12855 19876 12900 19904
rect 12894 19864 12900 19876
rect 12952 19864 12958 19916
rect 13357 19907 13415 19913
rect 13357 19873 13369 19907
rect 13403 19873 13415 19907
rect 13538 19904 13544 19916
rect 13499 19876 13544 19904
rect 13357 19867 13415 19873
rect 8202 19836 8208 19848
rect 7576 19808 8208 19836
rect 8202 19796 8208 19808
rect 8260 19836 8266 19848
rect 9030 19836 9036 19848
rect 8260 19808 9036 19836
rect 8260 19796 8266 19808
rect 9030 19796 9036 19808
rect 9088 19796 9094 19848
rect 9306 19796 9312 19848
rect 9364 19836 9370 19848
rect 10410 19836 10416 19848
rect 9364 19808 10416 19836
rect 9364 19796 9370 19808
rect 10410 19796 10416 19808
rect 10468 19796 10474 19848
rect 10594 19836 10600 19848
rect 10555 19808 10600 19836
rect 10594 19796 10600 19808
rect 10652 19796 10658 19848
rect 13372 19836 13400 19867
rect 13538 19864 13544 19876
rect 13596 19864 13602 19916
rect 14458 19904 14464 19916
rect 14419 19876 14464 19904
rect 14458 19864 14464 19876
rect 14516 19904 14522 19916
rect 14516 19876 14596 19904
rect 14516 19864 14522 19876
rect 13446 19836 13452 19848
rect 13372 19808 13452 19836
rect 13446 19796 13452 19808
rect 13504 19796 13510 19848
rect 14568 19836 14596 19876
rect 14642 19864 14648 19916
rect 14700 19904 14706 19916
rect 15102 19904 15108 19916
rect 14700 19876 15108 19904
rect 14700 19864 14706 19876
rect 15102 19864 15108 19876
rect 15160 19904 15166 19916
rect 15289 19907 15347 19913
rect 15289 19904 15301 19907
rect 15160 19876 15301 19904
rect 15160 19864 15166 19876
rect 15289 19873 15301 19876
rect 15335 19873 15347 19907
rect 15289 19867 15347 19873
rect 15396 19836 15424 19944
rect 15473 19907 15531 19913
rect 15473 19873 15485 19907
rect 15519 19873 15531 19907
rect 16942 19904 16948 19916
rect 16903 19876 16948 19904
rect 15473 19867 15531 19873
rect 14568 19808 15424 19836
rect 15488 19768 15516 19867
rect 16942 19864 16948 19876
rect 17000 19864 17006 19916
rect 17052 19836 17080 19944
rect 19168 19944 19248 19972
rect 17129 19907 17187 19913
rect 17129 19873 17141 19907
rect 17175 19904 17187 19907
rect 17494 19904 17500 19916
rect 17175 19876 17500 19904
rect 17175 19873 17187 19876
rect 17129 19867 17187 19873
rect 17494 19864 17500 19876
rect 17552 19864 17558 19916
rect 17586 19864 17592 19916
rect 17644 19904 17650 19916
rect 19168 19913 19196 19944
rect 19242 19932 19248 19944
rect 19300 19932 19306 19984
rect 17681 19907 17739 19913
rect 17681 19904 17693 19907
rect 17644 19876 17693 19904
rect 17644 19864 17650 19876
rect 17681 19873 17693 19876
rect 17727 19873 17739 19907
rect 17681 19867 17739 19873
rect 18049 19907 18107 19913
rect 18049 19873 18061 19907
rect 18095 19873 18107 19907
rect 18049 19867 18107 19873
rect 19153 19907 19211 19913
rect 19153 19873 19165 19907
rect 19199 19873 19211 19907
rect 19334 19904 19340 19916
rect 19295 19876 19340 19904
rect 19153 19867 19211 19873
rect 17770 19836 17776 19848
rect 17052 19808 17776 19836
rect 17770 19796 17776 19808
rect 17828 19836 17834 19848
rect 18064 19836 18092 19867
rect 19334 19864 19340 19876
rect 19392 19864 19398 19916
rect 19444 19904 19472 20012
rect 20916 20012 21956 20040
rect 19613 19907 19671 19913
rect 19613 19904 19625 19907
rect 19444 19876 19625 19904
rect 19613 19873 19625 19876
rect 19659 19873 19671 19907
rect 20254 19904 20260 19916
rect 20215 19876 20260 19904
rect 19613 19867 19671 19873
rect 20254 19864 20260 19876
rect 20312 19864 20318 19916
rect 20916 19913 20944 20012
rect 21928 19972 21956 20012
rect 22002 20000 22008 20052
rect 22060 20040 22066 20052
rect 22281 20043 22339 20049
rect 22281 20040 22293 20043
rect 22060 20012 22293 20040
rect 22060 20000 22066 20012
rect 22281 20009 22293 20012
rect 22327 20009 22339 20043
rect 25958 20040 25964 20052
rect 22281 20003 22339 20009
rect 25056 20012 25964 20040
rect 25056 19972 25084 20012
rect 25958 20000 25964 20012
rect 26016 20000 26022 20052
rect 26510 20000 26516 20052
rect 26568 20040 26574 20052
rect 26789 20043 26847 20049
rect 26789 20040 26801 20043
rect 26568 20012 26801 20040
rect 26568 20000 26574 20012
rect 26789 20009 26801 20012
rect 26835 20009 26847 20043
rect 26789 20003 26847 20009
rect 27430 20000 27436 20052
rect 27488 20040 27494 20052
rect 30006 20040 30012 20052
rect 27488 20012 30012 20040
rect 27488 20000 27494 20012
rect 30006 20000 30012 20012
rect 30064 20000 30070 20052
rect 31772 20012 34652 20040
rect 31772 19972 31800 20012
rect 34330 19972 34336 19984
rect 21928 19944 25084 19972
rect 25148 19944 31800 19972
rect 33336 19944 34336 19972
rect 25148 19916 25176 19944
rect 20901 19907 20959 19913
rect 20901 19873 20913 19907
rect 20947 19873 20959 19907
rect 20901 19867 20959 19873
rect 21634 19864 21640 19916
rect 21692 19904 21698 19916
rect 21818 19904 21824 19916
rect 21692 19876 21824 19904
rect 21692 19864 21698 19876
rect 21818 19864 21824 19876
rect 21876 19904 21882 19916
rect 23017 19907 23075 19913
rect 23017 19904 23029 19907
rect 21876 19876 23029 19904
rect 21876 19864 21882 19876
rect 23017 19873 23029 19876
rect 23063 19873 23075 19907
rect 23017 19867 23075 19873
rect 24673 19907 24731 19913
rect 24673 19873 24685 19907
rect 24719 19904 24731 19907
rect 25130 19904 25136 19916
rect 24719 19876 24808 19904
rect 25043 19876 25136 19904
rect 24719 19873 24731 19876
rect 24673 19867 24731 19873
rect 18969 19839 19027 19845
rect 18969 19836 18981 19839
rect 17828 19808 18981 19836
rect 17828 19796 17834 19808
rect 18969 19805 18981 19808
rect 19015 19805 19027 19839
rect 18969 19799 19027 19805
rect 21177 19839 21235 19845
rect 21177 19805 21189 19839
rect 21223 19836 21235 19839
rect 21223 19808 24072 19836
rect 21223 19805 21235 19808
rect 21177 19799 21235 19805
rect 11716 19740 15516 19768
rect 8110 19700 8116 19712
rect 4203 19672 8116 19700
rect 4203 19669 4215 19672
rect 4157 19663 4215 19669
rect 8110 19660 8116 19672
rect 8168 19660 8174 19712
rect 9769 19703 9827 19709
rect 9769 19669 9781 19703
rect 9815 19700 9827 19703
rect 9858 19700 9864 19712
rect 9815 19672 9864 19700
rect 9815 19669 9827 19672
rect 9769 19663 9827 19669
rect 9858 19660 9864 19672
rect 9916 19700 9922 19712
rect 11716 19700 11744 19740
rect 16022 19728 16028 19780
rect 16080 19768 16086 19780
rect 19426 19768 19432 19780
rect 16080 19740 19432 19768
rect 16080 19728 16086 19740
rect 19426 19728 19432 19740
rect 19484 19728 19490 19780
rect 23842 19728 23848 19780
rect 23900 19768 23906 19780
rect 24044 19777 24072 19808
rect 23937 19771 23995 19777
rect 23937 19768 23949 19771
rect 23900 19740 23949 19768
rect 23900 19728 23906 19740
rect 23937 19737 23949 19740
rect 23983 19737 23995 19771
rect 23937 19731 23995 19737
rect 24029 19771 24087 19777
rect 24029 19737 24041 19771
rect 24075 19737 24087 19771
rect 24029 19731 24087 19737
rect 24670 19728 24676 19780
rect 24728 19768 24734 19780
rect 24780 19768 24808 19876
rect 25130 19864 25136 19876
rect 25188 19864 25194 19916
rect 25406 19904 25412 19916
rect 25367 19876 25412 19904
rect 25406 19864 25412 19876
rect 25464 19864 25470 19916
rect 25498 19864 25504 19916
rect 25556 19904 25562 19916
rect 25593 19907 25651 19913
rect 25593 19904 25605 19907
rect 25556 19876 25605 19904
rect 25556 19864 25562 19876
rect 25593 19873 25605 19876
rect 25639 19873 25651 19907
rect 25593 19867 25651 19873
rect 26513 19907 26571 19913
rect 26513 19873 26525 19907
rect 26559 19904 26571 19907
rect 26602 19904 26608 19916
rect 26559 19876 26608 19904
rect 26559 19873 26571 19876
rect 26513 19867 26571 19873
rect 26602 19864 26608 19876
rect 26660 19864 26666 19916
rect 26697 19907 26755 19913
rect 26697 19873 26709 19907
rect 26743 19873 26755 19907
rect 26697 19867 26755 19873
rect 26712 19836 26740 19867
rect 27430 19864 27436 19916
rect 27488 19904 27494 19916
rect 27525 19907 27583 19913
rect 27525 19904 27537 19907
rect 27488 19876 27537 19904
rect 27488 19864 27494 19876
rect 27525 19873 27537 19876
rect 27571 19873 27583 19907
rect 27525 19867 27583 19873
rect 28445 19907 28503 19913
rect 28445 19873 28457 19907
rect 28491 19904 28503 19907
rect 28534 19904 28540 19916
rect 28491 19876 28540 19904
rect 28491 19873 28503 19876
rect 28445 19867 28503 19873
rect 28534 19864 28540 19876
rect 28592 19864 28598 19916
rect 28994 19904 29000 19916
rect 28955 19876 29000 19904
rect 28994 19864 29000 19876
rect 29052 19904 29058 19916
rect 29733 19907 29791 19913
rect 29733 19904 29745 19907
rect 29052 19876 29745 19904
rect 29052 19864 29058 19876
rect 29733 19873 29745 19876
rect 29779 19873 29791 19907
rect 29733 19867 29791 19873
rect 30837 19907 30895 19913
rect 30837 19873 30849 19907
rect 30883 19904 30895 19907
rect 32030 19904 32036 19916
rect 30883 19876 32036 19904
rect 30883 19873 30895 19876
rect 30837 19867 30895 19873
rect 32030 19864 32036 19876
rect 32088 19864 32094 19916
rect 33336 19913 33364 19944
rect 34330 19932 34336 19944
rect 34388 19932 34394 19984
rect 34624 19981 34652 20012
rect 35618 20000 35624 20052
rect 35676 20000 35682 20052
rect 34609 19975 34667 19981
rect 34609 19941 34621 19975
rect 34655 19941 34667 19975
rect 35636 19972 35664 20000
rect 34609 19935 34667 19941
rect 35360 19944 35664 19972
rect 32953 19907 33011 19913
rect 32953 19873 32965 19907
rect 32999 19904 33011 19907
rect 33321 19907 33379 19913
rect 32999 19876 33272 19904
rect 32999 19873 33011 19876
rect 32953 19867 33011 19873
rect 27614 19836 27620 19848
rect 26712 19808 27620 19836
rect 27614 19796 27620 19808
rect 27672 19796 27678 19848
rect 29086 19836 29092 19848
rect 29047 19808 29092 19836
rect 29086 19796 29092 19808
rect 29144 19796 29150 19848
rect 24728 19740 30696 19768
rect 24728 19728 24734 19740
rect 30668 19712 30696 19740
rect 14642 19700 14648 19712
rect 9916 19672 11744 19700
rect 14603 19672 14648 19700
rect 9916 19660 9922 19672
rect 14642 19660 14648 19672
rect 14700 19660 14706 19712
rect 14826 19660 14832 19712
rect 14884 19700 14890 19712
rect 15565 19703 15623 19709
rect 15565 19700 15577 19703
rect 14884 19672 15577 19700
rect 14884 19660 14890 19672
rect 15565 19669 15577 19672
rect 15611 19669 15623 19703
rect 15565 19663 15623 19669
rect 16114 19660 16120 19712
rect 16172 19700 16178 19712
rect 18690 19700 18696 19712
rect 16172 19672 18696 19700
rect 16172 19660 16178 19672
rect 18690 19660 18696 19672
rect 18748 19660 18754 19712
rect 22554 19660 22560 19712
rect 22612 19700 22618 19712
rect 22922 19700 22928 19712
rect 22612 19672 22928 19700
rect 22612 19660 22618 19672
rect 22922 19660 22928 19672
rect 22980 19700 22986 19712
rect 23201 19703 23259 19709
rect 23201 19700 23213 19703
rect 22980 19672 23213 19700
rect 22980 19660 22986 19672
rect 23201 19669 23213 19672
rect 23247 19669 23259 19703
rect 23201 19663 23259 19669
rect 25958 19660 25964 19712
rect 26016 19700 26022 19712
rect 27062 19700 27068 19712
rect 26016 19672 27068 19700
rect 26016 19660 26022 19672
rect 27062 19660 27068 19672
rect 27120 19660 27126 19712
rect 27706 19700 27712 19712
rect 27667 19672 27712 19700
rect 27706 19660 27712 19672
rect 27764 19660 27770 19712
rect 28445 19703 28503 19709
rect 28445 19669 28457 19703
rect 28491 19700 28503 19703
rect 29638 19700 29644 19712
rect 28491 19672 29644 19700
rect 28491 19669 28503 19672
rect 28445 19663 28503 19669
rect 29638 19660 29644 19672
rect 29696 19660 29702 19712
rect 29822 19700 29828 19712
rect 29783 19672 29828 19700
rect 29822 19660 29828 19672
rect 29880 19660 29886 19712
rect 30650 19660 30656 19712
rect 30708 19700 30714 19712
rect 31021 19703 31079 19709
rect 31021 19700 31033 19703
rect 30708 19672 31033 19700
rect 30708 19660 30714 19672
rect 31021 19669 31033 19672
rect 31067 19669 31079 19703
rect 31021 19663 31079 19669
rect 32030 19660 32036 19712
rect 32088 19700 32094 19712
rect 32769 19703 32827 19709
rect 32769 19700 32781 19703
rect 32088 19672 32781 19700
rect 32088 19660 32094 19672
rect 32769 19669 32781 19672
rect 32815 19669 32827 19703
rect 33244 19700 33272 19876
rect 33321 19873 33333 19907
rect 33367 19873 33379 19907
rect 33502 19904 33508 19916
rect 33463 19876 33508 19904
rect 33321 19867 33379 19873
rect 33502 19864 33508 19876
rect 33560 19864 33566 19916
rect 33962 19904 33968 19916
rect 33923 19876 33968 19904
rect 33962 19864 33968 19876
rect 34020 19864 34026 19916
rect 35360 19913 35388 19944
rect 35161 19907 35219 19913
rect 35161 19873 35173 19907
rect 35207 19873 35219 19907
rect 35161 19867 35219 19873
rect 35345 19907 35403 19913
rect 35345 19873 35357 19907
rect 35391 19873 35403 19907
rect 35345 19867 35403 19873
rect 35176 19836 35204 19867
rect 35434 19864 35440 19916
rect 35492 19904 35498 19916
rect 35621 19907 35679 19913
rect 35492 19876 35537 19904
rect 35492 19864 35498 19876
rect 35621 19873 35633 19907
rect 35667 19873 35679 19907
rect 35621 19867 35679 19873
rect 35897 19907 35955 19913
rect 35897 19873 35909 19907
rect 35943 19873 35955 19907
rect 35897 19867 35955 19873
rect 35526 19836 35532 19848
rect 35176 19808 35532 19836
rect 35526 19796 35532 19808
rect 35584 19796 35590 19848
rect 33962 19728 33968 19780
rect 34020 19768 34026 19780
rect 35636 19768 35664 19867
rect 34020 19740 35664 19768
rect 34020 19728 34026 19740
rect 35342 19700 35348 19712
rect 33244 19672 35348 19700
rect 32769 19663 32827 19669
rect 35342 19660 35348 19672
rect 35400 19700 35406 19712
rect 35912 19700 35940 19867
rect 35986 19864 35992 19916
rect 36044 19904 36050 19916
rect 36909 19907 36967 19913
rect 36909 19904 36921 19907
rect 36044 19876 36921 19904
rect 36044 19864 36050 19876
rect 36909 19873 36921 19876
rect 36955 19873 36967 19907
rect 38102 19904 38108 19916
rect 38063 19876 38108 19904
rect 36909 19867 36967 19873
rect 38102 19864 38108 19876
rect 38160 19864 38166 19916
rect 38470 19904 38476 19916
rect 38431 19876 38476 19904
rect 38470 19864 38476 19876
rect 38528 19864 38534 19916
rect 38654 19904 38660 19916
rect 38615 19876 38660 19904
rect 38654 19864 38660 19876
rect 38712 19864 38718 19916
rect 35400 19672 35940 19700
rect 35400 19660 35406 19672
rect 36998 19660 37004 19712
rect 37056 19700 37062 19712
rect 37093 19703 37151 19709
rect 37093 19700 37105 19703
rect 37056 19672 37105 19700
rect 37056 19660 37062 19672
rect 37093 19669 37105 19672
rect 37139 19669 37151 19703
rect 37093 19663 37151 19669
rect 1104 19610 39836 19632
rect 1104 19558 4246 19610
rect 4298 19558 4310 19610
rect 4362 19558 4374 19610
rect 4426 19558 4438 19610
rect 4490 19558 34966 19610
rect 35018 19558 35030 19610
rect 35082 19558 35094 19610
rect 35146 19558 35158 19610
rect 35210 19558 39836 19610
rect 1104 19536 39836 19558
rect 1581 19499 1639 19505
rect 1581 19465 1593 19499
rect 1627 19496 1639 19499
rect 1670 19496 1676 19508
rect 1627 19468 1676 19496
rect 1627 19465 1639 19468
rect 1581 19459 1639 19465
rect 1670 19456 1676 19468
rect 1728 19456 1734 19508
rect 4062 19456 4068 19508
rect 4120 19496 4126 19508
rect 9766 19496 9772 19508
rect 4120 19468 9772 19496
rect 4120 19456 4126 19468
rect 9766 19456 9772 19468
rect 9824 19456 9830 19508
rect 11330 19456 11336 19508
rect 11388 19496 11394 19508
rect 11517 19499 11575 19505
rect 11517 19496 11529 19499
rect 11388 19468 11529 19496
rect 11388 19456 11394 19468
rect 11517 19465 11529 19468
rect 11563 19465 11575 19499
rect 11517 19459 11575 19465
rect 15194 19456 15200 19508
rect 15252 19496 15258 19508
rect 15565 19499 15623 19505
rect 15565 19496 15577 19499
rect 15252 19468 15577 19496
rect 15252 19456 15258 19468
rect 15565 19465 15577 19468
rect 15611 19465 15623 19499
rect 15565 19459 15623 19465
rect 16666 19456 16672 19508
rect 16724 19496 16730 19508
rect 18046 19496 18052 19508
rect 16724 19468 18052 19496
rect 16724 19456 16730 19468
rect 18046 19456 18052 19468
rect 18104 19456 18110 19508
rect 27062 19456 27068 19508
rect 27120 19496 27126 19508
rect 27120 19468 28396 19496
rect 27120 19456 27126 19468
rect 3050 19428 3056 19440
rect 1688 19400 3056 19428
rect 1489 19295 1547 19301
rect 1489 19261 1501 19295
rect 1535 19292 1547 19295
rect 1688 19292 1716 19400
rect 3050 19388 3056 19400
rect 3108 19388 3114 19440
rect 7282 19388 7288 19440
rect 7340 19428 7346 19440
rect 9306 19428 9312 19440
rect 7340 19400 9312 19428
rect 7340 19388 7346 19400
rect 9306 19388 9312 19400
rect 9364 19388 9370 19440
rect 24026 19428 24032 19440
rect 23987 19400 24032 19428
rect 24026 19388 24032 19400
rect 24084 19388 24090 19440
rect 28368 19428 28396 19468
rect 28534 19456 28540 19508
rect 28592 19496 28598 19508
rect 31481 19499 31539 19505
rect 31481 19496 31493 19499
rect 28592 19468 31493 19496
rect 28592 19456 28598 19468
rect 31481 19465 31493 19468
rect 31527 19465 31539 19499
rect 31481 19459 31539 19465
rect 34790 19456 34796 19508
rect 34848 19496 34854 19508
rect 35069 19499 35127 19505
rect 35069 19496 35081 19499
rect 34848 19468 35081 19496
rect 34848 19456 34854 19468
rect 35069 19465 35081 19468
rect 35115 19496 35127 19499
rect 35526 19496 35532 19508
rect 35115 19468 35532 19496
rect 35115 19465 35127 19468
rect 35069 19459 35127 19465
rect 35526 19456 35532 19468
rect 35584 19456 35590 19508
rect 28368 19400 28580 19428
rect 7834 19360 7840 19372
rect 7795 19332 7840 19360
rect 7834 19320 7840 19332
rect 7892 19320 7898 19372
rect 9416 19332 9720 19360
rect 1535 19264 1716 19292
rect 2121 19295 2179 19301
rect 1535 19261 1547 19264
rect 1489 19255 1547 19261
rect 2121 19261 2133 19295
rect 2167 19261 2179 19295
rect 2121 19255 2179 19261
rect 3145 19295 3203 19301
rect 3145 19261 3157 19295
rect 3191 19292 3203 19295
rect 3234 19292 3240 19304
rect 3191 19264 3240 19292
rect 3191 19261 3203 19264
rect 3145 19255 3203 19261
rect 2148 19224 2176 19255
rect 3234 19252 3240 19264
rect 3292 19252 3298 19304
rect 3326 19252 3332 19304
rect 3384 19292 3390 19304
rect 3694 19292 3700 19304
rect 3384 19264 3429 19292
rect 3655 19264 3700 19292
rect 3384 19252 3390 19264
rect 3694 19252 3700 19264
rect 3752 19252 3758 19304
rect 4246 19292 4252 19304
rect 4159 19264 4252 19292
rect 4246 19252 4252 19264
rect 4304 19292 4310 19304
rect 4890 19292 4896 19304
rect 4304 19264 4896 19292
rect 4304 19252 4310 19264
rect 4890 19252 4896 19264
rect 4948 19252 4954 19304
rect 5445 19295 5503 19301
rect 5445 19261 5457 19295
rect 5491 19292 5503 19295
rect 5534 19292 5540 19304
rect 5491 19264 5540 19292
rect 5491 19261 5503 19264
rect 5445 19255 5503 19261
rect 5534 19252 5540 19264
rect 5592 19252 5598 19304
rect 5810 19292 5816 19304
rect 5771 19264 5816 19292
rect 5810 19252 5816 19264
rect 5868 19252 5874 19304
rect 7098 19292 7104 19304
rect 7059 19264 7104 19292
rect 7098 19252 7104 19264
rect 7156 19252 7162 19304
rect 7653 19295 7711 19301
rect 7653 19261 7665 19295
rect 7699 19261 7711 19295
rect 7653 19255 7711 19261
rect 2774 19224 2780 19236
rect 2148 19196 2780 19224
rect 2774 19184 2780 19196
rect 2832 19184 2838 19236
rect 5994 19224 6000 19236
rect 5955 19196 6000 19224
rect 5994 19184 6000 19196
rect 6052 19184 6058 19236
rect 7668 19224 7696 19255
rect 7742 19252 7748 19304
rect 7800 19292 7806 19304
rect 7800 19264 7845 19292
rect 7800 19252 7806 19264
rect 8294 19252 8300 19304
rect 8352 19292 8358 19304
rect 8481 19295 8539 19301
rect 8481 19292 8493 19295
rect 8352 19264 8493 19292
rect 8352 19252 8358 19264
rect 8481 19261 8493 19264
rect 8527 19292 8539 19295
rect 9122 19292 9128 19304
rect 8527 19264 9128 19292
rect 8527 19261 8539 19264
rect 8481 19255 8539 19261
rect 9122 19252 9128 19264
rect 9180 19252 9186 19304
rect 9309 19295 9367 19301
rect 9309 19261 9321 19295
rect 9355 19292 9367 19295
rect 9416 19292 9444 19332
rect 9582 19292 9588 19304
rect 9355 19264 9444 19292
rect 9543 19264 9588 19292
rect 9355 19261 9367 19264
rect 9309 19255 9367 19261
rect 9582 19252 9588 19264
rect 9640 19252 9646 19304
rect 9692 19292 9720 19332
rect 10594 19320 10600 19372
rect 10652 19360 10658 19372
rect 13722 19360 13728 19372
rect 10652 19332 11560 19360
rect 13683 19332 13728 19360
rect 10652 19320 10658 19332
rect 9950 19292 9956 19304
rect 9692 19264 9956 19292
rect 9950 19252 9956 19264
rect 10008 19252 10014 19304
rect 10962 19292 10968 19304
rect 10923 19264 10968 19292
rect 10962 19252 10968 19264
rect 11020 19252 11026 19304
rect 11425 19295 11483 19301
rect 11425 19292 11437 19295
rect 11072 19264 11437 19292
rect 7668 19196 7788 19224
rect 7760 19168 7788 19196
rect 2317 19159 2375 19165
rect 2317 19125 2329 19159
rect 2363 19156 2375 19159
rect 3050 19156 3056 19168
rect 2363 19128 3056 19156
rect 2363 19125 2375 19128
rect 2317 19119 2375 19125
rect 3050 19116 3056 19128
rect 3108 19116 3114 19168
rect 3970 19116 3976 19168
rect 4028 19156 4034 19168
rect 4065 19159 4123 19165
rect 4065 19156 4077 19159
rect 4028 19128 4077 19156
rect 4028 19116 4034 19128
rect 4065 19125 4077 19128
rect 4111 19156 4123 19159
rect 7558 19156 7564 19168
rect 4111 19128 7564 19156
rect 4111 19125 4123 19128
rect 4065 19119 4123 19125
rect 7558 19116 7564 19128
rect 7616 19116 7622 19168
rect 7742 19156 7748 19168
rect 7655 19128 7748 19156
rect 7742 19116 7748 19128
rect 7800 19156 7806 19168
rect 8386 19156 8392 19168
rect 7800 19128 8392 19156
rect 7800 19116 7806 19128
rect 8386 19116 8392 19128
rect 8444 19156 8450 19168
rect 11072 19156 11100 19264
rect 11425 19261 11437 19264
rect 11471 19261 11483 19295
rect 11425 19255 11483 19261
rect 8444 19128 11100 19156
rect 11532 19156 11560 19332
rect 13722 19320 13728 19332
rect 13780 19320 13786 19372
rect 14826 19360 14832 19372
rect 14108 19332 14832 19360
rect 12250 19292 12256 19304
rect 12211 19264 12256 19292
rect 12250 19252 12256 19264
rect 12308 19252 12314 19304
rect 12802 19292 12808 19304
rect 12763 19264 12808 19292
rect 12802 19252 12808 19264
rect 12860 19252 12866 19304
rect 13170 19292 13176 19304
rect 13131 19264 13176 19292
rect 13170 19252 13176 19264
rect 13228 19252 13234 19304
rect 13541 19295 13599 19301
rect 13541 19261 13553 19295
rect 13587 19292 13599 19295
rect 14108 19292 14136 19332
rect 14826 19320 14832 19332
rect 14884 19320 14890 19372
rect 21266 19360 21272 19372
rect 16316 19332 16620 19360
rect 13587 19264 14136 19292
rect 14185 19295 14243 19301
rect 13587 19261 13599 19264
rect 13541 19255 13599 19261
rect 14185 19261 14197 19295
rect 14231 19261 14243 19295
rect 14185 19255 14243 19261
rect 14461 19295 14519 19301
rect 14461 19261 14473 19295
rect 14507 19292 14519 19295
rect 16206 19292 16212 19304
rect 14507 19264 16212 19292
rect 14507 19261 14519 19264
rect 14461 19255 14519 19261
rect 12434 19184 12440 19236
rect 12492 19224 12498 19236
rect 14200 19224 14228 19255
rect 16206 19252 16212 19264
rect 16264 19252 16270 19304
rect 16316 19301 16344 19332
rect 16301 19295 16359 19301
rect 16301 19261 16313 19295
rect 16347 19261 16359 19295
rect 16301 19255 16359 19261
rect 16393 19295 16451 19301
rect 16393 19261 16405 19295
rect 16439 19292 16451 19295
rect 16482 19292 16488 19304
rect 16439 19264 16488 19292
rect 16439 19261 16451 19264
rect 16393 19255 16451 19261
rect 16482 19252 16488 19264
rect 16540 19252 16546 19304
rect 16592 19292 16620 19332
rect 17972 19332 19748 19360
rect 16666 19292 16672 19304
rect 16592 19264 16672 19292
rect 16666 19252 16672 19264
rect 16724 19252 16730 19304
rect 17313 19295 17371 19301
rect 17313 19261 17325 19295
rect 17359 19261 17371 19295
rect 17313 19255 17371 19261
rect 17405 19295 17463 19301
rect 17405 19261 17417 19295
rect 17451 19292 17463 19295
rect 17972 19292 18000 19332
rect 17451 19264 18000 19292
rect 18049 19295 18107 19301
rect 17451 19261 17463 19264
rect 17405 19255 17463 19261
rect 18049 19261 18061 19295
rect 18095 19292 18107 19295
rect 18138 19292 18144 19304
rect 18095 19264 18144 19292
rect 18095 19261 18107 19264
rect 18049 19255 18107 19261
rect 12492 19196 14228 19224
rect 12492 19184 12498 19196
rect 15194 19184 15200 19236
rect 15252 19224 15258 19236
rect 16853 19227 16911 19233
rect 16853 19224 16865 19227
rect 15252 19196 16865 19224
rect 15252 19184 15258 19196
rect 16853 19193 16865 19196
rect 16899 19193 16911 19227
rect 17328 19224 17356 19255
rect 18138 19252 18144 19264
rect 18196 19252 18202 19304
rect 18690 19292 18696 19304
rect 18651 19264 18696 19292
rect 18690 19252 18696 19264
rect 18748 19252 18754 19304
rect 18966 19292 18972 19304
rect 18927 19264 18972 19292
rect 18966 19252 18972 19264
rect 19024 19252 19030 19304
rect 19058 19252 19064 19304
rect 19116 19292 19122 19304
rect 19720 19292 19748 19332
rect 20732 19332 21272 19360
rect 20732 19292 20760 19332
rect 21266 19320 21272 19332
rect 21324 19320 21330 19372
rect 21542 19320 21548 19372
rect 21600 19360 21606 19372
rect 22557 19363 22615 19369
rect 22557 19360 22569 19363
rect 21600 19332 22569 19360
rect 21600 19320 21606 19332
rect 22557 19329 22569 19332
rect 22603 19360 22615 19363
rect 28442 19360 28448 19372
rect 22603 19332 28448 19360
rect 22603 19329 22615 19332
rect 22557 19323 22615 19329
rect 28442 19320 28448 19332
rect 28500 19320 28506 19372
rect 28552 19360 28580 19400
rect 28552 19332 29316 19360
rect 19116 19264 19656 19292
rect 19720 19264 20760 19292
rect 20809 19295 20867 19301
rect 19116 19252 19122 19264
rect 19628 19224 19656 19264
rect 20809 19261 20821 19295
rect 20855 19292 20867 19295
rect 20898 19292 20904 19304
rect 20855 19264 20904 19292
rect 20855 19261 20867 19264
rect 20809 19255 20867 19261
rect 20898 19252 20904 19264
rect 20956 19252 20962 19304
rect 21082 19252 21088 19304
rect 21140 19292 21146 19304
rect 22649 19295 22707 19301
rect 22649 19292 22661 19295
rect 21140 19264 22661 19292
rect 21140 19252 21146 19264
rect 22649 19261 22661 19264
rect 22695 19261 22707 19295
rect 22649 19255 22707 19261
rect 22741 19295 22799 19301
rect 22741 19261 22753 19295
rect 22787 19261 22799 19295
rect 22741 19255 22799 19261
rect 22756 19224 22784 19255
rect 23842 19252 23848 19304
rect 23900 19292 23906 19304
rect 23937 19295 23995 19301
rect 23937 19292 23949 19295
rect 23900 19264 23949 19292
rect 23900 19252 23906 19264
rect 23937 19261 23949 19264
rect 23983 19261 23995 19295
rect 24670 19292 24676 19304
rect 24631 19264 24676 19292
rect 23937 19255 23995 19261
rect 24670 19252 24676 19264
rect 24728 19252 24734 19304
rect 25130 19292 25136 19304
rect 25091 19264 25136 19292
rect 25130 19252 25136 19264
rect 25188 19252 25194 19304
rect 25406 19292 25412 19304
rect 25319 19264 25412 19292
rect 25406 19252 25412 19264
rect 25464 19252 25470 19304
rect 25498 19252 25504 19304
rect 25556 19292 25562 19304
rect 25593 19295 25651 19301
rect 25593 19292 25605 19295
rect 25556 19264 25605 19292
rect 25556 19252 25562 19264
rect 25593 19261 25605 19264
rect 25639 19261 25651 19295
rect 26326 19292 26332 19304
rect 26287 19264 26332 19292
rect 25593 19255 25651 19261
rect 26326 19252 26332 19264
rect 26384 19252 26390 19304
rect 27062 19292 27068 19304
rect 27023 19264 27068 19292
rect 27062 19252 27068 19264
rect 27120 19252 27126 19304
rect 27154 19252 27160 19304
rect 27212 19292 27218 19304
rect 27341 19295 27399 19301
rect 27341 19292 27353 19295
rect 27212 19264 27353 19292
rect 27212 19252 27218 19264
rect 27341 19261 27353 19264
rect 27387 19261 27399 19295
rect 27341 19255 27399 19261
rect 28721 19295 28779 19301
rect 28721 19261 28733 19295
rect 28767 19292 28779 19295
rect 28994 19292 29000 19304
rect 28767 19264 29000 19292
rect 28767 19261 28779 19264
rect 28721 19255 28779 19261
rect 28994 19252 29000 19264
rect 29052 19252 29058 19304
rect 29288 19301 29316 19332
rect 29454 19320 29460 19372
rect 29512 19360 29518 19372
rect 29549 19363 29607 19369
rect 29549 19360 29561 19363
rect 29512 19332 29561 19360
rect 29512 19320 29518 19332
rect 29549 19329 29561 19332
rect 29595 19329 29607 19363
rect 29549 19323 29607 19329
rect 32490 19320 32496 19372
rect 32548 19360 32554 19372
rect 33962 19360 33968 19372
rect 32548 19332 33968 19360
rect 32548 19320 32554 19332
rect 33962 19320 33968 19332
rect 34020 19360 34026 19372
rect 34020 19332 34100 19360
rect 34020 19320 34026 19332
rect 29273 19295 29331 19301
rect 29273 19261 29285 19295
rect 29319 19292 29331 19295
rect 30006 19292 30012 19304
rect 29319 19264 30012 19292
rect 29319 19261 29331 19264
rect 29273 19255 29331 19261
rect 30006 19252 30012 19264
rect 30064 19252 30070 19304
rect 31665 19295 31723 19301
rect 31665 19261 31677 19295
rect 31711 19292 31723 19295
rect 31846 19292 31852 19304
rect 31711 19264 31852 19292
rect 31711 19261 31723 19264
rect 31665 19255 31723 19261
rect 31846 19252 31852 19264
rect 31904 19252 31910 19304
rect 32030 19292 32036 19304
rect 31991 19264 32036 19292
rect 32030 19252 32036 19264
rect 32088 19252 32094 19304
rect 32401 19295 32459 19301
rect 32401 19261 32413 19295
rect 32447 19292 32459 19295
rect 32950 19292 32956 19304
rect 32447 19264 32956 19292
rect 32447 19261 32459 19264
rect 32401 19255 32459 19261
rect 32950 19252 32956 19264
rect 33008 19252 33014 19304
rect 34072 19301 34100 19332
rect 34514 19320 34520 19372
rect 34572 19360 34578 19372
rect 34572 19332 35664 19360
rect 34572 19320 34578 19332
rect 35636 19301 35664 19332
rect 36078 19320 36084 19372
rect 36136 19360 36142 19372
rect 37274 19360 37280 19372
rect 36136 19332 37280 19360
rect 36136 19320 36142 19332
rect 33873 19295 33931 19301
rect 33873 19261 33885 19295
rect 33919 19261 33931 19295
rect 33873 19255 33931 19261
rect 34057 19295 34115 19301
rect 34057 19261 34069 19295
rect 34103 19261 34115 19295
rect 34057 19255 34115 19261
rect 34885 19295 34943 19301
rect 34885 19261 34897 19295
rect 34931 19261 34943 19295
rect 34885 19255 34943 19261
rect 35621 19295 35679 19301
rect 35621 19261 35633 19295
rect 35667 19261 35679 19295
rect 35621 19255 35679 19261
rect 36173 19295 36231 19301
rect 36173 19261 36185 19295
rect 36219 19292 36231 19295
rect 36262 19292 36268 19304
rect 36219 19264 36268 19292
rect 36219 19261 36231 19264
rect 36173 19255 36231 19261
rect 23198 19224 23204 19236
rect 17328 19196 18828 19224
rect 19628 19196 22784 19224
rect 23159 19196 23204 19224
rect 16853 19187 16911 19193
rect 12069 19159 12127 19165
rect 12069 19156 12081 19159
rect 11532 19128 12081 19156
rect 8444 19116 8450 19128
rect 12069 19125 12081 19128
rect 12115 19125 12127 19159
rect 12069 19119 12127 19125
rect 18233 19159 18291 19165
rect 18233 19125 18245 19159
rect 18279 19156 18291 19159
rect 18414 19156 18420 19168
rect 18279 19128 18420 19156
rect 18279 19125 18291 19128
rect 18233 19119 18291 19125
rect 18414 19116 18420 19128
rect 18472 19116 18478 19168
rect 18800 19156 18828 19196
rect 23198 19184 23204 19196
rect 23256 19184 23262 19236
rect 25424 19224 25452 19252
rect 26050 19224 26056 19236
rect 25424 19196 26056 19224
rect 26050 19184 26056 19196
rect 26108 19184 26114 19236
rect 33134 19184 33140 19236
rect 33192 19224 33198 19236
rect 33888 19224 33916 19255
rect 34900 19224 34928 19255
rect 36262 19252 36268 19264
rect 36320 19252 36326 19304
rect 36924 19301 36952 19332
rect 37274 19320 37280 19332
rect 37332 19320 37338 19372
rect 36909 19295 36967 19301
rect 36909 19261 36921 19295
rect 36955 19261 36967 19295
rect 37182 19292 37188 19304
rect 37143 19264 37188 19292
rect 36909 19255 36967 19261
rect 37182 19252 37188 19264
rect 37240 19252 37246 19304
rect 38378 19252 38384 19304
rect 38436 19292 38442 19304
rect 38565 19295 38623 19301
rect 38565 19292 38577 19295
rect 38436 19264 38577 19292
rect 38436 19252 38442 19264
rect 38565 19261 38577 19264
rect 38611 19261 38623 19295
rect 38565 19255 38623 19261
rect 33192 19196 34928 19224
rect 35728 19196 36308 19224
rect 33192 19184 33198 19196
rect 19242 19156 19248 19168
rect 18800 19128 19248 19156
rect 19242 19116 19248 19128
rect 19300 19116 19306 19168
rect 19334 19116 19340 19168
rect 19392 19156 19398 19168
rect 20073 19159 20131 19165
rect 20073 19156 20085 19159
rect 19392 19128 20085 19156
rect 19392 19116 19398 19128
rect 20073 19125 20085 19128
rect 20119 19125 20131 19159
rect 20073 19119 20131 19125
rect 21818 19116 21824 19168
rect 21876 19156 21882 19168
rect 22922 19156 22928 19168
rect 21876 19128 22928 19156
rect 21876 19116 21882 19128
rect 22922 19116 22928 19128
rect 22980 19156 22986 19168
rect 26513 19159 26571 19165
rect 26513 19156 26525 19159
rect 22980 19128 26525 19156
rect 22980 19116 22986 19128
rect 26513 19125 26525 19128
rect 26559 19125 26571 19159
rect 26513 19119 26571 19125
rect 27614 19116 27620 19168
rect 27672 19156 27678 19168
rect 28074 19156 28080 19168
rect 27672 19128 28080 19156
rect 27672 19116 27678 19128
rect 28074 19116 28080 19128
rect 28132 19116 28138 19168
rect 29638 19116 29644 19168
rect 29696 19156 29702 19168
rect 30653 19159 30711 19165
rect 30653 19156 30665 19159
rect 29696 19128 30665 19156
rect 29696 19116 29702 19128
rect 30653 19125 30665 19128
rect 30699 19125 30711 19159
rect 30653 19119 30711 19125
rect 33873 19159 33931 19165
rect 33873 19125 33885 19159
rect 33919 19156 33931 19159
rect 35728 19156 35756 19196
rect 33919 19128 35756 19156
rect 33919 19125 33931 19128
rect 33873 19119 33931 19125
rect 35802 19116 35808 19168
rect 35860 19156 35866 19168
rect 35897 19159 35955 19165
rect 35897 19156 35909 19159
rect 35860 19128 35909 19156
rect 35860 19116 35866 19128
rect 35897 19125 35909 19128
rect 35943 19125 35955 19159
rect 36280 19156 36308 19196
rect 38930 19156 38936 19168
rect 36280 19128 38936 19156
rect 35897 19119 35955 19125
rect 38930 19116 38936 19128
rect 38988 19116 38994 19168
rect 1104 19066 39836 19088
rect 1104 19014 19606 19066
rect 19658 19014 19670 19066
rect 19722 19014 19734 19066
rect 19786 19014 19798 19066
rect 19850 19014 39836 19066
rect 1104 18992 39836 19014
rect 3234 18912 3240 18964
rect 3292 18952 3298 18964
rect 4801 18955 4859 18961
rect 4801 18952 4813 18955
rect 3292 18924 4813 18952
rect 3292 18912 3298 18924
rect 2774 18884 2780 18896
rect 2608 18856 2780 18884
rect 2608 18825 2636 18856
rect 2774 18844 2780 18856
rect 2832 18884 2838 18896
rect 3418 18884 3424 18896
rect 2832 18856 3424 18884
rect 2832 18844 2838 18856
rect 3418 18844 3424 18856
rect 3476 18844 3482 18896
rect 3528 18828 3556 18924
rect 4801 18921 4813 18924
rect 4847 18952 4859 18955
rect 5626 18952 5632 18964
rect 4847 18924 5632 18952
rect 4847 18921 4859 18924
rect 4801 18915 4859 18921
rect 5626 18912 5632 18924
rect 5684 18912 5690 18964
rect 9766 18912 9772 18964
rect 9824 18912 9830 18964
rect 9858 18912 9864 18964
rect 9916 18952 9922 18964
rect 9916 18924 9996 18952
rect 9916 18912 9922 18924
rect 8757 18887 8815 18893
rect 8757 18884 8769 18887
rect 4632 18856 8769 18884
rect 2593 18819 2651 18825
rect 2593 18785 2605 18819
rect 2639 18785 2651 18819
rect 2593 18779 2651 18785
rect 2685 18819 2743 18825
rect 2685 18785 2697 18819
rect 2731 18785 2743 18819
rect 2866 18816 2872 18828
rect 2827 18788 2872 18816
rect 2685 18779 2743 18785
rect 2700 18748 2728 18779
rect 2866 18776 2872 18788
rect 2924 18776 2930 18828
rect 2958 18776 2964 18828
rect 3016 18816 3022 18828
rect 3237 18819 3295 18825
rect 3237 18816 3249 18819
rect 3016 18788 3249 18816
rect 3016 18776 3022 18788
rect 3237 18785 3249 18788
rect 3283 18816 3295 18819
rect 3326 18816 3332 18828
rect 3283 18788 3332 18816
rect 3283 18785 3295 18788
rect 3237 18779 3295 18785
rect 3326 18776 3332 18788
rect 3384 18776 3390 18828
rect 3510 18776 3516 18828
rect 3568 18816 3574 18828
rect 4632 18825 4660 18856
rect 8757 18853 8769 18856
rect 8803 18853 8815 18887
rect 8757 18847 8815 18853
rect 4617 18819 4675 18825
rect 3568 18788 3661 18816
rect 3568 18776 3574 18788
rect 4617 18785 4629 18819
rect 4663 18785 4675 18819
rect 4617 18779 4675 18785
rect 5445 18819 5503 18825
rect 5445 18785 5457 18819
rect 5491 18816 5503 18819
rect 5718 18816 5724 18828
rect 5491 18788 5580 18816
rect 5679 18788 5724 18816
rect 5491 18785 5503 18788
rect 5445 18779 5503 18785
rect 4246 18748 4252 18760
rect 2700 18720 4252 18748
rect 4246 18708 4252 18720
rect 4304 18708 4310 18760
rect 5350 18640 5356 18692
rect 5408 18680 5414 18692
rect 5552 18680 5580 18788
rect 5718 18776 5724 18788
rect 5776 18776 5782 18828
rect 5994 18776 6000 18828
rect 6052 18816 6058 18828
rect 6089 18819 6147 18825
rect 6089 18816 6101 18819
rect 6052 18788 6101 18816
rect 6052 18776 6058 18788
rect 6089 18785 6101 18788
rect 6135 18785 6147 18819
rect 6089 18779 6147 18785
rect 6825 18819 6883 18825
rect 6825 18785 6837 18819
rect 6871 18816 6883 18819
rect 7742 18816 7748 18828
rect 6871 18788 7748 18816
rect 6871 18785 6883 18788
rect 6825 18779 6883 18785
rect 7742 18776 7748 18788
rect 7800 18776 7806 18828
rect 8205 18819 8263 18825
rect 8205 18785 8217 18819
rect 8251 18816 8263 18819
rect 8294 18816 8300 18828
rect 8251 18788 8300 18816
rect 8251 18785 8263 18788
rect 8205 18779 8263 18785
rect 8294 18776 8300 18788
rect 8352 18776 8358 18828
rect 8665 18819 8723 18825
rect 8665 18785 8677 18819
rect 8711 18785 8723 18819
rect 8665 18779 8723 18785
rect 5902 18748 5908 18760
rect 5863 18720 5908 18748
rect 5902 18708 5908 18720
rect 5960 18708 5966 18760
rect 7837 18751 7895 18757
rect 7837 18717 7849 18751
rect 7883 18748 7895 18751
rect 8570 18748 8576 18760
rect 7883 18720 8576 18748
rect 7883 18717 7895 18720
rect 7837 18711 7895 18717
rect 8570 18708 8576 18720
rect 8628 18708 8634 18760
rect 8680 18680 8708 18779
rect 8772 18748 8800 18847
rect 9582 18844 9588 18896
rect 9640 18884 9646 18896
rect 9674 18884 9680 18896
rect 9640 18856 9680 18884
rect 9640 18844 9646 18856
rect 9674 18844 9680 18856
rect 9732 18844 9738 18896
rect 9784 18825 9812 18912
rect 9968 18884 9996 18924
rect 10042 18912 10048 18964
rect 10100 18952 10106 18964
rect 14734 18952 14740 18964
rect 10100 18924 14740 18952
rect 10100 18912 10106 18924
rect 14734 18912 14740 18924
rect 14792 18912 14798 18964
rect 15562 18952 15568 18964
rect 15523 18924 15568 18952
rect 15562 18912 15568 18924
rect 15620 18912 15626 18964
rect 16206 18912 16212 18964
rect 16264 18952 16270 18964
rect 23198 18952 23204 18964
rect 16264 18924 23204 18952
rect 16264 18912 16270 18924
rect 23198 18912 23204 18924
rect 23256 18912 23262 18964
rect 26694 18952 26700 18964
rect 26655 18924 26700 18952
rect 26694 18912 26700 18924
rect 26752 18912 26758 18964
rect 27890 18912 27896 18964
rect 27948 18952 27954 18964
rect 34146 18952 34152 18964
rect 27948 18924 34152 18952
rect 27948 18912 27954 18924
rect 34146 18912 34152 18924
rect 34204 18912 34210 18964
rect 36740 18924 38516 18952
rect 10229 18887 10287 18893
rect 10229 18884 10241 18887
rect 9968 18856 10241 18884
rect 10229 18853 10241 18856
rect 10275 18853 10287 18887
rect 10229 18847 10287 18853
rect 12802 18844 12808 18896
rect 12860 18884 12866 18896
rect 14001 18887 14059 18893
rect 14001 18884 14013 18887
rect 12860 18856 14013 18884
rect 12860 18844 12866 18856
rect 14001 18853 14013 18856
rect 14047 18853 14059 18887
rect 14001 18847 14059 18853
rect 14090 18844 14096 18896
rect 14148 18884 14154 18896
rect 14642 18884 14648 18896
rect 14148 18856 14648 18884
rect 14148 18844 14154 18856
rect 14642 18844 14648 18856
rect 14700 18884 14706 18896
rect 15289 18887 15347 18893
rect 15289 18884 15301 18887
rect 14700 18856 15301 18884
rect 14700 18844 14706 18856
rect 15289 18853 15301 18856
rect 15335 18853 15347 18887
rect 15289 18847 15347 18853
rect 18966 18844 18972 18896
rect 19024 18884 19030 18896
rect 20533 18887 20591 18893
rect 20533 18884 20545 18887
rect 19024 18856 20545 18884
rect 19024 18844 19030 18856
rect 20533 18853 20545 18856
rect 20579 18853 20591 18887
rect 21082 18884 21088 18896
rect 20533 18847 20591 18853
rect 20640 18856 21088 18884
rect 9784 18819 9847 18825
rect 9784 18788 9801 18819
rect 9789 18785 9801 18788
rect 9835 18785 9847 18819
rect 9789 18779 9847 18785
rect 12437 18819 12495 18825
rect 12437 18785 12449 18819
rect 12483 18816 12495 18819
rect 13265 18819 13323 18825
rect 13265 18816 13277 18819
rect 12483 18788 13277 18816
rect 12483 18785 12495 18788
rect 12437 18779 12495 18785
rect 13265 18785 13277 18788
rect 13311 18785 13323 18819
rect 13265 18779 13323 18785
rect 13354 18776 13360 18828
rect 13412 18816 13418 18828
rect 13814 18816 13820 18828
rect 13412 18788 13820 18816
rect 13412 18776 13418 18788
rect 13814 18776 13820 18788
rect 13872 18776 13878 18828
rect 14458 18816 14464 18828
rect 14419 18788 14464 18816
rect 14458 18776 14464 18788
rect 14516 18776 14522 18828
rect 15473 18819 15531 18825
rect 15473 18785 15485 18819
rect 15519 18785 15531 18819
rect 15473 18779 15531 18785
rect 9677 18751 9735 18757
rect 8772 18720 8892 18748
rect 5408 18652 8708 18680
rect 5408 18640 5414 18652
rect 2133 18615 2191 18621
rect 2133 18581 2145 18615
rect 2179 18612 2191 18615
rect 2222 18612 2228 18624
rect 2179 18584 2228 18612
rect 2179 18581 2191 18584
rect 2133 18575 2191 18581
rect 2222 18572 2228 18584
rect 2280 18572 2286 18624
rect 3878 18572 3884 18624
rect 3936 18612 3942 18624
rect 5718 18612 5724 18624
rect 3936 18584 5724 18612
rect 3936 18572 3942 18584
rect 5718 18572 5724 18584
rect 5776 18612 5782 18624
rect 6086 18612 6092 18624
rect 5776 18584 6092 18612
rect 5776 18572 5782 18584
rect 6086 18572 6092 18584
rect 6144 18572 6150 18624
rect 8864 18612 8892 18720
rect 9677 18717 9689 18751
rect 9723 18748 9735 18751
rect 10042 18748 10048 18760
rect 9723 18720 10048 18748
rect 9723 18717 9735 18720
rect 9677 18711 9735 18717
rect 10042 18708 10048 18720
rect 10100 18708 10106 18760
rect 10781 18751 10839 18757
rect 10781 18717 10793 18751
rect 10827 18717 10839 18751
rect 11054 18748 11060 18760
rect 11015 18720 11060 18748
rect 10781 18711 10839 18717
rect 9858 18640 9864 18692
rect 9916 18680 9922 18692
rect 10594 18680 10600 18692
rect 9916 18652 10600 18680
rect 9916 18640 9922 18652
rect 10594 18640 10600 18652
rect 10652 18680 10658 18692
rect 10796 18680 10824 18711
rect 11054 18708 11060 18720
rect 11112 18708 11118 18760
rect 12710 18708 12716 18760
rect 12768 18748 12774 18760
rect 12989 18751 13047 18757
rect 12989 18748 13001 18751
rect 12768 18720 13001 18748
rect 12768 18708 12774 18720
rect 12989 18717 13001 18720
rect 13035 18748 13047 18751
rect 13078 18748 13084 18760
rect 13035 18720 13084 18748
rect 13035 18717 13047 18720
rect 12989 18711 13047 18717
rect 13078 18708 13084 18720
rect 13136 18708 13142 18760
rect 13906 18708 13912 18760
rect 13964 18748 13970 18760
rect 15488 18748 15516 18779
rect 15930 18776 15936 18828
rect 15988 18816 15994 18828
rect 16761 18819 16819 18825
rect 16761 18816 16773 18819
rect 15988 18788 16773 18816
rect 15988 18776 15994 18788
rect 16761 18785 16773 18788
rect 16807 18785 16819 18819
rect 16761 18779 16819 18785
rect 18417 18819 18475 18825
rect 18417 18785 18429 18819
rect 18463 18816 18475 18819
rect 19058 18816 19064 18828
rect 18463 18788 19064 18816
rect 18463 18785 18475 18788
rect 18417 18779 18475 18785
rect 19058 18776 19064 18788
rect 19116 18776 19122 18828
rect 19334 18816 19340 18828
rect 19295 18788 19340 18816
rect 19334 18776 19340 18788
rect 19392 18776 19398 18828
rect 19518 18776 19524 18828
rect 19576 18816 19582 18828
rect 19613 18819 19671 18825
rect 19613 18816 19625 18819
rect 19576 18788 19625 18816
rect 19576 18776 19582 18788
rect 19613 18785 19625 18788
rect 19659 18785 19671 18819
rect 19613 18779 19671 18785
rect 19702 18776 19708 18828
rect 19760 18816 19766 18828
rect 20073 18819 20131 18825
rect 20073 18816 20085 18819
rect 19760 18788 20085 18816
rect 19760 18776 19766 18788
rect 20073 18785 20085 18788
rect 20119 18785 20131 18819
rect 20073 18779 20131 18785
rect 13964 18720 15516 18748
rect 17037 18751 17095 18757
rect 13964 18708 13970 18720
rect 17037 18717 17049 18751
rect 17083 18748 17095 18751
rect 17954 18748 17960 18760
rect 17083 18720 17960 18748
rect 17083 18717 17095 18720
rect 17037 18711 17095 18717
rect 17954 18708 17960 18720
rect 18012 18708 18018 18760
rect 18322 18708 18328 18760
rect 18380 18748 18386 18760
rect 18877 18751 18935 18757
rect 18877 18748 18889 18751
rect 18380 18720 18889 18748
rect 18380 18708 18386 18720
rect 18877 18717 18889 18720
rect 18923 18717 18935 18751
rect 18877 18711 18935 18717
rect 19242 18708 19248 18760
rect 19300 18748 19306 18760
rect 19300 18720 19932 18748
rect 19300 18708 19306 18720
rect 10652 18652 10824 18680
rect 10652 18640 10658 18652
rect 18046 18640 18052 18692
rect 18104 18680 18110 18692
rect 19613 18683 19671 18689
rect 19613 18680 19625 18683
rect 18104 18652 19625 18680
rect 18104 18640 18110 18652
rect 19613 18649 19625 18652
rect 19659 18649 19671 18683
rect 19904 18680 19932 18720
rect 19978 18708 19984 18760
rect 20036 18748 20042 18760
rect 20640 18748 20668 18856
rect 21082 18844 21088 18856
rect 21140 18844 21146 18896
rect 21358 18844 21364 18896
rect 21416 18884 21422 18896
rect 21453 18887 21511 18893
rect 21453 18884 21465 18887
rect 21416 18856 21465 18884
rect 21416 18844 21422 18856
rect 21453 18853 21465 18856
rect 21499 18853 21511 18887
rect 21453 18847 21511 18853
rect 21637 18887 21695 18893
rect 21637 18853 21649 18887
rect 21683 18884 21695 18887
rect 21818 18884 21824 18896
rect 21683 18856 21824 18884
rect 21683 18853 21695 18856
rect 21637 18847 21695 18853
rect 21818 18844 21824 18856
rect 21876 18844 21882 18896
rect 22002 18884 22008 18896
rect 21963 18856 22008 18884
rect 22002 18844 22008 18856
rect 22060 18844 22066 18896
rect 22097 18887 22155 18893
rect 22097 18853 22109 18887
rect 22143 18884 22155 18887
rect 23842 18884 23848 18896
rect 22143 18856 23848 18884
rect 22143 18853 22155 18856
rect 22097 18847 22155 18853
rect 23842 18844 23848 18856
rect 23900 18844 23906 18896
rect 24854 18884 24860 18896
rect 23952 18856 24860 18884
rect 20901 18819 20959 18825
rect 20901 18785 20913 18819
rect 20947 18785 20959 18819
rect 20901 18779 20959 18785
rect 21545 18819 21603 18825
rect 21545 18785 21557 18819
rect 21591 18816 21603 18819
rect 22462 18816 22468 18828
rect 21591 18788 22468 18816
rect 21591 18785 21603 18788
rect 21545 18779 21603 18785
rect 20036 18720 20668 18748
rect 20036 18708 20042 18720
rect 20916 18680 20944 18779
rect 22462 18776 22468 18788
rect 22520 18776 22526 18828
rect 22557 18819 22615 18825
rect 22557 18785 22569 18819
rect 22603 18785 22615 18819
rect 22557 18779 22615 18785
rect 22741 18819 22799 18825
rect 22741 18785 22753 18819
rect 22787 18816 22799 18819
rect 22830 18816 22836 18828
rect 22787 18788 22836 18816
rect 22787 18785 22799 18788
rect 22741 18779 22799 18785
rect 21269 18751 21327 18757
rect 21269 18717 21281 18751
rect 21315 18748 21327 18751
rect 22094 18748 22100 18760
rect 21315 18720 22100 18748
rect 21315 18717 21327 18720
rect 21269 18711 21327 18717
rect 22094 18708 22100 18720
rect 22152 18748 22158 18760
rect 22278 18748 22284 18760
rect 22152 18720 22284 18748
rect 22152 18708 22158 18720
rect 22278 18708 22284 18720
rect 22336 18708 22342 18760
rect 21174 18680 21180 18692
rect 19904 18652 21180 18680
rect 19613 18643 19671 18649
rect 21174 18640 21180 18652
rect 21232 18640 21238 18692
rect 22572 18680 22600 18779
rect 22830 18776 22836 18788
rect 22888 18776 22894 18828
rect 22925 18819 22983 18825
rect 22925 18785 22937 18819
rect 22971 18785 22983 18819
rect 22925 18779 22983 18785
rect 22940 18748 22968 18779
rect 23198 18776 23204 18828
rect 23256 18816 23262 18828
rect 23661 18819 23719 18825
rect 23661 18816 23673 18819
rect 23256 18788 23673 18816
rect 23256 18776 23262 18788
rect 23661 18785 23673 18788
rect 23707 18816 23719 18819
rect 23952 18816 23980 18856
rect 24854 18844 24860 18856
rect 24912 18844 24918 18896
rect 26712 18884 26740 18912
rect 34790 18884 34796 18896
rect 26712 18856 27844 18884
rect 23707 18788 23980 18816
rect 24029 18819 24087 18825
rect 23707 18785 23719 18788
rect 23661 18779 23719 18785
rect 24029 18785 24041 18819
rect 24075 18816 24087 18819
rect 24394 18816 24400 18828
rect 24075 18788 24400 18816
rect 24075 18785 24087 18788
rect 24029 18779 24087 18785
rect 24044 18748 24072 18779
rect 24394 18776 24400 18788
rect 24452 18776 24458 18828
rect 25222 18816 25228 18828
rect 25183 18788 25228 18816
rect 25222 18776 25228 18788
rect 25280 18776 25286 18828
rect 25593 18819 25651 18825
rect 25593 18785 25605 18819
rect 25639 18816 25651 18819
rect 26234 18816 26240 18828
rect 25639 18788 26240 18816
rect 25639 18785 25651 18788
rect 25593 18779 25651 18785
rect 26234 18776 26240 18788
rect 26292 18776 26298 18828
rect 27816 18825 27844 18856
rect 34348 18856 34796 18884
rect 26513 18819 26571 18825
rect 26513 18785 26525 18819
rect 26559 18785 26571 18819
rect 26513 18779 26571 18785
rect 27525 18819 27583 18825
rect 27525 18785 27537 18819
rect 27571 18785 27583 18819
rect 27525 18779 27583 18785
rect 27801 18819 27859 18825
rect 27801 18785 27813 18819
rect 27847 18785 27859 18819
rect 27801 18779 27859 18785
rect 22940 18720 24072 18748
rect 24121 18751 24179 18757
rect 24121 18717 24133 18751
rect 24167 18748 24179 18751
rect 24302 18748 24308 18760
rect 24167 18720 24308 18748
rect 24167 18717 24179 18720
rect 24121 18711 24179 18717
rect 24302 18708 24308 18720
rect 24360 18708 24366 18760
rect 24854 18748 24860 18760
rect 24815 18720 24860 18748
rect 24854 18708 24860 18720
rect 24912 18708 24918 18760
rect 26142 18708 26148 18760
rect 26200 18748 26206 18760
rect 26528 18748 26556 18779
rect 26200 18720 26556 18748
rect 27540 18748 27568 18779
rect 28074 18776 28080 18828
rect 28132 18816 28138 18828
rect 28445 18819 28503 18825
rect 28445 18816 28457 18819
rect 28132 18788 28457 18816
rect 28132 18776 28138 18788
rect 28445 18785 28457 18788
rect 28491 18816 28503 18819
rect 28534 18816 28540 18828
rect 28491 18788 28540 18816
rect 28491 18785 28503 18788
rect 28445 18779 28503 18785
rect 28534 18776 28540 18788
rect 28592 18776 28598 18828
rect 29730 18776 29736 18828
rect 29788 18816 29794 18828
rect 30009 18819 30067 18825
rect 30009 18816 30021 18819
rect 29788 18788 30021 18816
rect 29788 18776 29794 18788
rect 30009 18785 30021 18788
rect 30055 18785 30067 18819
rect 30190 18816 30196 18828
rect 30151 18788 30196 18816
rect 30009 18779 30067 18785
rect 30190 18776 30196 18788
rect 30248 18776 30254 18828
rect 30469 18819 30527 18825
rect 30469 18785 30481 18819
rect 30515 18785 30527 18819
rect 30650 18816 30656 18828
rect 30611 18788 30656 18816
rect 30469 18779 30527 18785
rect 29086 18748 29092 18760
rect 27540 18720 29092 18748
rect 26200 18708 26206 18720
rect 29086 18708 29092 18720
rect 29144 18708 29150 18760
rect 29546 18748 29552 18760
rect 29507 18720 29552 18748
rect 29546 18708 29552 18720
rect 29604 18708 29610 18760
rect 30484 18748 30512 18779
rect 30650 18776 30656 18788
rect 30708 18776 30714 18828
rect 30929 18819 30987 18825
rect 30929 18785 30941 18819
rect 30975 18816 30987 18819
rect 31846 18816 31852 18828
rect 30975 18788 31852 18816
rect 30975 18785 30987 18788
rect 30929 18779 30987 18785
rect 31846 18776 31852 18788
rect 31904 18776 31910 18828
rect 32030 18776 32036 18828
rect 32088 18816 32094 18828
rect 32125 18819 32183 18825
rect 32125 18816 32137 18819
rect 32088 18788 32137 18816
rect 32088 18776 32094 18788
rect 32125 18785 32137 18788
rect 32171 18785 32183 18819
rect 32490 18816 32496 18828
rect 32451 18788 32496 18816
rect 32125 18779 32183 18785
rect 32490 18776 32496 18788
rect 32548 18776 32554 18828
rect 32950 18816 32956 18828
rect 32911 18788 32956 18816
rect 32950 18776 32956 18788
rect 33008 18776 33014 18828
rect 33042 18776 33048 18828
rect 33100 18816 33106 18828
rect 34348 18825 34376 18856
rect 34790 18844 34796 18856
rect 34848 18844 34854 18896
rect 33781 18819 33839 18825
rect 33781 18816 33793 18819
rect 33100 18788 33793 18816
rect 33100 18776 33106 18788
rect 33781 18785 33793 18788
rect 33827 18785 33839 18819
rect 33781 18779 33839 18785
rect 34333 18819 34391 18825
rect 34333 18785 34345 18819
rect 34379 18785 34391 18819
rect 34514 18816 34520 18828
rect 34475 18788 34520 18816
rect 34333 18779 34391 18785
rect 34514 18776 34520 18788
rect 34572 18776 34578 18828
rect 34698 18776 34704 18828
rect 34756 18816 34762 18828
rect 35069 18819 35127 18825
rect 35069 18816 35081 18819
rect 34756 18788 35081 18816
rect 34756 18776 34762 18788
rect 35069 18785 35081 18788
rect 35115 18785 35127 18819
rect 35069 18779 35127 18785
rect 35805 18819 35863 18825
rect 35805 18785 35817 18819
rect 35851 18816 35863 18819
rect 35894 18816 35900 18828
rect 35851 18788 35900 18816
rect 35851 18785 35863 18788
rect 35805 18779 35863 18785
rect 35894 18776 35900 18788
rect 35952 18776 35958 18828
rect 36740 18825 36768 18924
rect 36906 18884 36912 18896
rect 36867 18856 36912 18884
rect 36906 18844 36912 18856
rect 36964 18844 36970 18896
rect 38378 18884 38384 18896
rect 37200 18856 38384 18884
rect 37200 18825 37228 18856
rect 38378 18844 38384 18856
rect 38436 18844 38442 18896
rect 38488 18828 38516 18924
rect 36357 18819 36415 18825
rect 36357 18785 36369 18819
rect 36403 18785 36415 18819
rect 36357 18779 36415 18785
rect 36725 18819 36783 18825
rect 36725 18785 36737 18819
rect 36771 18785 36783 18819
rect 36725 18779 36783 18785
rect 37185 18819 37243 18825
rect 37185 18785 37197 18819
rect 37231 18785 37243 18819
rect 37185 18779 37243 18785
rect 32968 18748 32996 18776
rect 34606 18748 34612 18760
rect 30484 18720 32996 18748
rect 34567 18720 34612 18748
rect 34606 18708 34612 18720
rect 34664 18708 34670 18760
rect 36372 18748 36400 18779
rect 38102 18776 38108 18828
rect 38160 18816 38166 18828
rect 38289 18819 38347 18825
rect 38289 18816 38301 18819
rect 38160 18788 38301 18816
rect 38160 18776 38166 18788
rect 38289 18785 38301 18788
rect 38335 18785 38347 18819
rect 38289 18779 38347 18785
rect 38470 18776 38476 18828
rect 38528 18816 38534 18828
rect 38657 18819 38715 18825
rect 38657 18816 38669 18819
rect 38528 18788 38669 18816
rect 38528 18776 38534 18788
rect 38657 18785 38669 18788
rect 38703 18785 38715 18819
rect 38657 18779 38715 18785
rect 38194 18748 38200 18760
rect 36372 18720 38200 18748
rect 38194 18708 38200 18720
rect 38252 18708 38258 18760
rect 38749 18751 38807 18757
rect 38749 18717 38761 18751
rect 38795 18717 38807 18751
rect 38749 18711 38807 18717
rect 23198 18680 23204 18692
rect 22572 18652 23204 18680
rect 23198 18640 23204 18652
rect 23256 18640 23262 18692
rect 23477 18683 23535 18689
rect 23477 18649 23489 18683
rect 23523 18680 23535 18683
rect 23842 18680 23848 18692
rect 23523 18652 23848 18680
rect 23523 18649 23535 18652
rect 23477 18643 23535 18649
rect 23842 18640 23848 18652
rect 23900 18640 23906 18692
rect 25498 18680 25504 18692
rect 25459 18652 25504 18680
rect 25498 18640 25504 18652
rect 25556 18640 25562 18692
rect 29362 18640 29368 18692
rect 29420 18680 29426 18692
rect 33042 18680 33048 18692
rect 29420 18652 33048 18680
rect 29420 18640 29426 18652
rect 33042 18640 33048 18652
rect 33100 18640 33106 18692
rect 38105 18683 38163 18689
rect 38105 18649 38117 18683
rect 38151 18680 38163 18683
rect 38654 18680 38660 18692
rect 38151 18652 38660 18680
rect 38151 18649 38163 18652
rect 38105 18643 38163 18649
rect 38654 18640 38660 18652
rect 38712 18640 38718 18692
rect 9766 18612 9772 18624
rect 8864 18584 9772 18612
rect 9766 18572 9772 18584
rect 9824 18572 9830 18624
rect 14645 18615 14703 18621
rect 14645 18581 14657 18615
rect 14691 18612 14703 18615
rect 17862 18612 17868 18624
rect 14691 18584 17868 18612
rect 14691 18581 14703 18584
rect 14645 18575 14703 18581
rect 17862 18572 17868 18584
rect 17920 18572 17926 18624
rect 18414 18572 18420 18624
rect 18472 18612 18478 18624
rect 19978 18612 19984 18624
rect 18472 18584 19984 18612
rect 18472 18572 18478 18584
rect 19978 18572 19984 18584
rect 20036 18572 20042 18624
rect 21085 18615 21143 18621
rect 21085 18581 21097 18615
rect 21131 18612 21143 18615
rect 21634 18612 21640 18624
rect 21131 18584 21640 18612
rect 21131 18581 21143 18584
rect 21085 18575 21143 18581
rect 21634 18572 21640 18584
rect 21692 18572 21698 18624
rect 27338 18612 27344 18624
rect 27299 18584 27344 18612
rect 27338 18572 27344 18584
rect 27396 18572 27402 18624
rect 27430 18572 27436 18624
rect 27488 18612 27494 18624
rect 28629 18615 28687 18621
rect 28629 18612 28641 18615
rect 27488 18584 28641 18612
rect 27488 18572 27494 18584
rect 28629 18581 28641 18584
rect 28675 18581 28687 18615
rect 28629 18575 28687 18581
rect 31938 18572 31944 18624
rect 31996 18612 32002 18624
rect 32217 18615 32275 18621
rect 32217 18612 32229 18615
rect 31996 18584 32229 18612
rect 31996 18572 32002 18584
rect 32217 18581 32229 18584
rect 32263 18581 32275 18615
rect 32217 18575 32275 18581
rect 35894 18572 35900 18624
rect 35952 18612 35958 18624
rect 38764 18612 38792 18711
rect 35952 18584 38792 18612
rect 35952 18572 35958 18584
rect 1104 18522 39836 18544
rect 1104 18470 4246 18522
rect 4298 18470 4310 18522
rect 4362 18470 4374 18522
rect 4426 18470 4438 18522
rect 4490 18470 34966 18522
rect 35018 18470 35030 18522
rect 35082 18470 35094 18522
rect 35146 18470 35158 18522
rect 35210 18470 39836 18522
rect 1104 18448 39836 18470
rect 9217 18411 9275 18417
rect 9217 18377 9229 18411
rect 9263 18408 9275 18411
rect 9766 18408 9772 18420
rect 9263 18380 9772 18408
rect 9263 18377 9275 18380
rect 9217 18371 9275 18377
rect 9766 18368 9772 18380
rect 9824 18368 9830 18420
rect 9950 18368 9956 18420
rect 10008 18408 10014 18420
rect 11425 18411 11483 18417
rect 11425 18408 11437 18411
rect 10008 18380 11437 18408
rect 10008 18368 10014 18380
rect 11425 18377 11437 18380
rect 11471 18408 11483 18411
rect 12342 18408 12348 18420
rect 11471 18380 12348 18408
rect 11471 18377 11483 18380
rect 11425 18371 11483 18377
rect 12342 18368 12348 18380
rect 12400 18368 12406 18420
rect 12437 18411 12495 18417
rect 12437 18377 12449 18411
rect 12483 18408 12495 18411
rect 12483 18380 17172 18408
rect 12483 18377 12495 18380
rect 12437 18371 12495 18377
rect 4614 18300 4620 18352
rect 4672 18340 4678 18352
rect 5537 18343 5595 18349
rect 5537 18340 5549 18343
rect 4672 18312 5549 18340
rect 4672 18300 4678 18312
rect 5537 18309 5549 18312
rect 5583 18309 5595 18343
rect 5537 18303 5595 18309
rect 6273 18343 6331 18349
rect 6273 18309 6285 18343
rect 6319 18340 6331 18343
rect 6822 18340 6828 18352
rect 6319 18312 6828 18340
rect 6319 18309 6331 18312
rect 6273 18303 6331 18309
rect 6822 18300 6828 18312
rect 6880 18340 6886 18352
rect 7834 18340 7840 18352
rect 6880 18312 7840 18340
rect 6880 18300 6886 18312
rect 7834 18300 7840 18312
rect 7892 18300 7898 18352
rect 10318 18300 10324 18352
rect 10376 18340 10382 18352
rect 13906 18340 13912 18352
rect 10376 18312 13912 18340
rect 10376 18300 10382 18312
rect 13906 18300 13912 18312
rect 13964 18300 13970 18352
rect 2866 18232 2872 18284
rect 2924 18272 2930 18284
rect 4893 18275 4951 18281
rect 4893 18272 4905 18275
rect 2924 18244 4905 18272
rect 2924 18232 2930 18244
rect 2774 18164 2780 18216
rect 2832 18204 2838 18216
rect 3510 18204 3516 18216
rect 2832 18176 2877 18204
rect 3471 18176 3516 18204
rect 2832 18164 2838 18176
rect 3510 18164 3516 18176
rect 3568 18164 3574 18216
rect 3804 18213 3832 18244
rect 4893 18241 4905 18244
rect 4939 18272 4951 18275
rect 5442 18272 5448 18284
rect 4939 18244 5448 18272
rect 4939 18241 4951 18244
rect 4893 18235 4951 18241
rect 5442 18232 5448 18244
rect 5500 18232 5506 18284
rect 10336 18272 10364 18300
rect 8220 18244 10364 18272
rect 11793 18275 11851 18281
rect 3789 18207 3847 18213
rect 3789 18173 3801 18207
rect 3835 18173 3847 18207
rect 3789 18167 3847 18173
rect 4157 18207 4215 18213
rect 4157 18173 4169 18207
rect 4203 18204 4215 18207
rect 5261 18207 5319 18213
rect 5261 18204 5273 18207
rect 4203 18176 5273 18204
rect 4203 18173 4215 18176
rect 4157 18167 4215 18173
rect 5261 18173 5273 18176
rect 5307 18173 5319 18207
rect 5626 18204 5632 18216
rect 5587 18176 5632 18204
rect 5261 18167 5319 18173
rect 4249 18139 4307 18145
rect 3528 18108 4200 18136
rect 3528 18080 3556 18108
rect 3510 18028 3516 18080
rect 3568 18028 3574 18080
rect 4172 18068 4200 18108
rect 4249 18105 4261 18139
rect 4295 18136 4307 18139
rect 4706 18136 4712 18148
rect 4295 18108 4712 18136
rect 4295 18105 4307 18108
rect 4249 18099 4307 18105
rect 4706 18096 4712 18108
rect 4764 18096 4770 18148
rect 5276 18136 5304 18167
rect 5626 18164 5632 18176
rect 5684 18164 5690 18216
rect 6457 18207 6515 18213
rect 6457 18204 6469 18207
rect 5920 18176 6469 18204
rect 5810 18136 5816 18148
rect 5276 18108 5816 18136
rect 5810 18096 5816 18108
rect 5868 18096 5874 18148
rect 5920 18068 5948 18176
rect 6457 18173 6469 18176
rect 6503 18173 6515 18207
rect 6457 18167 6515 18173
rect 7009 18207 7067 18213
rect 7009 18173 7021 18207
rect 7055 18173 7067 18207
rect 7190 18204 7196 18216
rect 7151 18176 7196 18204
rect 7009 18167 7067 18173
rect 6914 18096 6920 18148
rect 6972 18136 6978 18148
rect 7024 18136 7052 18167
rect 7190 18164 7196 18176
rect 7248 18164 7254 18216
rect 8220 18213 8248 18244
rect 11793 18241 11805 18275
rect 11839 18272 11851 18275
rect 14826 18272 14832 18284
rect 11839 18244 14832 18272
rect 11839 18241 11851 18244
rect 11793 18235 11851 18241
rect 14826 18232 14832 18244
rect 14884 18232 14890 18284
rect 15194 18272 15200 18284
rect 15155 18244 15200 18272
rect 15194 18232 15200 18244
rect 15252 18232 15258 18284
rect 7561 18207 7619 18213
rect 7561 18173 7573 18207
rect 7607 18173 7619 18207
rect 7561 18167 7619 18173
rect 8205 18207 8263 18213
rect 8205 18173 8217 18207
rect 8251 18173 8263 18207
rect 8386 18204 8392 18216
rect 8347 18176 8392 18204
rect 8205 18167 8263 18173
rect 7576 18136 7604 18167
rect 8386 18164 8392 18176
rect 8444 18164 8450 18216
rect 8573 18207 8631 18213
rect 8573 18173 8585 18207
rect 8619 18173 8631 18207
rect 8573 18167 8631 18173
rect 9217 18207 9275 18213
rect 9217 18173 9229 18207
rect 9263 18204 9275 18207
rect 9309 18207 9367 18213
rect 9309 18204 9321 18207
rect 9263 18176 9321 18204
rect 9263 18173 9275 18176
rect 9217 18167 9275 18173
rect 9309 18173 9321 18176
rect 9355 18173 9367 18207
rect 9309 18167 9367 18173
rect 9585 18207 9643 18213
rect 9585 18173 9597 18207
rect 9631 18204 9643 18207
rect 10226 18204 10232 18216
rect 9631 18176 10232 18204
rect 9631 18173 9643 18176
rect 9585 18167 9643 18173
rect 8110 18136 8116 18148
rect 6972 18108 7144 18136
rect 7576 18108 8116 18136
rect 6972 18096 6978 18108
rect 4172 18040 5948 18068
rect 7116 18068 7144 18108
rect 8110 18096 8116 18108
rect 8168 18096 8174 18148
rect 8294 18096 8300 18148
rect 8352 18136 8358 18148
rect 8588 18136 8616 18167
rect 10226 18164 10232 18176
rect 10284 18164 10290 18216
rect 11609 18207 11667 18213
rect 11609 18173 11621 18207
rect 11655 18173 11667 18207
rect 11609 18167 11667 18173
rect 11701 18207 11759 18213
rect 11701 18173 11713 18207
rect 11747 18204 11759 18207
rect 12345 18207 12403 18213
rect 12345 18204 12357 18207
rect 11747 18176 12357 18204
rect 11747 18173 11759 18176
rect 11701 18167 11759 18173
rect 12345 18173 12357 18176
rect 12391 18173 12403 18207
rect 12618 18204 12624 18216
rect 12579 18176 12624 18204
rect 12345 18167 12403 18173
rect 11624 18136 11652 18167
rect 12618 18164 12624 18176
rect 12676 18164 12682 18216
rect 13449 18207 13507 18213
rect 13449 18204 13461 18207
rect 12912 18176 13461 18204
rect 12250 18136 12256 18148
rect 8352 18108 8616 18136
rect 10244 18108 11560 18136
rect 11624 18108 12256 18136
rect 8352 18096 8358 18108
rect 10244 18068 10272 18108
rect 7116 18040 10272 18068
rect 10410 18028 10416 18080
rect 10468 18068 10474 18080
rect 10689 18071 10747 18077
rect 10689 18068 10701 18071
rect 10468 18040 10701 18068
rect 10468 18028 10474 18040
rect 10689 18037 10701 18040
rect 10735 18037 10747 18071
rect 11532 18068 11560 18108
rect 12250 18096 12256 18108
rect 12308 18096 12314 18148
rect 12912 18136 12940 18176
rect 13449 18173 13461 18176
rect 13495 18173 13507 18207
rect 14090 18204 14096 18216
rect 13449 18167 13507 18173
rect 13740 18176 14096 18204
rect 12360 18108 12940 18136
rect 13265 18139 13323 18145
rect 12360 18068 12388 18108
rect 13265 18105 13277 18139
rect 13311 18136 13323 18139
rect 13740 18136 13768 18176
rect 14090 18164 14096 18176
rect 14148 18164 14154 18216
rect 14277 18207 14335 18213
rect 14277 18173 14289 18207
rect 14323 18173 14335 18207
rect 14277 18167 14335 18173
rect 14921 18207 14979 18213
rect 14921 18173 14933 18207
rect 14967 18204 14979 18207
rect 15286 18204 15292 18216
rect 14967 18176 15292 18204
rect 14967 18173 14979 18176
rect 14921 18167 14979 18173
rect 13311 18108 13768 18136
rect 13817 18139 13875 18145
rect 13311 18105 13323 18108
rect 13265 18099 13323 18105
rect 13817 18105 13829 18139
rect 13863 18136 13875 18139
rect 14182 18136 14188 18148
rect 13863 18108 14188 18136
rect 13863 18105 13875 18108
rect 13817 18099 13875 18105
rect 14182 18096 14188 18108
rect 14240 18096 14246 18148
rect 14292 18136 14320 18167
rect 15286 18164 15292 18176
rect 15344 18204 15350 18216
rect 15930 18204 15936 18216
rect 15344 18176 15936 18204
rect 15344 18164 15350 18176
rect 15930 18164 15936 18176
rect 15988 18164 15994 18216
rect 17144 18136 17172 18380
rect 17862 18368 17868 18420
rect 17920 18408 17926 18420
rect 19518 18408 19524 18420
rect 17920 18380 19524 18408
rect 17920 18368 17926 18380
rect 19518 18368 19524 18380
rect 19576 18368 19582 18420
rect 19613 18411 19671 18417
rect 19613 18377 19625 18411
rect 19659 18408 19671 18411
rect 19702 18408 19708 18420
rect 19659 18380 19708 18408
rect 19659 18377 19671 18380
rect 19613 18371 19671 18377
rect 19702 18368 19708 18380
rect 19760 18368 19766 18420
rect 19981 18411 20039 18417
rect 19981 18377 19993 18411
rect 20027 18408 20039 18411
rect 22278 18408 22284 18420
rect 20027 18380 22284 18408
rect 20027 18377 20039 18380
rect 19981 18371 20039 18377
rect 22278 18368 22284 18380
rect 22336 18408 22342 18420
rect 22830 18408 22836 18420
rect 22336 18380 22836 18408
rect 22336 18368 22342 18380
rect 22830 18368 22836 18380
rect 22888 18368 22894 18420
rect 29270 18368 29276 18420
rect 29328 18408 29334 18420
rect 35710 18408 35716 18420
rect 29328 18380 35716 18408
rect 29328 18368 29334 18380
rect 35710 18368 35716 18380
rect 35768 18368 35774 18420
rect 36630 18368 36636 18420
rect 36688 18408 36694 18420
rect 39022 18408 39028 18420
rect 36688 18380 39028 18408
rect 36688 18368 36694 18380
rect 39022 18368 39028 18380
rect 39080 18368 39086 18420
rect 21174 18300 21180 18352
rect 21232 18340 21238 18352
rect 21545 18343 21603 18349
rect 21545 18340 21557 18343
rect 21232 18312 21557 18340
rect 21232 18300 21238 18312
rect 21545 18309 21557 18312
rect 21591 18309 21603 18343
rect 21545 18303 21603 18309
rect 22186 18300 22192 18352
rect 22244 18340 22250 18352
rect 22373 18343 22431 18349
rect 22373 18340 22385 18343
rect 22244 18312 22385 18340
rect 22244 18300 22250 18312
rect 22373 18309 22385 18312
rect 22419 18309 22431 18343
rect 23934 18340 23940 18352
rect 23895 18312 23940 18340
rect 22373 18303 22431 18309
rect 23934 18300 23940 18312
rect 23992 18300 23998 18352
rect 29454 18340 29460 18352
rect 29415 18312 29460 18340
rect 29454 18300 29460 18312
rect 29512 18300 29518 18352
rect 32950 18340 32956 18352
rect 32911 18312 32956 18340
rect 32950 18300 32956 18312
rect 33008 18300 33014 18352
rect 34330 18300 34336 18352
rect 34388 18340 34394 18352
rect 35069 18343 35127 18349
rect 35069 18340 35081 18343
rect 34388 18312 35081 18340
rect 34388 18300 34394 18312
rect 35069 18309 35081 18312
rect 35115 18309 35127 18343
rect 35069 18303 35127 18309
rect 18049 18275 18107 18281
rect 18049 18241 18061 18275
rect 18095 18272 18107 18275
rect 18690 18272 18696 18284
rect 18095 18244 18696 18272
rect 18095 18241 18107 18244
rect 18049 18235 18107 18241
rect 18690 18232 18696 18244
rect 18748 18232 18754 18284
rect 23842 18272 23848 18284
rect 19812 18244 21128 18272
rect 23803 18244 23848 18272
rect 17221 18207 17279 18213
rect 17221 18173 17233 18207
rect 17267 18204 17279 18207
rect 18138 18204 18144 18216
rect 17267 18176 18144 18204
rect 17267 18173 17279 18176
rect 17221 18167 17279 18173
rect 18138 18164 18144 18176
rect 18196 18164 18202 18216
rect 18322 18204 18328 18216
rect 18283 18176 18328 18204
rect 18322 18164 18328 18176
rect 18380 18164 18386 18216
rect 18708 18204 18736 18232
rect 19812 18213 19840 18244
rect 19797 18207 19855 18213
rect 18708 18176 19748 18204
rect 19720 18136 19748 18176
rect 19797 18173 19809 18207
rect 19843 18173 19855 18207
rect 19797 18167 19855 18173
rect 20165 18207 20223 18213
rect 20165 18173 20177 18207
rect 20211 18173 20223 18207
rect 20438 18204 20444 18216
rect 20399 18176 20444 18204
rect 20165 18167 20223 18173
rect 20180 18136 20208 18167
rect 20438 18164 20444 18176
rect 20496 18164 20502 18216
rect 14292 18108 15056 18136
rect 17144 18108 18184 18136
rect 19720 18108 20208 18136
rect 11532 18040 12388 18068
rect 10689 18031 10747 18037
rect 12434 18028 12440 18080
rect 12492 18068 12498 18080
rect 12713 18071 12771 18077
rect 12713 18068 12725 18071
rect 12492 18040 12725 18068
rect 12492 18028 12498 18040
rect 12713 18037 12725 18040
rect 12759 18037 12771 18071
rect 12713 18031 12771 18037
rect 14369 18071 14427 18077
rect 14369 18037 14381 18071
rect 14415 18068 14427 18071
rect 14918 18068 14924 18080
rect 14415 18040 14924 18068
rect 14415 18037 14427 18040
rect 14369 18031 14427 18037
rect 14918 18028 14924 18040
rect 14976 18028 14982 18080
rect 15028 18068 15056 18108
rect 16114 18068 16120 18080
rect 15028 18040 16120 18068
rect 16114 18028 16120 18040
rect 16172 18028 16178 18080
rect 16298 18068 16304 18080
rect 16259 18040 16304 18068
rect 16298 18028 16304 18040
rect 16356 18028 16362 18080
rect 17402 18068 17408 18080
rect 17363 18040 17408 18068
rect 17402 18028 17408 18040
rect 17460 18028 17466 18080
rect 18156 18068 18184 18108
rect 19334 18068 19340 18080
rect 18156 18040 19340 18068
rect 19334 18028 19340 18040
rect 19392 18028 19398 18080
rect 21100 18068 21128 18244
rect 23842 18232 23848 18244
rect 23900 18232 23906 18284
rect 27154 18272 27160 18284
rect 27115 18244 27160 18272
rect 27154 18232 27160 18244
rect 27212 18232 27218 18284
rect 30190 18272 30196 18284
rect 27816 18244 30196 18272
rect 22554 18204 22560 18216
rect 22515 18176 22560 18204
rect 22554 18164 22560 18176
rect 22612 18164 22618 18216
rect 22738 18164 22744 18216
rect 22796 18204 22802 18216
rect 22833 18207 22891 18213
rect 22833 18204 22845 18207
rect 22796 18176 22845 18204
rect 22796 18164 22802 18176
rect 22833 18173 22845 18176
rect 22879 18173 22891 18207
rect 22833 18167 22891 18173
rect 24581 18207 24639 18213
rect 24581 18173 24593 18207
rect 24627 18204 24639 18207
rect 24670 18204 24676 18216
rect 24627 18176 24676 18204
rect 24627 18173 24639 18176
rect 24581 18167 24639 18173
rect 24670 18164 24676 18176
rect 24728 18164 24734 18216
rect 25041 18207 25099 18213
rect 25041 18173 25053 18207
rect 25087 18204 25099 18207
rect 25130 18204 25136 18216
rect 25087 18176 25136 18204
rect 25087 18173 25099 18176
rect 25041 18167 25099 18173
rect 25130 18164 25136 18176
rect 25188 18164 25194 18216
rect 25314 18204 25320 18216
rect 25275 18176 25320 18204
rect 25314 18164 25320 18176
rect 25372 18164 25378 18216
rect 25498 18204 25504 18216
rect 25459 18176 25504 18204
rect 25498 18164 25504 18176
rect 25556 18164 25562 18216
rect 26510 18204 26516 18216
rect 26471 18176 26516 18204
rect 26510 18164 26516 18176
rect 26568 18164 26574 18216
rect 26697 18207 26755 18213
rect 26697 18173 26709 18207
rect 26743 18204 26755 18207
rect 27338 18204 27344 18216
rect 26743 18176 27344 18204
rect 26743 18173 26755 18176
rect 26697 18167 26755 18173
rect 27338 18164 27344 18176
rect 27396 18164 27402 18216
rect 27816 18213 27844 18244
rect 30190 18232 30196 18244
rect 30248 18232 30254 18284
rect 33594 18272 33600 18284
rect 31312 18244 33272 18272
rect 33507 18244 33600 18272
rect 27801 18207 27859 18213
rect 27801 18173 27813 18207
rect 27847 18173 27859 18207
rect 27801 18167 27859 18173
rect 28353 18207 28411 18213
rect 28353 18173 28365 18207
rect 28399 18173 28411 18207
rect 28626 18204 28632 18216
rect 28587 18176 28632 18204
rect 28353 18167 28411 18173
rect 22002 18096 22008 18148
rect 22060 18136 22066 18148
rect 23198 18136 23204 18148
rect 22060 18108 23204 18136
rect 22060 18096 22066 18108
rect 23198 18096 23204 18108
rect 23256 18096 23262 18148
rect 26605 18139 26663 18145
rect 26605 18105 26617 18139
rect 26651 18136 26663 18139
rect 28368 18136 28396 18167
rect 28626 18164 28632 18176
rect 28684 18164 28690 18216
rect 29270 18204 29276 18216
rect 29231 18176 29276 18204
rect 29270 18164 29276 18176
rect 29328 18164 29334 18216
rect 29546 18164 29552 18216
rect 29604 18204 29610 18216
rect 29825 18207 29883 18213
rect 29825 18204 29837 18207
rect 29604 18176 29837 18204
rect 29604 18164 29610 18176
rect 29825 18173 29837 18176
rect 29871 18173 29883 18207
rect 29825 18167 29883 18173
rect 30285 18207 30343 18213
rect 30285 18173 30297 18207
rect 30331 18204 30343 18207
rect 30834 18204 30840 18216
rect 30331 18176 30840 18204
rect 30331 18173 30343 18176
rect 30285 18167 30343 18173
rect 30834 18164 30840 18176
rect 30892 18164 30898 18216
rect 31312 18213 31340 18244
rect 31297 18207 31355 18213
rect 31297 18173 31309 18207
rect 31343 18173 31355 18207
rect 31297 18167 31355 18173
rect 32033 18207 32091 18213
rect 32033 18173 32045 18207
rect 32079 18173 32091 18207
rect 33134 18204 33140 18216
rect 33095 18176 33140 18204
rect 32033 18167 32091 18173
rect 29086 18136 29092 18148
rect 26651 18108 28304 18136
rect 28368 18108 29092 18136
rect 26651 18105 26663 18108
rect 26605 18099 26663 18105
rect 22094 18068 22100 18080
rect 21100 18040 22100 18068
rect 22094 18028 22100 18040
rect 22152 18028 22158 18080
rect 27709 18071 27767 18077
rect 27709 18037 27721 18071
rect 27755 18068 27767 18071
rect 27982 18068 27988 18080
rect 27755 18040 27988 18068
rect 27755 18037 27767 18040
rect 27709 18031 27767 18037
rect 27982 18028 27988 18040
rect 28040 18028 28046 18080
rect 28276 18068 28304 18108
rect 29086 18096 29092 18108
rect 29144 18096 29150 18148
rect 28718 18068 28724 18080
rect 28276 18040 28724 18068
rect 28718 18028 28724 18040
rect 28776 18028 28782 18080
rect 30282 18028 30288 18080
rect 30340 18068 30346 18080
rect 31481 18071 31539 18077
rect 31481 18068 31493 18071
rect 30340 18040 31493 18068
rect 30340 18028 30346 18040
rect 31481 18037 31493 18040
rect 31527 18037 31539 18071
rect 32048 18068 32076 18167
rect 33134 18164 33140 18176
rect 33192 18164 33198 18216
rect 33244 18204 33272 18244
rect 33594 18232 33600 18244
rect 33652 18272 33658 18284
rect 34241 18275 34299 18281
rect 34241 18272 34253 18275
rect 33652 18244 34253 18272
rect 33652 18232 33658 18244
rect 34241 18241 34253 18244
rect 34287 18241 34299 18275
rect 34241 18235 34299 18241
rect 34422 18232 34428 18284
rect 34480 18272 34486 18284
rect 35713 18275 35771 18281
rect 35713 18272 35725 18275
rect 34480 18244 35725 18272
rect 34480 18232 34486 18244
rect 35713 18241 35725 18244
rect 35759 18272 35771 18275
rect 36078 18272 36084 18284
rect 35759 18244 36084 18272
rect 35759 18241 35771 18244
rect 35713 18235 35771 18241
rect 36078 18232 36084 18244
rect 36136 18232 36142 18284
rect 38562 18272 38568 18284
rect 38523 18244 38568 18272
rect 38562 18232 38568 18244
rect 38620 18232 38626 18284
rect 33502 18204 33508 18216
rect 33244 18176 33508 18204
rect 33502 18164 33508 18176
rect 33560 18164 33566 18216
rect 33686 18164 33692 18216
rect 33744 18204 33750 18216
rect 34149 18207 34207 18213
rect 34149 18204 34161 18207
rect 33744 18176 34161 18204
rect 33744 18164 33750 18176
rect 34149 18173 34161 18176
rect 34195 18173 34207 18207
rect 34149 18167 34207 18173
rect 34790 18164 34796 18216
rect 34848 18204 34854 18216
rect 34885 18207 34943 18213
rect 34885 18204 34897 18207
rect 34848 18176 34897 18204
rect 34848 18164 34854 18176
rect 34885 18173 34897 18176
rect 34931 18173 34943 18207
rect 35986 18204 35992 18216
rect 35947 18176 35992 18204
rect 34885 18167 34943 18173
rect 35986 18164 35992 18176
rect 36044 18164 36050 18216
rect 38194 18204 38200 18216
rect 38155 18176 38200 18204
rect 38194 18164 38200 18176
rect 38252 18164 38258 18216
rect 38378 18204 38384 18216
rect 38339 18176 38384 18204
rect 38378 18164 38384 18176
rect 38436 18164 38442 18216
rect 38654 18204 38660 18216
rect 38615 18176 38660 18204
rect 38654 18164 38660 18176
rect 38712 18164 38718 18216
rect 32125 18139 32183 18145
rect 32125 18105 32137 18139
rect 32171 18136 32183 18139
rect 34514 18136 34520 18148
rect 32171 18108 34520 18136
rect 32171 18105 32183 18108
rect 32125 18099 32183 18105
rect 34514 18096 34520 18108
rect 34572 18096 34578 18148
rect 37369 18139 37427 18145
rect 34624 18108 35388 18136
rect 32858 18068 32864 18080
rect 32048 18040 32864 18068
rect 31481 18031 31539 18037
rect 32858 18028 32864 18040
rect 32916 18068 32922 18080
rect 34624 18068 34652 18108
rect 32916 18040 34652 18068
rect 35360 18068 35388 18108
rect 37369 18105 37381 18139
rect 37415 18136 37427 18139
rect 38562 18136 38568 18148
rect 37415 18108 38568 18136
rect 37415 18105 37427 18108
rect 37369 18099 37427 18105
rect 37384 18068 37412 18099
rect 38562 18096 38568 18108
rect 38620 18096 38626 18148
rect 35360 18040 37412 18068
rect 32916 18028 32922 18040
rect 1104 17978 39836 18000
rect 1104 17926 19606 17978
rect 19658 17926 19670 17978
rect 19722 17926 19734 17978
rect 19786 17926 19798 17978
rect 19850 17926 39836 17978
rect 1104 17904 39836 17926
rect 5442 17824 5448 17876
rect 5500 17864 5506 17876
rect 9769 17867 9827 17873
rect 5500 17836 7880 17864
rect 5500 17824 5506 17836
rect 3145 17799 3203 17805
rect 3145 17765 3157 17799
rect 3191 17796 3203 17799
rect 3878 17796 3884 17808
rect 3191 17768 3884 17796
rect 3191 17765 3203 17768
rect 3145 17759 3203 17765
rect 3878 17756 3884 17768
rect 3936 17756 3942 17808
rect 7852 17796 7880 17836
rect 9769 17833 9781 17867
rect 9815 17864 9827 17867
rect 10318 17864 10324 17876
rect 9815 17836 10324 17864
rect 9815 17833 9827 17836
rect 9769 17827 9827 17833
rect 10318 17824 10324 17836
rect 10376 17824 10382 17876
rect 13078 17824 13084 17876
rect 13136 17864 13142 17876
rect 24026 17864 24032 17876
rect 13136 17836 24032 17864
rect 13136 17824 13142 17836
rect 24026 17824 24032 17836
rect 24084 17824 24090 17876
rect 25774 17824 25780 17876
rect 25832 17864 25838 17876
rect 30929 17867 30987 17873
rect 30929 17864 30941 17867
rect 25832 17836 30941 17864
rect 25832 17824 25838 17836
rect 30929 17833 30941 17836
rect 30975 17833 30987 17867
rect 32398 17864 32404 17876
rect 32359 17836 32404 17864
rect 30929 17827 30987 17833
rect 32398 17824 32404 17836
rect 32456 17824 32462 17876
rect 33689 17867 33747 17873
rect 33689 17833 33701 17867
rect 33735 17864 33747 17867
rect 35342 17864 35348 17876
rect 33735 17836 35348 17864
rect 33735 17833 33747 17836
rect 33689 17827 33747 17833
rect 35342 17824 35348 17836
rect 35400 17824 35406 17876
rect 9214 17796 9220 17808
rect 4908 17768 6960 17796
rect 4908 17740 4936 17768
rect 1394 17688 1400 17740
rect 1452 17728 1458 17740
rect 1489 17731 1547 17737
rect 1489 17728 1501 17731
rect 1452 17700 1501 17728
rect 1452 17688 1458 17700
rect 1489 17697 1501 17700
rect 1535 17697 1547 17731
rect 1489 17691 1547 17697
rect 3970 17688 3976 17740
rect 4028 17728 4034 17740
rect 4065 17731 4123 17737
rect 4065 17728 4077 17731
rect 4028 17700 4077 17728
rect 4028 17688 4034 17700
rect 4065 17697 4077 17700
rect 4111 17697 4123 17731
rect 4890 17728 4896 17740
rect 4803 17700 4896 17728
rect 4065 17691 4123 17697
rect 4890 17688 4896 17700
rect 4948 17688 4954 17740
rect 5350 17728 5356 17740
rect 5311 17700 5356 17728
rect 5350 17688 5356 17700
rect 5408 17688 5414 17740
rect 5721 17731 5779 17737
rect 5721 17697 5733 17731
rect 5767 17728 5779 17731
rect 5902 17728 5908 17740
rect 5767 17700 5908 17728
rect 5767 17697 5779 17700
rect 5721 17691 5779 17697
rect 5902 17688 5908 17700
rect 5960 17688 5966 17740
rect 6086 17728 6092 17740
rect 6047 17700 6092 17728
rect 6086 17688 6092 17700
rect 6144 17688 6150 17740
rect 6932 17737 6960 17768
rect 7852 17768 9220 17796
rect 6917 17731 6975 17737
rect 6917 17697 6929 17731
rect 6963 17697 6975 17731
rect 7098 17728 7104 17740
rect 7059 17700 7104 17728
rect 6917 17691 6975 17697
rect 1762 17660 1768 17672
rect 1723 17632 1768 17660
rect 1762 17620 1768 17632
rect 1820 17620 1826 17672
rect 6932 17660 6960 17691
rect 7098 17688 7104 17700
rect 7156 17688 7162 17740
rect 7650 17728 7656 17740
rect 7611 17700 7656 17728
rect 7650 17688 7656 17700
rect 7708 17688 7714 17740
rect 7852 17728 7880 17768
rect 9214 17756 9220 17768
rect 9272 17796 9278 17808
rect 10873 17799 10931 17805
rect 9272 17768 9720 17796
rect 9272 17756 9278 17768
rect 7929 17731 7987 17737
rect 7929 17728 7941 17731
rect 7852 17700 7941 17728
rect 7929 17697 7941 17700
rect 7975 17697 7987 17731
rect 8570 17728 8576 17740
rect 8531 17700 8576 17728
rect 7929 17691 7987 17697
rect 8570 17688 8576 17700
rect 8628 17688 8634 17740
rect 9692 17737 9720 17768
rect 10873 17765 10885 17799
rect 10919 17796 10931 17799
rect 11054 17796 11060 17808
rect 10919 17768 11060 17796
rect 10919 17765 10931 17768
rect 10873 17759 10931 17765
rect 11054 17756 11060 17768
rect 11112 17756 11118 17808
rect 17954 17756 17960 17808
rect 18012 17796 18018 17808
rect 20165 17799 20223 17805
rect 20165 17796 20177 17799
rect 18012 17768 20177 17796
rect 18012 17756 18018 17768
rect 20165 17765 20177 17768
rect 20211 17765 20223 17799
rect 22738 17796 22744 17808
rect 20165 17759 20223 17765
rect 21652 17768 22416 17796
rect 9677 17731 9735 17737
rect 9677 17697 9689 17731
rect 9723 17697 9735 17731
rect 10410 17728 10416 17740
rect 10371 17700 10416 17728
rect 9677 17691 9735 17697
rect 10410 17688 10416 17700
rect 10468 17688 10474 17740
rect 13906 17728 13912 17740
rect 13867 17700 13912 17728
rect 13906 17688 13912 17700
rect 13964 17688 13970 17740
rect 14182 17688 14188 17740
rect 14240 17728 14246 17740
rect 14277 17731 14335 17737
rect 14277 17728 14289 17731
rect 14240 17700 14289 17728
rect 14240 17688 14246 17700
rect 14277 17697 14289 17700
rect 14323 17697 14335 17731
rect 15286 17728 15292 17740
rect 15247 17700 15292 17728
rect 14277 17691 14335 17697
rect 15286 17688 15292 17700
rect 15344 17688 15350 17740
rect 17586 17728 17592 17740
rect 17547 17700 17592 17728
rect 17586 17688 17592 17700
rect 17644 17688 17650 17740
rect 17681 17731 17739 17737
rect 17681 17697 17693 17731
rect 17727 17728 17739 17731
rect 17770 17728 17776 17740
rect 17727 17700 17776 17728
rect 17727 17697 17739 17700
rect 17681 17691 17739 17697
rect 17770 17688 17776 17700
rect 17828 17688 17834 17740
rect 18693 17731 18751 17737
rect 18693 17697 18705 17731
rect 18739 17728 18751 17731
rect 18874 17728 18880 17740
rect 18739 17700 18880 17728
rect 18739 17697 18751 17700
rect 18693 17691 18751 17697
rect 18874 17688 18880 17700
rect 18932 17688 18938 17740
rect 19705 17731 19763 17737
rect 19705 17697 19717 17731
rect 19751 17728 19763 17731
rect 20070 17728 20076 17740
rect 19751 17700 20076 17728
rect 19751 17697 19763 17700
rect 19705 17691 19763 17697
rect 20070 17688 20076 17700
rect 20128 17688 20134 17740
rect 8665 17663 8723 17669
rect 8665 17660 8677 17663
rect 6932 17632 8677 17660
rect 8665 17629 8677 17632
rect 8711 17629 8723 17663
rect 8665 17623 8723 17629
rect 10321 17663 10379 17669
rect 10321 17629 10333 17663
rect 10367 17660 10379 17663
rect 11238 17660 11244 17672
rect 10367 17632 11244 17660
rect 10367 17629 10379 17632
rect 10321 17623 10379 17629
rect 11238 17620 11244 17632
rect 11296 17620 11302 17672
rect 11333 17663 11391 17669
rect 11333 17629 11345 17663
rect 11379 17629 11391 17663
rect 11606 17660 11612 17672
rect 11567 17632 11612 17660
rect 11333 17623 11391 17629
rect 6089 17595 6147 17601
rect 6089 17561 6101 17595
rect 6135 17592 6147 17595
rect 8294 17592 8300 17604
rect 6135 17564 8300 17592
rect 6135 17561 6147 17564
rect 6089 17555 6147 17561
rect 8294 17552 8300 17564
rect 8352 17552 8358 17604
rect 9766 17552 9772 17604
rect 9824 17592 9830 17604
rect 11348 17592 11376 17623
rect 11606 17620 11612 17632
rect 11664 17620 11670 17672
rect 13630 17660 13636 17672
rect 13591 17632 13636 17660
rect 13630 17620 13636 17632
rect 13688 17620 13694 17672
rect 15562 17660 15568 17672
rect 15523 17632 15568 17660
rect 15562 17620 15568 17632
rect 15620 17620 15626 17672
rect 18598 17660 18604 17672
rect 18559 17632 18604 17660
rect 18598 17620 18604 17632
rect 18656 17620 18662 17672
rect 19613 17663 19671 17669
rect 19613 17660 19625 17663
rect 18708 17632 19625 17660
rect 9824 17564 11376 17592
rect 9824 17552 9830 17564
rect 13998 17552 14004 17604
rect 14056 17592 14062 17604
rect 14277 17595 14335 17601
rect 14277 17592 14289 17595
rect 14056 17564 14289 17592
rect 14056 17552 14062 17564
rect 14277 17561 14289 17564
rect 14323 17561 14335 17595
rect 14277 17555 14335 17561
rect 17402 17552 17408 17604
rect 17460 17592 17466 17604
rect 18708 17592 18736 17632
rect 19613 17629 19625 17632
rect 19659 17629 19671 17663
rect 19613 17623 19671 17629
rect 21082 17620 21088 17672
rect 21140 17660 21146 17672
rect 21361 17663 21419 17669
rect 21361 17660 21373 17663
rect 21140 17632 21373 17660
rect 21140 17620 21146 17632
rect 21361 17629 21373 17632
rect 21407 17629 21419 17663
rect 21361 17623 21419 17629
rect 17460 17564 18736 17592
rect 17460 17552 17466 17564
rect 19150 17552 19156 17604
rect 19208 17592 19214 17604
rect 21652 17592 21680 17768
rect 21726 17688 21732 17740
rect 21784 17728 21790 17740
rect 21821 17731 21879 17737
rect 21821 17728 21833 17731
rect 21784 17700 21833 17728
rect 21784 17688 21790 17700
rect 21821 17697 21833 17700
rect 21867 17697 21879 17731
rect 21821 17691 21879 17697
rect 22097 17731 22155 17737
rect 22097 17697 22109 17731
rect 22143 17728 22155 17731
rect 22281 17731 22339 17737
rect 22143 17700 22232 17728
rect 22143 17697 22155 17700
rect 22097 17691 22155 17697
rect 19208 17564 21680 17592
rect 19208 17552 19214 17564
rect 3970 17484 3976 17536
rect 4028 17524 4034 17536
rect 4157 17527 4215 17533
rect 4157 17524 4169 17527
rect 4028 17496 4169 17524
rect 4028 17484 4034 17496
rect 4157 17493 4169 17496
rect 4203 17493 4215 17527
rect 4157 17487 4215 17493
rect 8021 17527 8079 17533
rect 8021 17493 8033 17527
rect 8067 17524 8079 17527
rect 8110 17524 8116 17536
rect 8067 17496 8116 17524
rect 8067 17493 8079 17496
rect 8021 17487 8079 17493
rect 8110 17484 8116 17496
rect 8168 17484 8174 17536
rect 12894 17524 12900 17536
rect 12855 17496 12900 17524
rect 12894 17484 12900 17496
rect 12952 17484 12958 17536
rect 16666 17524 16672 17536
rect 16627 17496 16672 17524
rect 16666 17484 16672 17496
rect 16724 17484 16730 17536
rect 17862 17524 17868 17536
rect 17823 17496 17868 17524
rect 17862 17484 17868 17496
rect 17920 17484 17926 17536
rect 18322 17484 18328 17536
rect 18380 17524 18386 17536
rect 18877 17527 18935 17533
rect 18877 17524 18889 17527
rect 18380 17496 18889 17524
rect 18380 17484 18386 17496
rect 18877 17493 18889 17496
rect 18923 17493 18935 17527
rect 18877 17487 18935 17493
rect 22094 17484 22100 17536
rect 22152 17524 22158 17536
rect 22204 17524 22232 17700
rect 22281 17697 22293 17731
rect 22327 17697 22339 17731
rect 22281 17691 22339 17697
rect 22296 17592 22324 17691
rect 22388 17660 22416 17768
rect 22480 17768 22744 17796
rect 22480 17737 22508 17768
rect 22738 17756 22744 17768
rect 22796 17756 22802 17808
rect 24210 17756 24216 17808
rect 24268 17796 24274 17808
rect 30009 17799 30067 17805
rect 24268 17768 27476 17796
rect 24268 17756 24274 17768
rect 22465 17731 22523 17737
rect 22465 17697 22477 17731
rect 22511 17697 22523 17731
rect 22465 17691 22523 17697
rect 22649 17731 22707 17737
rect 22649 17697 22661 17731
rect 22695 17728 22707 17731
rect 22922 17728 22928 17740
rect 22695 17700 22928 17728
rect 22695 17697 22707 17700
rect 22649 17691 22707 17697
rect 22922 17688 22928 17700
rect 22980 17688 22986 17740
rect 23842 17728 23848 17740
rect 23803 17700 23848 17728
rect 23842 17688 23848 17700
rect 23900 17688 23906 17740
rect 24581 17731 24639 17737
rect 24581 17697 24593 17731
rect 24627 17728 24639 17731
rect 24670 17728 24676 17740
rect 24627 17700 24676 17728
rect 24627 17697 24639 17700
rect 24581 17691 24639 17697
rect 24670 17688 24676 17700
rect 24728 17688 24734 17740
rect 25041 17731 25099 17737
rect 25041 17697 25053 17731
rect 25087 17728 25099 17731
rect 25130 17728 25136 17740
rect 25087 17700 25136 17728
rect 25087 17697 25099 17700
rect 25041 17691 25099 17697
rect 25130 17688 25136 17700
rect 25188 17688 25194 17740
rect 25314 17728 25320 17740
rect 25227 17700 25320 17728
rect 25314 17688 25320 17700
rect 25372 17688 25378 17740
rect 25498 17728 25504 17740
rect 25459 17700 25504 17728
rect 25498 17688 25504 17700
rect 25556 17688 25562 17740
rect 26786 17728 26792 17740
rect 26747 17700 26792 17728
rect 26786 17688 26792 17700
rect 26844 17688 26850 17740
rect 26970 17688 26976 17740
rect 27028 17728 27034 17740
rect 27065 17731 27123 17737
rect 27065 17728 27077 17731
rect 27028 17700 27077 17728
rect 27028 17688 27034 17700
rect 27065 17697 27077 17700
rect 27111 17697 27123 17731
rect 27065 17691 27123 17697
rect 25332 17660 25360 17688
rect 26418 17660 26424 17672
rect 22388 17632 23980 17660
rect 25332 17632 26424 17660
rect 23750 17592 23756 17604
rect 22296 17564 23756 17592
rect 23750 17552 23756 17564
rect 23808 17552 23814 17604
rect 23952 17601 23980 17632
rect 26418 17620 26424 17632
rect 26476 17620 26482 17672
rect 27448 17660 27476 17768
rect 27540 17768 29776 17796
rect 27540 17737 27568 17768
rect 27525 17731 27583 17737
rect 27525 17697 27537 17731
rect 27571 17697 27583 17731
rect 27525 17691 27583 17697
rect 27709 17731 27767 17737
rect 27709 17697 27721 17731
rect 27755 17697 27767 17731
rect 28169 17731 28227 17737
rect 28169 17728 28181 17731
rect 27709 17691 27767 17697
rect 27816 17700 28181 17728
rect 27724 17660 27752 17691
rect 27448 17632 27752 17660
rect 23937 17595 23995 17601
rect 23937 17561 23949 17595
rect 23983 17561 23995 17595
rect 23937 17555 23995 17561
rect 26602 17552 26608 17604
rect 26660 17592 26666 17604
rect 26660 17564 26705 17592
rect 26660 17552 26666 17564
rect 27062 17552 27068 17604
rect 27120 17592 27126 17604
rect 27706 17592 27712 17604
rect 27120 17564 27712 17592
rect 27120 17552 27126 17564
rect 27706 17552 27712 17564
rect 27764 17552 27770 17604
rect 24118 17524 24124 17536
rect 22152 17496 24124 17524
rect 22152 17484 22158 17496
rect 24118 17484 24124 17496
rect 24176 17524 24182 17536
rect 24302 17524 24308 17536
rect 24176 17496 24308 17524
rect 24176 17484 24182 17496
rect 24302 17484 24308 17496
rect 24360 17484 24366 17536
rect 25222 17484 25228 17536
rect 25280 17524 25286 17536
rect 27816 17524 27844 17700
rect 28169 17697 28181 17700
rect 28215 17697 28227 17731
rect 28169 17691 28227 17697
rect 28626 17688 28632 17740
rect 28684 17728 28690 17740
rect 28810 17728 28816 17740
rect 28684 17700 28816 17728
rect 28684 17688 28690 17700
rect 28810 17688 28816 17700
rect 28868 17728 28874 17740
rect 29748 17737 29776 17768
rect 30009 17765 30021 17799
rect 30055 17796 30067 17799
rect 30190 17796 30196 17808
rect 30055 17768 30196 17796
rect 30055 17765 30067 17768
rect 30009 17759 30067 17765
rect 30190 17756 30196 17768
rect 30248 17756 30254 17808
rect 31404 17768 33732 17796
rect 29273 17731 29331 17737
rect 29273 17728 29285 17731
rect 28868 17700 29285 17728
rect 28868 17688 28874 17700
rect 29273 17697 29285 17700
rect 29319 17697 29331 17731
rect 29273 17691 29331 17697
rect 29733 17731 29791 17737
rect 29733 17697 29745 17731
rect 29779 17697 29791 17731
rect 31110 17728 31116 17740
rect 31071 17700 31116 17728
rect 29733 17691 29791 17697
rect 29086 17660 29092 17672
rect 29047 17632 29092 17660
rect 29086 17620 29092 17632
rect 29144 17620 29150 17672
rect 29748 17660 29776 17691
rect 31110 17688 31116 17700
rect 31168 17688 31174 17740
rect 31404 17737 31432 17768
rect 33704 17740 33732 17768
rect 34514 17756 34520 17808
rect 34572 17796 34578 17808
rect 36446 17796 36452 17808
rect 34572 17768 35664 17796
rect 34572 17756 34578 17768
rect 31389 17731 31447 17737
rect 31389 17697 31401 17731
rect 31435 17697 31447 17731
rect 32306 17728 32312 17740
rect 32267 17700 32312 17728
rect 31389 17691 31447 17697
rect 32306 17688 32312 17700
rect 32364 17688 32370 17740
rect 32674 17728 32680 17740
rect 32635 17700 32680 17728
rect 32674 17688 32680 17700
rect 32732 17688 32738 17740
rect 33505 17731 33563 17737
rect 33505 17697 33517 17731
rect 33551 17728 33563 17731
rect 33594 17728 33600 17740
rect 33551 17700 33600 17728
rect 33551 17697 33563 17700
rect 33505 17691 33563 17697
rect 33594 17688 33600 17700
rect 33652 17688 33658 17740
rect 33686 17688 33692 17740
rect 33744 17688 33750 17740
rect 34606 17728 34612 17740
rect 34567 17700 34612 17728
rect 34606 17688 34612 17700
rect 34664 17688 34670 17740
rect 34790 17728 34796 17740
rect 34751 17700 34796 17728
rect 34790 17688 34796 17700
rect 34848 17688 34854 17740
rect 35636 17737 35664 17768
rect 36280 17768 36452 17796
rect 36280 17737 36308 17768
rect 36446 17756 36452 17768
rect 36504 17756 36510 17808
rect 35345 17731 35403 17737
rect 35345 17697 35357 17731
rect 35391 17697 35403 17731
rect 35345 17691 35403 17697
rect 35621 17731 35679 17737
rect 35621 17697 35633 17731
rect 35667 17697 35679 17731
rect 35621 17691 35679 17697
rect 36265 17731 36323 17737
rect 36265 17697 36277 17731
rect 36311 17697 36323 17731
rect 36265 17691 36323 17697
rect 29748 17632 29868 17660
rect 25280 17496 27844 17524
rect 29840 17524 29868 17632
rect 30006 17620 30012 17672
rect 30064 17660 30070 17672
rect 30190 17660 30196 17672
rect 30064 17632 30196 17660
rect 30064 17620 30070 17632
rect 30190 17620 30196 17632
rect 30248 17620 30254 17672
rect 35360 17592 35388 17691
rect 36354 17688 36360 17740
rect 36412 17728 36418 17740
rect 36817 17731 36875 17737
rect 36817 17728 36829 17731
rect 36412 17700 36829 17728
rect 36412 17688 36418 17700
rect 36817 17697 36829 17700
rect 36863 17697 36875 17731
rect 36817 17691 36875 17697
rect 38289 17731 38347 17737
rect 38289 17697 38301 17731
rect 38335 17697 38347 17731
rect 38562 17728 38568 17740
rect 38523 17700 38568 17728
rect 38289 17691 38347 17697
rect 35802 17620 35808 17672
rect 35860 17660 35866 17672
rect 37829 17663 37887 17669
rect 37829 17660 37841 17663
rect 35860 17632 37841 17660
rect 35860 17620 35866 17632
rect 37829 17629 37841 17632
rect 37875 17629 37887 17663
rect 38304 17660 38332 17691
rect 38562 17688 38568 17700
rect 38620 17688 38626 17740
rect 38838 17660 38844 17672
rect 38304 17632 38844 17660
rect 37829 17623 37887 17629
rect 38838 17620 38844 17632
rect 38896 17620 38902 17672
rect 35360 17564 36492 17592
rect 32490 17524 32496 17536
rect 29840 17496 32496 17524
rect 25280 17484 25286 17496
rect 32490 17484 32496 17496
rect 32548 17524 32554 17536
rect 34790 17524 34796 17536
rect 32548 17496 34796 17524
rect 32548 17484 32554 17496
rect 34790 17484 34796 17496
rect 34848 17524 34854 17536
rect 35526 17524 35532 17536
rect 34848 17496 35532 17524
rect 34848 17484 34854 17496
rect 35526 17484 35532 17496
rect 35584 17484 35590 17536
rect 35710 17524 35716 17536
rect 35671 17496 35716 17524
rect 35710 17484 35716 17496
rect 35768 17484 35774 17536
rect 36262 17484 36268 17536
rect 36320 17524 36326 17536
rect 36357 17527 36415 17533
rect 36357 17524 36369 17527
rect 36320 17496 36369 17524
rect 36320 17484 36326 17496
rect 36357 17493 36369 17496
rect 36403 17493 36415 17527
rect 36464 17524 36492 17564
rect 36538 17552 36544 17604
rect 36596 17592 36602 17604
rect 38565 17595 38623 17601
rect 38565 17592 38577 17595
rect 36596 17564 38577 17592
rect 36596 17552 36602 17564
rect 38565 17561 38577 17564
rect 38611 17561 38623 17595
rect 38565 17555 38623 17561
rect 37550 17524 37556 17536
rect 36464 17496 37556 17524
rect 36357 17487 36415 17493
rect 37550 17484 37556 17496
rect 37608 17484 37614 17536
rect 1104 17434 39836 17456
rect 1104 17382 4246 17434
rect 4298 17382 4310 17434
rect 4362 17382 4374 17434
rect 4426 17382 4438 17434
rect 4490 17382 34966 17434
rect 35018 17382 35030 17434
rect 35082 17382 35094 17434
rect 35146 17382 35158 17434
rect 35210 17382 39836 17434
rect 1104 17360 39836 17382
rect 2774 17280 2780 17332
rect 2832 17320 2838 17332
rect 4706 17320 4712 17332
rect 2832 17292 4712 17320
rect 2832 17280 2838 17292
rect 4706 17280 4712 17292
rect 4764 17280 4770 17332
rect 6914 17320 6920 17332
rect 6875 17292 6920 17320
rect 6914 17280 6920 17292
rect 6972 17280 6978 17332
rect 9214 17320 9220 17332
rect 9175 17292 9220 17320
rect 9214 17280 9220 17292
rect 9272 17280 9278 17332
rect 10226 17320 10232 17332
rect 10187 17292 10232 17320
rect 10226 17280 10232 17292
rect 10284 17280 10290 17332
rect 11606 17320 11612 17332
rect 11567 17292 11612 17320
rect 11606 17280 11612 17292
rect 11664 17280 11670 17332
rect 14734 17280 14740 17332
rect 14792 17320 14798 17332
rect 14792 17292 15976 17320
rect 14792 17280 14798 17292
rect 10042 17212 10048 17264
rect 10100 17212 10106 17264
rect 13814 17252 13820 17264
rect 13464 17224 13820 17252
rect 3050 17184 3056 17196
rect 3011 17156 3056 17184
rect 3050 17144 3056 17156
rect 3108 17144 3114 17196
rect 4614 17184 4620 17196
rect 3252 17156 4620 17184
rect 1673 17119 1731 17125
rect 1673 17085 1685 17119
rect 1719 17116 1731 17119
rect 1946 17116 1952 17128
rect 1719 17088 1952 17116
rect 1719 17085 1731 17088
rect 1673 17079 1731 17085
rect 1946 17076 1952 17088
rect 2004 17076 2010 17128
rect 2222 17116 2228 17128
rect 2183 17088 2228 17116
rect 2222 17076 2228 17088
rect 2280 17076 2286 17128
rect 2409 17119 2467 17125
rect 2409 17085 2421 17119
rect 2455 17116 2467 17119
rect 2774 17116 2780 17128
rect 2455 17088 2780 17116
rect 2455 17085 2467 17088
rect 2409 17079 2467 17085
rect 2774 17076 2780 17088
rect 2832 17076 2838 17128
rect 3252 17125 3280 17156
rect 4614 17144 4620 17156
rect 4672 17144 4678 17196
rect 4706 17144 4712 17196
rect 4764 17184 4770 17196
rect 6178 17184 6184 17196
rect 4764 17156 5580 17184
rect 6139 17156 6184 17184
rect 4764 17144 4770 17156
rect 3237 17119 3295 17125
rect 3237 17085 3249 17119
rect 3283 17085 3295 17119
rect 3418 17116 3424 17128
rect 3379 17088 3424 17116
rect 3237 17079 3295 17085
rect 3418 17076 3424 17088
rect 3476 17076 3482 17128
rect 3970 17116 3976 17128
rect 3931 17088 3976 17116
rect 3970 17076 3976 17088
rect 4028 17076 4034 17128
rect 4890 17116 4896 17128
rect 4851 17088 4896 17116
rect 4890 17076 4896 17088
rect 4948 17076 4954 17128
rect 5442 17116 5448 17128
rect 5403 17088 5448 17116
rect 5442 17076 5448 17088
rect 5500 17076 5506 17128
rect 5552 17125 5580 17156
rect 6178 17144 6184 17156
rect 6236 17144 6242 17196
rect 9953 17187 10011 17193
rect 9953 17153 9965 17187
rect 9999 17184 10011 17187
rect 10060 17184 10088 17212
rect 9999 17156 10088 17184
rect 9999 17153 10011 17156
rect 9953 17147 10011 17153
rect 11238 17144 11244 17196
rect 11296 17184 11302 17196
rect 11333 17187 11391 17193
rect 11333 17184 11345 17187
rect 11296 17156 11345 17184
rect 11296 17144 11302 17156
rect 11333 17153 11345 17156
rect 11379 17153 11391 17187
rect 11333 17147 11391 17153
rect 5537 17119 5595 17125
rect 5537 17085 5549 17119
rect 5583 17085 5595 17119
rect 6270 17116 6276 17128
rect 6231 17088 6276 17116
rect 5537 17079 5595 17085
rect 6270 17076 6276 17088
rect 6328 17116 6334 17128
rect 6825 17119 6883 17125
rect 6825 17116 6837 17119
rect 6328 17088 6837 17116
rect 6328 17076 6334 17088
rect 6825 17085 6837 17088
rect 6871 17085 6883 17119
rect 7834 17116 7840 17128
rect 7795 17088 7840 17116
rect 6825 17079 6883 17085
rect 7834 17076 7840 17088
rect 7892 17076 7898 17128
rect 8113 17119 8171 17125
rect 8113 17085 8125 17119
rect 8159 17116 8171 17119
rect 8570 17116 8576 17128
rect 8159 17088 8576 17116
rect 8159 17085 8171 17088
rect 8113 17079 8171 17085
rect 8570 17076 8576 17088
rect 8628 17076 8634 17128
rect 10045 17119 10103 17125
rect 10045 17085 10057 17119
rect 10091 17116 10103 17119
rect 10686 17116 10692 17128
rect 10091 17088 10692 17116
rect 10091 17085 10103 17088
rect 10045 17079 10103 17085
rect 10686 17076 10692 17088
rect 10744 17076 10750 17128
rect 11422 17076 11428 17128
rect 11480 17116 11486 17128
rect 12710 17116 12716 17128
rect 11480 17088 11525 17116
rect 12671 17088 12716 17116
rect 11480 17076 11486 17088
rect 12710 17076 12716 17088
rect 12768 17076 12774 17128
rect 12894 17116 12900 17128
rect 12855 17088 12900 17116
rect 12894 17076 12900 17088
rect 12952 17076 12958 17128
rect 13464 17125 13492 17224
rect 13814 17212 13820 17224
rect 13872 17252 13878 17264
rect 15838 17252 15844 17264
rect 13872 17224 15516 17252
rect 15799 17224 15844 17252
rect 13872 17212 13878 17224
rect 13630 17184 13636 17196
rect 13591 17156 13636 17184
rect 13630 17144 13636 17156
rect 13688 17144 13694 17196
rect 15286 17184 15292 17196
rect 14200 17156 15292 17184
rect 14200 17125 14228 17156
rect 15286 17144 15292 17156
rect 15344 17144 15350 17196
rect 13449 17119 13507 17125
rect 13449 17085 13461 17119
rect 13495 17085 13507 17119
rect 13449 17079 13507 17085
rect 14185 17119 14243 17125
rect 14185 17085 14197 17119
rect 14231 17085 14243 17119
rect 14918 17116 14924 17128
rect 14879 17088 14924 17116
rect 14185 17079 14243 17085
rect 14918 17076 14924 17088
rect 14976 17076 14982 17128
rect 15194 17076 15200 17128
rect 15252 17116 15258 17128
rect 15381 17119 15439 17125
rect 15381 17116 15393 17119
rect 15252 17088 15393 17116
rect 15252 17076 15258 17088
rect 15381 17085 15393 17088
rect 15427 17085 15439 17119
rect 15488 17116 15516 17224
rect 15838 17212 15844 17224
rect 15896 17212 15902 17264
rect 15948 17252 15976 17292
rect 16114 17280 16120 17332
rect 16172 17320 16178 17332
rect 16577 17323 16635 17329
rect 16577 17320 16589 17323
rect 16172 17292 16589 17320
rect 16172 17280 16178 17292
rect 16577 17289 16589 17292
rect 16623 17289 16635 17323
rect 23474 17320 23480 17332
rect 16577 17283 16635 17289
rect 19812 17292 23480 17320
rect 18233 17255 18291 17261
rect 18233 17252 18245 17255
rect 15948 17224 18245 17252
rect 18233 17221 18245 17224
rect 18279 17252 18291 17255
rect 18598 17252 18604 17264
rect 18279 17224 18604 17252
rect 18279 17221 18291 17224
rect 18233 17215 18291 17221
rect 18598 17212 18604 17224
rect 18656 17212 18662 17264
rect 18690 17144 18696 17196
rect 18748 17184 18754 17196
rect 18877 17187 18935 17193
rect 18877 17184 18889 17187
rect 18748 17156 18889 17184
rect 18748 17144 18754 17156
rect 18877 17153 18889 17156
rect 18923 17153 18935 17187
rect 19150 17184 19156 17196
rect 19111 17156 19156 17184
rect 18877 17147 18935 17153
rect 19150 17144 19156 17156
rect 19208 17144 19214 17196
rect 15749 17119 15807 17125
rect 15749 17116 15761 17119
rect 15488 17088 15761 17116
rect 15381 17079 15439 17085
rect 15749 17085 15761 17088
rect 15795 17085 15807 17119
rect 16666 17116 16672 17128
rect 16627 17088 16672 17116
rect 15749 17079 15807 17085
rect 16666 17076 16672 17088
rect 16724 17076 16730 17128
rect 17218 17116 17224 17128
rect 17179 17088 17224 17116
rect 17218 17076 17224 17088
rect 17276 17076 17282 17128
rect 18049 17119 18107 17125
rect 18049 17085 18061 17119
rect 18095 17116 18107 17119
rect 18138 17116 18144 17128
rect 18095 17088 18144 17116
rect 18095 17085 18107 17088
rect 18049 17079 18107 17085
rect 18138 17076 18144 17088
rect 18196 17116 18202 17128
rect 19812 17116 19840 17292
rect 23474 17280 23480 17292
rect 23532 17280 23538 17332
rect 26510 17280 26516 17332
rect 26568 17320 26574 17332
rect 27433 17323 27491 17329
rect 27433 17320 27445 17323
rect 26568 17292 27445 17320
rect 26568 17280 26574 17292
rect 27433 17289 27445 17292
rect 27479 17289 27491 17323
rect 27433 17283 27491 17289
rect 27522 17280 27528 17332
rect 27580 17320 27586 17332
rect 28350 17320 28356 17332
rect 27580 17292 28356 17320
rect 27580 17280 27586 17292
rect 28350 17280 28356 17292
rect 28408 17320 28414 17332
rect 28408 17292 33088 17320
rect 28408 17280 28414 17292
rect 22646 17252 22652 17264
rect 22607 17224 22652 17252
rect 22646 17212 22652 17224
rect 22704 17212 22710 17264
rect 24026 17212 24032 17264
rect 24084 17252 24090 17264
rect 25682 17252 25688 17264
rect 24084 17224 25688 17252
rect 24084 17212 24090 17224
rect 25682 17212 25688 17224
rect 25740 17212 25746 17264
rect 31573 17255 31631 17261
rect 31573 17221 31585 17255
rect 31619 17221 31631 17255
rect 33060 17252 33088 17292
rect 33134 17280 33140 17332
rect 33192 17320 33198 17332
rect 33505 17323 33563 17329
rect 33505 17320 33517 17323
rect 33192 17292 33517 17320
rect 33192 17280 33198 17292
rect 33505 17289 33517 17292
rect 33551 17289 33563 17323
rect 33505 17283 33563 17289
rect 34606 17280 34612 17332
rect 34664 17320 34670 17332
rect 38102 17320 38108 17332
rect 34664 17292 38108 17320
rect 34664 17280 34670 17292
rect 38102 17280 38108 17292
rect 38160 17320 38166 17332
rect 38562 17320 38568 17332
rect 38160 17292 38568 17320
rect 38160 17280 38166 17292
rect 38562 17280 38568 17292
rect 38620 17320 38626 17332
rect 38841 17323 38899 17329
rect 38841 17320 38853 17323
rect 38620 17292 38853 17320
rect 38620 17280 38626 17292
rect 38841 17289 38853 17292
rect 38887 17289 38899 17323
rect 38841 17283 38899 17289
rect 34330 17252 34336 17264
rect 33060 17224 34336 17252
rect 31573 17215 31631 17221
rect 21358 17144 21364 17196
rect 21416 17184 21422 17196
rect 22738 17184 22744 17196
rect 21416 17156 22744 17184
rect 21416 17144 21422 17156
rect 18196 17088 19840 17116
rect 21545 17119 21603 17125
rect 18196 17076 18202 17088
rect 21545 17085 21557 17119
rect 21591 17116 21603 17119
rect 21634 17116 21640 17128
rect 21591 17088 21640 17116
rect 21591 17085 21603 17088
rect 21545 17079 21603 17085
rect 21634 17076 21640 17088
rect 21692 17076 21698 17128
rect 21744 17125 21772 17156
rect 22738 17144 22744 17156
rect 22796 17144 22802 17196
rect 24486 17144 24492 17196
rect 24544 17184 24550 17196
rect 24544 17156 26556 17184
rect 24544 17144 24550 17156
rect 21729 17119 21787 17125
rect 21729 17085 21741 17119
rect 21775 17116 21787 17119
rect 21775 17088 21809 17116
rect 21775 17085 21787 17088
rect 21729 17079 21787 17085
rect 22002 17076 22008 17128
rect 22060 17116 22066 17128
rect 22097 17119 22155 17125
rect 22097 17116 22109 17119
rect 22060 17088 22109 17116
rect 22060 17076 22066 17088
rect 22097 17085 22109 17088
rect 22143 17085 22155 17119
rect 22097 17079 22155 17085
rect 22186 17076 22192 17128
rect 22244 17116 22250 17128
rect 22465 17119 22523 17125
rect 22465 17116 22477 17119
rect 22244 17088 22477 17116
rect 22244 17076 22250 17088
rect 22465 17085 22477 17088
rect 22511 17085 22523 17119
rect 22465 17079 22523 17085
rect 23566 17076 23572 17128
rect 23624 17116 23630 17128
rect 24121 17119 24179 17125
rect 24121 17116 24133 17119
rect 23624 17088 24133 17116
rect 23624 17076 23630 17088
rect 24121 17085 24133 17088
rect 24167 17085 24179 17119
rect 24121 17079 24179 17085
rect 24394 17076 24400 17128
rect 24452 17116 24458 17128
rect 24857 17119 24915 17125
rect 24857 17116 24869 17119
rect 24452 17088 24869 17116
rect 24452 17076 24458 17088
rect 24857 17085 24869 17088
rect 24903 17116 24915 17119
rect 26142 17116 26148 17128
rect 24903 17088 25636 17116
rect 26103 17088 26148 17116
rect 24903 17085 24915 17088
rect 24857 17079 24915 17085
rect 3436 17048 3464 17076
rect 6546 17048 6552 17060
rect 3436 17020 6552 17048
rect 6546 17008 6552 17020
rect 6604 17008 6610 17060
rect 15470 17048 15476 17060
rect 13464 17020 15476 17048
rect 1673 16983 1731 16989
rect 1673 16949 1685 16983
rect 1719 16980 1731 16983
rect 1762 16980 1768 16992
rect 1719 16952 1768 16980
rect 1719 16949 1731 16952
rect 1673 16943 1731 16949
rect 1762 16940 1768 16952
rect 1820 16940 1826 16992
rect 11238 16940 11244 16992
rect 11296 16980 11302 16992
rect 13464 16980 13492 17020
rect 15470 17008 15476 17020
rect 15528 17048 15534 17060
rect 17402 17048 17408 17060
rect 15528 17020 17408 17048
rect 15528 17008 15534 17020
rect 17402 17008 17408 17020
rect 17460 17008 17466 17060
rect 20162 17008 20168 17060
rect 20220 17048 20226 17060
rect 25501 17051 25559 17057
rect 25501 17048 25513 17051
rect 20220 17020 25513 17048
rect 20220 17008 20226 17020
rect 25501 17017 25513 17020
rect 25547 17017 25559 17051
rect 25608 17048 25636 17088
rect 26142 17076 26148 17088
rect 26200 17076 26206 17128
rect 26234 17076 26240 17128
rect 26292 17116 26298 17128
rect 26528 17125 26556 17156
rect 26786 17144 26792 17196
rect 26844 17184 26850 17196
rect 26844 17156 28488 17184
rect 26844 17144 26850 17156
rect 28460 17128 28488 17156
rect 28810 17144 28816 17196
rect 28868 17184 28874 17196
rect 31588 17184 31616 17215
rect 34330 17212 34336 17224
rect 34388 17212 34394 17264
rect 32398 17184 32404 17196
rect 28868 17156 30512 17184
rect 31588 17156 32260 17184
rect 32359 17156 32404 17184
rect 28868 17144 28874 17156
rect 26513 17119 26571 17125
rect 26292 17088 26337 17116
rect 26292 17076 26298 17088
rect 26513 17085 26525 17119
rect 26559 17085 26571 17119
rect 26513 17079 26571 17085
rect 26697 17119 26755 17125
rect 26697 17085 26709 17119
rect 26743 17116 26755 17119
rect 27522 17116 27528 17128
rect 26743 17088 27528 17116
rect 26743 17085 26755 17088
rect 26697 17079 26755 17085
rect 27522 17076 27528 17088
rect 27580 17076 27586 17128
rect 27982 17116 27988 17128
rect 27943 17088 27988 17116
rect 27982 17076 27988 17088
rect 28040 17076 28046 17128
rect 28074 17076 28080 17128
rect 28132 17116 28138 17128
rect 28353 17119 28411 17125
rect 28132 17088 28177 17116
rect 28132 17076 28138 17088
rect 28353 17085 28365 17119
rect 28399 17085 28411 17119
rect 28353 17079 28411 17085
rect 27430 17048 27436 17060
rect 25608 17020 27436 17048
rect 25501 17011 25559 17017
rect 27430 17008 27436 17020
rect 27488 17008 27494 17060
rect 27706 17008 27712 17060
rect 27764 17048 27770 17060
rect 28368 17048 28396 17079
rect 28442 17076 28448 17128
rect 28500 17116 28506 17128
rect 29546 17116 29552 17128
rect 28500 17088 28545 17116
rect 29507 17088 29552 17116
rect 28500 17076 28506 17088
rect 29546 17076 29552 17088
rect 29604 17076 29610 17128
rect 30006 17116 30012 17128
rect 29967 17088 30012 17116
rect 30006 17076 30012 17088
rect 30064 17076 30070 17128
rect 30282 17116 30288 17128
rect 30243 17088 30288 17116
rect 30282 17076 30288 17088
rect 30340 17076 30346 17128
rect 30484 17125 30512 17156
rect 30469 17119 30527 17125
rect 30469 17085 30481 17119
rect 30515 17085 30527 17119
rect 30469 17079 30527 17085
rect 31389 17119 31447 17125
rect 31389 17085 31401 17119
rect 31435 17116 31447 17119
rect 31938 17116 31944 17128
rect 31435 17088 31944 17116
rect 31435 17085 31447 17088
rect 31389 17079 31447 17085
rect 31938 17076 31944 17088
rect 31996 17076 32002 17128
rect 32122 17116 32128 17128
rect 32083 17088 32128 17116
rect 32122 17076 32128 17088
rect 32180 17076 32186 17128
rect 32232 17116 32260 17156
rect 32398 17144 32404 17156
rect 32456 17144 32462 17196
rect 35802 17184 35808 17196
rect 34256 17156 35808 17184
rect 32766 17116 32772 17128
rect 32232 17088 32772 17116
rect 32766 17076 32772 17088
rect 32824 17116 32830 17128
rect 34256 17116 34284 17156
rect 35802 17144 35808 17156
rect 35860 17144 35866 17196
rect 35989 17187 36047 17193
rect 35989 17153 36001 17187
rect 36035 17184 36047 17187
rect 36354 17184 36360 17196
rect 36035 17156 36360 17184
rect 36035 17153 36047 17156
rect 35989 17147 36047 17153
rect 36354 17144 36360 17156
rect 36412 17144 36418 17196
rect 37182 17184 37188 17196
rect 36556 17156 37188 17184
rect 32824 17088 34284 17116
rect 32824 17076 32830 17088
rect 34514 17076 34520 17128
rect 34572 17116 34578 17128
rect 34885 17119 34943 17125
rect 34885 17116 34897 17119
rect 34572 17088 34897 17116
rect 34572 17076 34578 17088
rect 34885 17085 34897 17088
rect 34931 17085 34943 17119
rect 35342 17116 35348 17128
rect 35303 17088 35348 17116
rect 34885 17079 34943 17085
rect 35342 17076 35348 17088
rect 35400 17076 35406 17128
rect 35710 17116 35716 17128
rect 35671 17088 35716 17116
rect 35710 17076 35716 17088
rect 35768 17076 35774 17128
rect 36078 17076 36084 17128
rect 36136 17116 36142 17128
rect 36556 17125 36584 17156
rect 37182 17144 37188 17156
rect 37240 17144 37246 17196
rect 36541 17119 36599 17125
rect 36541 17116 36553 17119
rect 36136 17088 36553 17116
rect 36136 17076 36142 17088
rect 36541 17085 36553 17088
rect 36587 17085 36599 17119
rect 36541 17079 36599 17085
rect 36817 17119 36875 17125
rect 36817 17085 36829 17119
rect 36863 17116 36875 17119
rect 37826 17116 37832 17128
rect 36863 17088 37832 17116
rect 36863 17085 36875 17088
rect 36817 17079 36875 17085
rect 37826 17076 37832 17088
rect 37884 17076 37890 17128
rect 38654 17116 38660 17128
rect 38615 17088 38660 17116
rect 38654 17076 38660 17088
rect 38712 17076 38718 17128
rect 27764 17020 28396 17048
rect 30300 17048 30328 17076
rect 30300 17020 32260 17048
rect 27764 17008 27770 17020
rect 11296 16952 13492 16980
rect 11296 16940 11302 16952
rect 13538 16940 13544 16992
rect 13596 16980 13602 16992
rect 14369 16983 14427 16989
rect 14369 16980 14381 16983
rect 13596 16952 14381 16980
rect 13596 16940 13602 16952
rect 14369 16949 14381 16952
rect 14415 16980 14427 16983
rect 17494 16980 17500 16992
rect 14415 16952 17500 16980
rect 14415 16949 14427 16952
rect 14369 16943 14427 16949
rect 17494 16940 17500 16952
rect 17552 16940 17558 16992
rect 20441 16983 20499 16989
rect 20441 16949 20453 16983
rect 20487 16980 20499 16983
rect 20622 16980 20628 16992
rect 20487 16952 20628 16980
rect 20487 16949 20499 16952
rect 20441 16943 20499 16949
rect 20622 16940 20628 16952
rect 20680 16940 20686 16992
rect 24302 16980 24308 16992
rect 24263 16952 24308 16980
rect 24302 16940 24308 16952
rect 24360 16980 24366 16992
rect 24762 16980 24768 16992
rect 24360 16952 24768 16980
rect 24360 16940 24366 16952
rect 24762 16940 24768 16952
rect 24820 16940 24826 16992
rect 24946 16980 24952 16992
rect 24907 16952 24952 16980
rect 24946 16940 24952 16952
rect 25004 16940 25010 16992
rect 25682 16940 25688 16992
rect 25740 16980 25746 16992
rect 27522 16980 27528 16992
rect 25740 16952 27528 16980
rect 25740 16940 25746 16952
rect 27522 16940 27528 16952
rect 27580 16940 27586 16992
rect 30374 16940 30380 16992
rect 30432 16980 30438 16992
rect 30469 16983 30527 16989
rect 30469 16980 30481 16983
rect 30432 16952 30481 16980
rect 30432 16940 30438 16952
rect 30469 16949 30481 16952
rect 30515 16949 30527 16983
rect 32232 16980 32260 17020
rect 33962 16980 33968 16992
rect 32232 16952 33968 16980
rect 30469 16943 30527 16949
rect 33962 16940 33968 16952
rect 34020 16980 34026 16992
rect 34606 16980 34612 16992
rect 34020 16952 34612 16980
rect 34020 16940 34026 16952
rect 34606 16940 34612 16952
rect 34664 16940 34670 16992
rect 36446 16940 36452 16992
rect 36504 16980 36510 16992
rect 37921 16983 37979 16989
rect 37921 16980 37933 16983
rect 36504 16952 37933 16980
rect 36504 16940 36510 16952
rect 37921 16949 37933 16952
rect 37967 16949 37979 16983
rect 37921 16943 37979 16949
rect 1104 16890 39836 16912
rect 1104 16838 19606 16890
rect 19658 16838 19670 16890
rect 19722 16838 19734 16890
rect 19786 16838 19798 16890
rect 19850 16838 39836 16890
rect 1104 16816 39836 16838
rect 3421 16779 3479 16785
rect 3421 16745 3433 16779
rect 3467 16776 3479 16779
rect 4798 16776 4804 16788
rect 3467 16748 4804 16776
rect 3467 16745 3479 16748
rect 3421 16739 3479 16745
rect 4798 16736 4804 16748
rect 4856 16736 4862 16788
rect 5350 16736 5356 16788
rect 5408 16776 5414 16788
rect 5445 16779 5503 16785
rect 5445 16776 5457 16779
rect 5408 16748 5457 16776
rect 5408 16736 5414 16748
rect 5445 16745 5457 16748
rect 5491 16745 5503 16779
rect 8202 16776 8208 16788
rect 5445 16739 5503 16745
rect 8036 16748 8208 16776
rect 8036 16717 8064 16748
rect 8202 16736 8208 16748
rect 8260 16736 8266 16788
rect 11422 16736 11428 16788
rect 11480 16776 11486 16788
rect 11517 16779 11575 16785
rect 11517 16776 11529 16779
rect 11480 16748 11529 16776
rect 11480 16736 11486 16748
rect 11517 16745 11529 16748
rect 11563 16745 11575 16779
rect 11517 16739 11575 16745
rect 12710 16736 12716 16788
rect 12768 16776 12774 16788
rect 12768 16748 13768 16776
rect 12768 16736 12774 16748
rect 2777 16711 2835 16717
rect 2777 16677 2789 16711
rect 2823 16708 2835 16711
rect 8021 16711 8079 16717
rect 2823 16680 4016 16708
rect 2823 16677 2835 16680
rect 2777 16671 2835 16677
rect 2585 16643 2643 16649
rect 2585 16609 2597 16643
rect 2631 16609 2643 16643
rect 2585 16603 2643 16609
rect 2685 16643 2743 16649
rect 2685 16609 2697 16643
rect 2731 16640 2743 16643
rect 3050 16640 3056 16652
rect 2731 16612 3056 16640
rect 2731 16609 2743 16612
rect 2685 16603 2743 16609
rect 2608 16572 2636 16603
rect 3050 16600 3056 16612
rect 3108 16600 3114 16652
rect 3326 16640 3332 16652
rect 3287 16612 3332 16640
rect 3326 16600 3332 16612
rect 3384 16600 3390 16652
rect 3988 16640 4016 16680
rect 8021 16677 8033 16711
rect 8067 16677 8079 16711
rect 8570 16708 8576 16720
rect 8531 16680 8576 16708
rect 8021 16671 8079 16677
rect 8570 16668 8576 16680
rect 8628 16668 8634 16720
rect 13740 16708 13768 16748
rect 13998 16736 14004 16788
rect 14056 16776 14062 16788
rect 14185 16779 14243 16785
rect 14185 16776 14197 16779
rect 14056 16748 14197 16776
rect 14056 16736 14062 16748
rect 14185 16745 14197 16748
rect 14231 16745 14243 16779
rect 18601 16779 18659 16785
rect 18601 16776 18613 16779
rect 14185 16739 14243 16745
rect 14292 16748 18613 16776
rect 14292 16708 14320 16748
rect 18601 16745 18613 16748
rect 18647 16776 18659 16779
rect 19978 16776 19984 16788
rect 18647 16748 19984 16776
rect 18647 16745 18659 16748
rect 18601 16739 18659 16745
rect 19978 16736 19984 16748
rect 20036 16736 20042 16788
rect 20714 16736 20720 16788
rect 20772 16776 20778 16788
rect 21269 16779 21327 16785
rect 21269 16776 21281 16779
rect 20772 16748 21281 16776
rect 20772 16736 20778 16748
rect 21269 16745 21281 16748
rect 21315 16745 21327 16779
rect 21269 16739 21327 16745
rect 22002 16736 22008 16788
rect 22060 16776 22066 16788
rect 22060 16748 22508 16776
rect 22060 16736 22066 16748
rect 17862 16708 17868 16720
rect 13740 16680 14320 16708
rect 15120 16680 17868 16708
rect 4341 16643 4399 16649
rect 4341 16640 4353 16643
rect 3988 16612 4353 16640
rect 4341 16609 4353 16612
rect 4387 16609 4399 16643
rect 6178 16640 6184 16652
rect 6139 16612 6184 16640
rect 4341 16603 4399 16609
rect 6178 16600 6184 16612
rect 6236 16600 6242 16652
rect 6546 16640 6552 16652
rect 6507 16612 6552 16640
rect 6546 16600 6552 16612
rect 6604 16600 6610 16652
rect 7190 16640 7196 16652
rect 7151 16612 7196 16640
rect 7190 16600 7196 16612
rect 7248 16600 7254 16652
rect 7929 16643 7987 16649
rect 7929 16609 7941 16643
rect 7975 16609 7987 16643
rect 8110 16640 8116 16652
rect 8071 16612 8116 16640
rect 7929 16603 7987 16609
rect 3510 16572 3516 16584
rect 2608 16544 3516 16572
rect 3510 16532 3516 16544
rect 3568 16532 3574 16584
rect 4065 16575 4123 16581
rect 4065 16541 4077 16575
rect 4111 16541 4123 16575
rect 4065 16535 4123 16541
rect 3970 16464 3976 16516
rect 4028 16504 4034 16516
rect 4080 16504 4108 16535
rect 4430 16532 4436 16584
rect 4488 16572 4494 16584
rect 6273 16575 6331 16581
rect 6273 16572 6285 16575
rect 4488 16544 6285 16572
rect 4488 16532 4494 16544
rect 6273 16541 6285 16544
rect 6319 16541 6331 16575
rect 7944 16572 7972 16603
rect 8110 16600 8116 16612
rect 8168 16600 8174 16652
rect 8386 16640 8392 16652
rect 8220 16612 8392 16640
rect 8220 16572 8248 16612
rect 8386 16600 8392 16612
rect 8444 16600 8450 16652
rect 9950 16600 9956 16652
rect 10008 16640 10014 16652
rect 10137 16643 10195 16649
rect 10137 16640 10149 16643
rect 10008 16612 10149 16640
rect 10008 16600 10014 16612
rect 10137 16609 10149 16612
rect 10183 16609 10195 16643
rect 10137 16603 10195 16609
rect 10413 16643 10471 16649
rect 10413 16609 10425 16643
rect 10459 16640 10471 16643
rect 15120 16640 15148 16680
rect 17862 16668 17868 16680
rect 17920 16668 17926 16720
rect 22480 16708 22508 16748
rect 28994 16736 29000 16788
rect 29052 16776 29058 16788
rect 33686 16776 33692 16788
rect 29052 16748 32168 16776
rect 29052 16736 29058 16748
rect 24026 16708 24032 16720
rect 19812 16680 22416 16708
rect 22480 16680 24032 16708
rect 15470 16640 15476 16652
rect 10459 16612 15148 16640
rect 15431 16612 15476 16640
rect 10459 16609 10471 16612
rect 10413 16603 10471 16609
rect 15470 16600 15476 16612
rect 15528 16600 15534 16652
rect 15565 16643 15623 16649
rect 15565 16609 15577 16643
rect 15611 16640 15623 16643
rect 16298 16640 16304 16652
rect 15611 16612 16304 16640
rect 15611 16609 15623 16612
rect 15565 16603 15623 16609
rect 16298 16600 16304 16612
rect 16356 16600 16362 16652
rect 17405 16643 17463 16649
rect 17405 16609 17417 16643
rect 17451 16640 17463 16643
rect 17494 16640 17500 16652
rect 17451 16612 17500 16640
rect 17451 16609 17463 16612
rect 17405 16603 17463 16609
rect 17494 16600 17500 16612
rect 17552 16600 17558 16652
rect 17678 16640 17684 16652
rect 17639 16612 17684 16640
rect 17678 16600 17684 16612
rect 17736 16600 17742 16652
rect 18414 16640 18420 16652
rect 18375 16612 18420 16640
rect 18414 16600 18420 16612
rect 18472 16600 18478 16652
rect 18506 16600 18512 16652
rect 18564 16640 18570 16652
rect 19812 16649 19840 16680
rect 19153 16643 19211 16649
rect 19153 16640 19165 16643
rect 18564 16612 19165 16640
rect 18564 16600 18570 16612
rect 19153 16609 19165 16612
rect 19199 16609 19211 16643
rect 19153 16603 19211 16609
rect 19797 16643 19855 16649
rect 19797 16609 19809 16643
rect 19843 16609 19855 16643
rect 20162 16640 20168 16652
rect 20123 16612 20168 16640
rect 19797 16603 19855 16609
rect 20162 16600 20168 16612
rect 20220 16600 20226 16652
rect 21453 16643 21511 16649
rect 21453 16609 21465 16643
rect 21499 16640 21511 16643
rect 21634 16640 21640 16652
rect 21499 16612 21640 16640
rect 21499 16609 21511 16612
rect 21453 16603 21511 16609
rect 21634 16600 21640 16612
rect 21692 16600 21698 16652
rect 22002 16640 22008 16652
rect 21915 16612 22008 16640
rect 22002 16600 22008 16612
rect 22060 16600 22066 16652
rect 7944 16544 8248 16572
rect 6273 16535 6331 16541
rect 12526 16532 12532 16584
rect 12584 16572 12590 16584
rect 12805 16575 12863 16581
rect 12805 16572 12817 16575
rect 12584 16544 12817 16572
rect 12584 16532 12590 16544
rect 12805 16541 12817 16544
rect 12851 16541 12863 16575
rect 13078 16572 13084 16584
rect 13039 16544 13084 16572
rect 12805 16535 12863 16541
rect 13078 16532 13084 16544
rect 13136 16532 13142 16584
rect 15286 16532 15292 16584
rect 15344 16572 15350 16584
rect 16945 16575 17003 16581
rect 16945 16572 16957 16575
rect 15344 16544 16957 16572
rect 15344 16532 15350 16544
rect 16945 16541 16957 16544
rect 16991 16572 17003 16575
rect 17034 16572 17040 16584
rect 16991 16544 17040 16572
rect 16991 16541 17003 16544
rect 16945 16535 17003 16541
rect 17034 16532 17040 16544
rect 17092 16532 17098 16584
rect 17957 16575 18015 16581
rect 17957 16541 17969 16575
rect 18003 16572 18015 16575
rect 18322 16572 18328 16584
rect 18003 16544 18328 16572
rect 18003 16541 18015 16544
rect 17957 16535 18015 16541
rect 18322 16532 18328 16544
rect 18380 16532 18386 16584
rect 19334 16572 19340 16584
rect 19295 16544 19340 16572
rect 19334 16532 19340 16544
rect 19392 16532 19398 16584
rect 20714 16532 20720 16584
rect 20772 16572 20778 16584
rect 22020 16572 22048 16600
rect 20772 16544 22048 16572
rect 22097 16575 22155 16581
rect 20772 16532 20778 16544
rect 22097 16541 22109 16575
rect 22143 16572 22155 16575
rect 22388 16572 22416 16680
rect 24026 16668 24032 16680
rect 24084 16668 24090 16720
rect 24946 16668 24952 16720
rect 25004 16708 25010 16720
rect 32140 16717 32168 16748
rect 32968 16748 33692 16776
rect 32125 16711 32183 16717
rect 25004 16680 30880 16708
rect 25004 16668 25010 16680
rect 22738 16640 22744 16652
rect 22699 16612 22744 16640
rect 22738 16600 22744 16612
rect 22796 16600 22802 16652
rect 23750 16640 23756 16652
rect 23711 16612 23756 16640
rect 23750 16600 23756 16612
rect 23808 16600 23814 16652
rect 24305 16643 24363 16649
rect 24305 16609 24317 16643
rect 24351 16640 24363 16643
rect 24394 16640 24400 16652
rect 24351 16612 24400 16640
rect 24351 16609 24363 16612
rect 24305 16603 24363 16609
rect 24394 16600 24400 16612
rect 24452 16600 24458 16652
rect 24854 16640 24860 16652
rect 24815 16612 24860 16640
rect 24854 16600 24860 16612
rect 24912 16600 24918 16652
rect 25314 16640 25320 16652
rect 25275 16612 25320 16640
rect 25314 16600 25320 16612
rect 25372 16600 25378 16652
rect 25774 16640 25780 16652
rect 25735 16612 25780 16640
rect 25774 16600 25780 16612
rect 25832 16600 25838 16652
rect 25869 16643 25927 16649
rect 25869 16609 25881 16643
rect 25915 16640 25927 16643
rect 26786 16640 26792 16652
rect 25915 16612 26792 16640
rect 25915 16609 25927 16612
rect 25869 16603 25927 16609
rect 26786 16600 26792 16612
rect 26844 16600 26850 16652
rect 27062 16640 27068 16652
rect 27023 16612 27068 16640
rect 27062 16600 27068 16612
rect 27120 16600 27126 16652
rect 27249 16643 27307 16649
rect 27249 16609 27261 16643
rect 27295 16609 27307 16643
rect 27430 16640 27436 16652
rect 27391 16612 27436 16640
rect 27249 16603 27307 16609
rect 23768 16572 23796 16600
rect 24486 16572 24492 16584
rect 22143 16544 22324 16572
rect 22388 16544 23704 16572
rect 23768 16544 24492 16572
rect 22143 16541 22155 16544
rect 22097 16535 22155 16541
rect 21450 16504 21456 16516
rect 4028 16476 4108 16504
rect 13740 16476 21456 16504
rect 4028 16464 4034 16476
rect 1486 16396 1492 16448
rect 1544 16436 1550 16448
rect 2409 16439 2467 16445
rect 2409 16436 2421 16439
rect 1544 16408 2421 16436
rect 1544 16396 1550 16408
rect 2409 16405 2421 16408
rect 2455 16405 2467 16439
rect 2409 16399 2467 16405
rect 4062 16396 4068 16448
rect 4120 16436 4126 16448
rect 10042 16436 10048 16448
rect 4120 16408 10048 16436
rect 4120 16396 4126 16408
rect 10042 16396 10048 16408
rect 10100 16396 10106 16448
rect 10778 16396 10784 16448
rect 10836 16436 10842 16448
rect 13740 16436 13768 16476
rect 21450 16464 21456 16476
rect 21508 16464 21514 16516
rect 22296 16504 22324 16544
rect 22554 16504 22560 16516
rect 22296 16476 22560 16504
rect 22554 16464 22560 16476
rect 22612 16504 22618 16516
rect 22925 16507 22983 16513
rect 22925 16504 22937 16507
rect 22612 16476 22937 16504
rect 22612 16464 22618 16476
rect 22925 16473 22937 16476
rect 22971 16504 22983 16507
rect 23566 16504 23572 16516
rect 22971 16476 23572 16504
rect 22971 16473 22983 16476
rect 22925 16467 22983 16473
rect 23566 16464 23572 16476
rect 23624 16464 23630 16516
rect 23676 16513 23704 16544
rect 24486 16532 24492 16544
rect 24544 16532 24550 16584
rect 24670 16532 24676 16584
rect 24728 16572 24734 16584
rect 24765 16575 24823 16581
rect 24765 16572 24777 16575
rect 24728 16544 24777 16572
rect 24728 16532 24734 16544
rect 24765 16541 24777 16544
rect 24811 16572 24823 16575
rect 25038 16572 25044 16584
rect 24811 16544 25044 16572
rect 24811 16541 24823 16544
rect 24765 16535 24823 16541
rect 25038 16532 25044 16544
rect 25096 16532 25102 16584
rect 26602 16532 26608 16584
rect 26660 16572 26666 16584
rect 27264 16572 27292 16603
rect 27430 16600 27436 16612
rect 27488 16600 27494 16652
rect 27614 16600 27620 16652
rect 27672 16640 27678 16652
rect 28166 16640 28172 16652
rect 27672 16612 28172 16640
rect 27672 16600 27678 16612
rect 28166 16600 28172 16612
rect 28224 16600 28230 16652
rect 28350 16600 28356 16652
rect 28408 16640 28414 16652
rect 28629 16643 28687 16649
rect 28629 16640 28641 16643
rect 28408 16612 28641 16640
rect 28408 16600 28414 16612
rect 28629 16609 28641 16612
rect 28675 16609 28687 16643
rect 28810 16640 28816 16652
rect 28771 16612 28816 16640
rect 28629 16603 28687 16609
rect 28810 16600 28816 16612
rect 28868 16600 28874 16652
rect 28997 16643 29055 16649
rect 28997 16609 29009 16643
rect 29043 16640 29055 16643
rect 29086 16640 29092 16652
rect 29043 16612 29092 16640
rect 29043 16609 29055 16612
rect 28997 16603 29055 16609
rect 26660 16544 27292 16572
rect 26660 16532 26666 16544
rect 23661 16507 23719 16513
rect 23661 16473 23673 16507
rect 23707 16473 23719 16507
rect 23661 16467 23719 16473
rect 26881 16507 26939 16513
rect 26881 16473 26893 16507
rect 26927 16504 26939 16507
rect 27154 16504 27160 16516
rect 26927 16476 27160 16504
rect 26927 16473 26939 16476
rect 26881 16467 26939 16473
rect 27154 16464 27160 16476
rect 27212 16464 27218 16516
rect 29012 16504 29040 16603
rect 29086 16600 29092 16612
rect 29144 16600 29150 16652
rect 29181 16643 29239 16649
rect 29181 16609 29193 16643
rect 29227 16609 29239 16643
rect 29362 16640 29368 16652
rect 29323 16612 29368 16640
rect 29181 16603 29239 16609
rect 29196 16572 29224 16603
rect 29362 16600 29368 16612
rect 29420 16600 29426 16652
rect 30193 16643 30251 16649
rect 30193 16609 30205 16643
rect 30239 16640 30251 16643
rect 30239 16612 30328 16640
rect 30239 16609 30251 16612
rect 30193 16603 30251 16609
rect 29730 16572 29736 16584
rect 29196 16544 29736 16572
rect 29730 16532 29736 16544
rect 29788 16532 29794 16584
rect 30300 16572 30328 16612
rect 30374 16600 30380 16652
rect 30432 16640 30438 16652
rect 30852 16649 30880 16680
rect 32125 16677 32137 16711
rect 32171 16677 32183 16711
rect 32125 16671 32183 16677
rect 32214 16668 32220 16720
rect 32272 16708 32278 16720
rect 32968 16708 32996 16748
rect 33686 16736 33692 16748
rect 33744 16736 33750 16788
rect 34974 16776 34980 16788
rect 34935 16748 34980 16776
rect 34974 16736 34980 16748
rect 35032 16736 35038 16788
rect 35621 16779 35679 16785
rect 35621 16745 35633 16779
rect 35667 16776 35679 16779
rect 35986 16776 35992 16788
rect 35667 16748 35992 16776
rect 35667 16745 35679 16748
rect 35621 16739 35679 16745
rect 35986 16736 35992 16748
rect 36044 16736 36050 16788
rect 37829 16779 37887 16785
rect 37829 16745 37841 16779
rect 37875 16776 37887 16779
rect 38838 16776 38844 16788
rect 37875 16748 38844 16776
rect 37875 16745 37887 16748
rect 37829 16739 37887 16745
rect 38838 16736 38844 16748
rect 38896 16736 38902 16788
rect 34054 16708 34060 16720
rect 32272 16680 32996 16708
rect 32272 16668 32278 16680
rect 30837 16643 30895 16649
rect 30432 16612 30477 16640
rect 30432 16600 30438 16612
rect 30837 16609 30849 16643
rect 30883 16609 30895 16643
rect 30837 16603 30895 16609
rect 31110 16600 31116 16652
rect 31168 16640 31174 16652
rect 32968 16649 32996 16680
rect 33060 16680 34060 16708
rect 32815 16643 32873 16649
rect 32815 16640 32827 16643
rect 31168 16612 32827 16640
rect 31168 16600 31174 16612
rect 32815 16609 32827 16612
rect 32861 16609 32873 16643
rect 32815 16603 32873 16609
rect 32953 16643 33011 16649
rect 32953 16609 32965 16643
rect 32999 16609 33011 16643
rect 32953 16603 33011 16609
rect 30466 16572 30472 16584
rect 30300 16544 30472 16572
rect 30466 16532 30472 16544
rect 30524 16532 30530 16584
rect 32677 16575 32735 16581
rect 32677 16541 32689 16575
rect 32723 16572 32735 16575
rect 33060 16572 33088 16680
rect 34054 16668 34060 16680
rect 34112 16668 34118 16720
rect 34808 16680 37780 16708
rect 33226 16600 33232 16652
rect 33284 16640 33290 16652
rect 33597 16643 33655 16649
rect 33597 16640 33609 16643
rect 33284 16612 33609 16640
rect 33284 16600 33290 16612
rect 33597 16609 33609 16612
rect 33643 16609 33655 16643
rect 33597 16603 33655 16609
rect 34606 16600 34612 16652
rect 34664 16640 34670 16652
rect 34808 16649 34836 16680
rect 34793 16643 34851 16649
rect 34793 16640 34805 16643
rect 34664 16612 34805 16640
rect 34664 16600 34670 16612
rect 34793 16609 34805 16612
rect 34839 16609 34851 16643
rect 35618 16640 35624 16652
rect 35579 16612 35624 16640
rect 34793 16603 34851 16609
rect 35618 16600 35624 16612
rect 35676 16600 35682 16652
rect 36262 16640 36268 16652
rect 36223 16612 36268 16640
rect 36262 16600 36268 16612
rect 36320 16600 36326 16652
rect 36538 16640 36544 16652
rect 36499 16612 36544 16640
rect 36538 16600 36544 16612
rect 36596 16600 36602 16652
rect 37752 16649 37780 16680
rect 37737 16643 37795 16649
rect 37737 16609 37749 16643
rect 37783 16609 37795 16643
rect 37737 16603 37795 16609
rect 38289 16643 38347 16649
rect 38289 16609 38301 16643
rect 38335 16609 38347 16643
rect 38562 16640 38568 16652
rect 38523 16612 38568 16640
rect 38289 16603 38347 16609
rect 32723 16544 33088 16572
rect 32723 16541 32735 16544
rect 32677 16535 32735 16541
rect 33502 16532 33508 16584
rect 33560 16572 33566 16584
rect 36078 16572 36084 16584
rect 33560 16544 36084 16572
rect 33560 16532 33566 16544
rect 36078 16532 36084 16544
rect 36136 16532 36142 16584
rect 37550 16532 37556 16584
rect 37608 16572 37614 16584
rect 38304 16572 38332 16603
rect 38562 16600 38568 16612
rect 38620 16600 38626 16652
rect 37608 16544 38332 16572
rect 37608 16532 37614 16544
rect 30006 16504 30012 16516
rect 29012 16476 30012 16504
rect 30006 16464 30012 16476
rect 30064 16464 30070 16516
rect 30834 16504 30840 16516
rect 30795 16476 30840 16504
rect 30834 16464 30840 16476
rect 30892 16464 30898 16516
rect 36630 16504 36636 16516
rect 33428 16476 36636 16504
rect 10836 16408 13768 16436
rect 10836 16396 10842 16408
rect 15562 16396 15568 16448
rect 15620 16436 15626 16448
rect 15749 16439 15807 16445
rect 15749 16436 15761 16439
rect 15620 16408 15761 16436
rect 15620 16396 15626 16408
rect 15749 16405 15761 16408
rect 15795 16405 15807 16439
rect 15749 16399 15807 16405
rect 19334 16396 19340 16448
rect 19392 16436 19398 16448
rect 21174 16436 21180 16448
rect 19392 16408 21180 16436
rect 19392 16396 19398 16408
rect 21174 16396 21180 16408
rect 21232 16396 21238 16448
rect 23584 16436 23612 16464
rect 24210 16436 24216 16448
rect 23584 16408 24216 16436
rect 24210 16396 24216 16408
rect 24268 16436 24274 16448
rect 24670 16436 24676 16448
rect 24268 16408 24676 16436
rect 24268 16396 24274 16408
rect 24670 16396 24676 16408
rect 24728 16396 24734 16448
rect 28166 16436 28172 16448
rect 28127 16408 28172 16436
rect 28166 16396 28172 16408
rect 28224 16396 28230 16448
rect 28902 16396 28908 16448
rect 28960 16436 28966 16448
rect 33428 16436 33456 16476
rect 36630 16464 36636 16476
rect 36688 16464 36694 16516
rect 28960 16408 33456 16436
rect 28960 16396 28966 16408
rect 33502 16396 33508 16448
rect 33560 16436 33566 16448
rect 33781 16439 33839 16445
rect 33781 16436 33793 16439
rect 33560 16408 33793 16436
rect 33560 16396 33566 16408
rect 33781 16405 33793 16408
rect 33827 16436 33839 16439
rect 36354 16436 36360 16448
rect 33827 16408 36360 16436
rect 33827 16405 33839 16408
rect 33781 16399 33839 16405
rect 36354 16396 36360 16408
rect 36412 16396 36418 16448
rect 1104 16346 39836 16368
rect 1104 16294 4246 16346
rect 4298 16294 4310 16346
rect 4362 16294 4374 16346
rect 4426 16294 4438 16346
rect 4490 16294 34966 16346
rect 35018 16294 35030 16346
rect 35082 16294 35094 16346
rect 35146 16294 35158 16346
rect 35210 16294 39836 16346
rect 1104 16272 39836 16294
rect 2961 16235 3019 16241
rect 2961 16201 2973 16235
rect 3007 16232 3019 16235
rect 3142 16232 3148 16244
rect 3007 16204 3148 16232
rect 3007 16201 3019 16204
rect 2961 16195 3019 16201
rect 3142 16192 3148 16204
rect 3200 16192 3206 16244
rect 3970 16192 3976 16244
rect 4028 16232 4034 16244
rect 6181 16235 6239 16241
rect 4028 16204 5580 16232
rect 4028 16192 4034 16204
rect 3418 16056 3424 16108
rect 3476 16096 3482 16108
rect 4632 16105 4660 16204
rect 5552 16164 5580 16204
rect 6181 16201 6193 16235
rect 6227 16232 6239 16235
rect 6270 16232 6276 16244
rect 6227 16204 6276 16232
rect 6227 16201 6239 16204
rect 6181 16195 6239 16201
rect 6270 16192 6276 16204
rect 6328 16192 6334 16244
rect 7101 16235 7159 16241
rect 7101 16201 7113 16235
rect 7147 16232 7159 16235
rect 13722 16232 13728 16244
rect 7147 16204 13728 16232
rect 7147 16201 7159 16204
rect 7101 16195 7159 16201
rect 13722 16192 13728 16204
rect 13780 16192 13786 16244
rect 26510 16232 26516 16244
rect 21008 16204 26516 16232
rect 5552 16136 7880 16164
rect 7852 16108 7880 16136
rect 13078 16124 13084 16176
rect 13136 16164 13142 16176
rect 13541 16167 13599 16173
rect 13541 16164 13553 16167
rect 13136 16136 13553 16164
rect 13136 16124 13142 16136
rect 13541 16133 13553 16136
rect 13587 16133 13599 16167
rect 13541 16127 13599 16133
rect 3605 16099 3663 16105
rect 3605 16096 3617 16099
rect 3476 16068 3617 16096
rect 3476 16056 3482 16068
rect 3605 16065 3617 16068
rect 3651 16065 3663 16099
rect 3605 16059 3663 16065
rect 4617 16099 4675 16105
rect 4617 16065 4629 16099
rect 4663 16065 4675 16099
rect 4617 16059 4675 16065
rect 4798 16056 4804 16108
rect 4856 16096 4862 16108
rect 4893 16099 4951 16105
rect 4893 16096 4905 16099
rect 4856 16068 4905 16096
rect 4856 16056 4862 16068
rect 4893 16065 4905 16068
rect 4939 16065 4951 16099
rect 4893 16059 4951 16065
rect 6546 16056 6552 16108
rect 6604 16096 6610 16108
rect 6825 16099 6883 16105
rect 6825 16096 6837 16099
rect 6604 16068 6837 16096
rect 6604 16056 6610 16068
rect 6825 16065 6837 16068
rect 6871 16065 6883 16099
rect 6825 16059 6883 16065
rect 7834 16056 7840 16108
rect 7892 16096 7898 16108
rect 8389 16099 8447 16105
rect 8389 16096 8401 16099
rect 7892 16068 8401 16096
rect 7892 16056 7898 16068
rect 8389 16065 8401 16068
rect 8435 16065 8447 16099
rect 8389 16059 8447 16065
rect 10505 16099 10563 16105
rect 10505 16065 10517 16099
rect 10551 16096 10563 16099
rect 10778 16096 10784 16108
rect 10551 16068 10784 16096
rect 10551 16065 10563 16068
rect 10505 16059 10563 16065
rect 1397 16031 1455 16037
rect 1397 15997 1409 16031
rect 1443 16028 1455 16031
rect 1486 16028 1492 16040
rect 1443 16000 1492 16028
rect 1443 15997 1455 16000
rect 1397 15991 1455 15997
rect 1486 15988 1492 16000
rect 1544 15988 1550 16040
rect 1670 16028 1676 16040
rect 1631 16000 1676 16028
rect 1670 15988 1676 16000
rect 1728 15988 1734 16040
rect 3694 16028 3700 16040
rect 3655 16000 3700 16028
rect 3694 15988 3700 16000
rect 3752 15988 3758 16040
rect 5166 16028 5172 16040
rect 4724 16000 5172 16028
rect 4157 15963 4215 15969
rect 4157 15929 4169 15963
rect 4203 15960 4215 15963
rect 4724 15960 4752 16000
rect 5166 15988 5172 16000
rect 5224 15988 5230 16040
rect 6917 16031 6975 16037
rect 6917 15997 6929 16031
rect 6963 16028 6975 16031
rect 7006 16028 7012 16040
rect 6963 16000 7012 16028
rect 6963 15997 6975 16000
rect 6917 15991 6975 15997
rect 7006 15988 7012 16000
rect 7064 15988 7070 16040
rect 8662 16028 8668 16040
rect 8623 16000 8668 16028
rect 8662 15988 8668 16000
rect 8720 15988 8726 16040
rect 10520 16028 10548 16059
rect 10778 16056 10784 16068
rect 10836 16056 10842 16108
rect 11057 16099 11115 16105
rect 11057 16065 11069 16099
rect 11103 16096 11115 16099
rect 18322 16096 18328 16108
rect 11103 16068 18000 16096
rect 18283 16068 18328 16096
rect 11103 16065 11115 16068
rect 11057 16059 11115 16065
rect 9324 16000 10548 16028
rect 10597 16031 10655 16037
rect 4203 15932 4752 15960
rect 4203 15929 4215 15932
rect 4157 15923 4215 15929
rect 3786 15852 3792 15904
rect 3844 15892 3850 15904
rect 9324 15892 9352 16000
rect 10597 15997 10609 16031
rect 10643 15997 10655 16031
rect 11514 16028 11520 16040
rect 11475 16000 11520 16028
rect 10597 15991 10655 15997
rect 10045 15963 10103 15969
rect 10045 15929 10057 15963
rect 10091 15960 10103 15963
rect 10612 15960 10640 15991
rect 11514 15988 11520 16000
rect 11572 15988 11578 16040
rect 12894 15988 12900 16040
rect 12952 16028 12958 16040
rect 13078 16028 13084 16040
rect 12952 16000 13084 16028
rect 12952 15988 12958 16000
rect 13078 15988 13084 16000
rect 13136 15988 13142 16040
rect 13265 16031 13323 16037
rect 13265 15997 13277 16031
rect 13311 16028 13323 16031
rect 13538 16028 13544 16040
rect 13311 16000 13544 16028
rect 13311 15997 13323 16000
rect 13265 15991 13323 15997
rect 13538 15988 13544 16000
rect 13596 15988 13602 16040
rect 13633 16031 13691 16037
rect 13633 15997 13645 16031
rect 13679 16028 13691 16031
rect 13814 16028 13820 16040
rect 13679 16000 13820 16028
rect 13679 15997 13691 16000
rect 13633 15991 13691 15997
rect 13814 15988 13820 16000
rect 13872 15988 13878 16040
rect 14553 16031 14611 16037
rect 14553 15997 14565 16031
rect 14599 15997 14611 16031
rect 14826 16028 14832 16040
rect 14787 16000 14832 16028
rect 14553 15991 14611 15997
rect 10091 15932 10640 15960
rect 10091 15929 10103 15932
rect 10045 15923 10103 15929
rect 12526 15920 12532 15972
rect 12584 15960 12590 15972
rect 14568 15960 14596 15991
rect 14826 15988 14832 16000
rect 14884 15988 14890 16040
rect 15470 15988 15476 16040
rect 15528 16028 15534 16040
rect 16669 16031 16727 16037
rect 16669 16028 16681 16031
rect 15528 16000 16681 16028
rect 15528 15988 15534 16000
rect 16669 15997 16681 16000
rect 16715 15997 16727 16031
rect 16669 15991 16727 15997
rect 12584 15932 14596 15960
rect 12584 15920 12590 15932
rect 11606 15892 11612 15904
rect 3844 15864 9352 15892
rect 11567 15864 11612 15892
rect 3844 15852 3850 15864
rect 11606 15852 11612 15864
rect 11664 15852 11670 15904
rect 15930 15892 15936 15904
rect 15891 15864 15936 15892
rect 15930 15852 15936 15864
rect 15988 15852 15994 15904
rect 16666 15852 16672 15904
rect 16724 15892 16730 15904
rect 16853 15895 16911 15901
rect 16853 15892 16865 15895
rect 16724 15864 16865 15892
rect 16724 15852 16730 15864
rect 16853 15861 16865 15864
rect 16899 15861 16911 15895
rect 17972 15892 18000 16068
rect 18322 16056 18328 16068
rect 18380 16056 18386 16108
rect 21008 16105 21036 16204
rect 26510 16192 26516 16204
rect 26568 16192 26574 16244
rect 28994 16192 29000 16244
rect 29052 16232 29058 16244
rect 29917 16235 29975 16241
rect 29917 16232 29929 16235
rect 29052 16204 29929 16232
rect 29052 16192 29058 16204
rect 29917 16201 29929 16204
rect 29963 16232 29975 16235
rect 30190 16232 30196 16244
rect 29963 16204 30196 16232
rect 29963 16201 29975 16204
rect 29917 16195 29975 16201
rect 30190 16192 30196 16204
rect 30248 16192 30254 16244
rect 35526 16192 35532 16244
rect 35584 16232 35590 16244
rect 36909 16235 36967 16241
rect 36909 16232 36921 16235
rect 35584 16204 36921 16232
rect 35584 16192 35590 16204
rect 36909 16201 36921 16204
rect 36955 16201 36967 16235
rect 36909 16195 36967 16201
rect 38194 16192 38200 16244
rect 38252 16232 38258 16244
rect 38841 16235 38899 16241
rect 38841 16232 38853 16235
rect 38252 16204 38853 16232
rect 38252 16192 38258 16204
rect 38841 16201 38853 16204
rect 38887 16201 38899 16235
rect 38841 16195 38899 16201
rect 26418 16164 26424 16176
rect 21100 16136 25728 16164
rect 26379 16136 26424 16164
rect 20993 16099 21051 16105
rect 18984 16068 20852 16096
rect 18049 16031 18107 16037
rect 18049 15997 18061 16031
rect 18095 16028 18107 16031
rect 18690 16028 18696 16040
rect 18095 16000 18696 16028
rect 18095 15997 18107 16000
rect 18049 15991 18107 15997
rect 18690 15988 18696 16000
rect 18748 15988 18754 16040
rect 18984 15892 19012 16068
rect 20533 16031 20591 16037
rect 20533 15997 20545 16031
rect 20579 15997 20591 16031
rect 20714 16028 20720 16040
rect 20675 16000 20720 16028
rect 20533 15991 20591 15997
rect 19886 15920 19892 15972
rect 19944 15920 19950 15972
rect 19426 15892 19432 15904
rect 17972 15864 19012 15892
rect 19387 15864 19432 15892
rect 16853 15855 16911 15861
rect 19426 15852 19432 15864
rect 19484 15892 19490 15904
rect 19904 15892 19932 15920
rect 19484 15864 19932 15892
rect 20548 15892 20576 15991
rect 20714 15988 20720 16000
rect 20772 15988 20778 16040
rect 20824 16028 20852 16068
rect 20993 16065 21005 16099
rect 21039 16065 21051 16099
rect 20993 16059 21051 16065
rect 21100 16028 21128 16136
rect 21266 16056 21272 16108
rect 21324 16096 21330 16108
rect 21324 16068 24164 16096
rect 21324 16056 21330 16068
rect 21928 16037 21956 16068
rect 24136 16040 24164 16068
rect 20824 16000 21128 16028
rect 21913 16031 21971 16037
rect 21913 15997 21925 16031
rect 21959 16028 21971 16031
rect 22094 16028 22100 16040
rect 21959 16000 21993 16028
rect 22055 16000 22100 16028
rect 21959 15997 21971 16000
rect 21913 15991 21971 15997
rect 22094 15988 22100 16000
rect 22152 15988 22158 16040
rect 22278 16028 22284 16040
rect 22239 16000 22284 16028
rect 22278 15988 22284 16000
rect 22336 15988 22342 16040
rect 22557 16031 22615 16037
rect 22557 15997 22569 16031
rect 22603 16028 22615 16031
rect 22646 16028 22652 16040
rect 22603 16000 22652 16028
rect 22603 15997 22615 16000
rect 22557 15991 22615 15997
rect 22646 15988 22652 16000
rect 22704 15988 22710 16040
rect 22833 16031 22891 16037
rect 22833 15997 22845 16031
rect 22879 16028 22891 16031
rect 22922 16028 22928 16040
rect 22879 16000 22928 16028
rect 22879 15997 22891 16000
rect 22833 15991 22891 15997
rect 22922 15988 22928 16000
rect 22980 15988 22986 16040
rect 23474 15988 23480 16040
rect 23532 16028 23538 16040
rect 23842 16028 23848 16040
rect 23532 16000 23848 16028
rect 23532 15988 23538 16000
rect 23842 15988 23848 16000
rect 23900 15988 23906 16040
rect 24118 16028 24124 16040
rect 24031 16000 24124 16028
rect 24118 15988 24124 16000
rect 24176 15988 24182 16040
rect 24394 16028 24400 16040
rect 24355 16000 24400 16028
rect 24394 15988 24400 16000
rect 24452 15988 24458 16040
rect 24486 15988 24492 16040
rect 24544 16028 24550 16040
rect 24670 16028 24676 16040
rect 24544 16000 24589 16028
rect 24631 16000 24676 16028
rect 24544 15988 24550 16000
rect 24670 15988 24676 16000
rect 24728 15988 24734 16040
rect 24946 16028 24952 16040
rect 24907 16000 24952 16028
rect 24946 15988 24952 16000
rect 25004 15988 25010 16040
rect 20806 15920 20812 15972
rect 20864 15960 20870 15972
rect 21453 15963 21511 15969
rect 21453 15960 21465 15963
rect 20864 15932 21465 15960
rect 20864 15920 20870 15932
rect 21453 15929 21465 15932
rect 21499 15929 21511 15963
rect 22296 15960 22324 15988
rect 23661 15963 23719 15969
rect 22296 15932 23612 15960
rect 21453 15923 21511 15929
rect 22094 15892 22100 15904
rect 20548 15864 22100 15892
rect 19484 15852 19490 15864
rect 22094 15852 22100 15864
rect 22152 15892 22158 15904
rect 23014 15892 23020 15904
rect 22152 15864 23020 15892
rect 22152 15852 22158 15864
rect 23014 15852 23020 15864
rect 23072 15852 23078 15904
rect 23584 15892 23612 15932
rect 23661 15929 23673 15963
rect 23707 15960 23719 15963
rect 25130 15960 25136 15972
rect 23707 15932 25136 15960
rect 23707 15929 23719 15932
rect 23661 15923 23719 15929
rect 25130 15920 25136 15932
rect 25188 15920 25194 15972
rect 24394 15892 24400 15904
rect 23584 15864 24400 15892
rect 24394 15852 24400 15864
rect 24452 15852 24458 15904
rect 25700 15892 25728 16136
rect 26418 16124 26424 16136
rect 26476 16124 26482 16176
rect 35618 16164 35624 16176
rect 32876 16136 35624 16164
rect 25777 16099 25835 16105
rect 25777 16065 25789 16099
rect 25823 16096 25835 16099
rect 27338 16096 27344 16108
rect 25823 16068 27344 16096
rect 25823 16065 25835 16068
rect 25777 16059 25835 16065
rect 27338 16056 27344 16068
rect 27396 16056 27402 16108
rect 27985 16099 28043 16105
rect 27985 16096 27997 16099
rect 27448 16068 27997 16096
rect 26142 16028 26148 16040
rect 26103 16000 26148 16028
rect 26142 15988 26148 16000
rect 26200 15988 26206 16040
rect 26326 15988 26332 16040
rect 26384 16028 26390 16040
rect 26421 16031 26479 16037
rect 26421 16028 26433 16031
rect 26384 16000 26433 16028
rect 26384 15988 26390 16000
rect 26421 15997 26433 16000
rect 26467 15997 26479 16031
rect 27448 16028 27476 16068
rect 27985 16065 27997 16068
rect 28031 16065 28043 16099
rect 27985 16059 28043 16065
rect 28350 16056 28356 16108
rect 28408 16096 28414 16108
rect 29270 16096 29276 16108
rect 28408 16068 29276 16096
rect 28408 16056 28414 16068
rect 29270 16056 29276 16068
rect 29328 16056 29334 16108
rect 30466 16096 30472 16108
rect 30427 16068 30472 16096
rect 30466 16056 30472 16068
rect 30524 16056 30530 16108
rect 31110 16056 31116 16108
rect 31168 16105 31174 16108
rect 31168 16099 31217 16105
rect 31168 16065 31171 16099
rect 31205 16065 31217 16099
rect 31168 16059 31217 16065
rect 31168 16056 31174 16059
rect 26421 15991 26479 15997
rect 26528 16000 27476 16028
rect 27709 16031 27767 16037
rect 26050 15920 26056 15972
rect 26108 15960 26114 15972
rect 26528 15960 26556 16000
rect 27709 15997 27721 16031
rect 27755 16028 27767 16031
rect 27798 16028 27804 16040
rect 27755 16000 27804 16028
rect 27755 15997 27767 16000
rect 27709 15991 27767 15997
rect 27798 15988 27804 16000
rect 27856 15988 27862 16040
rect 28077 16031 28135 16037
rect 28077 15997 28089 16031
rect 28123 15997 28135 16031
rect 28077 15991 28135 15997
rect 26108 15932 26556 15960
rect 26108 15920 26114 15932
rect 27246 15920 27252 15972
rect 27304 15960 27310 15972
rect 28092 15960 28120 15991
rect 29178 15988 29184 16040
rect 29236 16028 29242 16040
rect 29733 16031 29791 16037
rect 29733 16028 29745 16031
rect 29236 16000 29745 16028
rect 29236 15988 29242 16000
rect 29733 15997 29745 16000
rect 29779 16028 29791 16031
rect 30282 16028 30288 16040
rect 29779 16000 30288 16028
rect 29779 15997 29791 16000
rect 29733 15991 29791 15997
rect 30282 15988 30288 16000
rect 30340 15988 30346 16040
rect 31018 16028 31024 16040
rect 30979 16000 31024 16028
rect 31018 15988 31024 16000
rect 31076 15988 31082 16040
rect 31297 16031 31355 16037
rect 31297 15997 31309 16031
rect 31343 16028 31355 16031
rect 31941 16031 31999 16037
rect 31941 16028 31953 16031
rect 31343 16000 31953 16028
rect 31343 15997 31355 16000
rect 31297 15991 31355 15997
rect 31941 15997 31953 16000
rect 31987 16028 31999 16031
rect 32214 16028 32220 16040
rect 31987 16000 32220 16028
rect 31987 15997 31999 16000
rect 31941 15991 31999 15997
rect 32214 15988 32220 16000
rect 32272 15988 32278 16040
rect 32876 16037 32904 16136
rect 35618 16124 35624 16136
rect 35676 16124 35682 16176
rect 34330 16056 34336 16108
rect 34388 16096 34394 16108
rect 34388 16068 36032 16096
rect 34388 16056 34394 16068
rect 32861 16031 32919 16037
rect 32861 15997 32873 16031
rect 32907 15997 32919 16031
rect 32861 15991 32919 15997
rect 32950 15988 32956 16040
rect 33008 16028 33014 16040
rect 33413 16031 33471 16037
rect 33413 16028 33425 16031
rect 33008 16000 33425 16028
rect 33008 15988 33014 16000
rect 33413 15997 33425 16000
rect 33459 15997 33471 16031
rect 33686 16028 33692 16040
rect 33647 16000 33692 16028
rect 33413 15991 33471 15997
rect 33686 15988 33692 16000
rect 33744 15988 33750 16040
rect 35434 16028 35440 16040
rect 33796 16000 35440 16028
rect 33796 15960 33824 16000
rect 35434 15988 35440 16000
rect 35492 15988 35498 16040
rect 35802 16028 35808 16040
rect 35763 16000 35808 16028
rect 35802 15988 35808 16000
rect 35860 15988 35866 16040
rect 36004 16037 36032 16068
rect 36078 16056 36084 16108
rect 36136 16096 36142 16108
rect 36136 16068 36860 16096
rect 36136 16056 36142 16068
rect 35989 16031 36047 16037
rect 35989 15997 36001 16031
rect 36035 15997 36047 16031
rect 35989 15991 36047 15997
rect 36173 16031 36231 16037
rect 36173 15997 36185 16031
rect 36219 16028 36231 16031
rect 36354 16028 36360 16040
rect 36219 16000 36360 16028
rect 36219 15997 36231 16000
rect 36173 15991 36231 15997
rect 36354 15988 36360 16000
rect 36412 15988 36418 16040
rect 36832 16037 36860 16068
rect 37182 16056 37188 16108
rect 37240 16096 37246 16108
rect 37461 16099 37519 16105
rect 37461 16096 37473 16099
rect 37240 16068 37473 16096
rect 37240 16056 37246 16068
rect 37461 16065 37473 16068
rect 37507 16065 37519 16099
rect 37461 16059 37519 16065
rect 36817 16031 36875 16037
rect 36817 15997 36829 16031
rect 36863 15997 36875 16031
rect 36817 15991 36875 15997
rect 37737 16031 37795 16037
rect 37737 15997 37749 16031
rect 37783 16028 37795 16031
rect 38746 16028 38752 16040
rect 37783 16000 38752 16028
rect 37783 15997 37795 16000
rect 37737 15991 37795 15997
rect 38746 15988 38752 16000
rect 38804 15988 38810 16040
rect 27304 15932 28120 15960
rect 28368 15932 33824 15960
rect 35345 15963 35403 15969
rect 27304 15920 27310 15932
rect 28368 15892 28396 15932
rect 35345 15929 35357 15963
rect 35391 15960 35403 15963
rect 36538 15960 36544 15972
rect 35391 15932 36544 15960
rect 35391 15929 35403 15932
rect 35345 15923 35403 15929
rect 36538 15920 36544 15932
rect 36596 15920 36602 15972
rect 25700 15864 28396 15892
rect 32030 15852 32036 15904
rect 32088 15892 32094 15904
rect 32125 15895 32183 15901
rect 32125 15892 32137 15895
rect 32088 15864 32137 15892
rect 32088 15852 32094 15864
rect 32125 15861 32137 15864
rect 32171 15861 32183 15895
rect 32125 15855 32183 15861
rect 32953 15895 33011 15901
rect 32953 15861 32965 15895
rect 32999 15892 33011 15895
rect 33778 15892 33784 15904
rect 32999 15864 33784 15892
rect 32999 15861 33011 15864
rect 32953 15855 33011 15861
rect 33778 15852 33784 15864
rect 33836 15852 33842 15904
rect 1104 15802 39836 15824
rect 1104 15750 19606 15802
rect 19658 15750 19670 15802
rect 19722 15750 19734 15802
rect 19786 15750 19798 15802
rect 19850 15750 39836 15802
rect 1104 15728 39836 15750
rect 3694 15648 3700 15700
rect 3752 15688 3758 15700
rect 5445 15691 5503 15697
rect 5445 15688 5457 15691
rect 3752 15660 5457 15688
rect 3752 15648 3758 15660
rect 5445 15657 5457 15660
rect 5491 15657 5503 15691
rect 5445 15651 5503 15657
rect 9674 15648 9680 15700
rect 9732 15688 9738 15700
rect 9732 15660 10916 15688
rect 9732 15648 9738 15660
rect 1670 15580 1676 15632
rect 1728 15620 1734 15632
rect 2961 15623 3019 15629
rect 2961 15620 2973 15623
rect 1728 15592 2973 15620
rect 1728 15580 1734 15592
rect 2961 15589 2973 15592
rect 3007 15589 3019 15623
rect 2961 15583 3019 15589
rect 10888 15620 10916 15660
rect 12618 15648 12624 15700
rect 12676 15688 12682 15700
rect 13630 15688 13636 15700
rect 12676 15660 13636 15688
rect 12676 15648 12682 15660
rect 13630 15648 13636 15660
rect 13688 15688 13694 15700
rect 14093 15691 14151 15697
rect 14093 15688 14105 15691
rect 13688 15660 14105 15688
rect 13688 15648 13694 15660
rect 14093 15657 14105 15660
rect 14139 15657 14151 15691
rect 14093 15651 14151 15657
rect 14458 15648 14464 15700
rect 14516 15688 14522 15700
rect 20806 15688 20812 15700
rect 14516 15660 20812 15688
rect 14516 15648 14522 15660
rect 20806 15648 20812 15660
rect 20864 15648 20870 15700
rect 21085 15691 21143 15697
rect 21085 15657 21097 15691
rect 21131 15688 21143 15691
rect 25222 15688 25228 15700
rect 21131 15660 25228 15688
rect 21131 15657 21143 15660
rect 21085 15651 21143 15657
rect 25222 15648 25228 15660
rect 25280 15648 25286 15700
rect 26602 15688 26608 15700
rect 26563 15660 26608 15688
rect 26602 15648 26608 15660
rect 26660 15648 26666 15700
rect 29270 15688 29276 15700
rect 29231 15660 29276 15688
rect 29270 15648 29276 15660
rect 29328 15648 29334 15700
rect 29638 15648 29644 15700
rect 29696 15688 29702 15700
rect 29914 15688 29920 15700
rect 29696 15660 29920 15688
rect 29696 15648 29702 15660
rect 29914 15648 29920 15660
rect 29972 15648 29978 15700
rect 30006 15648 30012 15700
rect 30064 15688 30070 15700
rect 31113 15691 31171 15697
rect 31113 15688 31125 15691
rect 30064 15660 31125 15688
rect 30064 15648 30070 15660
rect 31113 15657 31125 15660
rect 31159 15657 31171 15691
rect 31113 15651 31171 15657
rect 32306 15648 32312 15700
rect 32364 15688 32370 15700
rect 37826 15688 37832 15700
rect 32364 15660 36400 15688
rect 37787 15660 37832 15688
rect 32364 15648 32370 15660
rect 11606 15620 11612 15632
rect 10888 15592 11612 15620
rect 2501 15555 2559 15561
rect 2501 15521 2513 15555
rect 2547 15552 2559 15555
rect 2774 15552 2780 15564
rect 2547 15524 2780 15552
rect 2547 15521 2559 15524
rect 2501 15515 2559 15521
rect 2774 15512 2780 15524
rect 2832 15512 2838 15564
rect 3878 15552 3884 15564
rect 3839 15524 3884 15552
rect 3878 15512 3884 15524
rect 3936 15512 3942 15564
rect 6457 15555 6515 15561
rect 6457 15521 6469 15555
rect 6503 15552 6515 15555
rect 6503 15524 8064 15552
rect 6503 15521 6515 15524
rect 6457 15515 6515 15521
rect 2409 15487 2467 15493
rect 2409 15453 2421 15487
rect 2455 15484 2467 15487
rect 2682 15484 2688 15496
rect 2455 15456 2688 15484
rect 2455 15453 2467 15456
rect 2409 15447 2467 15453
rect 2682 15444 2688 15456
rect 2740 15484 2746 15496
rect 3786 15484 3792 15496
rect 2740 15456 3792 15484
rect 2740 15444 2746 15456
rect 3786 15444 3792 15456
rect 3844 15444 3850 15496
rect 4062 15484 4068 15496
rect 4023 15456 4068 15484
rect 4062 15444 4068 15456
rect 4120 15444 4126 15496
rect 4341 15487 4399 15493
rect 4341 15453 4353 15487
rect 4387 15484 4399 15487
rect 4798 15484 4804 15496
rect 4387 15456 4804 15484
rect 4387 15453 4399 15456
rect 4341 15447 4399 15453
rect 4798 15444 4804 15456
rect 4856 15444 4862 15496
rect 6733 15487 6791 15493
rect 6733 15453 6745 15487
rect 6779 15484 6791 15487
rect 6914 15484 6920 15496
rect 6779 15456 6920 15484
rect 6779 15453 6791 15456
rect 6733 15447 6791 15453
rect 6914 15444 6920 15456
rect 6972 15444 6978 15496
rect 3510 15376 3516 15428
rect 3568 15416 3574 15428
rect 3697 15419 3755 15425
rect 3697 15416 3709 15419
rect 3568 15388 3709 15416
rect 3568 15376 3574 15388
rect 3697 15385 3709 15388
rect 3743 15385 3755 15419
rect 8036 15416 8064 15524
rect 8478 15512 8484 15564
rect 8536 15552 8542 15564
rect 8573 15555 8631 15561
rect 8573 15552 8585 15555
rect 8536 15524 8585 15552
rect 8536 15512 8542 15524
rect 8573 15521 8585 15524
rect 8619 15521 8631 15555
rect 8573 15515 8631 15521
rect 9677 15555 9735 15561
rect 9677 15521 9689 15555
rect 9723 15521 9735 15555
rect 10410 15552 10416 15564
rect 10323 15524 10416 15552
rect 9677 15515 9735 15521
rect 8113 15487 8171 15493
rect 8113 15453 8125 15487
rect 8159 15484 8171 15487
rect 8846 15484 8852 15496
rect 8159 15456 8852 15484
rect 8159 15453 8171 15456
rect 8113 15447 8171 15453
rect 8846 15444 8852 15456
rect 8904 15484 8910 15496
rect 9692 15484 9720 15515
rect 10410 15512 10416 15524
rect 10468 15552 10474 15564
rect 10888 15561 10916 15592
rect 11606 15580 11612 15592
rect 11664 15580 11670 15632
rect 12802 15620 12808 15632
rect 12268 15592 12808 15620
rect 10873 15555 10931 15561
rect 10468 15524 10640 15552
rect 10468 15512 10474 15524
rect 8904 15456 9720 15484
rect 8904 15444 8910 15456
rect 9766 15444 9772 15496
rect 9824 15444 9830 15496
rect 10502 15484 10508 15496
rect 10463 15456 10508 15484
rect 10502 15444 10508 15456
rect 10560 15444 10566 15496
rect 10612 15484 10640 15524
rect 10873 15521 10885 15555
rect 10919 15521 10931 15555
rect 11054 15552 11060 15564
rect 11015 15524 11060 15552
rect 10873 15515 10931 15521
rect 11054 15512 11060 15524
rect 11112 15512 11118 15564
rect 11698 15552 11704 15564
rect 11659 15524 11704 15552
rect 11698 15512 11704 15524
rect 11756 15512 11762 15564
rect 12268 15561 12296 15592
rect 12802 15580 12808 15592
rect 12860 15580 12866 15632
rect 17586 15620 17592 15632
rect 13648 15592 17172 15620
rect 12253 15555 12311 15561
rect 12253 15521 12265 15555
rect 12299 15521 12311 15555
rect 12253 15515 12311 15521
rect 12526 15512 12532 15564
rect 12584 15552 12590 15564
rect 12713 15555 12771 15561
rect 12713 15552 12725 15555
rect 12584 15524 12725 15552
rect 12584 15512 12590 15524
rect 12713 15521 12725 15524
rect 12759 15521 12771 15555
rect 12986 15552 12992 15564
rect 12947 15524 12992 15552
rect 12713 15515 12771 15521
rect 12986 15512 12992 15524
rect 13044 15512 13050 15564
rect 13078 15512 13084 15564
rect 13136 15552 13142 15564
rect 13648 15552 13676 15592
rect 13136 15524 13676 15552
rect 16025 15555 16083 15561
rect 13136 15512 13142 15524
rect 16025 15521 16037 15555
rect 16071 15521 16083 15555
rect 16390 15552 16396 15564
rect 16351 15524 16396 15552
rect 16025 15515 16083 15521
rect 14458 15484 14464 15496
rect 10612 15456 14464 15484
rect 14458 15444 14464 15456
rect 14516 15444 14522 15496
rect 15657 15487 15715 15493
rect 15657 15453 15669 15487
rect 15703 15453 15715 15487
rect 16040 15484 16068 15515
rect 16390 15512 16396 15524
rect 16448 15512 16454 15564
rect 16482 15512 16488 15564
rect 16540 15552 16546 15564
rect 16577 15555 16635 15561
rect 16577 15552 16589 15555
rect 16540 15524 16589 15552
rect 16540 15512 16546 15524
rect 16577 15521 16589 15524
rect 16623 15521 16635 15555
rect 16577 15515 16635 15521
rect 16666 15484 16672 15496
rect 16040 15456 16672 15484
rect 15657 15447 15715 15453
rect 9784 15416 9812 15444
rect 10226 15416 10232 15428
rect 8036 15388 10232 15416
rect 3697 15379 3755 15385
rect 10226 15376 10232 15388
rect 10284 15376 10290 15428
rect 3234 15308 3240 15360
rect 3292 15348 3298 15360
rect 8757 15351 8815 15357
rect 8757 15348 8769 15351
rect 3292 15320 8769 15348
rect 3292 15308 3298 15320
rect 8757 15317 8769 15320
rect 8803 15317 8815 15351
rect 8757 15311 8815 15317
rect 9030 15308 9036 15360
rect 9088 15348 9094 15360
rect 9769 15351 9827 15357
rect 9769 15348 9781 15351
rect 9088 15320 9781 15348
rect 9088 15308 9094 15320
rect 9769 15317 9781 15320
rect 9815 15317 9827 15351
rect 9769 15311 9827 15317
rect 10134 15308 10140 15360
rect 10192 15348 10198 15360
rect 15286 15348 15292 15360
rect 10192 15320 15292 15348
rect 10192 15308 10198 15320
rect 15286 15308 15292 15320
rect 15344 15308 15350 15360
rect 15672 15348 15700 15447
rect 16666 15444 16672 15456
rect 16724 15444 16730 15496
rect 16942 15348 16948 15360
rect 15672 15320 16948 15348
rect 16942 15308 16948 15320
rect 17000 15308 17006 15360
rect 17144 15348 17172 15592
rect 17328 15592 17592 15620
rect 17328 15561 17356 15592
rect 17586 15580 17592 15592
rect 17644 15580 17650 15632
rect 18506 15620 18512 15632
rect 17788 15592 18512 15620
rect 17313 15555 17371 15561
rect 17313 15521 17325 15555
rect 17359 15521 17371 15555
rect 17313 15515 17371 15521
rect 17497 15555 17555 15561
rect 17497 15521 17509 15555
rect 17543 15552 17555 15555
rect 17788 15552 17816 15592
rect 18506 15580 18512 15592
rect 18564 15580 18570 15632
rect 22186 15620 22192 15632
rect 21008 15592 22192 15620
rect 17954 15552 17960 15564
rect 17543 15524 17816 15552
rect 17915 15524 17960 15552
rect 17543 15521 17555 15524
rect 17497 15515 17555 15521
rect 17954 15512 17960 15524
rect 18012 15512 18018 15564
rect 18690 15552 18696 15564
rect 18651 15524 18696 15552
rect 18690 15512 18696 15524
rect 18748 15512 18754 15564
rect 20530 15552 20536 15564
rect 18800 15524 20536 15552
rect 17678 15484 17684 15496
rect 17639 15456 17684 15484
rect 17678 15444 17684 15456
rect 17736 15444 17742 15496
rect 18138 15444 18144 15496
rect 18196 15484 18202 15496
rect 18800 15484 18828 15524
rect 20530 15512 20536 15524
rect 20588 15512 20594 15564
rect 21008 15561 21036 15592
rect 22186 15580 22192 15592
rect 22244 15580 22250 15632
rect 24394 15580 24400 15632
rect 24452 15620 24458 15632
rect 26620 15620 26648 15648
rect 29362 15620 29368 15632
rect 24452 15592 24532 15620
rect 26620 15592 29368 15620
rect 24452 15580 24458 15592
rect 20993 15555 21051 15561
rect 20993 15521 21005 15555
rect 21039 15521 21051 15555
rect 20993 15515 21051 15521
rect 22094 15512 22100 15564
rect 22152 15552 22158 15564
rect 22278 15552 22284 15564
rect 22152 15524 22197 15552
rect 22239 15524 22284 15552
rect 22152 15512 22158 15524
rect 22278 15512 22284 15524
rect 22336 15512 22342 15564
rect 22554 15552 22560 15564
rect 22515 15524 22560 15552
rect 22554 15512 22560 15524
rect 22612 15512 22618 15564
rect 22646 15512 22652 15564
rect 22704 15552 22710 15564
rect 23017 15555 23075 15561
rect 22704 15524 22749 15552
rect 22704 15512 22710 15524
rect 23017 15521 23029 15555
rect 23063 15552 23075 15555
rect 23290 15552 23296 15564
rect 23063 15524 23296 15552
rect 23063 15521 23075 15524
rect 23017 15515 23075 15521
rect 23290 15512 23296 15524
rect 23348 15512 23354 15564
rect 24118 15552 24124 15564
rect 24079 15524 24124 15552
rect 24118 15512 24124 15524
rect 24176 15512 24182 15564
rect 24504 15561 24532 15592
rect 24213 15555 24271 15561
rect 24213 15521 24225 15555
rect 24259 15521 24271 15555
rect 24213 15515 24271 15521
rect 24489 15555 24547 15561
rect 24489 15521 24501 15555
rect 24535 15521 24547 15555
rect 24489 15515 24547 15521
rect 24581 15555 24639 15561
rect 24581 15521 24593 15555
rect 24627 15521 24639 15555
rect 24946 15552 24952 15564
rect 24907 15524 24952 15552
rect 24581 15515 24639 15521
rect 18966 15484 18972 15496
rect 18196 15456 18828 15484
rect 18927 15456 18972 15484
rect 18196 15444 18202 15456
rect 18966 15444 18972 15456
rect 19024 15444 19030 15496
rect 20806 15444 20812 15496
rect 20864 15484 20870 15496
rect 21637 15487 21695 15493
rect 21637 15484 21649 15487
rect 20864 15456 21649 15484
rect 20864 15444 20870 15456
rect 21637 15453 21649 15456
rect 21683 15453 21695 15487
rect 21637 15447 21695 15453
rect 23569 15487 23627 15493
rect 23569 15453 23581 15487
rect 23615 15453 23627 15487
rect 23569 15447 23627 15453
rect 20714 15416 20720 15428
rect 19904 15388 20720 15416
rect 19904 15348 19932 15388
rect 20714 15376 20720 15388
rect 20772 15376 20778 15428
rect 23584 15416 23612 15447
rect 24026 15444 24032 15496
rect 24084 15484 24090 15496
rect 24228 15484 24256 15515
rect 24084 15456 24256 15484
rect 24084 15444 24090 15456
rect 24394 15444 24400 15496
rect 24452 15484 24458 15496
rect 24596 15484 24624 15515
rect 24946 15512 24952 15524
rect 25004 15552 25010 15564
rect 25501 15555 25559 15561
rect 25501 15552 25513 15555
rect 25004 15524 25513 15552
rect 25004 15512 25010 15524
rect 25501 15521 25513 15524
rect 25547 15521 25559 15555
rect 25501 15515 25559 15521
rect 26513 15555 26571 15561
rect 26513 15521 26525 15555
rect 26559 15552 26571 15555
rect 26878 15552 26884 15564
rect 26559 15524 26884 15552
rect 26559 15521 26571 15524
rect 26513 15515 26571 15521
rect 26878 15512 26884 15524
rect 26936 15512 26942 15564
rect 27154 15552 27160 15564
rect 27115 15524 27160 15552
rect 27154 15512 27160 15524
rect 27212 15512 27218 15564
rect 27890 15552 27896 15564
rect 27851 15524 27896 15552
rect 27890 15512 27896 15524
rect 27948 15512 27954 15564
rect 29012 15561 29040 15592
rect 29362 15580 29368 15592
rect 29420 15580 29426 15632
rect 29730 15620 29736 15632
rect 29656 15592 29736 15620
rect 29656 15561 29684 15592
rect 29730 15580 29736 15592
rect 29788 15580 29794 15632
rect 33502 15620 33508 15632
rect 29840 15592 30972 15620
rect 29840 15564 29868 15592
rect 28997 15555 29055 15561
rect 28997 15521 29009 15555
rect 29043 15521 29055 15555
rect 28997 15515 29055 15521
rect 29641 15555 29699 15561
rect 29641 15521 29653 15555
rect 29687 15521 29699 15555
rect 29822 15552 29828 15564
rect 29783 15524 29828 15552
rect 29641 15515 29699 15521
rect 29822 15512 29828 15524
rect 29880 15512 29886 15564
rect 30190 15552 30196 15564
rect 30151 15524 30196 15552
rect 30190 15512 30196 15524
rect 30248 15512 30254 15564
rect 30944 15561 30972 15592
rect 32600 15592 33508 15620
rect 32600 15561 32628 15592
rect 33502 15580 33508 15592
rect 33560 15580 33566 15632
rect 36262 15620 36268 15632
rect 35820 15592 36268 15620
rect 30929 15555 30987 15561
rect 30929 15521 30941 15555
rect 30975 15521 30987 15555
rect 30929 15515 30987 15521
rect 32585 15555 32643 15561
rect 32585 15521 32597 15555
rect 32631 15521 32643 15555
rect 32585 15515 32643 15521
rect 32677 15555 32735 15561
rect 32677 15521 32689 15555
rect 32723 15552 32735 15555
rect 32950 15552 32956 15564
rect 32723 15524 32956 15552
rect 32723 15521 32735 15524
rect 32677 15515 32735 15521
rect 32950 15512 32956 15524
rect 33008 15512 33014 15564
rect 33045 15555 33103 15561
rect 33045 15521 33057 15555
rect 33091 15552 33103 15555
rect 33134 15552 33140 15564
rect 33091 15524 33140 15552
rect 33091 15521 33103 15524
rect 33045 15515 33103 15521
rect 33134 15512 33140 15524
rect 33192 15512 33198 15564
rect 33778 15552 33784 15564
rect 33739 15524 33784 15552
rect 33778 15512 33784 15524
rect 33836 15512 33842 15564
rect 35820 15561 35848 15592
rect 36262 15580 36268 15592
rect 36320 15580 36326 15632
rect 36372 15620 36400 15660
rect 37826 15648 37832 15660
rect 37884 15648 37890 15700
rect 39022 15688 39028 15700
rect 38983 15660 39028 15688
rect 39022 15648 39028 15660
rect 39080 15648 39086 15700
rect 36372 15592 37780 15620
rect 35805 15555 35863 15561
rect 35805 15521 35817 15555
rect 35851 15521 35863 15555
rect 36170 15552 36176 15564
rect 36131 15524 36176 15552
rect 35805 15515 35863 15521
rect 36170 15512 36176 15524
rect 36228 15512 36234 15564
rect 36446 15552 36452 15564
rect 36407 15524 36452 15552
rect 36446 15512 36452 15524
rect 36504 15512 36510 15564
rect 36538 15512 36544 15564
rect 36596 15552 36602 15564
rect 37752 15561 37780 15592
rect 36817 15555 36875 15561
rect 36817 15552 36829 15555
rect 36596 15524 36829 15552
rect 36596 15512 36602 15524
rect 36817 15521 36829 15524
rect 36863 15521 36875 15555
rect 36817 15515 36875 15521
rect 37737 15555 37795 15561
rect 37737 15521 37749 15555
rect 37783 15521 37795 15555
rect 37737 15515 37795 15521
rect 38197 15555 38255 15561
rect 38197 15521 38209 15555
rect 38243 15521 38255 15555
rect 38930 15552 38936 15564
rect 38891 15524 38936 15552
rect 38197 15515 38255 15521
rect 24452 15456 24624 15484
rect 24452 15444 24458 15456
rect 26142 15444 26148 15496
rect 26200 15484 26206 15496
rect 27982 15484 27988 15496
rect 26200 15456 27844 15484
rect 27943 15456 27988 15484
rect 26200 15444 26206 15456
rect 27816 15428 27844 15456
rect 27982 15444 27988 15456
rect 28040 15444 28046 15496
rect 32122 15444 32128 15496
rect 32180 15484 32186 15496
rect 33505 15487 33563 15493
rect 33505 15484 33517 15487
rect 32180 15456 33517 15484
rect 32180 15444 32186 15456
rect 33505 15453 33517 15456
rect 33551 15484 33563 15487
rect 34238 15484 34244 15496
rect 33551 15456 34244 15484
rect 33551 15453 33563 15456
rect 33505 15447 33563 15453
rect 34238 15444 34244 15456
rect 34296 15484 34302 15496
rect 34422 15484 34428 15496
rect 34296 15456 34428 15484
rect 34296 15444 34302 15456
rect 34422 15444 34428 15456
rect 34480 15444 34486 15496
rect 36081 15487 36139 15493
rect 36081 15453 36093 15487
rect 36127 15484 36139 15487
rect 38212 15484 38240 15515
rect 38930 15512 38936 15524
rect 38988 15512 38994 15564
rect 36127 15456 38240 15484
rect 36127 15453 36139 15456
rect 36081 15447 36139 15453
rect 24670 15416 24676 15428
rect 23584 15388 24676 15416
rect 24670 15376 24676 15388
rect 24728 15376 24734 15428
rect 27430 15416 27436 15428
rect 27391 15388 27436 15416
rect 27430 15376 27436 15388
rect 27488 15376 27494 15428
rect 27798 15376 27804 15428
rect 27856 15416 27862 15428
rect 30926 15416 30932 15428
rect 27856 15388 30932 15416
rect 27856 15376 27862 15388
rect 30926 15376 30932 15388
rect 30984 15416 30990 15428
rect 32030 15416 32036 15428
rect 30984 15388 32036 15416
rect 30984 15376 30990 15388
rect 32030 15376 32036 15388
rect 32088 15376 32094 15428
rect 17144 15320 19932 15348
rect 20257 15351 20315 15357
rect 20257 15317 20269 15351
rect 20303 15348 20315 15351
rect 20530 15348 20536 15360
rect 20303 15320 20536 15348
rect 20303 15317 20315 15320
rect 20257 15311 20315 15317
rect 20530 15308 20536 15320
rect 20588 15308 20594 15360
rect 22922 15308 22928 15360
rect 22980 15348 22986 15360
rect 23382 15348 23388 15360
rect 22980 15320 23388 15348
rect 22980 15308 22986 15320
rect 23382 15308 23388 15320
rect 23440 15348 23446 15360
rect 24486 15348 24492 15360
rect 23440 15320 24492 15348
rect 23440 15308 23446 15320
rect 24486 15308 24492 15320
rect 24544 15308 24550 15360
rect 25682 15348 25688 15360
rect 25595 15320 25688 15348
rect 25682 15308 25688 15320
rect 25740 15348 25746 15360
rect 30558 15348 30564 15360
rect 25740 15320 30564 15348
rect 25740 15308 25746 15320
rect 30558 15308 30564 15320
rect 30616 15308 30622 15360
rect 35069 15351 35127 15357
rect 35069 15317 35081 15351
rect 35115 15348 35127 15351
rect 35342 15348 35348 15360
rect 35115 15320 35348 15348
rect 35115 15317 35127 15320
rect 35069 15311 35127 15317
rect 35342 15308 35348 15320
rect 35400 15308 35406 15360
rect 1104 15258 39836 15280
rect 1104 15206 4246 15258
rect 4298 15206 4310 15258
rect 4362 15206 4374 15258
rect 4426 15206 4438 15258
rect 4490 15206 34966 15258
rect 35018 15206 35030 15258
rect 35082 15206 35094 15258
rect 35146 15206 35158 15258
rect 35210 15206 39836 15258
rect 1104 15184 39836 15206
rect 2774 15104 2780 15156
rect 2832 15144 2838 15156
rect 5629 15147 5687 15153
rect 2832 15116 2877 15144
rect 2832 15104 2838 15116
rect 5629 15113 5641 15147
rect 5675 15144 5687 15147
rect 7006 15144 7012 15156
rect 5675 15116 7012 15144
rect 5675 15113 5687 15116
rect 5629 15107 5687 15113
rect 7006 15104 7012 15116
rect 7064 15104 7070 15156
rect 9214 15104 9220 15156
rect 9272 15144 9278 15156
rect 11054 15144 11060 15156
rect 9272 15116 11060 15144
rect 9272 15104 9278 15116
rect 11054 15104 11060 15116
rect 11112 15144 11118 15156
rect 11790 15144 11796 15156
rect 11112 15116 11796 15144
rect 11112 15104 11118 15116
rect 11790 15104 11796 15116
rect 11848 15104 11854 15156
rect 16022 15144 16028 15156
rect 13648 15116 16028 15144
rect 6914 15036 6920 15088
rect 6972 15076 6978 15088
rect 8481 15079 8539 15085
rect 8481 15076 8493 15079
rect 6972 15048 8493 15076
rect 6972 15036 6978 15048
rect 8481 15045 8493 15048
rect 8527 15045 8539 15079
rect 11698 15076 11704 15088
rect 8481 15039 8539 15045
rect 9600 15048 11704 15076
rect 1673 15011 1731 15017
rect 1673 14977 1685 15011
rect 1719 15008 1731 15011
rect 7561 15011 7619 15017
rect 7561 15008 7573 15011
rect 1719 14980 7573 15008
rect 1719 14977 1731 14980
rect 1673 14971 1731 14977
rect 7561 14977 7573 14980
rect 7607 14977 7619 15011
rect 9490 15008 9496 15020
rect 7561 14971 7619 14977
rect 8496 14980 9496 15008
rect 1397 14943 1455 14949
rect 1397 14909 1409 14943
rect 1443 14940 1455 14943
rect 1486 14940 1492 14952
rect 1443 14912 1492 14940
rect 1443 14909 1455 14912
rect 1397 14903 1455 14909
rect 1486 14900 1492 14912
rect 1544 14940 1550 14952
rect 4062 14940 4068 14952
rect 1544 14912 4068 14940
rect 1544 14900 1550 14912
rect 4062 14900 4068 14912
rect 4120 14900 4126 14952
rect 4341 14943 4399 14949
rect 4341 14909 4353 14943
rect 4387 14940 4399 14943
rect 4614 14940 4620 14952
rect 4387 14912 4620 14940
rect 4387 14909 4399 14912
rect 4341 14903 4399 14909
rect 4614 14900 4620 14912
rect 4672 14900 4678 14952
rect 7285 14943 7343 14949
rect 7285 14909 7297 14943
rect 7331 14940 7343 14943
rect 7469 14943 7527 14949
rect 7331 14912 7420 14940
rect 7331 14909 7343 14912
rect 7285 14903 7343 14909
rect 7098 14764 7104 14816
rect 7156 14804 7162 14816
rect 7392 14804 7420 14912
rect 7469 14909 7481 14943
rect 7515 14940 7527 14943
rect 8496 14940 8524 14980
rect 9490 14968 9496 14980
rect 9548 14968 9554 15020
rect 9600 14952 9628 15048
rect 11698 15036 11704 15048
rect 11756 15036 11762 15088
rect 13354 15076 13360 15088
rect 13315 15048 13360 15076
rect 13354 15036 13360 15048
rect 13412 15036 13418 15088
rect 13648 15008 13676 15116
rect 16022 15104 16028 15116
rect 16080 15104 16086 15156
rect 19426 15144 19432 15156
rect 17144 15116 19432 15144
rect 15654 15036 15660 15088
rect 15712 15076 15718 15088
rect 17144 15076 17172 15116
rect 19426 15104 19432 15116
rect 19484 15104 19490 15156
rect 20438 15104 20444 15156
rect 20496 15144 20502 15156
rect 21269 15147 21327 15153
rect 21269 15144 21281 15147
rect 20496 15116 21281 15144
rect 20496 15104 20502 15116
rect 21269 15113 21281 15116
rect 21315 15113 21327 15147
rect 38746 15144 38752 15156
rect 21269 15107 21327 15113
rect 22848 15116 28580 15144
rect 38707 15116 38752 15144
rect 15712 15048 17172 15076
rect 15712 15036 15718 15048
rect 17218 15036 17224 15088
rect 17276 15076 17282 15088
rect 17862 15076 17868 15088
rect 17276 15048 17868 15076
rect 17276 15036 17282 15048
rect 17862 15036 17868 15048
rect 17920 15076 17926 15088
rect 17920 15048 19104 15076
rect 17920 15036 17926 15048
rect 13814 15008 13820 15020
rect 13556 14980 13676 15008
rect 13775 14980 13820 15008
rect 7515 14912 8524 14940
rect 8573 14943 8631 14949
rect 7515 14909 7527 14912
rect 7469 14903 7527 14909
rect 8573 14909 8585 14943
rect 8619 14909 8631 14943
rect 9030 14940 9036 14952
rect 8991 14912 9036 14940
rect 8573 14903 8631 14909
rect 8110 14804 8116 14816
rect 7156 14776 8116 14804
rect 7156 14764 7162 14776
rect 8110 14764 8116 14776
rect 8168 14764 8174 14816
rect 8202 14764 8208 14816
rect 8260 14804 8266 14816
rect 8588 14804 8616 14903
rect 9030 14900 9036 14912
rect 9088 14900 9094 14952
rect 9214 14940 9220 14952
rect 9175 14912 9220 14940
rect 9214 14900 9220 14912
rect 9272 14900 9278 14952
rect 9582 14940 9588 14952
rect 9543 14912 9588 14940
rect 9582 14900 9588 14912
rect 9640 14900 9646 14952
rect 10321 14943 10379 14949
rect 10321 14909 10333 14943
rect 10367 14940 10379 14943
rect 10594 14940 10600 14952
rect 10367 14912 10600 14940
rect 10367 14909 10379 14912
rect 10321 14903 10379 14909
rect 10594 14900 10600 14912
rect 10652 14900 10658 14952
rect 10778 14940 10784 14952
rect 10739 14912 10784 14940
rect 10778 14900 10784 14912
rect 10836 14900 10842 14952
rect 11422 14900 11428 14952
rect 11480 14940 11486 14952
rect 11517 14943 11575 14949
rect 11517 14940 11529 14943
rect 11480 14912 11529 14940
rect 11480 14900 11486 14912
rect 11517 14909 11529 14912
rect 11563 14909 11575 14943
rect 11517 14903 11575 14909
rect 12437 14943 12495 14949
rect 12437 14909 12449 14943
rect 12483 14940 12495 14943
rect 12618 14940 12624 14952
rect 12483 14912 12624 14940
rect 12483 14909 12495 14912
rect 12437 14903 12495 14909
rect 12618 14900 12624 14912
rect 12676 14900 12682 14952
rect 13556 14949 13584 14980
rect 13814 14968 13820 14980
rect 13872 14968 13878 15020
rect 15286 15008 15292 15020
rect 14292 14980 15292 15008
rect 13541 14943 13599 14949
rect 13541 14909 13553 14943
rect 13587 14909 13599 14943
rect 13541 14903 13599 14909
rect 13630 14900 13636 14952
rect 13688 14940 13694 14952
rect 14292 14949 14320 14980
rect 15286 14968 15292 14980
rect 15344 15008 15350 15020
rect 16390 15008 16396 15020
rect 15344 14980 16252 15008
rect 16351 14980 16396 15008
rect 15344 14968 15350 14980
rect 14277 14943 14335 14949
rect 13688 14912 13733 14940
rect 13688 14900 13694 14912
rect 14277 14909 14289 14943
rect 14323 14909 14335 14943
rect 14277 14903 14335 14909
rect 14645 14943 14703 14949
rect 14645 14909 14657 14943
rect 14691 14940 14703 14943
rect 15378 14940 15384 14952
rect 14691 14912 15384 14940
rect 14691 14909 14703 14912
rect 14645 14903 14703 14909
rect 15378 14900 15384 14912
rect 15436 14900 15442 14952
rect 15562 14900 15568 14952
rect 15620 14940 15626 14952
rect 15841 14943 15899 14949
rect 15841 14940 15853 14943
rect 15620 14912 15853 14940
rect 15620 14900 15626 14912
rect 15841 14909 15853 14912
rect 15887 14909 15899 14943
rect 16224 14940 16252 14980
rect 16390 14968 16396 14980
rect 16448 14968 16454 15020
rect 18506 15008 18512 15020
rect 16500 14980 18512 15008
rect 16500 14949 16528 14980
rect 18506 14968 18512 14980
rect 18564 14968 18570 15020
rect 18966 15008 18972 15020
rect 18927 14980 18972 15008
rect 18966 14968 18972 14980
rect 19024 14968 19030 15020
rect 19076 15008 19104 15048
rect 19334 15036 19340 15088
rect 19392 15076 19398 15088
rect 22738 15076 22744 15088
rect 19392 15048 22744 15076
rect 19392 15036 19398 15048
rect 22738 15036 22744 15048
rect 22796 15036 22802 15088
rect 22848 15008 22876 15116
rect 23014 15036 23020 15088
rect 23072 15076 23078 15088
rect 24946 15076 24952 15088
rect 23072 15048 24952 15076
rect 23072 15036 23078 15048
rect 19076 14980 22876 15008
rect 16485 14943 16543 14949
rect 16485 14940 16497 14943
rect 16224 14912 16497 14940
rect 15841 14903 15899 14909
rect 16485 14909 16497 14912
rect 16531 14909 16543 14943
rect 16485 14903 16543 14909
rect 16853 14943 16911 14949
rect 16853 14909 16865 14943
rect 16899 14940 16911 14943
rect 17954 14940 17960 14952
rect 16899 14912 17960 14940
rect 16899 14909 16911 14912
rect 16853 14903 16911 14909
rect 17954 14900 17960 14912
rect 18012 14900 18018 14952
rect 18049 14943 18107 14949
rect 18049 14909 18061 14943
rect 18095 14909 18107 14943
rect 18049 14903 18107 14909
rect 18877 14943 18935 14949
rect 18877 14909 18889 14943
rect 18923 14909 18935 14943
rect 19334 14940 19340 14952
rect 19295 14912 19340 14940
rect 18877 14903 18935 14909
rect 8938 14832 8944 14884
rect 8996 14872 9002 14884
rect 17678 14872 17684 14884
rect 8996 14844 17684 14872
rect 8996 14832 9002 14844
rect 17678 14832 17684 14844
rect 17736 14832 17742 14884
rect 18064 14872 18092 14903
rect 17880 14844 18092 14872
rect 10410 14804 10416 14816
rect 8260 14776 10416 14804
rect 8260 14764 8266 14776
rect 10410 14764 10416 14776
rect 10468 14764 10474 14816
rect 10962 14804 10968 14816
rect 10923 14776 10968 14804
rect 10962 14764 10968 14776
rect 11020 14764 11026 14816
rect 11698 14804 11704 14816
rect 11659 14776 11704 14804
rect 11698 14764 11704 14776
rect 11756 14764 11762 14816
rect 11790 14764 11796 14816
rect 11848 14804 11854 14816
rect 12621 14807 12679 14813
rect 12621 14804 12633 14807
rect 11848 14776 12633 14804
rect 11848 14764 11854 14776
rect 12621 14773 12633 14776
rect 12667 14804 12679 14807
rect 15102 14804 15108 14816
rect 12667 14776 15108 14804
rect 12667 14773 12679 14776
rect 12621 14767 12679 14773
rect 15102 14764 15108 14776
rect 15160 14764 15166 14816
rect 15378 14764 15384 14816
rect 15436 14804 15442 14816
rect 17880 14804 17908 14844
rect 15436 14776 17908 14804
rect 15436 14764 15442 14776
rect 17954 14764 17960 14816
rect 18012 14804 18018 14816
rect 18233 14807 18291 14813
rect 18233 14804 18245 14807
rect 18012 14776 18245 14804
rect 18012 14764 18018 14776
rect 18233 14773 18245 14776
rect 18279 14773 18291 14807
rect 18233 14767 18291 14773
rect 18414 14764 18420 14816
rect 18472 14804 18478 14816
rect 18892 14804 18920 14903
rect 19334 14900 19340 14912
rect 19392 14900 19398 14952
rect 19797 14943 19855 14949
rect 19797 14909 19809 14943
rect 19843 14909 19855 14943
rect 19978 14940 19984 14952
rect 19939 14912 19984 14940
rect 19797 14903 19855 14909
rect 19812 14872 19840 14903
rect 19978 14900 19984 14912
rect 20036 14900 20042 14952
rect 20714 14940 20720 14952
rect 20675 14912 20720 14940
rect 20714 14900 20720 14912
rect 20772 14900 20778 14952
rect 21174 14940 21180 14952
rect 21135 14912 21180 14940
rect 21174 14900 21180 14912
rect 21232 14900 21238 14952
rect 21450 14900 21456 14952
rect 21508 14940 21514 14952
rect 21821 14943 21879 14949
rect 21821 14940 21833 14943
rect 21508 14912 21833 14940
rect 21508 14900 21514 14912
rect 21821 14909 21833 14912
rect 21867 14909 21879 14943
rect 21821 14903 21879 14909
rect 22281 14943 22339 14949
rect 22281 14909 22293 14943
rect 22327 14909 22339 14943
rect 22281 14903 22339 14909
rect 20898 14872 20904 14884
rect 19812 14844 20904 14872
rect 20898 14832 20904 14844
rect 20956 14832 20962 14884
rect 21266 14832 21272 14884
rect 21324 14872 21330 14884
rect 22296 14872 22324 14903
rect 23106 14900 23112 14952
rect 23164 14940 23170 14952
rect 23661 14943 23719 14949
rect 23661 14940 23673 14943
rect 23164 14912 23673 14940
rect 23164 14900 23170 14912
rect 23661 14909 23673 14912
rect 23707 14909 23719 14943
rect 23661 14903 23719 14909
rect 24013 14943 24071 14949
rect 24013 14909 24025 14943
rect 24059 14940 24071 14943
rect 24136 14940 24164 15048
rect 24946 15036 24952 15048
rect 25004 15076 25010 15088
rect 25041 15079 25099 15085
rect 25041 15076 25053 15079
rect 25004 15048 25053 15076
rect 25004 15036 25010 15048
rect 25041 15045 25053 15048
rect 25087 15045 25099 15079
rect 25041 15039 25099 15045
rect 27890 15036 27896 15088
rect 27948 15076 27954 15088
rect 28445 15079 28503 15085
rect 28445 15076 28457 15079
rect 27948 15048 28457 15076
rect 27948 15036 27954 15048
rect 28445 15045 28457 15048
rect 28491 15045 28503 15079
rect 28445 15039 28503 15045
rect 24059 14912 24164 14940
rect 24059 14909 24071 14912
rect 24013 14903 24071 14909
rect 24486 14900 24492 14952
rect 24544 14940 24550 14952
rect 24857 14943 24915 14949
rect 24857 14940 24869 14943
rect 24544 14912 24869 14940
rect 24544 14900 24550 14912
rect 24857 14909 24869 14912
rect 24903 14909 24915 14943
rect 25590 14940 25596 14952
rect 25551 14912 25596 14940
rect 24857 14903 24915 14909
rect 25590 14900 25596 14912
rect 25648 14900 25654 14952
rect 26329 14943 26387 14949
rect 26329 14909 26341 14943
rect 26375 14940 26387 14943
rect 26418 14940 26424 14952
rect 26375 14912 26424 14940
rect 26375 14909 26387 14912
rect 26329 14903 26387 14909
rect 26418 14900 26424 14912
rect 26476 14900 26482 14952
rect 26602 14940 26608 14952
rect 26563 14912 26608 14940
rect 26602 14900 26608 14912
rect 26660 14900 26666 14952
rect 26878 14900 26884 14952
rect 26936 14940 26942 14952
rect 27522 14940 27528 14952
rect 26936 14912 27528 14940
rect 26936 14900 26942 14912
rect 27522 14900 27528 14912
rect 27580 14940 27586 14952
rect 27617 14943 27675 14949
rect 27617 14940 27629 14943
rect 27580 14912 27629 14940
rect 27580 14900 27586 14912
rect 27617 14909 27629 14912
rect 27663 14909 27675 14943
rect 27617 14903 27675 14909
rect 28077 14943 28135 14949
rect 28077 14909 28089 14943
rect 28123 14909 28135 14943
rect 28077 14903 28135 14909
rect 22554 14872 22560 14884
rect 21324 14844 22324 14872
rect 22515 14844 22560 14872
rect 21324 14832 21330 14844
rect 22554 14832 22560 14844
rect 22612 14832 22618 14884
rect 23845 14875 23903 14881
rect 23845 14872 23857 14875
rect 23676 14844 23857 14872
rect 23676 14816 23704 14844
rect 23845 14841 23857 14844
rect 23891 14872 23903 14875
rect 23891 14844 24056 14872
rect 23891 14841 23903 14844
rect 23845 14835 23903 14841
rect 20806 14804 20812 14816
rect 18472 14776 20812 14804
rect 18472 14764 18478 14776
rect 20806 14764 20812 14776
rect 20864 14764 20870 14816
rect 23658 14764 23664 14816
rect 23716 14764 23722 14816
rect 23934 14804 23940 14816
rect 23895 14776 23940 14804
rect 23934 14764 23940 14776
rect 23992 14764 23998 14816
rect 24028 14804 24056 14844
rect 24118 14832 24124 14884
rect 24176 14872 24182 14884
rect 24397 14875 24455 14881
rect 24397 14872 24409 14875
rect 24176 14844 24409 14872
rect 24176 14832 24182 14844
rect 24397 14841 24409 14844
rect 24443 14841 24455 14875
rect 28092 14872 28120 14903
rect 28166 14900 28172 14952
rect 28224 14940 28230 14952
rect 28445 14943 28503 14949
rect 28445 14940 28457 14943
rect 28224 14912 28457 14940
rect 28224 14900 28230 14912
rect 28445 14909 28457 14912
rect 28491 14909 28503 14943
rect 28445 14903 28503 14909
rect 28552 14872 28580 15116
rect 38746 15104 38752 15116
rect 38804 15104 38810 15156
rect 33134 15076 33140 15088
rect 33095 15048 33140 15076
rect 33134 15036 33140 15048
rect 33192 15036 33198 15088
rect 29546 14968 29552 15020
rect 29604 15008 29610 15020
rect 36170 15008 36176 15020
rect 29604 14980 31432 15008
rect 29604 14968 29610 14980
rect 29730 14940 29736 14952
rect 29691 14912 29736 14940
rect 29730 14900 29736 14912
rect 29788 14900 29794 14952
rect 29822 14900 29828 14952
rect 29880 14940 29886 14952
rect 29917 14943 29975 14949
rect 29917 14940 29929 14943
rect 29880 14912 29929 14940
rect 29880 14900 29886 14912
rect 29917 14909 29929 14912
rect 29963 14909 29975 14943
rect 30282 14940 30288 14952
rect 30243 14912 30288 14940
rect 29917 14903 29975 14909
rect 30282 14900 30288 14912
rect 30340 14900 30346 14952
rect 31404 14884 31432 14980
rect 32876 14980 35296 15008
rect 36131 14980 36176 15008
rect 31478 14900 31484 14952
rect 31536 14940 31542 14952
rect 32876 14949 32904 14980
rect 35268 14952 35296 14980
rect 36170 14968 36176 14980
rect 36228 14968 36234 15020
rect 36630 14968 36636 15020
rect 36688 15008 36694 15020
rect 38473 15011 38531 15017
rect 38473 15008 38485 15011
rect 36688 14980 38485 15008
rect 36688 14968 36694 14980
rect 38473 14977 38485 14980
rect 38519 14977 38531 15011
rect 38473 14971 38531 14977
rect 32309 14943 32367 14949
rect 32309 14940 32321 14943
rect 31536 14912 32321 14940
rect 31536 14900 31542 14912
rect 32309 14909 32321 14912
rect 32355 14909 32367 14943
rect 32309 14903 32367 14909
rect 32861 14943 32919 14949
rect 32861 14909 32873 14943
rect 32907 14909 32919 14943
rect 33134 14940 33140 14952
rect 33095 14912 33140 14940
rect 32861 14903 32919 14909
rect 33134 14900 33140 14912
rect 33192 14900 33198 14952
rect 34057 14943 34115 14949
rect 34057 14909 34069 14943
rect 34103 14940 34115 14943
rect 34422 14940 34428 14952
rect 34103 14912 34428 14940
rect 34103 14909 34115 14912
rect 34057 14903 34115 14909
rect 34422 14900 34428 14912
rect 34480 14900 34486 14952
rect 35250 14940 35256 14952
rect 35211 14912 35256 14940
rect 35250 14900 35256 14912
rect 35308 14900 35314 14952
rect 35710 14940 35716 14952
rect 35671 14912 35716 14940
rect 35710 14900 35716 14912
rect 35768 14900 35774 14952
rect 36265 14943 36323 14949
rect 36265 14909 36277 14943
rect 36311 14940 36323 14943
rect 36354 14940 36360 14952
rect 36311 14912 36360 14940
rect 36311 14909 36323 14912
rect 36265 14903 36323 14909
rect 36354 14900 36360 14912
rect 36412 14900 36418 14952
rect 36449 14943 36507 14949
rect 36449 14909 36461 14943
rect 36495 14909 36507 14943
rect 36449 14903 36507 14909
rect 28718 14872 28724 14884
rect 28092 14844 28488 14872
rect 28552 14844 28724 14872
rect 24397 14835 24455 14841
rect 25406 14804 25412 14816
rect 24028 14776 25412 14804
rect 25406 14764 25412 14776
rect 25464 14764 25470 14816
rect 25685 14807 25743 14813
rect 25685 14773 25697 14807
rect 25731 14804 25743 14807
rect 26050 14804 26056 14816
rect 25731 14776 26056 14804
rect 25731 14773 25743 14776
rect 25685 14767 25743 14773
rect 26050 14764 26056 14776
rect 26108 14764 26114 14816
rect 28460 14804 28488 14844
rect 28718 14832 28724 14844
rect 28776 14872 28782 14884
rect 28776 14844 30420 14872
rect 28776 14832 28782 14844
rect 29549 14807 29607 14813
rect 29549 14804 29561 14807
rect 28460 14776 29561 14804
rect 29549 14773 29561 14776
rect 29595 14804 29607 14807
rect 30282 14804 30288 14816
rect 29595 14776 30288 14804
rect 29595 14773 29607 14776
rect 29549 14767 29607 14773
rect 30282 14764 30288 14776
rect 30340 14764 30346 14816
rect 30392 14804 30420 14844
rect 30558 14832 30564 14884
rect 30616 14872 30622 14884
rect 31021 14875 31079 14881
rect 31021 14872 31033 14875
rect 30616 14844 31033 14872
rect 30616 14832 30622 14844
rect 31021 14841 31033 14844
rect 31067 14841 31079 14875
rect 31021 14835 31079 14841
rect 31110 14832 31116 14884
rect 31168 14872 31174 14884
rect 31297 14875 31355 14881
rect 31297 14872 31309 14875
rect 31168 14844 31309 14872
rect 31168 14832 31174 14844
rect 31297 14841 31309 14844
rect 31343 14841 31355 14875
rect 31297 14835 31355 14841
rect 31386 14832 31392 14884
rect 31444 14872 31450 14884
rect 31757 14875 31815 14881
rect 31444 14844 31489 14872
rect 31444 14832 31450 14844
rect 31757 14841 31769 14875
rect 31803 14872 31815 14875
rect 32214 14872 32220 14884
rect 31803 14844 32220 14872
rect 31803 14841 31815 14844
rect 31757 14835 31815 14841
rect 32214 14832 32220 14844
rect 32272 14832 32278 14884
rect 33962 14832 33968 14884
rect 34020 14872 34026 14884
rect 36464 14872 36492 14903
rect 36538 14900 36544 14952
rect 36596 14940 36602 14952
rect 36909 14943 36967 14949
rect 36909 14940 36921 14943
rect 36596 14912 36921 14940
rect 36596 14900 36602 14912
rect 36909 14909 36921 14912
rect 36955 14909 36967 14943
rect 37734 14940 37740 14952
rect 37695 14912 37740 14940
rect 36909 14903 36967 14909
rect 37734 14900 37740 14912
rect 37792 14900 37798 14952
rect 38562 14900 38568 14952
rect 38620 14940 38626 14952
rect 38620 14912 38665 14940
rect 38620 14900 38626 14912
rect 34020 14844 36492 14872
rect 34020 14832 34026 14844
rect 31205 14807 31263 14813
rect 31205 14804 31217 14807
rect 30392 14776 31217 14804
rect 31205 14773 31217 14776
rect 31251 14773 31263 14807
rect 31205 14767 31263 14773
rect 34241 14807 34299 14813
rect 34241 14773 34253 14807
rect 34287 14804 34299 14807
rect 34330 14804 34336 14816
rect 34287 14776 34336 14804
rect 34287 14773 34299 14776
rect 34241 14767 34299 14773
rect 34330 14764 34336 14776
rect 34388 14764 34394 14816
rect 37826 14764 37832 14816
rect 37884 14804 37890 14816
rect 37921 14807 37979 14813
rect 37921 14804 37933 14807
rect 37884 14776 37933 14804
rect 37884 14764 37890 14776
rect 37921 14773 37933 14776
rect 37967 14773 37979 14807
rect 37921 14767 37979 14773
rect 1104 14714 39836 14736
rect 1104 14662 19606 14714
rect 19658 14662 19670 14714
rect 19722 14662 19734 14714
rect 19786 14662 19798 14714
rect 19850 14662 39836 14714
rect 1104 14640 39836 14662
rect 1854 14560 1860 14612
rect 1912 14600 1918 14612
rect 2041 14603 2099 14609
rect 2041 14600 2053 14603
rect 1912 14572 2053 14600
rect 1912 14560 1918 14572
rect 2041 14569 2053 14572
rect 2087 14569 2099 14603
rect 2041 14563 2099 14569
rect 3970 14560 3976 14612
rect 4028 14600 4034 14612
rect 4028 14572 11192 14600
rect 4028 14560 4034 14572
rect 4798 14532 4804 14544
rect 4759 14504 4804 14532
rect 4798 14492 4804 14504
rect 4856 14492 4862 14544
rect 8110 14492 8116 14544
rect 8168 14532 8174 14544
rect 10318 14532 10324 14544
rect 8168 14504 10324 14532
rect 8168 14492 8174 14504
rect 1946 14424 1952 14476
rect 2004 14464 2010 14476
rect 2225 14467 2283 14473
rect 2225 14464 2237 14467
rect 2004 14436 2237 14464
rect 2004 14424 2010 14436
rect 2225 14433 2237 14436
rect 2271 14433 2283 14467
rect 2498 14464 2504 14476
rect 2459 14436 2504 14464
rect 2225 14427 2283 14433
rect 2240 14396 2268 14427
rect 2498 14424 2504 14436
rect 2556 14424 2562 14476
rect 3234 14464 3240 14476
rect 3195 14436 3240 14464
rect 3234 14424 3240 14436
rect 3292 14424 3298 14476
rect 4341 14467 4399 14473
rect 4341 14433 4353 14467
rect 4387 14433 4399 14467
rect 4341 14427 4399 14433
rect 4617 14467 4675 14473
rect 4617 14433 4629 14467
rect 4663 14464 4675 14467
rect 5442 14464 5448 14476
rect 4663 14436 5448 14464
rect 4663 14433 4675 14436
rect 4617 14427 4675 14433
rect 4062 14396 4068 14408
rect 2240 14368 4068 14396
rect 4062 14356 4068 14368
rect 4120 14396 4126 14408
rect 4356 14396 4384 14427
rect 5442 14424 5448 14436
rect 5500 14424 5506 14476
rect 8404 14473 8432 14504
rect 10318 14492 10324 14504
rect 10376 14492 10382 14544
rect 11164 14532 11192 14572
rect 11514 14560 11520 14612
rect 11572 14600 11578 14612
rect 11609 14603 11667 14609
rect 11609 14600 11621 14603
rect 11572 14572 11621 14600
rect 11572 14560 11578 14572
rect 11609 14569 11621 14572
rect 11655 14569 11667 14603
rect 11609 14563 11667 14569
rect 11882 14560 11888 14612
rect 11940 14600 11946 14612
rect 15654 14600 15660 14612
rect 11940 14572 15660 14600
rect 11940 14560 11946 14572
rect 15654 14560 15660 14572
rect 15712 14560 15718 14612
rect 15838 14560 15844 14612
rect 15896 14600 15902 14612
rect 16669 14603 16727 14609
rect 16669 14600 16681 14603
rect 15896 14572 16681 14600
rect 15896 14560 15902 14572
rect 16669 14569 16681 14572
rect 16715 14569 16727 14603
rect 16669 14563 16727 14569
rect 18506 14560 18512 14612
rect 18564 14600 18570 14612
rect 20073 14603 20131 14609
rect 20073 14600 20085 14603
rect 18564 14572 20085 14600
rect 18564 14560 18570 14572
rect 20073 14569 20085 14572
rect 20119 14569 20131 14603
rect 22002 14600 22008 14612
rect 20073 14563 20131 14569
rect 21008 14572 22008 14600
rect 13354 14532 13360 14544
rect 11164 14504 13360 14532
rect 13354 14492 13360 14504
rect 13412 14492 13418 14544
rect 18874 14492 18880 14544
rect 18932 14532 18938 14544
rect 21008 14532 21036 14572
rect 22002 14560 22008 14572
rect 22060 14560 22066 14612
rect 23658 14560 23664 14612
rect 23716 14600 23722 14612
rect 23937 14603 23995 14609
rect 23937 14600 23949 14603
rect 23716 14572 23949 14600
rect 23716 14560 23722 14572
rect 23937 14569 23949 14572
rect 23983 14569 23995 14603
rect 23937 14563 23995 14569
rect 24029 14603 24087 14609
rect 24029 14569 24041 14603
rect 24075 14600 24087 14603
rect 24210 14600 24216 14612
rect 24075 14572 24216 14600
rect 24075 14569 24087 14572
rect 24029 14563 24087 14569
rect 24210 14560 24216 14572
rect 24268 14560 24274 14612
rect 26602 14600 26608 14612
rect 26563 14572 26608 14600
rect 26602 14560 26608 14572
rect 26660 14560 26666 14612
rect 28261 14603 28319 14609
rect 28261 14569 28273 14603
rect 28307 14600 28319 14603
rect 28810 14600 28816 14612
rect 28307 14572 28816 14600
rect 28307 14569 28319 14572
rect 28261 14563 28319 14569
rect 28810 14560 28816 14572
rect 28868 14560 28874 14612
rect 30558 14600 30564 14612
rect 30519 14572 30564 14600
rect 30558 14560 30564 14572
rect 30616 14560 30622 14612
rect 37093 14603 37151 14609
rect 37093 14569 37105 14603
rect 37139 14600 37151 14603
rect 38562 14600 38568 14612
rect 37139 14572 38568 14600
rect 37139 14569 37151 14572
rect 37093 14563 37151 14569
rect 38562 14560 38568 14572
rect 38620 14560 38626 14612
rect 18932 14504 21036 14532
rect 18932 14492 18938 14504
rect 23382 14492 23388 14544
rect 23440 14532 23446 14544
rect 24121 14535 24179 14541
rect 24121 14532 24133 14535
rect 23440 14504 24133 14532
rect 23440 14492 23446 14504
rect 24121 14501 24133 14504
rect 24167 14501 24179 14535
rect 24121 14495 24179 14501
rect 26418 14492 26424 14544
rect 26476 14532 26482 14544
rect 30009 14535 30067 14541
rect 30009 14532 30021 14535
rect 26476 14504 30021 14532
rect 26476 14492 26482 14504
rect 30009 14501 30021 14504
rect 30055 14501 30067 14535
rect 30009 14495 30067 14501
rect 30742 14492 30748 14544
rect 30800 14532 30806 14544
rect 32858 14532 32864 14544
rect 30800 14504 32864 14532
rect 30800 14492 30806 14504
rect 32858 14492 32864 14504
rect 32916 14492 32922 14544
rect 33318 14492 33324 14544
rect 33376 14532 33382 14544
rect 34330 14532 34336 14544
rect 33376 14504 34336 14532
rect 33376 14492 33382 14504
rect 34330 14492 34336 14504
rect 34388 14532 34394 14544
rect 37734 14532 37740 14544
rect 34388 14504 34468 14532
rect 34388 14492 34394 14504
rect 8389 14467 8447 14473
rect 8389 14433 8401 14467
rect 8435 14433 8447 14467
rect 8389 14427 8447 14433
rect 8573 14467 8631 14473
rect 8573 14433 8585 14467
rect 8619 14464 8631 14467
rect 9030 14464 9036 14476
rect 8619 14436 9036 14464
rect 8619 14433 8631 14436
rect 8573 14427 8631 14433
rect 9030 14424 9036 14436
rect 9088 14424 9094 14476
rect 10226 14464 10232 14476
rect 10187 14436 10232 14464
rect 10226 14424 10232 14436
rect 10284 14424 10290 14476
rect 10502 14464 10508 14476
rect 10463 14436 10508 14464
rect 10502 14424 10508 14436
rect 10560 14424 10566 14476
rect 10594 14424 10600 14476
rect 10652 14464 10658 14476
rect 13449 14467 13507 14473
rect 10652 14436 13124 14464
rect 10652 14424 10658 14436
rect 5074 14396 5080 14408
rect 4120 14368 5080 14396
rect 4120 14356 4126 14368
rect 5074 14356 5080 14368
rect 5132 14356 5138 14408
rect 5905 14399 5963 14405
rect 5905 14365 5917 14399
rect 5951 14365 5963 14399
rect 6178 14396 6184 14408
rect 6139 14368 6184 14396
rect 5905 14359 5963 14365
rect 3418 14260 3424 14272
rect 3379 14232 3424 14260
rect 3418 14220 3424 14232
rect 3476 14220 3482 14272
rect 5920 14260 5948 14359
rect 6178 14356 6184 14368
rect 6236 14356 6242 14408
rect 8662 14396 8668 14408
rect 8623 14368 8668 14396
rect 8662 14356 8668 14368
rect 8720 14356 8726 14408
rect 13096 14405 13124 14436
rect 13449 14433 13461 14467
rect 13495 14464 13507 14467
rect 13538 14464 13544 14476
rect 13495 14436 13544 14464
rect 13495 14433 13507 14436
rect 13449 14427 13507 14433
rect 13538 14424 13544 14436
rect 13596 14424 13602 14476
rect 13814 14464 13820 14476
rect 13775 14436 13820 14464
rect 13814 14424 13820 14436
rect 13872 14424 13878 14476
rect 14458 14464 14464 14476
rect 14419 14436 14464 14464
rect 14458 14424 14464 14436
rect 14516 14424 14522 14476
rect 15565 14467 15623 14473
rect 15565 14433 15577 14467
rect 15611 14464 15623 14467
rect 16482 14464 16488 14476
rect 15611 14436 16488 14464
rect 15611 14433 15623 14436
rect 15565 14427 15623 14433
rect 16482 14424 16488 14436
rect 16540 14424 16546 14476
rect 17880 14436 18276 14464
rect 13081 14399 13139 14405
rect 13081 14365 13093 14399
rect 13127 14396 13139 14399
rect 15289 14399 15347 14405
rect 13127 14368 14136 14396
rect 13127 14365 13139 14368
rect 13081 14359 13139 14365
rect 9950 14328 9956 14340
rect 7392 14300 9956 14328
rect 7392 14260 7420 14300
rect 9950 14288 9956 14300
rect 10008 14288 10014 14340
rect 12526 14288 12532 14340
rect 12584 14328 12590 14340
rect 12986 14328 12992 14340
rect 12584 14300 12992 14328
rect 12584 14288 12590 14300
rect 12986 14288 12992 14300
rect 13044 14288 13050 14340
rect 13262 14288 13268 14340
rect 13320 14328 13326 14340
rect 13725 14331 13783 14337
rect 13725 14328 13737 14331
rect 13320 14300 13737 14328
rect 13320 14288 13326 14300
rect 13725 14297 13737 14300
rect 13771 14297 13783 14331
rect 14108 14328 14136 14368
rect 15289 14365 15301 14399
rect 15335 14396 15347 14399
rect 17773 14399 17831 14405
rect 17773 14396 17785 14399
rect 15335 14368 17785 14396
rect 15335 14365 15347 14368
rect 15289 14359 15347 14365
rect 17773 14365 17785 14368
rect 17819 14396 17831 14399
rect 17880 14396 17908 14436
rect 18046 14396 18052 14408
rect 17819 14368 17908 14396
rect 18007 14368 18052 14396
rect 17819 14365 17831 14368
rect 17773 14359 17831 14365
rect 18046 14356 18052 14368
rect 18104 14356 18110 14408
rect 18248 14396 18276 14436
rect 19702 14424 19708 14476
rect 19760 14464 19766 14476
rect 19877 14467 19935 14473
rect 19877 14464 19889 14467
rect 19760 14436 19889 14464
rect 19760 14424 19766 14436
rect 19877 14433 19889 14436
rect 19923 14433 19935 14467
rect 23014 14464 23020 14476
rect 22975 14436 23020 14464
rect 19877 14427 19935 14433
rect 23014 14424 23020 14436
rect 23072 14424 23078 14476
rect 23106 14424 23112 14476
rect 23164 14464 23170 14476
rect 23753 14467 23811 14473
rect 23753 14464 23765 14467
rect 23164 14436 23765 14464
rect 23164 14424 23170 14436
rect 23753 14433 23765 14436
rect 23799 14433 23811 14467
rect 24946 14464 24952 14476
rect 23753 14427 23811 14433
rect 23860 14436 24952 14464
rect 18690 14396 18696 14408
rect 18248 14368 18696 14396
rect 18690 14356 18696 14368
rect 18748 14396 18754 14408
rect 20901 14399 20959 14405
rect 20901 14396 20913 14399
rect 18748 14368 20913 14396
rect 18748 14356 18754 14368
rect 20901 14365 20913 14368
rect 20947 14365 20959 14399
rect 21174 14396 21180 14408
rect 21135 14368 21180 14396
rect 20901 14359 20959 14365
rect 21174 14356 21180 14368
rect 21232 14356 21238 14408
rect 22738 14356 22744 14408
rect 22796 14396 22802 14408
rect 23860 14396 23888 14436
rect 24946 14424 24952 14436
rect 25004 14424 25010 14476
rect 25409 14467 25467 14473
rect 25409 14433 25421 14467
rect 25455 14433 25467 14467
rect 25409 14427 25467 14433
rect 24486 14396 24492 14408
rect 22796 14368 23888 14396
rect 24447 14368 24492 14396
rect 22796 14356 22802 14368
rect 24486 14356 24492 14368
rect 24544 14356 24550 14408
rect 25424 14396 25452 14427
rect 25498 14424 25504 14476
rect 25556 14464 25562 14476
rect 25593 14467 25651 14473
rect 25593 14464 25605 14467
rect 25556 14436 25605 14464
rect 25556 14424 25562 14436
rect 25593 14433 25605 14436
rect 25639 14433 25651 14467
rect 25593 14427 25651 14433
rect 25777 14467 25835 14473
rect 25777 14433 25789 14467
rect 25823 14464 25835 14467
rect 26694 14464 26700 14476
rect 25823 14436 26700 14464
rect 25823 14433 25835 14436
rect 25777 14427 25835 14433
rect 26694 14424 26700 14436
rect 26752 14424 26758 14476
rect 27065 14467 27123 14473
rect 27065 14433 27077 14467
rect 27111 14433 27123 14467
rect 27065 14427 27123 14433
rect 25424 14368 25912 14396
rect 20162 14328 20168 14340
rect 14108 14300 15332 14328
rect 13725 14291 13783 14297
rect 5920 14232 7420 14260
rect 7469 14263 7527 14269
rect 7469 14229 7481 14263
rect 7515 14260 7527 14263
rect 7558 14260 7564 14272
rect 7515 14232 7564 14260
rect 7515 14229 7527 14232
rect 7469 14223 7527 14229
rect 7558 14220 7564 14232
rect 7616 14220 7622 14272
rect 14645 14263 14703 14269
rect 14645 14229 14657 14263
rect 14691 14260 14703 14263
rect 15194 14260 15200 14272
rect 14691 14232 15200 14260
rect 14691 14229 14703 14232
rect 14645 14223 14703 14229
rect 15194 14220 15200 14232
rect 15252 14220 15258 14272
rect 15304 14260 15332 14300
rect 18708 14300 20168 14328
rect 18708 14260 18736 14300
rect 20162 14288 20168 14300
rect 20220 14288 20226 14340
rect 25225 14331 25283 14337
rect 25225 14297 25237 14331
rect 25271 14328 25283 14331
rect 25590 14328 25596 14340
rect 25271 14300 25596 14328
rect 25271 14297 25283 14300
rect 25225 14291 25283 14297
rect 25590 14288 25596 14300
rect 25648 14288 25654 14340
rect 25884 14328 25912 14368
rect 25958 14356 25964 14408
rect 26016 14396 26022 14408
rect 27080 14396 27108 14427
rect 27890 14424 27896 14476
rect 27948 14464 27954 14476
rect 28077 14467 28135 14473
rect 28077 14464 28089 14467
rect 27948 14436 28089 14464
rect 27948 14424 27954 14436
rect 28077 14433 28089 14436
rect 28123 14433 28135 14467
rect 29270 14464 29276 14476
rect 29231 14436 29276 14464
rect 28077 14427 28135 14433
rect 29270 14424 29276 14436
rect 29328 14424 29334 14476
rect 29822 14464 29828 14476
rect 29783 14436 29828 14464
rect 29822 14424 29828 14436
rect 29880 14424 29886 14476
rect 29914 14424 29920 14476
rect 29972 14464 29978 14476
rect 30469 14467 30527 14473
rect 30469 14464 30481 14467
rect 29972 14436 30481 14464
rect 29972 14424 29978 14436
rect 30469 14433 30481 14436
rect 30515 14433 30527 14467
rect 30469 14427 30527 14433
rect 30929 14467 30987 14473
rect 30929 14433 30941 14467
rect 30975 14433 30987 14467
rect 32582 14464 32588 14476
rect 32543 14436 32588 14464
rect 30929 14427 30987 14433
rect 26016 14368 27108 14396
rect 27525 14399 27583 14405
rect 26016 14356 26022 14368
rect 27525 14365 27537 14399
rect 27571 14396 27583 14399
rect 27614 14396 27620 14408
rect 27571 14368 27620 14396
rect 27571 14365 27583 14368
rect 27525 14359 27583 14365
rect 27614 14356 27620 14368
rect 27672 14396 27678 14408
rect 28442 14396 28448 14408
rect 27672 14368 28448 14396
rect 27672 14356 27678 14368
rect 28442 14356 28448 14368
rect 28500 14356 28506 14408
rect 29089 14399 29147 14405
rect 29089 14365 29101 14399
rect 29135 14396 29147 14399
rect 29730 14396 29736 14408
rect 29135 14368 29736 14396
rect 29135 14365 29147 14368
rect 29089 14359 29147 14365
rect 29730 14356 29736 14368
rect 29788 14356 29794 14408
rect 30190 14356 30196 14408
rect 30248 14396 30254 14408
rect 30944 14396 30972 14427
rect 32582 14424 32588 14436
rect 32640 14424 32646 14476
rect 32953 14467 33011 14473
rect 32953 14433 32965 14467
rect 32999 14464 33011 14467
rect 32999 14436 33640 14464
rect 32999 14433 33011 14436
rect 32953 14427 33011 14433
rect 33612 14408 33640 14436
rect 33962 14424 33968 14476
rect 34020 14464 34026 14476
rect 34440 14473 34468 14504
rect 36464 14504 37740 14532
rect 34057 14467 34115 14473
rect 34057 14464 34069 14467
rect 34020 14436 34069 14464
rect 34020 14424 34026 14436
rect 34057 14433 34069 14436
rect 34103 14433 34115 14467
rect 34241 14467 34299 14473
rect 34241 14464 34253 14467
rect 34057 14427 34115 14433
rect 34164 14436 34253 14464
rect 30248 14368 30972 14396
rect 33045 14399 33103 14405
rect 30248 14356 30254 14368
rect 33045 14365 33057 14399
rect 33091 14396 33103 14399
rect 33226 14396 33232 14408
rect 33091 14368 33232 14396
rect 33091 14365 33103 14368
rect 33045 14359 33103 14365
rect 33226 14356 33232 14368
rect 33284 14356 33290 14408
rect 33594 14396 33600 14408
rect 33555 14368 33600 14396
rect 33594 14356 33600 14368
rect 33652 14356 33658 14408
rect 27062 14328 27068 14340
rect 25884 14300 27068 14328
rect 27062 14288 27068 14300
rect 27120 14288 27126 14340
rect 32401 14331 32459 14337
rect 32401 14297 32413 14331
rect 32447 14328 32459 14331
rect 33686 14328 33692 14340
rect 32447 14300 33692 14328
rect 32447 14297 32459 14300
rect 32401 14291 32459 14297
rect 33686 14288 33692 14300
rect 33744 14288 33750 14340
rect 15304 14232 18736 14260
rect 19337 14263 19395 14269
rect 19337 14229 19349 14263
rect 19383 14260 19395 14263
rect 19426 14260 19432 14272
rect 19383 14232 19432 14260
rect 19383 14229 19395 14232
rect 19337 14223 19395 14229
rect 19426 14220 19432 14232
rect 19484 14220 19490 14272
rect 21358 14220 21364 14272
rect 21416 14260 21422 14272
rect 22281 14263 22339 14269
rect 22281 14260 22293 14263
rect 21416 14232 22293 14260
rect 21416 14220 21422 14232
rect 22281 14229 22293 14232
rect 22327 14229 22339 14263
rect 22281 14223 22339 14229
rect 23201 14263 23259 14269
rect 23201 14229 23213 14263
rect 23247 14260 23259 14263
rect 23290 14260 23296 14272
rect 23247 14232 23296 14260
rect 23247 14229 23259 14232
rect 23201 14223 23259 14229
rect 23290 14220 23296 14232
rect 23348 14260 23354 14272
rect 23566 14260 23572 14272
rect 23348 14232 23572 14260
rect 23348 14220 23354 14232
rect 23566 14220 23572 14232
rect 23624 14220 23630 14272
rect 29270 14220 29276 14272
rect 29328 14260 29334 14272
rect 34164 14260 34192 14436
rect 34241 14433 34253 14436
rect 34287 14433 34299 14467
rect 34241 14427 34299 14433
rect 34425 14467 34483 14473
rect 34425 14433 34437 14467
rect 34471 14433 34483 14467
rect 34606 14464 34612 14476
rect 34567 14436 34612 14464
rect 34425 14427 34483 14433
rect 34606 14424 34612 14436
rect 34664 14424 34670 14476
rect 34790 14424 34796 14476
rect 34848 14464 34854 14476
rect 34885 14467 34943 14473
rect 34885 14464 34897 14467
rect 34848 14436 34897 14464
rect 34848 14424 34854 14436
rect 34885 14433 34897 14436
rect 34931 14433 34943 14467
rect 34885 14427 34943 14433
rect 36170 14424 36176 14476
rect 36228 14464 36234 14476
rect 36464 14464 36492 14504
rect 37734 14492 37740 14504
rect 37792 14532 37798 14544
rect 38105 14535 38163 14541
rect 38105 14532 38117 14535
rect 37792 14504 38117 14532
rect 37792 14492 37798 14504
rect 38105 14501 38117 14504
rect 38151 14501 38163 14535
rect 38105 14495 38163 14501
rect 38473 14535 38531 14541
rect 38473 14501 38485 14535
rect 38519 14532 38531 14535
rect 38654 14532 38660 14544
rect 38519 14504 38660 14532
rect 38519 14501 38531 14504
rect 38473 14495 38531 14501
rect 38654 14492 38660 14504
rect 38712 14492 38718 14544
rect 37918 14464 37924 14476
rect 36228 14436 36492 14464
rect 37879 14436 37924 14464
rect 36228 14424 36234 14436
rect 37918 14424 37924 14436
rect 37976 14424 37982 14476
rect 38010 14424 38016 14476
rect 38068 14464 38074 14476
rect 38930 14464 38936 14476
rect 38068 14436 38113 14464
rect 38891 14436 38936 14464
rect 38068 14424 38074 14436
rect 38930 14424 38936 14436
rect 38988 14424 38994 14476
rect 34330 14356 34336 14408
rect 34388 14396 34394 14408
rect 35529 14399 35587 14405
rect 35529 14396 35541 14399
rect 34388 14368 35541 14396
rect 34388 14356 34394 14368
rect 35529 14365 35541 14368
rect 35575 14365 35587 14399
rect 35529 14359 35587 14365
rect 35805 14399 35863 14405
rect 35805 14365 35817 14399
rect 35851 14396 35863 14399
rect 36906 14396 36912 14408
rect 35851 14368 36912 14396
rect 35851 14365 35863 14368
rect 35805 14359 35863 14365
rect 36906 14356 36912 14368
rect 36964 14356 36970 14408
rect 37734 14396 37740 14408
rect 37695 14368 37740 14396
rect 37734 14356 37740 14368
rect 37792 14356 37798 14408
rect 35434 14260 35440 14272
rect 29328 14232 35440 14260
rect 29328 14220 29334 14232
rect 35434 14220 35440 14232
rect 35492 14220 35498 14272
rect 35526 14220 35532 14272
rect 35584 14260 35590 14272
rect 39025 14263 39083 14269
rect 39025 14260 39037 14263
rect 35584 14232 39037 14260
rect 35584 14220 35590 14232
rect 39025 14229 39037 14232
rect 39071 14229 39083 14263
rect 39025 14223 39083 14229
rect 1104 14170 39836 14192
rect 1104 14118 4246 14170
rect 4298 14118 4310 14170
rect 4362 14118 4374 14170
rect 4426 14118 4438 14170
rect 4490 14118 34966 14170
rect 35018 14118 35030 14170
rect 35082 14118 35094 14170
rect 35146 14118 35158 14170
rect 35210 14118 39836 14170
rect 1104 14096 39836 14118
rect 4908 14028 8524 14056
rect 3789 13991 3847 13997
rect 3789 13957 3801 13991
rect 3835 13988 3847 13991
rect 3878 13988 3884 14000
rect 3835 13960 3884 13988
rect 3835 13957 3847 13960
rect 3789 13951 3847 13957
rect 3878 13948 3884 13960
rect 3936 13948 3942 14000
rect 1486 13880 1492 13932
rect 1544 13920 1550 13932
rect 1581 13923 1639 13929
rect 1581 13920 1593 13923
rect 1544 13892 1593 13920
rect 1544 13880 1550 13892
rect 1581 13889 1593 13892
rect 1627 13889 1639 13923
rect 1854 13920 1860 13932
rect 1815 13892 1860 13920
rect 1581 13883 1639 13889
rect 1854 13880 1860 13892
rect 1912 13880 1918 13932
rect 4614 13920 4620 13932
rect 4575 13892 4620 13920
rect 4614 13880 4620 13892
rect 4672 13880 4678 13932
rect 3970 13852 3976 13864
rect 3931 13824 3976 13852
rect 3970 13812 3976 13824
rect 4028 13812 4034 13864
rect 4154 13852 4160 13864
rect 4115 13824 4160 13852
rect 4154 13812 4160 13824
rect 4212 13812 4218 13864
rect 4525 13855 4583 13861
rect 4525 13821 4537 13855
rect 4571 13852 4583 13855
rect 4908 13852 4936 14028
rect 6178 13948 6184 14000
rect 6236 13988 6242 14000
rect 8297 13991 8355 13997
rect 8297 13988 8309 13991
rect 6236 13960 8309 13988
rect 6236 13948 6242 13960
rect 8297 13957 8309 13960
rect 8343 13957 8355 13991
rect 8496 13988 8524 14028
rect 8938 14016 8944 14068
rect 8996 14056 9002 14068
rect 9306 14056 9312 14068
rect 8996 14028 9312 14056
rect 8996 14016 9002 14028
rect 9306 14016 9312 14028
rect 9364 14056 9370 14068
rect 11422 14056 11428 14068
rect 9364 14028 11428 14056
rect 9364 14016 9370 14028
rect 11422 14016 11428 14028
rect 11480 14016 11486 14068
rect 13814 14016 13820 14068
rect 13872 14056 13878 14068
rect 14737 14059 14795 14065
rect 14737 14056 14749 14059
rect 13872 14028 14749 14056
rect 13872 14016 13878 14028
rect 14737 14025 14749 14028
rect 14783 14025 14795 14059
rect 14737 14019 14795 14025
rect 19242 14016 19248 14068
rect 19300 14056 19306 14068
rect 20898 14056 20904 14068
rect 19300 14028 20904 14056
rect 19300 14016 19306 14028
rect 20898 14016 20904 14028
rect 20956 14016 20962 14068
rect 24854 14016 24860 14068
rect 24912 14056 24918 14068
rect 25041 14059 25099 14065
rect 25041 14056 25053 14059
rect 24912 14028 25053 14056
rect 24912 14016 24918 14028
rect 25041 14025 25053 14028
rect 25087 14025 25099 14059
rect 25041 14019 25099 14025
rect 27522 14016 27528 14068
rect 27580 14056 27586 14068
rect 28629 14059 28687 14065
rect 28629 14056 28641 14059
rect 27580 14028 28641 14056
rect 27580 14016 27586 14028
rect 28629 14025 28641 14028
rect 28675 14025 28687 14059
rect 28629 14019 28687 14025
rect 29273 14059 29331 14065
rect 29273 14025 29285 14059
rect 29319 14056 29331 14059
rect 30374 14056 30380 14068
rect 29319 14028 30380 14056
rect 29319 14025 29331 14028
rect 29273 14019 29331 14025
rect 12434 13988 12440 14000
rect 8496 13960 12440 13988
rect 8297 13951 8355 13957
rect 12434 13948 12440 13960
rect 12492 13948 12498 14000
rect 16482 13948 16488 14000
rect 16540 13988 16546 14000
rect 17954 13988 17960 14000
rect 16540 13960 16585 13988
rect 16684 13960 17960 13988
rect 16540 13948 16546 13960
rect 5258 13920 5264 13932
rect 5219 13892 5264 13920
rect 5258 13880 5264 13892
rect 5316 13880 5322 13932
rect 10042 13880 10048 13932
rect 10100 13920 10106 13932
rect 15562 13920 15568 13932
rect 10100 13892 15568 13920
rect 10100 13880 10106 13892
rect 15562 13880 15568 13892
rect 15620 13880 15626 13932
rect 16684 13920 16712 13960
rect 17954 13948 17960 13960
rect 18012 13948 18018 14000
rect 18046 13948 18052 14000
rect 18104 13988 18110 14000
rect 18325 13991 18383 13997
rect 18325 13988 18337 13991
rect 18104 13960 18337 13988
rect 18104 13948 18110 13960
rect 18325 13957 18337 13960
rect 18371 13957 18383 13991
rect 18325 13951 18383 13957
rect 19610 13948 19616 14000
rect 19668 13988 19674 14000
rect 19978 13988 19984 14000
rect 19668 13960 19984 13988
rect 19668 13948 19674 13960
rect 19978 13948 19984 13960
rect 20036 13988 20042 14000
rect 28644 13988 28672 14019
rect 30374 14016 30380 14028
rect 30432 14056 30438 14068
rect 31478 14056 31484 14068
rect 30432 14028 31484 14056
rect 30432 14016 30438 14028
rect 31478 14016 31484 14028
rect 31536 14016 31542 14068
rect 34330 14016 34336 14068
rect 34388 14056 34394 14068
rect 34425 14059 34483 14065
rect 34425 14056 34437 14059
rect 34388 14028 34437 14056
rect 34388 14016 34394 14028
rect 34425 14025 34437 14028
rect 34471 14025 34483 14059
rect 34425 14019 34483 14025
rect 35526 14016 35532 14068
rect 35584 14016 35590 14068
rect 37826 14056 37832 14068
rect 35728 14028 37832 14056
rect 31110 13988 31116 14000
rect 20036 13960 21956 13988
rect 28644 13960 31116 13988
rect 20036 13948 20042 13960
rect 15672 13892 16712 13920
rect 17313 13923 17371 13929
rect 5350 13852 5356 13864
rect 4571 13824 4936 13852
rect 5311 13824 5356 13852
rect 4571 13821 4583 13824
rect 4525 13815 4583 13821
rect 5350 13812 5356 13824
rect 5408 13812 5414 13864
rect 5810 13852 5816 13864
rect 5771 13824 5816 13852
rect 5810 13812 5816 13824
rect 5868 13812 5874 13864
rect 7193 13855 7251 13861
rect 7193 13821 7205 13855
rect 7239 13821 7251 13855
rect 7374 13852 7380 13864
rect 7335 13824 7380 13852
rect 7193 13815 7251 13821
rect 2958 13716 2964 13728
rect 2919 13688 2964 13716
rect 2958 13676 2964 13688
rect 3016 13676 3022 13728
rect 7208 13716 7236 13815
rect 7374 13812 7380 13824
rect 7432 13812 7438 13864
rect 7558 13852 7564 13864
rect 7519 13824 7564 13852
rect 7558 13812 7564 13824
rect 7616 13812 7622 13864
rect 8202 13852 8208 13864
rect 8163 13824 8208 13852
rect 8202 13812 8208 13824
rect 8260 13812 8266 13864
rect 8665 13855 8723 13861
rect 8665 13852 8677 13855
rect 8312 13824 8677 13852
rect 7650 13744 7656 13796
rect 7708 13784 7714 13796
rect 8312 13784 8340 13824
rect 8665 13821 8677 13824
rect 8711 13821 8723 13855
rect 9214 13852 9220 13864
rect 9175 13824 9220 13852
rect 8665 13815 8723 13821
rect 9214 13812 9220 13824
rect 9272 13812 9278 13864
rect 9582 13852 9588 13864
rect 9543 13824 9588 13852
rect 9582 13812 9588 13824
rect 9640 13812 9646 13864
rect 10134 13852 10140 13864
rect 10095 13824 10140 13852
rect 10134 13812 10140 13824
rect 10192 13812 10198 13864
rect 11149 13855 11207 13861
rect 11149 13821 11161 13855
rect 11195 13821 11207 13855
rect 11514 13852 11520 13864
rect 11475 13824 11520 13852
rect 11149 13815 11207 13821
rect 7708 13756 8340 13784
rect 7708 13744 7714 13756
rect 9858 13744 9864 13796
rect 9916 13784 9922 13796
rect 10962 13784 10968 13796
rect 9916 13756 10968 13784
rect 9916 13744 9922 13756
rect 10962 13744 10968 13756
rect 11020 13784 11026 13796
rect 11164 13784 11192 13815
rect 11514 13812 11520 13824
rect 11572 13812 11578 13864
rect 11882 13852 11888 13864
rect 11843 13824 11888 13852
rect 11882 13812 11888 13824
rect 11940 13812 11946 13864
rect 12526 13852 12532 13864
rect 12487 13824 12532 13852
rect 12526 13812 12532 13824
rect 12584 13812 12590 13864
rect 12805 13855 12863 13861
rect 12805 13821 12817 13855
rect 12851 13852 12863 13855
rect 13262 13852 13268 13864
rect 12851 13824 13268 13852
rect 12851 13821 12863 13824
rect 12805 13815 12863 13821
rect 13262 13812 13268 13824
rect 13320 13812 13326 13864
rect 13630 13812 13636 13864
rect 13688 13852 13694 13864
rect 14185 13855 14243 13861
rect 14185 13852 14197 13855
rect 13688 13824 14197 13852
rect 13688 13812 13694 13824
rect 14185 13821 14197 13824
rect 14231 13852 14243 13855
rect 14645 13855 14703 13861
rect 14645 13852 14657 13855
rect 14231 13824 14657 13852
rect 14231 13821 14243 13824
rect 14185 13815 14243 13821
rect 14645 13821 14657 13824
rect 14691 13821 14703 13855
rect 15286 13852 15292 13864
rect 15247 13824 15292 13852
rect 14645 13815 14703 13821
rect 15286 13812 15292 13824
rect 15344 13812 15350 13864
rect 15672 13861 15700 13892
rect 17313 13889 17325 13923
rect 17359 13920 17371 13923
rect 21174 13920 21180 13932
rect 17359 13892 19104 13920
rect 21135 13892 21180 13920
rect 17359 13889 17371 13892
rect 17313 13883 17371 13889
rect 15657 13855 15715 13861
rect 15657 13821 15669 13855
rect 15703 13821 15715 13855
rect 15657 13815 15715 13821
rect 16485 13855 16543 13861
rect 16485 13821 16497 13855
rect 16531 13852 16543 13855
rect 16531 13824 16620 13852
rect 16531 13821 16543 13824
rect 16485 13815 16543 13821
rect 11020 13756 11192 13784
rect 16592 13784 16620 13824
rect 16666 13812 16672 13864
rect 16724 13852 16730 13864
rect 16853 13855 16911 13861
rect 16853 13852 16865 13855
rect 16724 13824 16865 13852
rect 16724 13812 16730 13824
rect 16853 13821 16865 13824
rect 16899 13821 16911 13855
rect 16853 13815 16911 13821
rect 17678 13812 17684 13864
rect 17736 13852 17742 13864
rect 18414 13852 18420 13864
rect 17736 13824 18276 13852
rect 18375 13824 18420 13852
rect 17736 13812 17742 13824
rect 16758 13784 16764 13796
rect 16592 13756 16764 13784
rect 11020 13744 11026 13756
rect 16758 13744 16764 13756
rect 16816 13744 16822 13796
rect 18248 13784 18276 13824
rect 18414 13812 18420 13824
rect 18472 13812 18478 13864
rect 18693 13855 18751 13861
rect 18693 13852 18705 13855
rect 18524 13824 18705 13852
rect 18524 13784 18552 13824
rect 18693 13821 18705 13824
rect 18739 13852 18751 13855
rect 18874 13852 18880 13864
rect 18739 13824 18880 13852
rect 18739 13821 18751 13824
rect 18693 13815 18751 13821
rect 18874 13812 18880 13824
rect 18932 13812 18938 13864
rect 18248 13756 18552 13784
rect 8294 13716 8300 13728
rect 7208 13688 8300 13716
rect 8294 13676 8300 13688
rect 8352 13676 8358 13728
rect 9582 13676 9588 13728
rect 9640 13716 9646 13728
rect 14734 13716 14740 13728
rect 9640 13688 14740 13716
rect 9640 13676 9646 13688
rect 14734 13676 14740 13688
rect 14792 13676 14798 13728
rect 19076 13716 19104 13892
rect 21174 13880 21180 13892
rect 21232 13880 21238 13932
rect 19242 13852 19248 13864
rect 19203 13824 19248 13852
rect 19242 13812 19248 13824
rect 19300 13812 19306 13864
rect 19610 13852 19616 13864
rect 19571 13824 19616 13852
rect 19610 13812 19616 13824
rect 19668 13812 19674 13864
rect 20073 13855 20131 13861
rect 20073 13821 20085 13855
rect 20119 13852 20131 13855
rect 20162 13852 20168 13864
rect 20119 13824 20168 13852
rect 20119 13821 20131 13824
rect 20073 13815 20131 13821
rect 20162 13812 20168 13824
rect 20220 13812 20226 13864
rect 20806 13852 20812 13864
rect 20767 13824 20812 13852
rect 20806 13812 20812 13824
rect 20864 13812 20870 13864
rect 21266 13852 21272 13864
rect 21227 13824 21272 13852
rect 21266 13812 21272 13824
rect 21324 13812 21330 13864
rect 21928 13861 21956 13960
rect 22554 13880 22560 13932
rect 22612 13920 22618 13932
rect 23937 13923 23995 13929
rect 23937 13920 23949 13923
rect 22612 13892 23949 13920
rect 22612 13880 22618 13892
rect 23937 13889 23949 13892
rect 23983 13889 23995 13923
rect 26050 13920 26056 13932
rect 26011 13892 26056 13920
rect 23937 13883 23995 13889
rect 26050 13880 26056 13892
rect 26108 13880 26114 13932
rect 26142 13880 26148 13932
rect 26200 13920 26206 13932
rect 29273 13923 29331 13929
rect 29273 13920 29285 13923
rect 26200 13892 29285 13920
rect 26200 13880 26206 13892
rect 29273 13889 29285 13892
rect 29319 13889 29331 13923
rect 29822 13920 29828 13932
rect 29783 13892 29828 13920
rect 29273 13883 29331 13889
rect 29822 13880 29828 13892
rect 29880 13880 29886 13932
rect 21637 13855 21695 13861
rect 21637 13821 21649 13855
rect 21683 13821 21695 13855
rect 21637 13815 21695 13821
rect 21913 13855 21971 13861
rect 21913 13821 21925 13855
rect 21959 13821 21971 13855
rect 21913 13815 21971 13821
rect 19150 13744 19156 13796
rect 19208 13784 19214 13796
rect 19208 13756 20852 13784
rect 19208 13744 19214 13756
rect 19978 13716 19984 13728
rect 19076 13688 19984 13716
rect 19978 13676 19984 13688
rect 20036 13676 20042 13728
rect 20824 13716 20852 13756
rect 20898 13744 20904 13796
rect 20956 13784 20962 13796
rect 21652 13784 21680 13815
rect 20956 13756 21680 13784
rect 21928 13784 21956 13815
rect 22186 13812 22192 13864
rect 22244 13852 22250 13864
rect 22281 13855 22339 13861
rect 22281 13852 22293 13855
rect 22244 13824 22293 13852
rect 22244 13812 22250 13824
rect 22281 13821 22293 13824
rect 22327 13821 22339 13855
rect 23658 13852 23664 13864
rect 23619 13824 23664 13852
rect 22281 13815 22339 13821
rect 23658 13812 23664 13824
rect 23716 13812 23722 13864
rect 25590 13812 25596 13864
rect 25648 13852 25654 13864
rect 25777 13855 25835 13861
rect 25777 13852 25789 13855
rect 25648 13824 25789 13852
rect 25648 13812 25654 13824
rect 25777 13821 25789 13824
rect 25823 13821 25835 13855
rect 28442 13852 28448 13864
rect 28403 13824 28448 13852
rect 25777 13815 25835 13821
rect 28442 13812 28448 13824
rect 28500 13812 28506 13864
rect 29638 13852 29644 13864
rect 29599 13824 29644 13852
rect 29638 13812 29644 13824
rect 29696 13812 29702 13864
rect 29730 13812 29736 13864
rect 29788 13852 29794 13864
rect 29917 13855 29975 13861
rect 29917 13852 29929 13855
rect 29788 13824 29929 13852
rect 29788 13812 29794 13824
rect 29917 13821 29929 13824
rect 29963 13821 29975 13855
rect 30558 13852 30564 13864
rect 30519 13824 30564 13852
rect 29917 13815 29975 13821
rect 22462 13784 22468 13796
rect 21928 13756 22468 13784
rect 20956 13744 20962 13756
rect 21450 13716 21456 13728
rect 20824 13688 21456 13716
rect 21450 13676 21456 13688
rect 21508 13676 21514 13728
rect 21652 13716 21680 13756
rect 22462 13744 22468 13756
rect 22520 13744 22526 13796
rect 29932 13784 29960 13815
rect 30558 13812 30564 13824
rect 30616 13812 30622 13864
rect 30668 13852 30696 13960
rect 31110 13948 31116 13960
rect 31168 13948 31174 14000
rect 32582 13948 32588 14000
rect 32640 13988 32646 14000
rect 35544 13988 35572 14016
rect 32640 13960 35572 13988
rect 32640 13948 32646 13960
rect 33134 13920 33140 13932
rect 33095 13892 33140 13920
rect 33134 13880 33140 13892
rect 33192 13880 33198 13932
rect 30745 13855 30803 13861
rect 30745 13852 30757 13855
rect 30668 13824 30757 13852
rect 30745 13821 30757 13824
rect 30791 13821 30803 13855
rect 31386 13852 31392 13864
rect 31347 13824 31392 13852
rect 30745 13815 30803 13821
rect 31386 13812 31392 13824
rect 31444 13812 31450 13864
rect 31849 13855 31907 13861
rect 31849 13821 31861 13855
rect 31895 13852 31907 13855
rect 31938 13852 31944 13864
rect 31895 13824 31944 13852
rect 31895 13821 31907 13824
rect 31849 13815 31907 13821
rect 31938 13812 31944 13824
rect 31996 13812 32002 13864
rect 32490 13852 32496 13864
rect 32451 13824 32496 13852
rect 32490 13812 32496 13824
rect 32548 13812 32554 13864
rect 33045 13855 33103 13861
rect 33045 13821 33057 13855
rect 33091 13852 33103 13855
rect 33318 13852 33324 13864
rect 33091 13824 33324 13852
rect 33091 13821 33103 13824
rect 33045 13815 33103 13821
rect 33318 13812 33324 13824
rect 33376 13812 33382 13864
rect 33502 13852 33508 13864
rect 33463 13824 33508 13852
rect 33502 13812 33508 13824
rect 33560 13812 33566 13864
rect 33796 13861 33824 13960
rect 35434 13920 35440 13932
rect 35395 13892 35440 13920
rect 35434 13880 35440 13892
rect 35492 13880 35498 13932
rect 33781 13855 33839 13861
rect 33781 13821 33793 13855
rect 33827 13821 33839 13855
rect 33781 13815 33839 13821
rect 33870 13812 33876 13864
rect 33928 13852 33934 13864
rect 34609 13855 34667 13861
rect 34609 13852 34621 13855
rect 33928 13824 34621 13852
rect 33928 13812 33934 13824
rect 34609 13821 34621 13824
rect 34655 13821 34667 13855
rect 35618 13852 35624 13864
rect 35531 13824 35624 13852
rect 34609 13815 34667 13821
rect 35618 13812 35624 13824
rect 35676 13852 35682 13864
rect 35728 13852 35756 14028
rect 37826 14016 37832 14028
rect 37884 14016 37890 14068
rect 38102 13988 38108 14000
rect 36188 13960 38108 13988
rect 36188 13929 36216 13960
rect 38102 13948 38108 13960
rect 38160 13948 38166 14000
rect 36173 13923 36231 13929
rect 36173 13889 36185 13923
rect 36219 13889 36231 13923
rect 36173 13883 36231 13889
rect 37001 13923 37059 13929
rect 37001 13889 37013 13923
rect 37047 13920 37059 13923
rect 38562 13920 38568 13932
rect 37047 13892 38568 13920
rect 37047 13889 37059 13892
rect 37001 13883 37059 13889
rect 38562 13880 38568 13892
rect 38620 13880 38626 13932
rect 35676 13824 35756 13852
rect 35676 13812 35682 13824
rect 36078 13812 36084 13864
rect 36136 13852 36142 13864
rect 36633 13855 36691 13861
rect 36633 13852 36645 13855
rect 36136 13824 36645 13852
rect 36136 13812 36142 13824
rect 36633 13821 36645 13824
rect 36679 13821 36691 13855
rect 37366 13852 37372 13864
rect 37327 13824 37372 13852
rect 36633 13815 36691 13821
rect 37366 13812 37372 13824
rect 37424 13812 37430 13864
rect 37550 13852 37556 13864
rect 37511 13824 37556 13852
rect 37550 13812 37556 13824
rect 37608 13812 37614 13864
rect 37826 13812 37832 13864
rect 37884 13852 37890 13864
rect 37921 13855 37979 13861
rect 37921 13852 37933 13855
rect 37884 13824 37933 13852
rect 37884 13812 37890 13824
rect 37921 13821 37933 13824
rect 37967 13821 37979 13855
rect 37921 13815 37979 13821
rect 38289 13855 38347 13861
rect 38289 13821 38301 13855
rect 38335 13821 38347 13855
rect 38289 13815 38347 13821
rect 34790 13784 34796 13796
rect 29932 13756 34796 13784
rect 34790 13744 34796 13756
rect 34848 13784 34854 13796
rect 35713 13787 35771 13793
rect 35713 13784 35725 13787
rect 34848 13756 35725 13784
rect 34848 13744 34854 13756
rect 35713 13753 35725 13756
rect 35759 13753 35771 13787
rect 35713 13747 35771 13753
rect 35805 13787 35863 13793
rect 35805 13753 35817 13787
rect 35851 13784 35863 13787
rect 36538 13784 36544 13796
rect 35851 13756 36544 13784
rect 35851 13753 35863 13756
rect 35805 13747 35863 13753
rect 36538 13744 36544 13756
rect 36596 13784 36602 13796
rect 37274 13784 37280 13796
rect 36596 13756 37280 13784
rect 36596 13744 36602 13756
rect 37274 13744 37280 13756
rect 37332 13784 37338 13796
rect 37734 13784 37740 13796
rect 37332 13756 37740 13784
rect 37332 13744 37338 13756
rect 37734 13744 37740 13756
rect 37792 13784 37798 13796
rect 38304 13784 38332 13815
rect 37792 13756 38332 13784
rect 37792 13744 37798 13756
rect 22186 13716 22192 13728
rect 21652 13688 22192 13716
rect 22186 13676 22192 13688
rect 22244 13676 22250 13728
rect 24762 13676 24768 13728
rect 24820 13716 24826 13728
rect 27157 13719 27215 13725
rect 27157 13716 27169 13719
rect 24820 13688 27169 13716
rect 24820 13676 24826 13688
rect 27157 13685 27169 13688
rect 27203 13716 27215 13719
rect 27522 13716 27528 13728
rect 27203 13688 27528 13716
rect 27203 13685 27215 13688
rect 27157 13679 27215 13685
rect 27522 13676 27528 13688
rect 27580 13676 27586 13728
rect 31941 13719 31999 13725
rect 31941 13685 31953 13719
rect 31987 13716 31999 13719
rect 32950 13716 32956 13728
rect 31987 13688 32956 13716
rect 31987 13685 31999 13688
rect 31941 13679 31999 13685
rect 32950 13676 32956 13688
rect 33008 13676 33014 13728
rect 33134 13676 33140 13728
rect 33192 13716 33198 13728
rect 33778 13716 33784 13728
rect 33192 13688 33784 13716
rect 33192 13676 33198 13688
rect 33778 13676 33784 13688
rect 33836 13676 33842 13728
rect 34330 13676 34336 13728
rect 34388 13716 34394 13728
rect 34606 13716 34612 13728
rect 34388 13688 34612 13716
rect 34388 13676 34394 13688
rect 34606 13676 34612 13688
rect 34664 13676 34670 13728
rect 1104 13626 39836 13648
rect 1104 13574 19606 13626
rect 19658 13574 19670 13626
rect 19722 13574 19734 13626
rect 19786 13574 19798 13626
rect 19850 13574 39836 13626
rect 1104 13552 39836 13574
rect 1670 13472 1676 13524
rect 1728 13512 1734 13524
rect 7193 13515 7251 13521
rect 7193 13512 7205 13515
rect 1728 13484 7205 13512
rect 1728 13472 1734 13484
rect 7193 13481 7205 13484
rect 7239 13481 7251 13515
rect 15838 13512 15844 13524
rect 7193 13475 7251 13481
rect 11808 13484 15844 13512
rect 2958 13444 2964 13456
rect 1780 13416 2964 13444
rect 1780 13385 1808 13416
rect 2958 13404 2964 13416
rect 3016 13404 3022 13456
rect 3237 13447 3295 13453
rect 3237 13413 3249 13447
rect 3283 13444 3295 13447
rect 5074 13444 5080 13456
rect 3283 13416 5080 13444
rect 3283 13413 3295 13416
rect 3237 13407 3295 13413
rect 5074 13404 5080 13416
rect 5132 13404 5138 13456
rect 11238 13404 11244 13456
rect 11296 13444 11302 13456
rect 11808 13444 11836 13484
rect 15838 13472 15844 13484
rect 15896 13472 15902 13524
rect 16669 13515 16727 13521
rect 16669 13481 16681 13515
rect 16715 13512 16727 13515
rect 16850 13512 16856 13524
rect 16715 13484 16856 13512
rect 16715 13481 16727 13484
rect 16669 13475 16727 13481
rect 16850 13472 16856 13484
rect 16908 13472 16914 13524
rect 18230 13512 18236 13524
rect 18191 13484 18236 13512
rect 18230 13472 18236 13484
rect 18288 13472 18294 13524
rect 18322 13472 18328 13524
rect 18380 13512 18386 13524
rect 19150 13512 19156 13524
rect 18380 13484 19156 13512
rect 18380 13472 18386 13484
rect 19150 13472 19156 13484
rect 19208 13512 19214 13524
rect 19797 13515 19855 13521
rect 19797 13512 19809 13515
rect 19208 13484 19809 13512
rect 19208 13472 19214 13484
rect 19797 13481 19809 13484
rect 19843 13481 19855 13515
rect 19797 13475 19855 13481
rect 21266 13472 21272 13524
rect 21324 13512 21330 13524
rect 21453 13515 21511 13521
rect 21453 13512 21465 13515
rect 21324 13484 21465 13512
rect 21324 13472 21330 13484
rect 21453 13481 21465 13484
rect 21499 13481 21511 13515
rect 21453 13475 21511 13481
rect 23750 13472 23756 13524
rect 23808 13512 23814 13524
rect 24397 13515 24455 13521
rect 24397 13512 24409 13515
rect 23808 13484 24409 13512
rect 23808 13472 23814 13484
rect 24397 13481 24409 13484
rect 24443 13481 24455 13515
rect 28442 13512 28448 13524
rect 24397 13475 24455 13481
rect 24872 13484 28448 13512
rect 11296 13416 11836 13444
rect 11296 13404 11302 13416
rect 1765 13379 1823 13385
rect 1765 13345 1777 13379
rect 1811 13345 1823 13379
rect 1765 13339 1823 13345
rect 2774 13336 2780 13388
rect 2832 13376 2838 13388
rect 2832 13348 2877 13376
rect 2832 13336 2838 13348
rect 3326 13336 3332 13388
rect 3384 13376 3390 13388
rect 4249 13379 4307 13385
rect 4249 13376 4261 13379
rect 3384 13348 4261 13376
rect 3384 13336 3390 13348
rect 4249 13345 4261 13348
rect 4295 13376 4307 13379
rect 4798 13376 4804 13388
rect 4295 13348 4804 13376
rect 4295 13345 4307 13348
rect 4249 13339 4307 13345
rect 4798 13336 4804 13348
rect 4856 13336 4862 13388
rect 7098 13376 7104 13388
rect 7059 13348 7104 13376
rect 7098 13336 7104 13348
rect 7156 13336 7162 13388
rect 7190 13336 7196 13388
rect 7248 13376 7254 13388
rect 7650 13376 7656 13388
rect 7248 13348 7656 13376
rect 7248 13336 7254 13348
rect 7650 13336 7656 13348
rect 7708 13336 7714 13388
rect 8294 13376 8300 13388
rect 8255 13348 8300 13376
rect 8294 13336 8300 13348
rect 8352 13336 8358 13388
rect 8846 13376 8852 13388
rect 8807 13348 8852 13376
rect 8846 13336 8852 13348
rect 8904 13336 8910 13388
rect 9858 13376 9864 13388
rect 9819 13348 9864 13376
rect 9858 13336 9864 13348
rect 9916 13336 9922 13388
rect 10042 13336 10048 13388
rect 10100 13376 10106 13388
rect 10229 13379 10287 13385
rect 10229 13376 10241 13379
rect 10100 13348 10241 13376
rect 10100 13336 10106 13348
rect 10229 13345 10241 13348
rect 10275 13345 10287 13379
rect 11514 13376 11520 13388
rect 11475 13348 11520 13376
rect 10229 13339 10287 13345
rect 11514 13336 11520 13348
rect 11572 13336 11578 13388
rect 11808 13385 11836 13416
rect 12526 13404 12532 13456
rect 12584 13444 12590 13456
rect 24762 13444 24768 13456
rect 12584 13416 18736 13444
rect 12584 13404 12590 13416
rect 11793 13379 11851 13385
rect 11793 13345 11805 13379
rect 11839 13345 11851 13379
rect 11974 13376 11980 13388
rect 11935 13348 11980 13376
rect 11793 13339 11851 13345
rect 11974 13336 11980 13348
rect 12032 13336 12038 13388
rect 12897 13379 12955 13385
rect 12897 13376 12909 13379
rect 12084 13348 12909 13376
rect 1673 13311 1731 13317
rect 1673 13277 1685 13311
rect 1719 13277 1731 13311
rect 2682 13308 2688 13320
rect 2643 13280 2688 13308
rect 1673 13271 1731 13277
rect 1688 13240 1716 13271
rect 2682 13268 2688 13280
rect 2740 13308 2746 13320
rect 4985 13311 5043 13317
rect 2740 13280 4476 13308
rect 2740 13268 2746 13280
rect 3418 13240 3424 13252
rect 1688 13212 3424 13240
rect 3418 13200 3424 13212
rect 3476 13200 3482 13252
rect 4448 13249 4476 13280
rect 4985 13277 4997 13311
rect 5031 13308 5043 13311
rect 5166 13308 5172 13320
rect 5031 13280 5172 13308
rect 5031 13277 5043 13280
rect 4985 13271 5043 13277
rect 5166 13268 5172 13280
rect 5224 13268 5230 13320
rect 5261 13311 5319 13317
rect 5261 13277 5273 13311
rect 5307 13308 5319 13311
rect 9306 13308 9312 13320
rect 5307 13280 9312 13308
rect 5307 13277 5319 13280
rect 5261 13271 5319 13277
rect 9306 13268 9312 13280
rect 9364 13268 9370 13320
rect 10962 13268 10968 13320
rect 11020 13308 11026 13320
rect 12084 13308 12112 13348
rect 12897 13345 12909 13348
rect 12943 13345 12955 13379
rect 13630 13376 13636 13388
rect 13591 13348 13636 13376
rect 12897 13339 12955 13345
rect 13630 13336 13636 13348
rect 13688 13336 13694 13388
rect 13722 13336 13728 13388
rect 13780 13376 13786 13388
rect 14093 13379 14151 13385
rect 14093 13376 14105 13379
rect 13780 13348 14105 13376
rect 13780 13336 13786 13348
rect 14093 13345 14105 13348
rect 14139 13345 14151 13379
rect 15286 13376 15292 13388
rect 15199 13348 15292 13376
rect 14093 13339 14151 13345
rect 15286 13336 15292 13348
rect 15344 13376 15350 13388
rect 15930 13376 15936 13388
rect 15344 13348 15936 13376
rect 15344 13336 15350 13348
rect 15930 13336 15936 13348
rect 15988 13336 15994 13388
rect 16209 13379 16267 13385
rect 16209 13345 16221 13379
rect 16255 13345 16267 13379
rect 16758 13376 16764 13388
rect 16671 13348 16764 13376
rect 16209 13339 16267 13345
rect 12250 13308 12256 13320
rect 11020 13280 12112 13308
rect 12211 13280 12256 13308
rect 11020 13268 11026 13280
rect 12250 13268 12256 13280
rect 12308 13268 12314 13320
rect 4433 13243 4491 13249
rect 4433 13209 4445 13243
rect 4479 13209 4491 13243
rect 4433 13203 4491 13209
rect 9214 13200 9220 13252
rect 9272 13240 9278 13252
rect 15470 13240 15476 13252
rect 9272 13212 15476 13240
rect 9272 13200 9278 13212
rect 15470 13200 15476 13212
rect 15528 13200 15534 13252
rect 1946 13172 1952 13184
rect 1907 13144 1952 13172
rect 1946 13132 1952 13144
rect 2004 13132 2010 13184
rect 6549 13175 6607 13181
rect 6549 13141 6561 13175
rect 6595 13172 6607 13175
rect 6822 13172 6828 13184
rect 6595 13144 6828 13172
rect 6595 13141 6607 13144
rect 6549 13135 6607 13141
rect 6822 13132 6828 13144
rect 6880 13132 6886 13184
rect 7650 13132 7656 13184
rect 7708 13172 7714 13184
rect 8389 13175 8447 13181
rect 8389 13172 8401 13175
rect 7708 13144 8401 13172
rect 7708 13132 7714 13144
rect 8389 13141 8401 13144
rect 8435 13141 8447 13175
rect 8389 13135 8447 13141
rect 9674 13132 9680 13184
rect 9732 13172 9738 13184
rect 9769 13175 9827 13181
rect 9769 13172 9781 13175
rect 9732 13144 9781 13172
rect 9732 13132 9738 13144
rect 9769 13141 9781 13144
rect 9815 13141 9827 13175
rect 9769 13135 9827 13141
rect 10962 13132 10968 13184
rect 11020 13172 11026 13184
rect 12989 13175 13047 13181
rect 12989 13172 13001 13175
rect 11020 13144 13001 13172
rect 11020 13132 11026 13144
rect 12989 13141 13001 13144
rect 13035 13141 13047 13175
rect 12989 13135 13047 13141
rect 13630 13132 13636 13184
rect 13688 13172 13694 13184
rect 14277 13175 14335 13181
rect 14277 13172 14289 13175
rect 13688 13144 14289 13172
rect 13688 13132 13694 13144
rect 14277 13141 14289 13144
rect 14323 13141 14335 13175
rect 14277 13135 14335 13141
rect 14550 13132 14556 13184
rect 14608 13172 14614 13184
rect 15010 13172 15016 13184
rect 14608 13144 15016 13172
rect 14608 13132 14614 13144
rect 15010 13132 15016 13144
rect 15068 13172 15074 13184
rect 16025 13175 16083 13181
rect 16025 13172 16037 13175
rect 15068 13144 16037 13172
rect 15068 13132 15074 13144
rect 16025 13141 16037 13144
rect 16071 13141 16083 13175
rect 16224 13172 16252 13339
rect 16758 13336 16764 13348
rect 16816 13336 16822 13388
rect 17126 13376 17132 13388
rect 17087 13348 17132 13376
rect 17126 13336 17132 13348
rect 17184 13336 17190 13388
rect 17862 13376 17868 13388
rect 17236 13348 17868 13376
rect 16776 13308 16804 13336
rect 17236 13308 17264 13348
rect 17862 13336 17868 13348
rect 17920 13376 17926 13388
rect 18141 13379 18199 13385
rect 18141 13376 18153 13379
rect 17920 13348 18153 13376
rect 17920 13336 17926 13348
rect 18141 13345 18153 13348
rect 18187 13345 18199 13379
rect 18141 13339 18199 13345
rect 18230 13336 18236 13388
rect 18288 13336 18294 13388
rect 18708 13385 18736 13416
rect 19720 13416 24768 13444
rect 19720 13385 19748 13416
rect 18693 13379 18751 13385
rect 18693 13345 18705 13379
rect 18739 13345 18751 13379
rect 18693 13339 18751 13345
rect 19705 13379 19763 13385
rect 19705 13345 19717 13379
rect 19751 13345 19763 13379
rect 21358 13376 21364 13388
rect 21319 13348 21364 13376
rect 19705 13339 19763 13345
rect 21358 13336 21364 13348
rect 21416 13336 21422 13388
rect 21450 13336 21456 13388
rect 21508 13376 21514 13388
rect 22005 13379 22063 13385
rect 22005 13376 22017 13379
rect 21508 13348 22017 13376
rect 21508 13336 21514 13348
rect 22005 13345 22017 13348
rect 22051 13345 22063 13379
rect 22554 13376 22560 13388
rect 22515 13348 22560 13376
rect 22005 13339 22063 13345
rect 22554 13336 22560 13348
rect 22612 13336 22618 13388
rect 24320 13385 24348 13416
rect 24762 13404 24768 13416
rect 24820 13404 24826 13456
rect 24872 13385 24900 13484
rect 28442 13472 28448 13484
rect 28500 13512 28506 13524
rect 28537 13515 28595 13521
rect 28537 13512 28549 13515
rect 28500 13484 28549 13512
rect 28500 13472 28506 13484
rect 28537 13481 28549 13484
rect 28583 13481 28595 13515
rect 33686 13512 33692 13524
rect 28537 13475 28595 13481
rect 30300 13484 32536 13512
rect 33599 13484 33692 13512
rect 24946 13404 24952 13456
rect 25004 13444 25010 13456
rect 25593 13447 25651 13453
rect 25593 13444 25605 13447
rect 25004 13416 25605 13444
rect 25004 13404 25010 13416
rect 25593 13413 25605 13416
rect 25639 13413 25651 13447
rect 30300 13444 30328 13484
rect 30834 13444 30840 13456
rect 25593 13407 25651 13413
rect 28092 13416 29040 13444
rect 23201 13379 23259 13385
rect 23201 13376 23213 13379
rect 22664 13348 23213 13376
rect 16776 13280 17264 13308
rect 17589 13311 17647 13317
rect 17589 13277 17601 13311
rect 17635 13308 17647 13311
rect 18248 13308 18276 13336
rect 17635 13280 18276 13308
rect 17635 13277 17647 13280
rect 17589 13271 17647 13277
rect 18322 13268 18328 13320
rect 18380 13308 18386 13320
rect 18969 13311 19027 13317
rect 18969 13308 18981 13311
rect 18380 13280 18981 13308
rect 18380 13268 18386 13280
rect 18969 13277 18981 13280
rect 19015 13277 19027 13311
rect 18969 13271 19027 13277
rect 19426 13268 19432 13320
rect 19484 13308 19490 13320
rect 22664 13308 22692 13348
rect 23201 13345 23213 13348
rect 23247 13345 23259 13379
rect 23201 13339 23259 13345
rect 24305 13379 24363 13385
rect 24305 13345 24317 13379
rect 24351 13345 24363 13379
rect 24305 13339 24363 13345
rect 24857 13379 24915 13385
rect 24857 13345 24869 13379
rect 24903 13345 24915 13379
rect 24857 13339 24915 13345
rect 25501 13379 25559 13385
rect 25501 13345 25513 13379
rect 25547 13345 25559 13379
rect 25501 13339 25559 13345
rect 19484 13280 22692 13308
rect 22741 13311 22799 13317
rect 19484 13268 19490 13280
rect 22741 13277 22753 13311
rect 22787 13308 22799 13311
rect 23934 13308 23940 13320
rect 22787 13280 23940 13308
rect 22787 13277 22799 13280
rect 22741 13271 22799 13277
rect 23934 13268 23940 13280
rect 23992 13268 23998 13320
rect 20530 13200 20536 13252
rect 20588 13240 20594 13252
rect 25516 13240 25544 13339
rect 26234 13336 26240 13388
rect 26292 13376 26298 13388
rect 26513 13379 26571 13385
rect 26513 13376 26525 13379
rect 26292 13348 26525 13376
rect 26292 13336 26298 13348
rect 26513 13345 26525 13348
rect 26559 13345 26571 13379
rect 27430 13376 27436 13388
rect 27391 13348 27436 13376
rect 26513 13339 26571 13345
rect 27430 13336 27436 13348
rect 27488 13336 27494 13388
rect 26602 13268 26608 13320
rect 26660 13308 26666 13320
rect 27157 13311 27215 13317
rect 27157 13308 27169 13311
rect 26660 13280 27169 13308
rect 26660 13268 26666 13280
rect 27157 13277 27169 13280
rect 27203 13308 27215 13311
rect 28092 13308 28120 13416
rect 27203 13280 28120 13308
rect 29012 13308 29040 13416
rect 29656 13416 30328 13444
rect 30392 13416 30840 13444
rect 29656 13388 29684 13416
rect 29086 13336 29092 13388
rect 29144 13376 29150 13388
rect 29457 13379 29515 13385
rect 29457 13376 29469 13379
rect 29144 13348 29469 13376
rect 29144 13336 29150 13348
rect 29457 13345 29469 13348
rect 29503 13345 29515 13379
rect 29638 13376 29644 13388
rect 29599 13348 29644 13376
rect 29457 13339 29515 13345
rect 29638 13336 29644 13348
rect 29696 13336 29702 13388
rect 30392 13385 30420 13416
rect 30834 13404 30840 13416
rect 30892 13444 30898 13456
rect 32122 13444 32128 13456
rect 30892 13416 32128 13444
rect 30892 13404 30898 13416
rect 32122 13404 32128 13416
rect 32180 13404 32186 13456
rect 30377 13379 30435 13385
rect 30377 13345 30389 13379
rect 30423 13345 30435 13379
rect 30377 13339 30435 13345
rect 30561 13379 30619 13385
rect 30561 13345 30573 13379
rect 30607 13345 30619 13379
rect 30561 13339 30619 13345
rect 30929 13379 30987 13385
rect 30929 13345 30941 13379
rect 30975 13345 30987 13379
rect 30929 13339 30987 13345
rect 29012 13280 29316 13308
rect 27203 13277 27215 13280
rect 27157 13271 27215 13277
rect 29288 13249 29316 13280
rect 29730 13268 29736 13320
rect 29788 13268 29794 13320
rect 30009 13311 30067 13317
rect 30009 13277 30021 13311
rect 30055 13308 30067 13311
rect 30190 13308 30196 13320
rect 30055 13280 30196 13308
rect 30055 13277 30067 13280
rect 30009 13271 30067 13277
rect 30190 13268 30196 13280
rect 30248 13268 30254 13320
rect 30282 13268 30288 13320
rect 30340 13308 30346 13320
rect 30576 13308 30604 13339
rect 30340 13280 30604 13308
rect 30340 13268 30346 13280
rect 20588 13212 25544 13240
rect 29273 13243 29331 13249
rect 20588 13200 20594 13212
rect 29273 13209 29285 13243
rect 29319 13240 29331 13243
rect 29748 13240 29776 13268
rect 30944 13240 30972 13339
rect 31110 13336 31116 13388
rect 31168 13376 31174 13388
rect 31297 13379 31355 13385
rect 31297 13376 31309 13379
rect 31168 13348 31309 13376
rect 31168 13336 31174 13348
rect 31297 13345 31309 13348
rect 31343 13345 31355 13379
rect 31297 13339 31355 13345
rect 32122 13268 32128 13320
rect 32180 13308 32186 13320
rect 32217 13311 32275 13317
rect 32217 13308 32229 13311
rect 32180 13280 32229 13308
rect 32180 13268 32186 13280
rect 32217 13277 32229 13280
rect 32263 13277 32275 13311
rect 32508 13308 32536 13484
rect 33686 13472 33692 13484
rect 33744 13512 33750 13524
rect 33870 13512 33876 13524
rect 33744 13484 33876 13512
rect 33744 13472 33750 13484
rect 33870 13472 33876 13484
rect 33928 13472 33934 13524
rect 34606 13472 34612 13524
rect 34664 13512 34670 13524
rect 36170 13512 36176 13524
rect 34664 13484 36176 13512
rect 34664 13472 34670 13484
rect 36170 13472 36176 13484
rect 36228 13512 36234 13524
rect 36633 13515 36691 13521
rect 36228 13484 36492 13512
rect 36228 13472 36234 13484
rect 32858 13404 32864 13456
rect 32916 13444 32922 13456
rect 32916 13416 33088 13444
rect 32916 13404 32922 13416
rect 32677 13379 32735 13385
rect 32677 13345 32689 13379
rect 32723 13376 32735 13379
rect 32950 13376 32956 13388
rect 32723 13348 32956 13376
rect 32723 13345 32735 13348
rect 32677 13339 32735 13345
rect 32950 13336 32956 13348
rect 33008 13336 33014 13388
rect 33060 13385 33088 13416
rect 33502 13404 33508 13456
rect 33560 13444 33566 13456
rect 33962 13444 33968 13456
rect 33560 13416 33968 13444
rect 33560 13404 33566 13416
rect 33962 13404 33968 13416
rect 34020 13444 34026 13456
rect 34020 13416 35020 13444
rect 34020 13404 34026 13416
rect 33045 13379 33103 13385
rect 33045 13345 33057 13379
rect 33091 13345 33103 13379
rect 33045 13339 33103 13345
rect 33778 13336 33784 13388
rect 33836 13376 33842 13388
rect 33873 13379 33931 13385
rect 33873 13376 33885 13379
rect 33836 13348 33885 13376
rect 33836 13336 33842 13348
rect 33873 13345 33885 13348
rect 33919 13345 33931 13379
rect 33873 13339 33931 13345
rect 34793 13379 34851 13385
rect 34793 13345 34805 13379
rect 34839 13376 34851 13379
rect 34882 13376 34888 13388
rect 34839 13348 34888 13376
rect 34839 13345 34851 13348
rect 34793 13339 34851 13345
rect 34882 13336 34888 13348
rect 34940 13336 34946 13388
rect 34992 13385 35020 13416
rect 34977 13379 35035 13385
rect 34977 13345 34989 13379
rect 35023 13345 35035 13379
rect 35434 13376 35440 13388
rect 35395 13348 35440 13376
rect 34977 13339 35035 13345
rect 35434 13336 35440 13348
rect 35492 13336 35498 13388
rect 35713 13379 35771 13385
rect 35713 13345 35725 13379
rect 35759 13345 35771 13379
rect 36464 13376 36492 13484
rect 36633 13481 36645 13515
rect 36679 13512 36691 13515
rect 37366 13512 37372 13524
rect 36679 13484 37372 13512
rect 36679 13481 36691 13484
rect 36633 13475 36691 13481
rect 37366 13472 37372 13484
rect 37424 13472 37430 13524
rect 36538 13404 36544 13456
rect 36596 13444 36602 13456
rect 36817 13447 36875 13453
rect 36817 13444 36829 13447
rect 36596 13416 36829 13444
rect 36596 13404 36602 13416
rect 36817 13413 36829 13416
rect 36863 13413 36875 13447
rect 37550 13444 37556 13456
rect 36817 13407 36875 13413
rect 36924 13416 37556 13444
rect 36725 13379 36783 13385
rect 36725 13376 36737 13379
rect 36464 13348 36737 13376
rect 35713 13339 35771 13345
rect 36725 13345 36737 13348
rect 36771 13345 36783 13379
rect 36725 13339 36783 13345
rect 34057 13311 34115 13317
rect 34057 13308 34069 13311
rect 32508 13280 34069 13308
rect 32217 13271 32275 13277
rect 34057 13277 34069 13280
rect 34103 13277 34115 13311
rect 34057 13271 34115 13277
rect 34425 13311 34483 13317
rect 34425 13277 34437 13311
rect 34471 13308 34483 13311
rect 34606 13308 34612 13320
rect 34471 13280 34612 13308
rect 34471 13277 34483 13280
rect 34425 13271 34483 13277
rect 29319 13212 29684 13240
rect 29748 13212 30972 13240
rect 29319 13209 29331 13212
rect 29273 13203 29331 13209
rect 21542 13172 21548 13184
rect 16224 13144 21548 13172
rect 16025 13135 16083 13141
rect 21542 13132 21548 13144
rect 21600 13132 21606 13184
rect 22002 13132 22008 13184
rect 22060 13172 22066 13184
rect 23293 13175 23351 13181
rect 23293 13172 23305 13175
rect 22060 13144 23305 13172
rect 22060 13132 22066 13144
rect 23293 13141 23305 13144
rect 23339 13141 23351 13175
rect 23293 13135 23351 13141
rect 26605 13175 26663 13181
rect 26605 13141 26617 13175
rect 26651 13172 26663 13175
rect 28074 13172 28080 13184
rect 26651 13144 28080 13172
rect 26651 13141 26663 13144
rect 26605 13135 26663 13141
rect 28074 13132 28080 13144
rect 28132 13132 28138 13184
rect 29656 13172 29684 13212
rect 30466 13172 30472 13184
rect 29656 13144 30472 13172
rect 30466 13132 30472 13144
rect 30524 13132 30530 13184
rect 32232 13172 32260 13271
rect 32950 13240 32956 13252
rect 32911 13212 32956 13240
rect 32950 13200 32956 13212
rect 33008 13200 33014 13252
rect 34072 13240 34100 13271
rect 34606 13268 34612 13280
rect 34664 13268 34670 13320
rect 35250 13268 35256 13320
rect 35308 13308 35314 13320
rect 35728 13308 35756 13339
rect 35308 13280 35756 13308
rect 35308 13268 35314 13280
rect 36170 13268 36176 13320
rect 36228 13308 36234 13320
rect 36449 13311 36507 13317
rect 36449 13308 36461 13311
rect 36228 13280 36461 13308
rect 36228 13268 36234 13280
rect 36449 13277 36461 13280
rect 36495 13308 36507 13311
rect 36924 13308 36952 13416
rect 37550 13404 37556 13416
rect 37608 13404 37614 13456
rect 37366 13336 37372 13388
rect 37424 13376 37430 13388
rect 37737 13379 37795 13385
rect 37737 13376 37749 13379
rect 37424 13348 37749 13376
rect 37424 13336 37430 13348
rect 37737 13345 37749 13348
rect 37783 13345 37795 13379
rect 38102 13376 38108 13388
rect 38063 13348 38108 13376
rect 37737 13339 37795 13345
rect 38102 13336 38108 13348
rect 38160 13336 38166 13388
rect 38562 13376 38568 13388
rect 38523 13348 38568 13376
rect 38562 13336 38568 13348
rect 38620 13336 38626 13388
rect 37182 13308 37188 13320
rect 36495 13280 36952 13308
rect 37143 13280 37188 13308
rect 36495 13277 36507 13280
rect 36449 13271 36507 13277
rect 37182 13268 37188 13280
rect 37240 13268 37246 13320
rect 36078 13240 36084 13252
rect 34072 13212 36084 13240
rect 36078 13200 36084 13212
rect 36136 13200 36142 13252
rect 38470 13200 38476 13252
rect 38528 13240 38534 13252
rect 38565 13243 38623 13249
rect 38565 13240 38577 13243
rect 38528 13212 38577 13240
rect 38528 13200 38534 13212
rect 38565 13209 38577 13212
rect 38611 13209 38623 13243
rect 38565 13203 38623 13209
rect 35618 13172 35624 13184
rect 32232 13144 35624 13172
rect 35618 13132 35624 13144
rect 35676 13132 35682 13184
rect 1104 13082 39836 13104
rect 1104 13030 4246 13082
rect 4298 13030 4310 13082
rect 4362 13030 4374 13082
rect 4426 13030 4438 13082
rect 4490 13030 34966 13082
rect 35018 13030 35030 13082
rect 35082 13030 35094 13082
rect 35146 13030 35158 13082
rect 35210 13030 39836 13082
rect 1104 13008 39836 13030
rect 2774 12928 2780 12980
rect 2832 12968 2838 12980
rect 5077 12971 5135 12977
rect 2832 12940 2877 12968
rect 2832 12928 2838 12940
rect 5077 12937 5089 12971
rect 5123 12968 5135 12971
rect 5350 12968 5356 12980
rect 5123 12940 5356 12968
rect 5123 12937 5135 12940
rect 5077 12931 5135 12937
rect 5350 12928 5356 12940
rect 5408 12928 5414 12980
rect 5905 12971 5963 12977
rect 5905 12937 5917 12971
rect 5951 12968 5963 12971
rect 5951 12940 15332 12968
rect 5951 12937 5963 12940
rect 5905 12931 5963 12937
rect 8294 12860 8300 12912
rect 8352 12900 8358 12912
rect 9217 12903 9275 12909
rect 9217 12900 9229 12903
rect 8352 12872 9229 12900
rect 8352 12860 8358 12872
rect 9217 12869 9229 12872
rect 9263 12869 9275 12903
rect 9217 12863 9275 12869
rect 9306 12860 9312 12912
rect 9364 12900 9370 12912
rect 14369 12903 14427 12909
rect 14369 12900 14381 12903
rect 9364 12872 14381 12900
rect 9364 12860 9370 12872
rect 14369 12869 14381 12872
rect 14415 12869 14427 12903
rect 14369 12863 14427 12869
rect 1670 12832 1676 12844
rect 1631 12804 1676 12832
rect 1670 12792 1676 12804
rect 1728 12792 1734 12844
rect 2866 12792 2872 12844
rect 2924 12832 2930 12844
rect 5258 12832 5264 12844
rect 2924 12804 5264 12832
rect 2924 12792 2930 12804
rect 5258 12792 5264 12804
rect 5316 12832 5322 12844
rect 5629 12835 5687 12841
rect 5629 12832 5641 12835
rect 5316 12804 5641 12832
rect 5316 12792 5322 12804
rect 5629 12801 5641 12804
rect 5675 12801 5687 12835
rect 5629 12795 5687 12801
rect 6917 12835 6975 12841
rect 6917 12801 6929 12835
rect 6963 12832 6975 12835
rect 9582 12832 9588 12844
rect 6963 12804 9588 12832
rect 6963 12801 6975 12804
rect 6917 12795 6975 12801
rect 9582 12792 9588 12804
rect 9640 12792 9646 12844
rect 11885 12835 11943 12841
rect 9876 12804 11836 12832
rect 1397 12767 1455 12773
rect 1397 12733 1409 12767
rect 1443 12764 1455 12767
rect 3510 12764 3516 12776
rect 1443 12736 3516 12764
rect 1443 12733 1455 12736
rect 1397 12727 1455 12733
rect 3510 12724 3516 12736
rect 3568 12724 3574 12776
rect 3786 12764 3792 12776
rect 3747 12736 3792 12764
rect 3786 12724 3792 12736
rect 3844 12724 3850 12776
rect 5718 12724 5724 12776
rect 5776 12764 5782 12776
rect 6822 12764 6828 12776
rect 5776 12736 5821 12764
rect 6783 12736 6828 12764
rect 5776 12724 5782 12736
rect 6822 12724 6828 12736
rect 6880 12724 6886 12776
rect 7650 12764 7656 12776
rect 7611 12736 7656 12764
rect 7650 12724 7656 12736
rect 7708 12724 7714 12776
rect 7926 12764 7932 12776
rect 7887 12736 7932 12764
rect 7926 12724 7932 12736
rect 7984 12724 7990 12776
rect 8202 12764 8208 12776
rect 8163 12736 8208 12764
rect 8202 12724 8208 12736
rect 8260 12724 8266 12776
rect 8386 12724 8392 12776
rect 8444 12764 8450 12776
rect 9125 12767 9183 12773
rect 9125 12764 9137 12767
rect 8444 12736 9137 12764
rect 8444 12724 8450 12736
rect 9125 12733 9137 12736
rect 9171 12764 9183 12767
rect 9214 12764 9220 12776
rect 9171 12736 9220 12764
rect 9171 12733 9183 12736
rect 9125 12727 9183 12733
rect 9214 12724 9220 12736
rect 9272 12724 9278 12776
rect 9876 12773 9904 12804
rect 9861 12767 9919 12773
rect 9861 12733 9873 12767
rect 9907 12733 9919 12767
rect 10962 12764 10968 12776
rect 10923 12736 10968 12764
rect 9861 12727 9919 12733
rect 10962 12724 10968 12736
rect 11020 12724 11026 12776
rect 11238 12764 11244 12776
rect 11199 12736 11244 12764
rect 11238 12724 11244 12736
rect 11296 12724 11302 12776
rect 11422 12764 11428 12776
rect 11383 12736 11428 12764
rect 11422 12724 11428 12736
rect 11480 12724 11486 12776
rect 11808 12764 11836 12804
rect 11885 12801 11897 12835
rect 11931 12832 11943 12835
rect 15194 12832 15200 12844
rect 11931 12804 13308 12832
rect 11931 12801 11943 12804
rect 11885 12795 11943 12801
rect 12342 12764 12348 12776
rect 11808 12736 12348 12764
rect 12342 12724 12348 12736
rect 12400 12724 12406 12776
rect 12437 12767 12495 12773
rect 12437 12733 12449 12767
rect 12483 12764 12495 12767
rect 12526 12764 12532 12776
rect 12483 12736 12532 12764
rect 12483 12733 12495 12736
rect 12437 12727 12495 12733
rect 12526 12724 12532 12736
rect 12584 12724 12590 12776
rect 12894 12764 12900 12776
rect 12855 12736 12900 12764
rect 12894 12724 12900 12736
rect 12952 12724 12958 12776
rect 13280 12773 13308 12804
rect 14476 12804 15200 12832
rect 14476 12773 14504 12804
rect 15194 12792 15200 12804
rect 15252 12792 15258 12844
rect 15304 12832 15332 12940
rect 15838 12928 15844 12980
rect 15896 12968 15902 12980
rect 16853 12971 16911 12977
rect 16853 12968 16865 12971
rect 15896 12940 16865 12968
rect 15896 12928 15902 12940
rect 16853 12937 16865 12940
rect 16899 12937 16911 12971
rect 18322 12968 18328 12980
rect 18283 12940 18328 12968
rect 16853 12931 16911 12937
rect 18322 12928 18328 12940
rect 18380 12928 18386 12980
rect 19334 12928 19340 12980
rect 19392 12968 19398 12980
rect 19978 12968 19984 12980
rect 19392 12940 19984 12968
rect 19392 12928 19398 12940
rect 19978 12928 19984 12940
rect 20036 12928 20042 12980
rect 20714 12928 20720 12980
rect 20772 12968 20778 12980
rect 26050 12968 26056 12980
rect 20772 12940 26056 12968
rect 20772 12928 20778 12940
rect 26050 12928 26056 12940
rect 26108 12928 26114 12980
rect 30190 12928 30196 12980
rect 30248 12968 30254 12980
rect 31386 12968 31392 12980
rect 30248 12940 31392 12968
rect 30248 12928 30254 12940
rect 31386 12928 31392 12940
rect 31444 12928 31450 12980
rect 32122 12928 32128 12980
rect 32180 12968 32186 12980
rect 32953 12971 33011 12977
rect 32953 12968 32965 12971
rect 32180 12940 32965 12968
rect 32180 12928 32186 12940
rect 32953 12937 32965 12940
rect 32999 12968 33011 12971
rect 33778 12968 33784 12980
rect 32999 12940 33784 12968
rect 32999 12937 33011 12940
rect 32953 12931 33011 12937
rect 33778 12928 33784 12940
rect 33836 12928 33842 12980
rect 36354 12968 36360 12980
rect 36315 12940 36360 12968
rect 36354 12928 36360 12940
rect 36412 12928 36418 12980
rect 36906 12928 36912 12980
rect 36964 12968 36970 12980
rect 37185 12971 37243 12977
rect 37185 12968 37197 12971
rect 36964 12940 37197 12968
rect 36964 12928 36970 12940
rect 37185 12937 37197 12940
rect 37231 12937 37243 12971
rect 37185 12931 37243 12937
rect 16206 12860 16212 12912
rect 16264 12900 16270 12912
rect 16264 12872 20116 12900
rect 16264 12860 16270 12872
rect 17310 12832 17316 12844
rect 15304 12804 17316 12832
rect 17310 12792 17316 12804
rect 17368 12792 17374 12844
rect 19058 12792 19064 12844
rect 19116 12832 19122 12844
rect 19337 12835 19395 12841
rect 19337 12832 19349 12835
rect 19116 12804 19349 12832
rect 19116 12792 19122 12804
rect 19337 12801 19349 12804
rect 19383 12801 19395 12835
rect 19337 12795 19395 12801
rect 13081 12767 13139 12773
rect 13081 12733 13093 12767
rect 13127 12733 13139 12767
rect 13081 12727 13139 12733
rect 13265 12767 13323 12773
rect 13265 12733 13277 12767
rect 13311 12733 13323 12767
rect 13265 12727 13323 12733
rect 14461 12767 14519 12773
rect 14461 12733 14473 12767
rect 14507 12733 14519 12767
rect 14734 12764 14740 12776
rect 14695 12736 14740 12764
rect 14461 12727 14519 12733
rect 8665 12699 8723 12705
rect 8665 12665 8677 12699
rect 8711 12696 8723 12699
rect 13096 12696 13124 12727
rect 14734 12724 14740 12736
rect 14792 12724 14798 12776
rect 15102 12764 15108 12776
rect 15063 12736 15108 12764
rect 15102 12724 15108 12736
rect 15160 12724 15166 12776
rect 15657 12767 15715 12773
rect 15657 12733 15669 12767
rect 15703 12733 15715 12767
rect 16206 12764 16212 12776
rect 16167 12736 16212 12764
rect 15657 12727 15715 12733
rect 8711 12668 13124 12696
rect 15672 12696 15700 12727
rect 16206 12724 16212 12736
rect 16264 12724 16270 12776
rect 16669 12767 16727 12773
rect 16669 12733 16681 12767
rect 16715 12764 16727 12767
rect 18874 12764 18880 12776
rect 16715 12736 16896 12764
rect 18835 12736 18880 12764
rect 16715 12733 16727 12736
rect 16669 12727 16727 12733
rect 16758 12696 16764 12708
rect 15672 12668 16764 12696
rect 8711 12665 8723 12668
rect 8665 12659 8723 12665
rect 16758 12656 16764 12668
rect 16816 12656 16822 12708
rect 13998 12588 14004 12640
rect 14056 12628 14062 12640
rect 16868 12628 16896 12736
rect 18874 12724 18880 12736
rect 18932 12724 18938 12776
rect 18969 12767 19027 12773
rect 18969 12733 18981 12767
rect 19015 12733 19027 12767
rect 18969 12727 19027 12733
rect 19245 12767 19303 12773
rect 19245 12733 19257 12767
rect 19291 12764 19303 12767
rect 19426 12764 19432 12776
rect 19291 12736 19432 12764
rect 19291 12733 19303 12736
rect 19245 12727 19303 12733
rect 18984 12696 19012 12727
rect 19426 12724 19432 12736
rect 19484 12724 19490 12776
rect 19978 12764 19984 12776
rect 19939 12736 19984 12764
rect 19978 12724 19984 12736
rect 20036 12724 20042 12776
rect 19886 12696 19892 12708
rect 18984 12668 19892 12696
rect 19886 12656 19892 12668
rect 19944 12656 19950 12708
rect 14056 12600 16896 12628
rect 14056 12588 14062 12600
rect 19426 12588 19432 12640
rect 19484 12628 19490 12640
rect 19981 12631 20039 12637
rect 19981 12628 19993 12631
rect 19484 12600 19993 12628
rect 19484 12588 19490 12600
rect 19981 12597 19993 12600
rect 20027 12597 20039 12631
rect 20088 12628 20116 12872
rect 25498 12860 25504 12912
rect 25556 12900 25562 12912
rect 25866 12900 25872 12912
rect 25556 12872 25872 12900
rect 25556 12860 25562 12872
rect 25866 12860 25872 12872
rect 25924 12860 25930 12912
rect 27525 12903 27583 12909
rect 27525 12869 27537 12903
rect 27571 12900 27583 12903
rect 27982 12900 27988 12912
rect 27571 12872 27988 12900
rect 27571 12869 27583 12872
rect 27525 12863 27583 12869
rect 27982 12860 27988 12872
rect 28040 12860 28046 12912
rect 30742 12860 30748 12912
rect 30800 12900 30806 12912
rect 31481 12903 31539 12909
rect 31481 12900 31493 12903
rect 30800 12872 31493 12900
rect 30800 12860 30806 12872
rect 31481 12869 31493 12872
rect 31527 12869 31539 12903
rect 31481 12863 31539 12869
rect 33962 12860 33968 12912
rect 34020 12900 34026 12912
rect 34020 12872 35756 12900
rect 34020 12860 34026 12872
rect 23934 12832 23940 12844
rect 20456 12804 23612 12832
rect 23895 12804 23940 12832
rect 20456 12773 20484 12804
rect 20441 12767 20499 12773
rect 20441 12733 20453 12767
rect 20487 12733 20499 12767
rect 21266 12764 21272 12776
rect 21227 12736 21272 12764
rect 20441 12727 20499 12733
rect 21266 12724 21272 12736
rect 21324 12724 21330 12776
rect 21542 12764 21548 12776
rect 21503 12736 21548 12764
rect 21542 12724 21548 12736
rect 21600 12724 21606 12776
rect 23290 12696 23296 12708
rect 22480 12668 23296 12696
rect 22480 12628 22508 12668
rect 23290 12656 23296 12668
rect 23348 12656 23354 12708
rect 22646 12628 22652 12640
rect 20088 12600 22508 12628
rect 22607 12600 22652 12628
rect 19981 12591 20039 12597
rect 22646 12588 22652 12600
rect 22704 12628 22710 12640
rect 23382 12628 23388 12640
rect 22704 12600 23388 12628
rect 22704 12588 22710 12600
rect 23382 12588 23388 12600
rect 23440 12588 23446 12640
rect 23584 12628 23612 12804
rect 23934 12792 23940 12804
rect 23992 12792 23998 12844
rect 27614 12792 27620 12844
rect 27672 12832 27678 12844
rect 28077 12835 28135 12841
rect 28077 12832 28089 12835
rect 27672 12804 28089 12832
rect 27672 12792 27678 12804
rect 28077 12801 28089 12804
rect 28123 12801 28135 12835
rect 28077 12795 28135 12801
rect 29273 12835 29331 12841
rect 29273 12801 29285 12835
rect 29319 12832 29331 12835
rect 30282 12832 30288 12844
rect 29319 12804 30288 12832
rect 29319 12801 29331 12804
rect 29273 12795 29331 12801
rect 30282 12792 30288 12804
rect 30340 12792 30346 12844
rect 30834 12832 30840 12844
rect 30795 12804 30840 12832
rect 30834 12792 30840 12804
rect 30892 12792 30898 12844
rect 33229 12835 33287 12841
rect 33229 12832 33241 12835
rect 32232 12804 33241 12832
rect 32232 12776 32260 12804
rect 33229 12801 33241 12804
rect 33275 12801 33287 12835
rect 33229 12795 33287 12801
rect 33318 12792 33324 12844
rect 33376 12832 33382 12844
rect 33502 12832 33508 12844
rect 33376 12804 33508 12832
rect 33376 12792 33382 12804
rect 33502 12792 33508 12804
rect 33560 12832 33566 12844
rect 33560 12804 34468 12832
rect 33560 12792 33566 12804
rect 23658 12724 23664 12776
rect 23716 12764 23722 12776
rect 24210 12764 24216 12776
rect 23716 12736 24216 12764
rect 23716 12724 23722 12736
rect 24210 12724 24216 12736
rect 24268 12724 24274 12776
rect 25777 12767 25835 12773
rect 25777 12733 25789 12767
rect 25823 12764 25835 12767
rect 25866 12764 25872 12776
rect 25823 12736 25872 12764
rect 25823 12733 25835 12736
rect 25777 12727 25835 12733
rect 25866 12724 25872 12736
rect 25924 12724 25930 12776
rect 26421 12767 26479 12773
rect 26421 12733 26433 12767
rect 26467 12764 26479 12767
rect 26510 12764 26516 12776
rect 26467 12736 26516 12764
rect 26467 12733 26479 12736
rect 26421 12727 26479 12733
rect 26510 12724 26516 12736
rect 26568 12724 26574 12776
rect 26694 12724 26700 12776
rect 26752 12764 26758 12776
rect 27249 12767 27307 12773
rect 27249 12764 27261 12767
rect 26752 12736 27261 12764
rect 26752 12724 26758 12736
rect 27249 12733 27261 12736
rect 27295 12733 27307 12767
rect 27249 12727 27307 12733
rect 27985 12767 28043 12773
rect 27985 12733 27997 12767
rect 28031 12733 28043 12767
rect 27985 12727 28043 12733
rect 28000 12696 28028 12727
rect 28442 12724 28448 12776
rect 28500 12764 28506 12776
rect 29457 12767 29515 12773
rect 28500 12736 29408 12764
rect 28500 12724 28506 12736
rect 28626 12696 28632 12708
rect 28000 12668 28632 12696
rect 28626 12656 28632 12668
rect 28684 12656 28690 12708
rect 29380 12696 29408 12736
rect 29457 12733 29469 12767
rect 29503 12764 29515 12767
rect 29914 12764 29920 12776
rect 29503 12736 29920 12764
rect 29503 12733 29515 12736
rect 29457 12727 29515 12733
rect 29914 12724 29920 12736
rect 29972 12724 29978 12776
rect 31110 12764 31116 12776
rect 31071 12736 31116 12764
rect 31110 12724 31116 12736
rect 31168 12724 31174 12776
rect 31386 12724 31392 12776
rect 31444 12764 31450 12776
rect 31481 12767 31539 12773
rect 31481 12764 31493 12767
rect 31444 12736 31493 12764
rect 31444 12724 31450 12736
rect 31481 12733 31493 12736
rect 31527 12733 31539 12767
rect 32214 12764 32220 12776
rect 32175 12736 32220 12764
rect 31481 12727 31539 12733
rect 32214 12724 32220 12736
rect 32272 12724 32278 12776
rect 33134 12764 33140 12776
rect 33095 12736 33140 12764
rect 33134 12724 33140 12736
rect 33192 12724 33198 12776
rect 33413 12767 33471 12773
rect 33413 12733 33425 12767
rect 33459 12764 33471 12767
rect 34440 12764 34468 12804
rect 34514 12792 34520 12844
rect 34572 12832 34578 12844
rect 34790 12832 34796 12844
rect 34572 12804 34796 12832
rect 34572 12792 34578 12804
rect 34790 12792 34796 12804
rect 34848 12832 34854 12844
rect 34848 12804 35572 12832
rect 34848 12792 34854 12804
rect 35250 12764 35256 12776
rect 33459 12736 34376 12764
rect 34440 12736 35256 12764
rect 33459 12733 33471 12736
rect 33413 12727 33471 12733
rect 29641 12699 29699 12705
rect 29641 12696 29653 12699
rect 29380 12668 29653 12696
rect 29641 12665 29653 12668
rect 29687 12665 29699 12699
rect 29641 12659 29699 12665
rect 30009 12699 30067 12705
rect 30009 12665 30021 12699
rect 30055 12696 30067 12699
rect 31662 12696 31668 12708
rect 30055 12668 31668 12696
rect 30055 12665 30067 12668
rect 30009 12659 30067 12665
rect 31662 12656 31668 12668
rect 31720 12656 31726 12708
rect 24026 12628 24032 12640
rect 23584 12600 24032 12628
rect 24026 12588 24032 12600
rect 24084 12588 24090 12640
rect 25038 12628 25044 12640
rect 24999 12600 25044 12628
rect 25038 12588 25044 12600
rect 25096 12588 25102 12640
rect 25314 12588 25320 12640
rect 25372 12628 25378 12640
rect 26513 12631 26571 12637
rect 26513 12628 26525 12631
rect 25372 12600 26525 12628
rect 25372 12588 25378 12600
rect 26513 12597 26525 12600
rect 26559 12597 26571 12631
rect 26513 12591 26571 12597
rect 27522 12588 27528 12640
rect 27580 12628 27586 12640
rect 29549 12631 29607 12637
rect 29549 12628 29561 12631
rect 27580 12600 29561 12628
rect 27580 12588 27586 12600
rect 29549 12597 29561 12600
rect 29595 12597 29607 12631
rect 29549 12591 29607 12597
rect 30558 12588 30564 12640
rect 30616 12628 30622 12640
rect 32122 12628 32128 12640
rect 30616 12600 32128 12628
rect 30616 12588 30622 12600
rect 32122 12588 32128 12600
rect 32180 12588 32186 12640
rect 32398 12628 32404 12640
rect 32359 12600 32404 12628
rect 32398 12588 32404 12600
rect 32456 12588 32462 12640
rect 33134 12588 33140 12640
rect 33192 12628 33198 12640
rect 33428 12628 33456 12727
rect 33597 12699 33655 12705
rect 33597 12665 33609 12699
rect 33643 12696 33655 12699
rect 33778 12696 33784 12708
rect 33643 12668 33784 12696
rect 33643 12665 33655 12668
rect 33597 12659 33655 12665
rect 33778 12656 33784 12668
rect 33836 12656 33842 12708
rect 33962 12696 33968 12708
rect 33923 12668 33968 12696
rect 33962 12656 33968 12668
rect 34020 12656 34026 12708
rect 34348 12696 34376 12736
rect 35250 12724 35256 12736
rect 35308 12724 35314 12776
rect 35434 12764 35440 12776
rect 35395 12736 35440 12764
rect 35434 12724 35440 12736
rect 35492 12724 35498 12776
rect 34348 12668 34468 12696
rect 34440 12640 34468 12668
rect 33192 12600 33456 12628
rect 33192 12588 33198 12600
rect 33502 12588 33508 12640
rect 33560 12628 33566 12640
rect 33560 12600 33605 12628
rect 33560 12588 33566 12600
rect 34422 12588 34428 12640
rect 34480 12628 34486 12640
rect 35452 12628 35480 12724
rect 35544 12696 35572 12804
rect 35728 12773 35756 12872
rect 38562 12860 38568 12912
rect 38620 12900 38626 12912
rect 38749 12903 38807 12909
rect 38749 12900 38761 12903
rect 38620 12872 38761 12900
rect 38620 12860 38626 12872
rect 38749 12869 38761 12872
rect 38795 12869 38807 12903
rect 38749 12863 38807 12869
rect 36630 12792 36636 12844
rect 36688 12832 36694 12844
rect 36909 12835 36967 12841
rect 36909 12832 36921 12835
rect 36688 12804 36921 12832
rect 36688 12792 36694 12804
rect 36909 12801 36921 12804
rect 36955 12801 36967 12835
rect 36909 12795 36967 12801
rect 37182 12792 37188 12844
rect 37240 12832 37246 12844
rect 37240 12804 38332 12832
rect 37240 12792 37246 12804
rect 35713 12767 35771 12773
rect 35713 12733 35725 12767
rect 35759 12733 35771 12767
rect 35713 12727 35771 12733
rect 36265 12767 36323 12773
rect 36265 12733 36277 12767
rect 36311 12733 36323 12767
rect 36265 12727 36323 12733
rect 36280 12696 36308 12727
rect 36998 12724 37004 12776
rect 37056 12764 37062 12776
rect 37918 12764 37924 12776
rect 37056 12736 37101 12764
rect 37879 12736 37924 12764
rect 37056 12724 37062 12736
rect 37918 12724 37924 12736
rect 37976 12724 37982 12776
rect 38304 12773 38332 12804
rect 38289 12767 38347 12773
rect 38289 12733 38301 12767
rect 38335 12733 38347 12767
rect 38838 12764 38844 12776
rect 38799 12736 38844 12764
rect 38289 12727 38347 12733
rect 38838 12724 38844 12736
rect 38896 12724 38902 12776
rect 35544 12668 36308 12696
rect 34480 12600 35480 12628
rect 34480 12588 34486 12600
rect 1104 12538 39836 12560
rect 1104 12486 19606 12538
rect 19658 12486 19670 12538
rect 19722 12486 19734 12538
rect 19786 12486 19798 12538
rect 19850 12486 39836 12538
rect 1104 12464 39836 12486
rect 12894 12424 12900 12436
rect 11808 12396 12900 12424
rect 3513 12359 3571 12365
rect 3513 12325 3525 12359
rect 3559 12356 3571 12359
rect 3786 12356 3792 12368
rect 3559 12328 3792 12356
rect 3559 12325 3571 12328
rect 3513 12319 3571 12325
rect 3786 12316 3792 12328
rect 3844 12316 3850 12368
rect 8573 12359 8631 12365
rect 8573 12325 8585 12359
rect 8619 12356 8631 12359
rect 8619 12328 10732 12356
rect 8619 12325 8631 12328
rect 8573 12319 8631 12325
rect 2038 12288 2044 12300
rect 1999 12260 2044 12288
rect 2038 12248 2044 12260
rect 2096 12248 2102 12300
rect 2314 12248 2320 12300
rect 2372 12288 2378 12300
rect 2777 12291 2835 12297
rect 2777 12288 2789 12291
rect 2372 12260 2789 12288
rect 2372 12248 2378 12260
rect 2777 12257 2789 12260
rect 2823 12257 2835 12291
rect 2777 12251 2835 12257
rect 3329 12291 3387 12297
rect 3329 12257 3341 12291
rect 3375 12288 3387 12291
rect 6178 12288 6184 12300
rect 3375 12260 6184 12288
rect 3375 12257 3387 12260
rect 3329 12251 3387 12257
rect 6178 12248 6184 12260
rect 6236 12248 6242 12300
rect 7374 12288 7380 12300
rect 7335 12260 7380 12288
rect 7374 12248 7380 12260
rect 7432 12248 7438 12300
rect 7926 12288 7932 12300
rect 7887 12260 7932 12288
rect 7926 12248 7932 12260
rect 7984 12248 7990 12300
rect 8018 12248 8024 12300
rect 8076 12288 8082 12300
rect 8113 12291 8171 12297
rect 8113 12288 8125 12291
rect 8076 12260 8125 12288
rect 8076 12248 8082 12260
rect 8113 12257 8125 12260
rect 8159 12257 8171 12291
rect 10134 12288 10140 12300
rect 10095 12260 10140 12288
rect 8113 12251 8171 12257
rect 10134 12248 10140 12260
rect 10192 12248 10198 12300
rect 10318 12288 10324 12300
rect 10279 12260 10324 12288
rect 10318 12248 10324 12260
rect 10376 12248 10382 12300
rect 10502 12288 10508 12300
rect 10463 12260 10508 12288
rect 10502 12248 10508 12260
rect 10560 12248 10566 12300
rect 5166 12220 5172 12232
rect 5127 12192 5172 12220
rect 5166 12180 5172 12192
rect 5224 12180 5230 12232
rect 5442 12220 5448 12232
rect 5403 12192 5448 12220
rect 5442 12180 5448 12192
rect 5500 12180 5506 12232
rect 10704 12220 10732 12328
rect 11808 12297 11836 12396
rect 12894 12384 12900 12396
rect 12952 12384 12958 12436
rect 17865 12427 17923 12433
rect 17865 12393 17877 12427
rect 17911 12393 17923 12427
rect 17865 12387 17923 12393
rect 18601 12427 18659 12433
rect 18601 12393 18613 12427
rect 18647 12424 18659 12427
rect 19058 12424 19064 12436
rect 18647 12396 19064 12424
rect 18647 12393 18659 12396
rect 18601 12387 18659 12393
rect 12250 12316 12256 12368
rect 12308 12316 12314 12368
rect 15102 12316 15108 12368
rect 15160 12356 15166 12368
rect 16758 12356 16764 12368
rect 15160 12328 16068 12356
rect 16671 12328 16764 12356
rect 15160 12316 15166 12328
rect 11793 12291 11851 12297
rect 11793 12257 11805 12291
rect 11839 12257 11851 12291
rect 11793 12251 11851 12257
rect 11977 12291 12035 12297
rect 11977 12257 11989 12291
rect 12023 12257 12035 12291
rect 11977 12251 12035 12257
rect 12161 12291 12219 12297
rect 12161 12257 12173 12291
rect 12207 12288 12219 12291
rect 12268 12288 12296 12316
rect 12207 12260 12296 12288
rect 12207 12257 12219 12260
rect 12161 12251 12219 12257
rect 11992 12220 12020 12251
rect 12894 12248 12900 12300
rect 12952 12288 12958 12300
rect 13722 12288 13728 12300
rect 12952 12260 13728 12288
rect 12952 12248 12958 12260
rect 13722 12248 13728 12260
rect 13780 12248 13786 12300
rect 15194 12248 15200 12300
rect 15252 12288 15258 12300
rect 16040 12297 16068 12328
rect 16684 12297 16712 12328
rect 16758 12316 16764 12328
rect 16816 12356 16822 12368
rect 17880 12356 17908 12387
rect 19058 12384 19064 12396
rect 19116 12424 19122 12436
rect 22554 12424 22560 12436
rect 19116 12396 20024 12424
rect 19116 12384 19122 12396
rect 18138 12356 18144 12368
rect 16816 12328 17908 12356
rect 17972 12328 18144 12356
rect 16816 12316 16822 12328
rect 15289 12291 15347 12297
rect 15289 12288 15301 12291
rect 15252 12260 15301 12288
rect 15252 12248 15258 12260
rect 15289 12257 15301 12260
rect 15335 12257 15347 12291
rect 15289 12251 15347 12257
rect 15841 12291 15899 12297
rect 15841 12257 15853 12291
rect 15887 12257 15899 12291
rect 15841 12251 15899 12257
rect 16025 12291 16083 12297
rect 16025 12257 16037 12291
rect 16071 12257 16083 12291
rect 16025 12251 16083 12257
rect 16669 12291 16727 12297
rect 16669 12257 16681 12291
rect 16715 12257 16727 12291
rect 16669 12251 16727 12257
rect 10704 12192 12020 12220
rect 13081 12223 13139 12229
rect 13081 12189 13093 12223
rect 13127 12189 13139 12223
rect 13081 12183 13139 12189
rect 13357 12223 13415 12229
rect 13357 12189 13369 12223
rect 13403 12220 13415 12223
rect 15381 12223 15439 12229
rect 15381 12220 15393 12223
rect 13403 12192 15393 12220
rect 13403 12189 13415 12192
rect 13357 12183 13415 12189
rect 15381 12189 15393 12192
rect 15427 12189 15439 12223
rect 15856 12220 15884 12251
rect 16942 12248 16948 12300
rect 17000 12288 17006 12300
rect 17221 12291 17279 12297
rect 17221 12288 17233 12291
rect 17000 12260 17233 12288
rect 17000 12248 17006 12260
rect 17221 12257 17233 12260
rect 17267 12288 17279 12291
rect 17681 12291 17739 12297
rect 17267 12260 17540 12288
rect 17267 12257 17279 12260
rect 17221 12251 17279 12257
rect 15856 12192 16804 12220
rect 15381 12183 15439 12189
rect 9950 12152 9956 12164
rect 9911 12124 9956 12152
rect 9950 12112 9956 12124
rect 10008 12112 10014 12164
rect 11609 12155 11667 12161
rect 11609 12121 11621 12155
rect 11655 12152 11667 12155
rect 11655 12124 12848 12152
rect 11655 12121 11667 12124
rect 11609 12115 11667 12121
rect 2225 12087 2283 12093
rect 2225 12053 2237 12087
rect 2271 12084 2283 12087
rect 2314 12084 2320 12096
rect 2271 12056 2320 12084
rect 2271 12053 2283 12056
rect 2225 12047 2283 12053
rect 2314 12044 2320 12056
rect 2372 12044 2378 12096
rect 6733 12087 6791 12093
rect 6733 12053 6745 12087
rect 6779 12084 6791 12087
rect 6914 12084 6920 12096
rect 6779 12056 6920 12084
rect 6779 12053 6791 12056
rect 6733 12047 6791 12053
rect 6914 12044 6920 12056
rect 6972 12044 6978 12096
rect 12820 12084 12848 12124
rect 12894 12112 12900 12164
rect 12952 12152 12958 12164
rect 13096 12152 13124 12183
rect 16666 12152 16672 12164
rect 12952 12124 13124 12152
rect 14292 12124 16672 12152
rect 12952 12112 12958 12124
rect 14292 12084 14320 12124
rect 16666 12112 16672 12124
rect 16724 12112 16730 12164
rect 14458 12084 14464 12096
rect 12820 12056 14320 12084
rect 14419 12056 14464 12084
rect 14458 12044 14464 12056
rect 14516 12044 14522 12096
rect 14642 12044 14648 12096
rect 14700 12084 14706 12096
rect 16776 12084 16804 12192
rect 17512 12152 17540 12260
rect 17681 12257 17693 12291
rect 17727 12288 17739 12291
rect 17972 12288 18000 12328
rect 18138 12316 18144 12328
rect 18196 12316 18202 12368
rect 19153 12359 19211 12365
rect 19153 12325 19165 12359
rect 19199 12356 19211 12359
rect 19334 12356 19340 12368
rect 19199 12328 19340 12356
rect 19199 12325 19211 12328
rect 19153 12319 19211 12325
rect 19334 12316 19340 12328
rect 19392 12316 19398 12368
rect 18414 12288 18420 12300
rect 17727 12260 18000 12288
rect 18375 12260 18420 12288
rect 17727 12257 17739 12260
rect 17681 12251 17739 12257
rect 18414 12248 18420 12260
rect 18472 12248 18478 12300
rect 19242 12248 19248 12300
rect 19300 12288 19306 12300
rect 19797 12291 19855 12297
rect 19797 12288 19809 12291
rect 19300 12260 19809 12288
rect 19300 12248 19306 12260
rect 19797 12257 19809 12260
rect 19843 12257 19855 12291
rect 19797 12251 19855 12257
rect 19886 12220 19892 12232
rect 19847 12192 19892 12220
rect 19886 12180 19892 12192
rect 19944 12180 19950 12232
rect 19996 12220 20024 12396
rect 22112 12396 22560 12424
rect 21358 12356 21364 12368
rect 20180 12328 21364 12356
rect 20180 12297 20208 12328
rect 21358 12316 21364 12328
rect 21416 12316 21422 12368
rect 20165 12291 20223 12297
rect 20165 12257 20177 12291
rect 20211 12257 20223 12291
rect 20349 12291 20407 12297
rect 20349 12288 20361 12291
rect 20165 12251 20223 12257
rect 20272 12260 20361 12288
rect 20272 12220 20300 12260
rect 20349 12257 20361 12260
rect 20395 12288 20407 12291
rect 20714 12288 20720 12300
rect 20395 12260 20720 12288
rect 20395 12257 20407 12260
rect 20349 12251 20407 12257
rect 20714 12248 20720 12260
rect 20772 12248 20778 12300
rect 20806 12248 20812 12300
rect 20864 12288 20870 12300
rect 21269 12291 21327 12297
rect 21269 12288 21281 12291
rect 20864 12260 21281 12288
rect 20864 12248 20870 12260
rect 21269 12257 21281 12260
rect 21315 12257 21327 12291
rect 21269 12251 21327 12257
rect 21913 12291 21971 12297
rect 21913 12257 21925 12291
rect 21959 12288 21971 12291
rect 22112 12288 22140 12396
rect 22554 12384 22560 12396
rect 22612 12424 22618 12436
rect 23753 12427 23811 12433
rect 23753 12424 23765 12427
rect 22612 12396 23765 12424
rect 22612 12384 22618 12396
rect 23753 12393 23765 12396
rect 23799 12393 23811 12427
rect 25314 12424 25320 12436
rect 23753 12387 23811 12393
rect 23860 12396 25320 12424
rect 22462 12316 22468 12368
rect 22520 12356 22526 12368
rect 23860 12356 23888 12396
rect 25314 12384 25320 12396
rect 25372 12384 25378 12436
rect 26050 12384 26056 12436
rect 26108 12424 26114 12436
rect 26605 12427 26663 12433
rect 26605 12424 26617 12427
rect 26108 12396 26617 12424
rect 26108 12384 26114 12396
rect 26605 12393 26617 12396
rect 26651 12393 26663 12427
rect 28718 12424 28724 12436
rect 28679 12396 28724 12424
rect 26605 12387 26663 12393
rect 28718 12384 28724 12396
rect 28776 12384 28782 12436
rect 29457 12427 29515 12433
rect 29457 12393 29469 12427
rect 29503 12424 29515 12427
rect 29730 12424 29736 12436
rect 29503 12396 29736 12424
rect 29503 12393 29515 12396
rect 29457 12387 29515 12393
rect 29730 12384 29736 12396
rect 29788 12384 29794 12436
rect 31386 12384 31392 12436
rect 31444 12424 31450 12436
rect 32125 12427 32183 12433
rect 32125 12424 32137 12427
rect 31444 12396 32137 12424
rect 31444 12384 31450 12396
rect 32125 12393 32137 12396
rect 32171 12393 32183 12427
rect 32125 12387 32183 12393
rect 33137 12427 33195 12433
rect 33137 12393 33149 12427
rect 33183 12424 33195 12427
rect 33778 12424 33784 12436
rect 33183 12396 33784 12424
rect 33183 12393 33195 12396
rect 33137 12387 33195 12393
rect 33778 12384 33784 12396
rect 33836 12424 33842 12436
rect 34330 12424 34336 12436
rect 33836 12396 34336 12424
rect 33836 12384 33842 12396
rect 34330 12384 34336 12396
rect 34388 12384 34394 12436
rect 34422 12384 34428 12436
rect 34480 12424 34486 12436
rect 38930 12424 38936 12436
rect 34480 12396 38936 12424
rect 34480 12384 34486 12396
rect 38930 12384 38936 12396
rect 38988 12384 38994 12436
rect 24946 12356 24952 12368
rect 22520 12328 23888 12356
rect 24688 12328 24952 12356
rect 22520 12316 22526 12328
rect 22278 12288 22284 12300
rect 21959 12260 22140 12288
rect 22239 12260 22284 12288
rect 21959 12257 21971 12260
rect 21913 12251 21971 12257
rect 22278 12248 22284 12260
rect 22336 12248 22342 12300
rect 22664 12297 22692 12328
rect 22649 12291 22707 12297
rect 22649 12257 22661 12291
rect 22695 12257 22707 12291
rect 22649 12251 22707 12257
rect 23201 12291 23259 12297
rect 23201 12257 23213 12291
rect 23247 12257 23259 12291
rect 23201 12251 23259 12257
rect 23216 12220 23244 12251
rect 23382 12248 23388 12300
rect 23440 12288 23446 12300
rect 24688 12297 24716 12328
rect 24946 12316 24952 12328
rect 25004 12316 25010 12368
rect 25225 12359 25283 12365
rect 25225 12325 25237 12359
rect 25271 12356 25283 12359
rect 30098 12356 30104 12368
rect 25271 12328 30104 12356
rect 25271 12325 25283 12328
rect 25225 12319 25283 12325
rect 30098 12316 30104 12328
rect 30156 12316 30162 12368
rect 30558 12356 30564 12368
rect 30208 12328 30564 12356
rect 23661 12291 23719 12297
rect 23661 12288 23673 12291
rect 23440 12260 23673 12288
rect 23440 12248 23446 12260
rect 23661 12257 23673 12260
rect 23707 12257 23719 12291
rect 23661 12251 23719 12257
rect 24673 12291 24731 12297
rect 24673 12257 24685 12291
rect 24719 12257 24731 12291
rect 24673 12251 24731 12257
rect 24765 12291 24823 12297
rect 24765 12257 24777 12291
rect 24811 12288 24823 12291
rect 25038 12288 25044 12300
rect 24811 12260 25044 12288
rect 24811 12257 24823 12260
rect 24765 12251 24823 12257
rect 25038 12248 25044 12260
rect 25096 12248 25102 12300
rect 25685 12291 25743 12297
rect 25685 12257 25697 12291
rect 25731 12288 25743 12291
rect 26050 12288 26056 12300
rect 25731 12260 26056 12288
rect 25731 12257 25743 12260
rect 25685 12251 25743 12257
rect 26050 12248 26056 12260
rect 26108 12248 26114 12300
rect 26510 12288 26516 12300
rect 26471 12260 26516 12288
rect 26510 12248 26516 12260
rect 26568 12248 26574 12300
rect 27154 12288 27160 12300
rect 27115 12260 27160 12288
rect 27154 12248 27160 12260
rect 27212 12248 27218 12300
rect 27522 12248 27528 12300
rect 27580 12288 27586 12300
rect 30208 12297 30236 12328
rect 30558 12316 30564 12328
rect 30616 12316 30622 12368
rect 30926 12316 30932 12368
rect 30984 12356 30990 12368
rect 32674 12356 32680 12368
rect 30984 12328 32680 12356
rect 30984 12316 30990 12328
rect 32674 12316 32680 12328
rect 32732 12316 32738 12368
rect 36265 12359 36323 12365
rect 36265 12356 36277 12359
rect 35728 12328 36277 12356
rect 27801 12291 27859 12297
rect 27801 12288 27813 12291
rect 27580 12260 27813 12288
rect 27580 12248 27586 12260
rect 27801 12257 27813 12260
rect 27847 12288 27859 12291
rect 28537 12291 28595 12297
rect 28537 12288 28549 12291
rect 27847 12260 28549 12288
rect 27847 12257 27859 12260
rect 27801 12251 27859 12257
rect 28537 12257 28549 12260
rect 28583 12257 28595 12291
rect 28537 12251 28595 12257
rect 29273 12291 29331 12297
rect 29273 12257 29285 12291
rect 29319 12257 29331 12291
rect 29273 12251 29331 12257
rect 30193 12291 30251 12297
rect 30193 12257 30205 12291
rect 30239 12257 30251 12291
rect 30650 12288 30656 12300
rect 30611 12260 30656 12288
rect 30193 12251 30251 12257
rect 25777 12223 25835 12229
rect 25777 12220 25789 12223
rect 19996 12192 20300 12220
rect 20364 12192 25789 12220
rect 20364 12152 20392 12192
rect 25777 12189 25789 12192
rect 25823 12189 25835 12223
rect 29288 12220 29316 12251
rect 30650 12248 30656 12260
rect 30708 12248 30714 12300
rect 30742 12248 30748 12300
rect 30800 12288 30806 12300
rect 31021 12291 31079 12297
rect 31021 12288 31033 12291
rect 30800 12260 31033 12288
rect 30800 12248 30806 12260
rect 31021 12257 31033 12260
rect 31067 12257 31079 12291
rect 31021 12251 31079 12257
rect 31662 12248 31668 12300
rect 31720 12288 31726 12300
rect 32217 12291 32275 12297
rect 32217 12288 32229 12291
rect 31720 12260 32229 12288
rect 31720 12248 31726 12260
rect 32217 12257 32229 12260
rect 32263 12257 32275 12291
rect 32217 12251 32275 12257
rect 32490 12248 32496 12300
rect 32548 12288 32554 12300
rect 32953 12291 33011 12297
rect 32953 12288 32965 12291
rect 32548 12260 32965 12288
rect 32548 12248 32554 12260
rect 32953 12257 32965 12260
rect 32999 12257 33011 12291
rect 32953 12251 33011 12257
rect 33962 12248 33968 12300
rect 34020 12288 34026 12300
rect 34149 12291 34207 12297
rect 34149 12288 34161 12291
rect 34020 12260 34161 12288
rect 34020 12248 34026 12260
rect 34149 12257 34161 12260
rect 34195 12257 34207 12291
rect 34606 12288 34612 12300
rect 34567 12260 34612 12288
rect 34149 12251 34207 12257
rect 34606 12248 34612 12260
rect 34664 12248 34670 12300
rect 35728 12288 35756 12328
rect 36265 12325 36277 12328
rect 36311 12325 36323 12359
rect 36265 12319 36323 12325
rect 36633 12359 36691 12365
rect 36633 12325 36645 12359
rect 36679 12356 36691 12359
rect 37274 12356 37280 12368
rect 36679 12328 37280 12356
rect 36679 12325 36691 12328
rect 36633 12319 36691 12325
rect 37274 12316 37280 12328
rect 37332 12316 37338 12368
rect 36078 12288 36084 12300
rect 34808 12260 35756 12288
rect 36039 12260 36084 12288
rect 34808 12232 34836 12260
rect 36078 12248 36084 12260
rect 36136 12248 36142 12300
rect 36173 12291 36231 12297
rect 36173 12257 36185 12291
rect 36219 12288 36231 12291
rect 37826 12288 37832 12300
rect 36219 12260 37832 12288
rect 36219 12257 36231 12260
rect 36173 12251 36231 12257
rect 25777 12183 25835 12189
rect 28000 12192 29316 12220
rect 29380 12192 30880 12220
rect 17512 12124 20392 12152
rect 20622 12112 20628 12164
rect 20680 12152 20686 12164
rect 21358 12152 21364 12164
rect 20680 12124 21364 12152
rect 20680 12112 20686 12124
rect 21358 12112 21364 12124
rect 21416 12112 21422 12164
rect 21542 12152 21548 12164
rect 21503 12124 21548 12152
rect 21542 12112 21548 12124
rect 21600 12112 21606 12164
rect 23474 12112 23480 12164
rect 23532 12152 23538 12164
rect 28000 12161 28028 12192
rect 27985 12155 28043 12161
rect 27985 12152 27997 12155
rect 23532 12124 27997 12152
rect 23532 12112 23538 12124
rect 27985 12121 27997 12124
rect 28031 12121 28043 12155
rect 29380 12152 29408 12192
rect 30742 12152 30748 12164
rect 27985 12115 28043 12121
rect 28092 12124 29408 12152
rect 30703 12124 30748 12152
rect 17678 12084 17684 12096
rect 14700 12056 17684 12084
rect 14700 12044 14706 12056
rect 17678 12044 17684 12056
rect 17736 12044 17742 12096
rect 17770 12044 17776 12096
rect 17828 12084 17834 12096
rect 21634 12084 21640 12096
rect 17828 12056 21640 12084
rect 17828 12044 17834 12056
rect 21634 12044 21640 12056
rect 21692 12044 21698 12096
rect 23382 12044 23388 12096
rect 23440 12084 23446 12096
rect 24946 12084 24952 12096
rect 23440 12056 24952 12084
rect 23440 12044 23446 12056
rect 24946 12044 24952 12056
rect 25004 12084 25010 12096
rect 27249 12087 27307 12093
rect 27249 12084 27261 12087
rect 25004 12056 27261 12084
rect 25004 12044 25010 12056
rect 27249 12053 27261 12056
rect 27295 12084 27307 12087
rect 28092 12084 28120 12124
rect 30742 12112 30748 12124
rect 30800 12112 30806 12164
rect 30852 12152 30880 12192
rect 31386 12180 31392 12232
rect 31444 12220 31450 12232
rect 33873 12223 33931 12229
rect 31444 12192 31489 12220
rect 31444 12180 31450 12192
rect 33873 12189 33885 12223
rect 33919 12189 33931 12223
rect 33873 12183 33931 12189
rect 31662 12152 31668 12164
rect 30852 12124 31668 12152
rect 31662 12112 31668 12124
rect 31720 12112 31726 12164
rect 32125 12155 32183 12161
rect 32125 12121 32137 12155
rect 32171 12152 32183 12155
rect 33778 12152 33784 12164
rect 32171 12124 33784 12152
rect 32171 12121 32183 12124
rect 32125 12115 32183 12121
rect 33778 12112 33784 12124
rect 33836 12112 33842 12164
rect 27295 12056 28120 12084
rect 27295 12053 27307 12056
rect 27249 12047 27307 12053
rect 29086 12044 29092 12096
rect 29144 12084 29150 12096
rect 30009 12087 30067 12093
rect 30009 12084 30021 12087
rect 29144 12056 30021 12084
rect 29144 12044 29150 12056
rect 30009 12053 30021 12056
rect 30055 12053 30067 12087
rect 30009 12047 30067 12053
rect 30190 12044 30196 12096
rect 30248 12084 30254 12096
rect 32401 12087 32459 12093
rect 32401 12084 32413 12087
rect 30248 12056 32413 12084
rect 30248 12044 30254 12056
rect 32401 12053 32413 12056
rect 32447 12084 32459 12087
rect 33502 12084 33508 12096
rect 32447 12056 33508 12084
rect 32447 12053 32459 12056
rect 32401 12047 32459 12053
rect 33502 12044 33508 12056
rect 33560 12044 33566 12096
rect 33888 12084 33916 12183
rect 34422 12180 34428 12232
rect 34480 12220 34486 12232
rect 34790 12220 34796 12232
rect 34480 12192 34796 12220
rect 34480 12180 34486 12192
rect 34790 12180 34796 12192
rect 34848 12180 34854 12232
rect 35897 12223 35955 12229
rect 35897 12189 35909 12223
rect 35943 12220 35955 12223
rect 35986 12220 35992 12232
rect 35943 12192 35992 12220
rect 35943 12189 35955 12192
rect 35897 12183 35955 12189
rect 35986 12180 35992 12192
rect 36044 12220 36050 12232
rect 36446 12220 36452 12232
rect 36044 12192 36452 12220
rect 36044 12180 36050 12192
rect 36446 12180 36452 12192
rect 36504 12180 36510 12232
rect 33962 12112 33968 12164
rect 34020 12152 34026 12164
rect 34609 12155 34667 12161
rect 34609 12152 34621 12155
rect 34020 12124 34621 12152
rect 34020 12112 34026 12124
rect 34609 12121 34621 12124
rect 34655 12121 34667 12155
rect 34609 12115 34667 12121
rect 34514 12084 34520 12096
rect 33888 12056 34520 12084
rect 34514 12044 34520 12056
rect 34572 12044 34578 12096
rect 35342 12044 35348 12096
rect 35400 12084 35406 12096
rect 36556 12084 36584 12260
rect 37826 12248 37832 12260
rect 37884 12248 37890 12300
rect 38105 12291 38163 12297
rect 38105 12257 38117 12291
rect 38151 12288 38163 12291
rect 38194 12288 38200 12300
rect 38151 12260 38200 12288
rect 38151 12257 38163 12260
rect 38105 12251 38163 12257
rect 38194 12248 38200 12260
rect 38252 12248 38258 12300
rect 38562 12288 38568 12300
rect 38523 12260 38568 12288
rect 38562 12248 38568 12260
rect 38620 12248 38626 12300
rect 38746 12220 38752 12232
rect 38707 12192 38752 12220
rect 38746 12180 38752 12192
rect 38804 12180 38810 12232
rect 37734 12112 37740 12164
rect 37792 12152 37798 12164
rect 38013 12155 38071 12161
rect 38013 12152 38025 12155
rect 37792 12124 38025 12152
rect 37792 12112 37798 12124
rect 38013 12121 38025 12124
rect 38059 12121 38071 12155
rect 38013 12115 38071 12121
rect 35400 12056 36584 12084
rect 35400 12044 35406 12056
rect 1104 11994 39836 12016
rect 1104 11942 4246 11994
rect 4298 11942 4310 11994
rect 4362 11942 4374 11994
rect 4426 11942 4438 11994
rect 4490 11942 34966 11994
rect 35018 11942 35030 11994
rect 35082 11942 35094 11994
rect 35146 11942 35158 11994
rect 35210 11942 39836 11994
rect 1104 11920 39836 11942
rect 4617 11883 4675 11889
rect 4617 11849 4629 11883
rect 4663 11880 4675 11883
rect 5718 11880 5724 11892
rect 4663 11852 5724 11880
rect 4663 11849 4675 11852
rect 4617 11843 4675 11849
rect 5718 11840 5724 11852
rect 5776 11840 5782 11892
rect 6178 11880 6184 11892
rect 6139 11852 6184 11880
rect 6178 11840 6184 11852
rect 6236 11840 6242 11892
rect 7190 11880 7196 11892
rect 7151 11852 7196 11880
rect 7190 11840 7196 11852
rect 7248 11840 7254 11892
rect 12342 11840 12348 11892
rect 12400 11880 12406 11892
rect 14458 11880 14464 11892
rect 12400 11852 14464 11880
rect 12400 11840 12406 11852
rect 14458 11840 14464 11852
rect 14516 11840 14522 11892
rect 15562 11840 15568 11892
rect 15620 11880 15626 11892
rect 15620 11852 17908 11880
rect 15620 11840 15626 11852
rect 10134 11772 10140 11824
rect 10192 11812 10198 11824
rect 12710 11812 12716 11824
rect 10192 11784 12388 11812
rect 12671 11784 12716 11812
rect 10192 11772 10198 11784
rect 3053 11747 3111 11753
rect 3053 11713 3065 11747
rect 3099 11744 3111 11747
rect 3510 11744 3516 11756
rect 3099 11716 3516 11744
rect 3099 11713 3111 11716
rect 3053 11707 3111 11713
rect 3510 11704 3516 11716
rect 3568 11704 3574 11756
rect 8294 11744 8300 11756
rect 8036 11716 8300 11744
rect 3326 11676 3332 11688
rect 3287 11648 3332 11676
rect 3326 11636 3332 11648
rect 3384 11636 3390 11688
rect 6089 11679 6147 11685
rect 6089 11645 6101 11679
rect 6135 11676 6147 11679
rect 6914 11676 6920 11688
rect 6135 11648 6920 11676
rect 6135 11645 6147 11648
rect 6089 11639 6147 11645
rect 6914 11636 6920 11648
rect 6972 11636 6978 11688
rect 7101 11679 7159 11685
rect 7101 11645 7113 11679
rect 7147 11676 7159 11679
rect 7558 11676 7564 11688
rect 7147 11648 7564 11676
rect 7147 11645 7159 11648
rect 7101 11639 7159 11645
rect 7558 11636 7564 11648
rect 7616 11636 7622 11688
rect 8036 11685 8064 11716
rect 8294 11704 8300 11716
rect 8352 11704 8358 11756
rect 8941 11747 8999 11753
rect 8941 11713 8953 11747
rect 8987 11744 8999 11747
rect 10318 11744 10324 11756
rect 8987 11716 10324 11744
rect 8987 11713 8999 11716
rect 8941 11707 8999 11713
rect 10318 11704 10324 11716
rect 10376 11704 10382 11756
rect 10502 11744 10508 11756
rect 10463 11716 10508 11744
rect 10502 11704 10508 11716
rect 10560 11704 10566 11756
rect 11422 11744 11428 11756
rect 11383 11716 11428 11744
rect 11422 11704 11428 11716
rect 11480 11704 11486 11756
rect 12360 11744 12388 11784
rect 12710 11772 12716 11784
rect 12768 11772 12774 11824
rect 14366 11772 14372 11824
rect 14424 11812 14430 11824
rect 14645 11815 14703 11821
rect 14645 11812 14657 11815
rect 14424 11784 14657 11812
rect 14424 11772 14430 11784
rect 14645 11781 14657 11784
rect 14691 11781 14703 11815
rect 17770 11812 17776 11824
rect 14645 11775 14703 11781
rect 14752 11784 17776 11812
rect 12360 11716 12940 11744
rect 8021 11679 8079 11685
rect 8021 11645 8033 11679
rect 8067 11645 8079 11679
rect 8021 11639 8079 11645
rect 8205 11679 8263 11685
rect 8205 11645 8217 11679
rect 8251 11645 8263 11679
rect 8478 11676 8484 11688
rect 8439 11648 8484 11676
rect 8205 11639 8263 11645
rect 7926 11568 7932 11620
rect 7984 11608 7990 11620
rect 8220 11608 8248 11639
rect 8478 11636 8484 11648
rect 8536 11636 8542 11688
rect 9585 11679 9643 11685
rect 9585 11645 9597 11679
rect 9631 11676 9643 11679
rect 9674 11676 9680 11688
rect 9631 11648 9680 11676
rect 9631 11645 9643 11648
rect 9585 11639 9643 11645
rect 9674 11636 9680 11648
rect 9732 11636 9738 11688
rect 9861 11679 9919 11685
rect 9861 11645 9873 11679
rect 9907 11645 9919 11679
rect 9861 11639 9919 11645
rect 7984 11580 8248 11608
rect 7984 11568 7990 11580
rect 8220 11540 8248 11580
rect 9674 11540 9680 11552
rect 8220 11512 9680 11540
rect 9674 11500 9680 11512
rect 9732 11500 9738 11552
rect 9876 11540 9904 11639
rect 10042 11636 10048 11688
rect 10100 11676 10106 11688
rect 10137 11679 10195 11685
rect 10137 11676 10149 11679
rect 10100 11648 10149 11676
rect 10100 11636 10106 11648
rect 10137 11645 10149 11648
rect 10183 11645 10195 11679
rect 11330 11676 11336 11688
rect 11291 11648 11336 11676
rect 10137 11639 10195 11645
rect 11330 11636 11336 11648
rect 11388 11636 11394 11688
rect 11698 11676 11704 11688
rect 11659 11648 11704 11676
rect 11698 11636 11704 11648
rect 11756 11636 11762 11688
rect 12912 11685 12940 11716
rect 13538 11704 13544 11756
rect 13596 11744 13602 11756
rect 14752 11744 14780 11784
rect 17770 11772 17776 11784
rect 17828 11772 17834 11824
rect 17880 11812 17908 11852
rect 18230 11840 18236 11892
rect 18288 11880 18294 11892
rect 19797 11883 19855 11889
rect 19797 11880 19809 11883
rect 18288 11852 19809 11880
rect 18288 11840 18294 11852
rect 19797 11849 19809 11852
rect 19843 11849 19855 11883
rect 19797 11843 19855 11849
rect 19886 11840 19892 11892
rect 19944 11880 19950 11892
rect 21453 11883 21511 11889
rect 21453 11880 21465 11883
rect 19944 11852 21465 11880
rect 19944 11840 19950 11852
rect 21453 11849 21465 11852
rect 21499 11849 21511 11883
rect 21453 11843 21511 11849
rect 21634 11840 21640 11892
rect 21692 11880 21698 11892
rect 23474 11880 23480 11892
rect 21692 11852 23480 11880
rect 21692 11840 21698 11852
rect 23474 11840 23480 11852
rect 23532 11840 23538 11892
rect 23750 11880 23756 11892
rect 23711 11852 23756 11880
rect 23750 11840 23756 11852
rect 23808 11840 23814 11892
rect 23934 11840 23940 11892
rect 23992 11880 23998 11892
rect 24210 11880 24216 11892
rect 23992 11852 24216 11880
rect 23992 11840 23998 11852
rect 24210 11840 24216 11852
rect 24268 11840 24274 11892
rect 26326 11880 26332 11892
rect 24412 11852 26332 11880
rect 23382 11812 23388 11824
rect 17880 11784 18552 11812
rect 13596 11716 14780 11744
rect 13596 11704 13602 11716
rect 12897 11679 12955 11685
rect 12897 11645 12909 11679
rect 12943 11645 12955 11679
rect 13078 11676 13084 11688
rect 13039 11648 13084 11676
rect 12897 11639 12955 11645
rect 12912 11608 12940 11639
rect 13078 11636 13084 11648
rect 13136 11636 13142 11688
rect 13262 11676 13268 11688
rect 13223 11648 13268 11676
rect 13262 11636 13268 11648
rect 13320 11636 13326 11688
rect 14752 11685 14780 11716
rect 15565 11747 15623 11753
rect 15565 11713 15577 11747
rect 15611 11744 15623 11747
rect 17862 11744 17868 11756
rect 15611 11716 17868 11744
rect 15611 11713 15623 11716
rect 15565 11707 15623 11713
rect 17862 11704 17868 11716
rect 17920 11704 17926 11756
rect 18524 11688 18552 11784
rect 19076 11784 23388 11812
rect 13909 11679 13967 11685
rect 13909 11645 13921 11679
rect 13955 11676 13967 11679
rect 14737 11679 14795 11685
rect 13955 11648 14688 11676
rect 13955 11645 13967 11648
rect 13909 11639 13967 11645
rect 13630 11608 13636 11620
rect 12912 11580 13636 11608
rect 13630 11568 13636 11580
rect 13688 11568 13694 11620
rect 9950 11540 9956 11552
rect 9863 11512 9956 11540
rect 9950 11500 9956 11512
rect 10008 11540 10014 11552
rect 11238 11540 11244 11552
rect 10008 11512 11244 11540
rect 10008 11500 10014 11512
rect 11238 11500 11244 11512
rect 11296 11500 11302 11552
rect 14001 11543 14059 11549
rect 14001 11509 14013 11543
rect 14047 11540 14059 11543
rect 14090 11540 14096 11552
rect 14047 11512 14096 11540
rect 14047 11509 14059 11512
rect 14001 11503 14059 11509
rect 14090 11500 14096 11512
rect 14148 11500 14154 11552
rect 14660 11540 14688 11648
rect 14737 11645 14749 11679
rect 14783 11645 14795 11679
rect 15102 11676 15108 11688
rect 15063 11648 15108 11676
rect 14737 11639 14795 11645
rect 15102 11636 15108 11648
rect 15160 11636 15166 11688
rect 16206 11676 16212 11688
rect 16167 11648 16212 11676
rect 16206 11636 16212 11648
rect 16264 11636 16270 11688
rect 16574 11676 16580 11688
rect 16535 11648 16580 11676
rect 16574 11636 16580 11648
rect 16632 11636 16638 11688
rect 17126 11676 17132 11688
rect 17087 11648 17132 11676
rect 17126 11636 17132 11648
rect 17184 11636 17190 11688
rect 18506 11676 18512 11688
rect 18467 11648 18512 11676
rect 18506 11636 18512 11648
rect 18564 11636 18570 11688
rect 19076 11685 19104 11784
rect 23382 11772 23388 11784
rect 23440 11772 23446 11824
rect 19242 11744 19248 11756
rect 19203 11716 19248 11744
rect 19242 11704 19248 11716
rect 19300 11704 19306 11756
rect 19886 11704 19892 11756
rect 19944 11744 19950 11756
rect 20257 11747 20315 11753
rect 20257 11744 20269 11747
rect 19944 11716 20269 11744
rect 19944 11704 19950 11716
rect 20257 11713 20269 11716
rect 20303 11713 20315 11747
rect 22646 11744 22652 11756
rect 20257 11707 20315 11713
rect 20732 11716 22652 11744
rect 19061 11679 19119 11685
rect 19061 11645 19073 11679
rect 19107 11645 19119 11679
rect 20346 11676 20352 11688
rect 20307 11648 20352 11676
rect 19061 11639 19119 11645
rect 20346 11636 20352 11648
rect 20404 11636 20410 11688
rect 20732 11685 20760 11716
rect 22646 11704 22652 11716
rect 22704 11704 22710 11756
rect 24412 11753 24440 11852
rect 26326 11840 26332 11852
rect 26384 11880 26390 11892
rect 26384 11852 27108 11880
rect 26384 11840 26390 11852
rect 27080 11812 27108 11852
rect 27154 11840 27160 11892
rect 27212 11880 27218 11892
rect 27525 11883 27583 11889
rect 27525 11880 27537 11883
rect 27212 11852 27537 11880
rect 27212 11840 27218 11852
rect 27525 11849 27537 11852
rect 27571 11849 27583 11883
rect 27525 11843 27583 11849
rect 30377 11883 30435 11889
rect 30377 11849 30389 11883
rect 30423 11880 30435 11883
rect 30466 11880 30472 11892
rect 30423 11852 30472 11880
rect 30423 11849 30435 11852
rect 30377 11843 30435 11849
rect 30466 11840 30472 11852
rect 30524 11840 30530 11892
rect 38930 11880 38936 11892
rect 30668 11852 34008 11880
rect 38891 11852 38936 11880
rect 29733 11815 29791 11821
rect 27080 11784 28948 11812
rect 28920 11756 28948 11784
rect 29733 11781 29745 11815
rect 29779 11812 29791 11815
rect 30668 11812 30696 11852
rect 29779 11784 30696 11812
rect 29779 11781 29791 11784
rect 29733 11775 29791 11781
rect 30742 11772 30748 11824
rect 30800 11812 30806 11824
rect 32490 11812 32496 11824
rect 30800 11784 30972 11812
rect 32451 11784 32496 11812
rect 30800 11772 30806 11784
rect 24397 11747 24455 11753
rect 24397 11713 24409 11747
rect 24443 11713 24455 11747
rect 24397 11707 24455 11713
rect 25593 11747 25651 11753
rect 25593 11713 25605 11747
rect 25639 11744 25651 11747
rect 26421 11747 26479 11753
rect 26421 11744 26433 11747
rect 25639 11716 26433 11744
rect 25639 11713 25651 11716
rect 25593 11707 25651 11713
rect 26421 11713 26433 11716
rect 26467 11713 26479 11747
rect 26421 11707 26479 11713
rect 28902 11704 28908 11756
rect 28960 11744 28966 11756
rect 30944 11744 30972 11784
rect 32490 11772 32496 11784
rect 32548 11772 32554 11824
rect 33318 11772 33324 11824
rect 33376 11812 33382 11824
rect 33870 11812 33876 11824
rect 33376 11784 33876 11812
rect 33376 11772 33382 11784
rect 31205 11747 31263 11753
rect 31205 11744 31217 11747
rect 28960 11716 30328 11744
rect 30944 11716 31217 11744
rect 28960 11704 28966 11716
rect 20717 11679 20775 11685
rect 20717 11645 20729 11679
rect 20763 11645 20775 11679
rect 20717 11639 20775 11645
rect 20901 11679 20959 11685
rect 20901 11645 20913 11679
rect 20947 11676 20959 11679
rect 20990 11676 20996 11688
rect 20947 11648 20996 11676
rect 20947 11645 20959 11648
rect 20901 11639 20959 11645
rect 20990 11636 20996 11648
rect 21048 11636 21054 11688
rect 21358 11676 21364 11688
rect 21319 11648 21364 11676
rect 21358 11636 21364 11648
rect 21416 11636 21422 11688
rect 22557 11679 22615 11685
rect 22557 11645 22569 11679
rect 22603 11676 22615 11679
rect 23290 11676 23296 11688
rect 22603 11648 23296 11676
rect 22603 11645 22615 11648
rect 22557 11639 22615 11645
rect 23290 11636 23296 11648
rect 23348 11636 23354 11688
rect 23661 11679 23719 11685
rect 23661 11645 23673 11679
rect 23707 11676 23719 11679
rect 24210 11676 24216 11688
rect 23707 11648 24216 11676
rect 23707 11645 23719 11648
rect 23661 11639 23719 11645
rect 24210 11636 24216 11648
rect 24268 11636 24274 11688
rect 24486 11676 24492 11688
rect 24399 11648 24492 11676
rect 24486 11636 24492 11648
rect 24544 11636 24550 11688
rect 24946 11676 24952 11688
rect 24907 11648 24952 11676
rect 24946 11636 24952 11648
rect 25004 11636 25010 11688
rect 25041 11679 25099 11685
rect 25041 11645 25053 11679
rect 25087 11676 25099 11679
rect 25130 11676 25136 11688
rect 25087 11648 25136 11676
rect 25087 11645 25099 11648
rect 25041 11639 25099 11645
rect 25130 11636 25136 11648
rect 25188 11676 25194 11688
rect 26145 11679 26203 11685
rect 25188 11648 25360 11676
rect 25188 11636 25194 11648
rect 16482 11568 16488 11620
rect 16540 11608 16546 11620
rect 17313 11611 17371 11617
rect 17313 11608 17325 11611
rect 16540 11580 17325 11608
rect 16540 11568 16546 11580
rect 17313 11577 17325 11580
rect 17359 11577 17371 11611
rect 17313 11571 17371 11577
rect 20162 11568 20168 11620
rect 20220 11608 20226 11620
rect 24504 11608 24532 11636
rect 25332 11620 25360 11648
rect 26145 11645 26157 11679
rect 26191 11645 26203 11679
rect 27614 11676 27620 11688
rect 26145 11639 26203 11645
rect 26252 11648 27620 11676
rect 24762 11608 24768 11620
rect 20220 11580 24440 11608
rect 24504 11580 24768 11608
rect 20220 11568 20226 11580
rect 22002 11540 22008 11552
rect 14660 11512 22008 11540
rect 22002 11500 22008 11512
rect 22060 11500 22066 11552
rect 22278 11500 22284 11552
rect 22336 11540 22342 11552
rect 22741 11543 22799 11549
rect 22741 11540 22753 11543
rect 22336 11512 22753 11540
rect 22336 11500 22342 11512
rect 22741 11509 22753 11512
rect 22787 11540 22799 11543
rect 23382 11540 23388 11552
rect 22787 11512 23388 11540
rect 22787 11509 22799 11512
rect 22741 11503 22799 11509
rect 23382 11500 23388 11512
rect 23440 11500 23446 11552
rect 24412 11540 24440 11580
rect 24762 11568 24768 11580
rect 24820 11568 24826 11620
rect 25314 11568 25320 11620
rect 25372 11568 25378 11620
rect 25590 11568 25596 11620
rect 25648 11608 25654 11620
rect 26160 11608 26188 11639
rect 25648 11580 26188 11608
rect 25648 11568 25654 11580
rect 26252 11540 26280 11648
rect 27614 11636 27620 11648
rect 27672 11636 27678 11688
rect 28534 11676 28540 11688
rect 28495 11648 28540 11676
rect 28534 11636 28540 11648
rect 28592 11636 28598 11688
rect 29641 11679 29699 11685
rect 29641 11645 29653 11679
rect 29687 11676 29699 11679
rect 30190 11676 30196 11688
rect 29687 11648 30196 11676
rect 29687 11645 29699 11648
rect 29641 11639 29699 11645
rect 30190 11636 30196 11648
rect 30248 11636 30254 11688
rect 30300 11685 30328 11716
rect 31205 11713 31217 11716
rect 31251 11713 31263 11747
rect 31205 11707 31263 11713
rect 30285 11679 30343 11685
rect 30285 11645 30297 11679
rect 30331 11645 30343 11679
rect 30285 11639 30343 11645
rect 30558 11636 30564 11688
rect 30616 11676 30622 11688
rect 30929 11679 30987 11685
rect 30929 11676 30941 11679
rect 30616 11648 30941 11676
rect 30616 11636 30622 11648
rect 30929 11645 30941 11648
rect 30975 11645 30987 11679
rect 30929 11639 30987 11645
rect 31478 11636 31484 11688
rect 31536 11676 31542 11688
rect 33594 11676 33600 11688
rect 31536 11648 33456 11676
rect 33555 11648 33600 11676
rect 31536 11636 31542 11648
rect 30742 11608 30748 11620
rect 28644 11580 30748 11608
rect 24412 11512 26280 11540
rect 26694 11500 26700 11552
rect 26752 11540 26758 11552
rect 28644 11549 28672 11580
rect 30742 11568 30748 11580
rect 30800 11568 30806 11620
rect 33137 11611 33195 11617
rect 33137 11577 33149 11611
rect 33183 11608 33195 11611
rect 33226 11608 33232 11620
rect 33183 11580 33232 11608
rect 33183 11577 33195 11580
rect 33137 11571 33195 11577
rect 33226 11568 33232 11580
rect 33284 11568 33290 11620
rect 33428 11608 33456 11648
rect 33594 11636 33600 11648
rect 33652 11636 33658 11688
rect 33796 11685 33824 11784
rect 33870 11772 33876 11784
rect 33928 11772 33934 11824
rect 33980 11685 34008 11852
rect 38930 11840 38936 11852
rect 38988 11840 38994 11892
rect 34422 11772 34428 11824
rect 34480 11812 34486 11824
rect 34480 11784 37504 11812
rect 34480 11772 34486 11784
rect 33781 11679 33839 11685
rect 33781 11645 33793 11679
rect 33827 11645 33839 11679
rect 33781 11639 33839 11645
rect 33965 11679 34023 11685
rect 33965 11645 33977 11679
rect 34011 11645 34023 11679
rect 35342 11676 35348 11688
rect 35303 11648 35348 11676
rect 33965 11639 34023 11645
rect 35342 11636 35348 11648
rect 35400 11636 35406 11688
rect 35526 11676 35532 11688
rect 35487 11648 35532 11676
rect 35526 11636 35532 11648
rect 35584 11636 35590 11688
rect 35802 11636 35808 11688
rect 35860 11676 35866 11688
rect 35897 11679 35955 11685
rect 35897 11676 35909 11679
rect 35860 11648 35909 11676
rect 35860 11636 35866 11648
rect 35897 11645 35909 11648
rect 35943 11645 35955 11679
rect 35897 11639 35955 11645
rect 35986 11636 35992 11688
rect 36044 11676 36050 11688
rect 36814 11676 36820 11688
rect 36044 11648 36089 11676
rect 36775 11648 36820 11676
rect 36044 11636 36050 11648
rect 36814 11636 36820 11648
rect 36872 11636 36878 11688
rect 37001 11679 37059 11685
rect 37001 11645 37013 11679
rect 37047 11645 37059 11679
rect 37366 11676 37372 11688
rect 37327 11648 37372 11676
rect 37001 11639 37059 11645
rect 37016 11608 37044 11639
rect 37366 11636 37372 11648
rect 37424 11636 37430 11688
rect 37476 11676 37504 11784
rect 37553 11679 37611 11685
rect 37553 11676 37565 11679
rect 37476 11648 37565 11676
rect 37553 11645 37565 11648
rect 37599 11645 37611 11679
rect 37553 11639 37611 11645
rect 37737 11679 37795 11685
rect 37737 11645 37749 11679
rect 37783 11645 37795 11679
rect 37737 11639 37795 11645
rect 33428 11580 37044 11608
rect 37182 11568 37188 11620
rect 37240 11608 37246 11620
rect 37752 11608 37780 11639
rect 37826 11636 37832 11688
rect 37884 11676 37890 11688
rect 38749 11679 38807 11685
rect 38749 11676 38761 11679
rect 37884 11648 38761 11676
rect 37884 11636 37890 11648
rect 38749 11645 38761 11648
rect 38795 11645 38807 11679
rect 38749 11639 38807 11645
rect 37240 11580 37780 11608
rect 38289 11611 38347 11617
rect 37240 11568 37246 11580
rect 38289 11577 38301 11611
rect 38335 11608 38347 11611
rect 38378 11608 38384 11620
rect 38335 11580 38384 11608
rect 38335 11577 38347 11580
rect 38289 11571 38347 11577
rect 38378 11568 38384 11580
rect 38436 11568 38442 11620
rect 28629 11543 28687 11549
rect 28629 11540 28641 11543
rect 26752 11512 28641 11540
rect 26752 11500 26758 11512
rect 28629 11509 28641 11512
rect 28675 11509 28687 11543
rect 28629 11503 28687 11509
rect 29914 11500 29920 11552
rect 29972 11540 29978 11552
rect 32490 11540 32496 11552
rect 29972 11512 32496 11540
rect 29972 11500 29978 11512
rect 32490 11500 32496 11512
rect 32548 11500 32554 11552
rect 35161 11543 35219 11549
rect 35161 11509 35173 11543
rect 35207 11540 35219 11543
rect 36170 11540 36176 11552
rect 35207 11512 36176 11540
rect 35207 11509 35219 11512
rect 35161 11503 35219 11509
rect 36170 11500 36176 11512
rect 36228 11500 36234 11552
rect 1104 11450 39836 11472
rect 1104 11398 19606 11450
rect 19658 11398 19670 11450
rect 19722 11398 19734 11450
rect 19786 11398 19798 11450
rect 19850 11398 39836 11450
rect 1104 11376 39836 11398
rect 10318 11336 10324 11348
rect 6656 11308 10324 11336
rect 6178 11268 6184 11280
rect 5920 11240 6184 11268
rect 2314 11160 2320 11212
rect 2372 11200 2378 11212
rect 2777 11203 2835 11209
rect 2777 11200 2789 11203
rect 2372 11172 2789 11200
rect 2372 11160 2378 11172
rect 2777 11169 2789 11172
rect 2823 11169 2835 11203
rect 3234 11200 3240 11212
rect 3195 11172 3240 11200
rect 2777 11163 2835 11169
rect 3234 11160 3240 11172
rect 3292 11160 3298 11212
rect 3878 11160 3884 11212
rect 3936 11200 3942 11212
rect 4617 11203 4675 11209
rect 4617 11200 4629 11203
rect 3936 11172 4629 11200
rect 3936 11160 3942 11172
rect 4617 11169 4629 11172
rect 4663 11169 4675 11203
rect 5350 11200 5356 11212
rect 5311 11172 5356 11200
rect 4617 11163 4675 11169
rect 5350 11160 5356 11172
rect 5408 11160 5414 11212
rect 5920 11209 5948 11240
rect 6178 11228 6184 11240
rect 6236 11228 6242 11280
rect 6656 11209 6684 11308
rect 10318 11296 10324 11308
rect 10376 11296 10382 11348
rect 13722 11296 13728 11348
rect 13780 11336 13786 11348
rect 18693 11339 18751 11345
rect 13780 11308 17172 11336
rect 13780 11296 13786 11308
rect 7098 11268 7104 11280
rect 6748 11240 7104 11268
rect 5905 11203 5963 11209
rect 5905 11169 5917 11203
rect 5951 11169 5963 11203
rect 5905 11163 5963 11169
rect 6273 11203 6331 11209
rect 6273 11169 6285 11203
rect 6319 11169 6331 11203
rect 6273 11163 6331 11169
rect 6641 11203 6699 11209
rect 6641 11169 6653 11203
rect 6687 11169 6699 11203
rect 6641 11163 6699 11169
rect 3326 11132 3332 11144
rect 3287 11104 3332 11132
rect 3326 11092 3332 11104
rect 3384 11092 3390 11144
rect 5442 11132 5448 11144
rect 5403 11104 5448 11132
rect 5442 11092 5448 11104
rect 5500 11092 5506 11144
rect 6288 11132 6316 11163
rect 6748 11132 6776 11240
rect 7098 11228 7104 11240
rect 7156 11228 7162 11280
rect 9030 11268 9036 11280
rect 8404 11240 9036 11268
rect 6917 11203 6975 11209
rect 6917 11200 6929 11203
rect 6288 11104 6776 11132
rect 6840 11172 6929 11200
rect 6840 11064 6868 11172
rect 6917 11169 6929 11172
rect 6963 11169 6975 11203
rect 6917 11163 6975 11169
rect 7006 11160 7012 11212
rect 7064 11200 7070 11212
rect 7653 11203 7711 11209
rect 7653 11200 7665 11203
rect 7064 11172 7665 11200
rect 7064 11160 7070 11172
rect 7653 11169 7665 11172
rect 7699 11169 7711 11203
rect 8018 11200 8024 11212
rect 7979 11172 8024 11200
rect 7653 11163 7711 11169
rect 8018 11160 8024 11172
rect 8076 11160 8082 11212
rect 8404 11209 8432 11240
rect 9030 11228 9036 11240
rect 9088 11268 9094 11280
rect 11698 11268 11704 11280
rect 9088 11240 11704 11268
rect 9088 11228 9094 11240
rect 8389 11203 8447 11209
rect 8389 11169 8401 11203
rect 8435 11169 8447 11203
rect 9766 11200 9772 11212
rect 9727 11172 9772 11200
rect 8389 11163 8447 11169
rect 9766 11160 9772 11172
rect 9824 11160 9830 11212
rect 10042 11200 10048 11212
rect 10003 11172 10048 11200
rect 10042 11160 10048 11172
rect 10100 11160 10106 11212
rect 10428 11209 10456 11240
rect 11698 11228 11704 11240
rect 11756 11228 11762 11280
rect 12621 11271 12679 11277
rect 12621 11237 12633 11271
rect 12667 11268 12679 11271
rect 13078 11268 13084 11280
rect 12667 11240 13084 11268
rect 12667 11237 12679 11240
rect 12621 11231 12679 11237
rect 13078 11228 13084 11240
rect 13136 11228 13142 11280
rect 17144 11268 17172 11308
rect 18693 11305 18705 11339
rect 18739 11336 18751 11339
rect 18874 11336 18880 11348
rect 18739 11308 18880 11336
rect 18739 11305 18751 11308
rect 18693 11299 18751 11305
rect 18874 11296 18880 11308
rect 18932 11296 18938 11348
rect 20622 11336 20628 11348
rect 18984 11308 20628 11336
rect 18984 11268 19012 11308
rect 20622 11296 20628 11308
rect 20680 11296 20686 11348
rect 30190 11296 30196 11348
rect 30248 11336 30254 11348
rect 31202 11336 31208 11348
rect 30248 11308 31208 11336
rect 30248 11296 30254 11308
rect 31202 11296 31208 11308
rect 31260 11296 31266 11348
rect 31481 11339 31539 11345
rect 31481 11305 31493 11339
rect 31527 11336 31539 11339
rect 31570 11336 31576 11348
rect 31527 11308 31576 11336
rect 31527 11305 31539 11308
rect 31481 11299 31539 11305
rect 31570 11296 31576 11308
rect 31628 11296 31634 11348
rect 32217 11339 32275 11345
rect 32217 11305 32229 11339
rect 32263 11336 32275 11339
rect 35526 11336 35532 11348
rect 32263 11308 35532 11336
rect 32263 11305 32275 11308
rect 32217 11299 32275 11305
rect 35526 11296 35532 11308
rect 35584 11296 35590 11348
rect 35894 11296 35900 11348
rect 35952 11336 35958 11348
rect 35952 11308 36952 11336
rect 35952 11296 35958 11308
rect 20346 11268 20352 11280
rect 13372 11240 15332 11268
rect 17144 11240 19012 11268
rect 20307 11240 20352 11268
rect 10413 11203 10471 11209
rect 10413 11169 10425 11203
rect 10459 11169 10471 11203
rect 10413 11163 10471 11169
rect 10778 11160 10784 11212
rect 10836 11200 10842 11212
rect 10873 11203 10931 11209
rect 10873 11200 10885 11203
rect 10836 11172 10885 11200
rect 10836 11160 10842 11172
rect 10873 11169 10885 11172
rect 10919 11169 10931 11203
rect 11606 11200 11612 11212
rect 11567 11172 11612 11200
rect 10873 11163 10931 11169
rect 10888 11132 10916 11163
rect 11606 11160 11612 11172
rect 11664 11160 11670 11212
rect 12066 11200 12072 11212
rect 12027 11172 12072 11200
rect 12066 11160 12072 11172
rect 12124 11160 12130 11212
rect 12158 11160 12164 11212
rect 12216 11200 12222 11212
rect 12345 11203 12403 11209
rect 12345 11200 12357 11203
rect 12216 11172 12357 11200
rect 12216 11160 12222 11172
rect 12345 11169 12357 11172
rect 12391 11169 12403 11203
rect 12345 11163 12403 11169
rect 13372 11132 13400 11240
rect 15304 11212 15332 11240
rect 20346 11228 20352 11240
rect 20404 11228 20410 11280
rect 22462 11228 22468 11280
rect 22520 11268 22526 11280
rect 26694 11268 26700 11280
rect 22520 11240 22968 11268
rect 22520 11228 22526 11240
rect 13538 11200 13544 11212
rect 13499 11172 13544 11200
rect 13538 11160 13544 11172
rect 13596 11160 13602 11212
rect 13906 11200 13912 11212
rect 13867 11172 13912 11200
rect 13906 11160 13912 11172
rect 13964 11160 13970 11212
rect 14458 11160 14464 11212
rect 14516 11200 14522 11212
rect 14553 11203 14611 11209
rect 14553 11200 14565 11203
rect 14516 11172 14565 11200
rect 14516 11160 14522 11172
rect 14553 11169 14565 11172
rect 14599 11169 14611 11203
rect 14553 11163 14611 11169
rect 14642 11160 14648 11212
rect 14700 11200 14706 11212
rect 15286 11200 15292 11212
rect 14700 11172 14745 11200
rect 15247 11172 15292 11200
rect 14700 11160 14706 11172
rect 15286 11160 15292 11172
rect 15344 11160 15350 11212
rect 16209 11203 16267 11209
rect 16209 11169 16221 11203
rect 16255 11200 16267 11203
rect 16942 11200 16948 11212
rect 16255 11172 16948 11200
rect 16255 11169 16267 11172
rect 16209 11163 16267 11169
rect 16942 11160 16948 11172
rect 17000 11160 17006 11212
rect 18506 11200 18512 11212
rect 18467 11172 18512 11200
rect 18506 11160 18512 11172
rect 18564 11160 18570 11212
rect 18969 11203 19027 11209
rect 18969 11169 18981 11203
rect 19015 11169 19027 11203
rect 18969 11163 19027 11169
rect 10888 11104 13400 11132
rect 14001 11135 14059 11141
rect 14001 11101 14013 11135
rect 14047 11132 14059 11135
rect 16114 11132 16120 11144
rect 14047 11104 16120 11132
rect 14047 11101 14059 11104
rect 14001 11095 14059 11101
rect 16114 11092 16120 11104
rect 16172 11092 16178 11144
rect 16482 11092 16488 11144
rect 16540 11132 16546 11144
rect 16540 11104 16585 11132
rect 16540 11092 16546 11104
rect 10962 11064 10968 11076
rect 6840 11036 6960 11064
rect 10923 11036 10968 11064
rect 4433 10999 4491 11005
rect 4433 10965 4445 10999
rect 4479 10996 4491 10999
rect 4614 10996 4620 11008
rect 4479 10968 4620 10996
rect 4479 10965 4491 10968
rect 4433 10959 4491 10965
rect 4614 10956 4620 10968
rect 4672 10956 4678 11008
rect 6932 10996 6960 11036
rect 10962 11024 10968 11036
rect 11020 11024 11026 11076
rect 13357 11067 13415 11073
rect 13357 11033 13369 11067
rect 13403 11064 13415 11067
rect 13446 11064 13452 11076
rect 13403 11036 13452 11064
rect 13403 11033 13415 11036
rect 13357 11027 13415 11033
rect 13446 11024 13452 11036
rect 13504 11024 13510 11076
rect 15473 11067 15531 11073
rect 15473 11033 15485 11067
rect 15519 11064 15531 11067
rect 15562 11064 15568 11076
rect 15519 11036 15568 11064
rect 15519 11033 15531 11036
rect 15473 11027 15531 11033
rect 15562 11024 15568 11036
rect 15620 11064 15626 11076
rect 16206 11064 16212 11076
rect 15620 11036 16212 11064
rect 15620 11024 15626 11036
rect 16206 11024 16212 11036
rect 16264 11024 16270 11076
rect 18984 11064 19012 11163
rect 19334 11160 19340 11212
rect 19392 11200 19398 11212
rect 19889 11203 19947 11209
rect 19889 11200 19901 11203
rect 19392 11172 19901 11200
rect 19392 11160 19398 11172
rect 19889 11169 19901 11172
rect 19935 11200 19947 11203
rect 19978 11200 19984 11212
rect 19935 11172 19984 11200
rect 19935 11169 19947 11172
rect 19889 11163 19947 11169
rect 19978 11160 19984 11172
rect 20036 11160 20042 11212
rect 20162 11200 20168 11212
rect 20123 11172 20168 11200
rect 20162 11160 20168 11172
rect 20220 11160 20226 11212
rect 21542 11200 21548 11212
rect 21503 11172 21548 11200
rect 21542 11160 21548 11172
rect 21600 11160 21606 11212
rect 21910 11160 21916 11212
rect 21968 11209 21974 11212
rect 21968 11203 22017 11209
rect 21968 11169 21971 11203
rect 22005 11169 22017 11203
rect 22830 11200 22836 11212
rect 22791 11172 22836 11200
rect 21968 11163 22017 11169
rect 21968 11160 21974 11163
rect 22830 11160 22836 11172
rect 22888 11160 22894 11212
rect 22940 11209 22968 11240
rect 23683 11240 26700 11268
rect 22925 11203 22983 11209
rect 22925 11169 22937 11203
rect 22971 11169 22983 11203
rect 23290 11200 23296 11212
rect 23251 11172 23296 11200
rect 22925 11163 22983 11169
rect 23290 11160 23296 11172
rect 23348 11160 23354 11212
rect 21634 11092 21640 11144
rect 21692 11132 21698 11144
rect 21821 11135 21879 11141
rect 21821 11132 21833 11135
rect 21692 11104 21833 11132
rect 21692 11092 21698 11104
rect 21821 11101 21833 11104
rect 21867 11101 21879 11135
rect 23683 11132 23711 11240
rect 24762 11200 24768 11212
rect 24723 11172 24768 11200
rect 24762 11160 24768 11172
rect 24820 11160 24826 11212
rect 25314 11200 25320 11212
rect 25275 11172 25320 11200
rect 25314 11160 25320 11172
rect 25372 11160 25378 11212
rect 25516 11209 25544 11240
rect 26694 11228 26700 11240
rect 26752 11228 26758 11280
rect 30653 11271 30711 11277
rect 30653 11237 30665 11271
rect 30699 11268 30711 11271
rect 31386 11268 31392 11280
rect 30699 11240 31392 11268
rect 30699 11237 30711 11240
rect 30653 11231 30711 11237
rect 31386 11228 31392 11240
rect 31444 11228 31450 11280
rect 31496 11240 33548 11268
rect 25501 11203 25559 11209
rect 25501 11169 25513 11203
rect 25547 11169 25559 11203
rect 26602 11200 26608 11212
rect 26563 11172 26608 11200
rect 25501 11163 25559 11169
rect 26602 11160 26608 11172
rect 26660 11160 26666 11212
rect 27338 11160 27344 11212
rect 27396 11200 27402 11212
rect 29365 11203 29423 11209
rect 29365 11200 29377 11203
rect 27396 11172 29377 11200
rect 27396 11160 27402 11172
rect 29365 11169 29377 11172
rect 29411 11169 29423 11203
rect 29914 11200 29920 11212
rect 29875 11172 29920 11200
rect 29365 11163 29423 11169
rect 29914 11160 29920 11172
rect 29972 11160 29978 11212
rect 30834 11160 30840 11212
rect 30892 11200 30898 11212
rect 31110 11200 31116 11212
rect 30892 11172 31116 11200
rect 30892 11160 30898 11172
rect 31110 11160 31116 11172
rect 31168 11200 31174 11212
rect 31297 11203 31355 11209
rect 31297 11200 31309 11203
rect 31168 11172 31309 11200
rect 31168 11160 31174 11172
rect 31297 11169 31309 11172
rect 31343 11169 31355 11203
rect 31496 11200 31524 11240
rect 31297 11163 31355 11169
rect 31404 11172 31524 11200
rect 32217 11203 32275 11209
rect 21821 11095 21879 11101
rect 21928 11104 23711 11132
rect 23753 11135 23811 11141
rect 21928 11064 21956 11104
rect 23753 11101 23765 11135
rect 23799 11101 23811 11135
rect 23753 11095 23811 11101
rect 24673 11135 24731 11141
rect 24673 11101 24685 11135
rect 24719 11101 24731 11135
rect 24673 11095 24731 11101
rect 25869 11135 25927 11141
rect 25869 11101 25881 11135
rect 25915 11132 25927 11135
rect 26881 11135 26939 11141
rect 26881 11132 26893 11135
rect 25915 11104 26893 11132
rect 25915 11101 25927 11104
rect 25869 11095 25927 11101
rect 26881 11101 26893 11104
rect 26927 11101 26939 11135
rect 31404 11132 31432 11172
rect 32217 11169 32229 11203
rect 32263 11200 32275 11203
rect 32309 11203 32367 11209
rect 32309 11200 32321 11203
rect 32263 11172 32321 11200
rect 32263 11169 32275 11172
rect 32217 11163 32275 11169
rect 32309 11169 32321 11172
rect 32355 11169 32367 11203
rect 32309 11163 32367 11169
rect 33045 11203 33103 11209
rect 33045 11169 33057 11203
rect 33091 11200 33103 11203
rect 33134 11200 33140 11212
rect 33091 11172 33140 11200
rect 33091 11169 33103 11172
rect 33045 11163 33103 11169
rect 33134 11160 33140 11172
rect 33192 11160 33198 11212
rect 33318 11200 33324 11212
rect 33279 11172 33324 11200
rect 33318 11160 33324 11172
rect 33376 11160 33382 11212
rect 33520 11209 33548 11240
rect 33778 11228 33784 11280
rect 33836 11268 33842 11280
rect 35802 11268 35808 11280
rect 33836 11240 35808 11268
rect 33836 11228 33842 11240
rect 33505 11203 33563 11209
rect 33505 11169 33517 11203
rect 33551 11169 33563 11203
rect 33505 11163 33563 11169
rect 34241 11203 34299 11209
rect 34241 11169 34253 11203
rect 34287 11169 34299 11203
rect 34241 11163 34299 11169
rect 26881 11095 26939 11101
rect 31220 11104 31432 11132
rect 18984 11036 21956 11064
rect 22002 11024 22008 11076
rect 22060 11064 22066 11076
rect 23106 11064 23112 11076
rect 22060 11036 23112 11064
rect 22060 11024 22066 11036
rect 23106 11024 23112 11036
rect 23164 11024 23170 11076
rect 7466 10996 7472 11008
rect 6932 10968 7472 10996
rect 7466 10956 7472 10968
rect 7524 10996 7530 11008
rect 14090 10996 14096 11008
rect 7524 10968 14096 10996
rect 7524 10956 7530 10968
rect 14090 10956 14096 10968
rect 14148 10956 14154 11008
rect 16574 10956 16580 11008
rect 16632 10996 16638 11008
rect 17589 10999 17647 11005
rect 17589 10996 17601 10999
rect 16632 10968 17601 10996
rect 16632 10956 16638 10968
rect 17589 10965 17601 10968
rect 17635 10965 17647 10999
rect 23768 10996 23796 11095
rect 24688 11064 24716 11095
rect 25130 11064 25136 11076
rect 24688 11036 25136 11064
rect 25130 11024 25136 11036
rect 25188 11064 25194 11076
rect 28169 11067 28227 11073
rect 25188 11036 25820 11064
rect 25188 11024 25194 11036
rect 25682 10996 25688 11008
rect 23768 10968 25688 10996
rect 17589 10959 17647 10965
rect 25682 10956 25688 10968
rect 25740 10956 25746 11008
rect 25792 10996 25820 11036
rect 28169 11033 28181 11067
rect 28215 11064 28227 11067
rect 28534 11064 28540 11076
rect 28215 11036 28540 11064
rect 28215 11033 28227 11036
rect 28169 11027 28227 11033
rect 28534 11024 28540 11036
rect 28592 11064 28598 11076
rect 31220 11064 31248 11104
rect 31478 11092 31484 11144
rect 31536 11132 31542 11144
rect 34256 11132 34284 11163
rect 34514 11160 34520 11212
rect 34572 11200 34578 11212
rect 34790 11200 34796 11212
rect 34572 11172 34796 11200
rect 34572 11160 34578 11172
rect 34790 11160 34796 11172
rect 34848 11160 34854 11212
rect 35084 11209 35112 11240
rect 35802 11228 35808 11240
rect 35860 11228 35866 11280
rect 36170 11268 36176 11280
rect 36131 11240 36176 11268
rect 36170 11228 36176 11240
rect 36228 11228 36234 11280
rect 36924 11277 36952 11308
rect 36357 11271 36415 11277
rect 36357 11268 36369 11271
rect 36280 11240 36369 11268
rect 35069 11203 35127 11209
rect 35069 11169 35081 11203
rect 35115 11169 35127 11203
rect 35069 11163 35127 11169
rect 35713 11203 35771 11209
rect 35713 11169 35725 11203
rect 35759 11200 35771 11203
rect 35986 11200 35992 11212
rect 35759 11172 35992 11200
rect 35759 11169 35771 11172
rect 35713 11163 35771 11169
rect 35986 11160 35992 11172
rect 36044 11160 36050 11212
rect 31536 11104 34284 11132
rect 34701 11135 34759 11141
rect 31536 11092 31542 11104
rect 34701 11101 34713 11135
rect 34747 11132 34759 11135
rect 36280 11132 36308 11240
rect 36357 11237 36369 11240
rect 36403 11237 36415 11271
rect 36357 11231 36415 11237
rect 36541 11271 36599 11277
rect 36541 11237 36553 11271
rect 36587 11237 36599 11271
rect 36541 11231 36599 11237
rect 36909 11271 36967 11277
rect 36909 11237 36921 11271
rect 36955 11237 36967 11271
rect 36909 11231 36967 11237
rect 36446 11200 36452 11212
rect 36407 11172 36452 11200
rect 36446 11160 36452 11172
rect 36504 11160 36510 11212
rect 34747 11104 36308 11132
rect 34747 11101 34759 11104
rect 34701 11095 34759 11101
rect 28592 11036 31248 11064
rect 31404 11036 31616 11064
rect 28592 11024 28598 11036
rect 27246 10996 27252 11008
rect 25792 10968 27252 10996
rect 27246 10956 27252 10968
rect 27304 10956 27310 11008
rect 27706 10956 27712 11008
rect 27764 10996 27770 11008
rect 27890 10996 27896 11008
rect 27764 10968 27896 10996
rect 27764 10956 27770 10968
rect 27890 10956 27896 10968
rect 27948 10956 27954 11008
rect 28074 10956 28080 11008
rect 28132 10996 28138 11008
rect 31404 10996 31432 11036
rect 28132 10968 31432 10996
rect 31588 10996 31616 11036
rect 31662 11024 31668 11076
rect 31720 11064 31726 11076
rect 32217 11067 32275 11073
rect 32217 11064 32229 11067
rect 31720 11036 32229 11064
rect 31720 11024 31726 11036
rect 32217 11033 32229 11036
rect 32263 11033 32275 11067
rect 32217 11027 32275 11033
rect 32401 11067 32459 11073
rect 32401 11033 32413 11067
rect 32447 11064 32459 11067
rect 36556 11064 36584 11231
rect 38194 11228 38200 11280
rect 38252 11268 38258 11280
rect 38841 11271 38899 11277
rect 38841 11268 38853 11271
rect 38252 11240 38853 11268
rect 38252 11228 38258 11240
rect 38841 11237 38853 11240
rect 38887 11237 38899 11271
rect 38841 11231 38899 11237
rect 38105 11203 38163 11209
rect 38105 11200 38117 11203
rect 32447 11036 36584 11064
rect 36924 11172 38117 11200
rect 32447 11033 32459 11036
rect 32401 11027 32459 11033
rect 35894 10996 35900 11008
rect 31588 10968 35900 10996
rect 28132 10956 28138 10968
rect 35894 10956 35900 10968
rect 35952 10956 35958 11008
rect 36354 10956 36360 11008
rect 36412 10996 36418 11008
rect 36924 10996 36952 11172
rect 38105 11169 38117 11172
rect 38151 11169 38163 11203
rect 38562 11200 38568 11212
rect 38523 11172 38568 11200
rect 38105 11163 38163 11169
rect 38562 11160 38568 11172
rect 38620 11160 38626 11212
rect 37826 11132 37832 11144
rect 37787 11104 37832 11132
rect 37826 11092 37832 11104
rect 37884 11092 37890 11144
rect 36412 10968 36952 10996
rect 36412 10956 36418 10968
rect 1104 10906 39836 10928
rect 1104 10854 4246 10906
rect 4298 10854 4310 10906
rect 4362 10854 4374 10906
rect 4426 10854 4438 10906
rect 4490 10854 34966 10906
rect 35018 10854 35030 10906
rect 35082 10854 35094 10906
rect 35146 10854 35158 10906
rect 35210 10854 39836 10906
rect 1104 10832 39836 10854
rect 2498 10792 2504 10804
rect 2459 10764 2504 10792
rect 2498 10752 2504 10764
rect 2556 10752 2562 10804
rect 3234 10752 3240 10804
rect 3292 10792 3298 10804
rect 3878 10792 3884 10804
rect 3292 10764 3884 10792
rect 3292 10752 3298 10764
rect 3878 10752 3884 10764
rect 3936 10792 3942 10804
rect 4341 10795 4399 10801
rect 4341 10792 4353 10795
rect 3936 10764 4353 10792
rect 3936 10752 3942 10764
rect 4341 10761 4353 10764
rect 4387 10761 4399 10795
rect 4341 10755 4399 10761
rect 7009 10795 7067 10801
rect 7009 10761 7021 10795
rect 7055 10792 7067 10795
rect 7098 10792 7104 10804
rect 7055 10764 7104 10792
rect 7055 10761 7067 10764
rect 7009 10755 7067 10761
rect 7098 10752 7104 10764
rect 7156 10792 7162 10804
rect 7558 10792 7564 10804
rect 7156 10764 7564 10792
rect 7156 10752 7162 10764
rect 7558 10752 7564 10764
rect 7616 10752 7622 10804
rect 9030 10792 9036 10804
rect 8991 10764 9036 10792
rect 9030 10752 9036 10764
rect 9088 10752 9094 10804
rect 10686 10752 10692 10804
rect 10744 10792 10750 10804
rect 28074 10792 28080 10804
rect 10744 10764 28080 10792
rect 10744 10752 10750 10764
rect 28074 10752 28080 10764
rect 28132 10752 28138 10804
rect 29089 10795 29147 10801
rect 29089 10761 29101 10795
rect 29135 10792 29147 10795
rect 31202 10792 31208 10804
rect 29135 10764 31208 10792
rect 29135 10761 29147 10764
rect 29089 10755 29147 10761
rect 31202 10752 31208 10764
rect 31260 10752 31266 10804
rect 38746 10792 38752 10804
rect 31404 10764 38752 10792
rect 12618 10724 12624 10736
rect 6840 10696 12624 10724
rect 2225 10659 2283 10665
rect 2225 10625 2237 10659
rect 2271 10656 2283 10659
rect 2866 10656 2872 10668
rect 2271 10628 2872 10656
rect 2271 10625 2283 10628
rect 2225 10619 2283 10625
rect 2866 10616 2872 10628
rect 2924 10616 2930 10668
rect 4614 10656 4620 10668
rect 3436 10628 4620 10656
rect 2317 10591 2375 10597
rect 2317 10557 2329 10591
rect 2363 10588 2375 10591
rect 2958 10588 2964 10600
rect 2363 10560 2964 10588
rect 2363 10557 2375 10560
rect 2317 10551 2375 10557
rect 2958 10548 2964 10560
rect 3016 10548 3022 10600
rect 3436 10597 3464 10628
rect 4614 10616 4620 10628
rect 4672 10616 4678 10668
rect 3421 10591 3479 10597
rect 3421 10557 3433 10591
rect 3467 10557 3479 10591
rect 3421 10551 3479 10557
rect 4249 10591 4307 10597
rect 4249 10557 4261 10591
rect 4295 10588 4307 10591
rect 4338 10588 4344 10600
rect 4295 10560 4344 10588
rect 4295 10557 4307 10560
rect 4249 10551 4307 10557
rect 4338 10548 4344 10560
rect 4396 10548 4402 10600
rect 6178 10548 6184 10600
rect 6236 10588 6242 10600
rect 6840 10597 6868 10696
rect 12618 10684 12624 10696
rect 12676 10684 12682 10736
rect 13262 10724 13268 10736
rect 13223 10696 13268 10724
rect 13262 10684 13268 10696
rect 13320 10684 13326 10736
rect 16114 10684 16120 10736
rect 16172 10724 16178 10736
rect 21085 10727 21143 10733
rect 21085 10724 21097 10727
rect 16172 10696 21097 10724
rect 16172 10684 16178 10696
rect 21085 10693 21097 10696
rect 21131 10693 21143 10727
rect 29454 10724 29460 10736
rect 21085 10687 21143 10693
rect 27080 10696 29460 10724
rect 8021 10659 8079 10665
rect 8021 10625 8033 10659
rect 8067 10656 8079 10659
rect 8478 10656 8484 10668
rect 8067 10628 8484 10656
rect 8067 10625 8079 10628
rect 8021 10619 8079 10625
rect 8478 10616 8484 10628
rect 8536 10616 8542 10668
rect 9030 10656 9036 10668
rect 8680 10628 9036 10656
rect 6825 10591 6883 10597
rect 6825 10588 6837 10591
rect 6236 10560 6837 10588
rect 6236 10548 6242 10560
rect 6825 10557 6837 10560
rect 6871 10557 6883 10591
rect 7650 10588 7656 10600
rect 7611 10560 7656 10588
rect 6825 10551 6883 10557
rect 7650 10548 7656 10560
rect 7708 10548 7714 10600
rect 8389 10591 8447 10597
rect 8389 10557 8401 10591
rect 8435 10588 8447 10591
rect 8680 10588 8708 10628
rect 9030 10616 9036 10628
rect 9088 10616 9094 10668
rect 10962 10656 10968 10668
rect 9140 10628 10968 10656
rect 8846 10588 8852 10600
rect 8435 10560 8708 10588
rect 8759 10560 8852 10588
rect 8435 10557 8447 10560
rect 8389 10551 8447 10557
rect 8846 10548 8852 10560
rect 8904 10588 8910 10600
rect 9140 10588 9168 10628
rect 10962 10616 10968 10628
rect 11020 10616 11026 10668
rect 11517 10659 11575 10665
rect 11517 10625 11529 10659
rect 11563 10656 11575 10659
rect 11974 10656 11980 10668
rect 11563 10628 11980 10656
rect 11563 10625 11575 10628
rect 11517 10619 11575 10625
rect 11974 10616 11980 10628
rect 12032 10616 12038 10668
rect 12066 10616 12072 10668
rect 12124 10656 12130 10668
rect 12124 10628 13032 10656
rect 12124 10616 12130 10628
rect 13004 10600 13032 10628
rect 13906 10616 13912 10668
rect 13964 10656 13970 10668
rect 14001 10659 14059 10665
rect 14001 10656 14013 10659
rect 13964 10628 14013 10656
rect 13964 10616 13970 10628
rect 14001 10625 14013 10628
rect 14047 10625 14059 10659
rect 17126 10656 17132 10668
rect 17087 10628 17132 10656
rect 14001 10619 14059 10625
rect 17126 10616 17132 10628
rect 17184 10616 17190 10668
rect 17862 10616 17868 10668
rect 17920 10656 17926 10668
rect 18877 10659 18935 10665
rect 18877 10656 18889 10659
rect 17920 10628 18889 10656
rect 17920 10616 17926 10628
rect 18877 10625 18889 10628
rect 18923 10625 18935 10659
rect 20530 10656 20536 10668
rect 18877 10619 18935 10625
rect 19904 10628 20536 10656
rect 9858 10588 9864 10600
rect 8904 10560 9168 10588
rect 9819 10560 9864 10588
rect 8904 10548 8910 10560
rect 9858 10548 9864 10560
rect 9916 10548 9922 10600
rect 10045 10591 10103 10597
rect 10045 10557 10057 10591
rect 10091 10557 10103 10591
rect 11422 10588 11428 10600
rect 11383 10560 11428 10588
rect 10045 10551 10103 10557
rect 3602 10480 3608 10532
rect 3660 10520 3666 10532
rect 3660 10492 7144 10520
rect 3660 10480 3666 10492
rect 1394 10412 1400 10464
rect 1452 10452 1458 10464
rect 3237 10455 3295 10461
rect 3237 10452 3249 10455
rect 1452 10424 3249 10452
rect 1452 10412 1458 10424
rect 3237 10421 3249 10424
rect 3283 10452 3295 10455
rect 3510 10452 3516 10464
rect 3283 10424 3516 10452
rect 3283 10421 3295 10424
rect 3237 10415 3295 10421
rect 3510 10412 3516 10424
rect 3568 10412 3574 10464
rect 7116 10452 7144 10492
rect 8662 10480 8668 10532
rect 8720 10520 8726 10532
rect 10060 10520 10088 10551
rect 11422 10548 11428 10560
rect 11480 10548 11486 10600
rect 11698 10588 11704 10600
rect 11659 10560 11704 10588
rect 11698 10548 11704 10560
rect 11756 10548 11762 10600
rect 12434 10548 12440 10600
rect 12492 10588 12498 10600
rect 12986 10588 12992 10600
rect 12492 10560 12537 10588
rect 12947 10560 12992 10588
rect 12492 10548 12498 10560
rect 12986 10548 12992 10560
rect 13044 10548 13050 10600
rect 13354 10588 13360 10600
rect 13315 10560 13360 10588
rect 13354 10548 13360 10560
rect 13412 10548 13418 10600
rect 13630 10548 13636 10600
rect 13688 10588 13694 10600
rect 14458 10588 14464 10600
rect 13688 10560 14464 10588
rect 13688 10548 13694 10560
rect 14458 10548 14464 10560
rect 14516 10548 14522 10600
rect 14645 10591 14703 10597
rect 14645 10557 14657 10591
rect 14691 10557 14703 10591
rect 14645 10551 14703 10557
rect 14829 10591 14887 10597
rect 14829 10557 14841 10591
rect 14875 10588 14887 10591
rect 15286 10588 15292 10600
rect 14875 10560 15292 10588
rect 14875 10557 14887 10560
rect 14829 10551 14887 10557
rect 8720 10492 10088 10520
rect 10321 10523 10379 10529
rect 8720 10480 8726 10492
rect 10321 10489 10333 10523
rect 10367 10520 10379 10523
rect 12342 10520 12348 10532
rect 10367 10492 12348 10520
rect 10367 10489 10379 10492
rect 10321 10483 10379 10489
rect 12342 10480 12348 10492
rect 12400 10480 12406 10532
rect 12710 10480 12716 10532
rect 12768 10520 12774 10532
rect 14660 10520 14688 10551
rect 15286 10548 15292 10560
rect 15344 10548 15350 10600
rect 15378 10548 15384 10600
rect 15436 10588 15442 10600
rect 15473 10591 15531 10597
rect 15473 10588 15485 10591
rect 15436 10560 15485 10588
rect 15436 10548 15442 10560
rect 15473 10557 15485 10560
rect 15519 10557 15531 10591
rect 15473 10551 15531 10557
rect 16485 10591 16543 10597
rect 16485 10557 16497 10591
rect 16531 10588 16543 10591
rect 16574 10588 16580 10600
rect 16531 10560 16580 10588
rect 16531 10557 16543 10560
rect 16485 10551 16543 10557
rect 16574 10548 16580 10560
rect 16632 10548 16638 10600
rect 16945 10591 17003 10597
rect 16945 10557 16957 10591
rect 16991 10588 17003 10591
rect 17218 10588 17224 10600
rect 16991 10560 17224 10588
rect 16991 10557 17003 10560
rect 16945 10551 17003 10557
rect 17218 10548 17224 10560
rect 17276 10548 17282 10600
rect 17313 10591 17371 10597
rect 17313 10557 17325 10591
rect 17359 10557 17371 10591
rect 17313 10551 17371 10557
rect 18049 10591 18107 10597
rect 18049 10557 18061 10591
rect 18095 10588 18107 10591
rect 18414 10588 18420 10600
rect 18095 10560 18420 10588
rect 18095 10557 18107 10560
rect 18049 10551 18107 10557
rect 12768 10492 14688 10520
rect 17328 10520 17356 10551
rect 18414 10548 18420 10560
rect 18472 10548 18478 10600
rect 19426 10548 19432 10600
rect 19484 10588 19490 10600
rect 19904 10597 19932 10628
rect 20530 10616 20536 10628
rect 20588 10616 20594 10668
rect 21450 10616 21456 10668
rect 21508 10656 21514 10668
rect 21545 10659 21603 10665
rect 21545 10656 21557 10659
rect 21508 10628 21557 10656
rect 21508 10616 21514 10628
rect 21545 10625 21557 10628
rect 21591 10625 21603 10659
rect 22830 10656 22836 10668
rect 21545 10619 21603 10625
rect 22020 10628 22836 10656
rect 19521 10591 19579 10597
rect 19521 10588 19533 10591
rect 19484 10560 19533 10588
rect 19484 10548 19490 10560
rect 19521 10557 19533 10560
rect 19567 10557 19579 10591
rect 19521 10551 19579 10557
rect 19613 10591 19671 10597
rect 19613 10557 19625 10591
rect 19659 10557 19671 10591
rect 19613 10551 19671 10557
rect 19889 10591 19947 10597
rect 19889 10557 19901 10591
rect 19935 10557 19947 10591
rect 19889 10551 19947 10557
rect 20073 10591 20131 10597
rect 20073 10557 20085 10591
rect 20119 10588 20131 10591
rect 20162 10588 20168 10600
rect 20119 10560 20168 10588
rect 20119 10557 20131 10560
rect 20073 10551 20131 10557
rect 17954 10520 17960 10532
rect 17328 10492 17960 10520
rect 12768 10480 12774 10492
rect 17954 10480 17960 10492
rect 18012 10480 18018 10532
rect 19628 10520 19656 10551
rect 20162 10548 20168 10560
rect 20220 10548 20226 10600
rect 21634 10588 21640 10600
rect 21595 10560 21640 10588
rect 21634 10548 21640 10560
rect 21692 10548 21698 10600
rect 22020 10597 22048 10628
rect 22830 10616 22836 10628
rect 22888 10616 22894 10668
rect 24578 10616 24584 10668
rect 24636 10656 24642 10668
rect 24673 10659 24731 10665
rect 24673 10656 24685 10659
rect 24636 10628 24685 10656
rect 24636 10616 24642 10628
rect 24673 10625 24685 10628
rect 24719 10656 24731 10659
rect 25590 10656 25596 10668
rect 24719 10628 25596 10656
rect 24719 10625 24731 10628
rect 24673 10619 24731 10625
rect 25590 10616 25596 10628
rect 25648 10616 25654 10668
rect 27080 10600 27108 10696
rect 29454 10684 29460 10696
rect 29512 10684 29518 10736
rect 31404 10733 31432 10764
rect 38746 10752 38752 10764
rect 38804 10752 38810 10804
rect 31389 10727 31447 10733
rect 29564 10696 30420 10724
rect 28074 10616 28080 10668
rect 28132 10656 28138 10668
rect 29089 10659 29147 10665
rect 29089 10656 29101 10659
rect 28132 10628 29101 10656
rect 28132 10616 28138 10628
rect 29089 10625 29101 10628
rect 29135 10656 29147 10659
rect 29273 10659 29331 10665
rect 29273 10656 29285 10659
rect 29135 10628 29285 10656
rect 29135 10625 29147 10628
rect 29089 10619 29147 10625
rect 29273 10625 29285 10628
rect 29319 10625 29331 10659
rect 29564 10656 29592 10696
rect 29273 10619 29331 10625
rect 29380 10628 29592 10656
rect 30392 10656 30420 10696
rect 31389 10693 31401 10727
rect 31435 10693 31447 10727
rect 37274 10724 37280 10736
rect 31389 10687 31447 10693
rect 36096 10696 37280 10724
rect 30392 10628 31708 10656
rect 22005 10591 22063 10597
rect 22005 10557 22017 10591
rect 22051 10557 22063 10591
rect 22005 10551 22063 10557
rect 22097 10591 22155 10597
rect 22097 10557 22109 10591
rect 22143 10557 22155 10591
rect 22646 10588 22652 10600
rect 22607 10560 22652 10588
rect 22097 10551 22155 10557
rect 19978 10520 19984 10532
rect 19628 10492 19984 10520
rect 19978 10480 19984 10492
rect 20036 10480 20042 10532
rect 21542 10480 21548 10532
rect 21600 10520 21606 10532
rect 22112 10520 22140 10551
rect 22646 10548 22652 10560
rect 22704 10548 22710 10600
rect 23198 10548 23204 10600
rect 23256 10588 23262 10600
rect 23661 10591 23719 10597
rect 23661 10588 23673 10591
rect 23256 10560 23673 10588
rect 23256 10548 23262 10560
rect 23661 10557 23673 10560
rect 23707 10557 23719 10591
rect 24946 10588 24952 10600
rect 24907 10560 24952 10588
rect 23661 10551 23719 10557
rect 24946 10548 24952 10560
rect 25004 10548 25010 10600
rect 27062 10588 27068 10600
rect 26975 10560 27068 10588
rect 27062 10548 27068 10560
rect 27120 10548 27126 10600
rect 27154 10548 27160 10600
rect 27212 10588 27218 10600
rect 27522 10588 27528 10600
rect 27212 10560 27257 10588
rect 27483 10560 27528 10588
rect 27212 10548 27218 10560
rect 27522 10548 27528 10560
rect 27580 10548 27586 10600
rect 27617 10591 27675 10597
rect 27617 10557 27629 10591
rect 27663 10588 27675 10591
rect 27982 10588 27988 10600
rect 27663 10560 27988 10588
rect 27663 10557 27675 10560
rect 27617 10551 27675 10557
rect 27982 10548 27988 10560
rect 28040 10588 28046 10600
rect 28040 10560 28580 10588
rect 28040 10548 28046 10560
rect 21600 10492 22140 10520
rect 22664 10520 22692 10548
rect 23290 10520 23296 10532
rect 22664 10492 23296 10520
rect 21600 10480 21606 10492
rect 22020 10464 22048 10492
rect 23290 10480 23296 10492
rect 23348 10520 23354 10532
rect 23753 10523 23811 10529
rect 23753 10520 23765 10523
rect 23348 10492 23765 10520
rect 23348 10480 23354 10492
rect 23753 10489 23765 10492
rect 23799 10489 23811 10523
rect 23753 10483 23811 10489
rect 26050 10480 26056 10532
rect 26108 10520 26114 10532
rect 28074 10520 28080 10532
rect 26108 10492 28080 10520
rect 26108 10480 26114 10492
rect 28074 10480 28080 10492
rect 28132 10480 28138 10532
rect 28169 10523 28227 10529
rect 28169 10489 28181 10523
rect 28215 10520 28227 10523
rect 28442 10520 28448 10532
rect 28215 10492 28448 10520
rect 28215 10489 28227 10492
rect 28169 10483 28227 10489
rect 28442 10480 28448 10492
rect 28500 10480 28506 10532
rect 28552 10520 28580 10560
rect 28626 10548 28632 10600
rect 28684 10588 28690 10600
rect 29380 10588 29408 10628
rect 28684 10560 29408 10588
rect 28684 10548 28690 10560
rect 29454 10548 29460 10600
rect 29512 10588 29518 10600
rect 30009 10591 30067 10597
rect 29512 10560 29557 10588
rect 29512 10548 29518 10560
rect 30009 10557 30021 10591
rect 30055 10557 30067 10591
rect 30009 10551 30067 10557
rect 30193 10591 30251 10597
rect 30193 10557 30205 10591
rect 30239 10557 30251 10591
rect 30193 10551 30251 10557
rect 31297 10591 31355 10597
rect 31297 10557 31309 10591
rect 31343 10588 31355 10591
rect 31386 10588 31392 10600
rect 31343 10560 31392 10588
rect 31343 10557 31355 10560
rect 31297 10551 31355 10557
rect 30024 10520 30052 10551
rect 28552 10492 30052 10520
rect 30208 10520 30236 10551
rect 31386 10548 31392 10560
rect 31444 10548 31450 10600
rect 31680 10597 31708 10628
rect 35618 10616 35624 10668
rect 35676 10656 35682 10668
rect 36096 10665 36124 10696
rect 37274 10684 37280 10696
rect 37332 10684 37338 10736
rect 36081 10659 36139 10665
rect 36081 10656 36093 10659
rect 35676 10628 36093 10656
rect 35676 10616 35682 10628
rect 36081 10625 36093 10628
rect 36127 10625 36139 10659
rect 36081 10619 36139 10625
rect 36354 10616 36360 10668
rect 36412 10616 36418 10668
rect 37734 10656 37740 10668
rect 37695 10628 37740 10656
rect 37734 10616 37740 10628
rect 37792 10616 37798 10668
rect 37826 10616 37832 10668
rect 37884 10656 37890 10668
rect 38841 10659 38899 10665
rect 38841 10656 38853 10659
rect 37884 10628 38853 10656
rect 37884 10616 37890 10628
rect 38841 10625 38853 10628
rect 38887 10625 38899 10659
rect 38841 10619 38899 10625
rect 31665 10591 31723 10597
rect 31665 10557 31677 10591
rect 31711 10557 31723 10591
rect 31665 10551 31723 10557
rect 31754 10548 31760 10600
rect 31812 10588 31818 10600
rect 32125 10591 32183 10597
rect 32125 10588 32137 10591
rect 31812 10560 32137 10588
rect 31812 10548 31818 10560
rect 32125 10557 32137 10560
rect 32171 10588 32183 10591
rect 32214 10588 32220 10600
rect 32171 10560 32220 10588
rect 32171 10557 32183 10560
rect 32125 10551 32183 10557
rect 32214 10548 32220 10560
rect 32272 10548 32278 10600
rect 32861 10591 32919 10597
rect 32861 10557 32873 10591
rect 32907 10557 32919 10591
rect 33226 10588 33232 10600
rect 33187 10560 33232 10588
rect 32861 10551 32919 10557
rect 31478 10520 31484 10532
rect 30208 10492 31484 10520
rect 12618 10452 12624 10464
rect 7116 10424 12624 10452
rect 12618 10412 12624 10424
rect 12676 10412 12682 10464
rect 13078 10412 13084 10464
rect 13136 10452 13142 10464
rect 13722 10452 13728 10464
rect 13136 10424 13728 10452
rect 13136 10412 13142 10424
rect 13722 10412 13728 10424
rect 13780 10412 13786 10464
rect 14182 10412 14188 10464
rect 14240 10452 14246 10464
rect 15470 10452 15476 10464
rect 14240 10424 15476 10452
rect 14240 10412 14246 10424
rect 15470 10412 15476 10424
rect 15528 10452 15534 10464
rect 15657 10455 15715 10461
rect 15657 10452 15669 10455
rect 15528 10424 15669 10452
rect 15528 10412 15534 10424
rect 15657 10421 15669 10424
rect 15703 10421 15715 10455
rect 15657 10415 15715 10421
rect 16390 10412 16396 10464
rect 16448 10452 16454 10464
rect 18233 10455 18291 10461
rect 18233 10452 18245 10455
rect 16448 10424 18245 10452
rect 16448 10412 16454 10424
rect 18233 10421 18245 10424
rect 18279 10452 18291 10455
rect 19334 10452 19340 10464
rect 18279 10424 19340 10452
rect 18279 10421 18291 10424
rect 18233 10415 18291 10421
rect 19334 10412 19340 10424
rect 19392 10412 19398 10464
rect 22002 10412 22008 10464
rect 22060 10412 22066 10464
rect 22278 10412 22284 10464
rect 22336 10452 22342 10464
rect 22833 10455 22891 10461
rect 22833 10452 22845 10455
rect 22336 10424 22845 10452
rect 22336 10412 22342 10424
rect 22833 10421 22845 10424
rect 22879 10421 22891 10455
rect 22833 10415 22891 10421
rect 26142 10412 26148 10464
rect 26200 10452 26206 10464
rect 26237 10455 26295 10461
rect 26237 10452 26249 10455
rect 26200 10424 26249 10452
rect 26200 10412 26206 10424
rect 26237 10421 26249 10424
rect 26283 10452 26295 10455
rect 27338 10452 27344 10464
rect 26283 10424 27344 10452
rect 26283 10421 26295 10424
rect 26237 10415 26295 10421
rect 27338 10412 27344 10424
rect 27396 10412 27402 10464
rect 27706 10412 27712 10464
rect 27764 10452 27770 10464
rect 30208 10452 30236 10492
rect 31478 10480 31484 10492
rect 31536 10480 31542 10532
rect 32876 10520 32904 10551
rect 33226 10548 33232 10560
rect 33284 10548 33290 10600
rect 33502 10588 33508 10600
rect 33463 10560 33508 10588
rect 33502 10548 33508 10560
rect 33560 10548 33566 10600
rect 33686 10548 33692 10600
rect 33744 10588 33750 10600
rect 34425 10591 34483 10597
rect 34425 10588 34437 10591
rect 33744 10560 34437 10588
rect 33744 10548 33750 10560
rect 34425 10557 34437 10560
rect 34471 10557 34483 10591
rect 34425 10551 34483 10557
rect 35161 10591 35219 10597
rect 35161 10557 35173 10591
rect 35207 10557 35219 10591
rect 36372 10588 36400 10616
rect 36449 10591 36507 10597
rect 36449 10588 36461 10591
rect 36372 10560 36461 10588
rect 35161 10551 35219 10557
rect 36449 10557 36461 10560
rect 36495 10557 36507 10591
rect 36722 10588 36728 10600
rect 36683 10560 36728 10588
rect 36449 10551 36507 10557
rect 35176 10520 35204 10551
rect 36722 10548 36728 10560
rect 36780 10548 36786 10600
rect 37458 10588 37464 10600
rect 37419 10560 37464 10588
rect 37458 10548 37464 10560
rect 37516 10548 37522 10600
rect 36078 10520 36084 10532
rect 32876 10492 33272 10520
rect 35176 10492 36084 10520
rect 33244 10464 33272 10492
rect 36078 10480 36084 10492
rect 36136 10520 36142 10532
rect 36354 10520 36360 10532
rect 36136 10492 36360 10520
rect 36136 10480 36142 10492
rect 36354 10480 36360 10492
rect 36412 10480 36418 10532
rect 37001 10523 37059 10529
rect 37001 10489 37013 10523
rect 37047 10520 37059 10523
rect 37550 10520 37556 10532
rect 37047 10492 37556 10520
rect 37047 10489 37059 10492
rect 37001 10483 37059 10489
rect 37550 10480 37556 10492
rect 37608 10480 37614 10532
rect 30466 10452 30472 10464
rect 27764 10424 30236 10452
rect 30427 10424 30472 10452
rect 27764 10412 27770 10424
rect 30466 10412 30472 10424
rect 30524 10412 30530 10464
rect 32769 10455 32827 10461
rect 32769 10421 32781 10455
rect 32815 10452 32827 10455
rect 33134 10452 33140 10464
rect 32815 10424 33140 10452
rect 32815 10421 32827 10424
rect 32769 10415 32827 10421
rect 33134 10412 33140 10424
rect 33192 10412 33198 10464
rect 33226 10412 33232 10464
rect 33284 10412 33290 10464
rect 34241 10455 34299 10461
rect 34241 10421 34253 10455
rect 34287 10452 34299 10455
rect 34330 10452 34336 10464
rect 34287 10424 34336 10452
rect 34287 10421 34299 10424
rect 34241 10415 34299 10421
rect 34330 10412 34336 10424
rect 34388 10412 34394 10464
rect 34790 10412 34796 10464
rect 34848 10452 34854 10464
rect 35345 10455 35403 10461
rect 35345 10452 35357 10455
rect 34848 10424 35357 10452
rect 34848 10412 34854 10424
rect 35345 10421 35357 10424
rect 35391 10452 35403 10455
rect 38930 10452 38936 10464
rect 35391 10424 38936 10452
rect 35391 10421 35403 10424
rect 35345 10415 35403 10421
rect 38930 10412 38936 10424
rect 38988 10412 38994 10464
rect 1104 10362 39836 10384
rect 1104 10310 19606 10362
rect 19658 10310 19670 10362
rect 19722 10310 19734 10362
rect 19786 10310 19798 10362
rect 19850 10310 39836 10362
rect 1104 10288 39836 10310
rect 4338 10208 4344 10260
rect 4396 10248 4402 10260
rect 5629 10251 5687 10257
rect 5629 10248 5641 10251
rect 4396 10220 5641 10248
rect 4396 10208 4402 10220
rect 5629 10217 5641 10220
rect 5675 10248 5687 10251
rect 7650 10248 7656 10260
rect 5675 10220 7656 10248
rect 5675 10217 5687 10220
rect 5629 10211 5687 10217
rect 7650 10208 7656 10220
rect 7708 10208 7714 10260
rect 13078 10248 13084 10260
rect 7760 10220 13084 10248
rect 5350 10140 5356 10192
rect 5408 10180 5414 10192
rect 7760 10180 7788 10220
rect 13078 10208 13084 10220
rect 13136 10208 13142 10260
rect 13170 10208 13176 10260
rect 13228 10248 13234 10260
rect 13357 10251 13415 10257
rect 13357 10248 13369 10251
rect 13228 10220 13369 10248
rect 13228 10208 13234 10220
rect 13357 10217 13369 10220
rect 13403 10217 13415 10251
rect 13357 10211 13415 10217
rect 13722 10208 13728 10260
rect 13780 10248 13786 10260
rect 13780 10220 21220 10248
rect 13780 10208 13786 10220
rect 5408 10152 7788 10180
rect 11057 10183 11115 10189
rect 5408 10140 5414 10152
rect 11057 10149 11069 10183
rect 11103 10180 11115 10183
rect 12710 10180 12716 10192
rect 11103 10152 12716 10180
rect 11103 10149 11115 10152
rect 11057 10143 11115 10149
rect 12710 10140 12716 10152
rect 12768 10140 12774 10192
rect 12805 10183 12863 10189
rect 12805 10149 12817 10183
rect 12851 10180 12863 10183
rect 15286 10180 15292 10192
rect 12851 10152 14412 10180
rect 15247 10152 15292 10180
rect 12851 10149 12863 10152
rect 12805 10143 12863 10149
rect 1673 10115 1731 10121
rect 1673 10081 1685 10115
rect 1719 10112 1731 10115
rect 2498 10112 2504 10124
rect 1719 10084 2504 10112
rect 1719 10081 1731 10084
rect 1673 10075 1731 10081
rect 2498 10072 2504 10084
rect 2556 10072 2562 10124
rect 4065 10115 4123 10121
rect 4065 10081 4077 10115
rect 4111 10112 4123 10115
rect 4982 10112 4988 10124
rect 4111 10084 4988 10112
rect 4111 10081 4123 10084
rect 4065 10075 4123 10081
rect 4982 10072 4988 10084
rect 5040 10112 5046 10124
rect 5166 10112 5172 10124
rect 5040 10084 5172 10112
rect 5040 10072 5046 10084
rect 5166 10072 5172 10084
rect 5224 10072 5230 10124
rect 6178 10112 6184 10124
rect 6139 10084 6184 10112
rect 6178 10072 6184 10084
rect 6236 10072 6242 10124
rect 6914 10072 6920 10124
rect 6972 10112 6978 10124
rect 7561 10115 7619 10121
rect 7561 10112 7573 10115
rect 6972 10084 7573 10112
rect 6972 10072 6978 10084
rect 7561 10081 7573 10084
rect 7607 10081 7619 10115
rect 7561 10075 7619 10081
rect 8297 10115 8355 10121
rect 8297 10081 8309 10115
rect 8343 10112 8355 10115
rect 8846 10112 8852 10124
rect 8904 10121 8910 10124
rect 8343 10084 8852 10112
rect 8343 10081 8355 10084
rect 8297 10075 8355 10081
rect 8846 10072 8852 10084
rect 8904 10112 8913 10121
rect 10502 10112 10508 10124
rect 8904 10084 8949 10112
rect 10463 10084 10508 10112
rect 8904 10075 8913 10084
rect 8904 10072 8910 10075
rect 10502 10072 10508 10084
rect 10560 10072 10566 10124
rect 10778 10112 10784 10124
rect 10739 10084 10784 10112
rect 10778 10072 10784 10084
rect 10836 10072 10842 10124
rect 12345 10115 12403 10121
rect 12345 10081 12357 10115
rect 12391 10081 12403 10115
rect 12526 10112 12532 10124
rect 12487 10084 12532 10112
rect 12345 10075 12403 10081
rect 1394 10044 1400 10056
rect 1355 10016 1400 10044
rect 1394 10004 1400 10016
rect 1452 10004 1458 10056
rect 2774 10004 2780 10056
rect 2832 10044 2838 10056
rect 4341 10047 4399 10053
rect 2832 10016 2877 10044
rect 2832 10004 2838 10016
rect 4341 10013 4353 10047
rect 4387 10044 4399 10047
rect 4706 10044 4712 10056
rect 4387 10016 4712 10044
rect 4387 10013 4399 10016
rect 4341 10007 4399 10013
rect 4706 10004 4712 10016
rect 4764 10004 4770 10056
rect 7929 10047 7987 10053
rect 7929 10013 7941 10047
rect 7975 10044 7987 10047
rect 8202 10044 8208 10056
rect 7975 10016 8208 10044
rect 7975 10013 7987 10016
rect 7929 10007 7987 10013
rect 8202 10004 8208 10016
rect 8260 10004 8266 10056
rect 8570 10004 8576 10056
rect 8628 10044 8634 10056
rect 9582 10044 9588 10056
rect 8628 10016 9588 10044
rect 8628 10004 8634 10016
rect 9582 10004 9588 10016
rect 9640 10044 9646 10056
rect 10045 10047 10103 10053
rect 10045 10044 10057 10047
rect 9640 10016 10057 10044
rect 9640 10004 9646 10016
rect 10045 10013 10057 10016
rect 10091 10013 10103 10047
rect 12360 10044 12388 10075
rect 12526 10072 12532 10084
rect 12584 10072 12590 10124
rect 13449 10115 13507 10121
rect 13449 10081 13461 10115
rect 13495 10112 13507 10115
rect 13538 10112 13544 10124
rect 13495 10084 13544 10112
rect 13495 10081 13507 10084
rect 13449 10075 13507 10081
rect 13538 10072 13544 10084
rect 13596 10072 13602 10124
rect 13906 10112 13912 10124
rect 13867 10084 13912 10112
rect 13906 10072 13912 10084
rect 13964 10072 13970 10124
rect 14384 10112 14412 10152
rect 15286 10140 15292 10152
rect 15344 10140 15350 10192
rect 15933 10115 15991 10121
rect 15933 10112 15945 10115
rect 14384 10084 15945 10112
rect 15933 10081 15945 10084
rect 15979 10081 15991 10115
rect 15933 10075 15991 10081
rect 16301 10115 16359 10121
rect 16301 10081 16313 10115
rect 16347 10112 16359 10115
rect 16574 10112 16580 10124
rect 16347 10084 16580 10112
rect 16347 10081 16359 10084
rect 16301 10075 16359 10081
rect 16574 10072 16580 10084
rect 16632 10072 16638 10124
rect 17129 10115 17187 10121
rect 17129 10081 17141 10115
rect 17175 10081 17187 10115
rect 17129 10075 17187 10081
rect 14182 10044 14188 10056
rect 12360 10016 14188 10044
rect 10045 10007 10103 10013
rect 14182 10004 14188 10016
rect 14240 10004 14246 10056
rect 14277 10047 14335 10053
rect 14277 10013 14289 10047
rect 14323 10013 14335 10047
rect 14277 10007 14335 10013
rect 9674 9936 9680 9988
rect 9732 9976 9738 9988
rect 12802 9976 12808 9988
rect 9732 9948 12808 9976
rect 9732 9936 9738 9948
rect 12802 9936 12808 9948
rect 12860 9936 12866 9988
rect 14292 9976 14320 10007
rect 15746 10004 15752 10056
rect 15804 10044 15810 10056
rect 15841 10047 15899 10053
rect 15841 10044 15853 10047
rect 15804 10016 15853 10044
rect 15804 10004 15810 10016
rect 15841 10013 15853 10016
rect 15887 10013 15899 10047
rect 16390 10044 16396 10056
rect 16351 10016 16396 10044
rect 15841 10007 15899 10013
rect 16390 10004 16396 10016
rect 16448 10004 16454 10056
rect 16945 10047 17003 10053
rect 16945 10013 16957 10047
rect 16991 10044 17003 10047
rect 17144 10044 17172 10075
rect 17218 10072 17224 10124
rect 17276 10112 17282 10124
rect 17405 10115 17463 10121
rect 17405 10112 17417 10115
rect 17276 10084 17417 10112
rect 17276 10072 17282 10084
rect 17405 10081 17417 10084
rect 17451 10081 17463 10115
rect 17954 10112 17960 10124
rect 17915 10084 17960 10112
rect 17405 10075 17463 10081
rect 17954 10072 17960 10084
rect 18012 10072 18018 10124
rect 18969 10115 19027 10121
rect 18969 10081 18981 10115
rect 19015 10112 19027 10115
rect 19150 10112 19156 10124
rect 19015 10084 19156 10112
rect 19015 10081 19027 10084
rect 18969 10075 19027 10081
rect 19150 10072 19156 10084
rect 19208 10072 19214 10124
rect 19334 10112 19340 10124
rect 19295 10084 19340 10112
rect 19334 10072 19340 10084
rect 19392 10072 19398 10124
rect 19886 10112 19892 10124
rect 19847 10084 19892 10112
rect 19886 10072 19892 10084
rect 19944 10072 19950 10124
rect 18322 10044 18328 10056
rect 16991 10016 18328 10044
rect 16991 10013 17003 10016
rect 16945 10007 17003 10013
rect 18322 10004 18328 10016
rect 18380 10004 18386 10056
rect 20993 9979 21051 9985
rect 20993 9976 21005 9979
rect 14292 9948 21005 9976
rect 20993 9945 21005 9948
rect 21039 9945 21051 9979
rect 20993 9939 21051 9945
rect 5442 9868 5448 9920
rect 5500 9908 5506 9920
rect 6365 9911 6423 9917
rect 6365 9908 6377 9911
rect 5500 9880 6377 9908
rect 5500 9868 5506 9880
rect 6365 9877 6377 9880
rect 6411 9877 6423 9911
rect 6365 9871 6423 9877
rect 9033 9911 9091 9917
rect 9033 9877 9045 9911
rect 9079 9908 9091 9911
rect 10502 9908 10508 9920
rect 9079 9880 10508 9908
rect 9079 9877 9091 9880
rect 9033 9871 9091 9877
rect 10502 9868 10508 9880
rect 10560 9908 10566 9920
rect 12066 9908 12072 9920
rect 10560 9880 12072 9908
rect 10560 9868 10566 9880
rect 12066 9868 12072 9880
rect 12124 9868 12130 9920
rect 12710 9868 12716 9920
rect 12768 9908 12774 9920
rect 16945 9911 17003 9917
rect 16945 9908 16957 9911
rect 12768 9880 16957 9908
rect 12768 9868 12774 9880
rect 16945 9877 16957 9880
rect 16991 9877 17003 9911
rect 16945 9871 17003 9877
rect 17129 9911 17187 9917
rect 17129 9877 17141 9911
rect 17175 9908 17187 9911
rect 17218 9908 17224 9920
rect 17175 9880 17224 9908
rect 17175 9877 17187 9880
rect 17129 9871 17187 9877
rect 17218 9868 17224 9880
rect 17276 9868 17282 9920
rect 18414 9868 18420 9920
rect 18472 9908 18478 9920
rect 18785 9911 18843 9917
rect 18785 9908 18797 9911
rect 18472 9880 18797 9908
rect 18472 9868 18478 9880
rect 18785 9877 18797 9880
rect 18831 9877 18843 9911
rect 18785 9871 18843 9877
rect 19978 9868 19984 9920
rect 20036 9908 20042 9920
rect 20073 9911 20131 9917
rect 20073 9908 20085 9911
rect 20036 9880 20085 9908
rect 20036 9868 20042 9880
rect 20073 9877 20085 9880
rect 20119 9877 20131 9911
rect 21192 9908 21220 10220
rect 22830 10208 22836 10260
rect 22888 10248 22894 10260
rect 24121 10251 24179 10257
rect 24121 10248 24133 10251
rect 22888 10220 24133 10248
rect 22888 10208 22894 10220
rect 24121 10217 24133 10220
rect 24167 10217 24179 10251
rect 24121 10211 24179 10217
rect 24210 10208 24216 10260
rect 24268 10248 24274 10260
rect 27154 10248 27160 10260
rect 24268 10220 27160 10248
rect 24268 10208 24274 10220
rect 27154 10208 27160 10220
rect 27212 10208 27218 10260
rect 27614 10248 27620 10260
rect 27575 10220 27620 10248
rect 27614 10208 27620 10220
rect 27672 10208 27678 10260
rect 30374 10248 30380 10260
rect 27724 10220 30380 10248
rect 23750 10140 23756 10192
rect 23808 10180 23814 10192
rect 24228 10180 24256 10208
rect 23808 10152 24256 10180
rect 23808 10140 23814 10152
rect 25314 10140 25320 10192
rect 25372 10180 25378 10192
rect 25372 10152 26556 10180
rect 25372 10140 25378 10152
rect 21542 10112 21548 10124
rect 21503 10084 21548 10112
rect 21542 10072 21548 10084
rect 21600 10072 21606 10124
rect 21910 10112 21916 10124
rect 21871 10084 21916 10112
rect 21910 10072 21916 10084
rect 21968 10072 21974 10124
rect 23382 10072 23388 10124
rect 23440 10112 23446 10124
rect 23440 10084 24440 10112
rect 23440 10072 23446 10084
rect 21450 10044 21456 10056
rect 21411 10016 21456 10044
rect 21450 10004 21456 10016
rect 21508 10004 21514 10056
rect 22002 10044 22008 10056
rect 21963 10016 22008 10044
rect 22002 10004 22008 10016
rect 22060 10004 22066 10056
rect 22738 10044 22744 10056
rect 22699 10016 22744 10044
rect 22738 10004 22744 10016
rect 22796 10004 22802 10056
rect 23017 10047 23075 10053
rect 23017 10013 23029 10047
rect 23063 10044 23075 10047
rect 24412 10044 24440 10084
rect 24854 10072 24860 10124
rect 24912 10112 24918 10124
rect 25225 10115 25283 10121
rect 25225 10112 25237 10115
rect 24912 10084 25237 10112
rect 24912 10072 24918 10084
rect 25225 10081 25237 10084
rect 25271 10081 25283 10115
rect 25682 10112 25688 10124
rect 25643 10084 25688 10112
rect 25225 10075 25283 10081
rect 25682 10072 25688 10084
rect 25740 10072 25746 10124
rect 26528 10121 26556 10152
rect 27246 10140 27252 10192
rect 27304 10180 27310 10192
rect 27724 10180 27752 10220
rect 30374 10208 30380 10220
rect 30432 10208 30438 10260
rect 30561 10251 30619 10257
rect 30561 10217 30573 10251
rect 30607 10248 30619 10251
rect 31294 10248 31300 10260
rect 30607 10220 31300 10248
rect 30607 10217 30619 10220
rect 30561 10211 30619 10217
rect 31294 10208 31300 10220
rect 31352 10208 31358 10260
rect 32217 10251 32275 10257
rect 32217 10217 32229 10251
rect 32263 10248 32275 10251
rect 33502 10248 33508 10260
rect 32263 10220 33508 10248
rect 32263 10217 32275 10220
rect 32217 10211 32275 10217
rect 33502 10208 33508 10220
rect 33560 10208 33566 10260
rect 34793 10251 34851 10257
rect 34793 10217 34805 10251
rect 34839 10248 34851 10251
rect 37093 10251 37151 10257
rect 34839 10220 36216 10248
rect 34839 10217 34851 10220
rect 34793 10211 34851 10217
rect 36188 10180 36216 10220
rect 37093 10217 37105 10251
rect 37139 10248 37151 10251
rect 37274 10248 37280 10260
rect 37139 10220 37280 10248
rect 37139 10217 37151 10220
rect 37093 10211 37151 10217
rect 37274 10208 37280 10220
rect 37332 10208 37338 10260
rect 37366 10208 37372 10260
rect 37424 10248 37430 10260
rect 37829 10251 37887 10257
rect 37829 10248 37841 10251
rect 37424 10220 37841 10248
rect 37424 10208 37430 10220
rect 37829 10217 37841 10220
rect 37875 10217 37887 10251
rect 37829 10211 37887 10217
rect 27304 10152 27752 10180
rect 30668 10152 36124 10180
rect 36188 10152 38240 10180
rect 27304 10140 27310 10152
rect 26513 10115 26571 10121
rect 26513 10081 26525 10115
rect 26559 10081 26571 10115
rect 26513 10075 26571 10081
rect 27525 10115 27583 10121
rect 27525 10081 27537 10115
rect 27571 10112 27583 10115
rect 28442 10112 28448 10124
rect 27571 10084 28304 10112
rect 28403 10084 28448 10112
rect 27571 10081 27583 10084
rect 27525 10075 27583 10081
rect 24949 10047 25007 10053
rect 24949 10044 24961 10047
rect 23063 10016 24348 10044
rect 24412 10016 24961 10044
rect 23063 10013 23075 10016
rect 23017 10007 23075 10013
rect 21266 9936 21272 9988
rect 21324 9976 21330 9988
rect 22756 9976 22784 10004
rect 21324 9948 22784 9976
rect 24320 9976 24348 10016
rect 24949 10013 24961 10016
rect 24995 10013 25007 10047
rect 24949 10007 25007 10013
rect 27154 10004 27160 10056
rect 27212 10044 27218 10056
rect 27890 10044 27896 10056
rect 27212 10016 27896 10044
rect 27212 10004 27218 10016
rect 27890 10004 27896 10016
rect 27948 10004 27954 10056
rect 27982 10004 27988 10056
rect 28040 10044 28046 10056
rect 28169 10047 28227 10053
rect 28169 10044 28181 10047
rect 28040 10016 28181 10044
rect 28040 10004 28046 10016
rect 28169 10013 28181 10016
rect 28215 10013 28227 10047
rect 28276 10044 28304 10084
rect 28442 10072 28448 10084
rect 28500 10072 28506 10124
rect 30558 10112 30564 10124
rect 30519 10084 30564 10112
rect 30558 10072 30564 10084
rect 30616 10072 30622 10124
rect 30668 10056 30696 10152
rect 30834 10072 30840 10124
rect 30892 10112 30898 10124
rect 31021 10115 31079 10121
rect 31021 10112 31033 10115
rect 30892 10084 31033 10112
rect 30892 10072 30898 10084
rect 31021 10081 31033 10084
rect 31067 10081 31079 10115
rect 31021 10075 31079 10081
rect 31110 10072 31116 10124
rect 31168 10112 31174 10124
rect 31297 10115 31355 10121
rect 31297 10112 31309 10115
rect 31168 10084 31309 10112
rect 31168 10072 31174 10084
rect 31297 10081 31309 10084
rect 31343 10081 31355 10115
rect 31297 10075 31355 10081
rect 30650 10044 30656 10056
rect 28276 10016 30656 10044
rect 28169 10007 28227 10013
rect 30650 10004 30656 10016
rect 30708 10004 30714 10056
rect 31312 10044 31340 10075
rect 32306 10072 32312 10124
rect 32364 10112 32370 10124
rect 32674 10112 32680 10124
rect 32364 10084 32409 10112
rect 32635 10084 32680 10112
rect 32364 10072 32370 10084
rect 32674 10072 32680 10084
rect 32732 10072 32738 10124
rect 32766 10072 32772 10124
rect 32824 10112 32830 10124
rect 33689 10115 33747 10121
rect 33689 10112 33701 10115
rect 32824 10084 33701 10112
rect 32824 10072 32830 10084
rect 33689 10081 33701 10084
rect 33735 10112 33747 10115
rect 33778 10112 33784 10124
rect 33735 10084 33784 10112
rect 33735 10081 33747 10084
rect 33689 10075 33747 10081
rect 33778 10072 33784 10084
rect 33836 10072 33842 10124
rect 34793 10115 34851 10121
rect 34793 10081 34805 10115
rect 34839 10112 34851 10115
rect 34885 10115 34943 10121
rect 34885 10112 34897 10115
rect 34839 10084 34897 10112
rect 34839 10081 34851 10084
rect 34793 10075 34851 10081
rect 34885 10081 34897 10084
rect 34931 10081 34943 10115
rect 35618 10112 35624 10124
rect 35579 10084 35624 10112
rect 34885 10075 34943 10081
rect 35618 10072 35624 10084
rect 35676 10072 35682 10124
rect 35802 10112 35808 10124
rect 35763 10084 35808 10112
rect 35802 10072 35808 10084
rect 35860 10072 35866 10124
rect 36096 10121 36124 10152
rect 36081 10115 36139 10121
rect 36081 10081 36093 10115
rect 36127 10081 36139 10115
rect 36081 10075 36139 10081
rect 36909 10115 36967 10121
rect 36909 10081 36921 10115
rect 36955 10112 36967 10115
rect 38010 10112 38016 10124
rect 36955 10084 38016 10112
rect 36955 10081 36967 10084
rect 36909 10075 36967 10081
rect 38010 10072 38016 10084
rect 38068 10072 38074 10124
rect 38212 10121 38240 10152
rect 38197 10115 38255 10121
rect 38197 10081 38209 10115
rect 38243 10081 38255 10115
rect 38930 10112 38936 10124
rect 38891 10084 38936 10112
rect 38197 10075 38255 10081
rect 38930 10072 38936 10084
rect 38988 10072 38994 10124
rect 32953 10047 33011 10053
rect 32953 10044 32965 10047
rect 31312 10016 32965 10044
rect 32953 10013 32965 10016
rect 32999 10013 33011 10047
rect 32953 10007 33011 10013
rect 35345 10047 35403 10053
rect 35345 10013 35357 10047
rect 35391 10044 35403 10047
rect 36446 10044 36452 10056
rect 35391 10016 36452 10044
rect 35391 10013 35403 10016
rect 35345 10007 35403 10013
rect 36446 10004 36452 10016
rect 36504 10004 36510 10056
rect 25685 9979 25743 9985
rect 25685 9976 25697 9979
rect 24320 9948 25697 9976
rect 21324 9936 21330 9948
rect 25685 9945 25697 9948
rect 25731 9945 25743 9979
rect 25685 9939 25743 9945
rect 26697 9979 26755 9985
rect 26697 9945 26709 9979
rect 26743 9976 26755 9979
rect 27522 9976 27528 9988
rect 26743 9948 27528 9976
rect 26743 9945 26755 9948
rect 26697 9939 26755 9945
rect 27522 9936 27528 9948
rect 27580 9976 27586 9988
rect 28074 9976 28080 9988
rect 27580 9948 28080 9976
rect 27580 9936 27586 9948
rect 28074 9936 28080 9948
rect 28132 9936 28138 9988
rect 29362 9936 29368 9988
rect 29420 9976 29426 9988
rect 29420 9948 30236 9976
rect 29420 9936 29426 9948
rect 24670 9908 24676 9920
rect 21192 9880 24676 9908
rect 20073 9871 20131 9877
rect 24670 9868 24676 9880
rect 24728 9868 24734 9920
rect 28166 9868 28172 9920
rect 28224 9908 28230 9920
rect 28626 9908 28632 9920
rect 28224 9880 28632 9908
rect 28224 9868 28230 9880
rect 28626 9868 28632 9880
rect 28684 9868 28690 9920
rect 29733 9911 29791 9917
rect 29733 9877 29745 9911
rect 29779 9908 29791 9911
rect 30098 9908 30104 9920
rect 29779 9880 30104 9908
rect 29779 9877 29791 9880
rect 29733 9871 29791 9877
rect 30098 9868 30104 9880
rect 30156 9868 30162 9920
rect 30208 9908 30236 9948
rect 30558 9936 30564 9988
rect 30616 9976 30622 9988
rect 31386 9976 31392 9988
rect 30616 9948 31392 9976
rect 30616 9936 30622 9948
rect 31386 9936 31392 9948
rect 31444 9976 31450 9988
rect 32306 9976 32312 9988
rect 31444 9948 32312 9976
rect 31444 9936 31450 9948
rect 32306 9936 32312 9948
rect 32364 9976 32370 9988
rect 33873 9979 33931 9985
rect 33873 9976 33885 9979
rect 32364 9948 33885 9976
rect 32364 9936 32370 9948
rect 33873 9945 33885 9948
rect 33919 9945 33931 9979
rect 33873 9939 33931 9945
rect 35802 9936 35808 9988
rect 35860 9976 35866 9988
rect 39025 9979 39083 9985
rect 39025 9976 39037 9979
rect 35860 9948 39037 9976
rect 35860 9936 35866 9948
rect 39025 9945 39037 9948
rect 39071 9945 39083 9979
rect 39025 9939 39083 9945
rect 34793 9911 34851 9917
rect 34793 9908 34805 9911
rect 30208 9880 34805 9908
rect 34793 9877 34805 9880
rect 34839 9877 34851 9911
rect 34793 9871 34851 9877
rect 1104 9818 39836 9840
rect 1104 9766 4246 9818
rect 4298 9766 4310 9818
rect 4362 9766 4374 9818
rect 4426 9766 4438 9818
rect 4490 9766 34966 9818
rect 35018 9766 35030 9818
rect 35082 9766 35094 9818
rect 35146 9766 35158 9818
rect 35210 9766 39836 9818
rect 1104 9744 39836 9766
rect 19981 9707 20039 9713
rect 19981 9673 19993 9707
rect 20027 9704 20039 9707
rect 20162 9704 20168 9716
rect 20027 9676 20168 9704
rect 20027 9673 20039 9676
rect 19981 9667 20039 9673
rect 20162 9664 20168 9676
rect 20220 9664 20226 9716
rect 22738 9664 22744 9716
rect 22796 9704 22802 9716
rect 24578 9704 24584 9716
rect 22796 9676 24584 9704
rect 22796 9664 22802 9676
rect 24578 9664 24584 9676
rect 24636 9664 24642 9716
rect 24872 9676 25268 9704
rect 4062 9596 4068 9648
rect 4120 9636 4126 9648
rect 4614 9636 4620 9648
rect 4120 9608 4620 9636
rect 4120 9596 4126 9608
rect 4614 9596 4620 9608
rect 4672 9596 4678 9648
rect 10229 9639 10287 9645
rect 10229 9605 10241 9639
rect 10275 9636 10287 9639
rect 10778 9636 10784 9648
rect 10275 9608 10784 9636
rect 10275 9605 10287 9608
rect 10229 9599 10287 9605
rect 10778 9596 10784 9608
rect 10836 9596 10842 9648
rect 12802 9636 12808 9648
rect 12763 9608 12808 9636
rect 12802 9596 12808 9608
rect 12860 9596 12866 9648
rect 13630 9636 13636 9648
rect 13591 9608 13636 9636
rect 13630 9596 13636 9608
rect 13688 9596 13694 9648
rect 14458 9596 14464 9648
rect 14516 9636 14522 9648
rect 17402 9636 17408 9648
rect 14516 9608 15424 9636
rect 14516 9596 14522 9608
rect 4249 9571 4307 9577
rect 4249 9537 4261 9571
rect 4295 9568 4307 9571
rect 4706 9568 4712 9580
rect 4295 9540 4712 9568
rect 4295 9537 4307 9540
rect 4249 9531 4307 9537
rect 4706 9528 4712 9540
rect 4764 9528 4770 9580
rect 4816 9540 7696 9568
rect 2314 9500 2320 9512
rect 2275 9472 2320 9500
rect 2314 9460 2320 9472
rect 2372 9460 2378 9512
rect 2777 9503 2835 9509
rect 2777 9469 2789 9503
rect 2823 9469 2835 9503
rect 2777 9463 2835 9469
rect 3605 9503 3663 9509
rect 3605 9469 3617 9503
rect 3651 9469 3663 9503
rect 3878 9500 3884 9512
rect 3839 9472 3884 9500
rect 3605 9463 3663 9469
rect 1670 9324 1676 9376
rect 1728 9364 1734 9376
rect 2317 9367 2375 9373
rect 2317 9364 2329 9367
rect 1728 9336 2329 9364
rect 1728 9324 1734 9336
rect 2317 9333 2329 9336
rect 2363 9333 2375 9367
rect 2792 9364 2820 9463
rect 3620 9432 3648 9463
rect 3878 9460 3884 9472
rect 3936 9460 3942 9512
rect 4816 9509 4844 9540
rect 4341 9503 4399 9509
rect 4341 9469 4353 9503
rect 4387 9500 4399 9503
rect 4801 9503 4859 9509
rect 4387 9472 4568 9500
rect 4387 9469 4399 9472
rect 4341 9463 4399 9469
rect 4430 9432 4436 9444
rect 3620 9404 4436 9432
rect 4430 9392 4436 9404
rect 4488 9392 4494 9444
rect 4540 9432 4568 9472
rect 4801 9469 4813 9503
rect 4847 9469 4859 9503
rect 4801 9463 4859 9469
rect 5353 9503 5411 9509
rect 5353 9469 5365 9503
rect 5399 9469 5411 9503
rect 5353 9463 5411 9469
rect 5813 9503 5871 9509
rect 5813 9469 5825 9503
rect 5859 9500 5871 9503
rect 7009 9503 7067 9509
rect 5859 9472 6408 9500
rect 5859 9469 5871 9472
rect 5813 9463 5871 9469
rect 5166 9432 5172 9444
rect 4540 9404 5172 9432
rect 5166 9392 5172 9404
rect 5224 9392 5230 9444
rect 5368 9432 5396 9463
rect 6086 9432 6092 9444
rect 5368 9404 6092 9432
rect 6086 9392 6092 9404
rect 6144 9392 6150 9444
rect 4154 9364 4160 9376
rect 2792 9336 4160 9364
rect 2317 9327 2375 9333
rect 4154 9324 4160 9336
rect 4212 9324 4218 9376
rect 4890 9324 4896 9376
rect 4948 9364 4954 9376
rect 5905 9367 5963 9373
rect 5905 9364 5917 9367
rect 4948 9336 5917 9364
rect 4948 9324 4954 9336
rect 5905 9333 5917 9336
rect 5951 9333 5963 9367
rect 5905 9327 5963 9333
rect 6178 9324 6184 9376
rect 6236 9364 6242 9376
rect 6380 9364 6408 9472
rect 7009 9469 7021 9503
rect 7055 9469 7067 9503
rect 7282 9500 7288 9512
rect 7243 9472 7288 9500
rect 7009 9463 7067 9469
rect 6454 9392 6460 9444
rect 6512 9432 6518 9444
rect 7024 9432 7052 9463
rect 7282 9460 7288 9472
rect 7340 9460 7346 9512
rect 7668 9500 7696 9540
rect 7742 9528 7748 9580
rect 7800 9568 7806 9580
rect 9217 9571 9275 9577
rect 9217 9568 9229 9571
rect 7800 9540 9229 9568
rect 7800 9528 7806 9540
rect 9217 9537 9229 9540
rect 9263 9568 9275 9571
rect 12526 9568 12532 9580
rect 9263 9540 12532 9568
rect 9263 9537 9275 9540
rect 9217 9531 9275 9537
rect 12526 9528 12532 9540
rect 12584 9528 12590 9580
rect 8665 9503 8723 9509
rect 7668 9472 8524 9500
rect 6512 9404 7052 9432
rect 8496 9432 8524 9472
rect 8665 9469 8677 9503
rect 8711 9500 8723 9503
rect 9125 9503 9183 9509
rect 9125 9500 9137 9503
rect 8711 9472 9137 9500
rect 8711 9469 8723 9472
rect 8665 9463 8723 9469
rect 9125 9469 9137 9472
rect 9171 9469 9183 9503
rect 9950 9500 9956 9512
rect 9911 9472 9956 9500
rect 9125 9463 9183 9469
rect 9950 9460 9956 9472
rect 10008 9460 10014 9512
rect 10689 9503 10747 9509
rect 10689 9469 10701 9503
rect 10735 9469 10747 9503
rect 10689 9463 10747 9469
rect 8754 9432 8760 9444
rect 8496 9404 8760 9432
rect 6512 9392 6518 9404
rect 8754 9392 8760 9404
rect 8812 9392 8818 9444
rect 10594 9364 10600 9376
rect 6236 9336 10600 9364
rect 6236 9324 6242 9336
rect 10594 9324 10600 9336
rect 10652 9324 10658 9376
rect 10704 9364 10732 9463
rect 10778 9460 10784 9512
rect 10836 9500 10842 9512
rect 10836 9472 10881 9500
rect 10836 9460 10842 9472
rect 10962 9460 10968 9512
rect 11020 9500 11026 9512
rect 11517 9503 11575 9509
rect 11517 9500 11529 9503
rect 11020 9472 11529 9500
rect 11020 9460 11026 9472
rect 11517 9469 11529 9472
rect 11563 9469 11575 9503
rect 11517 9463 11575 9469
rect 12250 9460 12256 9512
rect 12308 9500 12314 9512
rect 12621 9503 12679 9509
rect 12621 9500 12633 9503
rect 12308 9472 12633 9500
rect 12308 9460 12314 9472
rect 12621 9469 12633 9472
rect 12667 9500 12679 9503
rect 13262 9500 13268 9512
rect 12667 9472 13268 9500
rect 12667 9469 12679 9472
rect 12621 9463 12679 9469
rect 13262 9460 13268 9472
rect 13320 9460 13326 9512
rect 13538 9500 13544 9512
rect 13499 9472 13544 9500
rect 13538 9460 13544 9472
rect 13596 9460 13602 9512
rect 15396 9509 15424 9608
rect 16592 9608 17408 9636
rect 16592 9577 16620 9608
rect 17402 9596 17408 9608
rect 17460 9596 17466 9648
rect 18509 9639 18567 9645
rect 18509 9605 18521 9639
rect 18555 9636 18567 9639
rect 18598 9636 18604 9648
rect 18555 9608 18604 9636
rect 18555 9605 18567 9608
rect 18509 9599 18567 9605
rect 18598 9596 18604 9608
rect 18656 9596 18662 9648
rect 20180 9636 20208 9664
rect 22002 9636 22008 9648
rect 20180 9608 22008 9636
rect 16577 9571 16635 9577
rect 16577 9537 16589 9571
rect 16623 9537 16635 9571
rect 17310 9568 17316 9580
rect 17271 9540 17316 9568
rect 16577 9531 16635 9537
rect 17310 9528 17316 9540
rect 17368 9528 17374 9580
rect 19245 9571 19303 9577
rect 19245 9537 19257 9571
rect 19291 9568 19303 9571
rect 19978 9568 19984 9580
rect 19291 9540 19984 9568
rect 19291 9537 19303 9540
rect 19245 9531 19303 9537
rect 19978 9528 19984 9540
rect 20036 9568 20042 9580
rect 21177 9571 21235 9577
rect 21177 9568 21189 9571
rect 20036 9540 21189 9568
rect 20036 9528 20042 9540
rect 21177 9537 21189 9540
rect 21223 9568 21235 9571
rect 21450 9568 21456 9580
rect 21223 9540 21456 9568
rect 21223 9537 21235 9540
rect 21177 9531 21235 9537
rect 21450 9528 21456 9540
rect 21508 9528 21514 9580
rect 21744 9577 21772 9608
rect 22002 9596 22008 9608
rect 22060 9596 22066 9648
rect 23290 9596 23296 9648
rect 23348 9636 23354 9648
rect 24872 9636 24900 9676
rect 23348 9608 24900 9636
rect 23348 9596 23354 9608
rect 24946 9596 24952 9648
rect 25004 9636 25010 9648
rect 25133 9639 25191 9645
rect 25133 9636 25145 9639
rect 25004 9608 25145 9636
rect 25004 9596 25010 9608
rect 25133 9605 25145 9608
rect 25179 9605 25191 9639
rect 25133 9599 25191 9605
rect 21729 9571 21787 9577
rect 21729 9537 21741 9571
rect 21775 9537 21787 9571
rect 25240 9568 25268 9676
rect 27430 9664 27436 9716
rect 27488 9704 27494 9716
rect 30190 9704 30196 9716
rect 27488 9676 30196 9704
rect 27488 9664 27494 9676
rect 30190 9664 30196 9676
rect 30248 9664 30254 9716
rect 30374 9664 30380 9716
rect 30432 9704 30438 9716
rect 31846 9704 31852 9716
rect 30432 9676 31852 9704
rect 30432 9664 30438 9676
rect 31846 9664 31852 9676
rect 31904 9704 31910 9716
rect 32674 9704 32680 9716
rect 31904 9676 32680 9704
rect 31904 9664 31910 9676
rect 32674 9664 32680 9676
rect 32732 9664 32738 9716
rect 33778 9664 33784 9716
rect 33836 9704 33842 9716
rect 35710 9704 35716 9716
rect 33836 9676 35716 9704
rect 33836 9664 33842 9676
rect 35710 9664 35716 9676
rect 35768 9664 35774 9716
rect 38010 9664 38016 9716
rect 38068 9704 38074 9716
rect 38289 9707 38347 9713
rect 38289 9704 38301 9707
rect 38068 9676 38301 9704
rect 38068 9664 38074 9676
rect 38289 9673 38301 9676
rect 38335 9673 38347 9707
rect 38289 9667 38347 9673
rect 26053 9639 26111 9645
rect 26053 9605 26065 9639
rect 26099 9636 26111 9639
rect 26234 9636 26240 9648
rect 26099 9608 26240 9636
rect 26099 9605 26111 9608
rect 26053 9599 26111 9605
rect 26234 9596 26240 9608
rect 26292 9636 26298 9648
rect 27062 9636 27068 9648
rect 26292 9608 27068 9636
rect 26292 9596 26298 9608
rect 27062 9596 27068 9608
rect 27120 9596 27126 9648
rect 28994 9636 29000 9648
rect 27172 9608 29000 9636
rect 26881 9571 26939 9577
rect 26881 9568 26893 9571
rect 21729 9531 21787 9537
rect 24136 9540 24348 9568
rect 25240 9540 26893 9568
rect 14093 9503 14151 9509
rect 14093 9469 14105 9503
rect 14139 9469 14151 9503
rect 14093 9463 14151 9469
rect 14369 9503 14427 9509
rect 14369 9469 14381 9503
rect 14415 9500 14427 9503
rect 15381 9503 15439 9509
rect 14415 9472 15332 9500
rect 14415 9469 14427 9472
rect 14369 9463 14427 9469
rect 13722 9432 13728 9444
rect 12452 9404 13728 9432
rect 12452 9376 12480 9404
rect 13722 9392 13728 9404
rect 13780 9392 13786 9444
rect 14108 9432 14136 9463
rect 14921 9435 14979 9441
rect 14921 9432 14933 9435
rect 14108 9404 14933 9432
rect 14921 9401 14933 9404
rect 14967 9401 14979 9435
rect 15304 9432 15332 9472
rect 15381 9469 15393 9503
rect 15427 9469 15439 9503
rect 15562 9500 15568 9512
rect 15523 9472 15568 9500
rect 15381 9463 15439 9469
rect 15562 9460 15568 9472
rect 15620 9460 15626 9512
rect 15654 9460 15660 9512
rect 15712 9500 15718 9512
rect 15749 9503 15807 9509
rect 15749 9500 15761 9503
rect 15712 9472 15761 9500
rect 15712 9460 15718 9472
rect 15749 9469 15761 9472
rect 15795 9469 15807 9503
rect 15749 9463 15807 9469
rect 16666 9460 16672 9512
rect 16724 9500 16730 9512
rect 16761 9503 16819 9509
rect 16761 9500 16773 9503
rect 16724 9472 16773 9500
rect 16724 9460 16730 9472
rect 16761 9469 16773 9472
rect 16807 9469 16819 9503
rect 17218 9500 17224 9512
rect 17179 9472 17224 9500
rect 16761 9463 16819 9469
rect 17218 9460 17224 9472
rect 17276 9460 17282 9512
rect 18414 9500 18420 9512
rect 18375 9472 18420 9500
rect 18414 9460 18420 9472
rect 18472 9460 18478 9512
rect 18782 9500 18788 9512
rect 18743 9472 18788 9500
rect 18782 9460 18788 9472
rect 18840 9460 18846 9512
rect 19058 9460 19064 9512
rect 19116 9500 19122 9512
rect 19797 9503 19855 9509
rect 19797 9500 19809 9503
rect 19116 9472 19809 9500
rect 19116 9460 19122 9472
rect 19797 9469 19809 9472
rect 19843 9469 19855 9503
rect 19797 9463 19855 9469
rect 21269 9503 21327 9509
rect 21269 9469 21281 9503
rect 21315 9469 21327 9503
rect 21634 9500 21640 9512
rect 21595 9472 21640 9500
rect 21269 9463 21327 9469
rect 20625 9435 20683 9441
rect 20625 9432 20637 9435
rect 15304 9404 20637 9432
rect 14921 9395 14979 9401
rect 20625 9401 20637 9404
rect 20671 9401 20683 9435
rect 21284 9432 21312 9463
rect 21634 9460 21640 9472
rect 21692 9460 21698 9512
rect 21818 9460 21824 9512
rect 21876 9500 21882 9512
rect 22281 9503 22339 9509
rect 22281 9500 22293 9503
rect 21876 9472 22293 9500
rect 21876 9460 21882 9472
rect 22281 9469 22293 9472
rect 22327 9469 22339 9503
rect 22830 9500 22836 9512
rect 22791 9472 22836 9500
rect 22281 9463 22339 9469
rect 22830 9460 22836 9472
rect 22888 9460 22894 9512
rect 23106 9460 23112 9512
rect 23164 9500 23170 9512
rect 23658 9500 23664 9512
rect 23164 9472 23664 9500
rect 23164 9460 23170 9472
rect 23658 9460 23664 9472
rect 23716 9500 23722 9512
rect 24029 9503 24087 9509
rect 24029 9500 24041 9503
rect 23716 9472 24041 9500
rect 23716 9460 23722 9472
rect 24029 9469 24041 9472
rect 24075 9469 24087 9503
rect 24029 9463 24087 9469
rect 21284 9404 22416 9432
rect 20625 9395 20683 9401
rect 11701 9367 11759 9373
rect 11701 9364 11713 9367
rect 10704 9336 11713 9364
rect 11701 9333 11713 9336
rect 11747 9364 11759 9367
rect 12434 9364 12440 9376
rect 11747 9336 12440 9364
rect 11747 9333 11759 9336
rect 11701 9327 11759 9333
rect 12434 9324 12440 9336
rect 12492 9324 12498 9376
rect 12802 9324 12808 9376
rect 12860 9364 12866 9376
rect 15746 9364 15752 9376
rect 12860 9336 15752 9364
rect 12860 9324 12866 9336
rect 15746 9324 15752 9336
rect 15804 9364 15810 9376
rect 16022 9364 16028 9376
rect 15804 9336 16028 9364
rect 15804 9324 15810 9336
rect 16022 9324 16028 9336
rect 16080 9324 16086 9376
rect 20990 9324 20996 9376
rect 21048 9364 21054 9376
rect 21818 9364 21824 9376
rect 21048 9336 21824 9364
rect 21048 9324 21054 9336
rect 21818 9324 21824 9336
rect 21876 9324 21882 9376
rect 22388 9373 22416 9404
rect 22373 9367 22431 9373
rect 22373 9333 22385 9367
rect 22419 9333 22431 9367
rect 22373 9327 22431 9333
rect 24026 9324 24032 9376
rect 24084 9364 24090 9376
rect 24136 9364 24164 9540
rect 24213 9503 24271 9509
rect 24213 9469 24225 9503
rect 24259 9469 24271 9503
rect 24320 9500 24348 9540
rect 26881 9537 26893 9540
rect 26927 9568 26939 9571
rect 27172 9568 27200 9608
rect 28994 9596 29000 9608
rect 29052 9596 29058 9648
rect 30650 9636 30656 9648
rect 30611 9608 30656 9636
rect 30650 9596 30656 9608
rect 30708 9596 30714 9648
rect 34054 9596 34060 9648
rect 34112 9596 34118 9648
rect 34330 9596 34336 9648
rect 34388 9636 34394 9648
rect 34388 9608 36952 9636
rect 34388 9596 34394 9608
rect 29549 9571 29607 9577
rect 26927 9540 27200 9568
rect 28000 9540 29408 9568
rect 26927 9537 26939 9540
rect 26881 9531 26939 9537
rect 24673 9503 24731 9509
rect 24673 9500 24685 9503
rect 24320 9472 24685 9500
rect 24213 9463 24271 9469
rect 24673 9469 24685 9472
rect 24719 9469 24731 9503
rect 24673 9463 24731 9469
rect 24765 9503 24823 9509
rect 24765 9469 24777 9503
rect 24811 9500 24823 9503
rect 25314 9500 25320 9512
rect 24811 9472 25320 9500
rect 24811 9469 24823 9472
rect 24765 9463 24823 9469
rect 24084 9336 24164 9364
rect 24228 9364 24256 9463
rect 24688 9432 24716 9463
rect 25314 9460 25320 9472
rect 25372 9460 25378 9512
rect 25869 9503 25927 9509
rect 25869 9469 25881 9503
rect 25915 9469 25927 9503
rect 27062 9500 27068 9512
rect 27023 9472 27068 9500
rect 25869 9463 25927 9469
rect 25038 9432 25044 9444
rect 24688 9404 25044 9432
rect 25038 9392 25044 9404
rect 25096 9392 25102 9444
rect 24762 9364 24768 9376
rect 24228 9336 24768 9364
rect 24084 9324 24090 9336
rect 24762 9324 24768 9336
rect 24820 9364 24826 9376
rect 25884 9364 25912 9463
rect 27062 9460 27068 9472
rect 27120 9460 27126 9512
rect 27525 9503 27583 9509
rect 27525 9469 27537 9503
rect 27571 9469 27583 9503
rect 27525 9463 27583 9469
rect 26326 9392 26332 9444
rect 26384 9432 26390 9444
rect 27540 9432 27568 9463
rect 27614 9460 27620 9512
rect 27672 9500 27678 9512
rect 27672 9472 27717 9500
rect 27672 9460 27678 9472
rect 28000 9432 28028 9540
rect 29380 9512 29408 9540
rect 29549 9537 29561 9571
rect 29595 9568 29607 9571
rect 30466 9568 30472 9580
rect 29595 9540 30472 9568
rect 29595 9537 29607 9540
rect 29549 9531 29607 9537
rect 30466 9528 30472 9540
rect 30524 9528 30530 9580
rect 31662 9528 31668 9580
rect 31720 9568 31726 9580
rect 34072 9568 34100 9596
rect 34514 9568 34520 9580
rect 31720 9540 32076 9568
rect 34072 9540 34520 9568
rect 31720 9528 31726 9540
rect 29086 9500 29092 9512
rect 29047 9472 29092 9500
rect 29086 9460 29092 9472
rect 29144 9460 29150 9512
rect 29178 9460 29184 9512
rect 29236 9500 29242 9512
rect 29273 9503 29331 9509
rect 29273 9500 29285 9503
rect 29236 9472 29285 9500
rect 29236 9460 29242 9472
rect 29273 9469 29285 9472
rect 29319 9469 29331 9503
rect 29273 9463 29331 9469
rect 29362 9460 29368 9512
rect 29420 9460 29426 9512
rect 31386 9500 31392 9512
rect 31347 9472 31392 9500
rect 31386 9460 31392 9472
rect 31444 9460 31450 9512
rect 32048 9509 32076 9540
rect 34514 9528 34520 9540
rect 34572 9528 34578 9580
rect 35802 9568 35808 9580
rect 35763 9540 35808 9568
rect 35802 9528 35808 9540
rect 35860 9528 35866 9580
rect 36924 9577 36952 9608
rect 36909 9571 36967 9577
rect 36909 9537 36921 9571
rect 36955 9568 36967 9571
rect 37366 9568 37372 9580
rect 36955 9540 37372 9568
rect 36955 9537 36967 9540
rect 36909 9531 36967 9537
rect 37366 9528 37372 9540
rect 37424 9528 37430 9580
rect 32033 9503 32091 9509
rect 32033 9469 32045 9503
rect 32079 9469 32091 9503
rect 32214 9500 32220 9512
rect 32175 9472 32220 9500
rect 32033 9463 32091 9469
rect 32214 9460 32220 9472
rect 32272 9460 32278 9512
rect 33413 9503 33471 9509
rect 33413 9469 33425 9503
rect 33459 9469 33471 9503
rect 33962 9500 33968 9512
rect 33923 9472 33968 9500
rect 33413 9463 33471 9469
rect 26384 9404 28028 9432
rect 28169 9435 28227 9441
rect 26384 9392 26390 9404
rect 28169 9401 28181 9435
rect 28215 9432 28227 9435
rect 28258 9432 28264 9444
rect 28215 9404 28264 9432
rect 28215 9401 28227 9404
rect 28169 9395 28227 9401
rect 28258 9392 28264 9404
rect 28316 9392 28322 9444
rect 33428 9432 33456 9463
rect 33962 9460 33968 9472
rect 34020 9460 34026 9512
rect 34054 9460 34060 9512
rect 34112 9500 34118 9512
rect 34112 9472 34157 9500
rect 34112 9460 34118 9472
rect 35066 9460 35072 9512
rect 35124 9500 35130 9512
rect 35345 9503 35403 9509
rect 35345 9500 35357 9503
rect 35124 9472 35357 9500
rect 35124 9460 35130 9472
rect 35345 9469 35357 9472
rect 35391 9469 35403 9503
rect 35710 9500 35716 9512
rect 35671 9472 35716 9500
rect 35345 9463 35403 9469
rect 35710 9460 35716 9472
rect 35768 9460 35774 9512
rect 37182 9500 37188 9512
rect 37143 9472 37188 9500
rect 37182 9460 37188 9472
rect 37240 9460 37246 9512
rect 34885 9435 34943 9441
rect 34885 9432 34897 9435
rect 28368 9404 29408 9432
rect 33428 9404 34897 9432
rect 24820 9336 25912 9364
rect 24820 9324 24826 9336
rect 26510 9324 26516 9376
rect 26568 9364 26574 9376
rect 28368 9364 28396 9404
rect 26568 9336 28396 9364
rect 28905 9367 28963 9373
rect 26568 9324 26574 9336
rect 28905 9333 28917 9367
rect 28951 9364 28963 9367
rect 29178 9364 29184 9376
rect 28951 9336 29184 9364
rect 28951 9333 28963 9336
rect 28905 9327 28963 9333
rect 29178 9324 29184 9336
rect 29236 9324 29242 9376
rect 29380 9364 29408 9404
rect 34885 9401 34897 9404
rect 34931 9401 34943 9435
rect 34885 9395 34943 9401
rect 30834 9364 30840 9376
rect 29380 9336 30840 9364
rect 30834 9324 30840 9336
rect 30892 9324 30898 9376
rect 31478 9364 31484 9376
rect 31439 9336 31484 9364
rect 31478 9324 31484 9336
rect 31536 9324 31542 9376
rect 33321 9367 33379 9373
rect 33321 9333 33333 9367
rect 33367 9364 33379 9367
rect 35250 9364 35256 9376
rect 33367 9336 35256 9364
rect 33367 9333 33379 9336
rect 33321 9327 33379 9333
rect 35250 9324 35256 9336
rect 35308 9324 35314 9376
rect 1104 9274 39836 9296
rect 1104 9222 19606 9274
rect 19658 9222 19670 9274
rect 19722 9222 19734 9274
rect 19786 9222 19798 9274
rect 19850 9222 39836 9274
rect 1104 9200 39836 9222
rect 2958 9160 2964 9172
rect 2919 9132 2964 9160
rect 2958 9120 2964 9132
rect 3016 9120 3022 9172
rect 13354 9120 13360 9172
rect 13412 9160 13418 9172
rect 13449 9163 13507 9169
rect 13449 9160 13461 9163
rect 13412 9132 13461 9160
rect 13412 9120 13418 9132
rect 13449 9129 13461 9132
rect 13495 9129 13507 9163
rect 13449 9123 13507 9129
rect 15470 9120 15476 9172
rect 15528 9160 15534 9172
rect 18322 9160 18328 9172
rect 15528 9132 18184 9160
rect 18283 9132 18328 9160
rect 15528 9120 15534 9132
rect 18156 9092 18184 9132
rect 18322 9120 18328 9132
rect 18380 9120 18386 9172
rect 21358 9120 21364 9172
rect 21416 9160 21422 9172
rect 23382 9160 23388 9172
rect 21416 9132 23388 9160
rect 21416 9120 21422 9132
rect 23382 9120 23388 9132
rect 23440 9120 23446 9172
rect 24762 9160 24768 9172
rect 24136 9132 24768 9160
rect 19058 9092 19064 9104
rect 5828 9064 17080 9092
rect 18156 9064 19064 9092
rect 1670 9024 1676 9036
rect 1631 8996 1676 9024
rect 1670 8984 1676 8996
rect 1728 8984 1734 9036
rect 3881 9027 3939 9033
rect 3881 8993 3893 9027
rect 3927 9024 3939 9027
rect 4062 9024 4068 9036
rect 3927 8996 4068 9024
rect 3927 8993 3939 8996
rect 3881 8987 3939 8993
rect 4062 8984 4068 8996
rect 4120 8984 4126 9036
rect 4430 9024 4436 9036
rect 4391 8996 4436 9024
rect 4430 8984 4436 8996
rect 4488 8984 4494 9036
rect 4890 9024 4896 9036
rect 4851 8996 4896 9024
rect 4890 8984 4896 8996
rect 4948 8984 4954 9036
rect 5166 8984 5172 9036
rect 5224 9024 5230 9036
rect 5442 9024 5448 9036
rect 5224 8996 5448 9024
rect 5224 8984 5230 8996
rect 5442 8984 5448 8996
rect 5500 8984 5506 9036
rect 5828 9033 5856 9064
rect 5813 9027 5871 9033
rect 5813 8993 5825 9027
rect 5859 8993 5871 9027
rect 6086 9024 6092 9036
rect 6047 8996 6092 9024
rect 5813 8987 5871 8993
rect 6086 8984 6092 8996
rect 6144 8984 6150 9036
rect 7098 8984 7104 9036
rect 7156 9024 7162 9036
rect 7193 9027 7251 9033
rect 7193 9024 7205 9027
rect 7156 8996 7205 9024
rect 7156 8984 7162 8996
rect 7193 8993 7205 8996
rect 7239 8993 7251 9027
rect 7742 9024 7748 9036
rect 7703 8996 7748 9024
rect 7193 8987 7251 8993
rect 7742 8984 7748 8996
rect 7800 8984 7806 9036
rect 8110 9024 8116 9036
rect 8071 8996 8116 9024
rect 8110 8984 8116 8996
rect 8168 8984 8174 9036
rect 8588 9033 8616 9064
rect 8573 9027 8631 9033
rect 8573 8993 8585 9027
rect 8619 8993 8631 9027
rect 9030 9024 9036 9036
rect 8991 8996 9036 9024
rect 8573 8987 8631 8993
rect 9030 8984 9036 8996
rect 9088 8984 9094 9036
rect 10134 8984 10140 9036
rect 10192 9024 10198 9036
rect 10689 9027 10747 9033
rect 10689 9024 10701 9027
rect 10192 8996 10701 9024
rect 10192 8984 10198 8996
rect 10689 8993 10701 8996
rect 10735 8993 10747 9027
rect 10689 8987 10747 8993
rect 11057 9027 11115 9033
rect 11057 8993 11069 9027
rect 11103 9024 11115 9027
rect 11701 9027 11759 9033
rect 11701 9024 11713 9027
rect 11103 8996 11713 9024
rect 11103 8993 11115 8996
rect 11057 8987 11115 8993
rect 11701 8993 11713 8996
rect 11747 8993 11759 9027
rect 12342 9024 12348 9036
rect 12303 8996 12348 9024
rect 11701 8987 11759 8993
rect 12342 8984 12348 8996
rect 12400 8984 12406 9036
rect 12710 9024 12716 9036
rect 12671 8996 12716 9024
rect 12710 8984 12716 8996
rect 12768 8984 12774 9036
rect 13262 8984 13268 9036
rect 13320 9024 13326 9036
rect 13357 9027 13415 9033
rect 13357 9024 13369 9027
rect 13320 8996 13369 9024
rect 13320 8984 13326 8996
rect 13357 8993 13369 8996
rect 13403 8993 13415 9027
rect 13357 8987 13415 8993
rect 13722 8984 13728 9036
rect 13780 9024 13786 9036
rect 13909 9027 13967 9033
rect 13909 9024 13921 9027
rect 13780 8996 13921 9024
rect 13780 8984 13786 8996
rect 13909 8993 13921 8996
rect 13955 8993 13967 9027
rect 13909 8987 13967 8993
rect 15746 8984 15752 9036
rect 15804 9024 15810 9036
rect 15933 9027 15991 9033
rect 15933 9024 15945 9027
rect 15804 8996 15945 9024
rect 15804 8984 15810 8996
rect 15933 8993 15945 8996
rect 15979 8993 15991 9027
rect 16298 9024 16304 9036
rect 16259 8996 16304 9024
rect 15933 8987 15991 8993
rect 16298 8984 16304 8996
rect 16356 8984 16362 9036
rect 1394 8956 1400 8968
rect 1355 8928 1400 8956
rect 1394 8916 1400 8928
rect 1452 8916 1458 8968
rect 4798 8956 4804 8968
rect 4759 8928 4804 8956
rect 4798 8916 4804 8928
rect 4856 8916 4862 8968
rect 7282 8956 7288 8968
rect 7243 8928 7288 8956
rect 7282 8916 7288 8928
rect 7340 8916 7346 8968
rect 11146 8956 11152 8968
rect 11107 8928 11152 8956
rect 11146 8916 11152 8928
rect 11204 8916 11210 8968
rect 12250 8956 12256 8968
rect 12211 8928 12256 8956
rect 12250 8916 12256 8928
rect 12308 8916 12314 8968
rect 12805 8959 12863 8965
rect 12360 8928 12756 8956
rect 10505 8891 10563 8897
rect 10505 8857 10517 8891
rect 10551 8888 10563 8891
rect 12360 8888 12388 8928
rect 10551 8860 12388 8888
rect 10551 8857 10563 8860
rect 10505 8851 10563 8857
rect 3694 8820 3700 8832
rect 3655 8792 3700 8820
rect 3694 8780 3700 8792
rect 3752 8780 3758 8832
rect 12728 8820 12756 8928
rect 12805 8925 12817 8959
rect 12851 8925 12863 8959
rect 14182 8956 14188 8968
rect 12805 8919 12863 8925
rect 13004 8928 14188 8956
rect 12820 8888 12848 8919
rect 13004 8888 13032 8928
rect 14182 8916 14188 8928
rect 14240 8916 14246 8968
rect 14366 8956 14372 8968
rect 14327 8928 14372 8956
rect 14366 8916 14372 8928
rect 14424 8916 14430 8968
rect 15838 8956 15844 8968
rect 15799 8928 15844 8956
rect 15838 8916 15844 8928
rect 15896 8916 15902 8968
rect 16206 8916 16212 8968
rect 16264 8956 16270 8968
rect 16393 8959 16451 8965
rect 16393 8956 16405 8959
rect 16264 8928 16405 8956
rect 16264 8916 16270 8928
rect 16393 8925 16405 8928
rect 16439 8925 16451 8959
rect 16942 8956 16948 8968
rect 16903 8928 16948 8956
rect 16393 8919 16451 8925
rect 16942 8916 16948 8928
rect 17000 8916 17006 8968
rect 17052 8956 17080 9064
rect 19058 9052 19064 9064
rect 19116 9052 19122 9104
rect 19153 9095 19211 9101
rect 19153 9061 19165 9095
rect 19199 9092 19211 9095
rect 19334 9092 19340 9104
rect 19199 9064 19340 9092
rect 19199 9061 19211 9064
rect 19153 9055 19211 9061
rect 19334 9052 19340 9064
rect 19392 9052 19398 9104
rect 23750 9092 23756 9104
rect 23216 9064 23756 9092
rect 17221 9027 17279 9033
rect 17221 8993 17233 9027
rect 17267 9024 17279 9027
rect 17310 9024 17316 9036
rect 17267 8996 17316 9024
rect 17267 8993 17279 8996
rect 17221 8987 17279 8993
rect 17310 8984 17316 8996
rect 17368 8984 17374 9036
rect 19794 9024 19800 9036
rect 19755 8996 19800 9024
rect 19794 8984 19800 8996
rect 19852 8984 19858 9036
rect 19886 8984 19892 9036
rect 19944 9024 19950 9036
rect 20162 9024 20168 9036
rect 19944 8996 19989 9024
rect 20123 8996 20168 9024
rect 19944 8984 19950 8996
rect 20162 8984 20168 8996
rect 20220 8984 20226 9036
rect 21821 9027 21879 9033
rect 21821 8993 21833 9027
rect 21867 8993 21879 9027
rect 22186 9024 22192 9036
rect 22147 8996 22192 9024
rect 21821 8987 21879 8993
rect 17052 8928 18460 8956
rect 12820 8860 13032 8888
rect 13078 8848 13084 8900
rect 13136 8888 13142 8900
rect 15654 8888 15660 8900
rect 13136 8860 15660 8888
rect 13136 8848 13142 8860
rect 15654 8848 15660 8860
rect 15712 8848 15718 8900
rect 13906 8820 13912 8832
rect 12728 8792 13912 8820
rect 13906 8780 13912 8792
rect 13964 8780 13970 8832
rect 15381 8823 15439 8829
rect 15381 8789 15393 8823
rect 15427 8820 15439 8823
rect 18046 8820 18052 8832
rect 15427 8792 18052 8820
rect 15427 8789 15439 8792
rect 15381 8783 15439 8789
rect 18046 8780 18052 8792
rect 18104 8780 18110 8832
rect 18432 8820 18460 8928
rect 19426 8916 19432 8968
rect 19484 8956 19490 8968
rect 20257 8959 20315 8965
rect 20257 8956 20269 8959
rect 19484 8928 20269 8956
rect 19484 8916 19490 8928
rect 20257 8925 20269 8928
rect 20303 8925 20315 8959
rect 21358 8956 21364 8968
rect 21319 8928 21364 8956
rect 20257 8919 20315 8925
rect 21358 8916 21364 8928
rect 21416 8916 21422 8968
rect 21450 8916 21456 8968
rect 21508 8956 21514 8968
rect 21836 8956 21864 8987
rect 22186 8984 22192 8996
rect 22244 8984 22250 9036
rect 23216 9033 23244 9064
rect 23750 9052 23756 9064
rect 23808 9052 23814 9104
rect 24136 9101 24164 9132
rect 24762 9120 24768 9132
rect 24820 9120 24826 9172
rect 26234 9160 26240 9172
rect 25056 9132 26240 9160
rect 24121 9095 24179 9101
rect 24121 9061 24133 9095
rect 24167 9061 24179 9095
rect 24121 9055 24179 9061
rect 23201 9027 23259 9033
rect 23201 8993 23213 9027
rect 23247 8993 23259 9027
rect 23201 8987 23259 8993
rect 23474 8984 23480 9036
rect 23532 9024 23538 9036
rect 23569 9027 23627 9033
rect 23569 9024 23581 9027
rect 23532 8996 23581 9024
rect 23532 8984 23538 8996
rect 23569 8993 23581 8996
rect 23615 8993 23627 9027
rect 23842 9024 23848 9036
rect 23803 8996 23848 9024
rect 23569 8987 23627 8993
rect 23382 8956 23388 8968
rect 21508 8928 23388 8956
rect 21508 8916 21514 8928
rect 23382 8916 23388 8928
rect 23440 8916 23446 8968
rect 23584 8956 23612 8987
rect 23842 8984 23848 8996
rect 23900 8984 23906 9036
rect 24026 8956 24032 8968
rect 23584 8928 24032 8956
rect 24026 8916 24032 8928
rect 24084 8916 24090 8968
rect 22094 8848 22100 8900
rect 22152 8888 22158 8900
rect 22152 8860 22197 8888
rect 22152 8848 22158 8860
rect 24136 8820 24164 9055
rect 24765 9027 24823 9033
rect 24765 8993 24777 9027
rect 24811 9024 24823 9027
rect 25056 9024 25084 9132
rect 26234 9120 26240 9132
rect 26292 9120 26298 9172
rect 26878 9120 26884 9172
rect 26936 9160 26942 9172
rect 27433 9163 27491 9169
rect 27433 9160 27445 9163
rect 26936 9132 27445 9160
rect 26936 9120 26942 9132
rect 27433 9129 27445 9132
rect 27479 9129 27491 9163
rect 30190 9160 30196 9172
rect 30151 9132 30196 9160
rect 27433 9123 27491 9129
rect 30190 9120 30196 9132
rect 30248 9120 30254 9172
rect 31478 9120 31484 9172
rect 31536 9160 31542 9172
rect 36354 9160 36360 9172
rect 31536 9132 35940 9160
rect 36315 9132 36360 9160
rect 31536 9120 31542 9132
rect 26605 9095 26663 9101
rect 26605 9092 26617 9095
rect 25240 9064 26617 9092
rect 25240 9036 25268 9064
rect 26605 9061 26617 9064
rect 26651 9061 26663 9095
rect 26605 9055 26663 9061
rect 31202 9052 31208 9104
rect 31260 9092 31266 9104
rect 31938 9092 31944 9104
rect 31260 9064 31944 9092
rect 31260 9052 31266 9064
rect 31938 9052 31944 9064
rect 31996 9052 32002 9104
rect 34238 9052 34244 9104
rect 34296 9092 34302 9104
rect 35066 9092 35072 9104
rect 34296 9064 35072 9092
rect 34296 9052 34302 9064
rect 35066 9052 35072 9064
rect 35124 9052 35130 9104
rect 35912 9092 35940 9132
rect 36354 9120 36360 9132
rect 36412 9120 36418 9172
rect 37182 9120 37188 9172
rect 37240 9160 37246 9172
rect 37829 9163 37887 9169
rect 37829 9160 37841 9163
rect 37240 9132 37841 9160
rect 37240 9120 37246 9132
rect 37829 9129 37841 9132
rect 37875 9129 37887 9163
rect 37829 9123 37887 9129
rect 35912 9064 38608 9092
rect 25222 9024 25228 9036
rect 24811 8996 25084 9024
rect 25183 8996 25228 9024
rect 24811 8993 24823 8996
rect 24765 8987 24823 8993
rect 25222 8984 25228 8996
rect 25280 8984 25286 9036
rect 25317 9027 25375 9033
rect 25317 8993 25329 9027
rect 25363 9024 25375 9027
rect 25363 8996 26188 9024
rect 25363 8993 25375 8996
rect 25317 8987 25375 8993
rect 24673 8959 24731 8965
rect 24673 8925 24685 8959
rect 24719 8956 24731 8959
rect 24854 8956 24860 8968
rect 24719 8928 24860 8956
rect 24719 8925 24731 8928
rect 24673 8919 24731 8925
rect 24854 8916 24860 8928
rect 24912 8916 24918 8968
rect 26160 8956 26188 8996
rect 26234 8984 26240 9036
rect 26292 9024 26298 9036
rect 26513 9027 26571 9033
rect 26513 9024 26525 9027
rect 26292 8996 26525 9024
rect 26292 8984 26298 8996
rect 26513 8993 26525 8996
rect 26559 8993 26571 9027
rect 26513 8987 26571 8993
rect 27341 9027 27399 9033
rect 27341 8993 27353 9027
rect 27387 9024 27399 9027
rect 28261 9027 28319 9033
rect 27387 8996 28212 9024
rect 27387 8993 27399 8996
rect 27341 8987 27399 8993
rect 27430 8956 27436 8968
rect 26160 8928 27436 8956
rect 27430 8916 27436 8928
rect 27488 8916 27494 8968
rect 27982 8956 27988 8968
rect 27943 8928 27988 8956
rect 27982 8916 27988 8928
rect 28040 8916 28046 8968
rect 28184 8956 28212 8996
rect 28261 8993 28273 9027
rect 28307 9024 28319 9027
rect 28350 9024 28356 9036
rect 28307 8996 28356 9024
rect 28307 8993 28319 8996
rect 28261 8987 28319 8993
rect 28350 8984 28356 8996
rect 28408 8984 28414 9036
rect 30098 9024 30104 9036
rect 30059 8996 30104 9024
rect 30098 8984 30104 8996
rect 30156 8984 30162 9036
rect 30745 9027 30803 9033
rect 30745 8993 30757 9027
rect 30791 9024 30803 9027
rect 31018 9024 31024 9036
rect 30791 8996 31024 9024
rect 30791 8993 30803 8996
rect 30745 8987 30803 8993
rect 31018 8984 31024 8996
rect 31076 8984 31082 9036
rect 32125 9027 32183 9033
rect 32125 9024 32137 9027
rect 31312 8996 32137 9024
rect 31312 8968 31340 8996
rect 32125 8993 32137 8996
rect 32171 8993 32183 9027
rect 33134 9024 33140 9036
rect 33095 8996 33140 9024
rect 32125 8987 32183 8993
rect 33134 8984 33140 8996
rect 33192 8984 33198 9036
rect 35250 9024 35256 9036
rect 35211 8996 35256 9024
rect 35250 8984 35256 8996
rect 35308 8984 35314 9036
rect 37550 8984 37556 9036
rect 37608 9024 37614 9036
rect 37737 9027 37795 9033
rect 37737 9024 37749 9027
rect 37608 8996 37749 9024
rect 37608 8984 37614 8996
rect 37737 8993 37749 8996
rect 37783 8993 37795 9027
rect 38470 9024 38476 9036
rect 38431 8996 38476 9024
rect 37737 8987 37795 8993
rect 38470 8984 38476 8996
rect 38528 8984 38534 9036
rect 38580 9033 38608 9064
rect 38565 9027 38623 9033
rect 38565 8993 38577 9027
rect 38611 8993 38623 9027
rect 38565 8987 38623 8993
rect 31294 8956 31300 8968
rect 28184 8928 31300 8956
rect 31294 8916 31300 8928
rect 31352 8916 31358 8968
rect 32861 8959 32919 8965
rect 32861 8925 32873 8959
rect 32907 8956 32919 8959
rect 33502 8956 33508 8968
rect 32907 8928 33508 8956
rect 32907 8925 32919 8928
rect 32861 8919 32919 8925
rect 33502 8916 33508 8928
rect 33560 8956 33566 8968
rect 34330 8956 34336 8968
rect 33560 8928 34336 8956
rect 33560 8916 33566 8928
rect 34330 8916 34336 8928
rect 34388 8956 34394 8968
rect 34977 8959 35035 8965
rect 34977 8956 34989 8959
rect 34388 8928 34989 8956
rect 34388 8916 34394 8928
rect 34977 8925 34989 8928
rect 35023 8925 35035 8959
rect 34977 8919 35035 8925
rect 24946 8848 24952 8900
rect 25004 8888 25010 8900
rect 25685 8891 25743 8897
rect 25685 8888 25697 8891
rect 25004 8860 25697 8888
rect 25004 8848 25010 8860
rect 25685 8857 25697 8860
rect 25731 8857 25743 8891
rect 25685 8851 25743 8857
rect 28994 8848 29000 8900
rect 29052 8888 29058 8900
rect 29822 8888 29828 8900
rect 29052 8860 29828 8888
rect 29052 8848 29058 8860
rect 29822 8848 29828 8860
rect 29880 8888 29886 8900
rect 30929 8891 30987 8897
rect 30929 8888 30941 8891
rect 29880 8860 30941 8888
rect 29880 8848 29886 8860
rect 30929 8857 30941 8860
rect 30975 8888 30987 8891
rect 31662 8888 31668 8900
rect 30975 8860 31668 8888
rect 30975 8857 30987 8860
rect 30929 8851 30987 8857
rect 31662 8848 31668 8860
rect 31720 8848 31726 8900
rect 18432 8792 24164 8820
rect 24854 8780 24860 8832
rect 24912 8820 24918 8832
rect 25866 8820 25872 8832
rect 24912 8792 25872 8820
rect 24912 8780 24918 8792
rect 25866 8780 25872 8792
rect 25924 8780 25930 8832
rect 29270 8780 29276 8832
rect 29328 8820 29334 8832
rect 29365 8823 29423 8829
rect 29365 8820 29377 8823
rect 29328 8792 29377 8820
rect 29328 8780 29334 8792
rect 29365 8789 29377 8792
rect 29411 8789 29423 8823
rect 29365 8783 29423 8789
rect 31846 8780 31852 8832
rect 31904 8820 31910 8832
rect 32309 8823 32367 8829
rect 32309 8820 32321 8823
rect 31904 8792 32321 8820
rect 31904 8780 31910 8792
rect 32309 8789 32321 8792
rect 32355 8789 32367 8823
rect 34422 8820 34428 8832
rect 34383 8792 34428 8820
rect 32309 8783 32367 8789
rect 34422 8780 34428 8792
rect 34480 8780 34486 8832
rect 1104 8730 39836 8752
rect 1104 8678 4246 8730
rect 4298 8678 4310 8730
rect 4362 8678 4374 8730
rect 4426 8678 4438 8730
rect 4490 8678 34966 8730
rect 35018 8678 35030 8730
rect 35082 8678 35094 8730
rect 35146 8678 35158 8730
rect 35210 8678 39836 8730
rect 1104 8656 39836 8678
rect 4062 8616 4068 8628
rect 4023 8588 4068 8616
rect 4062 8576 4068 8588
rect 4120 8576 4126 8628
rect 6178 8616 6184 8628
rect 6139 8588 6184 8616
rect 6178 8576 6184 8588
rect 6236 8576 6242 8628
rect 11793 8619 11851 8625
rect 11793 8585 11805 8619
rect 11839 8616 11851 8619
rect 12250 8616 12256 8628
rect 11839 8588 12256 8616
rect 11839 8585 11851 8588
rect 11793 8579 11851 8585
rect 12250 8576 12256 8588
rect 12308 8576 12314 8628
rect 21450 8616 21456 8628
rect 13924 8588 21456 8616
rect 6454 8508 6460 8560
rect 6512 8548 6518 8560
rect 11241 8551 11299 8557
rect 11241 8548 11253 8551
rect 6512 8520 11253 8548
rect 6512 8508 6518 8520
rect 11241 8517 11253 8520
rect 11287 8548 11299 8551
rect 12342 8548 12348 8560
rect 11287 8520 12348 8548
rect 11287 8517 11299 8520
rect 11241 8511 11299 8517
rect 12342 8508 12348 8520
rect 12400 8548 12406 8560
rect 12894 8548 12900 8560
rect 12400 8520 12900 8548
rect 12400 8508 12406 8520
rect 12894 8508 12900 8520
rect 12952 8508 12958 8560
rect 13078 8548 13084 8560
rect 13039 8520 13084 8548
rect 13078 8508 13084 8520
rect 13136 8508 13142 8560
rect 2774 8440 2780 8492
rect 2832 8480 2838 8492
rect 2832 8452 2877 8480
rect 2832 8440 2838 8452
rect 4798 8440 4804 8492
rect 4856 8480 4862 8492
rect 4893 8483 4951 8489
rect 4893 8480 4905 8483
rect 4856 8452 4905 8480
rect 4856 8440 4862 8452
rect 4893 8449 4905 8452
rect 4939 8449 4951 8483
rect 7190 8480 7196 8492
rect 7151 8452 7196 8480
rect 4893 8443 4951 8449
rect 7190 8440 7196 8452
rect 7248 8440 7254 8492
rect 8662 8480 8668 8492
rect 7760 8452 8668 8480
rect 1394 8412 1400 8424
rect 1355 8384 1400 8412
rect 1394 8372 1400 8384
rect 1452 8372 1458 8424
rect 1670 8412 1676 8424
rect 1631 8384 1676 8412
rect 1670 8372 1676 8384
rect 1728 8372 1734 8424
rect 3973 8415 4031 8421
rect 3973 8381 3985 8415
rect 4019 8412 4031 8415
rect 4617 8415 4675 8421
rect 4019 8384 4568 8412
rect 4019 8381 4031 8384
rect 3973 8375 4031 8381
rect 4540 8276 4568 8384
rect 4617 8381 4629 8415
rect 4663 8412 4675 8415
rect 4982 8412 4988 8424
rect 4663 8384 4988 8412
rect 4663 8381 4675 8384
rect 4617 8375 4675 8381
rect 4982 8372 4988 8384
rect 5040 8412 5046 8424
rect 5166 8412 5172 8424
rect 5040 8384 5172 8412
rect 5040 8372 5046 8384
rect 5166 8372 5172 8384
rect 5224 8412 5230 8424
rect 6454 8412 6460 8424
rect 5224 8384 6460 8412
rect 5224 8372 5230 8384
rect 6454 8372 6460 8384
rect 6512 8372 6518 8424
rect 7098 8412 7104 8424
rect 7059 8384 7104 8412
rect 7098 8372 7104 8384
rect 7156 8372 7162 8424
rect 7760 8421 7788 8452
rect 8662 8440 8668 8452
rect 8720 8440 8726 8492
rect 13262 8440 13268 8492
rect 13320 8480 13326 8492
rect 13541 8483 13599 8489
rect 13541 8480 13553 8483
rect 13320 8452 13553 8480
rect 13320 8440 13326 8452
rect 13541 8449 13553 8452
rect 13587 8449 13599 8483
rect 13541 8443 13599 8449
rect 7745 8415 7803 8421
rect 7745 8381 7757 8415
rect 7791 8381 7803 8415
rect 8110 8412 8116 8424
rect 8071 8384 8116 8412
rect 7745 8375 7803 8381
rect 8110 8372 8116 8384
rect 8168 8372 8174 8424
rect 8297 8415 8355 8421
rect 8297 8381 8309 8415
rect 8343 8381 8355 8415
rect 9030 8412 9036 8424
rect 8991 8384 9036 8412
rect 8297 8375 8355 8381
rect 5902 8304 5908 8356
rect 5960 8344 5966 8356
rect 8312 8344 8340 8375
rect 9030 8372 9036 8384
rect 9088 8412 9094 8424
rect 9674 8412 9680 8424
rect 9088 8384 9680 8412
rect 9088 8372 9094 8384
rect 9674 8372 9680 8384
rect 9732 8372 9738 8424
rect 9858 8372 9864 8424
rect 9916 8412 9922 8424
rect 10045 8415 10103 8421
rect 10045 8412 10057 8415
rect 9916 8384 10057 8412
rect 9916 8372 9922 8384
rect 10045 8381 10057 8384
rect 10091 8381 10103 8415
rect 10594 8412 10600 8424
rect 10555 8384 10600 8412
rect 10045 8375 10103 8381
rect 10594 8372 10600 8384
rect 10652 8372 10658 8424
rect 11238 8372 11244 8424
rect 11296 8412 11302 8424
rect 11425 8415 11483 8421
rect 11425 8412 11437 8415
rect 11296 8384 11437 8412
rect 11296 8372 11302 8384
rect 11425 8381 11437 8384
rect 11471 8381 11483 8415
rect 11425 8375 11483 8381
rect 11701 8415 11759 8421
rect 11701 8381 11713 8415
rect 11747 8412 11759 8415
rect 12066 8412 12072 8424
rect 11747 8384 12072 8412
rect 11747 8381 11759 8384
rect 11701 8375 11759 8381
rect 12066 8372 12072 8384
rect 12124 8372 12130 8424
rect 12526 8372 12532 8424
rect 12584 8412 12590 8424
rect 13633 8415 13691 8421
rect 13633 8412 13645 8415
rect 12584 8384 13645 8412
rect 12584 8372 12590 8384
rect 13633 8381 13645 8384
rect 13679 8381 13691 8415
rect 13633 8375 13691 8381
rect 13924 8344 13952 8588
rect 21450 8576 21456 8588
rect 21508 8576 21514 8628
rect 23842 8576 23848 8628
rect 23900 8616 23906 8628
rect 24121 8619 24179 8625
rect 24121 8616 24133 8619
rect 23900 8588 24133 8616
rect 23900 8576 23906 8588
rect 24121 8585 24133 8588
rect 24167 8616 24179 8619
rect 24394 8616 24400 8628
rect 24167 8588 24400 8616
rect 24167 8585 24179 8588
rect 24121 8579 24179 8585
rect 24394 8576 24400 8588
rect 24452 8576 24458 8628
rect 26234 8616 26240 8628
rect 26195 8588 26240 8616
rect 26234 8576 26240 8588
rect 26292 8576 26298 8628
rect 30837 8619 30895 8625
rect 30837 8585 30849 8619
rect 30883 8616 30895 8619
rect 31018 8616 31024 8628
rect 30883 8588 31024 8616
rect 30883 8585 30895 8588
rect 30837 8579 30895 8585
rect 31018 8576 31024 8588
rect 31076 8576 31082 8628
rect 34054 8616 34060 8628
rect 31680 8588 34060 8616
rect 14182 8548 14188 8560
rect 14095 8520 14188 8548
rect 14108 8489 14136 8520
rect 14182 8508 14188 8520
rect 14240 8548 14246 8560
rect 16206 8548 16212 8560
rect 14240 8520 16212 8548
rect 14240 8508 14246 8520
rect 16206 8508 16212 8520
rect 16264 8508 16270 8560
rect 23290 8548 23296 8560
rect 17328 8520 23296 8548
rect 14093 8483 14151 8489
rect 14093 8449 14105 8483
rect 14139 8449 14151 8483
rect 16022 8480 16028 8492
rect 15983 8452 16028 8480
rect 14093 8443 14151 8449
rect 16022 8440 16028 8452
rect 16080 8440 16086 8492
rect 16390 8440 16396 8492
rect 16448 8480 16454 8492
rect 16577 8483 16635 8489
rect 16577 8480 16589 8483
rect 16448 8452 16589 8480
rect 16448 8440 16454 8452
rect 16577 8449 16589 8452
rect 16623 8449 16635 8483
rect 16577 8443 16635 8449
rect 14001 8415 14059 8421
rect 14001 8381 14013 8415
rect 14047 8381 14059 8415
rect 16114 8412 16120 8424
rect 16075 8384 16120 8412
rect 14001 8375 14059 8381
rect 5960 8316 13952 8344
rect 14016 8344 14044 8375
rect 16114 8372 16120 8384
rect 16172 8372 16178 8424
rect 16485 8415 16543 8421
rect 16485 8381 16497 8415
rect 16531 8412 16543 8415
rect 17126 8412 17132 8424
rect 16531 8384 17132 8412
rect 16531 8381 16543 8384
rect 16485 8375 16543 8381
rect 17126 8372 17132 8384
rect 17184 8372 17190 8424
rect 17328 8421 17356 8520
rect 23290 8508 23296 8520
rect 23348 8508 23354 8560
rect 31680 8557 31708 8588
rect 34054 8576 34060 8588
rect 34112 8576 34118 8628
rect 38286 8576 38292 8628
rect 38344 8616 38350 8628
rect 38473 8619 38531 8625
rect 38473 8616 38485 8619
rect 38344 8588 38485 8616
rect 38344 8576 38350 8588
rect 38473 8585 38485 8588
rect 38519 8585 38531 8619
rect 38473 8579 38531 8585
rect 31665 8551 31723 8557
rect 31665 8517 31677 8551
rect 31711 8517 31723 8551
rect 33226 8548 33232 8560
rect 33187 8520 33232 8548
rect 31665 8511 31723 8517
rect 33226 8508 33232 8520
rect 33284 8508 33290 8560
rect 18417 8483 18475 8489
rect 18417 8449 18429 8483
rect 18463 8480 18475 8483
rect 18782 8480 18788 8492
rect 18463 8452 18788 8480
rect 18463 8449 18475 8452
rect 18417 8443 18475 8449
rect 18782 8440 18788 8452
rect 18840 8440 18846 8492
rect 19794 8440 19800 8492
rect 19852 8480 19858 8492
rect 20073 8483 20131 8489
rect 20073 8480 20085 8483
rect 19852 8452 20085 8480
rect 19852 8440 19858 8452
rect 20073 8449 20085 8452
rect 20119 8449 20131 8483
rect 20073 8443 20131 8449
rect 21453 8483 21511 8489
rect 21453 8449 21465 8483
rect 21499 8480 21511 8483
rect 21542 8480 21548 8492
rect 21499 8452 21548 8480
rect 21499 8449 21511 8452
rect 21453 8443 21511 8449
rect 21542 8440 21548 8452
rect 21600 8440 21606 8492
rect 22186 8480 22192 8492
rect 22147 8452 22192 8480
rect 22186 8440 22192 8452
rect 22244 8440 22250 8492
rect 23860 8452 24532 8480
rect 17313 8415 17371 8421
rect 17313 8381 17325 8415
rect 17359 8381 17371 8415
rect 17313 8375 17371 8381
rect 17402 8372 17408 8424
rect 17460 8412 17466 8424
rect 18046 8412 18052 8424
rect 17460 8384 17505 8412
rect 18007 8384 18052 8412
rect 17460 8372 17466 8384
rect 18046 8372 18052 8384
rect 18104 8372 18110 8424
rect 18601 8415 18659 8421
rect 18601 8381 18613 8415
rect 18647 8381 18659 8415
rect 18601 8375 18659 8381
rect 15378 8344 15384 8356
rect 14016 8316 15384 8344
rect 5960 8304 5966 8316
rect 15378 8304 15384 8316
rect 15436 8304 15442 8356
rect 15473 8347 15531 8353
rect 15473 8313 15485 8347
rect 15519 8344 15531 8347
rect 18616 8344 18644 8375
rect 19058 8372 19064 8424
rect 19116 8412 19122 8424
rect 19521 8415 19579 8421
rect 19521 8412 19533 8415
rect 19116 8384 19533 8412
rect 19116 8372 19122 8384
rect 19521 8381 19533 8384
rect 19567 8381 19579 8415
rect 19521 8375 19579 8381
rect 19981 8415 20039 8421
rect 19981 8381 19993 8415
rect 20027 8381 20039 8415
rect 20990 8412 20996 8424
rect 20951 8384 20996 8412
rect 19981 8375 20039 8381
rect 15519 8316 18644 8344
rect 19996 8344 20024 8375
rect 20990 8372 20996 8384
rect 21048 8372 21054 8424
rect 21269 8415 21327 8421
rect 21269 8381 21281 8415
rect 21315 8412 21327 8415
rect 21910 8412 21916 8424
rect 21315 8384 21772 8412
rect 21871 8384 21916 8412
rect 21315 8381 21327 8384
rect 21269 8375 21327 8381
rect 21450 8344 21456 8356
rect 19996 8316 21456 8344
rect 15519 8313 15531 8316
rect 15473 8307 15531 8313
rect 21450 8304 21456 8316
rect 21508 8304 21514 8356
rect 21744 8344 21772 8384
rect 21910 8372 21916 8384
rect 21968 8372 21974 8424
rect 22462 8412 22468 8424
rect 22423 8384 22468 8412
rect 22462 8372 22468 8384
rect 22520 8372 22526 8424
rect 22646 8412 22652 8424
rect 22607 8384 22652 8412
rect 22646 8372 22652 8384
rect 22704 8372 22710 8424
rect 23860 8344 23888 8452
rect 23937 8415 23995 8421
rect 23937 8381 23949 8415
rect 23983 8381 23995 8415
rect 24504 8412 24532 8452
rect 24578 8440 24584 8492
rect 24636 8480 24642 8492
rect 24673 8483 24731 8489
rect 24673 8480 24685 8483
rect 24636 8452 24685 8480
rect 24636 8440 24642 8452
rect 24673 8449 24685 8452
rect 24719 8449 24731 8483
rect 24946 8480 24952 8492
rect 24907 8452 24952 8480
rect 24673 8443 24731 8449
rect 24946 8440 24952 8452
rect 25004 8440 25010 8492
rect 26789 8483 26847 8489
rect 26789 8449 26801 8483
rect 26835 8480 26847 8483
rect 27982 8480 27988 8492
rect 26835 8452 27988 8480
rect 26835 8449 26847 8452
rect 26789 8443 26847 8449
rect 27982 8440 27988 8452
rect 28040 8440 28046 8492
rect 28350 8440 28356 8492
rect 28408 8480 28414 8492
rect 28445 8483 28503 8489
rect 28445 8480 28457 8483
rect 28408 8452 28457 8480
rect 28408 8440 28414 8452
rect 28445 8449 28457 8452
rect 28491 8480 28503 8483
rect 28491 8452 36124 8480
rect 28491 8449 28503 8452
rect 28445 8443 28503 8449
rect 26326 8412 26332 8424
rect 24504 8384 26332 8412
rect 23937 8375 23995 8381
rect 21744 8316 23888 8344
rect 23952 8344 23980 8375
rect 26326 8372 26332 8384
rect 26384 8372 26390 8424
rect 27065 8415 27123 8421
rect 27065 8381 27077 8415
rect 27111 8412 27123 8415
rect 27706 8412 27712 8424
rect 27111 8384 27712 8412
rect 27111 8381 27123 8384
rect 27065 8375 27123 8381
rect 27706 8372 27712 8384
rect 27764 8372 27770 8424
rect 28000 8412 28028 8440
rect 29086 8412 29092 8424
rect 28000 8384 29092 8412
rect 29086 8372 29092 8384
rect 29144 8412 29150 8424
rect 29273 8415 29331 8421
rect 29273 8412 29285 8415
rect 29144 8384 29285 8412
rect 29144 8372 29150 8384
rect 29273 8381 29285 8384
rect 29319 8381 29331 8415
rect 29546 8412 29552 8424
rect 29507 8384 29552 8412
rect 29273 8375 29331 8381
rect 29546 8372 29552 8384
rect 29604 8372 29610 8424
rect 31386 8412 31392 8424
rect 31347 8384 31392 8412
rect 31386 8372 31392 8384
rect 31444 8372 31450 8424
rect 31938 8372 31944 8424
rect 31996 8412 32002 8424
rect 32033 8415 32091 8421
rect 32033 8412 32045 8415
rect 31996 8384 32045 8412
rect 31996 8372 32002 8384
rect 32033 8381 32045 8384
rect 32079 8381 32091 8415
rect 32214 8412 32220 8424
rect 32175 8384 32220 8412
rect 32033 8375 32091 8381
rect 32214 8372 32220 8384
rect 32272 8372 32278 8424
rect 33413 8415 33471 8421
rect 33413 8381 33425 8415
rect 33459 8381 33471 8415
rect 33778 8412 33784 8424
rect 33739 8384 33784 8412
rect 33413 8375 33471 8381
rect 33428 8344 33456 8375
rect 33778 8372 33784 8384
rect 33836 8372 33842 8424
rect 33870 8372 33876 8424
rect 33928 8412 33934 8424
rect 33928 8384 33973 8412
rect 33928 8372 33934 8384
rect 34330 8372 34336 8424
rect 34388 8412 34394 8424
rect 34514 8412 34520 8424
rect 34388 8384 34520 8412
rect 34388 8372 34394 8384
rect 34514 8372 34520 8384
rect 34572 8412 34578 8424
rect 34885 8415 34943 8421
rect 34885 8412 34897 8415
rect 34572 8384 34897 8412
rect 34572 8372 34578 8384
rect 34885 8381 34897 8384
rect 34931 8381 34943 8415
rect 36096 8412 36124 8452
rect 36541 8415 36599 8421
rect 36541 8412 36553 8415
rect 36096 8384 36553 8412
rect 34885 8375 34943 8381
rect 36541 8381 36553 8384
rect 36587 8381 36599 8415
rect 36541 8375 36599 8381
rect 37277 8415 37335 8421
rect 37277 8381 37289 8415
rect 37323 8412 37335 8415
rect 37826 8412 37832 8424
rect 37323 8384 37832 8412
rect 37323 8381 37335 8384
rect 37277 8375 37335 8381
rect 37826 8372 37832 8384
rect 37884 8372 37890 8424
rect 38378 8412 38384 8424
rect 38339 8384 38384 8412
rect 38378 8372 38384 8384
rect 38436 8372 38442 8424
rect 34238 8344 34244 8356
rect 23952 8316 24808 8344
rect 33428 8316 34244 8344
rect 4982 8276 4988 8288
rect 4540 8248 4988 8276
rect 4982 8236 4988 8248
rect 5040 8236 5046 8288
rect 10321 8279 10379 8285
rect 10321 8245 10333 8279
rect 10367 8276 10379 8279
rect 12526 8276 12532 8288
rect 10367 8248 12532 8276
rect 10367 8245 10379 8248
rect 10321 8239 10379 8245
rect 12526 8236 12532 8248
rect 12584 8236 12590 8288
rect 13446 8236 13452 8288
rect 13504 8276 13510 8288
rect 18782 8276 18788 8288
rect 13504 8248 18788 8276
rect 13504 8236 13510 8248
rect 18782 8236 18788 8248
rect 18840 8236 18846 8288
rect 24780 8276 24808 8316
rect 34238 8304 34244 8316
rect 34296 8304 34302 8356
rect 36814 8304 36820 8356
rect 36872 8344 36878 8356
rect 36872 8316 36938 8344
rect 36872 8304 36878 8316
rect 25866 8276 25872 8288
rect 24780 8248 25872 8276
rect 25866 8236 25872 8248
rect 25924 8236 25930 8288
rect 33318 8236 33324 8288
rect 33376 8276 33382 8288
rect 35069 8279 35127 8285
rect 35069 8276 35081 8279
rect 33376 8248 35081 8276
rect 33376 8236 33382 8248
rect 35069 8245 35081 8248
rect 35115 8245 35127 8279
rect 35069 8239 35127 8245
rect 1104 8186 39836 8208
rect 1104 8134 19606 8186
rect 19658 8134 19670 8186
rect 19722 8134 19734 8186
rect 19786 8134 19798 8186
rect 19850 8134 39836 8186
rect 1104 8112 39836 8134
rect 8662 8072 8668 8084
rect 8623 8044 8668 8072
rect 8662 8032 8668 8044
rect 8720 8032 8726 8084
rect 16666 8072 16672 8084
rect 8772 8044 15792 8072
rect 16579 8044 16672 8072
rect 4614 8004 4620 8016
rect 4080 7976 4620 8004
rect 4080 7945 4108 7976
rect 4614 7964 4620 7976
rect 4672 7964 4678 8016
rect 7834 7964 7840 8016
rect 7892 8004 7898 8016
rect 8772 8004 8800 8044
rect 7892 7976 8800 8004
rect 14461 8007 14519 8013
rect 7892 7964 7898 7976
rect 14461 7973 14473 8007
rect 14507 8004 14519 8007
rect 15562 8004 15568 8016
rect 14507 7976 15568 8004
rect 14507 7973 14519 7976
rect 14461 7967 14519 7973
rect 15562 7964 15568 7976
rect 15620 7964 15626 8016
rect 4065 7939 4123 7945
rect 4065 7905 4077 7939
rect 4111 7905 4123 7939
rect 4065 7899 4123 7905
rect 4154 7896 4160 7948
rect 4212 7936 4218 7948
rect 4525 7939 4583 7945
rect 4525 7936 4537 7939
rect 4212 7908 4537 7936
rect 4212 7896 4218 7908
rect 4525 7905 4537 7908
rect 4571 7905 4583 7939
rect 4798 7936 4804 7948
rect 4759 7908 4804 7936
rect 4525 7899 4583 7905
rect 4798 7896 4804 7908
rect 4856 7936 4862 7948
rect 5350 7936 5356 7948
rect 4856 7908 5356 7936
rect 4856 7896 4862 7908
rect 5350 7896 5356 7908
rect 5408 7896 5414 7948
rect 5445 7939 5503 7945
rect 5445 7905 5457 7939
rect 5491 7936 5503 7939
rect 5902 7936 5908 7948
rect 5491 7908 5908 7936
rect 5491 7905 5503 7908
rect 5445 7899 5503 7905
rect 5902 7896 5908 7908
rect 5960 7896 5966 7948
rect 5997 7939 6055 7945
rect 5997 7905 6009 7939
rect 6043 7936 6055 7939
rect 6086 7936 6092 7948
rect 6043 7908 6092 7936
rect 6043 7905 6055 7908
rect 5997 7899 6055 7905
rect 6086 7896 6092 7908
rect 6144 7896 6150 7948
rect 6454 7936 6460 7948
rect 6415 7908 6460 7936
rect 6454 7896 6460 7908
rect 6512 7896 6518 7948
rect 6733 7939 6791 7945
rect 6733 7905 6745 7939
rect 6779 7936 6791 7939
rect 7190 7936 7196 7948
rect 6779 7908 7196 7936
rect 6779 7905 6791 7908
rect 6733 7899 6791 7905
rect 7190 7896 7196 7908
rect 7248 7896 7254 7948
rect 8113 7939 8171 7945
rect 8113 7905 8125 7939
rect 8159 7936 8171 7939
rect 8573 7939 8631 7945
rect 8573 7936 8585 7939
rect 8159 7908 8585 7936
rect 8159 7905 8171 7908
rect 8113 7899 8171 7905
rect 8573 7905 8585 7908
rect 8619 7905 8631 7939
rect 8573 7899 8631 7905
rect 9677 7939 9735 7945
rect 9677 7905 9689 7939
rect 9723 7936 9735 7939
rect 10042 7936 10048 7948
rect 9723 7908 10048 7936
rect 9723 7905 9735 7908
rect 9677 7899 9735 7905
rect 10042 7896 10048 7908
rect 10100 7896 10106 7948
rect 11977 7939 12035 7945
rect 11977 7905 11989 7939
rect 12023 7936 12035 7939
rect 12066 7936 12072 7948
rect 12023 7908 12072 7936
rect 12023 7905 12035 7908
rect 11977 7899 12035 7905
rect 12066 7896 12072 7908
rect 12124 7896 12130 7948
rect 12434 7896 12440 7948
rect 12492 7936 12498 7948
rect 12492 7908 12537 7936
rect 12492 7896 12498 7908
rect 12986 7896 12992 7948
rect 13044 7936 13050 7948
rect 13725 7939 13783 7945
rect 13725 7936 13737 7939
rect 13044 7908 13737 7936
rect 13044 7896 13050 7908
rect 13725 7905 13737 7908
rect 13771 7905 13783 7939
rect 14182 7936 14188 7948
rect 14143 7908 14188 7936
rect 13725 7899 13783 7905
rect 14182 7896 14188 7908
rect 14240 7896 14246 7948
rect 15470 7936 15476 7948
rect 15431 7908 15476 7936
rect 15470 7896 15476 7908
rect 15528 7896 15534 7948
rect 15764 7945 15792 8044
rect 16666 8032 16672 8044
rect 16724 8072 16730 8084
rect 16942 8072 16948 8084
rect 16724 8044 16948 8072
rect 16724 8032 16730 8044
rect 16942 8032 16948 8044
rect 17000 8072 17006 8084
rect 18874 8072 18880 8084
rect 17000 8044 18880 8072
rect 17000 8032 17006 8044
rect 18874 8032 18880 8044
rect 18932 8032 18938 8084
rect 22002 8032 22008 8084
rect 22060 8072 22066 8084
rect 22465 8075 22523 8081
rect 22465 8072 22477 8075
rect 22060 8044 22477 8072
rect 22060 8032 22066 8044
rect 22465 8041 22477 8044
rect 22511 8041 22523 8075
rect 22465 8035 22523 8041
rect 25133 8075 25191 8081
rect 25133 8041 25145 8075
rect 25179 8041 25191 8075
rect 25866 8072 25872 8084
rect 25827 8044 25872 8072
rect 25133 8035 25191 8041
rect 16025 8007 16083 8013
rect 16025 7973 16037 8007
rect 16071 8004 16083 8007
rect 16114 8004 16120 8016
rect 16071 7976 16120 8004
rect 16071 7973 16083 7976
rect 16025 7967 16083 7973
rect 16114 7964 16120 7976
rect 16172 7964 16178 8016
rect 19150 8004 19156 8016
rect 16868 7976 19156 8004
rect 15749 7939 15807 7945
rect 15749 7905 15761 7939
rect 15795 7905 15807 7939
rect 15749 7899 15807 7905
rect 15930 7896 15936 7948
rect 15988 7936 15994 7948
rect 16868 7945 16896 7976
rect 19150 7964 19156 7976
rect 19208 7964 19214 8016
rect 24762 7964 24768 8016
rect 24820 8004 24826 8016
rect 25148 8004 25176 8035
rect 25866 8032 25872 8044
rect 25924 8032 25930 8084
rect 27522 8072 27528 8084
rect 26160 8044 27528 8072
rect 26160 8004 26188 8044
rect 27522 8032 27528 8044
rect 27580 8032 27586 8084
rect 27706 8072 27712 8084
rect 27667 8044 27712 8072
rect 27706 8032 27712 8044
rect 27764 8032 27770 8084
rect 29362 8072 29368 8084
rect 29323 8044 29368 8072
rect 29362 8032 29368 8044
rect 29420 8032 29426 8084
rect 31294 8072 31300 8084
rect 31255 8044 31300 8072
rect 31294 8032 31300 8044
rect 31352 8032 31358 8084
rect 33870 8032 33876 8084
rect 33928 8072 33934 8084
rect 35805 8075 35863 8081
rect 35805 8072 35817 8075
rect 33928 8044 35817 8072
rect 33928 8032 33934 8044
rect 35805 8041 35817 8044
rect 35851 8041 35863 8075
rect 35805 8035 35863 8041
rect 28445 8007 28503 8013
rect 28445 8004 28457 8007
rect 24820 7976 26188 8004
rect 26436 7976 28457 8004
rect 24820 7964 24826 7976
rect 16853 7939 16911 7945
rect 16853 7936 16865 7939
rect 15988 7908 16865 7936
rect 15988 7896 15994 7908
rect 16853 7905 16865 7908
rect 16899 7905 16911 7939
rect 16853 7899 16911 7905
rect 16945 7939 17003 7945
rect 16945 7905 16957 7939
rect 16991 7905 17003 7939
rect 16945 7899 17003 7905
rect 1394 7868 1400 7880
rect 1355 7840 1400 7868
rect 1394 7828 1400 7840
rect 1452 7828 1458 7880
rect 1673 7871 1731 7877
rect 1673 7837 1685 7871
rect 1719 7868 1731 7871
rect 2498 7868 2504 7880
rect 1719 7840 2504 7868
rect 1719 7837 1731 7840
rect 1673 7831 1731 7837
rect 2498 7828 2504 7840
rect 2556 7828 2562 7880
rect 9950 7868 9956 7880
rect 9911 7840 9956 7868
rect 9950 7828 9956 7840
rect 10008 7828 10014 7880
rect 12621 7871 12679 7877
rect 12621 7868 12633 7871
rect 10612 7840 12633 7868
rect 3510 7760 3516 7812
rect 3568 7800 3574 7812
rect 4157 7803 4215 7809
rect 4157 7800 4169 7803
rect 3568 7772 4169 7800
rect 3568 7760 3574 7772
rect 4157 7769 4169 7772
rect 4203 7769 4215 7803
rect 4157 7763 4215 7769
rect 2958 7732 2964 7744
rect 2919 7704 2964 7732
rect 2958 7692 2964 7704
rect 3016 7692 3022 7744
rect 4982 7692 4988 7744
rect 5040 7732 5046 7744
rect 10612 7732 10640 7840
rect 12621 7837 12633 7840
rect 12667 7837 12679 7871
rect 12621 7831 12679 7837
rect 13541 7871 13599 7877
rect 13541 7837 13553 7871
rect 13587 7868 13599 7871
rect 15286 7868 15292 7880
rect 13587 7840 15292 7868
rect 13587 7837 13599 7840
rect 13541 7831 13599 7837
rect 15286 7828 15292 7840
rect 15344 7828 15350 7880
rect 15378 7828 15384 7880
rect 15436 7868 15442 7880
rect 16482 7868 16488 7880
rect 15436 7840 16488 7868
rect 15436 7828 15442 7840
rect 16482 7828 16488 7840
rect 16540 7868 16546 7880
rect 16960 7868 16988 7899
rect 17218 7896 17224 7948
rect 17276 7936 17282 7948
rect 17313 7939 17371 7945
rect 17313 7936 17325 7939
rect 17276 7908 17325 7936
rect 17276 7896 17282 7908
rect 17313 7905 17325 7908
rect 17359 7905 17371 7939
rect 17313 7899 17371 7905
rect 17494 7896 17500 7948
rect 17552 7936 17558 7948
rect 17681 7939 17739 7945
rect 17681 7936 17693 7939
rect 17552 7908 17693 7936
rect 17552 7896 17558 7908
rect 17681 7905 17693 7908
rect 17727 7905 17739 7939
rect 18782 7936 18788 7948
rect 18743 7908 18788 7936
rect 17681 7899 17739 7905
rect 18782 7896 18788 7908
rect 18840 7896 18846 7948
rect 18874 7896 18880 7948
rect 18932 7936 18938 7948
rect 19613 7939 19671 7945
rect 18932 7908 19288 7936
rect 18932 7896 18938 7908
rect 16540 7840 16988 7868
rect 19153 7871 19211 7877
rect 16540 7828 16546 7840
rect 19153 7837 19165 7871
rect 19199 7837 19211 7871
rect 19260 7868 19288 7908
rect 19613 7905 19625 7939
rect 19659 7936 19671 7939
rect 19794 7936 19800 7948
rect 19659 7908 19800 7936
rect 19659 7905 19671 7908
rect 19613 7899 19671 7905
rect 19794 7896 19800 7908
rect 19852 7896 19858 7948
rect 19978 7936 19984 7948
rect 19939 7908 19984 7936
rect 19978 7896 19984 7908
rect 20036 7896 20042 7948
rect 21361 7939 21419 7945
rect 21361 7905 21373 7939
rect 21407 7936 21419 7939
rect 22094 7936 22100 7948
rect 21407 7908 22100 7936
rect 21407 7905 21419 7908
rect 21361 7899 21419 7905
rect 22094 7896 22100 7908
rect 22152 7896 22158 7948
rect 23290 7936 23296 7948
rect 23251 7908 23296 7936
rect 23290 7896 23296 7908
rect 23348 7896 23354 7948
rect 23937 7939 23995 7945
rect 23937 7905 23949 7939
rect 23983 7936 23995 7939
rect 24026 7936 24032 7948
rect 23983 7908 24032 7936
rect 23983 7905 23995 7908
rect 23937 7899 23995 7905
rect 24026 7896 24032 7908
rect 24084 7896 24090 7948
rect 24305 7939 24363 7945
rect 24305 7905 24317 7939
rect 24351 7936 24363 7939
rect 24670 7936 24676 7948
rect 24351 7908 24676 7936
rect 24351 7905 24363 7908
rect 24305 7899 24363 7905
rect 24670 7896 24676 7908
rect 24728 7896 24734 7948
rect 24949 7939 25007 7945
rect 24949 7905 24961 7939
rect 24995 7936 25007 7939
rect 25406 7936 25412 7948
rect 24995 7908 25412 7936
rect 24995 7905 25007 7908
rect 24949 7899 25007 7905
rect 25406 7896 25412 7908
rect 25464 7936 25470 7948
rect 25685 7939 25743 7945
rect 25685 7936 25697 7939
rect 25464 7908 25697 7936
rect 25464 7896 25470 7908
rect 25685 7905 25697 7908
rect 25731 7905 25743 7939
rect 25685 7899 25743 7905
rect 21085 7871 21143 7877
rect 21085 7868 21097 7871
rect 19260 7840 21097 7868
rect 19153 7831 19211 7837
rect 21085 7837 21097 7840
rect 21131 7868 21143 7871
rect 21266 7868 21272 7880
rect 21131 7840 21272 7868
rect 21131 7837 21143 7840
rect 21085 7831 21143 7837
rect 11054 7760 11060 7812
rect 11112 7800 11118 7812
rect 11885 7803 11943 7809
rect 11885 7800 11897 7803
rect 11112 7772 11897 7800
rect 11112 7760 11118 7772
rect 11885 7769 11897 7772
rect 11931 7769 11943 7803
rect 11885 7763 11943 7769
rect 11974 7760 11980 7812
rect 12032 7800 12038 7812
rect 19168 7800 19196 7831
rect 21266 7828 21272 7840
rect 21324 7828 21330 7880
rect 21450 7828 21456 7880
rect 21508 7868 21514 7880
rect 26436 7868 26464 7976
rect 26697 7939 26755 7945
rect 26697 7905 26709 7939
rect 26743 7936 26755 7939
rect 27062 7936 27068 7948
rect 26743 7908 27068 7936
rect 26743 7905 26755 7908
rect 26697 7899 26755 7905
rect 27062 7896 27068 7908
rect 27120 7896 27126 7948
rect 27172 7945 27200 7976
rect 28445 7973 28457 7976
rect 28491 7973 28503 8007
rect 28445 7967 28503 7973
rect 33781 8007 33839 8013
rect 33781 7973 33793 8007
rect 33827 8004 33839 8007
rect 34330 8004 34336 8016
rect 33827 7976 34336 8004
rect 33827 7973 33839 7976
rect 33781 7967 33839 7973
rect 34330 7964 34336 7976
rect 34388 7964 34394 8016
rect 34422 7964 34428 8016
rect 34480 8004 34486 8016
rect 34480 7976 35756 8004
rect 34480 7964 34486 7976
rect 27157 7939 27215 7945
rect 27157 7905 27169 7939
rect 27203 7905 27215 7939
rect 27157 7899 27215 7905
rect 27249 7939 27307 7945
rect 27249 7905 27261 7939
rect 27295 7936 27307 7939
rect 27430 7936 27436 7948
rect 27295 7908 27436 7936
rect 27295 7905 27307 7908
rect 27249 7899 27307 7905
rect 27430 7896 27436 7908
rect 27488 7896 27494 7948
rect 28350 7936 28356 7948
rect 28311 7908 28356 7936
rect 28350 7896 28356 7908
rect 28408 7896 28414 7948
rect 29270 7936 29276 7948
rect 29231 7908 29276 7936
rect 29270 7896 29276 7908
rect 29328 7896 29334 7948
rect 32125 7939 32183 7945
rect 32125 7905 32137 7939
rect 32171 7936 32183 7939
rect 33502 7936 33508 7948
rect 32171 7908 33508 7936
rect 32171 7905 32183 7908
rect 32125 7899 32183 7905
rect 33502 7896 33508 7908
rect 33560 7896 33566 7948
rect 35069 7939 35127 7945
rect 35069 7905 35081 7939
rect 35115 7936 35127 7939
rect 35342 7936 35348 7948
rect 35115 7908 35348 7936
rect 35115 7905 35127 7908
rect 35069 7899 35127 7905
rect 35342 7896 35348 7908
rect 35400 7896 35406 7948
rect 35728 7945 35756 7976
rect 35713 7939 35771 7945
rect 35713 7905 35725 7939
rect 35759 7905 35771 7939
rect 35713 7899 35771 7905
rect 21508 7840 26464 7868
rect 26605 7871 26663 7877
rect 21508 7828 21514 7840
rect 26605 7837 26617 7871
rect 26651 7837 26663 7871
rect 26605 7831 26663 7837
rect 12032 7772 19196 7800
rect 12032 7760 12038 7772
rect 5040 7704 10640 7732
rect 11241 7735 11299 7741
rect 5040 7692 5046 7704
rect 11241 7701 11253 7735
rect 11287 7732 11299 7735
rect 11514 7732 11520 7744
rect 11287 7704 11520 7732
rect 11287 7701 11299 7704
rect 11241 7695 11299 7701
rect 11514 7692 11520 7704
rect 11572 7692 11578 7744
rect 17034 7732 17040 7744
rect 16995 7704 17040 7732
rect 17034 7692 17040 7704
rect 17092 7692 17098 7744
rect 17586 7692 17592 7744
rect 17644 7732 17650 7744
rect 17862 7732 17868 7744
rect 17644 7704 17868 7732
rect 17644 7692 17650 7704
rect 17862 7692 17868 7704
rect 17920 7692 17926 7744
rect 18601 7735 18659 7741
rect 18601 7701 18613 7735
rect 18647 7732 18659 7735
rect 19058 7732 19064 7744
rect 18647 7704 19064 7732
rect 18647 7701 18659 7704
rect 18601 7695 18659 7701
rect 19058 7692 19064 7704
rect 19116 7692 19122 7744
rect 19168 7732 19196 7772
rect 19242 7760 19248 7812
rect 19300 7800 19306 7812
rect 19889 7803 19947 7809
rect 19889 7800 19901 7803
rect 19300 7772 19901 7800
rect 19300 7760 19306 7772
rect 19889 7769 19901 7772
rect 19935 7769 19947 7803
rect 23382 7800 23388 7812
rect 23343 7772 23388 7800
rect 19889 7763 19947 7769
rect 23382 7760 23388 7772
rect 23440 7760 23446 7812
rect 26620 7800 26648 7831
rect 29086 7828 29092 7880
rect 29144 7868 29150 7880
rect 29917 7871 29975 7877
rect 29917 7868 29929 7871
rect 29144 7840 29929 7868
rect 29144 7828 29150 7840
rect 29917 7837 29929 7840
rect 29963 7837 29975 7871
rect 29917 7831 29975 7837
rect 30193 7871 30251 7877
rect 30193 7837 30205 7871
rect 30239 7868 30251 7871
rect 30558 7868 30564 7880
rect 30239 7840 30564 7868
rect 30239 7837 30251 7840
rect 30193 7831 30251 7837
rect 30558 7828 30564 7840
rect 30616 7828 30622 7880
rect 32398 7868 32404 7880
rect 32359 7840 32404 7868
rect 32398 7828 32404 7840
rect 32456 7828 32462 7880
rect 33686 7828 33692 7880
rect 33744 7868 33750 7880
rect 34241 7871 34299 7877
rect 34241 7868 34253 7871
rect 33744 7840 34253 7868
rect 33744 7828 33750 7840
rect 34241 7837 34253 7840
rect 34287 7837 34299 7871
rect 34790 7868 34796 7880
rect 34751 7840 34796 7868
rect 34241 7831 34299 7837
rect 34790 7828 34796 7840
rect 34848 7828 34854 7880
rect 35253 7871 35311 7877
rect 35253 7837 35265 7871
rect 35299 7868 35311 7871
rect 36078 7868 36084 7880
rect 35299 7840 36084 7868
rect 35299 7837 35311 7840
rect 35253 7831 35311 7837
rect 36078 7828 36084 7840
rect 36136 7828 36142 7880
rect 28166 7800 28172 7812
rect 26620 7772 28172 7800
rect 28166 7760 28172 7772
rect 28224 7760 28230 7812
rect 21818 7732 21824 7744
rect 19168 7704 21824 7732
rect 21818 7692 21824 7704
rect 21876 7692 21882 7744
rect 22462 7692 22468 7744
rect 22520 7732 22526 7744
rect 25314 7732 25320 7744
rect 22520 7704 25320 7732
rect 22520 7692 22526 7704
rect 25314 7692 25320 7704
rect 25372 7692 25378 7744
rect 29454 7692 29460 7744
rect 29512 7732 29518 7744
rect 36262 7732 36268 7744
rect 29512 7704 36268 7732
rect 29512 7692 29518 7704
rect 36262 7692 36268 7704
rect 36320 7692 36326 7744
rect 1104 7642 39836 7664
rect 1104 7590 4246 7642
rect 4298 7590 4310 7642
rect 4362 7590 4374 7642
rect 4426 7590 4438 7642
rect 4490 7590 34966 7642
rect 35018 7590 35030 7642
rect 35082 7590 35094 7642
rect 35146 7590 35158 7642
rect 35210 7590 39836 7642
rect 1104 7568 39836 7590
rect 4890 7528 4896 7540
rect 2516 7500 4896 7528
rect 2314 7324 2320 7336
rect 2275 7296 2320 7324
rect 2314 7284 2320 7296
rect 2372 7284 2378 7336
rect 2516 7333 2544 7500
rect 4890 7488 4896 7500
rect 4948 7488 4954 7540
rect 6086 7488 6092 7540
rect 6144 7528 6150 7540
rect 6546 7528 6552 7540
rect 6144 7500 6552 7528
rect 6144 7488 6150 7500
rect 6546 7488 6552 7500
rect 6604 7528 6610 7540
rect 7009 7531 7067 7537
rect 7009 7528 7021 7531
rect 6604 7500 7021 7528
rect 6604 7488 6610 7500
rect 7009 7497 7021 7500
rect 7055 7497 7067 7531
rect 7009 7491 7067 7497
rect 7098 7488 7104 7540
rect 7156 7528 7162 7540
rect 8573 7531 8631 7537
rect 8573 7528 8585 7531
rect 7156 7500 8585 7528
rect 7156 7488 7162 7500
rect 8573 7497 8585 7500
rect 8619 7497 8631 7531
rect 8573 7491 8631 7497
rect 4614 7420 4620 7472
rect 4672 7460 4678 7472
rect 5537 7463 5595 7469
rect 5537 7460 5549 7463
rect 4672 7432 5549 7460
rect 4672 7420 4678 7432
rect 5537 7429 5549 7432
rect 5583 7429 5595 7463
rect 7834 7460 7840 7472
rect 7795 7432 7840 7460
rect 5537 7423 5595 7429
rect 7834 7420 7840 7432
rect 7892 7420 7898 7472
rect 3510 7392 3516 7404
rect 3471 7364 3516 7392
rect 3510 7352 3516 7364
rect 3568 7352 3574 7404
rect 4893 7395 4951 7401
rect 4893 7361 4905 7395
rect 4939 7392 4951 7395
rect 4982 7392 4988 7404
rect 4939 7364 4988 7392
rect 4939 7361 4951 7364
rect 4893 7355 4951 7361
rect 4982 7352 4988 7364
rect 5040 7352 5046 7404
rect 2501 7327 2559 7333
rect 2501 7293 2513 7327
rect 2547 7293 2559 7327
rect 2501 7287 2559 7293
rect 3237 7327 3295 7333
rect 3237 7293 3249 7327
rect 3283 7324 3295 7327
rect 5166 7324 5172 7336
rect 3283 7296 5172 7324
rect 3283 7293 3295 7296
rect 3237 7287 3295 7293
rect 5166 7284 5172 7296
rect 5224 7284 5230 7336
rect 5258 7284 5264 7336
rect 5316 7324 5322 7336
rect 5353 7327 5411 7333
rect 5353 7324 5365 7327
rect 5316 7296 5365 7324
rect 5316 7284 5322 7296
rect 5353 7293 5365 7296
rect 5399 7293 5411 7327
rect 5353 7287 5411 7293
rect 6825 7327 6883 7333
rect 6825 7293 6837 7327
rect 6871 7324 6883 7327
rect 7466 7324 7472 7336
rect 6871 7296 7472 7324
rect 6871 7293 6883 7296
rect 6825 7287 6883 7293
rect 7466 7284 7472 7296
rect 7524 7284 7530 7336
rect 7745 7327 7803 7333
rect 7745 7293 7757 7327
rect 7791 7324 7803 7327
rect 8294 7324 8300 7336
rect 7791 7296 8300 7324
rect 7791 7293 7803 7296
rect 7745 7287 7803 7293
rect 8294 7284 8300 7296
rect 8352 7284 8358 7336
rect 8386 7284 8392 7336
rect 8444 7324 8450 7336
rect 8588 7324 8616 7491
rect 11238 7488 11244 7540
rect 11296 7528 11302 7540
rect 12805 7531 12863 7537
rect 12805 7528 12817 7531
rect 11296 7500 12817 7528
rect 11296 7488 11302 7500
rect 12805 7497 12817 7500
rect 12851 7497 12863 7531
rect 12805 7491 12863 7497
rect 15473 7531 15531 7537
rect 15473 7497 15485 7531
rect 15519 7528 15531 7531
rect 15930 7528 15936 7540
rect 15519 7500 15936 7528
rect 15519 7497 15531 7500
rect 15473 7491 15531 7497
rect 15930 7488 15936 7500
rect 15988 7488 15994 7540
rect 16482 7488 16488 7540
rect 16540 7528 16546 7540
rect 17129 7531 17187 7537
rect 17129 7528 17141 7531
rect 16540 7500 17141 7528
rect 16540 7488 16546 7500
rect 17129 7497 17141 7500
rect 17175 7497 17187 7531
rect 24762 7528 24768 7540
rect 17129 7491 17187 7497
rect 18248 7500 24768 7528
rect 14182 7460 14188 7472
rect 14143 7432 14188 7460
rect 14182 7420 14188 7432
rect 14240 7420 14246 7472
rect 9950 7392 9956 7404
rect 9911 7364 9956 7392
rect 9950 7352 9956 7364
rect 10008 7352 10014 7404
rect 11974 7392 11980 7404
rect 10520 7364 11980 7392
rect 9125 7327 9183 7333
rect 9125 7324 9137 7327
rect 8444 7296 8489 7324
rect 8588 7296 9137 7324
rect 8444 7284 8450 7296
rect 9125 7293 9137 7296
rect 9171 7293 9183 7327
rect 9125 7287 9183 7293
rect 9769 7327 9827 7333
rect 9769 7293 9781 7327
rect 9815 7293 9827 7327
rect 9769 7287 9827 7293
rect 9784 7256 9812 7287
rect 9858 7284 9864 7336
rect 9916 7324 9922 7336
rect 10520 7333 10548 7364
rect 11974 7352 11980 7364
rect 12032 7352 12038 7404
rect 12066 7352 12072 7404
rect 12124 7392 12130 7404
rect 12124 7364 13216 7392
rect 12124 7352 12130 7364
rect 10505 7327 10563 7333
rect 9916 7296 9961 7324
rect 9916 7284 9922 7296
rect 10505 7293 10517 7327
rect 10551 7293 10563 7327
rect 10778 7324 10784 7336
rect 10739 7296 10784 7324
rect 10505 7287 10563 7293
rect 10778 7284 10784 7296
rect 10836 7284 10842 7336
rect 11514 7324 11520 7336
rect 11475 7296 11520 7324
rect 11514 7284 11520 7296
rect 11572 7284 11578 7336
rect 12989 7327 13047 7333
rect 12989 7293 13001 7327
rect 13035 7293 13047 7327
rect 13188 7324 13216 7364
rect 13722 7352 13728 7404
rect 13780 7392 13786 7404
rect 14921 7395 14979 7401
rect 13780 7364 14504 7392
rect 13780 7352 13786 7364
rect 13814 7324 13820 7336
rect 13188 7296 13820 7324
rect 12989 7287 13047 7293
rect 10594 7256 10600 7268
rect 9784 7228 10600 7256
rect 10594 7216 10600 7228
rect 10652 7256 10658 7268
rect 11609 7259 11667 7265
rect 11609 7256 11621 7259
rect 10652 7228 11621 7256
rect 10652 7216 10658 7228
rect 11609 7225 11621 7228
rect 11655 7225 11667 7259
rect 13004 7256 13032 7287
rect 13814 7284 13820 7296
rect 13872 7324 13878 7336
rect 13998 7324 14004 7336
rect 13872 7296 14004 7324
rect 13872 7284 13878 7296
rect 13998 7284 14004 7296
rect 14056 7284 14062 7336
rect 14476 7333 14504 7364
rect 14921 7361 14933 7395
rect 14967 7392 14979 7395
rect 18138 7392 18144 7404
rect 14967 7364 18144 7392
rect 14967 7361 14979 7364
rect 14921 7355 14979 7361
rect 18138 7352 18144 7364
rect 18196 7352 18202 7404
rect 14461 7327 14519 7333
rect 14461 7293 14473 7327
rect 14507 7293 14519 7327
rect 14461 7287 14519 7293
rect 15657 7327 15715 7333
rect 15657 7293 15669 7327
rect 15703 7293 15715 7327
rect 15657 7287 15715 7293
rect 15749 7327 15807 7333
rect 15749 7293 15761 7327
rect 15795 7324 15807 7327
rect 16025 7327 16083 7333
rect 15795 7296 15884 7324
rect 15795 7293 15807 7296
rect 15749 7287 15807 7293
rect 14274 7256 14280 7268
rect 13004 7228 14280 7256
rect 11609 7219 11667 7225
rect 14274 7216 14280 7228
rect 14332 7256 14338 7268
rect 15672 7256 15700 7287
rect 14332 7228 15700 7256
rect 14332 7216 14338 7228
rect 1670 7148 1676 7200
rect 1728 7188 1734 7200
rect 2133 7191 2191 7197
rect 2133 7188 2145 7191
rect 1728 7160 2145 7188
rect 1728 7148 1734 7160
rect 2133 7157 2145 7160
rect 2179 7157 2191 7191
rect 15856 7188 15884 7296
rect 16025 7293 16037 7327
rect 16071 7324 16083 7327
rect 16850 7324 16856 7336
rect 16071 7296 16856 7324
rect 16071 7293 16083 7296
rect 16025 7287 16083 7293
rect 16850 7284 16856 7296
rect 16908 7284 16914 7336
rect 18248 7333 18276 7500
rect 24762 7488 24768 7500
rect 24820 7488 24826 7540
rect 25314 7488 25320 7540
rect 25372 7528 25378 7540
rect 28445 7531 28503 7537
rect 28445 7528 28457 7531
rect 25372 7500 28457 7528
rect 25372 7488 25378 7500
rect 28445 7497 28457 7500
rect 28491 7528 28503 7531
rect 33410 7528 33416 7540
rect 28491 7500 33416 7528
rect 28491 7497 28503 7500
rect 28445 7491 28503 7497
rect 33410 7488 33416 7500
rect 33468 7488 33474 7540
rect 22370 7460 22376 7472
rect 21928 7432 22140 7460
rect 22331 7432 22376 7460
rect 18874 7352 18880 7404
rect 18932 7392 18938 7404
rect 18969 7395 19027 7401
rect 18969 7392 18981 7395
rect 18932 7364 18981 7392
rect 18932 7352 18938 7364
rect 18969 7361 18981 7364
rect 19015 7361 19027 7395
rect 19242 7392 19248 7404
rect 19203 7364 19248 7392
rect 18969 7355 19027 7361
rect 19242 7352 19248 7364
rect 19300 7352 19306 7404
rect 18233 7327 18291 7333
rect 18233 7293 18245 7327
rect 18279 7293 18291 7327
rect 18233 7287 18291 7293
rect 19058 7284 19064 7336
rect 19116 7324 19122 7336
rect 21269 7327 21327 7333
rect 21269 7324 21281 7327
rect 19116 7296 21281 7324
rect 19116 7284 19122 7296
rect 21269 7293 21281 7296
rect 21315 7293 21327 7327
rect 21542 7324 21548 7336
rect 21503 7296 21548 7324
rect 21269 7287 21327 7293
rect 21542 7284 21548 7296
rect 21600 7284 21606 7336
rect 21818 7284 21824 7336
rect 21876 7324 21882 7336
rect 21928 7333 21956 7432
rect 22112 7392 22140 7432
rect 22370 7420 22376 7432
rect 22428 7420 22434 7472
rect 23753 7463 23811 7469
rect 23753 7460 23765 7463
rect 22480 7432 23765 7460
rect 22480 7392 22508 7432
rect 23753 7429 23765 7432
rect 23799 7429 23811 7463
rect 23753 7423 23811 7429
rect 23842 7420 23848 7472
rect 23900 7460 23906 7472
rect 24854 7460 24860 7472
rect 23900 7432 24860 7460
rect 23900 7420 23906 7432
rect 24854 7420 24860 7432
rect 24912 7460 24918 7472
rect 28166 7460 28172 7472
rect 24912 7432 28172 7460
rect 24912 7420 24918 7432
rect 28166 7420 28172 7432
rect 28224 7420 28230 7472
rect 30834 7420 30840 7472
rect 30892 7460 30898 7472
rect 30892 7432 33180 7460
rect 30892 7420 30898 7432
rect 25409 7395 25467 7401
rect 25409 7392 25421 7395
rect 22112 7364 22508 7392
rect 22572 7364 25421 7392
rect 21913 7327 21971 7333
rect 21913 7324 21925 7327
rect 21876 7296 21925 7324
rect 21876 7284 21882 7296
rect 21913 7293 21925 7296
rect 21959 7293 21971 7327
rect 22462 7324 22468 7336
rect 22423 7296 22468 7324
rect 21913 7287 21971 7293
rect 22462 7284 22468 7296
rect 22520 7284 22526 7336
rect 20254 7216 20260 7268
rect 20312 7256 20318 7268
rect 22572 7256 22600 7364
rect 25409 7361 25421 7364
rect 25455 7361 25467 7395
rect 25409 7355 25467 7361
rect 29273 7395 29331 7401
rect 29273 7361 29285 7395
rect 29319 7392 29331 7395
rect 29546 7392 29552 7404
rect 29319 7364 29552 7392
rect 29319 7361 29331 7364
rect 29273 7355 29331 7361
rect 29546 7352 29552 7364
rect 29604 7352 29610 7404
rect 30285 7395 30343 7401
rect 30285 7361 30297 7395
rect 30331 7392 30343 7395
rect 31018 7392 31024 7404
rect 30331 7364 31024 7392
rect 30331 7361 30343 7364
rect 30285 7355 30343 7361
rect 31018 7352 31024 7364
rect 31076 7352 31082 7404
rect 31570 7392 31576 7404
rect 31531 7364 31576 7392
rect 31570 7352 31576 7364
rect 31628 7352 31634 7404
rect 23842 7324 23848 7336
rect 23803 7296 23848 7324
rect 23842 7284 23848 7296
rect 23900 7284 23906 7336
rect 24026 7324 24032 7336
rect 23987 7296 24032 7324
rect 24026 7284 24032 7296
rect 24084 7284 24090 7336
rect 24394 7324 24400 7336
rect 24355 7296 24400 7324
rect 24394 7284 24400 7296
rect 24452 7284 24458 7336
rect 25222 7284 25228 7336
rect 25280 7324 25286 7336
rect 25317 7327 25375 7333
rect 25317 7324 25329 7327
rect 25280 7296 25329 7324
rect 25280 7284 25286 7296
rect 25317 7293 25329 7296
rect 25363 7293 25375 7327
rect 25774 7324 25780 7336
rect 25735 7296 25780 7324
rect 25317 7287 25375 7293
rect 25774 7284 25780 7296
rect 25832 7284 25838 7336
rect 26326 7324 26332 7336
rect 26287 7296 26332 7324
rect 26326 7284 26332 7296
rect 26384 7284 26390 7336
rect 27525 7327 27583 7333
rect 27525 7293 27537 7327
rect 27571 7324 27583 7327
rect 27798 7324 27804 7336
rect 27571 7296 27804 7324
rect 27571 7293 27583 7296
rect 27525 7287 27583 7293
rect 27798 7284 27804 7296
rect 27856 7324 27862 7336
rect 28261 7327 28319 7333
rect 28261 7324 28273 7327
rect 27856 7296 28273 7324
rect 27856 7284 27862 7296
rect 28261 7293 28273 7296
rect 28307 7293 28319 7327
rect 28261 7287 28319 7293
rect 28994 7284 29000 7336
rect 29052 7324 29058 7336
rect 29825 7327 29883 7333
rect 29825 7324 29837 7327
rect 29052 7296 29837 7324
rect 29052 7284 29058 7296
rect 29825 7293 29837 7296
rect 29871 7293 29883 7327
rect 29825 7287 29883 7293
rect 30101 7327 30159 7333
rect 30101 7293 30113 7327
rect 30147 7293 30159 7327
rect 31846 7324 31852 7336
rect 31807 7296 31852 7324
rect 30101 7287 30159 7293
rect 29546 7256 29552 7268
rect 20312 7228 22600 7256
rect 24964 7228 29552 7256
rect 20312 7216 20318 7228
rect 16666 7188 16672 7200
rect 15856 7160 16672 7188
rect 2133 7151 2191 7157
rect 16666 7148 16672 7160
rect 16724 7148 16730 7200
rect 17218 7148 17224 7200
rect 17276 7188 17282 7200
rect 18417 7191 18475 7197
rect 18417 7188 18429 7191
rect 17276 7160 18429 7188
rect 17276 7148 17282 7160
rect 18417 7157 18429 7160
rect 18463 7157 18475 7191
rect 18417 7151 18475 7157
rect 19242 7148 19248 7200
rect 19300 7188 19306 7200
rect 20349 7191 20407 7197
rect 20349 7188 20361 7191
rect 19300 7160 20361 7188
rect 19300 7148 19306 7160
rect 20349 7157 20361 7160
rect 20395 7157 20407 7191
rect 20349 7151 20407 7157
rect 21085 7191 21143 7197
rect 21085 7157 21097 7191
rect 21131 7188 21143 7191
rect 21726 7188 21732 7200
rect 21131 7160 21732 7188
rect 21131 7157 21143 7160
rect 21085 7151 21143 7157
rect 21726 7148 21732 7160
rect 21784 7188 21790 7200
rect 22002 7188 22008 7200
rect 21784 7160 22008 7188
rect 21784 7148 21790 7160
rect 22002 7148 22008 7160
rect 22060 7148 22066 7200
rect 22646 7148 22652 7200
rect 22704 7188 22710 7200
rect 23934 7188 23940 7200
rect 22704 7160 23940 7188
rect 22704 7148 22710 7160
rect 23934 7148 23940 7160
rect 23992 7188 23998 7200
rect 24964 7188 24992 7228
rect 29546 7216 29552 7228
rect 29604 7216 29610 7268
rect 30116 7256 30144 7287
rect 31846 7284 31852 7296
rect 31904 7284 31910 7336
rect 32030 7324 32036 7336
rect 31991 7296 32036 7324
rect 32030 7284 32036 7296
rect 32088 7284 32094 7336
rect 33045 7327 33103 7333
rect 33045 7293 33057 7327
rect 33091 7293 33103 7327
rect 33152 7324 33180 7432
rect 35345 7395 35403 7401
rect 35345 7361 35357 7395
rect 35391 7392 35403 7395
rect 35434 7392 35440 7404
rect 35391 7364 35440 7392
rect 35391 7361 35403 7364
rect 35345 7355 35403 7361
rect 35434 7352 35440 7364
rect 35492 7352 35498 7404
rect 36722 7392 36728 7404
rect 36683 7364 36728 7392
rect 36722 7352 36728 7364
rect 36780 7352 36786 7404
rect 37366 7392 37372 7404
rect 37327 7364 37372 7392
rect 37366 7352 37372 7364
rect 37424 7352 37430 7404
rect 37642 7392 37648 7404
rect 37603 7364 37648 7392
rect 37642 7352 37648 7364
rect 37700 7352 37706 7404
rect 33318 7324 33324 7336
rect 33152 7296 33324 7324
rect 33045 7287 33103 7293
rect 30282 7256 30288 7268
rect 30116 7228 30288 7256
rect 30282 7216 30288 7228
rect 30340 7216 30346 7268
rect 31021 7259 31079 7265
rect 31021 7225 31033 7259
rect 31067 7256 31079 7259
rect 31110 7256 31116 7268
rect 31067 7228 31116 7256
rect 31067 7225 31079 7228
rect 31021 7219 31079 7225
rect 31110 7216 31116 7228
rect 31168 7216 31174 7268
rect 32493 7259 32551 7265
rect 32493 7225 32505 7259
rect 32539 7256 32551 7259
rect 32766 7256 32772 7268
rect 32539 7228 32772 7256
rect 32539 7225 32551 7228
rect 32493 7219 32551 7225
rect 32766 7216 32772 7228
rect 32824 7216 32830 7268
rect 23992 7160 24992 7188
rect 27709 7191 27767 7197
rect 23992 7148 23998 7160
rect 27709 7157 27721 7191
rect 27755 7188 27767 7191
rect 27982 7188 27988 7200
rect 27755 7160 27988 7188
rect 27755 7157 27767 7160
rect 27709 7151 27767 7157
rect 27982 7148 27988 7160
rect 28040 7188 28046 7200
rect 30926 7188 30932 7200
rect 28040 7160 30932 7188
rect 28040 7148 28046 7160
rect 30926 7148 30932 7160
rect 30984 7188 30990 7200
rect 31570 7188 31576 7200
rect 30984 7160 31576 7188
rect 30984 7148 30990 7160
rect 31570 7148 31576 7160
rect 31628 7188 31634 7200
rect 32674 7188 32680 7200
rect 31628 7160 32680 7188
rect 31628 7148 31634 7160
rect 32674 7148 32680 7160
rect 32732 7188 32738 7200
rect 33060 7188 33088 7287
rect 33318 7284 33324 7296
rect 33376 7284 33382 7336
rect 33505 7327 33563 7333
rect 33505 7293 33517 7327
rect 33551 7293 33563 7327
rect 35066 7324 35072 7336
rect 35027 7296 35072 7324
rect 33505 7287 33563 7293
rect 33520 7188 33548 7287
rect 35066 7284 35072 7296
rect 35124 7284 35130 7336
rect 33594 7188 33600 7200
rect 32732 7160 33088 7188
rect 33507 7160 33600 7188
rect 32732 7148 32738 7160
rect 33594 7148 33600 7160
rect 33652 7188 33658 7200
rect 38749 7191 38807 7197
rect 38749 7188 38761 7191
rect 33652 7160 38761 7188
rect 33652 7148 33658 7160
rect 38749 7157 38761 7160
rect 38795 7157 38807 7191
rect 38749 7151 38807 7157
rect 1104 7098 39836 7120
rect 1104 7046 19606 7098
rect 19658 7046 19670 7098
rect 19722 7046 19734 7098
rect 19786 7046 19798 7098
rect 19850 7046 39836 7098
rect 1104 7024 39836 7046
rect 8294 6944 8300 6996
rect 8352 6984 8358 6996
rect 8665 6987 8723 6993
rect 8665 6984 8677 6987
rect 8352 6956 8677 6984
rect 8352 6944 8358 6956
rect 8665 6953 8677 6956
rect 8711 6953 8723 6987
rect 8665 6947 8723 6953
rect 10318 6944 10324 6996
rect 10376 6984 10382 6996
rect 20254 6984 20260 6996
rect 10376 6956 20260 6984
rect 10376 6944 10382 6956
rect 20254 6944 20260 6956
rect 20312 6944 20318 6996
rect 22557 6987 22615 6993
rect 22557 6953 22569 6987
rect 22603 6984 22615 6987
rect 22646 6984 22652 6996
rect 22603 6956 22652 6984
rect 22603 6953 22615 6956
rect 22557 6947 22615 6953
rect 22646 6944 22652 6956
rect 22704 6944 22710 6996
rect 24670 6944 24676 6996
rect 24728 6984 24734 6996
rect 29454 6984 29460 6996
rect 24728 6956 29460 6984
rect 24728 6944 24734 6956
rect 29454 6944 29460 6956
rect 29512 6944 29518 6996
rect 29546 6944 29552 6996
rect 29604 6984 29610 6996
rect 35066 6984 35072 6996
rect 29604 6956 35072 6984
rect 29604 6944 29610 6956
rect 35066 6944 35072 6956
rect 35124 6944 35130 6996
rect 4982 6876 4988 6928
rect 5040 6916 5046 6928
rect 5040 6888 5672 6916
rect 5040 6876 5046 6888
rect 2317 6851 2375 6857
rect 2317 6817 2329 6851
rect 2363 6848 2375 6851
rect 2774 6848 2780 6860
rect 2363 6820 2780 6848
rect 2363 6817 2375 6820
rect 2317 6811 2375 6817
rect 2774 6808 2780 6820
rect 2832 6808 2838 6860
rect 4249 6851 4307 6857
rect 4249 6817 4261 6851
rect 4295 6817 4307 6851
rect 4249 6811 4307 6817
rect 2225 6783 2283 6789
rect 2225 6749 2237 6783
rect 2271 6780 2283 6783
rect 2866 6780 2872 6792
rect 2271 6752 2872 6780
rect 2271 6749 2283 6752
rect 2225 6743 2283 6749
rect 2866 6740 2872 6752
rect 2924 6740 2930 6792
rect 4264 6780 4292 6811
rect 4614 6808 4620 6860
rect 4672 6848 4678 6860
rect 5644 6857 5672 6888
rect 15286 6876 15292 6928
rect 15344 6916 15350 6928
rect 15654 6916 15660 6928
rect 15344 6888 15660 6916
rect 15344 6876 15350 6888
rect 15654 6876 15660 6888
rect 15712 6876 15718 6928
rect 16850 6916 16856 6928
rect 16811 6888 16856 6916
rect 16850 6876 16856 6888
rect 16908 6876 16914 6928
rect 17494 6876 17500 6928
rect 17552 6916 17558 6928
rect 18414 6916 18420 6928
rect 17552 6888 17816 6916
rect 18375 6888 18420 6916
rect 17552 6876 17558 6888
rect 4893 6851 4951 6857
rect 4893 6848 4905 6851
rect 4672 6820 4905 6848
rect 4672 6808 4678 6820
rect 4893 6817 4905 6820
rect 4939 6817 4951 6851
rect 4893 6811 4951 6817
rect 5537 6851 5595 6857
rect 5537 6817 5549 6851
rect 5583 6817 5595 6851
rect 5537 6811 5595 6817
rect 5629 6851 5687 6857
rect 5629 6817 5641 6851
rect 5675 6817 5687 6851
rect 6270 6848 6276 6860
rect 6231 6820 6276 6848
rect 5629 6811 5687 6817
rect 5552 6780 5580 6811
rect 6270 6808 6276 6820
rect 6328 6808 6334 6860
rect 6546 6848 6552 6860
rect 6507 6820 6552 6848
rect 6546 6808 6552 6820
rect 6604 6808 6610 6860
rect 10502 6808 10508 6860
rect 10560 6848 10566 6860
rect 10597 6851 10655 6857
rect 10597 6848 10609 6851
rect 10560 6820 10609 6848
rect 10560 6808 10566 6820
rect 10597 6817 10609 6820
rect 10643 6817 10655 6851
rect 11054 6848 11060 6860
rect 11015 6820 11060 6848
rect 10597 6811 10655 6817
rect 11054 6808 11060 6820
rect 11112 6808 11118 6860
rect 11793 6851 11851 6857
rect 11793 6817 11805 6851
rect 11839 6848 11851 6851
rect 12434 6848 12440 6860
rect 11839 6820 12440 6848
rect 11839 6817 11851 6820
rect 11793 6811 11851 6817
rect 12434 6808 12440 6820
rect 12492 6808 12498 6860
rect 13449 6851 13507 6857
rect 13449 6817 13461 6851
rect 13495 6848 13507 6851
rect 13538 6848 13544 6860
rect 13495 6820 13544 6848
rect 13495 6817 13507 6820
rect 13449 6811 13507 6817
rect 13538 6808 13544 6820
rect 13596 6848 13602 6860
rect 13909 6851 13967 6857
rect 13909 6848 13921 6851
rect 13596 6820 13921 6848
rect 13596 6808 13602 6820
rect 13909 6817 13921 6820
rect 13955 6817 13967 6851
rect 13909 6811 13967 6817
rect 14553 6851 14611 6857
rect 14553 6817 14565 6851
rect 14599 6817 14611 6851
rect 14553 6811 14611 6817
rect 16301 6851 16359 6857
rect 16301 6817 16313 6851
rect 16347 6848 16359 6851
rect 16574 6848 16580 6860
rect 16347 6820 16580 6848
rect 16347 6817 16359 6820
rect 16301 6811 16359 6817
rect 6178 6780 6184 6792
rect 4264 6752 5120 6780
rect 5552 6752 6184 6780
rect 4890 6672 4896 6724
rect 4948 6712 4954 6724
rect 4985 6715 5043 6721
rect 4985 6712 4997 6715
rect 4948 6684 4997 6712
rect 4948 6672 4954 6684
rect 4985 6681 4997 6684
rect 5031 6681 5043 6715
rect 5092 6712 5120 6752
rect 6178 6740 6184 6752
rect 6236 6740 6242 6792
rect 6822 6740 6828 6792
rect 6880 6780 6886 6792
rect 7285 6783 7343 6789
rect 7285 6780 7297 6783
rect 6880 6752 7297 6780
rect 6880 6740 6886 6752
rect 7285 6749 7297 6752
rect 7331 6749 7343 6783
rect 7285 6743 7343 6749
rect 7466 6740 7472 6792
rect 7524 6780 7530 6792
rect 7561 6783 7619 6789
rect 7561 6780 7573 6783
rect 7524 6752 7573 6780
rect 7524 6740 7530 6752
rect 7561 6749 7573 6752
rect 7607 6749 7619 6783
rect 7561 6743 7619 6749
rect 10413 6783 10471 6789
rect 10413 6749 10425 6783
rect 10459 6749 10471 6783
rect 11146 6780 11152 6792
rect 11107 6752 11152 6780
rect 10413 6743 10471 6749
rect 7006 6712 7012 6724
rect 5092 6684 7012 6712
rect 4985 6675 5043 6681
rect 7006 6672 7012 6684
rect 7064 6672 7070 6724
rect 10428 6712 10456 6743
rect 11146 6740 11152 6752
rect 11204 6740 11210 6792
rect 12066 6780 12072 6792
rect 12027 6752 12072 6780
rect 12066 6740 12072 6752
rect 12124 6740 12130 6792
rect 14568 6780 14596 6811
rect 16574 6808 16580 6820
rect 16632 6808 16638 6860
rect 16669 6851 16727 6857
rect 16669 6817 16681 6851
rect 16715 6848 16727 6851
rect 17034 6848 17040 6860
rect 16715 6820 17040 6848
rect 16715 6817 16727 6820
rect 16669 6811 16727 6817
rect 17034 6808 17040 6820
rect 17092 6808 17098 6860
rect 17126 6808 17132 6860
rect 17184 6848 17190 6860
rect 17586 6848 17592 6860
rect 17184 6820 17592 6848
rect 17184 6808 17190 6820
rect 17586 6808 17592 6820
rect 17644 6808 17650 6860
rect 17681 6851 17739 6857
rect 17681 6817 17693 6851
rect 17727 6817 17739 6851
rect 17788 6848 17816 6888
rect 18414 6876 18420 6888
rect 18472 6876 18478 6928
rect 19426 6876 19432 6928
rect 19484 6916 19490 6928
rect 21082 6916 21088 6928
rect 19484 6888 21088 6916
rect 19484 6876 19490 6888
rect 21082 6876 21088 6888
rect 21140 6876 21146 6928
rect 25774 6916 25780 6928
rect 23492 6888 25780 6916
rect 18049 6851 18107 6857
rect 18049 6848 18061 6851
rect 17788 6820 18061 6848
rect 17681 6811 17739 6817
rect 18049 6817 18061 6820
rect 18095 6817 18107 6851
rect 18049 6811 18107 6817
rect 15933 6783 15991 6789
rect 14568 6752 15700 6780
rect 11790 6712 11796 6724
rect 10428 6684 11796 6712
rect 11790 6672 11796 6684
rect 11848 6672 11854 6724
rect 13630 6672 13636 6724
rect 13688 6712 13694 6724
rect 14645 6715 14703 6721
rect 14645 6712 14657 6715
rect 13688 6684 14657 6712
rect 13688 6672 13694 6684
rect 14645 6681 14657 6684
rect 14691 6681 14703 6715
rect 14645 6675 14703 6681
rect 2498 6644 2504 6656
rect 2459 6616 2504 6644
rect 2498 6604 2504 6616
rect 2556 6604 2562 6656
rect 4341 6647 4399 6653
rect 4341 6613 4353 6647
rect 4387 6644 4399 6647
rect 4614 6644 4620 6656
rect 4387 6616 4620 6644
rect 4387 6613 4399 6616
rect 4341 6607 4399 6613
rect 4614 6604 4620 6616
rect 4672 6604 4678 6656
rect 7558 6604 7564 6656
rect 7616 6644 7622 6656
rect 13354 6644 13360 6656
rect 7616 6616 13360 6644
rect 7616 6604 7622 6616
rect 13354 6604 13360 6616
rect 13412 6604 13418 6656
rect 14001 6647 14059 6653
rect 14001 6613 14013 6647
rect 14047 6644 14059 6647
rect 14182 6644 14188 6656
rect 14047 6616 14188 6644
rect 14047 6613 14059 6616
rect 14001 6607 14059 6613
rect 14182 6604 14188 6616
rect 14240 6604 14246 6656
rect 15672 6644 15700 6752
rect 15933 6749 15945 6783
rect 15979 6780 15991 6783
rect 16758 6780 16764 6792
rect 15979 6752 16764 6780
rect 15979 6749 15991 6752
rect 15933 6743 15991 6749
rect 16758 6740 16764 6752
rect 16816 6740 16822 6792
rect 17218 6740 17224 6792
rect 17276 6780 17282 6792
rect 17696 6780 17724 6811
rect 18138 6808 18144 6860
rect 18196 6848 18202 6860
rect 19153 6851 19211 6857
rect 19153 6848 19165 6851
rect 18196 6820 19165 6848
rect 18196 6808 18202 6820
rect 19153 6817 19165 6820
rect 19199 6848 19211 6851
rect 19242 6848 19248 6860
rect 19199 6820 19248 6848
rect 19199 6817 19211 6820
rect 19153 6811 19211 6817
rect 19242 6808 19248 6820
rect 19300 6808 19306 6860
rect 19521 6851 19579 6857
rect 19521 6817 19533 6851
rect 19567 6817 19579 6851
rect 19521 6811 19579 6817
rect 19536 6780 19564 6811
rect 19886 6808 19892 6860
rect 19944 6848 19950 6860
rect 20073 6851 20131 6857
rect 20073 6848 20085 6851
rect 19944 6820 20085 6848
rect 19944 6808 19950 6820
rect 20073 6817 20085 6820
rect 20119 6817 20131 6851
rect 20073 6811 20131 6817
rect 19978 6780 19984 6792
rect 17276 6752 19564 6780
rect 19939 6752 19984 6780
rect 17276 6740 17282 6752
rect 19978 6740 19984 6752
rect 20036 6740 20042 6792
rect 20088 6780 20116 6811
rect 20162 6808 20168 6860
rect 20220 6848 20226 6860
rect 20622 6848 20628 6860
rect 20220 6820 20628 6848
rect 20220 6808 20226 6820
rect 20622 6808 20628 6820
rect 20680 6848 20686 6860
rect 20901 6851 20959 6857
rect 20901 6848 20913 6851
rect 20680 6820 20913 6848
rect 20680 6808 20686 6820
rect 20901 6817 20913 6820
rect 20947 6817 20959 6851
rect 20901 6811 20959 6817
rect 21545 6851 21603 6857
rect 21545 6817 21557 6851
rect 21591 6817 21603 6851
rect 21910 6848 21916 6860
rect 21871 6820 21916 6848
rect 21545 6811 21603 6817
rect 20254 6780 20260 6792
rect 20088 6752 20260 6780
rect 20254 6740 20260 6752
rect 20312 6740 20318 6792
rect 21450 6780 21456 6792
rect 21411 6752 21456 6780
rect 21450 6740 21456 6752
rect 21508 6740 21514 6792
rect 21560 6780 21588 6811
rect 21910 6808 21916 6820
rect 21968 6808 21974 6860
rect 22002 6808 22008 6860
rect 22060 6848 22066 6860
rect 22741 6851 22799 6857
rect 22741 6848 22753 6851
rect 22060 6820 22753 6848
rect 22060 6808 22066 6820
rect 22741 6817 22753 6820
rect 22787 6817 22799 6851
rect 23106 6848 23112 6860
rect 23067 6820 23112 6848
rect 22741 6811 22799 6817
rect 23106 6808 23112 6820
rect 23164 6808 23170 6860
rect 23492 6857 23520 6888
rect 25148 6860 25176 6888
rect 25774 6876 25780 6888
rect 25832 6876 25838 6928
rect 28994 6916 29000 6928
rect 28955 6888 29000 6916
rect 28994 6876 29000 6888
rect 29052 6876 29058 6928
rect 23477 6851 23535 6857
rect 23477 6817 23489 6851
rect 23523 6817 23535 6851
rect 23477 6811 23535 6817
rect 23845 6851 23903 6857
rect 23845 6817 23857 6851
rect 23891 6848 23903 6851
rect 24670 6848 24676 6860
rect 23891 6820 24676 6848
rect 23891 6817 23903 6820
rect 23845 6811 23903 6817
rect 24670 6808 24676 6820
rect 24728 6808 24734 6860
rect 24765 6851 24823 6857
rect 24765 6817 24777 6851
rect 24811 6817 24823 6851
rect 25130 6848 25136 6860
rect 25043 6820 25136 6848
rect 24765 6811 24823 6817
rect 22554 6780 22560 6792
rect 21560 6752 22560 6780
rect 22554 6740 22560 6752
rect 22612 6740 22618 6792
rect 15838 6672 15844 6724
rect 15896 6712 15902 6724
rect 22925 6715 22983 6721
rect 22925 6712 22937 6715
rect 15896 6684 22937 6712
rect 15896 6672 15902 6684
rect 22925 6681 22937 6684
rect 22971 6681 22983 6715
rect 22925 6675 22983 6681
rect 20346 6644 20352 6656
rect 15672 6616 20352 6644
rect 20346 6604 20352 6616
rect 20404 6604 20410 6656
rect 21910 6604 21916 6656
rect 21968 6644 21974 6656
rect 22186 6644 22192 6656
rect 21968 6616 22192 6644
rect 21968 6604 21974 6616
rect 22186 6604 22192 6616
rect 22244 6604 22250 6656
rect 24780 6644 24808 6811
rect 25130 6808 25136 6820
rect 25188 6808 25194 6860
rect 25501 6851 25559 6857
rect 25501 6817 25513 6851
rect 25547 6848 25559 6851
rect 26326 6848 26332 6860
rect 25547 6820 26332 6848
rect 25547 6817 25559 6820
rect 25501 6811 25559 6817
rect 26326 6808 26332 6820
rect 26384 6808 26390 6860
rect 26513 6851 26571 6857
rect 26513 6817 26525 6851
rect 26559 6817 26571 6851
rect 26513 6811 26571 6817
rect 24946 6780 24952 6792
rect 24907 6752 24952 6780
rect 24946 6740 24952 6752
rect 25004 6740 25010 6792
rect 25866 6740 25872 6792
rect 25924 6780 25930 6792
rect 26528 6780 26556 6811
rect 28166 6808 28172 6860
rect 28224 6848 28230 6860
rect 28353 6851 28411 6857
rect 28353 6848 28365 6851
rect 28224 6820 28365 6848
rect 28224 6808 28230 6820
rect 28353 6817 28365 6820
rect 28399 6817 28411 6851
rect 29822 6848 29828 6860
rect 28353 6811 28411 6817
rect 28460 6820 29592 6848
rect 29783 6820 29828 6848
rect 25924 6752 26556 6780
rect 27525 6783 27583 6789
rect 25924 6740 25930 6752
rect 27525 6749 27537 6783
rect 27571 6780 27583 6783
rect 27614 6780 27620 6792
rect 27571 6752 27620 6780
rect 27571 6749 27583 6752
rect 27525 6743 27583 6749
rect 27614 6740 27620 6752
rect 27672 6740 27678 6792
rect 28077 6783 28135 6789
rect 28077 6749 28089 6783
rect 28123 6780 28135 6783
rect 28460 6780 28488 6820
rect 28123 6752 28488 6780
rect 28537 6783 28595 6789
rect 28123 6749 28135 6752
rect 28077 6743 28135 6749
rect 28537 6749 28549 6783
rect 28583 6780 28595 6783
rect 28626 6780 28632 6792
rect 28583 6752 28632 6780
rect 28583 6749 28595 6752
rect 28537 6743 28595 6749
rect 28626 6740 28632 6752
rect 28684 6740 28690 6792
rect 29564 6789 29592 6820
rect 29822 6808 29828 6820
rect 29880 6808 29886 6860
rect 30558 6848 30564 6860
rect 30519 6820 30564 6848
rect 30558 6808 30564 6820
rect 30616 6808 30622 6860
rect 31110 6848 31116 6860
rect 31071 6820 31116 6848
rect 31110 6808 31116 6820
rect 31168 6808 31174 6860
rect 31389 6851 31447 6857
rect 31389 6817 31401 6851
rect 31435 6817 31447 6851
rect 31389 6811 31447 6817
rect 29549 6783 29607 6789
rect 29549 6749 29561 6783
rect 29595 6780 29607 6783
rect 29914 6780 29920 6792
rect 29595 6752 29920 6780
rect 29595 6749 29607 6752
rect 29549 6743 29607 6749
rect 29914 6740 29920 6752
rect 29972 6740 29978 6792
rect 30009 6783 30067 6789
rect 30009 6749 30021 6783
rect 30055 6749 30067 6783
rect 30009 6743 30067 6749
rect 28644 6712 28672 6740
rect 30024 6712 30052 6743
rect 28644 6684 30052 6712
rect 31404 6712 31432 6811
rect 32030 6808 32036 6860
rect 32088 6848 32094 6860
rect 32125 6851 32183 6857
rect 32125 6848 32137 6851
rect 32088 6820 32137 6848
rect 32088 6808 32094 6820
rect 32125 6817 32137 6820
rect 32171 6848 32183 6851
rect 33686 6848 33692 6860
rect 32171 6820 33548 6848
rect 33647 6820 33692 6848
rect 32171 6817 32183 6820
rect 32125 6811 32183 6817
rect 31573 6783 31631 6789
rect 31573 6749 31585 6783
rect 31619 6780 31631 6783
rect 31754 6780 31760 6792
rect 31619 6752 31760 6780
rect 31619 6749 31631 6752
rect 31573 6743 31631 6749
rect 31754 6740 31760 6752
rect 31812 6740 31818 6792
rect 33410 6780 33416 6792
rect 33371 6752 33416 6780
rect 33410 6740 33416 6752
rect 33468 6740 33474 6792
rect 33520 6780 33548 6820
rect 33686 6808 33692 6820
rect 33744 6808 33750 6860
rect 35805 6851 35863 6857
rect 35805 6817 35817 6851
rect 35851 6848 35863 6851
rect 36906 6848 36912 6860
rect 35851 6820 36912 6848
rect 35851 6817 35863 6820
rect 35805 6811 35863 6817
rect 36906 6808 36912 6820
rect 36964 6808 36970 6860
rect 33594 6780 33600 6792
rect 33520 6752 33600 6780
rect 33594 6740 33600 6752
rect 33652 6740 33658 6792
rect 34422 6740 34428 6792
rect 34480 6780 34486 6792
rect 35529 6783 35587 6789
rect 35529 6780 35541 6783
rect 34480 6752 35541 6780
rect 34480 6740 34486 6752
rect 35529 6749 35541 6752
rect 35575 6749 35587 6783
rect 35529 6743 35587 6749
rect 31404 6684 33456 6712
rect 26050 6644 26056 6656
rect 24780 6616 26056 6644
rect 26050 6604 26056 6616
rect 26108 6604 26114 6656
rect 26326 6604 26332 6656
rect 26384 6644 26390 6656
rect 26697 6647 26755 6653
rect 26697 6644 26709 6647
rect 26384 6616 26709 6644
rect 26384 6604 26390 6616
rect 26697 6613 26709 6616
rect 26743 6644 26755 6647
rect 27522 6644 27528 6656
rect 26743 6616 27528 6644
rect 26743 6613 26755 6616
rect 26697 6607 26755 6613
rect 27522 6604 27528 6616
rect 27580 6604 27586 6656
rect 30024 6644 30052 6684
rect 31478 6644 31484 6656
rect 30024 6616 31484 6644
rect 31478 6604 31484 6616
rect 31536 6644 31542 6656
rect 32309 6647 32367 6653
rect 32309 6644 32321 6647
rect 31536 6616 32321 6644
rect 31536 6604 31542 6616
rect 32309 6613 32321 6616
rect 32355 6613 32367 6647
rect 33428 6644 33456 6684
rect 34698 6644 34704 6656
rect 33428 6616 34704 6644
rect 32309 6607 32367 6613
rect 34698 6604 34704 6616
rect 34756 6644 34762 6656
rect 34793 6647 34851 6653
rect 34793 6644 34805 6647
rect 34756 6616 34805 6644
rect 34756 6604 34762 6616
rect 34793 6613 34805 6616
rect 34839 6613 34851 6647
rect 36906 6644 36912 6656
rect 36867 6616 36912 6644
rect 34793 6607 34851 6613
rect 36906 6604 36912 6616
rect 36964 6604 36970 6656
rect 1104 6554 39836 6576
rect 1104 6502 4246 6554
rect 4298 6502 4310 6554
rect 4362 6502 4374 6554
rect 4426 6502 4438 6554
rect 4490 6502 34966 6554
rect 35018 6502 35030 6554
rect 35082 6502 35094 6554
rect 35146 6502 35158 6554
rect 35210 6502 39836 6554
rect 1104 6480 39836 6502
rect 8110 6400 8116 6452
rect 8168 6440 8174 6452
rect 9858 6440 9864 6452
rect 8168 6412 9864 6440
rect 8168 6400 8174 6412
rect 9858 6400 9864 6412
rect 9916 6400 9922 6452
rect 10888 6412 15608 6440
rect 4706 6372 4712 6384
rect 4172 6344 4712 6372
rect 3881 6239 3939 6245
rect 3881 6205 3893 6239
rect 3927 6236 3939 6239
rect 4172 6236 4200 6344
rect 4706 6332 4712 6344
rect 4764 6332 4770 6384
rect 6270 6332 6276 6384
rect 6328 6372 6334 6384
rect 6328 6344 8248 6372
rect 6328 6332 6334 6344
rect 4338 6304 4344 6316
rect 4299 6276 4344 6304
rect 4338 6264 4344 6276
rect 4396 6264 4402 6316
rect 6546 6304 6552 6316
rect 5644 6276 6552 6304
rect 3927 6208 4200 6236
rect 4249 6239 4307 6245
rect 3927 6205 3939 6208
rect 3881 6199 3939 6205
rect 4249 6205 4261 6239
rect 4295 6205 4307 6239
rect 4249 6199 4307 6205
rect 4709 6239 4767 6245
rect 4709 6205 4721 6239
rect 4755 6236 4767 6239
rect 4982 6236 4988 6248
rect 4755 6208 4988 6236
rect 4755 6205 4767 6208
rect 4709 6199 4767 6205
rect 4264 6168 4292 6199
rect 4982 6196 4988 6208
rect 5040 6196 5046 6248
rect 5077 6239 5135 6245
rect 5077 6205 5089 6239
rect 5123 6236 5135 6239
rect 5534 6236 5540 6248
rect 5123 6208 5540 6236
rect 5123 6205 5135 6208
rect 5077 6199 5135 6205
rect 5534 6196 5540 6208
rect 5592 6196 5598 6248
rect 5644 6245 5672 6276
rect 6546 6264 6552 6276
rect 6604 6264 6610 6316
rect 7466 6304 7472 6316
rect 7427 6276 7472 6304
rect 7466 6264 7472 6276
rect 7524 6264 7530 6316
rect 5629 6239 5687 6245
rect 5629 6205 5641 6239
rect 5675 6205 5687 6239
rect 6086 6236 6092 6248
rect 6047 6208 6092 6236
rect 5629 6199 5687 6205
rect 6086 6196 6092 6208
rect 6144 6196 6150 6248
rect 7098 6236 7104 6248
rect 7059 6208 7104 6236
rect 7098 6196 7104 6208
rect 7156 6196 7162 6248
rect 7745 6239 7803 6245
rect 7745 6205 7757 6239
rect 7791 6236 7803 6239
rect 7834 6236 7840 6248
rect 7791 6208 7840 6236
rect 7791 6205 7803 6208
rect 7745 6199 7803 6205
rect 7834 6196 7840 6208
rect 7892 6196 7898 6248
rect 8110 6236 8116 6248
rect 8071 6208 8116 6236
rect 8110 6196 8116 6208
rect 8168 6196 8174 6248
rect 8220 6236 8248 6344
rect 9674 6332 9680 6384
rect 9732 6372 9738 6384
rect 10597 6375 10655 6381
rect 10597 6372 10609 6375
rect 9732 6344 10609 6372
rect 9732 6332 9738 6344
rect 10597 6341 10609 6344
rect 10643 6372 10655 6375
rect 10778 6372 10784 6384
rect 10643 6344 10784 6372
rect 10643 6341 10655 6344
rect 10597 6335 10655 6341
rect 10778 6332 10784 6344
rect 10836 6332 10842 6384
rect 9692 6304 9720 6332
rect 10888 6304 10916 6412
rect 12066 6332 12072 6384
rect 12124 6372 12130 6384
rect 12713 6375 12771 6381
rect 12713 6372 12725 6375
rect 12124 6344 12725 6372
rect 12124 6332 12130 6344
rect 12713 6341 12725 6344
rect 12759 6341 12771 6375
rect 12713 6335 12771 6341
rect 9048 6276 9720 6304
rect 9968 6276 10916 6304
rect 8294 6236 8300 6248
rect 8207 6208 8300 6236
rect 8294 6196 8300 6208
rect 8352 6196 8358 6248
rect 9048 6245 9076 6276
rect 9033 6239 9091 6245
rect 9033 6205 9045 6239
rect 9079 6205 9091 6239
rect 9033 6199 9091 6205
rect 9677 6239 9735 6245
rect 9677 6205 9689 6239
rect 9723 6236 9735 6239
rect 9858 6236 9864 6248
rect 9723 6208 9864 6236
rect 9723 6205 9735 6208
rect 9677 6199 9735 6205
rect 9858 6196 9864 6208
rect 9916 6196 9922 6248
rect 4614 6168 4620 6180
rect 4264 6140 4620 6168
rect 4614 6128 4620 6140
rect 4672 6128 4678 6180
rect 6178 6168 6184 6180
rect 6091 6140 6184 6168
rect 6178 6128 6184 6140
rect 6236 6168 6242 6180
rect 9968 6168 9996 6276
rect 10413 6239 10471 6245
rect 10413 6205 10425 6239
rect 10459 6236 10471 6239
rect 10594 6236 10600 6248
rect 10459 6208 10600 6236
rect 10459 6205 10471 6208
rect 10413 6199 10471 6205
rect 10594 6196 10600 6208
rect 10652 6196 10658 6248
rect 11146 6236 11152 6248
rect 11107 6208 11152 6236
rect 11146 6196 11152 6208
rect 11204 6196 11210 6248
rect 11241 6239 11299 6245
rect 11241 6205 11253 6239
rect 11287 6205 11299 6239
rect 11241 6199 11299 6205
rect 12805 6239 12863 6245
rect 12805 6205 12817 6239
rect 12851 6236 12863 6239
rect 13170 6236 13176 6248
rect 12851 6208 13176 6236
rect 12851 6205 12863 6208
rect 12805 6199 12863 6205
rect 6236 6140 9996 6168
rect 6236 6128 6242 6140
rect 10870 6128 10876 6180
rect 10928 6168 10934 6180
rect 11256 6168 11284 6199
rect 13170 6196 13176 6208
rect 13228 6196 13234 6248
rect 13265 6239 13323 6245
rect 13265 6205 13277 6239
rect 13311 6205 13323 6239
rect 13265 6199 13323 6205
rect 11698 6168 11704 6180
rect 10928 6140 11284 6168
rect 11659 6140 11704 6168
rect 10928 6128 10934 6140
rect 11698 6128 11704 6140
rect 11756 6128 11762 6180
rect 13280 6168 13308 6199
rect 13354 6196 13360 6248
rect 13412 6236 13418 6248
rect 13998 6236 14004 6248
rect 13412 6208 13457 6236
rect 13959 6208 14004 6236
rect 13412 6196 13418 6208
rect 13998 6196 14004 6208
rect 14056 6196 14062 6248
rect 14090 6196 14096 6248
rect 14148 6236 14154 6248
rect 14277 6239 14335 6245
rect 14277 6236 14289 6239
rect 14148 6208 14289 6236
rect 14148 6196 14154 6208
rect 14277 6205 14289 6208
rect 14323 6205 14335 6239
rect 14277 6199 14335 6205
rect 15289 6239 15347 6245
rect 15289 6205 15301 6239
rect 15335 6236 15347 6239
rect 15470 6236 15476 6248
rect 15335 6208 15476 6236
rect 15335 6205 15347 6208
rect 15289 6199 15347 6205
rect 15470 6196 15476 6208
rect 15528 6196 15534 6248
rect 15580 6245 15608 6412
rect 16040 6412 20484 6440
rect 15746 6304 15752 6316
rect 15707 6276 15752 6304
rect 15746 6264 15752 6276
rect 15804 6264 15810 6316
rect 15565 6239 15623 6245
rect 15565 6205 15577 6239
rect 15611 6205 15623 6239
rect 15565 6199 15623 6205
rect 14182 6168 14188 6180
rect 13280 6140 14188 6168
rect 14182 6128 14188 6140
rect 14240 6128 14246 6180
rect 16040 6168 16068 6412
rect 16114 6332 16120 6384
rect 16172 6372 16178 6384
rect 19426 6372 19432 6384
rect 16172 6344 19432 6372
rect 16172 6332 16178 6344
rect 19426 6332 19432 6344
rect 19484 6332 19490 6384
rect 20456 6372 20484 6412
rect 20622 6400 20628 6452
rect 20680 6440 20686 6452
rect 20901 6443 20959 6449
rect 20901 6440 20913 6443
rect 20680 6412 20913 6440
rect 20680 6400 20686 6412
rect 20901 6409 20913 6412
rect 20947 6409 20959 6443
rect 24302 6440 24308 6452
rect 20901 6403 20959 6409
rect 21008 6412 24308 6440
rect 20806 6372 20812 6384
rect 20456 6344 20812 6372
rect 20806 6332 20812 6344
rect 20864 6332 20870 6384
rect 16390 6264 16396 6316
rect 16448 6304 16454 6316
rect 21008 6304 21036 6412
rect 24302 6400 24308 6412
rect 24360 6400 24366 6452
rect 26050 6440 26056 6452
rect 26011 6412 26056 6440
rect 26050 6400 26056 6412
rect 26108 6400 26114 6452
rect 27522 6400 27528 6452
rect 27580 6400 27586 6452
rect 28166 6440 28172 6452
rect 28127 6412 28172 6440
rect 28166 6400 28172 6412
rect 28224 6400 28230 6452
rect 29454 6440 29460 6452
rect 29415 6412 29460 6440
rect 29454 6400 29460 6412
rect 29512 6400 29518 6452
rect 29914 6400 29920 6452
rect 29972 6440 29978 6452
rect 34606 6440 34612 6452
rect 29972 6412 34612 6440
rect 29972 6400 29978 6412
rect 34606 6400 34612 6412
rect 34664 6400 34670 6452
rect 23753 6375 23811 6381
rect 23753 6372 23765 6375
rect 16448 6276 21036 6304
rect 21100 6344 23765 6372
rect 16448 6264 16454 6276
rect 16574 6236 16580 6248
rect 16535 6208 16580 6236
rect 16574 6196 16580 6208
rect 16632 6196 16638 6248
rect 16666 6196 16672 6248
rect 16724 6236 16730 6248
rect 16761 6239 16819 6245
rect 16761 6236 16773 6239
rect 16724 6208 16773 6236
rect 16724 6196 16730 6208
rect 16761 6205 16773 6208
rect 16807 6205 16819 6239
rect 16761 6199 16819 6205
rect 17313 6239 17371 6245
rect 17313 6205 17325 6239
rect 17359 6236 17371 6239
rect 18414 6236 18420 6248
rect 17359 6208 18420 6236
rect 17359 6205 17371 6208
rect 17313 6199 17371 6205
rect 18414 6196 18420 6208
rect 18472 6196 18478 6248
rect 18601 6239 18659 6245
rect 18601 6205 18613 6239
rect 18647 6236 18659 6239
rect 19058 6236 19064 6248
rect 18647 6208 19064 6236
rect 18647 6205 18659 6208
rect 18601 6199 18659 6205
rect 19058 6196 19064 6208
rect 19116 6196 19122 6248
rect 19150 6196 19156 6248
rect 19208 6236 19214 6248
rect 19245 6239 19303 6245
rect 19245 6236 19257 6239
rect 19208 6208 19257 6236
rect 19208 6196 19214 6208
rect 19245 6205 19257 6208
rect 19291 6205 19303 6239
rect 19245 6199 19303 6205
rect 19521 6239 19579 6245
rect 19521 6205 19533 6239
rect 19567 6205 19579 6239
rect 19521 6199 19579 6205
rect 19797 6239 19855 6245
rect 19797 6205 19809 6239
rect 19843 6236 19855 6239
rect 20714 6236 20720 6248
rect 19843 6208 20720 6236
rect 19843 6205 19855 6208
rect 19797 6199 19855 6205
rect 14568 6140 16068 6168
rect 17497 6171 17555 6177
rect 8294 6060 8300 6112
rect 8352 6100 8358 6112
rect 14568 6100 14596 6140
rect 17497 6137 17509 6171
rect 17543 6168 17555 6171
rect 17954 6168 17960 6180
rect 17543 6140 17960 6168
rect 17543 6137 17555 6140
rect 17497 6131 17555 6137
rect 17954 6128 17960 6140
rect 18012 6128 18018 6180
rect 19536 6168 19564 6199
rect 20714 6196 20720 6208
rect 20772 6196 20778 6248
rect 20806 6196 20812 6248
rect 20864 6236 20870 6248
rect 21100 6236 21128 6344
rect 23753 6341 23765 6344
rect 23799 6341 23811 6375
rect 27540 6372 27568 6400
rect 34882 6372 34888 6384
rect 27540 6344 34888 6372
rect 23753 6335 23811 6341
rect 34882 6332 34888 6344
rect 34940 6332 34946 6384
rect 37090 6332 37096 6384
rect 37148 6372 37154 6384
rect 37148 6344 37872 6372
rect 37148 6332 37154 6344
rect 22094 6264 22100 6316
rect 22152 6304 22158 6316
rect 22462 6304 22468 6316
rect 22152 6276 22324 6304
rect 22423 6276 22468 6304
rect 22152 6264 22158 6276
rect 20864 6208 21128 6236
rect 20864 6196 20870 6208
rect 21634 6196 21640 6248
rect 21692 6236 21698 6248
rect 21821 6239 21879 6245
rect 21821 6236 21833 6239
rect 21692 6208 21833 6236
rect 21692 6196 21698 6208
rect 21821 6205 21833 6208
rect 21867 6205 21879 6239
rect 21821 6199 21879 6205
rect 22189 6239 22247 6245
rect 22189 6205 22201 6239
rect 22235 6205 22247 6239
rect 22296 6236 22324 6276
rect 22462 6264 22468 6276
rect 22520 6264 22526 6316
rect 26418 6304 26424 6316
rect 25884 6276 26424 6304
rect 22557 6239 22615 6245
rect 22557 6236 22569 6239
rect 22296 6208 22569 6236
rect 22189 6199 22247 6205
rect 22557 6205 22569 6208
rect 22603 6205 22615 6239
rect 23934 6236 23940 6248
rect 23895 6208 23940 6236
rect 22557 6199 22615 6205
rect 19076 6140 19564 6168
rect 22204 6168 22232 6199
rect 23934 6196 23940 6208
rect 23992 6196 23998 6248
rect 24026 6196 24032 6248
rect 24084 6236 24090 6248
rect 24670 6236 24676 6248
rect 24084 6208 24129 6236
rect 24631 6208 24676 6236
rect 24084 6196 24090 6208
rect 24670 6196 24676 6208
rect 24728 6196 24734 6248
rect 25884 6245 25912 6276
rect 26418 6264 26424 6276
rect 26476 6304 26482 6316
rect 26970 6304 26976 6316
rect 26476 6276 26976 6304
rect 26476 6264 26482 6276
rect 26970 6264 26976 6276
rect 27028 6264 27034 6316
rect 27890 6264 27896 6316
rect 27948 6304 27954 6316
rect 30098 6304 30104 6316
rect 27948 6276 30104 6304
rect 27948 6264 27954 6276
rect 30098 6264 30104 6276
rect 30156 6264 30162 6316
rect 30926 6264 30932 6316
rect 30984 6304 30990 6316
rect 31021 6307 31079 6313
rect 31021 6304 31033 6307
rect 30984 6276 31033 6304
rect 30984 6264 30990 6276
rect 31021 6273 31033 6276
rect 31067 6273 31079 6307
rect 31478 6304 31484 6316
rect 31439 6276 31484 6304
rect 31021 6267 31079 6273
rect 31478 6264 31484 6276
rect 31536 6264 31542 6316
rect 32217 6307 32275 6313
rect 32217 6273 32229 6307
rect 32263 6304 32275 6307
rect 32398 6304 32404 6316
rect 32263 6276 32404 6304
rect 32263 6273 32275 6276
rect 32217 6267 32275 6273
rect 32398 6264 32404 6276
rect 32456 6264 32462 6316
rect 32766 6304 32772 6316
rect 32727 6276 32772 6304
rect 32766 6264 32772 6276
rect 32824 6264 32830 6316
rect 36078 6304 36084 6316
rect 33060 6276 36084 6304
rect 25869 6239 25927 6245
rect 25869 6205 25881 6239
rect 25915 6205 25927 6239
rect 25869 6199 25927 6205
rect 26605 6239 26663 6245
rect 26605 6205 26617 6239
rect 26651 6205 26663 6239
rect 26878 6236 26884 6248
rect 26839 6208 26884 6236
rect 26605 6199 26663 6205
rect 22462 6168 22468 6180
rect 22204 6140 22468 6168
rect 19076 6112 19104 6140
rect 22462 6128 22468 6140
rect 22520 6128 22526 6180
rect 8352 6072 14596 6100
rect 8352 6060 8358 6072
rect 17770 6060 17776 6112
rect 17828 6100 17834 6112
rect 18417 6103 18475 6109
rect 18417 6100 18429 6103
rect 17828 6072 18429 6100
rect 17828 6060 17834 6072
rect 18417 6069 18429 6072
rect 18463 6069 18475 6103
rect 19058 6100 19064 6112
rect 19019 6072 19064 6100
rect 18417 6063 18475 6069
rect 19058 6060 19064 6072
rect 19116 6060 19122 6112
rect 26620 6100 26648 6199
rect 26878 6196 26884 6208
rect 26936 6196 26942 6248
rect 29270 6236 29276 6248
rect 29231 6208 29276 6236
rect 29270 6196 29276 6208
rect 29328 6196 29334 6248
rect 31297 6239 31355 6245
rect 31297 6205 31309 6239
rect 31343 6236 31355 6239
rect 31938 6236 31944 6248
rect 31343 6208 31944 6236
rect 31343 6205 31355 6208
rect 31297 6199 31355 6205
rect 31938 6196 31944 6208
rect 31996 6196 32002 6248
rect 33060 6245 33088 6276
rect 36078 6264 36084 6276
rect 36136 6304 36142 6316
rect 36265 6307 36323 6313
rect 36265 6304 36277 6307
rect 36136 6276 36277 6304
rect 36136 6264 36142 6276
rect 36265 6273 36277 6276
rect 36311 6273 36323 6307
rect 36265 6267 36323 6273
rect 33045 6239 33103 6245
rect 33045 6205 33057 6239
rect 33091 6205 33103 6239
rect 33045 6199 33103 6205
rect 33229 6239 33287 6245
rect 33229 6205 33241 6239
rect 33275 6205 33287 6239
rect 33229 6199 33287 6205
rect 30469 6171 30527 6177
rect 30469 6137 30481 6171
rect 30515 6168 30527 6171
rect 30926 6168 30932 6180
rect 30515 6140 30932 6168
rect 30515 6137 30527 6140
rect 30469 6131 30527 6137
rect 30926 6128 30932 6140
rect 30984 6128 30990 6180
rect 31754 6128 31760 6180
rect 31812 6168 31818 6180
rect 33244 6168 33272 6199
rect 33594 6196 33600 6248
rect 33652 6236 33658 6248
rect 33689 6239 33747 6245
rect 33689 6236 33701 6239
rect 33652 6208 33701 6236
rect 33652 6196 33658 6208
rect 33689 6205 33701 6208
rect 33735 6205 33747 6239
rect 34885 6239 34943 6245
rect 34885 6236 34897 6239
rect 33689 6199 33747 6205
rect 34808 6208 34897 6236
rect 33781 6171 33839 6177
rect 33781 6168 33793 6171
rect 31812 6140 33793 6168
rect 31812 6128 31818 6140
rect 33781 6137 33793 6140
rect 33827 6137 33839 6171
rect 33781 6131 33839 6137
rect 29086 6100 29092 6112
rect 26620 6072 29092 6100
rect 29086 6060 29092 6072
rect 29144 6060 29150 6112
rect 33502 6060 33508 6112
rect 33560 6100 33566 6112
rect 34422 6100 34428 6112
rect 33560 6072 34428 6100
rect 33560 6060 33566 6072
rect 34422 6060 34428 6072
rect 34480 6100 34486 6112
rect 34808 6100 34836 6208
rect 34885 6205 34897 6208
rect 34931 6205 34943 6239
rect 34885 6199 34943 6205
rect 35161 6239 35219 6245
rect 35161 6205 35173 6239
rect 35207 6236 35219 6239
rect 37001 6239 37059 6245
rect 37001 6236 37013 6239
rect 35207 6208 37013 6236
rect 35207 6205 35219 6208
rect 35161 6199 35219 6205
rect 37001 6205 37013 6208
rect 37047 6205 37059 6239
rect 37001 6199 37059 6205
rect 37090 6196 37096 6248
rect 37148 6236 37154 6248
rect 37844 6245 37872 6344
rect 37553 6239 37611 6245
rect 37553 6236 37565 6239
rect 37148 6208 37565 6236
rect 37148 6196 37154 6208
rect 37553 6205 37565 6208
rect 37599 6205 37611 6239
rect 37553 6199 37611 6205
rect 37829 6239 37887 6245
rect 37829 6205 37841 6239
rect 37875 6205 37887 6239
rect 37829 6199 37887 6205
rect 38013 6239 38071 6245
rect 38013 6205 38025 6239
rect 38059 6205 38071 6239
rect 38013 6199 38071 6205
rect 36722 6128 36728 6180
rect 36780 6168 36786 6180
rect 38028 6168 38056 6199
rect 36780 6140 38056 6168
rect 36780 6128 36786 6140
rect 34480 6072 34836 6100
rect 34480 6060 34486 6072
rect 1104 6010 39836 6032
rect 1104 5958 19606 6010
rect 19658 5958 19670 6010
rect 19722 5958 19734 6010
rect 19786 5958 19798 6010
rect 19850 5958 39836 6010
rect 1104 5936 39836 5958
rect 5534 5856 5540 5908
rect 5592 5896 5598 5908
rect 11514 5896 11520 5908
rect 5592 5868 11520 5896
rect 5592 5856 5598 5868
rect 11514 5856 11520 5868
rect 11572 5856 11578 5908
rect 12158 5856 12164 5908
rect 12216 5896 12222 5908
rect 12805 5899 12863 5905
rect 12805 5896 12817 5899
rect 12216 5868 12817 5896
rect 12216 5856 12222 5868
rect 12805 5865 12817 5868
rect 12851 5865 12863 5899
rect 13814 5896 13820 5908
rect 12805 5859 12863 5865
rect 13280 5868 13820 5896
rect 6733 5831 6791 5837
rect 6733 5797 6745 5831
rect 6779 5828 6791 5831
rect 8202 5828 8208 5840
rect 6779 5800 8208 5828
rect 6779 5797 6791 5800
rect 6733 5791 6791 5797
rect 8202 5788 8208 5800
rect 8260 5788 8266 5840
rect 8386 5788 8392 5840
rect 8444 5828 8450 5840
rect 8444 5800 10364 5828
rect 8444 5788 8450 5800
rect 4338 5760 4344 5772
rect 4299 5732 4344 5760
rect 4338 5720 4344 5732
rect 4396 5720 4402 5772
rect 6273 5763 6331 5769
rect 6273 5729 6285 5763
rect 6319 5760 6331 5763
rect 6914 5760 6920 5772
rect 6319 5732 6920 5760
rect 6319 5729 6331 5732
rect 6273 5723 6331 5729
rect 6914 5720 6920 5732
rect 6972 5720 6978 5772
rect 7098 5720 7104 5772
rect 7156 5760 7162 5772
rect 7193 5763 7251 5769
rect 7193 5760 7205 5763
rect 7156 5732 7205 5760
rect 7156 5720 7162 5732
rect 7193 5729 7205 5732
rect 7239 5729 7251 5763
rect 7193 5723 7251 5729
rect 7837 5763 7895 5769
rect 7837 5729 7849 5763
rect 7883 5729 7895 5763
rect 8110 5760 8116 5772
rect 8071 5732 8116 5760
rect 7837 5723 7895 5729
rect 4062 5692 4068 5704
rect 4023 5664 4068 5692
rect 4062 5652 4068 5664
rect 4120 5652 4126 5704
rect 6181 5695 6239 5701
rect 6181 5661 6193 5695
rect 6227 5692 6239 5695
rect 6546 5692 6552 5704
rect 6227 5664 6552 5692
rect 6227 5661 6239 5664
rect 6181 5655 6239 5661
rect 6546 5652 6552 5664
rect 6604 5652 6610 5704
rect 7852 5692 7880 5723
rect 8110 5720 8116 5732
rect 8168 5720 8174 5772
rect 8573 5763 8631 5769
rect 8573 5729 8585 5763
rect 8619 5760 8631 5763
rect 8754 5760 8760 5772
rect 8619 5732 8760 5760
rect 8619 5729 8631 5732
rect 8573 5723 8631 5729
rect 8754 5720 8760 5732
rect 8812 5720 8818 5772
rect 9125 5763 9183 5769
rect 9125 5729 9137 5763
rect 9171 5760 9183 5763
rect 9582 5760 9588 5772
rect 9171 5732 9588 5760
rect 9171 5729 9183 5732
rect 9125 5723 9183 5729
rect 9582 5720 9588 5732
rect 9640 5720 9646 5772
rect 9677 5763 9735 5769
rect 9677 5729 9689 5763
rect 9723 5760 9735 5763
rect 9766 5760 9772 5772
rect 9723 5732 9772 5760
rect 9723 5729 9735 5732
rect 9677 5723 9735 5729
rect 9766 5720 9772 5732
rect 9824 5720 9830 5772
rect 10336 5769 10364 5800
rect 10321 5763 10379 5769
rect 10321 5729 10333 5763
rect 10367 5729 10379 5763
rect 10321 5723 10379 5729
rect 10965 5763 11023 5769
rect 10965 5729 10977 5763
rect 11011 5760 11023 5763
rect 11054 5760 11060 5772
rect 11011 5732 11060 5760
rect 11011 5729 11023 5732
rect 10965 5723 11023 5729
rect 7852 5664 9812 5692
rect 5629 5627 5687 5633
rect 5629 5593 5641 5627
rect 5675 5624 5687 5627
rect 7006 5624 7012 5636
rect 5675 5596 7012 5624
rect 5675 5593 5687 5596
rect 5629 5587 5687 5593
rect 7006 5584 7012 5596
rect 7064 5584 7070 5636
rect 7282 5624 7288 5636
rect 7243 5596 7288 5624
rect 7282 5584 7288 5596
rect 7340 5584 7346 5636
rect 9784 5565 9812 5664
rect 9769 5559 9827 5565
rect 9769 5525 9781 5559
rect 9815 5556 9827 5559
rect 10134 5556 10140 5568
rect 9815 5528 10140 5556
rect 9815 5525 9827 5528
rect 9769 5519 9827 5525
rect 10134 5516 10140 5528
rect 10192 5516 10198 5568
rect 10336 5556 10364 5723
rect 11054 5720 11060 5732
rect 11112 5720 11118 5772
rect 11333 5763 11391 5769
rect 11333 5729 11345 5763
rect 11379 5729 11391 5763
rect 11514 5760 11520 5772
rect 11475 5732 11520 5760
rect 11333 5723 11391 5729
rect 10502 5692 10508 5704
rect 10463 5664 10508 5692
rect 10502 5652 10508 5664
rect 10560 5652 10566 5704
rect 10410 5584 10416 5636
rect 10468 5624 10474 5636
rect 11348 5624 11376 5723
rect 11514 5720 11520 5732
rect 11572 5720 11578 5772
rect 12250 5760 12256 5772
rect 12211 5732 12256 5760
rect 12250 5720 12256 5732
rect 12308 5720 12314 5772
rect 12897 5763 12955 5769
rect 12897 5729 12909 5763
rect 12943 5760 12955 5763
rect 13280 5760 13308 5868
rect 13814 5856 13820 5868
rect 13872 5856 13878 5908
rect 14274 5896 14280 5908
rect 14235 5868 14280 5896
rect 14274 5856 14280 5868
rect 14332 5856 14338 5908
rect 16114 5896 16120 5908
rect 14384 5868 16120 5896
rect 13722 5828 13728 5840
rect 13372 5800 13728 5828
rect 13372 5769 13400 5800
rect 13722 5788 13728 5800
rect 13780 5788 13786 5840
rect 12943 5732 13308 5760
rect 13357 5763 13415 5769
rect 12943 5729 12955 5732
rect 12897 5723 12955 5729
rect 13357 5729 13369 5763
rect 13403 5729 13415 5763
rect 13538 5760 13544 5772
rect 13499 5732 13544 5760
rect 13357 5723 13415 5729
rect 13538 5720 13544 5732
rect 13596 5720 13602 5772
rect 13814 5720 13820 5772
rect 13872 5760 13878 5772
rect 14384 5760 14412 5868
rect 16114 5856 16120 5868
rect 16172 5856 16178 5908
rect 17586 5856 17592 5908
rect 17644 5896 17650 5908
rect 19061 5899 19119 5905
rect 19061 5896 19073 5899
rect 17644 5868 19073 5896
rect 17644 5856 17650 5868
rect 19061 5865 19073 5868
rect 19107 5865 19119 5899
rect 19061 5859 19119 5865
rect 20254 5856 20260 5908
rect 20312 5896 20318 5908
rect 20993 5899 21051 5905
rect 20993 5896 21005 5899
rect 20312 5868 21005 5896
rect 20312 5856 20318 5868
rect 20993 5865 21005 5868
rect 21039 5865 21051 5899
rect 20993 5859 21051 5865
rect 21634 5856 21640 5908
rect 21692 5896 21698 5908
rect 23201 5899 23259 5905
rect 23201 5896 23213 5899
rect 21692 5868 23213 5896
rect 21692 5856 21698 5868
rect 23201 5865 23213 5868
rect 23247 5865 23259 5899
rect 23201 5859 23259 5865
rect 25866 5856 25872 5908
rect 25924 5896 25930 5908
rect 25924 5868 28028 5896
rect 25924 5856 25930 5868
rect 17770 5828 17776 5840
rect 15120 5800 17776 5828
rect 13872 5732 14412 5760
rect 14461 5763 14519 5769
rect 13872 5720 13878 5732
rect 14461 5729 14473 5763
rect 14507 5760 14519 5763
rect 14550 5760 14556 5772
rect 14507 5732 14556 5760
rect 14507 5729 14519 5732
rect 14461 5723 14519 5729
rect 14550 5720 14556 5732
rect 14608 5720 14614 5772
rect 15120 5769 15148 5800
rect 17770 5788 17776 5800
rect 17828 5788 17834 5840
rect 20916 5800 21956 5828
rect 15105 5763 15163 5769
rect 15105 5729 15117 5763
rect 15151 5729 15163 5763
rect 15105 5723 15163 5729
rect 15194 5720 15200 5772
rect 15252 5760 15258 5772
rect 15289 5763 15347 5769
rect 15289 5760 15301 5763
rect 15252 5732 15301 5760
rect 15252 5720 15258 5732
rect 15289 5729 15301 5732
rect 15335 5729 15347 5763
rect 15930 5760 15936 5772
rect 15891 5732 15936 5760
rect 15289 5723 15347 5729
rect 15930 5720 15936 5732
rect 15988 5720 15994 5772
rect 16022 5720 16028 5772
rect 16080 5760 16086 5772
rect 16485 5763 16543 5769
rect 16080 5732 16125 5760
rect 16080 5720 16086 5732
rect 16485 5729 16497 5763
rect 16531 5729 16543 5763
rect 16485 5723 16543 5729
rect 13630 5624 13636 5636
rect 10468 5596 13636 5624
rect 10468 5584 10474 5596
rect 13630 5584 13636 5596
rect 13688 5584 13694 5636
rect 14734 5584 14740 5636
rect 14792 5624 14798 5636
rect 15381 5627 15439 5633
rect 15381 5624 15393 5627
rect 14792 5596 15393 5624
rect 14792 5584 14798 5596
rect 15381 5593 15393 5596
rect 15427 5593 15439 5627
rect 16500 5624 16528 5723
rect 16574 5720 16580 5772
rect 16632 5760 16638 5772
rect 17221 5763 17279 5769
rect 17221 5760 17233 5763
rect 16632 5732 17233 5760
rect 16632 5720 16638 5732
rect 17221 5729 17233 5732
rect 17267 5760 17279 5763
rect 17954 5760 17960 5772
rect 17267 5732 17816 5760
rect 17915 5732 17960 5760
rect 17267 5729 17279 5732
rect 17221 5723 17279 5729
rect 17681 5695 17739 5701
rect 17681 5661 17693 5695
rect 17727 5661 17739 5695
rect 17788 5692 17816 5732
rect 17954 5720 17960 5732
rect 18012 5720 18018 5772
rect 20916 5769 20944 5800
rect 20901 5763 20959 5769
rect 20901 5729 20913 5763
rect 20947 5729 20959 5763
rect 21726 5760 21732 5772
rect 21687 5732 21732 5760
rect 20901 5723 20959 5729
rect 21726 5720 21732 5732
rect 21784 5720 21790 5772
rect 21634 5692 21640 5704
rect 17788 5664 21640 5692
rect 17681 5655 17739 5661
rect 16942 5624 16948 5636
rect 16500 5596 16948 5624
rect 15381 5587 15439 5593
rect 16942 5584 16948 5596
rect 17000 5584 17006 5636
rect 12802 5556 12808 5568
rect 10336 5528 12808 5556
rect 12802 5516 12808 5528
rect 12860 5556 12866 5568
rect 13446 5556 13452 5568
rect 12860 5528 13452 5556
rect 12860 5516 12866 5528
rect 13446 5516 13452 5528
rect 13504 5516 13510 5568
rect 13538 5516 13544 5568
rect 13596 5556 13602 5568
rect 14921 5559 14979 5565
rect 14921 5556 14933 5559
rect 13596 5528 14933 5556
rect 13596 5516 13602 5528
rect 14921 5525 14933 5528
rect 14967 5525 14979 5559
rect 14921 5519 14979 5525
rect 15930 5516 15936 5568
rect 15988 5556 15994 5568
rect 17586 5556 17592 5568
rect 15988 5528 17592 5556
rect 15988 5516 15994 5528
rect 17586 5516 17592 5528
rect 17644 5516 17650 5568
rect 17696 5556 17724 5655
rect 21634 5652 21640 5664
rect 21692 5652 21698 5704
rect 21818 5692 21824 5704
rect 21731 5664 21824 5692
rect 21744 5624 21772 5664
rect 21818 5652 21824 5664
rect 21876 5652 21882 5704
rect 21928 5692 21956 5800
rect 26878 5788 26884 5840
rect 26936 5828 26942 5840
rect 27065 5831 27123 5837
rect 27065 5828 27077 5831
rect 26936 5800 27077 5828
rect 26936 5788 26942 5800
rect 27065 5797 27077 5800
rect 27111 5797 27123 5831
rect 27065 5791 27123 5797
rect 22097 5763 22155 5769
rect 22097 5729 22109 5763
rect 22143 5760 22155 5763
rect 22370 5760 22376 5772
rect 22143 5732 22376 5760
rect 22143 5729 22155 5732
rect 22097 5723 22155 5729
rect 22370 5720 22376 5732
rect 22428 5720 22434 5772
rect 23937 5763 23995 5769
rect 23937 5729 23949 5763
rect 23983 5760 23995 5763
rect 24210 5760 24216 5772
rect 23983 5732 24216 5760
rect 23983 5729 23995 5732
rect 23937 5723 23995 5729
rect 24210 5720 24216 5732
rect 24268 5720 24274 5772
rect 24949 5763 25007 5769
rect 24949 5729 24961 5763
rect 24995 5729 25007 5763
rect 25130 5760 25136 5772
rect 25091 5732 25136 5760
rect 24949 5723 25007 5729
rect 24118 5692 24124 5704
rect 21928 5664 24124 5692
rect 24118 5652 24124 5664
rect 24176 5652 24182 5704
rect 24854 5624 24860 5636
rect 19076 5596 21772 5624
rect 24815 5596 24860 5624
rect 19076 5568 19104 5596
rect 24854 5584 24860 5596
rect 24912 5584 24918 5636
rect 17954 5556 17960 5568
rect 17696 5528 17960 5556
rect 17954 5516 17960 5528
rect 18012 5556 18018 5568
rect 19058 5556 19064 5568
rect 18012 5528 19064 5556
rect 18012 5516 18018 5528
rect 19058 5516 19064 5528
rect 19116 5516 19122 5568
rect 19978 5516 19984 5568
rect 20036 5556 20042 5568
rect 21545 5559 21603 5565
rect 21545 5556 21557 5559
rect 20036 5528 21557 5556
rect 20036 5516 20042 5528
rect 21545 5525 21557 5528
rect 21591 5525 21603 5559
rect 21545 5519 21603 5525
rect 21634 5516 21640 5568
rect 21692 5556 21698 5568
rect 24029 5559 24087 5565
rect 24029 5556 24041 5559
rect 21692 5528 24041 5556
rect 21692 5516 21698 5528
rect 24029 5525 24041 5528
rect 24075 5525 24087 5559
rect 24964 5556 24992 5723
rect 25130 5720 25136 5732
rect 25188 5720 25194 5772
rect 25777 5763 25835 5769
rect 25777 5729 25789 5763
rect 25823 5760 25835 5763
rect 26326 5760 26332 5772
rect 25823 5732 26332 5760
rect 25823 5729 25835 5732
rect 25777 5723 25835 5729
rect 26326 5720 26332 5732
rect 26384 5720 26390 5772
rect 27614 5760 27620 5772
rect 27575 5732 27620 5760
rect 27614 5720 27620 5732
rect 27672 5720 27678 5772
rect 27890 5760 27896 5772
rect 27851 5732 27896 5760
rect 27890 5720 27896 5732
rect 27948 5720 27954 5772
rect 28000 5760 28028 5868
rect 28166 5856 28172 5908
rect 28224 5896 28230 5908
rect 28721 5899 28779 5905
rect 28721 5896 28733 5899
rect 28224 5868 28733 5896
rect 28224 5856 28230 5868
rect 28721 5865 28733 5868
rect 28767 5896 28779 5899
rect 29914 5896 29920 5908
rect 28767 5868 29920 5896
rect 28767 5865 28779 5868
rect 28721 5859 28779 5865
rect 29914 5856 29920 5868
rect 29972 5856 29978 5908
rect 31018 5856 31024 5908
rect 31076 5896 31082 5908
rect 31481 5899 31539 5905
rect 31481 5896 31493 5899
rect 31076 5868 31493 5896
rect 31076 5856 31082 5868
rect 31481 5865 31493 5868
rect 31527 5865 31539 5899
rect 35342 5896 35348 5908
rect 31481 5859 31539 5865
rect 34624 5868 35348 5896
rect 28626 5788 28632 5840
rect 28684 5828 28690 5840
rect 34624 5828 34652 5868
rect 35342 5856 35348 5868
rect 35400 5896 35406 5908
rect 36722 5896 36728 5908
rect 35400 5868 36728 5896
rect 35400 5856 35406 5868
rect 36722 5856 36728 5868
rect 36780 5856 36786 5908
rect 28684 5800 30420 5828
rect 28684 5788 28690 5800
rect 28537 5763 28595 5769
rect 28537 5760 28549 5763
rect 28000 5732 28549 5760
rect 28537 5729 28549 5732
rect 28583 5760 28595 5763
rect 29270 5760 29276 5772
rect 28583 5732 29276 5760
rect 28583 5729 28595 5732
rect 28537 5723 28595 5729
rect 29270 5720 29276 5732
rect 29328 5720 29334 5772
rect 29914 5760 29920 5772
rect 29875 5732 29920 5760
rect 29914 5720 29920 5732
rect 29972 5720 29978 5772
rect 30098 5720 30104 5772
rect 30156 5760 30162 5772
rect 30392 5769 30420 5800
rect 34532 5800 34652 5828
rect 34532 5772 34560 5800
rect 34790 5788 34796 5840
rect 34848 5828 34854 5840
rect 35161 5831 35219 5837
rect 35161 5828 35173 5831
rect 34848 5800 35173 5828
rect 34848 5788 34854 5800
rect 35161 5797 35173 5800
rect 35207 5797 35219 5831
rect 35161 5791 35219 5797
rect 30193 5763 30251 5769
rect 30193 5760 30205 5763
rect 30156 5732 30205 5760
rect 30156 5720 30162 5732
rect 30193 5729 30205 5732
rect 30239 5729 30251 5763
rect 30193 5723 30251 5729
rect 30377 5763 30435 5769
rect 30377 5729 30389 5763
rect 30423 5729 30435 5763
rect 30377 5723 30435 5729
rect 31297 5763 31355 5769
rect 31297 5729 31309 5763
rect 31343 5760 31355 5763
rect 31754 5760 31760 5772
rect 31343 5732 31760 5760
rect 31343 5729 31355 5732
rect 31297 5723 31355 5729
rect 31754 5720 31760 5732
rect 31812 5720 31818 5772
rect 32674 5760 32680 5772
rect 32635 5732 32680 5760
rect 32674 5720 32680 5732
rect 32732 5720 32738 5772
rect 32953 5763 33011 5769
rect 32953 5729 32965 5763
rect 32999 5760 33011 5763
rect 33226 5760 33232 5772
rect 32999 5732 33232 5760
rect 32999 5729 33011 5732
rect 32953 5723 33011 5729
rect 28077 5695 28135 5701
rect 28077 5661 28089 5695
rect 28123 5661 28135 5695
rect 29362 5692 29368 5704
rect 29323 5664 29368 5692
rect 28077 5655 28135 5661
rect 28092 5624 28120 5655
rect 29362 5652 29368 5664
rect 29420 5652 29426 5704
rect 32125 5695 32183 5701
rect 32125 5661 32137 5695
rect 32171 5692 32183 5695
rect 32582 5692 32588 5704
rect 32171 5664 32588 5692
rect 32171 5661 32183 5664
rect 32125 5655 32183 5661
rect 32582 5652 32588 5664
rect 32640 5652 32646 5704
rect 28994 5624 29000 5636
rect 28092 5596 29000 5624
rect 28994 5584 29000 5596
rect 29052 5584 29058 5636
rect 28902 5556 28908 5568
rect 24964 5528 28908 5556
rect 24029 5519 24087 5525
rect 28902 5516 28908 5528
rect 28960 5556 28966 5568
rect 32968 5556 32996 5723
rect 33226 5720 33232 5732
rect 33284 5720 33290 5772
rect 33594 5760 33600 5772
rect 33520 5732 33600 5760
rect 33137 5695 33195 5701
rect 33137 5661 33149 5695
rect 33183 5692 33195 5695
rect 33520 5692 33548 5732
rect 33594 5720 33600 5732
rect 33652 5720 33658 5772
rect 34514 5760 34520 5772
rect 34427 5732 34520 5760
rect 34514 5720 34520 5732
rect 34572 5720 34578 5772
rect 34698 5760 34704 5772
rect 34659 5732 34704 5760
rect 34698 5720 34704 5732
rect 34756 5720 34762 5772
rect 34882 5720 34888 5772
rect 34940 5760 34946 5772
rect 35618 5760 35624 5772
rect 34940 5732 35624 5760
rect 34940 5720 34946 5732
rect 35618 5720 35624 5732
rect 35676 5760 35682 5772
rect 35713 5763 35771 5769
rect 35713 5760 35725 5763
rect 35676 5732 35725 5760
rect 35676 5720 35682 5732
rect 35713 5729 35725 5732
rect 35759 5729 35771 5763
rect 35713 5723 35771 5729
rect 35989 5763 36047 5769
rect 35989 5729 36001 5763
rect 36035 5760 36047 5763
rect 36538 5760 36544 5772
rect 36035 5732 36544 5760
rect 36035 5729 36047 5732
rect 35989 5723 36047 5729
rect 36538 5720 36544 5732
rect 36596 5760 36602 5772
rect 36906 5760 36912 5772
rect 36596 5732 36912 5760
rect 36596 5720 36602 5732
rect 36906 5720 36912 5732
rect 36964 5720 36970 5772
rect 33686 5692 33692 5704
rect 33183 5664 33548 5692
rect 33647 5664 33692 5692
rect 33183 5661 33195 5664
rect 33137 5655 33195 5661
rect 33686 5652 33692 5664
rect 33744 5652 33750 5704
rect 34241 5695 34299 5701
rect 34241 5661 34253 5695
rect 34287 5692 34299 5695
rect 34606 5692 34612 5704
rect 34287 5664 34612 5692
rect 34287 5661 34299 5664
rect 34241 5655 34299 5661
rect 34606 5652 34612 5664
rect 34664 5652 34670 5704
rect 34716 5692 34744 5720
rect 36173 5695 36231 5701
rect 36173 5692 36185 5695
rect 34716 5664 36185 5692
rect 36173 5661 36185 5664
rect 36219 5661 36231 5695
rect 36173 5655 36231 5661
rect 28960 5528 32996 5556
rect 28960 5516 28966 5528
rect 1104 5466 39836 5488
rect 1104 5414 4246 5466
rect 4298 5414 4310 5466
rect 4362 5414 4374 5466
rect 4426 5414 4438 5466
rect 4490 5414 34966 5466
rect 35018 5414 35030 5466
rect 35082 5414 35094 5466
rect 35146 5414 35158 5466
rect 35210 5414 39836 5466
rect 1104 5392 39836 5414
rect 5997 5355 6055 5361
rect 5997 5321 6009 5355
rect 6043 5352 6055 5355
rect 6086 5352 6092 5364
rect 6043 5324 6092 5352
rect 6043 5321 6055 5324
rect 5997 5315 6055 5321
rect 6086 5312 6092 5324
rect 6144 5312 6150 5364
rect 8573 5355 8631 5361
rect 8573 5321 8585 5355
rect 8619 5352 8631 5355
rect 9766 5352 9772 5364
rect 8619 5324 9772 5352
rect 8619 5321 8631 5324
rect 8573 5315 8631 5321
rect 9766 5312 9772 5324
rect 9824 5312 9830 5364
rect 11054 5312 11060 5364
rect 11112 5352 11118 5364
rect 11514 5352 11520 5364
rect 11112 5324 11520 5352
rect 11112 5312 11118 5324
rect 11514 5312 11520 5324
rect 11572 5352 11578 5364
rect 11609 5355 11667 5361
rect 11609 5352 11621 5355
rect 11572 5324 11621 5352
rect 11572 5312 11578 5324
rect 11609 5321 11621 5324
rect 11655 5321 11667 5355
rect 11609 5315 11667 5321
rect 13446 5312 13452 5364
rect 13504 5352 13510 5364
rect 13722 5352 13728 5364
rect 13504 5324 13728 5352
rect 13504 5312 13510 5324
rect 13722 5312 13728 5324
rect 13780 5312 13786 5364
rect 17586 5312 17592 5364
rect 17644 5352 17650 5364
rect 18141 5355 18199 5361
rect 18141 5352 18153 5355
rect 17644 5324 18153 5352
rect 17644 5312 17650 5324
rect 18141 5321 18153 5324
rect 18187 5321 18199 5355
rect 26418 5352 26424 5364
rect 26379 5324 26424 5352
rect 18141 5315 18199 5321
rect 12250 5244 12256 5296
rect 12308 5284 12314 5296
rect 16390 5284 16396 5296
rect 12308 5256 16396 5284
rect 12308 5244 12314 5256
rect 4062 5176 4068 5228
rect 4120 5216 4126 5228
rect 4617 5219 4675 5225
rect 4617 5216 4629 5219
rect 4120 5188 4629 5216
rect 4120 5176 4126 5188
rect 4617 5185 4629 5188
rect 4663 5185 4675 5219
rect 4890 5216 4896 5228
rect 4851 5188 4896 5216
rect 4617 5179 4675 5185
rect 2314 5108 2320 5160
rect 2372 5148 2378 5160
rect 3329 5151 3387 5157
rect 3329 5148 3341 5151
rect 2372 5120 3341 5148
rect 2372 5108 2378 5120
rect 3329 5117 3341 5120
rect 3375 5117 3387 5151
rect 3329 5111 3387 5117
rect 3881 5151 3939 5157
rect 3881 5117 3893 5151
rect 3927 5148 3939 5151
rect 4522 5148 4528 5160
rect 3927 5120 4528 5148
rect 3927 5117 3939 5120
rect 3881 5111 3939 5117
rect 4522 5108 4528 5120
rect 4580 5108 4586 5160
rect 4632 5148 4660 5179
rect 4890 5176 4896 5188
rect 4948 5176 4954 5228
rect 7282 5216 7288 5228
rect 7243 5188 7288 5216
rect 7282 5176 7288 5188
rect 7340 5176 7346 5228
rect 8478 5176 8484 5228
rect 8536 5216 8542 5228
rect 9217 5219 9275 5225
rect 9217 5216 9229 5219
rect 8536 5188 9229 5216
rect 8536 5176 8542 5188
rect 9217 5185 9229 5188
rect 9263 5185 9275 5219
rect 9217 5179 9275 5185
rect 9858 5176 9864 5228
rect 9916 5216 9922 5228
rect 10410 5216 10416 5228
rect 9916 5188 10416 5216
rect 9916 5176 9922 5188
rect 6822 5148 6828 5160
rect 4632 5120 6828 5148
rect 6822 5108 6828 5120
rect 6880 5148 6886 5160
rect 7009 5151 7067 5157
rect 7009 5148 7021 5151
rect 6880 5120 7021 5148
rect 6880 5108 6886 5120
rect 7009 5117 7021 5120
rect 7055 5148 7067 5151
rect 8110 5148 8116 5160
rect 7055 5120 8116 5148
rect 7055 5117 7067 5120
rect 7009 5111 7067 5117
rect 8110 5108 8116 5120
rect 8168 5108 8174 5160
rect 8386 5108 8392 5160
rect 8444 5148 8450 5160
rect 9125 5151 9183 5157
rect 9125 5148 9137 5151
rect 8444 5120 9137 5148
rect 8444 5108 8450 5120
rect 9125 5117 9137 5120
rect 9171 5117 9183 5151
rect 9125 5111 9183 5117
rect 9674 5108 9680 5160
rect 9732 5148 9738 5160
rect 10152 5157 10180 5188
rect 10410 5176 10416 5188
rect 10468 5176 10474 5228
rect 10594 5176 10600 5228
rect 10652 5216 10658 5228
rect 12268 5216 12296 5244
rect 12710 5216 12716 5228
rect 10652 5188 12296 5216
rect 12671 5188 12716 5216
rect 10652 5176 10658 5188
rect 10137 5151 10195 5157
rect 9732 5120 9777 5148
rect 9732 5108 9738 5120
rect 10137 5117 10149 5151
rect 10183 5117 10195 5151
rect 10318 5148 10324 5160
rect 10279 5120 10324 5148
rect 10137 5111 10195 5117
rect 10318 5108 10324 5120
rect 10376 5108 10382 5160
rect 11072 5157 11100 5188
rect 12710 5176 12716 5188
rect 12768 5176 12774 5228
rect 11057 5151 11115 5157
rect 11057 5117 11069 5151
rect 11103 5117 11115 5151
rect 11057 5111 11115 5117
rect 11422 5108 11428 5160
rect 11480 5148 11486 5160
rect 11517 5151 11575 5157
rect 11517 5148 11529 5151
rect 11480 5120 11529 5148
rect 11480 5108 11486 5120
rect 11517 5117 11529 5120
rect 11563 5117 11575 5151
rect 12802 5148 12808 5160
rect 12763 5120 12808 5148
rect 11517 5111 11575 5117
rect 12802 5108 12808 5120
rect 12860 5108 12866 5160
rect 13265 5151 13323 5157
rect 13265 5117 13277 5151
rect 13311 5117 13323 5151
rect 13630 5148 13636 5160
rect 13591 5120 13636 5148
rect 13265 5111 13323 5117
rect 4062 5080 4068 5092
rect 4023 5052 4068 5080
rect 4062 5040 4068 5052
rect 4120 5040 4126 5092
rect 13280 5080 13308 5111
rect 13630 5108 13636 5120
rect 13688 5108 13694 5160
rect 13998 5148 14004 5160
rect 13959 5120 14004 5148
rect 13998 5108 14004 5120
rect 14056 5108 14062 5160
rect 14553 5151 14611 5157
rect 14553 5117 14565 5151
rect 14599 5148 14611 5151
rect 14660 5148 14688 5256
rect 16390 5244 16396 5256
rect 16448 5244 16454 5296
rect 16206 5216 16212 5228
rect 16167 5188 16212 5216
rect 16206 5176 16212 5188
rect 16264 5176 16270 5228
rect 16298 5176 16304 5228
rect 16356 5216 16362 5228
rect 18156 5216 18184 5315
rect 26418 5312 26424 5324
rect 26476 5312 26482 5364
rect 33137 5355 33195 5361
rect 33137 5321 33149 5355
rect 33183 5352 33195 5355
rect 33226 5352 33232 5364
rect 33183 5324 33232 5352
rect 33183 5321 33195 5324
rect 33137 5315 33195 5321
rect 33226 5312 33232 5324
rect 33284 5312 33290 5364
rect 36633 5355 36691 5361
rect 36633 5321 36645 5355
rect 36679 5352 36691 5355
rect 36722 5352 36728 5364
rect 36679 5324 36728 5352
rect 36679 5321 36691 5324
rect 36633 5315 36691 5321
rect 36722 5312 36728 5324
rect 36780 5312 36786 5364
rect 19429 5219 19487 5225
rect 16356 5188 18092 5216
rect 18156 5188 19196 5216
rect 16356 5176 16362 5188
rect 14599 5120 14688 5148
rect 14599 5117 14611 5120
rect 14553 5111 14611 5117
rect 15194 5108 15200 5160
rect 15252 5148 15258 5160
rect 15289 5151 15347 5157
rect 15289 5148 15301 5151
rect 15252 5120 15301 5148
rect 15252 5108 15258 5120
rect 15289 5117 15301 5120
rect 15335 5117 15347 5151
rect 15289 5111 15347 5117
rect 15654 5108 15660 5160
rect 15712 5148 15718 5160
rect 15749 5151 15807 5157
rect 15749 5148 15761 5151
rect 15712 5120 15761 5148
rect 15712 5108 15718 5120
rect 15749 5117 15761 5120
rect 15795 5117 15807 5151
rect 16022 5148 16028 5160
rect 15983 5120 16028 5148
rect 15749 5111 15807 5117
rect 13446 5080 13452 5092
rect 13280 5052 13452 5080
rect 13446 5040 13452 5052
rect 13504 5040 13510 5092
rect 15764 5080 15792 5111
rect 16022 5108 16028 5120
rect 16080 5108 16086 5160
rect 16669 5151 16727 5157
rect 16669 5117 16681 5151
rect 16715 5117 16727 5151
rect 16669 5111 16727 5117
rect 16482 5080 16488 5092
rect 15764 5052 16488 5080
rect 16482 5040 16488 5052
rect 16540 5040 16546 5092
rect 16684 5080 16712 5111
rect 16758 5108 16764 5160
rect 16816 5148 16822 5160
rect 16945 5151 17003 5157
rect 16945 5148 16957 5151
rect 16816 5120 16957 5148
rect 16816 5108 16822 5120
rect 16945 5117 16957 5120
rect 16991 5117 17003 5151
rect 16945 5111 17003 5117
rect 17770 5108 17776 5160
rect 17828 5148 17834 5160
rect 18064 5157 18092 5188
rect 17865 5151 17923 5157
rect 17865 5148 17877 5151
rect 17828 5120 17877 5148
rect 17828 5108 17834 5120
rect 17865 5117 17877 5120
rect 17911 5117 17923 5151
rect 17865 5111 17923 5117
rect 18049 5151 18107 5157
rect 18049 5117 18061 5151
rect 18095 5117 18107 5151
rect 18690 5148 18696 5160
rect 18651 5120 18696 5148
rect 18049 5111 18107 5117
rect 18690 5108 18696 5120
rect 18748 5108 18754 5160
rect 19168 5157 19196 5188
rect 19429 5185 19441 5219
rect 19475 5216 19487 5219
rect 20165 5219 20223 5225
rect 20165 5216 20177 5219
rect 19475 5188 20177 5216
rect 19475 5185 19487 5188
rect 19429 5179 19487 5185
rect 20165 5185 20177 5188
rect 20211 5185 20223 5219
rect 20165 5179 20223 5185
rect 21726 5176 21732 5228
rect 21784 5216 21790 5228
rect 22005 5219 22063 5225
rect 22005 5216 22017 5219
rect 21784 5188 22017 5216
rect 21784 5176 21790 5188
rect 22005 5185 22017 5188
rect 22051 5185 22063 5219
rect 28166 5216 28172 5228
rect 28127 5188 28172 5216
rect 22005 5179 22063 5185
rect 28166 5176 28172 5188
rect 28224 5176 28230 5228
rect 28626 5216 28632 5228
rect 28587 5188 28632 5216
rect 28626 5176 28632 5188
rect 28684 5176 28690 5228
rect 31573 5219 31631 5225
rect 31573 5216 31585 5219
rect 29288 5188 31585 5216
rect 19153 5151 19211 5157
rect 19153 5117 19165 5151
rect 19199 5117 19211 5151
rect 19153 5111 19211 5117
rect 19889 5151 19947 5157
rect 19889 5117 19901 5151
rect 19935 5117 19947 5151
rect 19889 5111 19947 5117
rect 16850 5080 16856 5092
rect 16684 5052 16856 5080
rect 16850 5040 16856 5052
rect 16908 5040 16914 5092
rect 17681 5015 17739 5021
rect 17681 4981 17693 5015
rect 17727 5012 17739 5015
rect 18046 5012 18052 5024
rect 17727 4984 18052 5012
rect 17727 4981 17739 4984
rect 17681 4975 17739 4981
rect 18046 4972 18052 4984
rect 18104 5012 18110 5024
rect 19904 5012 19932 5111
rect 22094 5108 22100 5160
rect 22152 5148 22158 5160
rect 22152 5120 22197 5148
rect 22152 5108 22158 5120
rect 23934 5108 23940 5160
rect 23992 5148 23998 5160
rect 24029 5151 24087 5157
rect 24029 5148 24041 5151
rect 23992 5120 24041 5148
rect 23992 5108 23998 5120
rect 24029 5117 24041 5120
rect 24075 5148 24087 5151
rect 24302 5148 24308 5160
rect 24075 5120 24308 5148
rect 24075 5117 24087 5120
rect 24029 5111 24087 5117
rect 24302 5108 24308 5120
rect 24360 5108 24366 5160
rect 24854 5148 24860 5160
rect 24815 5120 24860 5148
rect 24854 5108 24860 5120
rect 24912 5108 24918 5160
rect 25133 5151 25191 5157
rect 25133 5117 25145 5151
rect 25179 5148 25191 5151
rect 27522 5148 27528 5160
rect 25179 5120 27528 5148
rect 25179 5117 25191 5120
rect 25133 5111 25191 5117
rect 27522 5108 27528 5120
rect 27580 5108 27586 5160
rect 28258 5108 28264 5160
rect 28316 5148 28322 5160
rect 28445 5151 28503 5157
rect 28445 5148 28457 5151
rect 28316 5120 28457 5148
rect 28316 5108 28322 5120
rect 28445 5117 28457 5120
rect 28491 5117 28503 5151
rect 28445 5111 28503 5117
rect 29086 5108 29092 5160
rect 29144 5148 29150 5160
rect 29288 5157 29316 5188
rect 31573 5185 31585 5188
rect 31619 5185 31631 5219
rect 31573 5179 31631 5185
rect 35069 5219 35127 5225
rect 35069 5185 35081 5219
rect 35115 5216 35127 5219
rect 37090 5216 37096 5228
rect 35115 5188 37096 5216
rect 35115 5185 35127 5188
rect 35069 5179 35127 5185
rect 37090 5176 37096 5188
rect 37148 5176 37154 5228
rect 29273 5151 29331 5157
rect 29273 5148 29285 5151
rect 29144 5120 29285 5148
rect 29144 5108 29150 5120
rect 29273 5117 29285 5120
rect 29319 5117 29331 5151
rect 29546 5148 29552 5160
rect 29507 5120 29552 5148
rect 29273 5111 29331 5117
rect 29546 5108 29552 5120
rect 29604 5108 29610 5160
rect 31849 5151 31907 5157
rect 31849 5117 31861 5151
rect 31895 5148 31907 5151
rect 32122 5148 32128 5160
rect 31895 5120 32128 5148
rect 31895 5117 31907 5120
rect 31849 5111 31907 5117
rect 32122 5108 32128 5120
rect 32180 5108 32186 5160
rect 33965 5151 34023 5157
rect 33965 5117 33977 5151
rect 34011 5148 34023 5151
rect 34514 5148 34520 5160
rect 34011 5120 34520 5148
rect 34011 5117 34023 5120
rect 33965 5111 34023 5117
rect 34514 5108 34520 5120
rect 34572 5108 34578 5160
rect 35618 5148 35624 5160
rect 35579 5120 35624 5148
rect 35618 5108 35624 5120
rect 35676 5108 35682 5160
rect 35897 5151 35955 5157
rect 35897 5117 35909 5151
rect 35943 5117 35955 5151
rect 36078 5148 36084 5160
rect 36039 5120 36084 5148
rect 35897 5111 35955 5117
rect 21545 5083 21603 5089
rect 21545 5049 21557 5083
rect 21591 5080 21603 5083
rect 22186 5080 22192 5092
rect 21591 5052 22192 5080
rect 21591 5049 21603 5052
rect 21545 5043 21603 5049
rect 22186 5040 22192 5052
rect 22244 5040 22250 5092
rect 22557 5083 22615 5089
rect 22557 5049 22569 5083
rect 22603 5080 22615 5083
rect 22830 5080 22836 5092
rect 22603 5052 22836 5080
rect 22603 5049 22615 5052
rect 22557 5043 22615 5049
rect 22830 5040 22836 5052
rect 22888 5040 22894 5092
rect 27614 5080 27620 5092
rect 27575 5052 27620 5080
rect 27614 5040 27620 5052
rect 27672 5040 27678 5092
rect 24210 5012 24216 5024
rect 18104 4984 19932 5012
rect 24123 4984 24216 5012
rect 18104 4972 18110 4984
rect 24210 4972 24216 4984
rect 24268 5012 24274 5024
rect 28276 5012 28304 5108
rect 35912 5080 35940 5111
rect 36078 5108 36084 5120
rect 36136 5108 36142 5160
rect 36538 5148 36544 5160
rect 36499 5120 36544 5148
rect 36538 5108 36544 5120
rect 36596 5108 36602 5160
rect 35986 5080 35992 5092
rect 35899 5052 35992 5080
rect 35986 5040 35992 5052
rect 36044 5080 36050 5092
rect 36556 5080 36584 5108
rect 36044 5052 36584 5080
rect 36044 5040 36050 5052
rect 24268 4984 28304 5012
rect 24268 4972 24274 4984
rect 30006 4972 30012 5024
rect 30064 5012 30070 5024
rect 30653 5015 30711 5021
rect 30653 5012 30665 5015
rect 30064 4984 30665 5012
rect 30064 4972 30070 4984
rect 30653 4981 30665 4984
rect 30699 4981 30711 5015
rect 30653 4975 30711 4981
rect 34149 5015 34207 5021
rect 34149 4981 34161 5015
rect 34195 5012 34207 5015
rect 34422 5012 34428 5024
rect 34195 4984 34428 5012
rect 34195 4981 34207 4984
rect 34149 4975 34207 4981
rect 34422 4972 34428 4984
rect 34480 4972 34486 5024
rect 1104 4922 39836 4944
rect 1104 4870 19606 4922
rect 19658 4870 19670 4922
rect 19722 4870 19734 4922
rect 19786 4870 19798 4922
rect 19850 4870 39836 4922
rect 1104 4848 39836 4870
rect 2866 4768 2872 4820
rect 2924 4808 2930 4820
rect 5166 4808 5172 4820
rect 2924 4780 5172 4808
rect 2924 4768 2930 4780
rect 5166 4768 5172 4780
rect 5224 4808 5230 4820
rect 5261 4811 5319 4817
rect 5261 4808 5273 4811
rect 5224 4780 5273 4808
rect 5224 4768 5230 4780
rect 5261 4777 5273 4780
rect 5307 4777 5319 4811
rect 5261 4771 5319 4777
rect 6914 4768 6920 4820
rect 6972 4808 6978 4820
rect 7193 4811 7251 4817
rect 7193 4808 7205 4811
rect 6972 4780 7205 4808
rect 6972 4768 6978 4780
rect 7193 4777 7205 4780
rect 7239 4777 7251 4811
rect 8110 4808 8116 4820
rect 8071 4780 8116 4808
rect 7193 4771 7251 4777
rect 8110 4768 8116 4780
rect 8168 4768 8174 4820
rect 11238 4808 11244 4820
rect 8312 4780 11244 4808
rect 4798 4632 4804 4684
rect 4856 4672 4862 4684
rect 5077 4675 5135 4681
rect 5077 4672 5089 4675
rect 4856 4644 5089 4672
rect 4856 4632 4862 4644
rect 5077 4641 5089 4644
rect 5123 4672 5135 4675
rect 6362 4672 6368 4684
rect 5123 4644 6368 4672
rect 5123 4641 5135 4644
rect 5077 4635 5135 4641
rect 6362 4632 6368 4644
rect 6420 4632 6426 4684
rect 8312 4681 8340 4780
rect 11238 4768 11244 4780
rect 11296 4768 11302 4820
rect 11422 4768 11428 4820
rect 11480 4808 11486 4820
rect 11609 4811 11667 4817
rect 11609 4808 11621 4811
rect 11480 4780 11621 4808
rect 11480 4768 11486 4780
rect 11609 4777 11621 4780
rect 11655 4777 11667 4811
rect 11609 4771 11667 4777
rect 11790 4768 11796 4820
rect 11848 4808 11854 4820
rect 19058 4808 19064 4820
rect 11848 4780 19064 4808
rect 11848 4768 11854 4780
rect 8297 4675 8355 4681
rect 8297 4641 8309 4675
rect 8343 4641 8355 4675
rect 8662 4672 8668 4684
rect 8623 4644 8668 4672
rect 8297 4635 8355 4641
rect 8662 4632 8668 4644
rect 8720 4632 8726 4684
rect 8941 4675 8999 4681
rect 8941 4641 8953 4675
rect 8987 4672 8999 4675
rect 9674 4672 9680 4684
rect 8987 4644 9680 4672
rect 8987 4641 8999 4644
rect 8941 4635 8999 4641
rect 9674 4632 9680 4644
rect 9732 4672 9738 4684
rect 10318 4672 10324 4684
rect 9732 4644 10324 4672
rect 9732 4632 9738 4644
rect 10318 4632 10324 4644
rect 10376 4632 10382 4684
rect 10502 4672 10508 4684
rect 10463 4644 10508 4672
rect 10502 4632 10508 4644
rect 10560 4632 10566 4684
rect 12621 4675 12679 4681
rect 12621 4641 12633 4675
rect 12667 4672 12679 4675
rect 12710 4672 12716 4684
rect 12667 4644 12716 4672
rect 12667 4641 12679 4644
rect 12621 4635 12679 4641
rect 12710 4632 12716 4644
rect 12768 4632 12774 4684
rect 14001 4675 14059 4681
rect 14001 4641 14013 4675
rect 14047 4672 14059 4675
rect 14366 4672 14372 4684
rect 14047 4644 14372 4672
rect 14047 4641 14059 4644
rect 14001 4635 14059 4641
rect 14366 4632 14372 4644
rect 14424 4672 14430 4684
rect 14461 4675 14519 4681
rect 14461 4672 14473 4675
rect 14424 4644 14473 4672
rect 14424 4632 14430 4644
rect 14461 4641 14473 4644
rect 14507 4641 14519 4675
rect 14461 4635 14519 4641
rect 15194 4632 15200 4684
rect 15252 4672 15258 4684
rect 15565 4675 15623 4681
rect 15565 4672 15577 4675
rect 15252 4644 15577 4672
rect 15252 4632 15258 4644
rect 15565 4641 15577 4644
rect 15611 4641 15623 4675
rect 15948 4672 15976 4780
rect 19058 4768 19064 4780
rect 19116 4808 19122 4820
rect 20165 4811 20223 4817
rect 20165 4808 20177 4811
rect 19116 4780 20177 4808
rect 19116 4768 19122 4780
rect 20165 4777 20177 4780
rect 20211 4777 20223 4811
rect 24302 4808 24308 4820
rect 24263 4780 24308 4808
rect 20165 4771 20223 4777
rect 24302 4768 24308 4780
rect 24360 4768 24366 4820
rect 25038 4768 25044 4820
rect 25096 4808 25102 4820
rect 25409 4811 25467 4817
rect 25409 4808 25421 4811
rect 25096 4780 25421 4808
rect 25096 4768 25102 4780
rect 25409 4777 25421 4780
rect 25455 4777 25467 4811
rect 36630 4808 36636 4820
rect 36591 4780 36636 4808
rect 25409 4771 25467 4777
rect 36630 4768 36636 4780
rect 36688 4768 36694 4820
rect 17402 4740 17408 4752
rect 17236 4712 17408 4740
rect 16025 4675 16083 4681
rect 16025 4672 16037 4675
rect 15948 4644 16037 4672
rect 15565 4635 15623 4641
rect 16025 4641 16037 4644
rect 16071 4641 16083 4675
rect 16025 4635 16083 4641
rect 16114 4632 16120 4684
rect 16172 4672 16178 4684
rect 16301 4675 16359 4681
rect 16301 4672 16313 4675
rect 16172 4644 16313 4672
rect 16172 4632 16178 4644
rect 16301 4641 16313 4644
rect 16347 4641 16359 4675
rect 16850 4672 16856 4684
rect 16811 4644 16856 4672
rect 16301 4635 16359 4641
rect 16850 4632 16856 4644
rect 16908 4632 16914 4684
rect 17236 4681 17264 4712
rect 17402 4700 17408 4712
rect 17460 4700 17466 4752
rect 29181 4743 29239 4749
rect 29181 4709 29193 4743
rect 29227 4740 29239 4743
rect 29546 4740 29552 4752
rect 29227 4712 29552 4740
rect 29227 4709 29239 4712
rect 29181 4703 29239 4709
rect 29546 4700 29552 4712
rect 29604 4700 29610 4752
rect 32122 4740 32128 4752
rect 32083 4712 32128 4740
rect 32122 4700 32128 4712
rect 32180 4700 32186 4752
rect 17221 4675 17279 4681
rect 17221 4641 17233 4675
rect 17267 4641 17279 4675
rect 18233 4675 18291 4681
rect 18233 4672 18245 4675
rect 17221 4635 17279 4641
rect 17328 4644 18245 4672
rect 3694 4564 3700 4616
rect 3752 4604 3758 4616
rect 5813 4607 5871 4613
rect 5813 4604 5825 4607
rect 3752 4576 5825 4604
rect 3752 4564 3758 4576
rect 5813 4573 5825 4576
rect 5859 4573 5871 4607
rect 5813 4567 5871 4573
rect 6089 4607 6147 4613
rect 6089 4573 6101 4607
rect 6135 4604 6147 4607
rect 6914 4604 6920 4616
rect 6135 4576 6920 4604
rect 6135 4573 6147 4576
rect 6089 4567 6147 4573
rect 5828 4468 5856 4567
rect 6914 4564 6920 4576
rect 6972 4564 6978 4616
rect 9122 4604 9128 4616
rect 9083 4576 9128 4604
rect 9122 4564 9128 4576
rect 9180 4564 9186 4616
rect 10229 4607 10287 4613
rect 10229 4573 10241 4607
rect 10275 4604 10287 4607
rect 12345 4607 12403 4613
rect 12345 4604 12357 4607
rect 10275 4576 12357 4604
rect 10275 4573 10287 4576
rect 10229 4567 10287 4573
rect 12345 4573 12357 4576
rect 12391 4573 12403 4607
rect 12345 4567 12403 4573
rect 16485 4607 16543 4613
rect 16485 4573 16497 4607
rect 16531 4604 16543 4607
rect 17328 4604 17356 4644
rect 18233 4641 18245 4644
rect 18279 4641 18291 4675
rect 18233 4635 18291 4641
rect 19613 4675 19671 4681
rect 19613 4641 19625 4675
rect 19659 4672 19671 4675
rect 20073 4675 20131 4681
rect 20073 4672 20085 4675
rect 19659 4644 20085 4672
rect 19659 4641 19671 4644
rect 19613 4635 19671 4641
rect 20073 4641 20085 4644
rect 20119 4641 20131 4675
rect 20073 4635 20131 4641
rect 20806 4632 20812 4684
rect 20864 4672 20870 4684
rect 21269 4675 21327 4681
rect 21269 4672 21281 4675
rect 20864 4644 21281 4672
rect 20864 4632 20870 4644
rect 21269 4641 21281 4644
rect 21315 4641 21327 4675
rect 21269 4635 21327 4641
rect 21450 4632 21456 4684
rect 21508 4672 21514 4684
rect 21729 4675 21787 4681
rect 21729 4672 21741 4675
rect 21508 4644 21741 4672
rect 21508 4632 21514 4644
rect 21729 4641 21741 4644
rect 21775 4641 21787 4675
rect 21729 4635 21787 4641
rect 21818 4632 21824 4684
rect 21876 4672 21882 4684
rect 22925 4675 22983 4681
rect 22925 4672 22937 4675
rect 21876 4644 22937 4672
rect 21876 4632 21882 4644
rect 22925 4641 22937 4644
rect 22971 4672 22983 4675
rect 24854 4672 24860 4684
rect 22971 4644 24860 4672
rect 22971 4641 22983 4644
rect 22925 4635 22983 4641
rect 24854 4632 24860 4644
rect 24912 4632 24918 4684
rect 25317 4675 25375 4681
rect 25317 4641 25329 4675
rect 25363 4672 25375 4675
rect 26142 4672 26148 4684
rect 25363 4644 26148 4672
rect 25363 4641 25375 4644
rect 25317 4635 25375 4641
rect 26142 4632 26148 4644
rect 26200 4632 26206 4684
rect 27614 4672 27620 4684
rect 27575 4644 27620 4672
rect 27614 4632 27620 4644
rect 27672 4632 27678 4684
rect 27798 4632 27804 4684
rect 27856 4672 27862 4684
rect 27893 4675 27951 4681
rect 27893 4672 27905 4675
rect 27856 4644 27905 4672
rect 27856 4632 27862 4644
rect 27893 4641 27905 4644
rect 27939 4641 27951 4675
rect 27893 4635 27951 4641
rect 29362 4632 29368 4684
rect 29420 4672 29426 4684
rect 29733 4675 29791 4681
rect 29733 4672 29745 4675
rect 29420 4644 29745 4672
rect 29420 4632 29426 4644
rect 29733 4641 29745 4644
rect 29779 4641 29791 4675
rect 29733 4635 29791 4641
rect 30009 4675 30067 4681
rect 30009 4641 30021 4675
rect 30055 4672 30067 4675
rect 31386 4672 31392 4684
rect 30055 4644 31392 4672
rect 30055 4641 30067 4644
rect 30009 4635 30067 4641
rect 31386 4632 31392 4644
rect 31444 4632 31450 4684
rect 32582 4632 32588 4684
rect 32640 4672 32646 4684
rect 34330 4681 34336 4684
rect 32677 4675 32735 4681
rect 32677 4672 32689 4675
rect 32640 4644 32689 4672
rect 32640 4632 32646 4644
rect 32677 4641 32689 4644
rect 32723 4641 32735 4675
rect 32677 4635 32735 4641
rect 32953 4675 33011 4681
rect 32953 4641 32965 4675
rect 32999 4672 33011 4675
rect 34287 4675 34336 4681
rect 34287 4672 34299 4675
rect 32999 4644 34299 4672
rect 32999 4641 33011 4644
rect 32953 4635 33011 4641
rect 34287 4641 34299 4644
rect 34333 4641 34336 4675
rect 34287 4635 34336 4641
rect 34330 4632 34336 4635
rect 34388 4632 34394 4684
rect 34422 4632 34428 4684
rect 34480 4672 34486 4684
rect 34480 4644 34525 4672
rect 34480 4632 34486 4644
rect 17954 4604 17960 4616
rect 16531 4576 17356 4604
rect 17915 4576 17960 4604
rect 16531 4573 16543 4576
rect 16485 4567 16543 4573
rect 8110 4496 8116 4548
rect 8168 4536 8174 4548
rect 10042 4536 10048 4548
rect 8168 4508 10048 4536
rect 8168 4496 8174 4508
rect 10042 4496 10048 4508
rect 10100 4536 10106 4548
rect 10244 4536 10272 4567
rect 17954 4564 17960 4576
rect 18012 4564 18018 4616
rect 21085 4607 21143 4613
rect 21085 4573 21097 4607
rect 21131 4604 21143 4607
rect 21542 4604 21548 4616
rect 21131 4576 21548 4604
rect 21131 4573 21143 4576
rect 21085 4567 21143 4573
rect 21542 4564 21548 4576
rect 21600 4564 21606 4616
rect 23201 4607 23259 4613
rect 23201 4573 23213 4607
rect 23247 4604 23259 4607
rect 27065 4607 27123 4613
rect 27065 4604 27077 4607
rect 23247 4576 27077 4604
rect 23247 4573 23259 4576
rect 23201 4567 23259 4573
rect 27065 4573 27077 4576
rect 27111 4573 27123 4607
rect 27065 4567 27123 4573
rect 28077 4607 28135 4613
rect 28077 4573 28089 4607
rect 28123 4604 28135 4607
rect 28994 4604 29000 4616
rect 28123 4576 29000 4604
rect 28123 4573 28135 4576
rect 28077 4567 28135 4573
rect 28994 4564 29000 4576
rect 29052 4604 29058 4616
rect 30193 4607 30251 4613
rect 30193 4604 30205 4607
rect 29052 4576 30205 4604
rect 29052 4564 29058 4576
rect 30193 4573 30205 4576
rect 30239 4604 30251 4607
rect 31018 4604 31024 4616
rect 30239 4576 31024 4604
rect 30239 4573 30251 4576
rect 30193 4567 30251 4573
rect 31018 4564 31024 4576
rect 31076 4564 31082 4616
rect 31754 4564 31760 4616
rect 31812 4604 31818 4616
rect 32815 4607 32873 4613
rect 32815 4604 32827 4607
rect 31812 4576 32827 4604
rect 31812 4564 31818 4576
rect 32815 4573 32827 4576
rect 32861 4573 32873 4607
rect 33594 4604 33600 4616
rect 33555 4576 33600 4604
rect 32815 4567 32873 4573
rect 33594 4564 33600 4576
rect 33652 4564 33658 4616
rect 34149 4607 34207 4613
rect 34149 4573 34161 4607
rect 34195 4604 34207 4607
rect 34514 4604 34520 4616
rect 34195 4576 34520 4604
rect 34195 4573 34207 4576
rect 34149 4567 34207 4573
rect 34514 4564 34520 4576
rect 34572 4564 34578 4616
rect 35069 4607 35127 4613
rect 35069 4573 35081 4607
rect 35115 4573 35127 4607
rect 35342 4604 35348 4616
rect 35303 4576 35348 4604
rect 35069 4567 35127 4573
rect 10100 4508 10272 4536
rect 10100 4496 10106 4508
rect 13446 4496 13452 4548
rect 13504 4536 13510 4548
rect 14553 4539 14611 4545
rect 14553 4536 14565 4539
rect 13504 4508 14565 4536
rect 13504 4496 13510 4508
rect 14553 4505 14565 4508
rect 14599 4505 14611 4539
rect 14553 4499 14611 4505
rect 20714 4496 20720 4548
rect 20772 4536 20778 4548
rect 21729 4539 21787 4545
rect 21729 4536 21741 4539
rect 20772 4508 21741 4536
rect 20772 4496 20778 4508
rect 21729 4505 21741 4508
rect 21775 4505 21787 4539
rect 21729 4499 21787 4505
rect 26878 4496 26884 4548
rect 26936 4536 26942 4548
rect 35084 4536 35112 4567
rect 35342 4564 35348 4576
rect 35400 4564 35406 4616
rect 26936 4508 35112 4536
rect 26936 4496 26942 4508
rect 7006 4468 7012 4480
rect 5828 4440 7012 4468
rect 7006 4428 7012 4440
rect 7064 4428 7070 4480
rect 1104 4378 39836 4400
rect 1104 4326 4246 4378
rect 4298 4326 4310 4378
rect 4362 4326 4374 4378
rect 4426 4326 4438 4378
rect 4490 4326 34966 4378
rect 35018 4326 35030 4378
rect 35082 4326 35094 4378
rect 35146 4326 35158 4378
rect 35210 4326 39836 4378
rect 1104 4304 39836 4326
rect 5810 4224 5816 4276
rect 5868 4264 5874 4276
rect 35894 4264 35900 4276
rect 5868 4236 35900 4264
rect 5868 4224 5874 4236
rect 35894 4224 35900 4236
rect 35952 4224 35958 4276
rect 8570 4196 8576 4208
rect 7392 4168 8576 4196
rect 3694 4128 3700 4140
rect 3655 4100 3700 4128
rect 3694 4088 3700 4100
rect 3752 4088 3758 4140
rect 3973 4131 4031 4137
rect 3973 4097 3985 4131
rect 4019 4128 4031 4131
rect 4062 4128 4068 4140
rect 4019 4100 4068 4128
rect 4019 4097 4031 4100
rect 3973 4091 4031 4097
rect 4062 4088 4068 4100
rect 4120 4088 4126 4140
rect 6362 4088 6368 4140
rect 6420 4128 6426 4140
rect 6420 4100 7236 4128
rect 6420 4088 6426 4100
rect 5994 4060 6000 4072
rect 5955 4032 6000 4060
rect 5994 4020 6000 4032
rect 6052 4020 6058 4072
rect 7098 4060 7104 4072
rect 7059 4032 7104 4060
rect 7098 4020 7104 4032
rect 7156 4020 7162 4072
rect 7116 3992 7144 4020
rect 6196 3964 7144 3992
rect 7208 3992 7236 4100
rect 7392 4069 7420 4168
rect 8570 4156 8576 4168
rect 8628 4156 8634 4208
rect 15396 4168 19196 4196
rect 15396 4140 15424 4168
rect 8110 4088 8116 4140
rect 8168 4128 8174 4140
rect 8764 4131 8822 4137
rect 8764 4128 8776 4131
rect 8168 4100 8776 4128
rect 8168 4088 8174 4100
rect 8764 4097 8776 4100
rect 8810 4097 8822 4131
rect 9027 4131 9085 4137
rect 9027 4128 9039 4131
rect 8764 4091 8822 4097
rect 8956 4100 9039 4128
rect 7377 4063 7435 4069
rect 7377 4029 7389 4063
rect 7423 4029 7435 4063
rect 7377 4023 7435 4029
rect 8021 4063 8079 4069
rect 8021 4029 8033 4063
rect 8067 4029 8079 4063
rect 8021 4023 8079 4029
rect 8036 3992 8064 4023
rect 8478 4020 8484 4072
rect 8536 4060 8542 4072
rect 8956 4060 8984 4100
rect 9027 4097 9039 4100
rect 9073 4097 9085 4131
rect 9027 4091 9085 4097
rect 9214 4088 9220 4140
rect 9272 4128 9278 4140
rect 12894 4128 12900 4140
rect 9272 4100 12900 4128
rect 9272 4088 9278 4100
rect 12894 4088 12900 4100
rect 12952 4088 12958 4140
rect 14734 4128 14740 4140
rect 14695 4100 14740 4128
rect 14734 4088 14740 4100
rect 14792 4088 14798 4140
rect 15378 4088 15384 4140
rect 15436 4088 15442 4140
rect 16117 4131 16175 4137
rect 16117 4097 16129 4131
rect 16163 4128 16175 4131
rect 16298 4128 16304 4140
rect 16163 4100 16304 4128
rect 16163 4097 16175 4100
rect 16117 4091 16175 4097
rect 16298 4088 16304 4100
rect 16356 4088 16362 4140
rect 17497 4131 17555 4137
rect 17497 4097 17509 4131
rect 17543 4128 17555 4131
rect 17770 4128 17776 4140
rect 17543 4100 17776 4128
rect 17543 4097 17555 4100
rect 17497 4091 17555 4097
rect 17770 4088 17776 4100
rect 17828 4088 17834 4140
rect 8536 4032 8984 4060
rect 8536 4020 8542 4032
rect 9306 4020 9312 4072
rect 9364 4060 9370 4072
rect 10413 4063 10471 4069
rect 9364 4032 10272 4060
rect 9364 4020 9370 4032
rect 7208 3964 8064 3992
rect 5258 3924 5264 3936
rect 5219 3896 5264 3924
rect 5258 3884 5264 3896
rect 5316 3884 5322 3936
rect 6196 3933 6224 3964
rect 6181 3927 6239 3933
rect 6181 3893 6193 3927
rect 6227 3893 6239 3927
rect 6914 3924 6920 3936
rect 6875 3896 6920 3924
rect 6181 3887 6239 3893
rect 6914 3884 6920 3896
rect 6972 3884 6978 3936
rect 8205 3927 8263 3933
rect 8205 3893 8217 3927
rect 8251 3924 8263 3927
rect 10042 3924 10048 3936
rect 8251 3896 10048 3924
rect 8251 3893 8263 3896
rect 8205 3887 8263 3893
rect 10042 3884 10048 3896
rect 10100 3884 10106 3936
rect 10244 3924 10272 4032
rect 10413 4029 10425 4063
rect 10459 4060 10471 4063
rect 11238 4060 11244 4072
rect 10459 4032 11244 4060
rect 10459 4029 10471 4032
rect 10413 4023 10471 4029
rect 11238 4020 11244 4032
rect 11296 4020 11302 4072
rect 11333 4063 11391 4069
rect 11333 4029 11345 4063
rect 11379 4029 11391 4063
rect 11514 4060 11520 4072
rect 11475 4032 11520 4060
rect 11333 4023 11391 4029
rect 10318 3952 10324 4004
rect 10376 3992 10382 4004
rect 11348 3992 11376 4023
rect 11514 4020 11520 4032
rect 11572 4020 11578 4072
rect 13262 4060 13268 4072
rect 11716 4032 13268 4060
rect 11716 3992 11744 4032
rect 13262 4020 13268 4032
rect 13320 4020 13326 4072
rect 13446 4060 13452 4072
rect 13407 4032 13452 4060
rect 13446 4020 13452 4032
rect 13504 4020 13510 4072
rect 14458 4060 14464 4072
rect 14419 4032 14464 4060
rect 14458 4020 14464 4032
rect 14516 4020 14522 4072
rect 16761 4063 16819 4069
rect 16761 4060 16773 4063
rect 16408 4032 16773 4060
rect 10376 3964 11744 3992
rect 11793 3995 11851 4001
rect 10376 3952 10382 3964
rect 11793 3961 11805 3995
rect 11839 3992 11851 3995
rect 11882 3992 11888 4004
rect 11839 3964 11888 3992
rect 11839 3961 11851 3964
rect 11793 3955 11851 3961
rect 11882 3952 11888 3964
rect 11940 3952 11946 4004
rect 13725 3995 13783 4001
rect 13725 3961 13737 3995
rect 13771 3992 13783 3995
rect 13814 3992 13820 4004
rect 13771 3964 13820 3992
rect 13771 3961 13783 3964
rect 13725 3955 13783 3961
rect 13814 3952 13820 3964
rect 13872 3952 13878 4004
rect 16408 3924 16436 4032
rect 16761 4029 16773 4032
rect 16807 4029 16819 4063
rect 17218 4060 17224 4072
rect 17179 4032 17224 4060
rect 16761 4023 16819 4029
rect 16776 3992 16804 4023
rect 17218 4020 17224 4032
rect 17276 4020 17282 4072
rect 18601 4063 18659 4069
rect 18601 4029 18613 4063
rect 18647 4060 18659 4063
rect 18690 4060 18696 4072
rect 18647 4032 18696 4060
rect 18647 4029 18659 4032
rect 18601 4023 18659 4029
rect 18138 3992 18144 4004
rect 16776 3964 18144 3992
rect 18138 3952 18144 3964
rect 18196 3992 18202 4004
rect 18616 3992 18644 4023
rect 18690 4020 18696 4032
rect 18748 4020 18754 4072
rect 19058 4060 19064 4072
rect 19019 4032 19064 4060
rect 19058 4020 19064 4032
rect 19116 4020 19122 4072
rect 19168 4060 19196 4168
rect 22094 4156 22100 4208
rect 22152 4156 22158 4208
rect 29196 4168 29408 4196
rect 19242 4088 19248 4140
rect 19300 4128 19306 4140
rect 20257 4131 20315 4137
rect 20257 4128 20269 4131
rect 19300 4100 20269 4128
rect 19300 4088 19306 4100
rect 20257 4097 20269 4100
rect 20303 4097 20315 4131
rect 20257 4091 20315 4097
rect 20438 4088 20444 4140
rect 20496 4088 20502 4140
rect 21637 4131 21695 4137
rect 21637 4097 21649 4131
rect 21683 4128 21695 4131
rect 22112 4128 22140 4156
rect 21683 4100 22140 4128
rect 22649 4131 22707 4137
rect 21683 4097 21695 4100
rect 21637 4091 21695 4097
rect 22649 4097 22661 4131
rect 22695 4128 22707 4131
rect 26418 4128 26424 4140
rect 22695 4100 26424 4128
rect 22695 4097 22707 4100
rect 22649 4091 22707 4097
rect 26418 4088 26424 4100
rect 26476 4088 26482 4140
rect 26694 4088 26700 4140
rect 26752 4128 26758 4140
rect 29196 4128 29224 4168
rect 26752 4100 29224 4128
rect 29380 4128 29408 4168
rect 29454 4156 29460 4208
rect 29512 4196 29518 4208
rect 33962 4196 33968 4208
rect 29512 4168 29557 4196
rect 31220 4168 33968 4196
rect 29512 4156 29518 4168
rect 30926 4128 30932 4140
rect 29380 4100 30512 4128
rect 30887 4100 30932 4128
rect 26752 4088 26758 4100
rect 19978 4060 19984 4072
rect 19168 4032 19840 4060
rect 19939 4032 19984 4060
rect 19334 3992 19340 4004
rect 18196 3964 18644 3992
rect 19295 3964 19340 3992
rect 18196 3952 18202 3964
rect 19334 3952 19340 3964
rect 19392 3952 19398 4004
rect 19812 3992 19840 4032
rect 19978 4020 19984 4032
rect 20036 4020 20042 4072
rect 20456 4060 20484 4088
rect 20088 4032 20484 4060
rect 20088 3992 20116 4032
rect 21726 4020 21732 4072
rect 21784 4060 21790 4072
rect 22097 4063 22155 4069
rect 22097 4060 22109 4063
rect 21784 4032 22109 4060
rect 21784 4020 21790 4032
rect 22097 4029 22109 4032
rect 22143 4029 22155 4063
rect 22097 4023 22155 4029
rect 22186 4020 22192 4072
rect 22244 4060 22250 4072
rect 25593 4063 25651 4069
rect 22244 4032 22289 4060
rect 22244 4020 22250 4032
rect 25593 4029 25605 4063
rect 25639 4029 25651 4063
rect 25866 4060 25872 4072
rect 25827 4032 25872 4060
rect 25593 4023 25651 4029
rect 19812 3964 20116 3992
rect 20990 3952 20996 4004
rect 21048 3992 21054 4004
rect 24486 3992 24492 4004
rect 21048 3964 24492 3992
rect 21048 3952 21054 3964
rect 24486 3952 24492 3964
rect 24544 3952 24550 4004
rect 25041 3995 25099 4001
rect 25041 3961 25053 3995
rect 25087 3961 25099 3995
rect 25608 3992 25636 4023
rect 25866 4020 25872 4032
rect 25924 4020 25930 4072
rect 26050 4060 26056 4072
rect 26011 4032 26056 4060
rect 26050 4020 26056 4032
rect 26108 4020 26114 4072
rect 26326 4020 26332 4072
rect 26384 4060 26390 4072
rect 26513 4063 26571 4069
rect 26513 4060 26525 4063
rect 26384 4032 26525 4060
rect 26384 4020 26390 4032
rect 26513 4029 26525 4032
rect 26559 4029 26571 4063
rect 26513 4023 26571 4029
rect 26789 4063 26847 4069
rect 26789 4029 26801 4063
rect 26835 4060 26847 4063
rect 27062 4060 27068 4072
rect 26835 4032 27068 4060
rect 26835 4029 26847 4032
rect 26789 4023 26847 4029
rect 27062 4020 27068 4032
rect 27120 4020 27126 4072
rect 29270 4020 29276 4072
rect 29328 4060 29334 4072
rect 29328 4032 29373 4060
rect 29328 4020 29334 4032
rect 25608 3964 26556 3992
rect 25041 3955 25099 3961
rect 10244 3896 16436 3924
rect 17862 3884 17868 3936
rect 17920 3924 17926 3936
rect 18414 3924 18420 3936
rect 17920 3896 18420 3924
rect 17920 3884 17926 3896
rect 18414 3884 18420 3896
rect 18472 3884 18478 3936
rect 18966 3884 18972 3936
rect 19024 3924 19030 3936
rect 23750 3924 23756 3936
rect 19024 3896 23756 3924
rect 19024 3884 19030 3896
rect 23750 3884 23756 3896
rect 23808 3884 23814 3936
rect 25056 3924 25084 3955
rect 26528 3936 26556 3964
rect 27522 3952 27528 4004
rect 27580 3992 27586 4004
rect 30377 3995 30435 4001
rect 30377 3992 30389 3995
rect 27580 3964 29224 3992
rect 27580 3952 27586 3964
rect 26418 3924 26424 3936
rect 25056 3896 26424 3924
rect 26418 3884 26424 3896
rect 26476 3884 26482 3936
rect 26510 3884 26516 3936
rect 26568 3884 26574 3936
rect 27890 3924 27896 3936
rect 27851 3896 27896 3924
rect 27890 3884 27896 3896
rect 27948 3884 27954 3936
rect 29196 3924 29224 3964
rect 29380 3964 30389 3992
rect 29380 3924 29408 3964
rect 30377 3961 30389 3964
rect 30423 3961 30435 3995
rect 30377 3955 30435 3961
rect 29196 3896 29408 3924
rect 30484 3924 30512 4100
rect 30926 4088 30932 4100
rect 30984 4088 30990 4140
rect 31220 4069 31248 4168
rect 33962 4156 33968 4168
rect 34020 4156 34026 4208
rect 34422 4196 34428 4208
rect 34164 4168 34428 4196
rect 31938 4088 31944 4140
rect 31996 4128 32002 4140
rect 32766 4128 32772 4140
rect 31996 4100 32772 4128
rect 31996 4088 32002 4100
rect 31205 4063 31263 4069
rect 31205 4029 31217 4063
rect 31251 4029 31263 4063
rect 31205 4023 31263 4029
rect 31389 4063 31447 4069
rect 31389 4029 31401 4063
rect 31435 4060 31447 4063
rect 31754 4060 31760 4072
rect 31435 4032 31760 4060
rect 31435 4029 31447 4032
rect 31389 4023 31447 4029
rect 31754 4020 31760 4032
rect 31812 4020 31818 4072
rect 32122 4020 32128 4072
rect 32180 4060 32186 4072
rect 32692 4069 32720 4100
rect 32766 4088 32772 4100
rect 32824 4088 32830 4140
rect 33042 4088 33048 4140
rect 33100 4128 33106 4140
rect 34164 4128 34192 4168
rect 34422 4156 34428 4168
rect 34480 4156 34486 4208
rect 33100 4100 34192 4128
rect 33100 4088 33106 4100
rect 32401 4063 32459 4069
rect 32401 4060 32413 4063
rect 32180 4032 32413 4060
rect 32180 4020 32186 4032
rect 32401 4029 32413 4032
rect 32447 4029 32459 4063
rect 32401 4023 32459 4029
rect 32677 4063 32735 4069
rect 32677 4029 32689 4063
rect 32723 4029 32735 4063
rect 32858 4060 32864 4072
rect 32819 4032 32864 4060
rect 32677 4023 32735 4029
rect 32858 4020 32864 4032
rect 32916 4020 32922 4072
rect 33870 4060 33876 4072
rect 33831 4032 33876 4060
rect 33870 4020 33876 4032
rect 33928 4020 33934 4072
rect 33962 4020 33968 4072
rect 34020 4069 34026 4072
rect 34164 4069 34192 4100
rect 34606 4088 34612 4140
rect 34664 4128 34670 4140
rect 34885 4131 34943 4137
rect 34885 4128 34897 4131
rect 34664 4100 34897 4128
rect 34664 4088 34670 4100
rect 34885 4097 34897 4100
rect 34931 4097 34943 4131
rect 35575 4131 35633 4137
rect 35575 4128 35587 4131
rect 34885 4091 34943 4097
rect 34992 4100 35587 4128
rect 34020 4063 34069 4069
rect 34020 4029 34023 4063
rect 34057 4029 34069 4063
rect 34020 4023 34069 4029
rect 34149 4063 34207 4069
rect 34149 4029 34161 4063
rect 34195 4029 34207 4063
rect 34149 4023 34207 4029
rect 34020 4020 34026 4023
rect 34422 4020 34428 4072
rect 34480 4060 34486 4072
rect 34992 4060 35020 4100
rect 35575 4097 35587 4100
rect 35621 4097 35633 4131
rect 35986 4128 35992 4140
rect 35575 4091 35633 4097
rect 35728 4100 35992 4128
rect 35434 4060 35440 4072
rect 34480 4032 35020 4060
rect 35395 4032 35440 4060
rect 34480 4020 34486 4032
rect 35434 4020 35440 4032
rect 35492 4020 35498 4072
rect 35728 4069 35756 4100
rect 35986 4088 35992 4100
rect 36044 4088 36050 4140
rect 35713 4063 35771 4069
rect 35713 4029 35725 4063
rect 35759 4029 35771 4063
rect 35713 4023 35771 4029
rect 31846 3992 31852 4004
rect 31807 3964 31852 3992
rect 31846 3952 31852 3964
rect 31904 3952 31910 4004
rect 32030 3952 32036 4004
rect 32088 3992 32094 4004
rect 33321 3995 33379 4001
rect 33321 3992 33333 3995
rect 32088 3964 33333 3992
rect 32088 3952 32094 3964
rect 33321 3961 33333 3964
rect 33367 3961 33379 3995
rect 33321 3955 33379 3961
rect 35342 3924 35348 3936
rect 30484 3896 35348 3924
rect 35342 3884 35348 3896
rect 35400 3884 35406 3936
rect 1104 3834 39836 3856
rect 1104 3782 19606 3834
rect 19658 3782 19670 3834
rect 19722 3782 19734 3834
rect 19786 3782 19798 3834
rect 19850 3782 39836 3834
rect 1104 3760 39836 3782
rect 7193 3723 7251 3729
rect 7193 3689 7205 3723
rect 7239 3720 7251 3723
rect 7374 3720 7380 3732
rect 7239 3692 7380 3720
rect 7239 3689 7251 3692
rect 7193 3683 7251 3689
rect 7374 3680 7380 3692
rect 7432 3680 7438 3732
rect 7466 3680 7472 3732
rect 7524 3720 7530 3732
rect 9769 3723 9827 3729
rect 9769 3720 9781 3723
rect 7524 3692 9781 3720
rect 7524 3680 7530 3692
rect 9769 3689 9781 3692
rect 9815 3689 9827 3723
rect 20990 3720 20996 3732
rect 9769 3683 9827 3689
rect 9876 3692 20996 3720
rect 5994 3612 6000 3664
rect 6052 3652 6058 3664
rect 6052 3624 8708 3652
rect 6052 3612 6058 3624
rect 5258 3584 5264 3596
rect 5219 3556 5264 3584
rect 5258 3544 5264 3556
rect 5316 3544 5322 3596
rect 6362 3584 6368 3596
rect 6323 3556 6368 3584
rect 6362 3544 6368 3556
rect 6420 3544 6426 3596
rect 7098 3584 7104 3596
rect 7059 3556 7104 3584
rect 7098 3544 7104 3556
rect 7156 3544 7162 3596
rect 7837 3587 7895 3593
rect 7837 3553 7849 3587
rect 7883 3584 7895 3587
rect 8570 3584 8576 3596
rect 7883 3556 8576 3584
rect 7883 3553 7895 3556
rect 7837 3547 7895 3553
rect 8570 3544 8576 3556
rect 8628 3544 8634 3596
rect 8680 3593 8708 3624
rect 8754 3612 8760 3664
rect 8812 3652 8818 3664
rect 9876 3652 9904 3692
rect 20990 3680 20996 3692
rect 21048 3680 21054 3732
rect 27062 3720 27068 3732
rect 24964 3692 27068 3720
rect 10318 3652 10324 3664
rect 8812 3624 9904 3652
rect 9968 3624 10324 3652
rect 8812 3612 8818 3624
rect 8665 3587 8723 3593
rect 8665 3553 8677 3587
rect 8711 3584 8723 3587
rect 8938 3584 8944 3596
rect 8711 3556 8944 3584
rect 8711 3553 8723 3556
rect 8665 3547 8723 3553
rect 8938 3544 8944 3556
rect 8996 3544 9002 3596
rect 9968 3593 9996 3624
rect 10318 3612 10324 3624
rect 10376 3612 10382 3664
rect 10410 3612 10416 3664
rect 10468 3652 10474 3664
rect 24964 3661 24992 3692
rect 27062 3680 27068 3692
rect 27120 3680 27126 3732
rect 27816 3692 30052 3720
rect 10965 3655 11023 3661
rect 10965 3652 10977 3655
rect 10468 3624 10977 3652
rect 10468 3612 10474 3624
rect 10965 3621 10977 3624
rect 11011 3621 11023 3655
rect 24949 3655 25007 3661
rect 10965 3615 11023 3621
rect 17880 3624 18184 3652
rect 9953 3587 10011 3593
rect 9953 3553 9965 3587
rect 9999 3553 10011 3587
rect 10134 3584 10140 3596
rect 10095 3556 10140 3584
rect 9953 3547 10011 3553
rect 5166 3516 5172 3528
rect 5127 3488 5172 3516
rect 5166 3476 5172 3488
rect 5224 3476 5230 3528
rect 5718 3516 5724 3528
rect 5679 3488 5724 3516
rect 5718 3476 5724 3488
rect 5776 3476 5782 3528
rect 7929 3519 7987 3525
rect 7929 3516 7941 3519
rect 7116 3488 7941 3516
rect 6086 3408 6092 3460
rect 6144 3448 6150 3460
rect 6822 3448 6828 3460
rect 6144 3420 6828 3448
rect 6144 3408 6150 3420
rect 6822 3408 6828 3420
rect 6880 3448 6886 3460
rect 7116 3448 7144 3488
rect 7929 3485 7941 3488
rect 7975 3485 7987 3519
rect 7929 3479 7987 3485
rect 6880 3420 7144 3448
rect 6880 3408 6886 3420
rect 8662 3408 8668 3460
rect 8720 3448 8726 3460
rect 8849 3451 8907 3457
rect 8849 3448 8861 3451
rect 8720 3420 8861 3448
rect 8720 3408 8726 3420
rect 8849 3417 8861 3420
rect 8895 3448 8907 3451
rect 9968 3448 9996 3547
rect 10134 3544 10140 3556
rect 10192 3544 10198 3596
rect 10873 3587 10931 3593
rect 10873 3553 10885 3587
rect 10919 3584 10931 3587
rect 11238 3584 11244 3596
rect 10919 3556 11244 3584
rect 10919 3553 10931 3556
rect 10873 3547 10931 3553
rect 11238 3544 11244 3556
rect 11296 3544 11302 3596
rect 11882 3584 11888 3596
rect 11843 3556 11888 3584
rect 11882 3544 11888 3556
rect 11940 3544 11946 3596
rect 13262 3544 13268 3596
rect 13320 3584 13326 3596
rect 13725 3587 13783 3593
rect 13725 3584 13737 3587
rect 13320 3556 13737 3584
rect 13320 3544 13326 3556
rect 13725 3553 13737 3556
rect 13771 3553 13783 3587
rect 14182 3584 14188 3596
rect 14143 3556 14188 3584
rect 13725 3547 13783 3553
rect 14182 3544 14188 3556
rect 14240 3544 14246 3596
rect 14458 3544 14464 3596
rect 14516 3584 14522 3596
rect 15933 3587 15991 3593
rect 15933 3584 15945 3587
rect 14516 3556 15945 3584
rect 14516 3544 14522 3556
rect 15933 3553 15945 3556
rect 15979 3553 15991 3587
rect 16206 3584 16212 3596
rect 16167 3556 16212 3584
rect 15933 3547 15991 3553
rect 10410 3476 10416 3528
rect 10468 3516 10474 3528
rect 11609 3519 11667 3525
rect 11609 3516 11621 3519
rect 10468 3488 11621 3516
rect 10468 3476 10474 3488
rect 11609 3485 11621 3488
rect 11655 3516 11667 3519
rect 13538 3516 13544 3528
rect 11655 3488 13544 3516
rect 11655 3485 11667 3488
rect 11609 3479 11667 3485
rect 13538 3476 13544 3488
rect 13596 3476 13602 3528
rect 14274 3516 14280 3528
rect 14235 3488 14280 3516
rect 14274 3476 14280 3488
rect 14332 3476 14338 3528
rect 15948 3516 15976 3547
rect 16206 3544 16212 3556
rect 16264 3544 16270 3596
rect 16298 3544 16304 3596
rect 16356 3584 16362 3596
rect 17880 3584 17908 3624
rect 18046 3584 18052 3596
rect 16356 3556 17908 3584
rect 18007 3556 18052 3584
rect 16356 3544 16362 3556
rect 18046 3544 18052 3556
rect 18104 3544 18110 3596
rect 18156 3584 18184 3624
rect 24949 3621 24961 3655
rect 24995 3621 25007 3655
rect 27433 3655 27491 3661
rect 27433 3652 27445 3655
rect 24949 3615 25007 3621
rect 25516 3624 27445 3652
rect 21358 3584 21364 3596
rect 18156 3556 20024 3584
rect 21319 3556 21364 3584
rect 17954 3516 17960 3528
rect 15948 3488 17960 3516
rect 17954 3476 17960 3488
rect 18012 3476 18018 3528
rect 18230 3476 18236 3528
rect 18288 3516 18294 3528
rect 18325 3519 18383 3525
rect 18325 3516 18337 3519
rect 18288 3488 18337 3516
rect 18288 3476 18294 3488
rect 18325 3485 18337 3488
rect 18371 3485 18383 3519
rect 18325 3479 18383 3485
rect 18414 3476 18420 3528
rect 18472 3516 18478 3528
rect 19886 3516 19892 3528
rect 18472 3488 19892 3516
rect 18472 3476 18478 3488
rect 19886 3476 19892 3488
rect 19944 3476 19950 3528
rect 19996 3516 20024 3556
rect 21358 3544 21364 3556
rect 21416 3544 21422 3596
rect 22557 3587 22615 3593
rect 22557 3553 22569 3587
rect 22603 3584 22615 3587
rect 22646 3584 22652 3596
rect 22603 3556 22652 3584
rect 22603 3553 22615 3556
rect 22557 3547 22615 3553
rect 22646 3544 22652 3556
rect 22704 3544 22710 3596
rect 22830 3584 22836 3596
rect 22791 3556 22836 3584
rect 22830 3544 22836 3556
rect 22888 3544 22894 3596
rect 25516 3593 25544 3624
rect 27433 3621 27445 3624
rect 27479 3621 27491 3655
rect 27433 3615 27491 3621
rect 25501 3587 25559 3593
rect 25501 3553 25513 3587
rect 25547 3553 25559 3587
rect 25501 3547 25559 3553
rect 25777 3587 25835 3593
rect 25777 3553 25789 3587
rect 25823 3584 25835 3587
rect 25866 3584 25872 3596
rect 25823 3556 25872 3584
rect 25823 3553 25835 3556
rect 25777 3547 25835 3553
rect 25866 3544 25872 3556
rect 25924 3584 25930 3596
rect 27816 3584 27844 3692
rect 27890 3612 27896 3664
rect 27948 3652 27954 3664
rect 30024 3652 30052 3692
rect 30098 3680 30104 3732
rect 30156 3720 30162 3732
rect 30282 3720 30288 3732
rect 30156 3692 30288 3720
rect 30156 3680 30162 3692
rect 30282 3680 30288 3692
rect 30340 3720 30346 3732
rect 30469 3723 30527 3729
rect 30469 3720 30481 3723
rect 30340 3692 30481 3720
rect 30340 3680 30346 3692
rect 30469 3689 30481 3692
rect 30515 3720 30527 3723
rect 30650 3720 30656 3732
rect 30515 3692 30656 3720
rect 30515 3689 30527 3692
rect 30469 3683 30527 3689
rect 30650 3680 30656 3692
rect 30708 3680 30714 3732
rect 31386 3680 31392 3732
rect 31444 3720 31450 3732
rect 32858 3720 32864 3732
rect 31444 3692 32864 3720
rect 31444 3680 31450 3692
rect 32858 3680 32864 3692
rect 32916 3680 32922 3732
rect 34330 3680 34336 3732
rect 34388 3720 34394 3732
rect 34977 3723 35035 3729
rect 34977 3720 34989 3723
rect 34388 3692 34989 3720
rect 34388 3680 34394 3692
rect 34977 3689 34989 3692
rect 35023 3689 35035 3723
rect 34977 3683 35035 3689
rect 31938 3652 31944 3664
rect 27948 3624 28488 3652
rect 30024 3624 31944 3652
rect 27948 3612 27954 3624
rect 27982 3584 27988 3596
rect 25924 3556 27844 3584
rect 27943 3556 27988 3584
rect 25924 3544 25930 3556
rect 27982 3544 27988 3556
rect 28040 3544 28046 3596
rect 28258 3584 28264 3596
rect 28219 3556 28264 3584
rect 28258 3544 28264 3556
rect 28316 3544 28322 3596
rect 28460 3593 28488 3624
rect 31938 3612 31944 3624
rect 31996 3612 32002 3664
rect 32122 3652 32128 3664
rect 32083 3624 32128 3652
rect 32122 3612 32128 3624
rect 32180 3612 32186 3664
rect 28445 3587 28503 3593
rect 28445 3553 28457 3587
rect 28491 3553 28503 3587
rect 28445 3547 28503 3553
rect 29181 3587 29239 3593
rect 29181 3553 29193 3587
rect 29227 3584 29239 3587
rect 31846 3584 31852 3596
rect 29227 3556 31852 3584
rect 29227 3553 29239 3556
rect 29181 3547 29239 3553
rect 31846 3544 31852 3556
rect 31904 3544 31910 3596
rect 32953 3587 33011 3593
rect 32953 3584 32965 3587
rect 32600 3556 32965 3584
rect 21269 3519 21327 3525
rect 21269 3516 21281 3519
rect 19996 3488 21281 3516
rect 21269 3485 21281 3488
rect 21315 3516 21327 3519
rect 21726 3516 21732 3528
rect 21315 3488 21732 3516
rect 21315 3485 21327 3488
rect 21269 3479 21327 3485
rect 21726 3476 21732 3488
rect 21784 3476 21790 3528
rect 21821 3519 21879 3525
rect 21821 3485 21833 3519
rect 21867 3516 21879 3519
rect 22094 3516 22100 3528
rect 21867 3488 22100 3516
rect 21867 3485 21879 3488
rect 21821 3479 21879 3485
rect 22094 3476 22100 3488
rect 22152 3476 22158 3528
rect 25961 3519 26019 3525
rect 25961 3485 25973 3519
rect 26007 3516 26019 3519
rect 27798 3516 27804 3528
rect 26007 3488 27804 3516
rect 26007 3485 26019 3488
rect 25961 3479 26019 3485
rect 27798 3476 27804 3488
rect 27856 3476 27862 3528
rect 28905 3519 28963 3525
rect 28905 3485 28917 3519
rect 28951 3516 28963 3519
rect 29086 3516 29092 3528
rect 28951 3488 29092 3516
rect 28951 3485 28963 3488
rect 28905 3479 28963 3485
rect 8895 3420 9996 3448
rect 8895 3417 8907 3420
rect 8849 3411 8907 3417
rect 10042 3408 10048 3460
rect 10100 3448 10106 3460
rect 11146 3448 11152 3460
rect 10100 3420 11152 3448
rect 10100 3408 10106 3420
rect 11146 3408 11152 3420
rect 11204 3408 11210 3460
rect 19058 3408 19064 3460
rect 19116 3448 19122 3460
rect 22278 3448 22284 3460
rect 19116 3420 22284 3448
rect 19116 3408 19122 3420
rect 22278 3408 22284 3420
rect 22336 3408 22342 3460
rect 23842 3408 23848 3460
rect 23900 3448 23906 3460
rect 26694 3448 26700 3460
rect 23900 3420 26700 3448
rect 23900 3408 23906 3420
rect 26694 3408 26700 3420
rect 26752 3408 26758 3460
rect 27062 3408 27068 3460
rect 27120 3448 27126 3460
rect 28920 3448 28948 3479
rect 29086 3476 29092 3488
rect 29144 3476 29150 3528
rect 29546 3476 29552 3528
rect 29604 3516 29610 3528
rect 29604 3488 30236 3516
rect 29604 3476 29610 3488
rect 27120 3420 28948 3448
rect 30208 3448 30236 3488
rect 30558 3476 30564 3528
rect 30616 3516 30622 3528
rect 32600 3516 32628 3556
rect 32953 3553 32965 3556
rect 32999 3584 33011 3587
rect 33410 3584 33416 3596
rect 32999 3556 33416 3584
rect 32999 3553 33011 3556
rect 32953 3547 33011 3553
rect 33410 3544 33416 3556
rect 33468 3544 33474 3596
rect 33686 3544 33692 3596
rect 33744 3584 33750 3596
rect 33873 3587 33931 3593
rect 33873 3584 33885 3587
rect 33744 3556 33885 3584
rect 33744 3544 33750 3556
rect 33873 3553 33885 3556
rect 33919 3553 33931 3587
rect 33873 3547 33931 3553
rect 35713 3587 35771 3593
rect 35713 3553 35725 3587
rect 35759 3584 35771 3587
rect 35986 3584 35992 3596
rect 35759 3556 35992 3584
rect 35759 3553 35771 3556
rect 35713 3547 35771 3553
rect 35986 3544 35992 3556
rect 36044 3544 36050 3596
rect 30616 3488 32628 3516
rect 30616 3476 30622 3488
rect 32674 3476 32680 3528
rect 32732 3516 32738 3528
rect 33137 3519 33195 3525
rect 33137 3516 33149 3519
rect 32732 3488 32777 3516
rect 32876 3488 33149 3516
rect 32732 3476 32738 3488
rect 32692 3448 32720 3476
rect 30208 3420 32720 3448
rect 27120 3408 27126 3420
rect 6546 3380 6552 3392
rect 6507 3352 6552 3380
rect 6546 3340 6552 3352
rect 6604 3340 6610 3392
rect 13173 3383 13231 3389
rect 13173 3349 13185 3383
rect 13219 3380 13231 3383
rect 16574 3380 16580 3392
rect 13219 3352 16580 3380
rect 13219 3349 13231 3352
rect 13173 3343 13231 3349
rect 16574 3340 16580 3352
rect 16632 3340 16638 3392
rect 17497 3383 17555 3389
rect 17497 3349 17509 3383
rect 17543 3380 17555 3383
rect 18322 3380 18328 3392
rect 17543 3352 18328 3380
rect 17543 3349 17555 3352
rect 17497 3343 17555 3349
rect 18322 3340 18328 3352
rect 18380 3340 18386 3392
rect 19613 3383 19671 3389
rect 19613 3349 19625 3383
rect 19659 3380 19671 3383
rect 21542 3380 21548 3392
rect 19659 3352 21548 3380
rect 19659 3349 19671 3352
rect 19613 3343 19671 3349
rect 21542 3340 21548 3352
rect 21600 3340 21606 3392
rect 24118 3380 24124 3392
rect 24079 3352 24124 3380
rect 24118 3340 24124 3352
rect 24176 3340 24182 3392
rect 24762 3340 24768 3392
rect 24820 3380 24826 3392
rect 26878 3380 26884 3392
rect 24820 3352 26884 3380
rect 24820 3340 24826 3352
rect 26878 3340 26884 3352
rect 26936 3340 26942 3392
rect 28258 3340 28264 3392
rect 28316 3380 28322 3392
rect 30558 3380 30564 3392
rect 28316 3352 30564 3380
rect 28316 3340 28322 3352
rect 30558 3340 30564 3352
rect 30616 3340 30622 3392
rect 30650 3340 30656 3392
rect 30708 3380 30714 3392
rect 32876 3380 32904 3488
rect 33137 3485 33149 3488
rect 33183 3485 33195 3519
rect 33137 3479 33195 3485
rect 33502 3476 33508 3528
rect 33560 3516 33566 3528
rect 33597 3519 33655 3525
rect 33597 3516 33609 3519
rect 33560 3488 33609 3516
rect 33560 3476 33566 3488
rect 33597 3485 33609 3488
rect 33643 3485 33655 3519
rect 33597 3479 33655 3485
rect 30708 3352 32904 3380
rect 30708 3340 30714 3352
rect 33410 3340 33416 3392
rect 33468 3380 33474 3392
rect 35710 3380 35716 3392
rect 33468 3352 35716 3380
rect 33468 3340 33474 3352
rect 35710 3340 35716 3352
rect 35768 3380 35774 3392
rect 35897 3383 35955 3389
rect 35897 3380 35909 3383
rect 35768 3352 35909 3380
rect 35768 3340 35774 3352
rect 35897 3349 35909 3352
rect 35943 3349 35955 3383
rect 35897 3343 35955 3349
rect 1104 3290 39836 3312
rect 1104 3238 4246 3290
rect 4298 3238 4310 3290
rect 4362 3238 4374 3290
rect 4426 3238 4438 3290
rect 4490 3238 34966 3290
rect 35018 3238 35030 3290
rect 35082 3238 35094 3290
rect 35146 3238 35158 3290
rect 35210 3238 39836 3290
rect 1104 3216 39836 3238
rect 6546 3136 6552 3188
rect 6604 3176 6610 3188
rect 10870 3176 10876 3188
rect 6604 3148 10272 3176
rect 10831 3148 10876 3176
rect 6604 3136 6610 3148
rect 1394 3000 1400 3052
rect 1452 3040 1458 3052
rect 1857 3043 1915 3049
rect 1857 3040 1869 3043
rect 1452 3012 1869 3040
rect 1452 3000 1458 3012
rect 1857 3009 1869 3012
rect 1903 3009 1915 3043
rect 1857 3003 1915 3009
rect 6273 3043 6331 3049
rect 6273 3009 6285 3043
rect 6319 3040 6331 3043
rect 7098 3040 7104 3052
rect 6319 3012 7104 3040
rect 6319 3009 6331 3012
rect 6273 3003 6331 3009
rect 7098 3000 7104 3012
rect 7156 3000 7162 3052
rect 7466 3040 7472 3052
rect 7427 3012 7472 3040
rect 7466 3000 7472 3012
rect 7524 3000 7530 3052
rect 9122 3000 9128 3052
rect 9180 3040 9186 3052
rect 9585 3043 9643 3049
rect 9585 3040 9597 3043
rect 9180 3012 9597 3040
rect 9180 3000 9186 3012
rect 9585 3009 9597 3012
rect 9631 3009 9643 3043
rect 10244 3040 10272 3148
rect 10870 3136 10876 3148
rect 10928 3136 10934 3188
rect 11054 3136 11060 3188
rect 11112 3176 11118 3188
rect 12713 3179 12771 3185
rect 12713 3176 12725 3179
rect 11112 3148 12725 3176
rect 11112 3136 11118 3148
rect 12713 3145 12725 3148
rect 12759 3145 12771 3179
rect 18230 3176 18236 3188
rect 12713 3139 12771 3145
rect 13556 3148 18236 3176
rect 11698 3068 11704 3120
rect 11756 3108 11762 3120
rect 13556 3108 13584 3148
rect 18230 3136 18236 3148
rect 18288 3136 18294 3188
rect 23842 3176 23848 3188
rect 19168 3148 23848 3176
rect 16114 3108 16120 3120
rect 11756 3080 13584 3108
rect 14936 3080 16120 3108
rect 11756 3068 11762 3080
rect 13538 3040 13544 3052
rect 10244 3012 13400 3040
rect 13499 3012 13544 3040
rect 9585 3003 9643 3009
rect 1946 2932 1952 2984
rect 2004 2972 2010 2984
rect 2133 2975 2191 2981
rect 2133 2972 2145 2975
rect 2004 2944 2145 2972
rect 2004 2932 2010 2944
rect 2133 2941 2145 2944
rect 2179 2941 2191 2975
rect 5810 2972 5816 2984
rect 5771 2944 5816 2972
rect 2133 2935 2191 2941
rect 5810 2932 5816 2944
rect 5868 2932 5874 2984
rect 6086 2972 6092 2984
rect 6047 2944 6092 2972
rect 6086 2932 6092 2944
rect 6144 2932 6150 2984
rect 6914 2932 6920 2984
rect 6972 2972 6978 2984
rect 7193 2975 7251 2981
rect 7193 2972 7205 2975
rect 6972 2944 7205 2972
rect 6972 2932 6978 2944
rect 7193 2941 7205 2944
rect 7239 2941 7251 2975
rect 7193 2935 7251 2941
rect 9309 2975 9367 2981
rect 9309 2941 9321 2975
rect 9355 2972 9367 2975
rect 10410 2972 10416 2984
rect 9355 2944 10416 2972
rect 9355 2941 9367 2944
rect 9309 2935 9367 2941
rect 10410 2932 10416 2944
rect 10468 2932 10474 2984
rect 11146 2932 11152 2984
rect 11204 2972 11210 2984
rect 12342 2972 12348 2984
rect 11204 2944 12348 2972
rect 11204 2932 11210 2944
rect 12342 2932 12348 2944
rect 12400 2972 12406 2984
rect 12437 2975 12495 2981
rect 12437 2972 12449 2975
rect 12400 2944 12449 2972
rect 12400 2932 12406 2944
rect 12437 2941 12449 2944
rect 12483 2941 12495 2975
rect 12437 2935 12495 2941
rect 12529 2975 12587 2981
rect 12529 2941 12541 2975
rect 12575 2941 12587 2975
rect 13372 2972 13400 3012
rect 13538 3000 13544 3012
rect 13596 3000 13602 3052
rect 13814 3040 13820 3052
rect 13775 3012 13820 3040
rect 13814 3000 13820 3012
rect 13872 3000 13878 3052
rect 14936 2972 14964 3080
rect 16114 3068 16120 3080
rect 16172 3068 16178 3120
rect 19168 3108 19196 3148
rect 23842 3136 23848 3148
rect 23900 3136 23906 3188
rect 26050 3136 26056 3188
rect 26108 3176 26114 3188
rect 27706 3176 27712 3188
rect 26108 3148 27712 3176
rect 26108 3136 26114 3148
rect 27706 3136 27712 3148
rect 27764 3136 27770 3188
rect 27798 3136 27804 3188
rect 27856 3176 27862 3188
rect 28445 3179 28503 3185
rect 28445 3176 28457 3179
rect 27856 3148 28457 3176
rect 27856 3136 27862 3148
rect 28445 3145 28457 3148
rect 28491 3176 28503 3179
rect 28718 3176 28724 3188
rect 28491 3148 28724 3176
rect 28491 3145 28503 3148
rect 28445 3139 28503 3145
rect 28718 3136 28724 3148
rect 28776 3136 28782 3188
rect 31386 3176 31392 3188
rect 31347 3148 31392 3176
rect 31386 3136 31392 3148
rect 31444 3136 31450 3188
rect 33689 3179 33747 3185
rect 33689 3145 33701 3179
rect 33735 3176 33747 3179
rect 33962 3176 33968 3188
rect 33735 3148 33968 3176
rect 33735 3145 33747 3148
rect 33689 3139 33747 3145
rect 33962 3136 33968 3148
rect 34020 3176 34026 3188
rect 34020 3148 35940 3176
rect 34020 3136 34026 3148
rect 16224 3080 19196 3108
rect 16224 3049 16252 3080
rect 15657 3043 15715 3049
rect 15657 3009 15669 3043
rect 15703 3040 15715 3043
rect 16209 3043 16267 3049
rect 15703 3012 16160 3040
rect 15703 3009 15715 3012
rect 15657 3003 15715 3009
rect 15672 2972 15700 3003
rect 13372 2944 14964 2972
rect 15028 2944 15700 2972
rect 15749 2975 15807 2981
rect 12529 2935 12587 2941
rect 12544 2904 12572 2935
rect 10520 2876 12572 2904
rect 2590 2796 2596 2848
rect 2648 2836 2654 2848
rect 3237 2839 3295 2845
rect 3237 2836 3249 2839
rect 2648 2808 3249 2836
rect 2648 2796 2654 2808
rect 3237 2805 3249 2808
rect 3283 2805 3295 2839
rect 3237 2799 3295 2805
rect 8757 2839 8815 2845
rect 8757 2805 8769 2839
rect 8803 2836 8815 2839
rect 10520 2836 10548 2876
rect 8803 2808 10548 2836
rect 8803 2805 8815 2808
rect 8757 2799 8815 2805
rect 12434 2796 12440 2848
rect 12492 2836 12498 2848
rect 15028 2836 15056 2944
rect 15749 2941 15761 2975
rect 15795 2941 15807 2975
rect 16132 2972 16160 3012
rect 16209 3009 16221 3043
rect 16255 3009 16267 3043
rect 16209 3003 16267 3009
rect 16574 3000 16580 3052
rect 16632 3040 16638 3052
rect 16632 3012 16804 3040
rect 16632 3000 16638 3012
rect 16776 2981 16804 3012
rect 16868 3012 19012 3040
rect 16669 2975 16727 2981
rect 16669 2972 16681 2975
rect 16132 2944 16681 2972
rect 15749 2935 15807 2941
rect 16669 2941 16681 2944
rect 16715 2941 16727 2975
rect 16669 2935 16727 2941
rect 16761 2975 16819 2981
rect 16761 2941 16773 2975
rect 16807 2941 16819 2975
rect 16761 2935 16819 2941
rect 15194 2864 15200 2916
rect 15252 2904 15258 2916
rect 15764 2904 15792 2935
rect 15252 2876 15792 2904
rect 16684 2904 16712 2935
rect 16868 2904 16896 3012
rect 18138 2972 18144 2984
rect 18099 2944 18144 2972
rect 18138 2932 18144 2944
rect 18196 2932 18202 2984
rect 18598 2972 18604 2984
rect 18559 2944 18604 2972
rect 18598 2932 18604 2944
rect 18656 2932 18662 2984
rect 17218 2904 17224 2916
rect 16684 2876 16896 2904
rect 17179 2876 17224 2904
rect 15252 2864 15258 2876
rect 17218 2864 17224 2876
rect 17276 2864 17282 2916
rect 18874 2904 18880 2916
rect 18835 2876 18880 2904
rect 18874 2864 18880 2876
rect 18932 2864 18938 2916
rect 18984 2904 19012 3012
rect 19334 3000 19340 3052
rect 19392 3040 19398 3052
rect 19797 3043 19855 3049
rect 19797 3040 19809 3043
rect 19392 3012 19809 3040
rect 19392 3000 19398 3012
rect 19797 3009 19809 3012
rect 19843 3009 19855 3043
rect 19797 3003 19855 3009
rect 21177 3043 21235 3049
rect 21177 3009 21189 3043
rect 21223 3040 21235 3043
rect 21223 3012 23796 3040
rect 21223 3009 21235 3012
rect 21177 3003 21235 3009
rect 19426 2932 19432 2984
rect 19484 2972 19490 2984
rect 19521 2975 19579 2981
rect 19521 2972 19533 2975
rect 19484 2944 19533 2972
rect 19484 2932 19490 2944
rect 19521 2941 19533 2944
rect 19567 2941 19579 2975
rect 21637 2975 21695 2981
rect 21637 2972 21649 2975
rect 19521 2935 19579 2941
rect 19628 2944 21649 2972
rect 19628 2904 19656 2944
rect 21637 2941 21649 2944
rect 21683 2941 21695 2975
rect 21637 2935 21695 2941
rect 21729 2975 21787 2981
rect 21729 2941 21741 2975
rect 21775 2941 21787 2975
rect 21729 2935 21787 2941
rect 18984 2876 19656 2904
rect 12492 2808 15056 2836
rect 15105 2839 15163 2845
rect 12492 2796 12498 2808
rect 15105 2805 15117 2839
rect 15151 2836 15163 2839
rect 21744 2836 21772 2935
rect 21818 2932 21824 2984
rect 21876 2972 21882 2984
rect 23768 2981 23796 3012
rect 24118 3000 24124 3052
rect 24176 3040 24182 3052
rect 32401 3043 32459 3049
rect 24176 3012 32352 3040
rect 24176 3000 24182 3012
rect 23661 2975 23719 2981
rect 23661 2972 23673 2975
rect 21876 2944 23673 2972
rect 21876 2932 21882 2944
rect 23661 2941 23673 2944
rect 23707 2941 23719 2975
rect 23661 2935 23719 2941
rect 23753 2975 23811 2981
rect 23753 2941 23765 2975
rect 23799 2941 23811 2975
rect 23753 2935 23811 2941
rect 24026 2932 24032 2984
rect 24084 2972 24090 2984
rect 24762 2972 24768 2984
rect 24084 2944 24768 2972
rect 24084 2932 24090 2944
rect 24762 2932 24768 2944
rect 24820 2972 24826 2984
rect 24949 2975 25007 2981
rect 24949 2972 24961 2975
rect 24820 2944 24961 2972
rect 24820 2932 24826 2944
rect 24949 2941 24961 2944
rect 24995 2941 25007 2975
rect 25225 2975 25283 2981
rect 25225 2972 25237 2975
rect 24949 2935 25007 2941
rect 25056 2944 25237 2972
rect 22189 2907 22247 2913
rect 22189 2873 22201 2907
rect 22235 2873 22247 2907
rect 22189 2867 22247 2873
rect 24213 2907 24271 2913
rect 24213 2873 24225 2907
rect 24259 2904 24271 2907
rect 24302 2904 24308 2916
rect 24259 2876 24308 2904
rect 24259 2873 24271 2876
rect 24213 2867 24271 2873
rect 15151 2808 21772 2836
rect 22204 2836 22232 2867
rect 24302 2864 24308 2876
rect 24360 2864 24366 2916
rect 25056 2836 25084 2944
rect 25225 2941 25237 2944
rect 25271 2941 25283 2975
rect 25225 2935 25283 2941
rect 26326 2932 26332 2984
rect 26384 2972 26390 2984
rect 27062 2972 27068 2984
rect 26384 2944 27068 2972
rect 26384 2932 26390 2944
rect 27062 2932 27068 2944
rect 27120 2932 27126 2984
rect 27341 2975 27399 2981
rect 27341 2972 27353 2975
rect 27172 2944 27353 2972
rect 26418 2864 26424 2916
rect 26476 2904 26482 2916
rect 27172 2904 27200 2944
rect 27341 2941 27353 2944
rect 27387 2941 27399 2975
rect 27341 2935 27399 2941
rect 27706 2932 27712 2984
rect 27764 2972 27770 2984
rect 27764 2944 29040 2972
rect 27764 2932 27770 2944
rect 26476 2876 27200 2904
rect 29012 2904 29040 2944
rect 29086 2932 29092 2984
rect 29144 2972 29150 2984
rect 30009 2975 30067 2981
rect 30009 2972 30021 2975
rect 29144 2944 30021 2972
rect 29144 2932 29150 2944
rect 30009 2941 30021 2944
rect 30055 2941 30067 2975
rect 30009 2935 30067 2941
rect 30285 2975 30343 2981
rect 30285 2941 30297 2975
rect 30331 2972 30343 2975
rect 32030 2972 32036 2984
rect 30331 2944 32036 2972
rect 30331 2941 30343 2944
rect 30285 2935 30343 2941
rect 32030 2932 32036 2944
rect 32088 2932 32094 2984
rect 32125 2975 32183 2981
rect 32125 2941 32137 2975
rect 32171 2941 32183 2975
rect 32324 2972 32352 3012
rect 32401 3009 32413 3043
rect 32447 3040 32459 3043
rect 33594 3040 33600 3052
rect 32447 3012 33600 3040
rect 32447 3009 32459 3012
rect 32401 3003 32459 3009
rect 33594 3000 33600 3012
rect 33652 3000 33658 3052
rect 34514 3000 34520 3052
rect 34572 3040 34578 3052
rect 34885 3043 34943 3049
rect 34885 3040 34897 3043
rect 34572 3012 34897 3040
rect 34572 3000 34578 3012
rect 34885 3009 34897 3012
rect 34931 3009 34943 3043
rect 35434 3040 35440 3052
rect 35395 3012 35440 3040
rect 34885 3003 34943 3009
rect 35434 3000 35440 3012
rect 35492 3000 35498 3052
rect 35912 3049 35940 3148
rect 35897 3043 35955 3049
rect 35897 3009 35909 3043
rect 35943 3009 35955 3043
rect 35897 3003 35955 3009
rect 32324 2944 33088 2972
rect 32125 2935 32183 2941
rect 30098 2904 30104 2916
rect 29012 2876 30104 2904
rect 26476 2864 26482 2876
rect 30098 2864 30104 2876
rect 30156 2864 30162 2916
rect 22204 2808 25084 2836
rect 26513 2839 26571 2845
rect 15151 2805 15163 2808
rect 15105 2799 15163 2805
rect 26513 2805 26525 2839
rect 26559 2836 26571 2839
rect 27982 2836 27988 2848
rect 26559 2808 27988 2836
rect 26559 2805 26571 2808
rect 26513 2799 26571 2805
rect 27982 2796 27988 2808
rect 28040 2796 28046 2848
rect 30282 2796 30288 2848
rect 30340 2836 30346 2848
rect 32030 2836 32036 2848
rect 30340 2808 32036 2836
rect 30340 2796 30346 2808
rect 32030 2796 32036 2808
rect 32088 2796 32094 2848
rect 32140 2836 32168 2935
rect 33060 2904 33088 2944
rect 33134 2932 33140 2984
rect 33192 2972 33198 2984
rect 35452 2972 35480 3000
rect 35710 2972 35716 2984
rect 33192 2944 35480 2972
rect 35671 2944 35716 2972
rect 33192 2932 33198 2944
rect 35710 2932 35716 2944
rect 35768 2932 35774 2984
rect 36354 2904 36360 2916
rect 33060 2876 36360 2904
rect 36354 2864 36360 2876
rect 36412 2864 36418 2916
rect 33502 2836 33508 2848
rect 32140 2808 33508 2836
rect 33502 2796 33508 2808
rect 33560 2796 33566 2848
rect 1104 2746 39836 2768
rect 1104 2694 19606 2746
rect 19658 2694 19670 2746
rect 19722 2694 19734 2746
rect 19786 2694 19798 2746
rect 19850 2694 39836 2746
rect 1104 2672 39836 2694
rect 8570 2592 8576 2644
rect 8628 2632 8634 2644
rect 9125 2635 9183 2641
rect 9125 2632 9137 2635
rect 8628 2604 9137 2632
rect 8628 2592 8634 2604
rect 9125 2601 9137 2604
rect 9171 2601 9183 2635
rect 9125 2595 9183 2601
rect 16482 2592 16488 2644
rect 16540 2632 16546 2644
rect 18417 2635 18475 2641
rect 18417 2632 18429 2635
rect 16540 2604 18429 2632
rect 16540 2592 16546 2604
rect 18417 2601 18429 2604
rect 18463 2632 18475 2635
rect 18598 2632 18604 2644
rect 18463 2604 18604 2632
rect 18463 2601 18475 2604
rect 18417 2595 18475 2601
rect 18598 2592 18604 2604
rect 18656 2592 18662 2644
rect 19978 2592 19984 2644
rect 20036 2632 20042 2644
rect 24026 2632 24032 2644
rect 20036 2604 24032 2632
rect 20036 2592 20042 2604
rect 24026 2592 24032 2604
rect 24084 2592 24090 2644
rect 28445 2635 28503 2641
rect 28445 2601 28457 2635
rect 28491 2632 28503 2635
rect 30282 2632 30288 2644
rect 28491 2604 30288 2632
rect 28491 2601 28503 2604
rect 28445 2595 28503 2601
rect 30282 2592 30288 2604
rect 30340 2592 30346 2644
rect 14921 2567 14979 2573
rect 14921 2533 14933 2567
rect 14967 2564 14979 2567
rect 15194 2564 15200 2576
rect 14967 2536 15200 2564
rect 14967 2533 14979 2536
rect 14921 2527 14979 2533
rect 15194 2524 15200 2536
rect 15252 2524 15258 2576
rect 3694 2456 3700 2508
rect 3752 2496 3758 2508
rect 4065 2499 4123 2505
rect 4065 2496 4077 2499
rect 3752 2468 4077 2496
rect 3752 2456 3758 2468
rect 4065 2465 4077 2468
rect 4111 2465 4123 2499
rect 4065 2459 4123 2465
rect 4341 2499 4399 2505
rect 4341 2465 4353 2499
rect 4387 2496 4399 2499
rect 4982 2496 4988 2508
rect 4387 2468 4988 2496
rect 4387 2465 4399 2468
rect 4341 2459 4399 2465
rect 4982 2456 4988 2468
rect 5040 2456 5046 2508
rect 6914 2456 6920 2508
rect 6972 2496 6978 2508
rect 6972 2468 7017 2496
rect 6972 2456 6978 2468
rect 8846 2456 8852 2508
rect 8904 2496 8910 2508
rect 9033 2499 9091 2505
rect 9033 2496 9045 2499
rect 8904 2468 9045 2496
rect 8904 2456 8910 2468
rect 9033 2465 9045 2468
rect 9079 2465 9091 2499
rect 10410 2496 10416 2508
rect 10371 2468 10416 2496
rect 9033 2459 9091 2465
rect 10410 2456 10416 2468
rect 10468 2456 10474 2508
rect 10689 2499 10747 2505
rect 10689 2465 10701 2499
rect 10735 2496 10747 2499
rect 11054 2496 11060 2508
rect 10735 2468 11060 2496
rect 10735 2465 10747 2468
rect 10689 2459 10747 2465
rect 11054 2456 11060 2468
rect 11112 2456 11118 2508
rect 13541 2499 13599 2505
rect 13541 2465 13553 2499
rect 13587 2496 13599 2499
rect 14274 2496 14280 2508
rect 13587 2468 14280 2496
rect 13587 2465 13599 2468
rect 13541 2459 13599 2465
rect 14274 2456 14280 2468
rect 14332 2456 14338 2508
rect 15841 2499 15899 2505
rect 15841 2465 15853 2499
rect 15887 2496 15899 2499
rect 17218 2496 17224 2508
rect 15887 2468 17224 2496
rect 15887 2465 15899 2468
rect 15841 2459 15899 2465
rect 17218 2456 17224 2468
rect 17276 2456 17282 2508
rect 18322 2496 18328 2508
rect 18283 2468 18328 2496
rect 18322 2456 18328 2468
rect 18380 2456 18386 2508
rect 18874 2456 18880 2508
rect 18932 2496 18938 2508
rect 19245 2499 19303 2505
rect 19245 2496 19257 2499
rect 18932 2468 19257 2496
rect 18932 2456 18938 2468
rect 19245 2465 19257 2468
rect 19291 2465 19303 2499
rect 19245 2459 19303 2465
rect 19518 2456 19524 2508
rect 19576 2496 19582 2508
rect 19996 2496 20024 2592
rect 20625 2567 20683 2573
rect 20625 2533 20637 2567
rect 20671 2564 20683 2567
rect 21358 2564 21364 2576
rect 20671 2536 21364 2564
rect 20671 2533 20683 2536
rect 20625 2527 20683 2533
rect 21358 2524 21364 2536
rect 21416 2524 21422 2576
rect 19576 2468 20024 2496
rect 19576 2456 19582 2468
rect 22094 2456 22100 2508
rect 22152 2496 22158 2508
rect 24044 2505 24072 2592
rect 26602 2524 26608 2576
rect 26660 2564 26666 2576
rect 26660 2536 27016 2564
rect 26660 2524 26666 2536
rect 24029 2499 24087 2505
rect 22152 2468 22197 2496
rect 22152 2456 22158 2468
rect 24029 2465 24041 2499
rect 24075 2465 24087 2499
rect 24302 2496 24308 2508
rect 24263 2468 24308 2496
rect 24029 2459 24087 2465
rect 24302 2456 24308 2468
rect 24360 2456 24366 2508
rect 26878 2496 26884 2508
rect 26839 2468 26884 2496
rect 26878 2456 26884 2468
rect 26936 2456 26942 2508
rect 26988 2496 27016 2536
rect 29454 2524 29460 2576
rect 29512 2564 29518 2576
rect 32585 2567 32643 2573
rect 29512 2536 30328 2564
rect 29512 2524 29518 2536
rect 28997 2499 29055 2505
rect 26988 2468 28212 2496
rect 5718 2388 5724 2440
rect 5776 2428 5782 2440
rect 7193 2431 7251 2437
rect 7193 2428 7205 2431
rect 5776 2400 7205 2428
rect 5776 2388 5782 2400
rect 7193 2397 7205 2400
rect 7239 2397 7251 2431
rect 7193 2391 7251 2397
rect 13265 2431 13323 2437
rect 13265 2397 13277 2431
rect 13311 2428 13323 2431
rect 15565 2431 15623 2437
rect 15565 2428 15577 2431
rect 13311 2400 15577 2428
rect 13311 2397 13323 2400
rect 13265 2391 13323 2397
rect 15565 2397 15577 2400
rect 15611 2428 15623 2431
rect 18046 2428 18052 2440
rect 15611 2400 18052 2428
rect 15611 2397 15623 2400
rect 15565 2391 15623 2397
rect 18046 2388 18052 2400
rect 18104 2388 18110 2440
rect 18969 2431 19027 2437
rect 18969 2397 18981 2431
rect 19015 2428 19027 2431
rect 19536 2428 19564 2456
rect 19015 2400 19564 2428
rect 21821 2431 21879 2437
rect 19015 2397 19027 2400
rect 18969 2391 19027 2397
rect 21821 2397 21833 2431
rect 21867 2428 21879 2431
rect 22554 2428 22560 2440
rect 21867 2400 22560 2428
rect 21867 2397 21879 2400
rect 21821 2391 21879 2397
rect 22554 2388 22560 2400
rect 22612 2388 22618 2440
rect 26694 2388 26700 2440
rect 26752 2428 26758 2440
rect 27157 2431 27215 2437
rect 27157 2428 27169 2431
rect 26752 2400 27169 2428
rect 26752 2388 26758 2400
rect 27157 2397 27169 2400
rect 27203 2397 27215 2431
rect 28184 2428 28212 2468
rect 28997 2465 29009 2499
rect 29043 2496 29055 2499
rect 30006 2496 30012 2508
rect 29043 2468 30012 2496
rect 29043 2465 29055 2468
rect 28997 2459 29055 2465
rect 30006 2456 30012 2468
rect 30064 2456 30070 2508
rect 30300 2505 30328 2536
rect 32585 2533 32597 2567
rect 32631 2564 32643 2567
rect 33870 2564 33876 2576
rect 32631 2536 33876 2564
rect 32631 2533 32643 2536
rect 32585 2527 32643 2533
rect 33870 2524 33876 2536
rect 33928 2524 33934 2576
rect 30285 2499 30343 2505
rect 30285 2465 30297 2499
rect 30331 2465 30343 2499
rect 30558 2496 30564 2508
rect 30519 2468 30564 2496
rect 30285 2459 30343 2465
rect 30558 2456 30564 2468
rect 30616 2456 30622 2508
rect 31386 2456 31392 2508
rect 31444 2496 31450 2508
rect 33410 2496 33416 2508
rect 31444 2468 33272 2496
rect 33371 2468 33416 2496
rect 31444 2456 31450 2468
rect 29733 2431 29791 2437
rect 29733 2428 29745 2431
rect 28184 2400 29745 2428
rect 27157 2391 27215 2397
rect 29733 2397 29745 2400
rect 29779 2397 29791 2431
rect 29733 2391 29791 2397
rect 30745 2431 30803 2437
rect 30745 2397 30757 2431
rect 30791 2397 30803 2431
rect 33134 2428 33140 2440
rect 33095 2400 33140 2428
rect 30745 2391 30803 2397
rect 8481 2363 8539 2369
rect 8481 2329 8493 2363
rect 8527 2360 8539 2363
rect 8527 2332 10456 2360
rect 8527 2329 8539 2332
rect 8481 2323 8539 2329
rect 4706 2252 4712 2304
rect 4764 2292 4770 2304
rect 5445 2295 5503 2301
rect 5445 2292 5457 2295
rect 4764 2264 5457 2292
rect 4764 2252 4770 2264
rect 5445 2261 5457 2264
rect 5491 2261 5503 2295
rect 10428 2292 10456 2332
rect 28718 2320 28724 2372
rect 28776 2360 28782 2372
rect 30760 2360 30788 2391
rect 33134 2388 33140 2400
rect 33192 2388 33198 2440
rect 33244 2428 33272 2468
rect 33410 2456 33416 2468
rect 33468 2456 33474 2508
rect 33597 2431 33655 2437
rect 33597 2428 33609 2431
rect 33244 2400 33609 2428
rect 33597 2397 33609 2400
rect 33643 2397 33655 2431
rect 33597 2391 33655 2397
rect 28776 2332 30788 2360
rect 28776 2320 28782 2332
rect 11054 2292 11060 2304
rect 10428 2264 11060 2292
rect 5445 2255 5503 2261
rect 11054 2252 11060 2264
rect 11112 2252 11118 2304
rect 11977 2295 12035 2301
rect 11977 2261 11989 2295
rect 12023 2292 12035 2295
rect 13078 2292 13084 2304
rect 12023 2264 13084 2292
rect 12023 2261 12035 2264
rect 11977 2255 12035 2261
rect 13078 2252 13084 2264
rect 13136 2252 13142 2304
rect 17129 2295 17187 2301
rect 17129 2261 17141 2295
rect 17175 2292 17187 2295
rect 17310 2292 17316 2304
rect 17175 2264 17316 2292
rect 17175 2261 17187 2264
rect 17129 2255 17187 2261
rect 17310 2252 17316 2264
rect 17368 2252 17374 2304
rect 23382 2292 23388 2304
rect 23343 2264 23388 2292
rect 23382 2252 23388 2264
rect 23440 2252 23446 2304
rect 25590 2292 25596 2304
rect 25551 2264 25596 2292
rect 25590 2252 25596 2264
rect 25648 2252 25654 2304
rect 38470 2292 38476 2304
rect 38431 2264 38476 2292
rect 38470 2252 38476 2264
rect 38528 2252 38534 2304
rect 1104 2202 39836 2224
rect 1104 2150 4246 2202
rect 4298 2150 4310 2202
rect 4362 2150 4374 2202
rect 4426 2150 4438 2202
rect 4490 2150 34966 2202
rect 35018 2150 35030 2202
rect 35082 2150 35094 2202
rect 35146 2150 35158 2202
rect 35210 2150 39836 2202
rect 1104 2128 39836 2150
rect 19518 2048 19524 2100
rect 19576 2088 19582 2100
rect 20070 2088 20076 2100
rect 19576 2060 20076 2088
rect 19576 2048 19582 2060
rect 20070 2048 20076 2060
rect 20128 2048 20134 2100
rect 23382 2048 23388 2100
rect 23440 2088 23446 2100
rect 34238 2088 34244 2100
rect 23440 2060 34244 2088
rect 23440 2048 23446 2060
rect 34238 2048 34244 2060
rect 34296 2048 34302 2100
rect 25590 1980 25596 2032
rect 25648 2020 25654 2032
rect 36446 2020 36452 2032
rect 25648 1992 36452 2020
rect 25648 1980 25654 1992
rect 36446 1980 36452 1992
rect 36504 1980 36510 2032
rect 19886 1912 19892 1964
rect 19944 1952 19950 1964
rect 25774 1952 25780 1964
rect 19944 1924 25780 1952
rect 19944 1912 19950 1924
rect 25774 1912 25780 1924
rect 25832 1912 25838 1964
rect 566 1776 572 1828
rect 624 1816 630 1828
rect 8754 1816 8760 1828
rect 624 1788 8760 1816
rect 624 1776 630 1788
rect 8754 1776 8760 1788
rect 8812 1776 8818 1828
<< via1 >>
rect 19606 38598 19658 38650
rect 19670 38598 19722 38650
rect 19734 38598 19786 38650
rect 19798 38598 19850 38650
rect 7564 38496 7616 38548
rect 19248 38496 19300 38548
rect 29828 38539 29880 38548
rect 1308 38360 1360 38412
rect 9680 38428 9732 38480
rect 29828 38505 29837 38539
rect 29837 38505 29871 38539
rect 29871 38505 29880 38539
rect 29828 38496 29880 38505
rect 9036 38403 9088 38412
rect 9036 38369 9045 38403
rect 9045 38369 9079 38403
rect 9079 38369 9088 38403
rect 9036 38360 9088 38369
rect 10968 38360 11020 38412
rect 11336 38403 11388 38412
rect 11336 38369 11345 38403
rect 11345 38369 11379 38403
rect 11379 38369 11388 38403
rect 11336 38360 11388 38369
rect 11428 38360 11480 38412
rect 13728 38360 13780 38412
rect 6092 38292 6144 38344
rect 7932 38292 7984 38344
rect 30472 38292 30524 38344
rect 25504 38224 25556 38276
rect 30656 38224 30708 38276
rect 8116 38156 8168 38208
rect 10784 38199 10836 38208
rect 10784 38165 10793 38199
rect 10793 38165 10827 38199
rect 10827 38165 10836 38199
rect 10784 38156 10836 38165
rect 11060 38156 11112 38208
rect 12716 38199 12768 38208
rect 12716 38165 12725 38199
rect 12725 38165 12759 38199
rect 12759 38165 12768 38199
rect 12716 38156 12768 38165
rect 26792 38156 26844 38208
rect 32956 38156 33008 38208
rect 4246 38054 4298 38106
rect 4310 38054 4362 38106
rect 4374 38054 4426 38106
rect 4438 38054 4490 38106
rect 34966 38054 35018 38106
rect 35030 38054 35082 38106
rect 35094 38054 35146 38106
rect 35158 38054 35210 38106
rect 9772 37952 9824 38004
rect 14004 37995 14056 38004
rect 14004 37961 14013 37995
rect 14013 37961 14047 37995
rect 14047 37961 14056 37995
rect 14004 37952 14056 37961
rect 26792 37952 26844 38004
rect 37188 37952 37240 38004
rect 3332 37816 3384 37868
rect 8116 37859 8168 37868
rect 5172 37748 5224 37800
rect 7472 37748 7524 37800
rect 7748 37748 7800 37800
rect 8116 37825 8125 37859
rect 8125 37825 8159 37859
rect 8159 37825 8168 37859
rect 8116 37816 8168 37825
rect 8208 37816 8260 37868
rect 15292 37816 15344 37868
rect 17224 37816 17276 37868
rect 25504 37816 25556 37868
rect 26700 37816 26752 37868
rect 34612 37816 34664 37868
rect 9680 37748 9732 37800
rect 10968 37791 11020 37800
rect 6092 37612 6144 37664
rect 6920 37655 6972 37664
rect 6920 37621 6929 37655
rect 6929 37621 6963 37655
rect 6963 37621 6972 37655
rect 6920 37612 6972 37621
rect 10968 37757 10977 37791
rect 10977 37757 11011 37791
rect 11011 37757 11020 37791
rect 10968 37748 11020 37757
rect 11428 37791 11480 37800
rect 11428 37757 11437 37791
rect 11437 37757 11471 37791
rect 11471 37757 11480 37791
rect 11428 37748 11480 37757
rect 12440 37791 12492 37800
rect 12440 37757 12449 37791
rect 12449 37757 12483 37791
rect 12483 37757 12492 37791
rect 12440 37748 12492 37757
rect 13544 37748 13596 37800
rect 15844 37748 15896 37800
rect 17960 37748 18012 37800
rect 14004 37612 14056 37664
rect 18788 37612 18840 37664
rect 21456 37791 21508 37800
rect 21456 37757 21465 37791
rect 21465 37757 21499 37791
rect 21499 37757 21508 37791
rect 21456 37748 21508 37757
rect 21824 37748 21876 37800
rect 24216 37791 24268 37800
rect 23296 37680 23348 37732
rect 21456 37612 21508 37664
rect 23020 37612 23072 37664
rect 24216 37757 24225 37791
rect 24225 37757 24259 37791
rect 24259 37757 24268 37791
rect 24216 37748 24268 37757
rect 24584 37612 24636 37664
rect 26424 37748 26476 37800
rect 29828 37791 29880 37800
rect 29828 37757 29837 37791
rect 29837 37757 29871 37791
rect 29871 37757 29880 37791
rect 29828 37748 29880 37757
rect 30472 37791 30524 37800
rect 30472 37757 30481 37791
rect 30481 37757 30515 37791
rect 30515 37757 30524 37791
rect 30472 37748 30524 37757
rect 31484 37748 31536 37800
rect 33600 37748 33652 37800
rect 31024 37680 31076 37732
rect 26792 37612 26844 37664
rect 19606 37510 19658 37562
rect 19670 37510 19722 37562
rect 19734 37510 19786 37562
rect 19798 37510 19850 37562
rect 17224 37408 17276 37460
rect 1860 37272 1912 37324
rect 5540 37340 5592 37392
rect 9036 37383 9088 37392
rect 8208 37315 8260 37324
rect 8208 37281 8217 37315
rect 8217 37281 8251 37315
rect 8251 37281 8260 37315
rect 8208 37272 8260 37281
rect 9036 37349 9045 37383
rect 9045 37349 9079 37383
rect 9079 37349 9088 37383
rect 9036 37340 9088 37349
rect 8668 37315 8720 37324
rect 8668 37281 8677 37315
rect 8677 37281 8711 37315
rect 8711 37281 8720 37315
rect 8668 37272 8720 37281
rect 9680 37315 9732 37324
rect 9680 37281 9689 37315
rect 9689 37281 9723 37315
rect 9723 37281 9732 37315
rect 9680 37272 9732 37281
rect 11060 37315 11112 37324
rect 11060 37281 11069 37315
rect 11069 37281 11103 37315
rect 11103 37281 11112 37315
rect 11060 37272 11112 37281
rect 14004 37340 14056 37392
rect 13728 37315 13780 37324
rect 13728 37281 13737 37315
rect 13737 37281 13771 37315
rect 13771 37281 13780 37315
rect 13728 37272 13780 37281
rect 14096 37315 14148 37324
rect 14096 37281 14105 37315
rect 14105 37281 14139 37315
rect 14139 37281 14148 37315
rect 14096 37272 14148 37281
rect 14372 37315 14424 37324
rect 14372 37281 14381 37315
rect 14381 37281 14415 37315
rect 14415 37281 14424 37315
rect 14372 37272 14424 37281
rect 6092 37204 6144 37256
rect 8484 37204 8536 37256
rect 9220 37204 9272 37256
rect 9864 37204 9916 37256
rect 12440 37204 12492 37256
rect 13912 37204 13964 37256
rect 15752 37272 15804 37324
rect 16028 37315 16080 37324
rect 16028 37281 16037 37315
rect 16037 37281 16071 37315
rect 16071 37281 16080 37315
rect 16028 37272 16080 37281
rect 15384 37204 15436 37256
rect 17960 37408 18012 37460
rect 21824 37408 21876 37460
rect 17500 37315 17552 37324
rect 17500 37281 17509 37315
rect 17509 37281 17543 37315
rect 17543 37281 17552 37315
rect 17500 37272 17552 37281
rect 24216 37408 24268 37460
rect 25320 37451 25372 37460
rect 25320 37417 25329 37451
rect 25329 37417 25363 37451
rect 25363 37417 25372 37451
rect 25320 37408 25372 37417
rect 28724 37408 28776 37460
rect 39396 37340 39448 37392
rect 23296 37315 23348 37324
rect 23296 37281 23305 37315
rect 23305 37281 23339 37315
rect 23339 37281 23348 37315
rect 23296 37272 23348 37281
rect 25504 37315 25556 37324
rect 25504 37281 25513 37315
rect 25513 37281 25547 37315
rect 25547 37281 25556 37315
rect 25504 37272 25556 37281
rect 26240 37272 26292 37324
rect 26424 37272 26476 37324
rect 26792 37315 26844 37324
rect 20168 37204 20220 37256
rect 21180 37247 21232 37256
rect 21180 37213 21189 37247
rect 21189 37213 21223 37247
rect 21223 37213 21232 37247
rect 21180 37204 21232 37213
rect 23020 37247 23072 37256
rect 23020 37213 23029 37247
rect 23029 37213 23063 37247
rect 23063 37213 23072 37247
rect 23020 37204 23072 37213
rect 26792 37281 26801 37315
rect 26801 37281 26835 37315
rect 26835 37281 26844 37315
rect 26792 37272 26844 37281
rect 33968 37272 34020 37324
rect 28908 37247 28960 37256
rect 28908 37213 28917 37247
rect 28917 37213 28951 37247
rect 28951 37213 28960 37247
rect 28908 37204 28960 37213
rect 33600 37247 33652 37256
rect 33600 37213 33609 37247
rect 33609 37213 33643 37247
rect 33643 37213 33652 37247
rect 33600 37204 33652 37213
rect 11888 37136 11940 37188
rect 14372 37136 14424 37188
rect 7196 37111 7248 37120
rect 7196 37077 7205 37111
rect 7205 37077 7239 37111
rect 7239 37077 7248 37111
rect 7196 37068 7248 37077
rect 9680 37068 9732 37120
rect 13176 37111 13228 37120
rect 13176 37077 13185 37111
rect 13185 37077 13219 37111
rect 13219 37077 13228 37111
rect 13176 37068 13228 37077
rect 13728 37068 13780 37120
rect 15016 37068 15068 37120
rect 15200 37068 15252 37120
rect 27712 37068 27764 37120
rect 30012 37111 30064 37120
rect 30012 37077 30021 37111
rect 30021 37077 30055 37111
rect 30055 37077 30064 37111
rect 30012 37068 30064 37077
rect 4246 36966 4298 37018
rect 4310 36966 4362 37018
rect 4374 36966 4426 37018
rect 4438 36966 4490 37018
rect 34966 36966 35018 37018
rect 35030 36966 35082 37018
rect 35094 36966 35146 37018
rect 35158 36966 35210 37018
rect 8668 36907 8720 36916
rect 8668 36873 8677 36907
rect 8677 36873 8711 36907
rect 8711 36873 8720 36907
rect 8668 36864 8720 36873
rect 5632 36796 5684 36848
rect 14372 36864 14424 36916
rect 15844 36907 15896 36916
rect 15844 36873 15853 36907
rect 15853 36873 15887 36907
rect 15887 36873 15896 36907
rect 15844 36864 15896 36873
rect 20352 36864 20404 36916
rect 9220 36796 9272 36848
rect 5540 36771 5592 36780
rect 5540 36737 5549 36771
rect 5549 36737 5583 36771
rect 5583 36737 5592 36771
rect 5540 36728 5592 36737
rect 8484 36728 8536 36780
rect 6920 36660 6972 36712
rect 7196 36703 7248 36712
rect 7196 36669 7205 36703
rect 7205 36669 7239 36703
rect 7239 36669 7248 36703
rect 7196 36660 7248 36669
rect 8576 36660 8628 36712
rect 9680 36728 9732 36780
rect 10048 36703 10100 36712
rect 5816 36592 5868 36644
rect 8116 36592 8168 36644
rect 10048 36669 10057 36703
rect 10057 36669 10091 36703
rect 10091 36669 10100 36703
rect 10048 36660 10100 36669
rect 22468 36796 22520 36848
rect 24216 36796 24268 36848
rect 24584 36839 24636 36848
rect 24584 36805 24593 36839
rect 24593 36805 24627 36839
rect 24627 36805 24636 36839
rect 24584 36796 24636 36805
rect 31484 36839 31536 36848
rect 31484 36805 31493 36839
rect 31493 36805 31527 36839
rect 31527 36805 31536 36839
rect 31484 36796 31536 36805
rect 33692 36796 33744 36848
rect 11336 36728 11388 36780
rect 10784 36703 10836 36712
rect 10784 36669 10793 36703
rect 10793 36669 10827 36703
rect 10827 36669 10836 36703
rect 10784 36660 10836 36669
rect 11888 36660 11940 36712
rect 13728 36660 13780 36712
rect 14004 36703 14056 36712
rect 14004 36669 14013 36703
rect 14013 36669 14047 36703
rect 14047 36669 14056 36703
rect 14004 36660 14056 36669
rect 15200 36728 15252 36780
rect 17960 36728 18012 36780
rect 20168 36771 20220 36780
rect 20168 36737 20177 36771
rect 20177 36737 20211 36771
rect 20211 36737 20220 36771
rect 20168 36728 20220 36737
rect 14280 36703 14332 36712
rect 14280 36669 14289 36703
rect 14289 36669 14323 36703
rect 14323 36669 14332 36703
rect 14464 36703 14516 36712
rect 14280 36660 14332 36669
rect 14464 36669 14473 36703
rect 14473 36669 14507 36703
rect 14507 36669 14516 36703
rect 14464 36660 14516 36669
rect 15016 36660 15068 36712
rect 13176 36592 13228 36644
rect 8024 36567 8076 36576
rect 8024 36533 8033 36567
rect 8033 36533 8067 36567
rect 8067 36533 8076 36567
rect 8024 36524 8076 36533
rect 11796 36567 11848 36576
rect 11796 36533 11805 36567
rect 11805 36533 11839 36567
rect 11839 36533 11848 36567
rect 11796 36524 11848 36533
rect 12900 36567 12952 36576
rect 12900 36533 12909 36567
rect 12909 36533 12943 36567
rect 12943 36533 12952 36567
rect 12900 36524 12952 36533
rect 18144 36660 18196 36712
rect 15936 36592 15988 36644
rect 20076 36592 20128 36644
rect 15752 36524 15804 36576
rect 24492 36728 24544 36780
rect 25504 36728 25556 36780
rect 26424 36728 26476 36780
rect 20444 36703 20496 36712
rect 20444 36669 20453 36703
rect 20453 36669 20487 36703
rect 20487 36669 20496 36703
rect 20444 36660 20496 36669
rect 20536 36660 20588 36712
rect 22468 36703 22520 36712
rect 22468 36669 22477 36703
rect 22477 36669 22511 36703
rect 22511 36669 22520 36703
rect 22468 36660 22520 36669
rect 22836 36703 22888 36712
rect 22836 36669 22845 36703
rect 22845 36669 22879 36703
rect 22879 36669 22888 36703
rect 22836 36660 22888 36669
rect 24676 36660 24728 36712
rect 25320 36703 25372 36712
rect 25320 36669 25329 36703
rect 25329 36669 25363 36703
rect 25363 36669 25372 36703
rect 25320 36660 25372 36669
rect 26608 36660 26660 36712
rect 27712 36728 27764 36780
rect 28908 36728 28960 36780
rect 30012 36728 30064 36780
rect 35256 36728 35308 36780
rect 31392 36703 31444 36712
rect 20904 36524 20956 36576
rect 21180 36524 21232 36576
rect 22376 36567 22428 36576
rect 22376 36533 22385 36567
rect 22385 36533 22419 36567
rect 22419 36533 22428 36567
rect 22376 36524 22428 36533
rect 25228 36567 25280 36576
rect 25228 36533 25237 36567
rect 25237 36533 25271 36567
rect 25271 36533 25280 36567
rect 25228 36524 25280 36533
rect 31392 36669 31401 36703
rect 31401 36669 31435 36703
rect 31435 36669 31444 36703
rect 31392 36660 31444 36669
rect 30012 36524 30064 36576
rect 19606 36422 19658 36474
rect 19670 36422 19722 36474
rect 19734 36422 19786 36474
rect 19798 36422 19850 36474
rect 7472 36363 7524 36372
rect 7472 36329 7481 36363
rect 7481 36329 7515 36363
rect 7515 36329 7524 36363
rect 7472 36320 7524 36329
rect 7840 36320 7892 36372
rect 5724 36252 5776 36304
rect 7196 36252 7248 36304
rect 12900 36320 12952 36372
rect 25504 36363 25556 36372
rect 25504 36329 25513 36363
rect 25513 36329 25547 36363
rect 25547 36329 25556 36363
rect 25504 36320 25556 36329
rect 5540 36184 5592 36236
rect 6736 36227 6788 36236
rect 6736 36193 6745 36227
rect 6745 36193 6779 36227
rect 6779 36193 6788 36227
rect 6736 36184 6788 36193
rect 7380 36227 7432 36236
rect 7380 36193 7389 36227
rect 7389 36193 7423 36227
rect 7423 36193 7432 36227
rect 7380 36184 7432 36193
rect 8576 36184 8628 36236
rect 9404 36184 9456 36236
rect 10324 36227 10376 36236
rect 10324 36193 10333 36227
rect 10333 36193 10367 36227
rect 10367 36193 10376 36227
rect 10324 36184 10376 36193
rect 7472 36159 7524 36168
rect 4988 36048 5040 36100
rect 5356 36048 5408 36100
rect 7472 36125 7481 36159
rect 7481 36125 7515 36159
rect 7515 36125 7524 36159
rect 7472 36116 7524 36125
rect 10784 36184 10836 36236
rect 11796 36227 11848 36236
rect 11796 36193 11805 36227
rect 11805 36193 11839 36227
rect 11839 36193 11848 36227
rect 11796 36184 11848 36193
rect 12716 36252 12768 36304
rect 14096 36252 14148 36304
rect 20444 36252 20496 36304
rect 12532 36227 12584 36236
rect 12532 36193 12541 36227
rect 12541 36193 12575 36227
rect 12575 36193 12584 36227
rect 12532 36184 12584 36193
rect 13728 36227 13780 36236
rect 13728 36193 13737 36227
rect 13737 36193 13771 36227
rect 13771 36193 13780 36227
rect 13728 36184 13780 36193
rect 13912 36227 13964 36236
rect 13912 36193 13921 36227
rect 13921 36193 13955 36227
rect 13955 36193 13964 36227
rect 13912 36184 13964 36193
rect 14280 36184 14332 36236
rect 17960 36184 18012 36236
rect 18696 36227 18748 36236
rect 18696 36193 18705 36227
rect 18705 36193 18739 36227
rect 18739 36193 18748 36227
rect 18696 36184 18748 36193
rect 20904 36227 20956 36236
rect 20904 36193 20913 36227
rect 20913 36193 20947 36227
rect 20947 36193 20956 36227
rect 20904 36184 20956 36193
rect 22652 36227 22704 36236
rect 22652 36193 22661 36227
rect 22661 36193 22695 36227
rect 22695 36193 22704 36227
rect 22652 36184 22704 36193
rect 23112 36227 23164 36236
rect 23112 36193 23121 36227
rect 23121 36193 23155 36227
rect 23155 36193 23164 36227
rect 23112 36184 23164 36193
rect 30012 36227 30064 36236
rect 30012 36193 30021 36227
rect 30021 36193 30055 36227
rect 30055 36193 30064 36227
rect 30012 36184 30064 36193
rect 32128 36227 32180 36236
rect 32128 36193 32137 36227
rect 32137 36193 32171 36227
rect 32171 36193 32180 36227
rect 32128 36184 32180 36193
rect 33600 36184 33652 36236
rect 11244 36116 11296 36168
rect 16672 36159 16724 36168
rect 10048 36048 10100 36100
rect 13820 36048 13872 36100
rect 15292 36048 15344 36100
rect 16672 36125 16681 36159
rect 16681 36125 16715 36159
rect 16715 36125 16724 36159
rect 16672 36116 16724 36125
rect 20076 36116 20128 36168
rect 24124 36159 24176 36168
rect 24124 36125 24133 36159
rect 24133 36125 24167 36159
rect 24167 36125 24176 36159
rect 24124 36116 24176 36125
rect 24400 36159 24452 36168
rect 24400 36125 24409 36159
rect 24409 36125 24443 36159
rect 24443 36125 24452 36159
rect 24400 36116 24452 36125
rect 26332 36116 26384 36168
rect 29644 36116 29696 36168
rect 29736 36159 29788 36168
rect 29736 36125 29745 36159
rect 29745 36125 29779 36159
rect 29779 36125 29788 36159
rect 32404 36159 32456 36168
rect 29736 36116 29788 36125
rect 32404 36125 32413 36159
rect 32413 36125 32447 36159
rect 32447 36125 32456 36159
rect 32404 36116 32456 36125
rect 34520 36159 34572 36168
rect 34520 36125 34529 36159
rect 34529 36125 34563 36159
rect 34563 36125 34572 36159
rect 34520 36116 34572 36125
rect 22836 36048 22888 36100
rect 9036 36023 9088 36032
rect 9036 35989 9045 36023
rect 9045 35989 9079 36023
rect 9079 35989 9088 36023
rect 9036 35980 9088 35989
rect 18144 35980 18196 36032
rect 18236 35980 18288 36032
rect 20812 35980 20864 36032
rect 20996 36023 21048 36032
rect 20996 35989 21005 36023
rect 21005 35989 21039 36023
rect 21039 35989 21048 36023
rect 20996 35980 21048 35989
rect 27344 35980 27396 36032
rect 31116 36023 31168 36032
rect 31116 35989 31125 36023
rect 31125 35989 31159 36023
rect 31159 35989 31168 36023
rect 31116 35980 31168 35989
rect 33508 36023 33560 36032
rect 33508 35989 33517 36023
rect 33517 35989 33551 36023
rect 33551 35989 33560 36023
rect 33508 35980 33560 35989
rect 35624 36023 35676 36032
rect 35624 35989 35633 36023
rect 35633 35989 35667 36023
rect 35667 35989 35676 36023
rect 35624 35980 35676 35989
rect 4246 35878 4298 35930
rect 4310 35878 4362 35930
rect 4374 35878 4426 35930
rect 4438 35878 4490 35930
rect 34966 35878 35018 35930
rect 35030 35878 35082 35930
rect 35094 35878 35146 35930
rect 35158 35878 35210 35930
rect 9404 35819 9456 35828
rect 9404 35785 9413 35819
rect 9413 35785 9447 35819
rect 9447 35785 9456 35819
rect 9404 35776 9456 35785
rect 15752 35776 15804 35828
rect 16672 35819 16724 35828
rect 16672 35785 16681 35819
rect 16681 35785 16715 35819
rect 16715 35785 16724 35819
rect 16672 35776 16724 35785
rect 18052 35776 18104 35828
rect 18696 35776 18748 35828
rect 22468 35776 22520 35828
rect 22652 35819 22704 35828
rect 22652 35785 22661 35819
rect 22661 35785 22695 35819
rect 22695 35785 22704 35819
rect 22652 35776 22704 35785
rect 5816 35751 5868 35760
rect 5816 35717 5825 35751
rect 5825 35717 5859 35751
rect 5859 35717 5868 35751
rect 5816 35708 5868 35717
rect 10968 35708 11020 35760
rect 5540 35640 5592 35692
rect 3792 35615 3844 35624
rect 3792 35581 3801 35615
rect 3801 35581 3835 35615
rect 3835 35581 3844 35615
rect 3792 35572 3844 35581
rect 4160 35572 4212 35624
rect 5356 35615 5408 35624
rect 5356 35581 5365 35615
rect 5365 35581 5399 35615
rect 5399 35581 5408 35615
rect 5356 35572 5408 35581
rect 7472 35640 7524 35692
rect 7748 35640 7800 35692
rect 9864 35640 9916 35692
rect 11244 35683 11296 35692
rect 11244 35649 11253 35683
rect 11253 35649 11287 35683
rect 11287 35649 11296 35683
rect 11244 35640 11296 35649
rect 13912 35708 13964 35760
rect 24400 35751 24452 35760
rect 12532 35640 12584 35692
rect 14924 35640 14976 35692
rect 6828 35615 6880 35624
rect 6828 35581 6837 35615
rect 6837 35581 6871 35615
rect 6871 35581 6880 35615
rect 6828 35572 6880 35581
rect 8300 35615 8352 35624
rect 8300 35581 8309 35615
rect 8309 35581 8343 35615
rect 8343 35581 8352 35615
rect 8300 35572 8352 35581
rect 10784 35572 10836 35624
rect 11612 35572 11664 35624
rect 12440 35615 12492 35624
rect 12440 35581 12449 35615
rect 12449 35581 12483 35615
rect 12483 35581 12492 35615
rect 12440 35572 12492 35581
rect 12900 35572 12952 35624
rect 14372 35615 14424 35624
rect 14372 35581 14381 35615
rect 14381 35581 14415 35615
rect 14415 35581 14424 35615
rect 15292 35615 15344 35624
rect 14372 35572 14424 35581
rect 15292 35581 15301 35615
rect 15301 35581 15335 35615
rect 15335 35581 15344 35615
rect 15292 35572 15344 35581
rect 16028 35640 16080 35692
rect 19248 35615 19300 35624
rect 14832 35547 14884 35556
rect 14832 35513 14841 35547
rect 14841 35513 14875 35547
rect 14875 35513 14884 35547
rect 14832 35504 14884 35513
rect 19248 35581 19257 35615
rect 19257 35581 19291 35615
rect 19291 35581 19300 35615
rect 19248 35572 19300 35581
rect 20444 35640 20496 35692
rect 21456 35640 21508 35692
rect 22376 35640 22428 35692
rect 24400 35717 24409 35751
rect 24409 35717 24443 35751
rect 24443 35717 24452 35751
rect 24400 35708 24452 35717
rect 25136 35708 25188 35760
rect 24768 35640 24820 35692
rect 27712 35708 27764 35760
rect 29644 35776 29696 35828
rect 32404 35819 32456 35828
rect 32404 35785 32413 35819
rect 32413 35785 32447 35819
rect 32447 35785 32456 35819
rect 32404 35776 32456 35785
rect 33232 35819 33284 35828
rect 33232 35785 33241 35819
rect 33241 35785 33275 35819
rect 33275 35785 33284 35819
rect 33232 35776 33284 35785
rect 30840 35708 30892 35760
rect 31116 35683 31168 35692
rect 20076 35572 20128 35624
rect 20996 35572 21048 35624
rect 23940 35615 23992 35624
rect 23940 35581 23949 35615
rect 23949 35581 23983 35615
rect 23983 35581 23992 35615
rect 23940 35572 23992 35581
rect 25228 35572 25280 35624
rect 25136 35504 25188 35556
rect 25504 35615 25556 35624
rect 25504 35581 25513 35615
rect 25513 35581 25547 35615
rect 25547 35581 25556 35615
rect 25504 35572 25556 35581
rect 26240 35572 26292 35624
rect 26792 35572 26844 35624
rect 27344 35615 27396 35624
rect 27344 35581 27353 35615
rect 27353 35581 27387 35615
rect 27387 35581 27396 35615
rect 27344 35572 27396 35581
rect 27068 35504 27120 35556
rect 27620 35572 27672 35624
rect 31116 35649 31125 35683
rect 31125 35649 31159 35683
rect 31159 35649 31168 35683
rect 31116 35640 31168 35649
rect 29736 35572 29788 35624
rect 32128 35572 32180 35624
rect 2872 35436 2924 35488
rect 4160 35436 4212 35488
rect 6736 35436 6788 35488
rect 13084 35436 13136 35488
rect 24124 35436 24176 35488
rect 26332 35436 26384 35488
rect 26608 35436 26660 35488
rect 30748 35436 30800 35488
rect 31576 35436 31628 35488
rect 33048 35615 33100 35624
rect 33048 35581 33057 35615
rect 33057 35581 33091 35615
rect 33091 35581 33100 35615
rect 33048 35572 33100 35581
rect 19606 35334 19658 35386
rect 19670 35334 19722 35386
rect 19734 35334 19786 35386
rect 19798 35334 19850 35386
rect 6644 35164 6696 35216
rect 1952 35096 2004 35148
rect 4160 35096 4212 35148
rect 4988 35139 5040 35148
rect 4988 35105 4997 35139
rect 4997 35105 5031 35139
rect 5031 35105 5040 35139
rect 4988 35096 5040 35105
rect 6828 35096 6880 35148
rect 7472 35139 7524 35148
rect 2136 35028 2188 35080
rect 2688 35028 2740 35080
rect 6092 35028 6144 35080
rect 7472 35105 7481 35139
rect 7481 35105 7515 35139
rect 7515 35105 7524 35139
rect 7472 35096 7524 35105
rect 8024 35139 8076 35148
rect 8024 35105 8033 35139
rect 8033 35105 8067 35139
rect 8067 35105 8076 35139
rect 8024 35096 8076 35105
rect 8208 35139 8260 35148
rect 8208 35105 8217 35139
rect 8217 35105 8251 35139
rect 8251 35105 8260 35139
rect 8208 35096 8260 35105
rect 10324 35096 10376 35148
rect 12532 35232 12584 35284
rect 24676 35232 24728 35284
rect 12440 35164 12492 35216
rect 11612 35139 11664 35148
rect 10784 35028 10836 35080
rect 7380 34960 7432 35012
rect 8208 34960 8260 35012
rect 8484 34960 8536 35012
rect 9588 34960 9640 35012
rect 11612 35105 11621 35139
rect 11621 35105 11655 35139
rect 11655 35105 11664 35139
rect 11612 35096 11664 35105
rect 13084 35139 13136 35148
rect 13084 35105 13093 35139
rect 13093 35105 13127 35139
rect 13127 35105 13136 35139
rect 13084 35096 13136 35105
rect 14832 35096 14884 35148
rect 18052 35139 18104 35148
rect 18052 35105 18061 35139
rect 18061 35105 18095 35139
rect 18095 35105 18104 35139
rect 18052 35096 18104 35105
rect 13176 35028 13228 35080
rect 15752 35028 15804 35080
rect 20904 35028 20956 35080
rect 22100 35071 22152 35080
rect 22100 35037 22109 35071
rect 22109 35037 22143 35071
rect 22143 35037 22152 35071
rect 22100 35028 22152 35037
rect 2780 34935 2832 34944
rect 2780 34901 2789 34935
rect 2789 34901 2823 34935
rect 2823 34901 2832 34935
rect 2780 34892 2832 34901
rect 5632 34892 5684 34944
rect 5908 34892 5960 34944
rect 9772 34892 9824 34944
rect 22284 34960 22336 35012
rect 22652 35096 22704 35148
rect 23112 35139 23164 35148
rect 23112 35105 23121 35139
rect 23121 35105 23155 35139
rect 23155 35105 23164 35139
rect 23112 35096 23164 35105
rect 23388 35139 23440 35148
rect 23388 35105 23397 35139
rect 23397 35105 23431 35139
rect 23431 35105 23440 35139
rect 23388 35096 23440 35105
rect 23940 35096 23992 35148
rect 24768 35139 24820 35148
rect 24768 35105 24777 35139
rect 24777 35105 24811 35139
rect 24811 35105 24820 35139
rect 24768 35096 24820 35105
rect 35992 35232 36044 35284
rect 30656 35164 30708 35216
rect 26792 35139 26844 35148
rect 26792 35105 26801 35139
rect 26801 35105 26835 35139
rect 26835 35105 26844 35139
rect 26792 35096 26844 35105
rect 27068 35139 27120 35148
rect 27068 35105 27077 35139
rect 27077 35105 27111 35139
rect 27111 35105 27120 35139
rect 27068 35096 27120 35105
rect 27252 35139 27304 35148
rect 27252 35105 27261 35139
rect 27261 35105 27295 35139
rect 27295 35105 27304 35139
rect 27252 35096 27304 35105
rect 27528 35096 27580 35148
rect 26608 35071 26660 35080
rect 26608 35037 26617 35071
rect 26617 35037 26651 35071
rect 26651 35037 26660 35071
rect 26608 35028 26660 35037
rect 29736 35096 29788 35148
rect 30748 35139 30800 35148
rect 30748 35105 30757 35139
rect 30757 35105 30791 35139
rect 30791 35105 30800 35139
rect 30748 35096 30800 35105
rect 34520 35164 34572 35216
rect 32036 35096 32088 35148
rect 32128 35096 32180 35148
rect 33508 35096 33560 35148
rect 31300 35071 31352 35080
rect 27712 34960 27764 35012
rect 14004 34892 14056 34944
rect 14280 34892 14332 34944
rect 17040 34892 17092 34944
rect 18972 34892 19024 34944
rect 24492 34892 24544 34944
rect 26332 34892 26384 34944
rect 29552 34892 29604 34944
rect 31300 35037 31309 35071
rect 31309 35037 31343 35071
rect 31343 35037 31352 35071
rect 31300 35028 31352 35037
rect 35624 34892 35676 34944
rect 4246 34790 4298 34842
rect 4310 34790 4362 34842
rect 4374 34790 4426 34842
rect 4438 34790 4490 34842
rect 34966 34790 35018 34842
rect 35030 34790 35082 34842
rect 35094 34790 35146 34842
rect 35158 34790 35210 34842
rect 2136 34731 2188 34740
rect 2136 34697 2145 34731
rect 2145 34697 2179 34731
rect 2179 34697 2188 34731
rect 2136 34688 2188 34697
rect 3792 34688 3844 34740
rect 5724 34620 5776 34672
rect 2688 34552 2740 34604
rect 1768 34527 1820 34536
rect 1768 34493 1777 34527
rect 1777 34493 1811 34527
rect 1811 34493 1820 34527
rect 1768 34484 1820 34493
rect 1952 34527 2004 34536
rect 1952 34493 1961 34527
rect 1961 34493 1995 34527
rect 1995 34493 2004 34527
rect 1952 34484 2004 34493
rect 4160 34484 4212 34536
rect 5356 34527 5408 34536
rect 5356 34493 5365 34527
rect 5365 34493 5399 34527
rect 5399 34493 5408 34527
rect 5356 34484 5408 34493
rect 5908 34527 5960 34536
rect 5908 34493 5917 34527
rect 5917 34493 5951 34527
rect 5951 34493 5960 34527
rect 5908 34484 5960 34493
rect 6736 34484 6788 34536
rect 8116 34688 8168 34740
rect 8760 34620 8812 34672
rect 11612 34688 11664 34740
rect 15016 34688 15068 34740
rect 17224 34731 17276 34740
rect 17224 34697 17233 34731
rect 17233 34697 17267 34731
rect 17267 34697 17276 34731
rect 17224 34688 17276 34697
rect 22100 34731 22152 34740
rect 22100 34697 22109 34731
rect 22109 34697 22143 34731
rect 22143 34697 22152 34731
rect 22100 34688 22152 34697
rect 24676 34688 24728 34740
rect 32036 34688 32088 34740
rect 23388 34620 23440 34672
rect 33048 34688 33100 34740
rect 7380 34527 7432 34536
rect 7380 34493 7389 34527
rect 7389 34493 7423 34527
rect 7423 34493 7432 34527
rect 7380 34484 7432 34493
rect 9588 34552 9640 34604
rect 8944 34527 8996 34536
rect 4712 34416 4764 34468
rect 8944 34493 8953 34527
rect 8953 34493 8987 34527
rect 8987 34493 8996 34527
rect 8944 34484 8996 34493
rect 8392 34416 8444 34468
rect 10232 34527 10284 34536
rect 10232 34493 10241 34527
rect 10241 34493 10275 34527
rect 10275 34493 10284 34527
rect 10232 34484 10284 34493
rect 13912 34552 13964 34604
rect 15292 34552 15344 34604
rect 20352 34552 20404 34604
rect 21640 34552 21692 34604
rect 36176 34620 36228 34672
rect 24492 34595 24544 34604
rect 5724 34348 5776 34400
rect 8852 34348 8904 34400
rect 9864 34348 9916 34400
rect 10508 34348 10560 34400
rect 11060 34484 11112 34536
rect 12624 34484 12676 34536
rect 11520 34416 11572 34468
rect 14004 34484 14056 34536
rect 14464 34484 14516 34536
rect 15108 34527 15160 34536
rect 15108 34493 15117 34527
rect 15117 34493 15151 34527
rect 15151 34493 15160 34527
rect 15108 34484 15160 34493
rect 17040 34527 17092 34536
rect 17040 34493 17049 34527
rect 17049 34493 17083 34527
rect 17083 34493 17092 34527
rect 17040 34484 17092 34493
rect 18972 34527 19024 34536
rect 18972 34493 18981 34527
rect 18981 34493 19015 34527
rect 19015 34493 19024 34527
rect 19892 34527 19944 34536
rect 18972 34484 19024 34493
rect 19892 34493 19901 34527
rect 19901 34493 19935 34527
rect 19935 34493 19944 34527
rect 19892 34484 19944 34493
rect 20168 34527 20220 34536
rect 20168 34493 20177 34527
rect 20177 34493 20211 34527
rect 20211 34493 20220 34527
rect 20168 34484 20220 34493
rect 22284 34527 22336 34536
rect 22284 34493 22293 34527
rect 22293 34493 22327 34527
rect 22327 34493 22336 34527
rect 22284 34484 22336 34493
rect 22744 34527 22796 34536
rect 22744 34493 22753 34527
rect 22753 34493 22787 34527
rect 22787 34493 22796 34527
rect 22744 34484 22796 34493
rect 24124 34484 24176 34536
rect 24492 34561 24501 34595
rect 24501 34561 24535 34595
rect 24535 34561 24544 34595
rect 24492 34552 24544 34561
rect 27252 34552 27304 34604
rect 29552 34595 29604 34604
rect 29552 34561 29561 34595
rect 29561 34561 29595 34595
rect 29595 34561 29604 34595
rect 29552 34552 29604 34561
rect 31300 34552 31352 34604
rect 34888 34595 34940 34604
rect 34888 34561 34897 34595
rect 34897 34561 34931 34595
rect 34931 34561 34940 34595
rect 34888 34552 34940 34561
rect 26332 34484 26384 34536
rect 28172 34484 28224 34536
rect 29368 34484 29420 34536
rect 19432 34459 19484 34468
rect 19432 34425 19441 34459
rect 19441 34425 19475 34459
rect 19475 34425 19484 34459
rect 19432 34416 19484 34425
rect 21824 34416 21876 34468
rect 12624 34348 12676 34400
rect 28356 34391 28408 34400
rect 28356 34357 28365 34391
rect 28365 34357 28399 34391
rect 28399 34357 28408 34391
rect 28356 34348 28408 34357
rect 30656 34391 30708 34400
rect 30656 34357 30665 34391
rect 30665 34357 30699 34391
rect 30699 34357 30708 34391
rect 30656 34348 30708 34357
rect 31300 34416 31352 34468
rect 33784 34527 33836 34536
rect 33784 34493 33793 34527
rect 33793 34493 33827 34527
rect 33827 34493 33836 34527
rect 33784 34484 33836 34493
rect 34796 34484 34848 34536
rect 34980 34527 35032 34536
rect 34980 34493 34989 34527
rect 34989 34493 35023 34527
rect 35023 34493 35032 34527
rect 34980 34484 35032 34493
rect 35256 34416 35308 34468
rect 32496 34348 32548 34400
rect 19606 34246 19658 34298
rect 19670 34246 19722 34298
rect 19734 34246 19786 34298
rect 19798 34246 19850 34298
rect 8300 34187 8352 34196
rect 8300 34153 8309 34187
rect 8309 34153 8343 34187
rect 8343 34153 8352 34187
rect 8300 34144 8352 34153
rect 11060 34144 11112 34196
rect 15108 34144 15160 34196
rect 27252 34144 27304 34196
rect 1768 34076 1820 34128
rect 2780 34076 2832 34128
rect 3056 34076 3108 34128
rect 4160 34076 4212 34128
rect 5632 34076 5684 34128
rect 3148 34051 3200 34060
rect 3148 34017 3157 34051
rect 3157 34017 3191 34051
rect 3191 34017 3200 34051
rect 3148 34008 3200 34017
rect 3332 34051 3384 34060
rect 3332 34017 3341 34051
rect 3341 34017 3375 34051
rect 3375 34017 3384 34051
rect 3332 34008 3384 34017
rect 3700 34008 3752 34060
rect 2964 33940 3016 33992
rect 4620 33983 4672 33992
rect 4620 33949 4629 33983
rect 4629 33949 4663 33983
rect 4663 33949 4672 33983
rect 4620 33940 4672 33949
rect 5080 33983 5132 33992
rect 5080 33949 5089 33983
rect 5089 33949 5123 33983
rect 5123 33949 5132 33983
rect 5080 33940 5132 33949
rect 5908 33983 5960 33992
rect 5908 33949 5917 33983
rect 5917 33949 5951 33983
rect 5951 33949 5960 33983
rect 5908 33940 5960 33949
rect 6092 33872 6144 33924
rect 6644 34008 6696 34060
rect 6920 34008 6972 34060
rect 8116 34076 8168 34128
rect 8576 34076 8628 34128
rect 9036 34076 9088 34128
rect 9588 34076 9640 34128
rect 10232 34076 10284 34128
rect 10968 34076 11020 34128
rect 12624 34119 12676 34128
rect 12624 34085 12633 34119
rect 12633 34085 12667 34119
rect 12667 34085 12676 34119
rect 12624 34076 12676 34085
rect 7196 34051 7248 34060
rect 7196 34017 7205 34051
rect 7205 34017 7239 34051
rect 7239 34017 7248 34051
rect 7196 34008 7248 34017
rect 8208 34051 8260 34060
rect 8208 34017 8217 34051
rect 8217 34017 8251 34051
rect 8251 34017 8260 34051
rect 8208 34008 8260 34017
rect 8484 34051 8536 34060
rect 8484 34017 8493 34051
rect 8493 34017 8527 34051
rect 8527 34017 8536 34051
rect 8484 34008 8536 34017
rect 8852 34051 8904 34060
rect 8852 34017 8861 34051
rect 8861 34017 8895 34051
rect 8895 34017 8904 34051
rect 8852 34008 8904 34017
rect 11520 34008 11572 34060
rect 13360 34051 13412 34060
rect 13360 34017 13369 34051
rect 13369 34017 13403 34051
rect 13403 34017 13412 34051
rect 13360 34008 13412 34017
rect 13912 34051 13964 34060
rect 13912 34017 13921 34051
rect 13921 34017 13955 34051
rect 13955 34017 13964 34051
rect 13912 34008 13964 34017
rect 17224 34008 17276 34060
rect 19432 34008 19484 34060
rect 20996 34008 21048 34060
rect 24216 34051 24268 34060
rect 24216 34017 24225 34051
rect 24225 34017 24259 34051
rect 24259 34017 24268 34051
rect 24216 34008 24268 34017
rect 25228 34051 25280 34060
rect 25228 34017 25237 34051
rect 25237 34017 25271 34051
rect 25271 34017 25280 34051
rect 25228 34008 25280 34017
rect 27068 34076 27120 34128
rect 28356 34076 28408 34128
rect 27252 34051 27304 34060
rect 27252 34017 27261 34051
rect 27261 34017 27295 34051
rect 27295 34017 27304 34051
rect 27252 34008 27304 34017
rect 27712 34051 27764 34060
rect 27712 34017 27721 34051
rect 27721 34017 27755 34051
rect 27755 34017 27764 34051
rect 27712 34008 27764 34017
rect 31392 34144 31444 34196
rect 7104 33940 7156 33992
rect 7840 33940 7892 33992
rect 10600 33940 10652 33992
rect 11244 33983 11296 33992
rect 8392 33872 8444 33924
rect 9864 33872 9916 33924
rect 10048 33872 10100 33924
rect 11244 33949 11253 33983
rect 11253 33949 11287 33983
rect 11287 33949 11296 33983
rect 11244 33940 11296 33949
rect 13820 33983 13872 33992
rect 13820 33949 13829 33983
rect 13829 33949 13863 33983
rect 13863 33949 13872 33983
rect 13820 33940 13872 33949
rect 15936 33940 15988 33992
rect 19892 33940 19944 33992
rect 22284 33983 22336 33992
rect 22284 33949 22293 33983
rect 22293 33949 22327 33983
rect 22327 33949 22336 33983
rect 22284 33940 22336 33949
rect 24124 33983 24176 33992
rect 24124 33949 24133 33983
rect 24133 33949 24167 33983
rect 24167 33949 24176 33983
rect 24124 33940 24176 33949
rect 25136 33983 25188 33992
rect 25136 33949 25145 33983
rect 25145 33949 25179 33983
rect 25179 33949 25188 33983
rect 25136 33940 25188 33949
rect 5724 33804 5776 33856
rect 8300 33804 8352 33856
rect 26240 33872 26292 33924
rect 29460 33940 29512 33992
rect 31576 33940 31628 33992
rect 34888 34144 34940 34196
rect 34980 34119 35032 34128
rect 34980 34085 34989 34119
rect 34989 34085 35023 34119
rect 35023 34085 35032 34119
rect 34980 34076 35032 34085
rect 32312 34008 32364 34060
rect 32496 34008 32548 34060
rect 34520 34008 34572 34060
rect 36084 34008 36136 34060
rect 13176 33804 13228 33856
rect 18420 33804 18472 33856
rect 20260 33847 20312 33856
rect 20260 33813 20269 33847
rect 20269 33813 20303 33847
rect 20303 33813 20312 33847
rect 20260 33804 20312 33813
rect 21640 33804 21692 33856
rect 23572 33847 23624 33856
rect 23572 33813 23581 33847
rect 23581 33813 23615 33847
rect 23615 33813 23624 33847
rect 23572 33804 23624 33813
rect 24400 33847 24452 33856
rect 24400 33813 24409 33847
rect 24409 33813 24443 33847
rect 24443 33813 24452 33847
rect 24400 33804 24452 33813
rect 24860 33804 24912 33856
rect 28172 33847 28224 33856
rect 28172 33813 28181 33847
rect 28181 33813 28215 33847
rect 28215 33813 28224 33847
rect 28172 33804 28224 33813
rect 4246 33702 4298 33754
rect 4310 33702 4362 33754
rect 4374 33702 4426 33754
rect 4438 33702 4490 33754
rect 34966 33702 35018 33754
rect 35030 33702 35082 33754
rect 35094 33702 35146 33754
rect 35158 33702 35210 33754
rect 3148 33600 3200 33652
rect 5080 33600 5132 33652
rect 7196 33600 7248 33652
rect 8576 33600 8628 33652
rect 11244 33600 11296 33652
rect 20168 33600 20220 33652
rect 3792 33507 3844 33516
rect 3792 33473 3801 33507
rect 3801 33473 3835 33507
rect 3835 33473 3844 33507
rect 3792 33464 3844 33473
rect 2780 33439 2832 33448
rect 2780 33405 2789 33439
rect 2789 33405 2823 33439
rect 2823 33405 2832 33439
rect 3332 33439 3384 33448
rect 2780 33396 2832 33405
rect 3332 33405 3341 33439
rect 3341 33405 3375 33439
rect 3375 33405 3384 33439
rect 3332 33396 3384 33405
rect 3700 33439 3752 33448
rect 3700 33405 3709 33439
rect 3709 33405 3743 33439
rect 3743 33405 3752 33439
rect 3700 33396 3752 33405
rect 4712 33439 4764 33448
rect 4712 33405 4721 33439
rect 4721 33405 4755 33439
rect 4755 33405 4764 33439
rect 4712 33396 4764 33405
rect 6736 33464 6788 33516
rect 6920 33507 6972 33516
rect 6920 33473 6929 33507
rect 6929 33473 6963 33507
rect 6963 33473 6972 33507
rect 6920 33464 6972 33473
rect 7104 33439 7156 33448
rect 7104 33405 7113 33439
rect 7113 33405 7147 33439
rect 7147 33405 7156 33439
rect 7104 33396 7156 33405
rect 8208 33532 8260 33584
rect 13360 33532 13412 33584
rect 16212 33464 16264 33516
rect 8116 33439 8168 33448
rect 7380 33328 7432 33380
rect 7196 33260 7248 33312
rect 8116 33405 8125 33439
rect 8125 33405 8159 33439
rect 8159 33405 8168 33439
rect 8116 33396 8168 33405
rect 8300 33396 8352 33448
rect 10324 33396 10376 33448
rect 10508 33439 10560 33448
rect 10508 33405 10517 33439
rect 10517 33405 10551 33439
rect 10551 33405 10560 33439
rect 10508 33396 10560 33405
rect 10600 33439 10652 33448
rect 10600 33405 10609 33439
rect 10609 33405 10643 33439
rect 10643 33405 10652 33439
rect 10600 33396 10652 33405
rect 11060 33439 11112 33448
rect 8852 33328 8904 33380
rect 9588 33328 9640 33380
rect 11060 33405 11069 33439
rect 11069 33405 11103 33439
rect 11103 33405 11112 33439
rect 11060 33396 11112 33405
rect 13636 33439 13688 33448
rect 10968 33328 11020 33380
rect 13636 33405 13645 33439
rect 13645 33405 13679 33439
rect 13679 33405 13688 33439
rect 13636 33396 13688 33405
rect 13912 33439 13964 33448
rect 13912 33405 13921 33439
rect 13921 33405 13955 33439
rect 13955 33405 13964 33439
rect 13912 33396 13964 33405
rect 14004 33396 14056 33448
rect 15108 33439 15160 33448
rect 15108 33405 15117 33439
rect 15117 33405 15151 33439
rect 15151 33405 15160 33439
rect 15108 33396 15160 33405
rect 16580 33396 16632 33448
rect 21640 33532 21692 33584
rect 20352 33464 20404 33516
rect 21088 33464 21140 33516
rect 24124 33600 24176 33652
rect 24492 33600 24544 33652
rect 29552 33600 29604 33652
rect 31576 33643 31628 33652
rect 22284 33507 22336 33516
rect 22284 33473 22293 33507
rect 22293 33473 22327 33507
rect 22327 33473 22336 33507
rect 22284 33464 22336 33473
rect 23204 33464 23256 33516
rect 24860 33507 24912 33516
rect 20536 33396 20588 33448
rect 20812 33439 20864 33448
rect 20812 33405 20821 33439
rect 20821 33405 20855 33439
rect 20855 33405 20864 33439
rect 20812 33396 20864 33405
rect 21824 33439 21876 33448
rect 21824 33405 21833 33439
rect 21833 33405 21867 33439
rect 21867 33405 21876 33439
rect 21824 33396 21876 33405
rect 24492 33396 24544 33448
rect 24860 33473 24869 33507
rect 24869 33473 24903 33507
rect 24903 33473 24912 33507
rect 24860 33464 24912 33473
rect 27160 33464 27212 33516
rect 29460 33464 29512 33516
rect 30656 33464 30708 33516
rect 27620 33396 27672 33448
rect 31576 33609 31585 33643
rect 31585 33609 31619 33643
rect 31619 33609 31628 33643
rect 31576 33600 31628 33609
rect 33784 33600 33836 33652
rect 32496 33464 32548 33516
rect 33232 33464 33284 33516
rect 35256 33464 35308 33516
rect 34520 33396 34572 33448
rect 13452 33328 13504 33380
rect 21180 33328 21232 33380
rect 37004 33328 37056 33380
rect 8760 33260 8812 33312
rect 15844 33260 15896 33312
rect 17132 33303 17184 33312
rect 17132 33269 17141 33303
rect 17141 33269 17175 33303
rect 17175 33269 17184 33303
rect 17132 33260 17184 33269
rect 17960 33260 18012 33312
rect 19248 33303 19300 33312
rect 19248 33269 19257 33303
rect 19257 33269 19291 33303
rect 19291 33269 19300 33303
rect 19248 33260 19300 33269
rect 23756 33260 23808 33312
rect 27896 33260 27948 33312
rect 31484 33260 31536 33312
rect 19606 33158 19658 33210
rect 19670 33158 19722 33210
rect 19734 33158 19786 33210
rect 19798 33158 19850 33210
rect 3332 32988 3384 33040
rect 2688 32920 2740 32972
rect 6000 33056 6052 33108
rect 8392 33056 8444 33108
rect 10968 33056 11020 33108
rect 4620 32988 4672 33040
rect 5080 32988 5132 33040
rect 4712 32963 4764 32972
rect 4712 32929 4721 32963
rect 4721 32929 4755 32963
rect 4755 32929 4764 32963
rect 4712 32920 4764 32929
rect 4988 32963 5040 32972
rect 4988 32929 4997 32963
rect 4997 32929 5031 32963
rect 5031 32929 5040 32963
rect 4988 32920 5040 32929
rect 8944 32988 8996 33040
rect 15108 33056 15160 33108
rect 13360 32988 13412 33040
rect 16672 33056 16724 33108
rect 25228 33056 25280 33108
rect 8576 32963 8628 32972
rect 1676 32895 1728 32904
rect 1676 32861 1685 32895
rect 1685 32861 1719 32895
rect 1719 32861 1728 32895
rect 1676 32852 1728 32861
rect 4068 32852 4120 32904
rect 8576 32929 8585 32963
rect 8585 32929 8619 32963
rect 8619 32929 8628 32963
rect 8576 32920 8628 32929
rect 9128 32920 9180 32972
rect 11336 32963 11388 32972
rect 6092 32852 6144 32904
rect 6460 32895 6512 32904
rect 6460 32861 6469 32895
rect 6469 32861 6503 32895
rect 6503 32861 6512 32895
rect 6460 32852 6512 32861
rect 6736 32895 6788 32904
rect 6736 32861 6745 32895
rect 6745 32861 6779 32895
rect 6779 32861 6788 32895
rect 6736 32852 6788 32861
rect 9680 32895 9732 32904
rect 9680 32861 9689 32895
rect 9689 32861 9723 32895
rect 9723 32861 9732 32895
rect 9680 32852 9732 32861
rect 10232 32895 10284 32904
rect 10232 32861 10241 32895
rect 10241 32861 10275 32895
rect 10275 32861 10284 32895
rect 10232 32852 10284 32861
rect 11060 32852 11112 32904
rect 11336 32929 11345 32963
rect 11345 32929 11379 32963
rect 11379 32929 11388 32963
rect 11336 32920 11388 32929
rect 11428 32963 11480 32972
rect 11428 32929 11437 32963
rect 11437 32929 11471 32963
rect 11471 32929 11480 32963
rect 11428 32920 11480 32929
rect 14464 32963 14516 32972
rect 14464 32929 14473 32963
rect 14473 32929 14507 32963
rect 14507 32929 14516 32963
rect 14464 32920 14516 32929
rect 15660 32963 15712 32972
rect 15660 32929 15669 32963
rect 15669 32929 15703 32963
rect 15703 32929 15712 32963
rect 15660 32920 15712 32929
rect 16580 32988 16632 33040
rect 31300 33056 31352 33108
rect 16120 32963 16172 32972
rect 16120 32929 16129 32963
rect 16129 32929 16163 32963
rect 16163 32929 16172 32963
rect 16120 32920 16172 32929
rect 16212 32920 16264 32972
rect 16396 32852 16448 32904
rect 17132 32920 17184 32972
rect 19892 32920 19944 32972
rect 20444 32920 20496 32972
rect 21180 32963 21232 32972
rect 18328 32852 18380 32904
rect 18972 32895 19024 32904
rect 18972 32861 18981 32895
rect 18981 32861 19015 32895
rect 19015 32861 19024 32895
rect 18972 32852 19024 32861
rect 21180 32929 21189 32963
rect 21189 32929 21223 32963
rect 21223 32929 21232 32963
rect 21180 32920 21232 32929
rect 23204 32895 23256 32904
rect 23204 32861 23213 32895
rect 23213 32861 23247 32895
rect 23247 32861 23256 32895
rect 23204 32852 23256 32861
rect 24400 32920 24452 32972
rect 25136 32852 25188 32904
rect 27160 32895 27212 32904
rect 27160 32861 27169 32895
rect 27169 32861 27203 32895
rect 27203 32861 27212 32895
rect 27436 32895 27488 32904
rect 27160 32852 27212 32861
rect 27436 32861 27445 32895
rect 27445 32861 27479 32895
rect 27479 32861 27488 32895
rect 27436 32852 27488 32861
rect 29276 32895 29328 32904
rect 29276 32861 29285 32895
rect 29285 32861 29319 32895
rect 29319 32861 29328 32895
rect 29552 32920 29604 32972
rect 30380 32920 30432 32972
rect 32864 32963 32916 32972
rect 32864 32929 32873 32963
rect 32873 32929 32907 32963
rect 32907 32929 32916 32963
rect 32864 32920 32916 32929
rect 33784 32920 33836 32972
rect 33876 32963 33928 32972
rect 33876 32929 33885 32963
rect 33885 32929 33919 32963
rect 33919 32929 33928 32963
rect 33876 32920 33928 32929
rect 34796 32920 34848 32972
rect 39120 32920 39172 32972
rect 29276 32852 29328 32861
rect 32772 32852 32824 32904
rect 34520 32852 34572 32904
rect 8116 32784 8168 32836
rect 11336 32784 11388 32836
rect 32404 32827 32456 32836
rect 32404 32793 32413 32827
rect 32413 32793 32447 32827
rect 32447 32793 32456 32827
rect 32404 32784 32456 32793
rect 7104 32716 7156 32768
rect 8208 32716 8260 32768
rect 8760 32759 8812 32768
rect 8760 32725 8769 32759
rect 8769 32725 8803 32759
rect 8803 32725 8812 32759
rect 8760 32716 8812 32725
rect 9588 32716 9640 32768
rect 17868 32716 17920 32768
rect 19156 32716 19208 32768
rect 25596 32759 25648 32768
rect 25596 32725 25605 32759
rect 25605 32725 25639 32759
rect 25639 32725 25648 32759
rect 25596 32716 25648 32725
rect 27620 32716 27672 32768
rect 33232 32716 33284 32768
rect 36268 32759 36320 32768
rect 36268 32725 36277 32759
rect 36277 32725 36311 32759
rect 36311 32725 36320 32759
rect 36268 32716 36320 32725
rect 38200 32716 38252 32768
rect 4246 32614 4298 32666
rect 4310 32614 4362 32666
rect 4374 32614 4426 32666
rect 4438 32614 4490 32666
rect 34966 32614 35018 32666
rect 35030 32614 35082 32666
rect 35094 32614 35146 32666
rect 35158 32614 35210 32666
rect 5908 32512 5960 32564
rect 15660 32512 15712 32564
rect 16212 32512 16264 32564
rect 18328 32512 18380 32564
rect 22652 32512 22704 32564
rect 27436 32512 27488 32564
rect 3056 32444 3108 32496
rect 3240 32487 3292 32496
rect 3240 32453 3249 32487
rect 3249 32453 3283 32487
rect 3283 32453 3292 32487
rect 3240 32444 3292 32453
rect 4160 32444 4212 32496
rect 4620 32444 4672 32496
rect 4988 32444 5040 32496
rect 10968 32444 11020 32496
rect 18972 32487 19024 32496
rect 2964 32376 3016 32428
rect 4068 32376 4120 32428
rect 3332 32351 3384 32360
rect 3332 32317 3341 32351
rect 3341 32317 3375 32351
rect 3375 32317 3384 32351
rect 3332 32308 3384 32317
rect 4160 32351 4212 32360
rect 3056 32240 3108 32292
rect 4160 32317 4169 32351
rect 4169 32317 4203 32351
rect 4203 32317 4212 32351
rect 4160 32308 4212 32317
rect 6736 32376 6788 32428
rect 7380 32376 7432 32428
rect 5080 32351 5132 32360
rect 5080 32317 5089 32351
rect 5089 32317 5123 32351
rect 5123 32317 5132 32351
rect 5080 32308 5132 32317
rect 5724 32351 5776 32360
rect 5724 32317 5733 32351
rect 5733 32317 5767 32351
rect 5767 32317 5776 32351
rect 5724 32308 5776 32317
rect 6920 32308 6972 32360
rect 8300 32351 8352 32360
rect 4712 32240 4764 32292
rect 6552 32240 6604 32292
rect 7288 32240 7340 32292
rect 8300 32317 8309 32351
rect 8309 32317 8343 32351
rect 8343 32317 8352 32351
rect 8300 32308 8352 32317
rect 10232 32376 10284 32428
rect 8760 32351 8812 32360
rect 8760 32317 8769 32351
rect 8769 32317 8803 32351
rect 8803 32317 8812 32351
rect 8760 32308 8812 32317
rect 9864 32351 9916 32360
rect 9864 32317 9873 32351
rect 9873 32317 9907 32351
rect 9907 32317 9916 32351
rect 9864 32308 9916 32317
rect 10600 32351 10652 32360
rect 9496 32240 9548 32292
rect 9588 32240 9640 32292
rect 10600 32317 10609 32351
rect 10609 32317 10643 32351
rect 10643 32317 10652 32351
rect 10600 32308 10652 32317
rect 11060 32351 11112 32360
rect 11060 32317 11069 32351
rect 11069 32317 11103 32351
rect 11103 32317 11112 32351
rect 11060 32308 11112 32317
rect 18972 32453 18981 32487
rect 18981 32453 19015 32487
rect 19015 32453 19024 32487
rect 18972 32444 19024 32453
rect 28080 32487 28132 32496
rect 28080 32453 28089 32487
rect 28089 32453 28123 32487
rect 28123 32453 28132 32487
rect 28080 32444 28132 32453
rect 32864 32444 32916 32496
rect 13176 32419 13228 32428
rect 13176 32385 13185 32419
rect 13185 32385 13219 32419
rect 13219 32385 13228 32419
rect 13176 32376 13228 32385
rect 13452 32419 13504 32428
rect 13452 32385 13461 32419
rect 13461 32385 13495 32419
rect 13495 32385 13504 32419
rect 13452 32376 13504 32385
rect 14556 32376 14608 32428
rect 15108 32308 15160 32360
rect 15844 32308 15896 32360
rect 16672 32376 16724 32428
rect 20444 32419 20496 32428
rect 11428 32240 11480 32292
rect 14832 32283 14884 32292
rect 14832 32249 14841 32283
rect 14841 32249 14875 32283
rect 14875 32249 14884 32283
rect 14832 32240 14884 32249
rect 17500 32308 17552 32360
rect 17960 32308 18012 32360
rect 20444 32385 20453 32419
rect 20453 32385 20487 32419
rect 20487 32385 20496 32419
rect 20444 32376 20496 32385
rect 21088 32376 21140 32428
rect 23204 32376 23256 32428
rect 18512 32351 18564 32360
rect 18512 32317 18521 32351
rect 18521 32317 18555 32351
rect 18555 32317 18564 32351
rect 18512 32308 18564 32317
rect 18880 32351 18932 32360
rect 18880 32317 18889 32351
rect 18889 32317 18923 32351
rect 18923 32317 18932 32351
rect 18880 32308 18932 32317
rect 20720 32351 20772 32360
rect 20720 32317 20729 32351
rect 20729 32317 20763 32351
rect 20763 32317 20772 32351
rect 20720 32308 20772 32317
rect 25596 32376 25648 32428
rect 29276 32419 29328 32428
rect 29276 32385 29285 32419
rect 29285 32385 29319 32419
rect 29319 32385 29328 32419
rect 29276 32376 29328 32385
rect 33876 32376 33928 32428
rect 25780 32351 25832 32360
rect 25780 32317 25789 32351
rect 25789 32317 25823 32351
rect 25823 32317 25832 32351
rect 25780 32308 25832 32317
rect 26056 32351 26108 32360
rect 26056 32317 26065 32351
rect 26065 32317 26099 32351
rect 26099 32317 26108 32351
rect 26056 32308 26108 32317
rect 28632 32308 28684 32360
rect 28816 32308 28868 32360
rect 30196 32308 30248 32360
rect 30840 32351 30892 32360
rect 17776 32240 17828 32292
rect 3148 32172 3200 32224
rect 16212 32172 16264 32224
rect 18512 32172 18564 32224
rect 24400 32172 24452 32224
rect 27160 32215 27212 32224
rect 27160 32181 27169 32215
rect 27169 32181 27203 32215
rect 27203 32181 27212 32215
rect 27160 32172 27212 32181
rect 30840 32317 30849 32351
rect 30849 32317 30883 32351
rect 30883 32317 30892 32351
rect 30840 32308 30892 32317
rect 32956 32351 33008 32360
rect 32956 32317 32965 32351
rect 32965 32317 32999 32351
rect 32999 32317 33008 32351
rect 32956 32308 33008 32317
rect 34796 32308 34848 32360
rect 36084 32308 36136 32360
rect 36268 32351 36320 32360
rect 36268 32317 36277 32351
rect 36277 32317 36311 32351
rect 36311 32317 36320 32351
rect 36268 32308 36320 32317
rect 38660 32351 38712 32360
rect 38660 32317 38669 32351
rect 38669 32317 38703 32351
rect 38703 32317 38712 32351
rect 38660 32308 38712 32317
rect 32220 32283 32272 32292
rect 32220 32249 32229 32283
rect 32229 32249 32263 32283
rect 32263 32249 32272 32283
rect 32220 32240 32272 32249
rect 33324 32240 33376 32292
rect 35808 32283 35860 32292
rect 32128 32172 32180 32224
rect 34520 32172 34572 32224
rect 35808 32249 35817 32283
rect 35817 32249 35851 32283
rect 35851 32249 35860 32283
rect 35808 32240 35860 32249
rect 36176 32172 36228 32224
rect 36544 32172 36596 32224
rect 38752 32215 38804 32224
rect 38752 32181 38761 32215
rect 38761 32181 38795 32215
rect 38795 32181 38804 32215
rect 38752 32172 38804 32181
rect 19606 32070 19658 32122
rect 19670 32070 19722 32122
rect 19734 32070 19786 32122
rect 19798 32070 19850 32122
rect 1676 31968 1728 32020
rect 4068 31968 4120 32020
rect 2504 31875 2556 31884
rect 2504 31841 2513 31875
rect 2513 31841 2547 31875
rect 2547 31841 2556 31875
rect 2504 31832 2556 31841
rect 3056 31875 3108 31884
rect 3056 31841 3065 31875
rect 3065 31841 3099 31875
rect 3099 31841 3108 31875
rect 3056 31832 3108 31841
rect 3240 31875 3292 31884
rect 3240 31841 3249 31875
rect 3249 31841 3283 31875
rect 3283 31841 3292 31875
rect 3240 31832 3292 31841
rect 4068 31875 4120 31884
rect 4068 31841 4077 31875
rect 4077 31841 4111 31875
rect 4111 31841 4120 31875
rect 4068 31832 4120 31841
rect 7196 31900 7248 31952
rect 7288 31832 7340 31884
rect 8760 31900 8812 31952
rect 8208 31875 8260 31884
rect 8208 31841 8217 31875
rect 8217 31841 8251 31875
rect 8251 31841 8260 31875
rect 8208 31832 8260 31841
rect 10600 31968 10652 32020
rect 11060 31968 11112 32020
rect 13636 31968 13688 32020
rect 14464 31968 14516 32020
rect 9588 31832 9640 31884
rect 9680 31832 9732 31884
rect 12256 31832 12308 31884
rect 12992 31875 13044 31884
rect 12992 31841 13001 31875
rect 13001 31841 13035 31875
rect 13035 31841 13044 31875
rect 12992 31832 13044 31841
rect 13636 31832 13688 31884
rect 13912 31900 13964 31952
rect 14004 31875 14056 31884
rect 14004 31841 14013 31875
rect 14013 31841 14047 31875
rect 14047 31841 14056 31875
rect 14004 31832 14056 31841
rect 15200 31832 15252 31884
rect 15844 31832 15896 31884
rect 16120 31900 16172 31952
rect 16212 31832 16264 31884
rect 16396 31832 16448 31884
rect 17868 31875 17920 31884
rect 17868 31841 17877 31875
rect 17877 31841 17911 31875
rect 17911 31841 17920 31875
rect 17868 31832 17920 31841
rect 10048 31764 10100 31816
rect 11336 31764 11388 31816
rect 15108 31764 15160 31816
rect 17224 31764 17276 31816
rect 17500 31764 17552 31816
rect 6000 31696 6052 31748
rect 15844 31696 15896 31748
rect 18880 31968 18932 32020
rect 25780 31968 25832 32020
rect 27252 31968 27304 32020
rect 18604 31875 18656 31884
rect 18604 31841 18613 31875
rect 18613 31841 18647 31875
rect 18647 31841 18656 31875
rect 18604 31832 18656 31841
rect 19156 31832 19208 31884
rect 18328 31807 18380 31816
rect 18328 31773 18337 31807
rect 18337 31773 18371 31807
rect 18371 31773 18380 31807
rect 18328 31764 18380 31773
rect 21456 31832 21508 31884
rect 22652 31875 22704 31884
rect 22652 31841 22661 31875
rect 22661 31841 22695 31875
rect 22695 31841 22704 31875
rect 22652 31832 22704 31841
rect 27344 31900 27396 31952
rect 33692 31968 33744 32020
rect 33876 31900 33928 31952
rect 36176 31900 36228 31952
rect 37096 31900 37148 31952
rect 21088 31764 21140 31816
rect 20444 31696 20496 31748
rect 23480 31764 23532 31816
rect 24400 31764 24452 31816
rect 24676 31764 24728 31816
rect 26056 31764 26108 31816
rect 5632 31671 5684 31680
rect 5632 31637 5641 31671
rect 5641 31637 5675 31671
rect 5675 31637 5684 31671
rect 5632 31628 5684 31637
rect 6092 31628 6144 31680
rect 9864 31628 9916 31680
rect 14648 31671 14700 31680
rect 14648 31637 14657 31671
rect 14657 31637 14691 31671
rect 14691 31637 14700 31671
rect 14648 31628 14700 31637
rect 20720 31628 20772 31680
rect 24032 31628 24084 31680
rect 27160 31832 27212 31884
rect 30012 31832 30064 31884
rect 30288 31875 30340 31884
rect 30288 31841 30297 31875
rect 30297 31841 30331 31875
rect 30331 31841 30340 31875
rect 30288 31832 30340 31841
rect 27252 31807 27304 31816
rect 27252 31773 27261 31807
rect 27261 31773 27295 31807
rect 27295 31773 27304 31807
rect 27252 31764 27304 31773
rect 27620 31764 27672 31816
rect 29460 31764 29512 31816
rect 29552 31764 29604 31816
rect 32128 31875 32180 31884
rect 32128 31841 32137 31875
rect 32137 31841 32171 31875
rect 32171 31841 32180 31875
rect 32128 31832 32180 31841
rect 32404 31875 32456 31884
rect 32404 31841 32413 31875
rect 32413 31841 32447 31875
rect 32447 31841 32456 31875
rect 32404 31832 32456 31841
rect 34520 31875 34572 31884
rect 34520 31841 34529 31875
rect 34529 31841 34563 31875
rect 34563 31841 34572 31875
rect 36636 31875 36688 31884
rect 34520 31832 34572 31841
rect 34704 31764 34756 31816
rect 36636 31841 36645 31875
rect 36645 31841 36679 31875
rect 36679 31841 36688 31875
rect 36636 31832 36688 31841
rect 36820 31764 36872 31816
rect 30472 31696 30524 31748
rect 28448 31628 28500 31680
rect 36084 31671 36136 31680
rect 36084 31637 36093 31671
rect 36093 31637 36127 31671
rect 36127 31637 36136 31671
rect 36084 31628 36136 31637
rect 36728 31671 36780 31680
rect 36728 31637 36737 31671
rect 36737 31637 36771 31671
rect 36771 31637 36780 31671
rect 36728 31628 36780 31637
rect 38016 31628 38068 31680
rect 38936 31671 38988 31680
rect 38936 31637 38945 31671
rect 38945 31637 38979 31671
rect 38979 31637 38988 31671
rect 38936 31628 38988 31637
rect 4246 31526 4298 31578
rect 4310 31526 4362 31578
rect 4374 31526 4426 31578
rect 4438 31526 4490 31578
rect 34966 31526 35018 31578
rect 35030 31526 35082 31578
rect 35094 31526 35146 31578
rect 35158 31526 35210 31578
rect 2872 31424 2924 31476
rect 4068 31424 4120 31476
rect 9496 31467 9548 31476
rect 9496 31433 9505 31467
rect 9505 31433 9539 31467
rect 9539 31433 9548 31467
rect 9496 31424 9548 31433
rect 15108 31424 15160 31476
rect 18512 31424 18564 31476
rect 27344 31467 27396 31476
rect 27344 31433 27353 31467
rect 27353 31433 27387 31467
rect 27387 31433 27396 31467
rect 27344 31424 27396 31433
rect 9864 31356 9916 31408
rect 2688 31288 2740 31340
rect 1676 31263 1728 31272
rect 1676 31229 1685 31263
rect 1685 31229 1719 31263
rect 1719 31229 1728 31263
rect 1676 31220 1728 31229
rect 3976 31220 4028 31272
rect 4620 31288 4672 31340
rect 8208 31288 8260 31340
rect 4712 31220 4764 31272
rect 4896 31220 4948 31272
rect 6092 31263 6144 31272
rect 6092 31229 6101 31263
rect 6101 31229 6135 31263
rect 6135 31229 6144 31263
rect 6092 31220 6144 31229
rect 6460 31220 6512 31272
rect 8760 31220 8812 31272
rect 18328 31288 18380 31340
rect 19432 31288 19484 31340
rect 23480 31356 23532 31408
rect 23572 31356 23624 31408
rect 24216 31356 24268 31408
rect 27712 31356 27764 31408
rect 30840 31356 30892 31408
rect 12900 31263 12952 31272
rect 7380 31152 7432 31204
rect 10876 31195 10928 31204
rect 10876 31161 10885 31195
rect 10885 31161 10919 31195
rect 10919 31161 10928 31195
rect 10876 31152 10928 31161
rect 3240 31084 3292 31136
rect 5816 31084 5868 31136
rect 12900 31229 12909 31263
rect 12909 31229 12943 31263
rect 12943 31229 12952 31263
rect 12900 31220 12952 31229
rect 13636 31263 13688 31272
rect 13636 31229 13645 31263
rect 13645 31229 13679 31263
rect 13679 31229 13688 31263
rect 13636 31220 13688 31229
rect 14004 31220 14056 31272
rect 14648 31220 14700 31272
rect 15384 31220 15436 31272
rect 15568 31263 15620 31272
rect 15568 31229 15577 31263
rect 15577 31229 15611 31263
rect 15611 31229 15620 31263
rect 15568 31220 15620 31229
rect 15660 31220 15712 31272
rect 15292 31152 15344 31204
rect 13360 31084 13412 31136
rect 14648 31084 14700 31136
rect 17316 31152 17368 31204
rect 17776 31220 17828 31272
rect 19156 31263 19208 31272
rect 19156 31229 19165 31263
rect 19165 31229 19199 31263
rect 19199 31229 19208 31263
rect 19156 31220 19208 31229
rect 19892 31220 19944 31272
rect 20444 31263 20496 31272
rect 20444 31229 20453 31263
rect 20453 31229 20487 31263
rect 20487 31229 20496 31263
rect 20444 31220 20496 31229
rect 21640 31263 21692 31272
rect 18604 31152 18656 31204
rect 21640 31229 21649 31263
rect 21649 31229 21683 31263
rect 21683 31229 21692 31263
rect 21640 31220 21692 31229
rect 23572 31220 23624 31272
rect 22560 31152 22612 31204
rect 24032 31220 24084 31272
rect 26240 31263 26292 31272
rect 26240 31229 26249 31263
rect 26249 31229 26283 31263
rect 26283 31229 26292 31263
rect 26240 31220 26292 31229
rect 26424 31263 26476 31272
rect 26424 31229 26433 31263
rect 26433 31229 26467 31263
rect 26467 31229 26476 31263
rect 26424 31220 26476 31229
rect 27160 31220 27212 31272
rect 27896 31152 27948 31204
rect 29000 31220 29052 31272
rect 29460 31263 29512 31272
rect 29460 31229 29469 31263
rect 29469 31229 29503 31263
rect 29503 31229 29512 31263
rect 29460 31220 29512 31229
rect 30472 31263 30524 31272
rect 28540 31152 28592 31204
rect 28816 31152 28868 31204
rect 30472 31229 30481 31263
rect 30481 31229 30515 31263
rect 30515 31229 30524 31263
rect 30472 31220 30524 31229
rect 34796 31424 34848 31476
rect 34888 31356 34940 31408
rect 31576 31220 31628 31272
rect 32220 31220 32272 31272
rect 33324 31288 33376 31340
rect 33232 31220 33284 31272
rect 34796 31220 34848 31272
rect 35808 31263 35860 31272
rect 33600 31152 33652 31204
rect 33784 31195 33836 31204
rect 33784 31161 33793 31195
rect 33793 31161 33827 31195
rect 33827 31161 33836 31195
rect 35808 31229 35817 31263
rect 35817 31229 35851 31263
rect 35851 31229 35860 31263
rect 35808 31220 35860 31229
rect 36084 31220 36136 31272
rect 36820 31220 36872 31272
rect 37740 31263 37792 31272
rect 37740 31229 37749 31263
rect 37749 31229 37783 31263
rect 37783 31229 37792 31263
rect 37740 31220 37792 31229
rect 33784 31152 33836 31161
rect 35900 31152 35952 31204
rect 18052 31084 18104 31136
rect 18328 31084 18380 31136
rect 21548 31084 21600 31136
rect 22376 31084 22428 31136
rect 28448 31127 28500 31136
rect 28448 31093 28457 31127
rect 28457 31093 28491 31127
rect 28491 31093 28500 31127
rect 28448 31084 28500 31093
rect 28908 31084 28960 31136
rect 33048 31084 33100 31136
rect 38660 31084 38712 31136
rect 19606 30982 19658 31034
rect 19670 30982 19722 31034
rect 19734 30982 19786 31034
rect 19798 30982 19850 31034
rect 1676 30880 1728 30932
rect 17776 30880 17828 30932
rect 34704 30880 34756 30932
rect 2872 30812 2924 30864
rect 7196 30855 7248 30864
rect 7196 30821 7205 30855
rect 7205 30821 7239 30855
rect 7239 30821 7248 30855
rect 7196 30812 7248 30821
rect 17500 30812 17552 30864
rect 30380 30812 30432 30864
rect 2688 30787 2740 30796
rect 2688 30753 2697 30787
rect 2697 30753 2731 30787
rect 2731 30753 2740 30787
rect 2688 30744 2740 30753
rect 3240 30787 3292 30796
rect 3240 30753 3249 30787
rect 3249 30753 3283 30787
rect 3283 30753 3292 30787
rect 3240 30744 3292 30753
rect 3700 30744 3752 30796
rect 4068 30787 4120 30796
rect 4068 30753 4077 30787
rect 4077 30753 4111 30787
rect 4111 30753 4120 30787
rect 4068 30744 4120 30753
rect 5632 30744 5684 30796
rect 7656 30787 7708 30796
rect 7656 30753 7665 30787
rect 7665 30753 7699 30787
rect 7699 30753 7708 30787
rect 7656 30744 7708 30753
rect 7840 30787 7892 30796
rect 7840 30753 7849 30787
rect 7849 30753 7883 30787
rect 7883 30753 7892 30787
rect 7840 30744 7892 30753
rect 5080 30719 5132 30728
rect 5080 30685 5089 30719
rect 5089 30685 5123 30719
rect 5123 30685 5132 30719
rect 5080 30676 5132 30685
rect 7012 30676 7064 30728
rect 8392 30744 8444 30796
rect 10416 30787 10468 30796
rect 10416 30753 10425 30787
rect 10425 30753 10459 30787
rect 10459 30753 10468 30787
rect 10416 30744 10468 30753
rect 10876 30744 10928 30796
rect 14280 30744 14332 30796
rect 11152 30676 11204 30728
rect 14188 30719 14240 30728
rect 14188 30685 14197 30719
rect 14197 30685 14231 30719
rect 14231 30685 14240 30719
rect 14188 30676 14240 30685
rect 14832 30744 14884 30796
rect 15844 30744 15896 30796
rect 16212 30787 16264 30796
rect 16212 30753 16221 30787
rect 16221 30753 16255 30787
rect 16255 30753 16264 30787
rect 16212 30744 16264 30753
rect 17132 30744 17184 30796
rect 17316 30744 17368 30796
rect 17960 30744 18012 30796
rect 19156 30787 19208 30796
rect 19156 30753 19165 30787
rect 19165 30753 19199 30787
rect 19199 30753 19208 30787
rect 19156 30744 19208 30753
rect 19432 30787 19484 30796
rect 19432 30753 19441 30787
rect 19441 30753 19475 30787
rect 19475 30753 19484 30787
rect 19432 30744 19484 30753
rect 19892 30787 19944 30796
rect 19892 30753 19901 30787
rect 19901 30753 19935 30787
rect 19935 30753 19944 30787
rect 19892 30744 19944 30753
rect 21548 30787 21600 30796
rect 21548 30753 21557 30787
rect 21557 30753 21591 30787
rect 21591 30753 21600 30787
rect 21548 30744 21600 30753
rect 23664 30787 23716 30796
rect 23664 30753 23673 30787
rect 23673 30753 23707 30787
rect 23707 30753 23716 30787
rect 23664 30744 23716 30753
rect 15476 30676 15528 30728
rect 18236 30676 18288 30728
rect 23020 30676 23072 30728
rect 24216 30787 24268 30796
rect 24216 30753 24225 30787
rect 24225 30753 24259 30787
rect 24259 30753 24268 30787
rect 24216 30744 24268 30753
rect 24584 30787 24636 30796
rect 24584 30753 24593 30787
rect 24593 30753 24627 30787
rect 24627 30753 24636 30787
rect 24584 30744 24636 30753
rect 25320 30787 25372 30796
rect 25320 30753 25329 30787
rect 25329 30753 25363 30787
rect 25363 30753 25372 30787
rect 25320 30744 25372 30753
rect 27712 30787 27764 30796
rect 27712 30753 27721 30787
rect 27721 30753 27755 30787
rect 27755 30753 27764 30787
rect 27712 30744 27764 30753
rect 28172 30744 28224 30796
rect 26884 30719 26936 30728
rect 26884 30685 26893 30719
rect 26893 30685 26927 30719
rect 26927 30685 26936 30719
rect 26884 30676 26936 30685
rect 26976 30676 27028 30728
rect 30288 30744 30340 30796
rect 30564 30787 30616 30796
rect 30564 30753 30573 30787
rect 30573 30753 30607 30787
rect 30607 30753 30616 30787
rect 30564 30744 30616 30753
rect 33324 30812 33376 30864
rect 30012 30676 30064 30728
rect 32220 30719 32272 30728
rect 7104 30608 7156 30660
rect 15200 30608 15252 30660
rect 27620 30651 27672 30660
rect 27620 30617 27629 30651
rect 27629 30617 27663 30651
rect 27663 30617 27672 30651
rect 27620 30608 27672 30617
rect 31116 30608 31168 30660
rect 32220 30685 32229 30719
rect 32229 30685 32263 30719
rect 32263 30685 32272 30719
rect 32220 30676 32272 30685
rect 33048 30787 33100 30796
rect 33048 30753 33057 30787
rect 33057 30753 33091 30787
rect 33091 30753 33100 30787
rect 33048 30744 33100 30753
rect 33140 30744 33192 30796
rect 34888 30787 34940 30796
rect 34888 30753 34897 30787
rect 34897 30753 34931 30787
rect 34931 30753 34940 30787
rect 34888 30744 34940 30753
rect 34244 30676 34296 30728
rect 36084 30719 36136 30728
rect 36084 30685 36093 30719
rect 36093 30685 36127 30719
rect 36127 30685 36136 30719
rect 36084 30676 36136 30685
rect 36728 30744 36780 30796
rect 37464 30744 37516 30796
rect 37924 30744 37976 30796
rect 38016 30676 38068 30728
rect 38844 30719 38896 30728
rect 38844 30685 38853 30719
rect 38853 30685 38887 30719
rect 38887 30685 38896 30719
rect 38844 30676 38896 30685
rect 2780 30540 2832 30592
rect 4712 30540 4764 30592
rect 8944 30540 8996 30592
rect 9220 30540 9272 30592
rect 9864 30583 9916 30592
rect 9864 30549 9873 30583
rect 9873 30549 9907 30583
rect 9907 30549 9916 30583
rect 9864 30540 9916 30549
rect 10140 30540 10192 30592
rect 10600 30583 10652 30592
rect 10600 30549 10609 30583
rect 10609 30549 10643 30583
rect 10643 30549 10652 30583
rect 10600 30540 10652 30549
rect 11704 30540 11756 30592
rect 15660 30540 15712 30592
rect 16120 30540 16172 30592
rect 22652 30583 22704 30592
rect 22652 30549 22661 30583
rect 22661 30549 22695 30583
rect 22695 30549 22704 30583
rect 22652 30540 22704 30549
rect 25596 30540 25648 30592
rect 29000 30540 29052 30592
rect 29276 30540 29328 30592
rect 31576 30540 31628 30592
rect 32772 30540 32824 30592
rect 34244 30540 34296 30592
rect 4246 30438 4298 30490
rect 4310 30438 4362 30490
rect 4374 30438 4426 30490
rect 4438 30438 4490 30490
rect 34966 30438 35018 30490
rect 35030 30438 35082 30490
rect 35094 30438 35146 30490
rect 35158 30438 35210 30490
rect 9864 30336 9916 30388
rect 10232 30336 10284 30388
rect 10416 30336 10468 30388
rect 10968 30336 11020 30388
rect 3700 30311 3752 30320
rect 3700 30277 3709 30311
rect 3709 30277 3743 30311
rect 3743 30277 3752 30311
rect 3700 30268 3752 30277
rect 7656 30311 7708 30320
rect 7656 30277 7665 30311
rect 7665 30277 7699 30311
rect 7699 30277 7708 30311
rect 7656 30268 7708 30277
rect 9956 30268 10008 30320
rect 10600 30268 10652 30320
rect 2412 30175 2464 30184
rect 2412 30141 2421 30175
rect 2421 30141 2455 30175
rect 2455 30141 2464 30175
rect 2412 30132 2464 30141
rect 2780 30175 2832 30184
rect 2780 30141 2789 30175
rect 2789 30141 2823 30175
rect 2823 30141 2832 30175
rect 2780 30132 2832 30141
rect 3056 30132 3108 30184
rect 4620 30200 4672 30252
rect 3240 30132 3292 30184
rect 4068 30132 4120 30184
rect 4528 30175 4580 30184
rect 4528 30141 4537 30175
rect 4537 30141 4571 30175
rect 4571 30141 4580 30175
rect 4528 30132 4580 30141
rect 4712 30175 4764 30184
rect 4712 30141 4721 30175
rect 4721 30141 4755 30175
rect 4755 30141 4764 30175
rect 5816 30175 5868 30184
rect 4712 30132 4764 30141
rect 5816 30141 5825 30175
rect 5825 30141 5859 30175
rect 5859 30141 5868 30175
rect 5816 30132 5868 30141
rect 7012 30175 7064 30184
rect 5448 30064 5500 30116
rect 7012 30141 7021 30175
rect 7021 30141 7055 30175
rect 7055 30141 7064 30175
rect 7012 30132 7064 30141
rect 7840 30200 7892 30252
rect 8300 30200 8352 30252
rect 8484 30200 8536 30252
rect 9588 30200 9640 30252
rect 8392 30175 8444 30184
rect 8392 30141 8401 30175
rect 8401 30141 8435 30175
rect 8435 30141 8444 30175
rect 8392 30132 8444 30141
rect 9312 30175 9364 30184
rect 9312 30141 9321 30175
rect 9321 30141 9355 30175
rect 9355 30141 9364 30175
rect 9312 30132 9364 30141
rect 10140 30132 10192 30184
rect 10232 30132 10284 30184
rect 11336 30175 11388 30184
rect 11336 30141 11345 30175
rect 11345 30141 11379 30175
rect 11379 30141 11388 30175
rect 11336 30132 11388 30141
rect 11704 30336 11756 30388
rect 12992 30336 13044 30388
rect 19340 30336 19392 30388
rect 20444 30336 20496 30388
rect 26240 30336 26292 30388
rect 26976 30336 27028 30388
rect 12440 30268 12492 30320
rect 17960 30268 18012 30320
rect 18052 30268 18104 30320
rect 14832 30200 14884 30252
rect 15568 30243 15620 30252
rect 12532 30175 12584 30184
rect 12532 30141 12541 30175
rect 12541 30141 12575 30175
rect 12575 30141 12584 30175
rect 12532 30132 12584 30141
rect 13912 30175 13964 30184
rect 8300 30064 8352 30116
rect 13912 30141 13921 30175
rect 13921 30141 13955 30175
rect 13955 30141 13964 30175
rect 13912 30132 13964 30141
rect 14464 30175 14516 30184
rect 14464 30141 14473 30175
rect 14473 30141 14507 30175
rect 14507 30141 14516 30175
rect 14464 30132 14516 30141
rect 15568 30209 15577 30243
rect 15577 30209 15611 30243
rect 15611 30209 15620 30243
rect 15568 30200 15620 30209
rect 15844 30132 15896 30184
rect 17224 30200 17276 30252
rect 16396 30175 16448 30184
rect 16396 30141 16405 30175
rect 16405 30141 16439 30175
rect 16439 30141 16448 30175
rect 16396 30132 16448 30141
rect 16764 30132 16816 30184
rect 14648 30064 14700 30116
rect 19248 30200 19300 30252
rect 19892 30200 19944 30252
rect 17868 30132 17920 30184
rect 18328 30175 18380 30184
rect 18328 30141 18337 30175
rect 18337 30141 18371 30175
rect 18371 30141 18380 30175
rect 18328 30132 18380 30141
rect 20168 30175 20220 30184
rect 20168 30141 20177 30175
rect 20177 30141 20211 30175
rect 20211 30141 20220 30175
rect 20168 30132 20220 30141
rect 21640 30200 21692 30252
rect 26056 30200 26108 30252
rect 29460 30243 29512 30252
rect 29460 30209 29469 30243
rect 29469 30209 29503 30243
rect 29503 30209 29512 30243
rect 29460 30200 29512 30209
rect 32036 30336 32088 30388
rect 32220 30379 32272 30388
rect 32220 30345 32229 30379
rect 32229 30345 32263 30379
rect 32263 30345 32272 30379
rect 32220 30336 32272 30345
rect 37464 30379 37516 30388
rect 37464 30345 37473 30379
rect 37473 30345 37507 30379
rect 37507 30345 37516 30379
rect 37464 30336 37516 30345
rect 35900 30268 35952 30320
rect 37740 30268 37792 30320
rect 31116 30243 31168 30252
rect 31116 30209 31125 30243
rect 31125 30209 31159 30243
rect 31159 30209 31168 30243
rect 31116 30200 31168 30209
rect 34244 30243 34296 30252
rect 34244 30209 34253 30243
rect 34253 30209 34287 30243
rect 34287 30209 34296 30243
rect 34244 30200 34296 30209
rect 3148 29996 3200 30048
rect 8760 29996 8812 30048
rect 9128 30039 9180 30048
rect 9128 30005 9137 30039
rect 9137 30005 9171 30039
rect 9171 30005 9180 30039
rect 9128 29996 9180 30005
rect 9220 29996 9272 30048
rect 13820 29996 13872 30048
rect 17960 29996 18012 30048
rect 19156 30064 19208 30116
rect 22008 30132 22060 30184
rect 21272 30107 21324 30116
rect 21272 30073 21281 30107
rect 21281 30073 21315 30107
rect 21315 30073 21324 30107
rect 22652 30132 22704 30184
rect 23204 30132 23256 30184
rect 23940 30175 23992 30184
rect 23940 30141 23949 30175
rect 23949 30141 23983 30175
rect 23983 30141 23992 30175
rect 23940 30132 23992 30141
rect 25228 30175 25280 30184
rect 21272 30064 21324 30073
rect 23296 30064 23348 30116
rect 25228 30141 25237 30175
rect 25237 30141 25271 30175
rect 25271 30141 25280 30175
rect 25228 30132 25280 30141
rect 27344 30175 27396 30184
rect 27344 30141 27353 30175
rect 27353 30141 27387 30175
rect 27387 30141 27396 30175
rect 27344 30132 27396 30141
rect 30012 30132 30064 30184
rect 30288 30132 30340 30184
rect 33140 30132 33192 30184
rect 36084 30200 36136 30252
rect 38844 30243 38896 30252
rect 38844 30209 38853 30243
rect 38853 30209 38887 30243
rect 38887 30209 38896 30243
rect 38844 30200 38896 30209
rect 28724 30107 28776 30116
rect 28724 30073 28733 30107
rect 28733 30073 28767 30107
rect 28767 30073 28776 30107
rect 28724 30064 28776 30073
rect 32496 30064 32548 30116
rect 35256 30132 35308 30184
rect 36820 30132 36872 30184
rect 38108 30175 38160 30184
rect 38108 30141 38117 30175
rect 38117 30141 38151 30175
rect 38151 30141 38160 30175
rect 38108 30132 38160 30141
rect 38752 30175 38804 30184
rect 38752 30141 38761 30175
rect 38761 30141 38795 30175
rect 38795 30141 38804 30175
rect 38752 30132 38804 30141
rect 34704 30064 34756 30116
rect 35716 30064 35768 30116
rect 21732 29996 21784 30048
rect 23664 29996 23716 30048
rect 33876 29996 33928 30048
rect 19606 29894 19658 29946
rect 19670 29894 19722 29946
rect 19734 29894 19786 29946
rect 19798 29894 19850 29946
rect 5540 29792 5592 29844
rect 6552 29792 6604 29844
rect 4528 29724 4580 29776
rect 9312 29792 9364 29844
rect 13636 29792 13688 29844
rect 14004 29792 14056 29844
rect 16304 29792 16356 29844
rect 4620 29699 4672 29708
rect 1400 29631 1452 29640
rect 1400 29597 1409 29631
rect 1409 29597 1443 29631
rect 1443 29597 1452 29631
rect 1400 29588 1452 29597
rect 1860 29588 1912 29640
rect 3148 29452 3200 29504
rect 3976 29452 4028 29504
rect 4620 29665 4629 29699
rect 4629 29665 4663 29699
rect 4663 29665 4672 29699
rect 4620 29656 4672 29665
rect 5448 29656 5500 29708
rect 4896 29631 4948 29640
rect 4896 29597 4905 29631
rect 4905 29597 4939 29631
rect 4939 29597 4948 29631
rect 4896 29588 4948 29597
rect 5816 29631 5868 29640
rect 5816 29597 5825 29631
rect 5825 29597 5859 29631
rect 5859 29597 5868 29631
rect 5816 29588 5868 29597
rect 4804 29520 4856 29572
rect 5632 29520 5684 29572
rect 7012 29656 7064 29708
rect 9588 29724 9640 29776
rect 9772 29724 9824 29776
rect 7380 29588 7432 29640
rect 8116 29656 8168 29708
rect 13912 29724 13964 29776
rect 15476 29724 15528 29776
rect 13360 29699 13412 29708
rect 11152 29588 11204 29640
rect 12532 29631 12584 29640
rect 12532 29597 12541 29631
rect 12541 29597 12575 29631
rect 12575 29597 12584 29631
rect 12532 29588 12584 29597
rect 9680 29520 9732 29572
rect 12256 29520 12308 29572
rect 13360 29665 13369 29699
rect 13369 29665 13403 29699
rect 13403 29665 13412 29699
rect 13360 29656 13412 29665
rect 14096 29656 14148 29708
rect 14280 29699 14332 29708
rect 14280 29665 14289 29699
rect 14289 29665 14323 29699
rect 14323 29665 14332 29699
rect 14280 29656 14332 29665
rect 15200 29656 15252 29708
rect 15844 29656 15896 29708
rect 16764 29724 16816 29776
rect 16120 29699 16172 29708
rect 16120 29665 16129 29699
rect 16129 29665 16163 29699
rect 16163 29665 16172 29699
rect 16120 29656 16172 29665
rect 16304 29656 16356 29708
rect 19064 29699 19116 29708
rect 19064 29665 19073 29699
rect 19073 29665 19107 29699
rect 19107 29665 19116 29699
rect 19064 29656 19116 29665
rect 25320 29792 25372 29844
rect 25412 29792 25464 29844
rect 22008 29767 22060 29776
rect 22008 29733 22017 29767
rect 22017 29733 22051 29767
rect 22051 29733 22060 29767
rect 22008 29724 22060 29733
rect 24584 29724 24636 29776
rect 19984 29656 20036 29708
rect 21272 29699 21324 29708
rect 21272 29665 21281 29699
rect 21281 29665 21315 29699
rect 21315 29665 21324 29699
rect 21272 29656 21324 29665
rect 21732 29699 21784 29708
rect 21732 29665 21741 29699
rect 21741 29665 21775 29699
rect 21775 29665 21784 29699
rect 21732 29656 21784 29665
rect 19340 29588 19392 29640
rect 22652 29588 22704 29640
rect 12900 29520 12952 29572
rect 15200 29520 15252 29572
rect 15292 29520 15344 29572
rect 17316 29520 17368 29572
rect 23388 29656 23440 29708
rect 24032 29699 24084 29708
rect 24032 29665 24041 29699
rect 24041 29665 24075 29699
rect 24075 29665 24084 29699
rect 24032 29656 24084 29665
rect 24216 29699 24268 29708
rect 24216 29665 24225 29699
rect 24225 29665 24259 29699
rect 24259 29665 24268 29699
rect 24216 29656 24268 29665
rect 25320 29656 25372 29708
rect 27344 29724 27396 29776
rect 28080 29656 28132 29708
rect 32956 29792 33008 29844
rect 34796 29792 34848 29844
rect 38476 29792 38528 29844
rect 29276 29724 29328 29776
rect 30564 29767 30616 29776
rect 29368 29656 29420 29708
rect 30012 29699 30064 29708
rect 30012 29665 30021 29699
rect 30021 29665 30055 29699
rect 30055 29665 30064 29699
rect 30012 29656 30064 29665
rect 30288 29699 30340 29708
rect 30288 29665 30297 29699
rect 30297 29665 30331 29699
rect 30331 29665 30340 29699
rect 30288 29656 30340 29665
rect 30564 29733 30573 29767
rect 30573 29733 30607 29767
rect 30607 29733 30616 29767
rect 30564 29724 30616 29733
rect 32220 29724 32272 29776
rect 26884 29588 26936 29640
rect 23664 29520 23716 29572
rect 30380 29588 30432 29640
rect 32588 29656 32640 29708
rect 33876 29699 33928 29708
rect 33876 29665 33885 29699
rect 33885 29665 33919 29699
rect 33919 29665 33928 29699
rect 33876 29656 33928 29665
rect 37464 29724 37516 29776
rect 33232 29588 33284 29640
rect 34520 29588 34572 29640
rect 36820 29656 36872 29708
rect 38108 29699 38160 29708
rect 27252 29520 27304 29572
rect 31576 29520 31628 29572
rect 38108 29665 38117 29699
rect 38117 29665 38151 29699
rect 38151 29665 38160 29699
rect 38108 29656 38160 29665
rect 38016 29588 38068 29640
rect 38752 29520 38804 29572
rect 7748 29452 7800 29504
rect 8392 29452 8444 29504
rect 10784 29452 10836 29504
rect 10876 29452 10928 29504
rect 14004 29452 14056 29504
rect 19156 29452 19208 29504
rect 28632 29495 28684 29504
rect 28632 29461 28641 29495
rect 28641 29461 28675 29495
rect 28675 29461 28684 29495
rect 28632 29452 28684 29461
rect 36544 29495 36596 29504
rect 36544 29461 36553 29495
rect 36553 29461 36587 29495
rect 36587 29461 36596 29495
rect 36544 29452 36596 29461
rect 39028 29495 39080 29504
rect 39028 29461 39037 29495
rect 39037 29461 39071 29495
rect 39071 29461 39080 29495
rect 39028 29452 39080 29461
rect 4246 29350 4298 29402
rect 4310 29350 4362 29402
rect 4374 29350 4426 29402
rect 4438 29350 4490 29402
rect 34966 29350 35018 29402
rect 35030 29350 35082 29402
rect 35094 29350 35146 29402
rect 35158 29350 35210 29402
rect 1860 29291 1912 29300
rect 1860 29257 1869 29291
rect 1869 29257 1903 29291
rect 1903 29257 1912 29291
rect 1860 29248 1912 29257
rect 5080 29248 5132 29300
rect 8484 29248 8536 29300
rect 2964 29180 3016 29232
rect 2412 29087 2464 29096
rect 2412 29053 2421 29087
rect 2421 29053 2455 29087
rect 2455 29053 2464 29087
rect 2412 29044 2464 29053
rect 3056 29087 3108 29096
rect 3056 29053 3065 29087
rect 3065 29053 3099 29087
rect 3099 29053 3108 29087
rect 3056 29044 3108 29053
rect 3240 29087 3292 29096
rect 3240 29053 3249 29087
rect 3249 29053 3283 29087
rect 3283 29053 3292 29087
rect 3240 29044 3292 29053
rect 4160 29087 4212 29096
rect 4160 29053 4169 29087
rect 4169 29053 4203 29087
rect 4203 29053 4212 29087
rect 4160 29044 4212 29053
rect 4620 29044 4672 29096
rect 4804 29087 4856 29096
rect 4804 29053 4813 29087
rect 4813 29053 4847 29087
rect 4847 29053 4856 29087
rect 4804 29044 4856 29053
rect 7012 29180 7064 29232
rect 8392 29180 8444 29232
rect 4896 28976 4948 29028
rect 7012 29044 7064 29096
rect 8116 29112 8168 29164
rect 8300 29155 8352 29164
rect 8300 29121 8309 29155
rect 8309 29121 8343 29155
rect 8343 29121 8352 29155
rect 8300 29112 8352 29121
rect 7564 29087 7616 29096
rect 7564 29053 7573 29087
rect 7573 29053 7607 29087
rect 7607 29053 7616 29087
rect 13820 29248 13872 29300
rect 13912 29248 13964 29300
rect 9772 29180 9824 29232
rect 10876 29180 10928 29232
rect 11336 29180 11388 29232
rect 13636 29180 13688 29232
rect 16120 29248 16172 29300
rect 16672 29248 16724 29300
rect 8852 29087 8904 29096
rect 7564 29044 7616 29053
rect 8852 29053 8861 29087
rect 8861 29053 8895 29087
rect 8895 29053 8904 29087
rect 8852 29044 8904 29053
rect 6920 28976 6972 29028
rect 7748 28951 7800 28960
rect 7748 28917 7757 28951
rect 7757 28917 7791 28951
rect 7791 28917 7800 28951
rect 9220 29044 9272 29096
rect 9956 29087 10008 29096
rect 9956 29053 9965 29087
rect 9965 29053 9999 29087
rect 9999 29053 10008 29087
rect 9956 29044 10008 29053
rect 10600 29087 10652 29096
rect 10600 29053 10609 29087
rect 10609 29053 10643 29087
rect 10643 29053 10652 29087
rect 10600 29044 10652 29053
rect 10784 29044 10836 29096
rect 10416 28976 10468 29028
rect 14096 29112 14148 29164
rect 14464 29112 14516 29164
rect 16396 29112 16448 29164
rect 18328 29248 18380 29300
rect 12716 29087 12768 29096
rect 7748 28908 7800 28917
rect 9588 28908 9640 28960
rect 11704 28908 11756 28960
rect 12716 29053 12725 29087
rect 12725 29053 12759 29087
rect 12759 29053 12768 29087
rect 12716 29044 12768 29053
rect 14188 29044 14240 29096
rect 14648 29044 14700 29096
rect 14096 29019 14148 29028
rect 14096 28985 14105 29019
rect 14105 28985 14139 29019
rect 14139 28985 14148 29019
rect 14096 28976 14148 28985
rect 15660 29019 15712 29028
rect 15660 28985 15669 29019
rect 15669 28985 15703 29019
rect 15703 28985 15712 29019
rect 15660 28976 15712 28985
rect 16304 29044 16356 29096
rect 17316 29087 17368 29096
rect 17316 29053 17325 29087
rect 17325 29053 17359 29087
rect 17359 29053 17368 29087
rect 17316 29044 17368 29053
rect 18972 29044 19024 29096
rect 19064 29087 19116 29096
rect 19064 29053 19073 29087
rect 19073 29053 19107 29087
rect 19107 29053 19116 29087
rect 19064 29044 19116 29053
rect 15844 28976 15896 29028
rect 16120 28976 16172 29028
rect 20996 29248 21048 29300
rect 21364 29248 21416 29300
rect 20168 29180 20220 29232
rect 21088 29112 21140 29164
rect 22836 29180 22888 29232
rect 20444 29087 20496 29096
rect 20444 29053 20453 29087
rect 20453 29053 20487 29087
rect 20487 29053 20496 29087
rect 20444 29044 20496 29053
rect 21548 29087 21600 29096
rect 19432 28976 19484 29028
rect 21548 29053 21557 29087
rect 21557 29053 21591 29087
rect 21591 29053 21600 29087
rect 21548 29044 21600 29053
rect 22100 29087 22152 29096
rect 22100 29053 22109 29087
rect 22109 29053 22143 29087
rect 22143 29053 22152 29087
rect 23664 29087 23716 29096
rect 22100 29044 22152 29053
rect 23664 29053 23673 29087
rect 23673 29053 23707 29087
rect 23707 29053 23716 29087
rect 23664 29044 23716 29053
rect 23020 28976 23072 29028
rect 30748 29248 30800 29300
rect 25228 29180 25280 29232
rect 24584 29112 24636 29164
rect 28080 29155 28132 29164
rect 24400 29044 24452 29096
rect 24768 29044 24820 29096
rect 25596 29087 25648 29096
rect 25596 29053 25605 29087
rect 25605 29053 25639 29087
rect 25639 29053 25648 29087
rect 25596 29044 25648 29053
rect 28080 29121 28089 29155
rect 28089 29121 28123 29155
rect 28123 29121 28132 29155
rect 28080 29112 28132 29121
rect 31576 29112 31628 29164
rect 26424 29087 26476 29096
rect 26424 29053 26433 29087
rect 26433 29053 26467 29087
rect 26467 29053 26476 29087
rect 26424 29044 26476 29053
rect 27252 29087 27304 29096
rect 27252 29053 27261 29087
rect 27261 29053 27295 29087
rect 27295 29053 27304 29087
rect 27252 29044 27304 29053
rect 28908 29087 28960 29096
rect 28908 29053 28917 29087
rect 28917 29053 28951 29087
rect 28951 29053 28960 29087
rect 28908 29044 28960 29053
rect 29552 29087 29604 29096
rect 29552 29053 29561 29087
rect 29561 29053 29595 29087
rect 29595 29053 29604 29087
rect 29552 29044 29604 29053
rect 31300 29044 31352 29096
rect 32312 29044 32364 29096
rect 33140 29180 33192 29232
rect 32588 29112 32640 29164
rect 34704 29180 34756 29232
rect 37096 29180 37148 29232
rect 38016 29155 38068 29164
rect 33232 29087 33284 29096
rect 33232 29053 33241 29087
rect 33241 29053 33275 29087
rect 33275 29053 33284 29087
rect 33232 29044 33284 29053
rect 29276 28976 29328 29028
rect 34796 29044 34848 29096
rect 38016 29121 38025 29155
rect 38025 29121 38059 29155
rect 38059 29121 38068 29155
rect 38016 29112 38068 29121
rect 35716 29087 35768 29096
rect 35716 29053 35725 29087
rect 35725 29053 35759 29087
rect 35759 29053 35768 29087
rect 35716 29044 35768 29053
rect 36820 29044 36872 29096
rect 37464 29087 37516 29096
rect 37464 29053 37473 29087
rect 37473 29053 37507 29087
rect 37507 29053 37516 29087
rect 37464 29044 37516 29053
rect 37924 29087 37976 29096
rect 37924 29053 37933 29087
rect 37933 29053 37967 29087
rect 37967 29053 37976 29087
rect 37924 29044 37976 29053
rect 38660 29087 38712 29096
rect 38660 29053 38669 29087
rect 38669 29053 38703 29087
rect 38703 29053 38712 29087
rect 38660 29044 38712 29053
rect 35900 28976 35952 29028
rect 15292 28908 15344 28960
rect 18512 28908 18564 28960
rect 18788 28908 18840 28960
rect 18880 28908 18932 28960
rect 20168 28908 20220 28960
rect 20628 28908 20680 28960
rect 27712 28908 27764 28960
rect 33600 28908 33652 28960
rect 36452 28908 36504 28960
rect 36728 28908 36780 28960
rect 19606 28806 19658 28858
rect 19670 28806 19722 28858
rect 19734 28806 19786 28858
rect 19798 28806 19850 28858
rect 4160 28704 4212 28756
rect 6920 28704 6972 28756
rect 5540 28636 5592 28688
rect 7380 28636 7432 28688
rect 2320 28568 2372 28620
rect 3148 28611 3200 28620
rect 3148 28577 3157 28611
rect 3157 28577 3191 28611
rect 3191 28577 3200 28611
rect 3148 28568 3200 28577
rect 5356 28568 5408 28620
rect 9128 28636 9180 28688
rect 11336 28636 11388 28688
rect 4712 28500 4764 28552
rect 5080 28500 5132 28552
rect 5724 28543 5776 28552
rect 5724 28509 5733 28543
rect 5733 28509 5767 28543
rect 5767 28509 5776 28543
rect 5724 28500 5776 28509
rect 8208 28543 8260 28552
rect 8208 28509 8217 28543
rect 8217 28509 8251 28543
rect 8251 28509 8260 28543
rect 8208 28500 8260 28509
rect 10140 28568 10192 28620
rect 10600 28611 10652 28620
rect 10600 28577 10609 28611
rect 10609 28577 10643 28611
rect 10643 28577 10652 28611
rect 10600 28568 10652 28577
rect 10876 28568 10928 28620
rect 15568 28704 15620 28756
rect 9128 28543 9180 28552
rect 9128 28509 9137 28543
rect 9137 28509 9171 28543
rect 9171 28509 9180 28543
rect 9128 28500 9180 28509
rect 20076 28636 20128 28688
rect 20352 28636 20404 28688
rect 13636 28568 13688 28620
rect 14096 28568 14148 28620
rect 15292 28611 15344 28620
rect 15292 28577 15301 28611
rect 15301 28577 15335 28611
rect 15335 28577 15344 28611
rect 15292 28568 15344 28577
rect 18052 28568 18104 28620
rect 18512 28611 18564 28620
rect 18512 28577 18521 28611
rect 18521 28577 18555 28611
rect 18555 28577 18564 28611
rect 18512 28568 18564 28577
rect 20996 28568 21048 28620
rect 21548 28568 21600 28620
rect 24216 28704 24268 28756
rect 24768 28704 24820 28756
rect 27252 28704 27304 28756
rect 30288 28704 30340 28756
rect 22100 28568 22152 28620
rect 23296 28611 23348 28620
rect 23296 28577 23305 28611
rect 23305 28577 23339 28611
rect 23339 28577 23348 28611
rect 23296 28568 23348 28577
rect 23848 28568 23900 28620
rect 24400 28611 24452 28620
rect 24400 28577 24409 28611
rect 24409 28577 24443 28611
rect 24443 28577 24452 28611
rect 24400 28568 24452 28577
rect 24768 28611 24820 28620
rect 24768 28577 24777 28611
rect 24777 28577 24811 28611
rect 24811 28577 24820 28611
rect 24768 28568 24820 28577
rect 25412 28568 25464 28620
rect 27252 28611 27304 28620
rect 11244 28432 11296 28484
rect 11612 28432 11664 28484
rect 14004 28500 14056 28552
rect 15476 28500 15528 28552
rect 15752 28500 15804 28552
rect 17960 28500 18012 28552
rect 18236 28543 18288 28552
rect 18236 28509 18245 28543
rect 18245 28509 18279 28543
rect 18279 28509 18288 28543
rect 18236 28500 18288 28509
rect 19248 28500 19300 28552
rect 24676 28543 24728 28552
rect 24676 28509 24685 28543
rect 24685 28509 24719 28543
rect 24719 28509 24728 28543
rect 24676 28500 24728 28509
rect 12624 28432 12676 28484
rect 1952 28407 2004 28416
rect 1952 28373 1961 28407
rect 1961 28373 1995 28407
rect 1995 28373 2004 28407
rect 1952 28364 2004 28373
rect 2412 28407 2464 28416
rect 2412 28373 2421 28407
rect 2421 28373 2455 28407
rect 2455 28373 2464 28407
rect 2412 28364 2464 28373
rect 4620 28364 4672 28416
rect 11152 28364 11204 28416
rect 11704 28364 11756 28416
rect 22284 28432 22336 28484
rect 23756 28432 23808 28484
rect 27252 28577 27261 28611
rect 27261 28577 27295 28611
rect 27295 28577 27304 28611
rect 27252 28568 27304 28577
rect 28080 28611 28132 28620
rect 28080 28577 28089 28611
rect 28089 28577 28123 28611
rect 28123 28577 28132 28611
rect 28080 28568 28132 28577
rect 28724 28568 28776 28620
rect 30380 28611 30432 28620
rect 30380 28577 30389 28611
rect 30389 28577 30423 28611
rect 30423 28577 30432 28611
rect 30380 28568 30432 28577
rect 32496 28636 32548 28688
rect 35624 28704 35676 28756
rect 35256 28679 35308 28688
rect 35256 28645 35265 28679
rect 35265 28645 35299 28679
rect 35299 28645 35308 28679
rect 35256 28636 35308 28645
rect 36636 28636 36688 28688
rect 35716 28611 35768 28620
rect 27620 28500 27672 28552
rect 27712 28500 27764 28552
rect 32772 28500 32824 28552
rect 33876 28543 33928 28552
rect 33876 28509 33885 28543
rect 33885 28509 33919 28543
rect 33919 28509 33928 28543
rect 33876 28500 33928 28509
rect 35716 28577 35725 28611
rect 35725 28577 35759 28611
rect 35759 28577 35768 28611
rect 35716 28568 35768 28577
rect 36360 28611 36412 28620
rect 36360 28577 36369 28611
rect 36369 28577 36403 28611
rect 36403 28577 36412 28611
rect 36360 28568 36412 28577
rect 36544 28611 36596 28620
rect 36544 28577 36553 28611
rect 36553 28577 36587 28611
rect 36587 28577 36596 28611
rect 36544 28568 36596 28577
rect 38292 28611 38344 28620
rect 38292 28577 38301 28611
rect 38301 28577 38335 28611
rect 38335 28577 38344 28611
rect 38292 28568 38344 28577
rect 38476 28611 38528 28620
rect 38476 28577 38485 28611
rect 38485 28577 38519 28611
rect 38519 28577 38528 28611
rect 38476 28568 38528 28577
rect 38844 28568 38896 28620
rect 33508 28432 33560 28484
rect 16580 28364 16632 28416
rect 16764 28364 16816 28416
rect 19248 28364 19300 28416
rect 19984 28364 20036 28416
rect 26608 28407 26660 28416
rect 26608 28373 26617 28407
rect 26617 28373 26651 28407
rect 26651 28373 26660 28407
rect 26608 28364 26660 28373
rect 29644 28364 29696 28416
rect 34244 28364 34296 28416
rect 4246 28262 4298 28314
rect 4310 28262 4362 28314
rect 4374 28262 4426 28314
rect 4438 28262 4490 28314
rect 34966 28262 35018 28314
rect 35030 28262 35082 28314
rect 35094 28262 35146 28314
rect 35158 28262 35210 28314
rect 2320 27956 2372 28008
rect 4068 28092 4120 28144
rect 3240 28067 3292 28076
rect 3240 28033 3249 28067
rect 3249 28033 3283 28067
rect 3283 28033 3292 28067
rect 3240 28024 3292 28033
rect 2964 27999 3016 28008
rect 2964 27965 2973 27999
rect 2973 27965 3007 27999
rect 3007 27965 3016 27999
rect 2964 27956 3016 27965
rect 3332 27999 3384 28008
rect 3332 27965 3341 27999
rect 3341 27965 3375 27999
rect 3375 27965 3384 27999
rect 3332 27956 3384 27965
rect 4436 27956 4488 28008
rect 15476 28203 15528 28212
rect 15476 28169 15485 28203
rect 15485 28169 15519 28203
rect 15519 28169 15528 28203
rect 15476 28160 15528 28169
rect 16120 28203 16172 28212
rect 16120 28169 16129 28203
rect 16129 28169 16163 28203
rect 16163 28169 16172 28203
rect 16120 28160 16172 28169
rect 16580 28160 16632 28212
rect 24768 28160 24820 28212
rect 31760 28160 31812 28212
rect 32772 28203 32824 28212
rect 32772 28169 32781 28203
rect 32781 28169 32815 28203
rect 32815 28169 32824 28203
rect 32772 28160 32824 28169
rect 35808 28160 35860 28212
rect 36820 28160 36872 28212
rect 5724 28092 5776 28144
rect 7104 28092 7156 28144
rect 11152 28092 11204 28144
rect 11336 28092 11388 28144
rect 5632 27956 5684 28008
rect 5816 27999 5868 28008
rect 5816 27965 5825 27999
rect 5825 27965 5859 27999
rect 5859 27965 5868 27999
rect 5816 27956 5868 27965
rect 6828 27999 6880 28008
rect 5448 27888 5500 27940
rect 6828 27965 6837 27999
rect 6837 27965 6871 27999
rect 6871 27965 6880 27999
rect 6828 27956 6880 27965
rect 9680 28024 9732 28076
rect 12164 28092 12216 28144
rect 16672 28135 16724 28144
rect 9128 27956 9180 28008
rect 16672 28101 16681 28135
rect 16681 28101 16715 28135
rect 16715 28101 16724 28135
rect 16672 28092 16724 28101
rect 18236 28092 18288 28144
rect 20536 28092 20588 28144
rect 24584 28092 24636 28144
rect 27804 28092 27856 28144
rect 33048 28092 33100 28144
rect 8944 27888 8996 27940
rect 11612 27956 11664 28008
rect 13636 27999 13688 28008
rect 13636 27965 13645 27999
rect 13645 27965 13679 27999
rect 13679 27965 13688 27999
rect 13636 27956 13688 27965
rect 14004 27999 14056 28008
rect 14004 27965 14013 27999
rect 14013 27965 14047 27999
rect 14047 27965 14056 27999
rect 14004 27956 14056 27965
rect 15384 27999 15436 28008
rect 15384 27965 15393 27999
rect 15393 27965 15427 27999
rect 15427 27965 15436 27999
rect 15384 27956 15436 27965
rect 16304 27999 16356 28008
rect 16304 27965 16313 27999
rect 16313 27965 16347 27999
rect 16347 27965 16356 27999
rect 16304 27956 16356 27965
rect 16396 27999 16448 28008
rect 16396 27965 16405 27999
rect 16405 27965 16439 27999
rect 16439 27965 16448 27999
rect 17040 27999 17092 28008
rect 16396 27956 16448 27965
rect 17040 27965 17049 27999
rect 17049 27965 17083 27999
rect 17083 27965 17092 27999
rect 17040 27956 17092 27965
rect 17224 27999 17276 28008
rect 17224 27965 17233 27999
rect 17233 27965 17267 27999
rect 17267 27965 17276 27999
rect 17224 27956 17276 27965
rect 15568 27888 15620 27940
rect 3884 27820 3936 27872
rect 9312 27863 9364 27872
rect 9312 27829 9321 27863
rect 9321 27829 9355 27863
rect 9355 27829 9364 27863
rect 9312 27820 9364 27829
rect 11612 27863 11664 27872
rect 11612 27829 11621 27863
rect 11621 27829 11655 27863
rect 11655 27829 11664 27863
rect 11612 27820 11664 27829
rect 14556 27820 14608 27872
rect 22836 28067 22888 28076
rect 22836 28033 22845 28067
rect 22845 28033 22879 28067
rect 22879 28033 22888 28067
rect 22836 28024 22888 28033
rect 24216 28024 24268 28076
rect 20352 27956 20404 28008
rect 22560 27999 22612 28008
rect 19432 27888 19484 27940
rect 20996 27888 21048 27940
rect 22560 27965 22569 27999
rect 22569 27965 22603 27999
rect 22603 27965 22612 27999
rect 22560 27956 22612 27965
rect 23756 27999 23808 28008
rect 23756 27965 23765 27999
rect 23765 27965 23799 27999
rect 23799 27965 23808 27999
rect 23756 27956 23808 27965
rect 24584 27999 24636 28008
rect 24032 27888 24084 27940
rect 24584 27965 24593 27999
rect 24593 27965 24627 27999
rect 24627 27965 24636 27999
rect 24584 27956 24636 27965
rect 26056 28024 26108 28076
rect 27252 28024 27304 28076
rect 26240 27956 26292 28008
rect 29644 27999 29696 28008
rect 24676 27888 24728 27940
rect 27620 27888 27672 27940
rect 29644 27965 29653 27999
rect 29653 27965 29687 27999
rect 29687 27965 29696 27999
rect 29644 27956 29696 27965
rect 30380 27956 30432 28008
rect 30748 27956 30800 28008
rect 30932 27956 30984 28008
rect 33140 28024 33192 28076
rect 32956 27999 33008 28008
rect 29368 27888 29420 27940
rect 32956 27965 32965 27999
rect 32965 27965 32999 27999
rect 32999 27965 33008 27999
rect 32956 27956 33008 27965
rect 33232 27999 33284 28008
rect 33232 27965 33241 27999
rect 33241 27965 33275 27999
rect 33275 27965 33284 27999
rect 33232 27956 33284 27965
rect 33600 27999 33652 28008
rect 33600 27965 33609 27999
rect 33609 27965 33643 27999
rect 33643 27965 33652 27999
rect 33600 27956 33652 27965
rect 34520 27956 34572 28008
rect 35348 28024 35400 28076
rect 38292 28092 38344 28144
rect 37924 28024 37976 28076
rect 38844 28024 38896 28076
rect 35532 27956 35584 28008
rect 37096 27956 37148 28008
rect 38476 27999 38528 28008
rect 38476 27965 38485 27999
rect 38485 27965 38519 27999
rect 38519 27965 38528 27999
rect 38476 27956 38528 27965
rect 38752 27999 38804 28008
rect 38752 27965 38761 27999
rect 38761 27965 38795 27999
rect 38795 27965 38804 27999
rect 38752 27956 38804 27965
rect 34060 27888 34112 27940
rect 34336 27931 34388 27940
rect 34336 27897 34345 27931
rect 34345 27897 34379 27931
rect 34379 27897 34388 27931
rect 34336 27888 34388 27897
rect 24400 27820 24452 27872
rect 31300 27863 31352 27872
rect 31300 27829 31309 27863
rect 31309 27829 31343 27863
rect 31343 27829 31352 27863
rect 31300 27820 31352 27829
rect 19606 27718 19658 27770
rect 19670 27718 19722 27770
rect 19734 27718 19786 27770
rect 19798 27718 19850 27770
rect 2964 27659 3016 27668
rect 2964 27625 2973 27659
rect 2973 27625 3007 27659
rect 3007 27625 3016 27659
rect 2964 27616 3016 27625
rect 2688 27548 2740 27600
rect 7104 27616 7156 27668
rect 8208 27616 8260 27668
rect 1400 27523 1452 27532
rect 1400 27489 1409 27523
rect 1409 27489 1443 27523
rect 1443 27489 1452 27523
rect 1400 27480 1452 27489
rect 2412 27480 2464 27532
rect 4620 27480 4672 27532
rect 2780 27412 2832 27464
rect 5080 27412 5132 27464
rect 7564 27480 7616 27532
rect 8668 27523 8720 27532
rect 8668 27489 8677 27523
rect 8677 27489 8711 27523
rect 8711 27489 8720 27523
rect 8668 27480 8720 27489
rect 9128 27523 9180 27532
rect 9128 27489 9137 27523
rect 9137 27489 9171 27523
rect 9171 27489 9180 27523
rect 9128 27480 9180 27489
rect 6828 27412 6880 27464
rect 7380 27412 7432 27464
rect 9680 27412 9732 27464
rect 10416 27523 10468 27532
rect 10416 27489 10425 27523
rect 10425 27489 10459 27523
rect 10459 27489 10468 27523
rect 10416 27480 10468 27489
rect 11152 27480 11204 27532
rect 11612 27480 11664 27532
rect 13636 27480 13688 27532
rect 14004 27548 14056 27600
rect 18328 27616 18380 27668
rect 19064 27659 19116 27668
rect 19064 27625 19073 27659
rect 19073 27625 19107 27659
rect 19107 27625 19116 27659
rect 19064 27616 19116 27625
rect 20628 27616 20680 27668
rect 20996 27616 21048 27668
rect 24676 27616 24728 27668
rect 33876 27659 33928 27668
rect 33876 27625 33885 27659
rect 33885 27625 33919 27659
rect 33919 27625 33928 27659
rect 33876 27616 33928 27625
rect 34520 27616 34572 27668
rect 36636 27616 36688 27668
rect 18144 27548 18196 27600
rect 23848 27591 23900 27600
rect 16120 27480 16172 27532
rect 17224 27480 17276 27532
rect 19156 27480 19208 27532
rect 10876 27412 10928 27464
rect 11428 27412 11480 27464
rect 15752 27412 15804 27464
rect 16396 27412 16448 27464
rect 19340 27480 19392 27532
rect 21640 27480 21692 27532
rect 22284 27523 22336 27532
rect 19892 27412 19944 27464
rect 22284 27489 22293 27523
rect 22293 27489 22327 27523
rect 22327 27489 22336 27523
rect 22284 27480 22336 27489
rect 22468 27523 22520 27532
rect 22468 27489 22477 27523
rect 22477 27489 22511 27523
rect 22511 27489 22520 27523
rect 22468 27480 22520 27489
rect 23020 27412 23072 27464
rect 23204 27412 23256 27464
rect 4068 27276 4120 27328
rect 6000 27276 6052 27328
rect 6460 27276 6512 27328
rect 8116 27276 8168 27328
rect 8392 27276 8444 27328
rect 13912 27344 13964 27396
rect 22928 27344 22980 27396
rect 12256 27276 12308 27328
rect 22836 27276 22888 27328
rect 23480 27276 23532 27328
rect 23848 27557 23857 27591
rect 23857 27557 23891 27591
rect 23891 27557 23900 27591
rect 23848 27548 23900 27557
rect 24032 27548 24084 27600
rect 24584 27548 24636 27600
rect 29368 27591 29420 27600
rect 29368 27557 29377 27591
rect 29377 27557 29411 27591
rect 29411 27557 29420 27591
rect 29368 27548 29420 27557
rect 30932 27591 30984 27600
rect 30932 27557 30941 27591
rect 30941 27557 30975 27591
rect 30975 27557 30984 27591
rect 30932 27548 30984 27557
rect 24400 27523 24452 27532
rect 24400 27489 24409 27523
rect 24409 27489 24443 27523
rect 24443 27489 24452 27523
rect 24400 27480 24452 27489
rect 24492 27480 24544 27532
rect 26608 27523 26660 27532
rect 26608 27489 26617 27523
rect 26617 27489 26651 27523
rect 26651 27489 26660 27523
rect 26608 27480 26660 27489
rect 27620 27480 27672 27532
rect 30748 27523 30800 27532
rect 27712 27455 27764 27464
rect 27712 27421 27721 27455
rect 27721 27421 27755 27455
rect 27755 27421 27764 27455
rect 27712 27412 27764 27421
rect 27988 27455 28040 27464
rect 27988 27421 27997 27455
rect 27997 27421 28031 27455
rect 28031 27421 28040 27455
rect 27988 27412 28040 27421
rect 30748 27489 30757 27523
rect 30757 27489 30791 27523
rect 30791 27489 30800 27523
rect 30748 27480 30800 27489
rect 31392 27523 31444 27532
rect 31392 27489 31401 27523
rect 31401 27489 31435 27523
rect 31435 27489 31444 27523
rect 31392 27480 31444 27489
rect 33232 27548 33284 27600
rect 35256 27548 35308 27600
rect 36728 27591 36780 27600
rect 32496 27523 32548 27532
rect 32496 27489 32505 27523
rect 32505 27489 32539 27523
rect 32539 27489 32548 27523
rect 32496 27480 32548 27489
rect 30380 27412 30432 27464
rect 31668 27412 31720 27464
rect 33048 27480 33100 27532
rect 34336 27523 34388 27532
rect 34336 27489 34345 27523
rect 34345 27489 34379 27523
rect 34379 27489 34388 27523
rect 34336 27480 34388 27489
rect 35348 27523 35400 27532
rect 35348 27489 35357 27523
rect 35357 27489 35391 27523
rect 35391 27489 35400 27523
rect 35348 27480 35400 27489
rect 36728 27557 36737 27591
rect 36737 27557 36771 27591
rect 36771 27557 36780 27591
rect 36728 27548 36780 27557
rect 37096 27591 37148 27600
rect 37096 27557 37105 27591
rect 37105 27557 37139 27591
rect 37139 27557 37148 27591
rect 37096 27548 37148 27557
rect 33600 27412 33652 27464
rect 34060 27412 34112 27464
rect 26240 27344 26292 27396
rect 23848 27276 23900 27328
rect 32220 27319 32272 27328
rect 32220 27285 32229 27319
rect 32229 27285 32263 27319
rect 32263 27285 32272 27319
rect 32220 27276 32272 27285
rect 33508 27344 33560 27396
rect 37924 27480 37976 27532
rect 36452 27412 36504 27464
rect 37188 27412 37240 27464
rect 35716 27276 35768 27328
rect 35808 27276 35860 27328
rect 37832 27319 37884 27328
rect 37832 27285 37841 27319
rect 37841 27285 37875 27319
rect 37875 27285 37884 27319
rect 37832 27276 37884 27285
rect 4246 27174 4298 27226
rect 4310 27174 4362 27226
rect 4374 27174 4426 27226
rect 4438 27174 4490 27226
rect 34966 27174 35018 27226
rect 35030 27174 35082 27226
rect 35094 27174 35146 27226
rect 35158 27174 35210 27226
rect 2320 27115 2372 27124
rect 2320 27081 2329 27115
rect 2329 27081 2363 27115
rect 2363 27081 2372 27115
rect 2320 27072 2372 27081
rect 8668 27072 8720 27124
rect 11336 27115 11388 27124
rect 11336 27081 11345 27115
rect 11345 27081 11379 27115
rect 11379 27081 11388 27115
rect 11336 27072 11388 27081
rect 12716 27072 12768 27124
rect 16396 27072 16448 27124
rect 21088 27115 21140 27124
rect 21088 27081 21097 27115
rect 21097 27081 21131 27115
rect 21131 27081 21140 27115
rect 21088 27072 21140 27081
rect 22928 27072 22980 27124
rect 24492 27115 24544 27124
rect 2964 27004 3016 27056
rect 4804 27004 4856 27056
rect 8576 27004 8628 27056
rect 3332 26936 3384 26988
rect 4712 26936 4764 26988
rect 2412 26911 2464 26920
rect 2412 26877 2421 26911
rect 2421 26877 2455 26911
rect 2455 26877 2464 26911
rect 2412 26868 2464 26877
rect 2872 26911 2924 26920
rect 2872 26877 2881 26911
rect 2881 26877 2915 26911
rect 2915 26877 2924 26911
rect 2872 26868 2924 26877
rect 3056 26911 3108 26920
rect 3056 26877 3065 26911
rect 3065 26877 3099 26911
rect 3099 26877 3108 26911
rect 3056 26868 3108 26877
rect 3884 26911 3936 26920
rect 3884 26877 3893 26911
rect 3893 26877 3927 26911
rect 3927 26877 3936 26911
rect 3884 26868 3936 26877
rect 4068 26911 4120 26920
rect 4068 26877 4077 26911
rect 4077 26877 4111 26911
rect 4111 26877 4120 26911
rect 4068 26868 4120 26877
rect 5540 26911 5592 26920
rect 5540 26877 5549 26911
rect 5549 26877 5583 26911
rect 5583 26877 5592 26911
rect 5540 26868 5592 26877
rect 7840 26911 7892 26920
rect 6184 26800 6236 26852
rect 4988 26775 5040 26784
rect 4988 26741 4997 26775
rect 4997 26741 5031 26775
rect 5031 26741 5040 26775
rect 4988 26732 5040 26741
rect 7840 26877 7849 26911
rect 7849 26877 7883 26911
rect 7883 26877 7892 26911
rect 7840 26868 7892 26877
rect 9312 26936 9364 26988
rect 14004 27004 14056 27056
rect 18144 27004 18196 27056
rect 20444 27004 20496 27056
rect 20628 27004 20680 27056
rect 24124 27047 24176 27056
rect 24124 27013 24133 27047
rect 24133 27013 24167 27047
rect 24167 27013 24176 27047
rect 24124 27004 24176 27013
rect 24492 27081 24501 27115
rect 24501 27081 24535 27115
rect 24535 27081 24544 27115
rect 24492 27072 24544 27081
rect 29276 27072 29328 27124
rect 30012 27072 30064 27124
rect 32496 27072 32548 27124
rect 33232 27072 33284 27124
rect 34520 27072 34572 27124
rect 35808 27072 35860 27124
rect 38844 27115 38896 27124
rect 38844 27081 38853 27115
rect 38853 27081 38887 27115
rect 38887 27081 38896 27115
rect 38844 27072 38896 27081
rect 10508 26911 10560 26920
rect 8116 26800 8168 26852
rect 10508 26877 10517 26911
rect 10517 26877 10551 26911
rect 10551 26877 10560 26911
rect 10508 26868 10560 26877
rect 12440 26911 12492 26920
rect 12440 26877 12449 26911
rect 12449 26877 12483 26911
rect 12483 26877 12492 26911
rect 13544 26911 13596 26920
rect 12440 26868 12492 26877
rect 13544 26877 13553 26911
rect 13553 26877 13587 26911
rect 13587 26877 13596 26911
rect 13544 26868 13596 26877
rect 13912 26868 13964 26920
rect 18972 26979 19024 26988
rect 18972 26945 18981 26979
rect 18981 26945 19015 26979
rect 19015 26945 19024 26979
rect 18972 26936 19024 26945
rect 15476 26868 15528 26920
rect 16120 26911 16172 26920
rect 16120 26877 16129 26911
rect 16129 26877 16163 26911
rect 16163 26877 16172 26911
rect 16120 26868 16172 26877
rect 11428 26800 11480 26852
rect 13820 26800 13872 26852
rect 16028 26800 16080 26852
rect 8852 26732 8904 26784
rect 10784 26732 10836 26784
rect 15568 26775 15620 26784
rect 15568 26741 15577 26775
rect 15577 26741 15611 26775
rect 15611 26741 15620 26775
rect 15568 26732 15620 26741
rect 16672 26868 16724 26920
rect 19064 26911 19116 26920
rect 19064 26877 19073 26911
rect 19073 26877 19107 26911
rect 19107 26877 19116 26911
rect 19064 26868 19116 26877
rect 19432 26868 19484 26920
rect 20536 26936 20588 26988
rect 20076 26911 20128 26920
rect 20076 26877 20085 26911
rect 20085 26877 20119 26911
rect 20119 26877 20128 26911
rect 20076 26868 20128 26877
rect 20444 26911 20496 26920
rect 20444 26877 20453 26911
rect 20453 26877 20487 26911
rect 20487 26877 20496 26911
rect 20444 26868 20496 26877
rect 20812 26868 20864 26920
rect 21916 26868 21968 26920
rect 22284 26911 22336 26920
rect 22284 26877 22293 26911
rect 22293 26877 22327 26911
rect 22327 26877 22336 26911
rect 22284 26868 22336 26877
rect 19984 26800 20036 26852
rect 22836 26868 22888 26920
rect 23848 26843 23900 26852
rect 23848 26809 23857 26843
rect 23857 26809 23891 26843
rect 23891 26809 23900 26843
rect 23848 26800 23900 26809
rect 17040 26732 17092 26784
rect 17500 26732 17552 26784
rect 18512 26732 18564 26784
rect 27988 26936 28040 26988
rect 25596 26911 25648 26920
rect 25596 26877 25605 26911
rect 25605 26877 25639 26911
rect 25639 26877 25648 26911
rect 25596 26868 25648 26877
rect 27804 26868 27856 26920
rect 28632 26936 28684 26988
rect 28540 26911 28592 26920
rect 28540 26877 28549 26911
rect 28549 26877 28583 26911
rect 28583 26877 28592 26911
rect 28540 26868 28592 26877
rect 29552 26911 29604 26920
rect 29552 26877 29561 26911
rect 29561 26877 29595 26911
rect 29595 26877 29604 26911
rect 29552 26868 29604 26877
rect 32312 26936 32364 26988
rect 34244 26936 34296 26988
rect 30840 26911 30892 26920
rect 30840 26877 30849 26911
rect 30849 26877 30883 26911
rect 30883 26877 30892 26911
rect 30840 26868 30892 26877
rect 31576 26911 31628 26920
rect 31576 26877 31585 26911
rect 31585 26877 31619 26911
rect 31619 26877 31628 26911
rect 31576 26868 31628 26877
rect 31852 26911 31904 26920
rect 31852 26877 31861 26911
rect 31861 26877 31895 26911
rect 31895 26877 31904 26911
rect 31852 26868 31904 26877
rect 33692 26911 33744 26920
rect 33692 26877 33701 26911
rect 33701 26877 33735 26911
rect 33735 26877 33744 26911
rect 33692 26868 33744 26877
rect 34796 26868 34848 26920
rect 36636 26868 36688 26920
rect 37464 26911 37516 26920
rect 37464 26877 37473 26911
rect 37473 26877 37507 26911
rect 37507 26877 37516 26911
rect 37464 26868 37516 26877
rect 25412 26732 25464 26784
rect 30104 26732 30156 26784
rect 33508 26732 33560 26784
rect 35808 26775 35860 26784
rect 35808 26741 35817 26775
rect 35817 26741 35851 26775
rect 35851 26741 35860 26775
rect 35808 26732 35860 26741
rect 19606 26630 19658 26682
rect 19670 26630 19722 26682
rect 19734 26630 19786 26682
rect 19798 26630 19850 26682
rect 7748 26528 7800 26580
rect 8760 26528 8812 26580
rect 9036 26528 9088 26580
rect 13820 26528 13872 26580
rect 14004 26528 14056 26580
rect 16212 26528 16264 26580
rect 1952 26503 2004 26512
rect 1952 26469 1961 26503
rect 1961 26469 1995 26503
rect 1995 26469 2004 26503
rect 1952 26460 2004 26469
rect 9128 26460 9180 26512
rect 12256 26460 12308 26512
rect 2412 26435 2464 26444
rect 2412 26401 2421 26435
rect 2421 26401 2455 26435
rect 2455 26401 2464 26435
rect 2412 26392 2464 26401
rect 2872 26435 2924 26444
rect 2872 26401 2881 26435
rect 2881 26401 2915 26435
rect 2915 26401 2924 26435
rect 2872 26392 2924 26401
rect 3976 26392 4028 26444
rect 4804 26435 4856 26444
rect 4804 26401 4813 26435
rect 4813 26401 4847 26435
rect 4847 26401 4856 26435
rect 4804 26392 4856 26401
rect 8208 26435 8260 26444
rect 8208 26401 8217 26435
rect 8217 26401 8251 26435
rect 8251 26401 8260 26435
rect 8208 26392 8260 26401
rect 8668 26392 8720 26444
rect 11060 26392 11112 26444
rect 11244 26435 11296 26444
rect 11244 26401 11253 26435
rect 11253 26401 11287 26435
rect 11287 26401 11296 26435
rect 11244 26392 11296 26401
rect 11428 26435 11480 26444
rect 11428 26401 11437 26435
rect 11437 26401 11471 26435
rect 11471 26401 11480 26435
rect 11428 26392 11480 26401
rect 11520 26392 11572 26444
rect 15384 26460 15436 26512
rect 2964 26324 3016 26376
rect 5080 26324 5132 26376
rect 5080 26188 5132 26240
rect 6828 26188 6880 26240
rect 10784 26324 10836 26376
rect 9772 26299 9824 26308
rect 9772 26265 9781 26299
rect 9781 26265 9815 26299
rect 9815 26265 9824 26299
rect 9772 26256 9824 26265
rect 11980 26299 12032 26308
rect 11980 26265 11989 26299
rect 11989 26265 12023 26299
rect 12023 26265 12032 26299
rect 11980 26256 12032 26265
rect 13268 26256 13320 26308
rect 20444 26528 20496 26580
rect 15292 26367 15344 26376
rect 15292 26333 15301 26367
rect 15301 26333 15335 26367
rect 15335 26333 15344 26367
rect 15292 26324 15344 26333
rect 15476 26256 15528 26308
rect 16948 26392 17000 26444
rect 17684 26392 17736 26444
rect 16028 26324 16080 26376
rect 16396 26256 16448 26308
rect 17500 26324 17552 26376
rect 18052 26367 18104 26376
rect 18052 26333 18061 26367
rect 18061 26333 18095 26367
rect 18095 26333 18104 26367
rect 18052 26324 18104 26333
rect 18328 26435 18380 26444
rect 18328 26401 18337 26435
rect 18337 26401 18371 26435
rect 18371 26401 18380 26435
rect 18328 26392 18380 26401
rect 18604 26392 18656 26444
rect 19064 26392 19116 26444
rect 20352 26503 20404 26512
rect 20352 26469 20361 26503
rect 20361 26469 20395 26503
rect 20395 26469 20404 26503
rect 20352 26460 20404 26469
rect 20812 26460 20864 26512
rect 19892 26435 19944 26444
rect 19892 26401 19901 26435
rect 19901 26401 19935 26435
rect 19935 26401 19944 26435
rect 19892 26392 19944 26401
rect 19984 26392 20036 26444
rect 21916 26392 21968 26444
rect 22836 26435 22888 26444
rect 18328 26256 18380 26308
rect 22100 26367 22152 26376
rect 22100 26333 22109 26367
rect 22109 26333 22143 26367
rect 22143 26333 22152 26367
rect 22836 26401 22845 26435
rect 22845 26401 22879 26435
rect 22879 26401 22888 26435
rect 22836 26392 22888 26401
rect 23480 26392 23532 26444
rect 24584 26528 24636 26580
rect 26608 26571 26660 26580
rect 26608 26537 26617 26571
rect 26617 26537 26651 26571
rect 26651 26537 26660 26571
rect 26608 26528 26660 26537
rect 37648 26528 37700 26580
rect 30840 26460 30892 26512
rect 24216 26435 24268 26444
rect 24216 26401 24225 26435
rect 24225 26401 24259 26435
rect 24259 26401 24268 26435
rect 24216 26392 24268 26401
rect 24952 26392 25004 26444
rect 26516 26435 26568 26444
rect 26516 26401 26525 26435
rect 26525 26401 26559 26435
rect 26559 26401 26568 26435
rect 26516 26392 26568 26401
rect 30564 26392 30616 26444
rect 32128 26392 32180 26444
rect 33324 26392 33376 26444
rect 33508 26435 33560 26444
rect 33508 26401 33517 26435
rect 33517 26401 33551 26435
rect 33551 26401 33560 26435
rect 33508 26392 33560 26401
rect 35532 26435 35584 26444
rect 35532 26401 35541 26435
rect 35541 26401 35575 26435
rect 35575 26401 35584 26435
rect 35532 26392 35584 26401
rect 35808 26435 35860 26444
rect 35808 26401 35817 26435
rect 35817 26401 35851 26435
rect 35851 26401 35860 26435
rect 35808 26392 35860 26401
rect 38016 26435 38068 26444
rect 38016 26401 38025 26435
rect 38025 26401 38059 26435
rect 38059 26401 38068 26435
rect 38016 26392 38068 26401
rect 39028 26392 39080 26444
rect 22100 26324 22152 26333
rect 7840 26188 7892 26240
rect 11428 26188 11480 26240
rect 18604 26188 18656 26240
rect 20076 26256 20128 26308
rect 24124 26324 24176 26376
rect 24400 26324 24452 26376
rect 23572 26256 23624 26308
rect 19432 26188 19484 26240
rect 23480 26188 23532 26240
rect 23848 26188 23900 26240
rect 24860 26231 24912 26240
rect 24860 26197 24869 26231
rect 24869 26197 24903 26231
rect 24903 26197 24912 26231
rect 24860 26188 24912 26197
rect 26148 26188 26200 26240
rect 27712 26256 27764 26308
rect 27988 26324 28040 26376
rect 29276 26324 29328 26376
rect 29644 26256 29696 26308
rect 30104 26256 30156 26308
rect 29184 26231 29236 26240
rect 29184 26197 29193 26231
rect 29193 26197 29227 26231
rect 29227 26197 29236 26231
rect 29184 26188 29236 26197
rect 29736 26188 29788 26240
rect 31576 26324 31628 26376
rect 31668 26256 31720 26308
rect 34612 26231 34664 26240
rect 34612 26197 34621 26231
rect 34621 26197 34655 26231
rect 34655 26197 34664 26231
rect 34612 26188 34664 26197
rect 36544 26188 36596 26240
rect 36728 26188 36780 26240
rect 4246 26086 4298 26138
rect 4310 26086 4362 26138
rect 4374 26086 4426 26138
rect 4438 26086 4490 26138
rect 34966 26086 35018 26138
rect 35030 26086 35082 26138
rect 35094 26086 35146 26138
rect 35158 26086 35210 26138
rect 4620 25984 4672 26036
rect 2780 25848 2832 25900
rect 10968 25916 11020 25968
rect 11060 25916 11112 25968
rect 11244 25916 11296 25968
rect 22468 25984 22520 26036
rect 25504 25984 25556 26036
rect 25780 25984 25832 26036
rect 32128 25984 32180 26036
rect 35624 25984 35676 26036
rect 39120 25984 39172 26036
rect 4160 25780 4212 25832
rect 4620 25780 4672 25832
rect 5724 25823 5776 25832
rect 5724 25789 5733 25823
rect 5733 25789 5767 25823
rect 5767 25789 5776 25823
rect 5724 25780 5776 25789
rect 7104 25823 7156 25832
rect 7104 25789 7113 25823
rect 7113 25789 7147 25823
rect 7147 25789 7156 25823
rect 7104 25780 7156 25789
rect 8208 25780 8260 25832
rect 8668 25823 8720 25832
rect 8668 25789 8677 25823
rect 8677 25789 8711 25823
rect 8711 25789 8720 25823
rect 8668 25780 8720 25789
rect 9404 25823 9456 25832
rect 7472 25712 7524 25764
rect 4068 25644 4120 25696
rect 5816 25644 5868 25696
rect 7656 25644 7708 25696
rect 8024 25644 8076 25696
rect 8576 25712 8628 25764
rect 9404 25789 9413 25823
rect 9413 25789 9447 25823
rect 9447 25789 9456 25823
rect 9404 25780 9456 25789
rect 11980 25848 12032 25900
rect 13084 25848 13136 25900
rect 10876 25823 10928 25832
rect 10876 25789 10885 25823
rect 10885 25789 10919 25823
rect 10919 25789 10928 25823
rect 10876 25780 10928 25789
rect 10968 25644 11020 25696
rect 12532 25780 12584 25832
rect 13820 25823 13872 25832
rect 13820 25789 13829 25823
rect 13829 25789 13863 25823
rect 13863 25789 13872 25823
rect 13820 25780 13872 25789
rect 14280 25823 14332 25832
rect 14280 25789 14289 25823
rect 14289 25789 14323 25823
rect 14323 25789 14332 25823
rect 14280 25780 14332 25789
rect 14556 25823 14608 25832
rect 14556 25789 14565 25823
rect 14565 25789 14599 25823
rect 14599 25789 14608 25823
rect 14556 25780 14608 25789
rect 15292 25823 15344 25832
rect 15292 25789 15301 25823
rect 15301 25789 15335 25823
rect 15335 25789 15344 25823
rect 15292 25780 15344 25789
rect 15752 25780 15804 25832
rect 16120 25823 16172 25832
rect 16120 25789 16129 25823
rect 16129 25789 16163 25823
rect 16163 25789 16172 25823
rect 16120 25780 16172 25789
rect 16948 25823 17000 25832
rect 16948 25789 16957 25823
rect 16957 25789 16991 25823
rect 16991 25789 17000 25823
rect 16948 25780 17000 25789
rect 17684 25780 17736 25832
rect 19340 25848 19392 25900
rect 19984 25848 20036 25900
rect 21364 25891 21416 25900
rect 21364 25857 21373 25891
rect 21373 25857 21407 25891
rect 21407 25857 21416 25891
rect 21364 25848 21416 25857
rect 22100 25891 22152 25900
rect 22100 25857 22109 25891
rect 22109 25857 22143 25891
rect 22143 25857 22152 25891
rect 22100 25848 22152 25857
rect 18696 25823 18748 25832
rect 18696 25789 18705 25823
rect 18705 25789 18739 25823
rect 18739 25789 18748 25823
rect 19156 25823 19208 25832
rect 18696 25780 18748 25789
rect 19156 25789 19165 25823
rect 19165 25789 19199 25823
rect 19199 25789 19208 25823
rect 19156 25780 19208 25789
rect 19616 25780 19668 25832
rect 19892 25780 19944 25832
rect 20444 25823 20496 25832
rect 20444 25789 20453 25823
rect 20453 25789 20487 25823
rect 20487 25789 20496 25823
rect 20444 25780 20496 25789
rect 21180 25823 21232 25832
rect 11428 25712 11480 25764
rect 13176 25755 13228 25764
rect 13176 25721 13185 25755
rect 13185 25721 13219 25755
rect 13219 25721 13228 25755
rect 13176 25712 13228 25721
rect 18052 25712 18104 25764
rect 19708 25712 19760 25764
rect 19984 25712 20036 25764
rect 21180 25789 21189 25823
rect 21189 25789 21223 25823
rect 21223 25789 21232 25823
rect 21180 25780 21232 25789
rect 31852 25959 31904 25968
rect 31852 25925 31861 25959
rect 31861 25925 31895 25959
rect 31895 25925 31904 25959
rect 31852 25916 31904 25925
rect 24676 25891 24728 25900
rect 24676 25857 24685 25891
rect 24685 25857 24719 25891
rect 24719 25857 24728 25891
rect 24676 25848 24728 25857
rect 25228 25848 25280 25900
rect 26148 25848 26200 25900
rect 29644 25891 29696 25900
rect 29644 25857 29653 25891
rect 29653 25857 29687 25891
rect 29687 25857 29696 25891
rect 29644 25848 29696 25857
rect 23664 25823 23716 25832
rect 23664 25789 23673 25823
rect 23673 25789 23707 25823
rect 23707 25789 23716 25823
rect 23664 25780 23716 25789
rect 24584 25823 24636 25832
rect 24584 25789 24593 25823
rect 24593 25789 24627 25823
rect 24627 25789 24636 25823
rect 24584 25780 24636 25789
rect 25320 25780 25372 25832
rect 26700 25823 26752 25832
rect 26700 25789 26709 25823
rect 26709 25789 26743 25823
rect 26743 25789 26752 25823
rect 26700 25780 26752 25789
rect 29184 25780 29236 25832
rect 32312 25848 32364 25900
rect 35532 25848 35584 25900
rect 37464 25891 37516 25900
rect 37464 25857 37473 25891
rect 37473 25857 37507 25891
rect 37507 25857 37516 25891
rect 37464 25848 37516 25857
rect 37832 25848 37884 25900
rect 32220 25823 32272 25832
rect 25136 25712 25188 25764
rect 28080 25755 28132 25764
rect 28080 25721 28089 25755
rect 28089 25721 28123 25755
rect 28123 25721 28132 25755
rect 28080 25712 28132 25721
rect 13728 25644 13780 25696
rect 22560 25644 22612 25696
rect 28632 25687 28684 25696
rect 28632 25653 28641 25687
rect 28641 25653 28675 25687
rect 28675 25653 28684 25687
rect 28632 25644 28684 25653
rect 32220 25789 32229 25823
rect 32229 25789 32263 25823
rect 32263 25789 32272 25823
rect 32220 25780 32272 25789
rect 32496 25823 32548 25832
rect 32496 25789 32505 25823
rect 32505 25789 32539 25823
rect 32539 25789 32548 25823
rect 32496 25780 32548 25789
rect 30380 25712 30432 25764
rect 34060 25780 34112 25832
rect 35164 25823 35216 25832
rect 35164 25789 35173 25823
rect 35173 25789 35207 25823
rect 35207 25789 35216 25823
rect 35164 25780 35216 25789
rect 29644 25644 29696 25696
rect 19606 25542 19658 25594
rect 19670 25542 19722 25594
rect 19734 25542 19786 25594
rect 19798 25542 19850 25594
rect 2872 25440 2924 25492
rect 4160 25483 4212 25492
rect 4160 25449 4169 25483
rect 4169 25449 4203 25483
rect 4203 25449 4212 25483
rect 4160 25440 4212 25449
rect 4068 25372 4120 25424
rect 2780 25304 2832 25356
rect 2964 25304 3016 25356
rect 7012 25440 7064 25492
rect 16120 25440 16172 25492
rect 19340 25440 19392 25492
rect 19432 25440 19484 25492
rect 23480 25483 23532 25492
rect 23480 25449 23489 25483
rect 23489 25449 23523 25483
rect 23523 25449 23532 25483
rect 23480 25440 23532 25449
rect 26700 25440 26752 25492
rect 28080 25440 28132 25492
rect 8116 25415 8168 25424
rect 8116 25381 8125 25415
rect 8125 25381 8159 25415
rect 8159 25381 8168 25415
rect 8116 25372 8168 25381
rect 11152 25372 11204 25424
rect 11520 25415 11572 25424
rect 11520 25381 11529 25415
rect 11529 25381 11563 25415
rect 11563 25381 11572 25415
rect 11520 25372 11572 25381
rect 11980 25372 12032 25424
rect 19248 25415 19300 25424
rect 5816 25347 5868 25356
rect 1676 25279 1728 25288
rect 1676 25245 1685 25279
rect 1685 25245 1719 25279
rect 1719 25245 1728 25279
rect 1676 25236 1728 25245
rect 5816 25313 5825 25347
rect 5825 25313 5859 25347
rect 5859 25313 5868 25347
rect 5816 25304 5868 25313
rect 6092 25347 6144 25356
rect 6092 25313 6101 25347
rect 6101 25313 6135 25347
rect 6135 25313 6144 25347
rect 6828 25347 6880 25356
rect 6092 25304 6144 25313
rect 6828 25313 6837 25347
rect 6837 25313 6871 25347
rect 6871 25313 6880 25347
rect 6828 25304 6880 25313
rect 7564 25347 7616 25356
rect 7564 25313 7573 25347
rect 7573 25313 7607 25347
rect 7607 25313 7616 25347
rect 7564 25304 7616 25313
rect 8576 25347 8628 25356
rect 5080 25236 5132 25288
rect 5540 25279 5592 25288
rect 5540 25245 5549 25279
rect 5549 25245 5583 25279
rect 5583 25245 5592 25279
rect 5540 25236 5592 25245
rect 7104 25236 7156 25288
rect 7748 25236 7800 25288
rect 8576 25313 8585 25347
rect 8585 25313 8619 25347
rect 8619 25313 8628 25347
rect 8576 25304 8628 25313
rect 11060 25304 11112 25356
rect 12808 25347 12860 25356
rect 12808 25313 12817 25347
rect 12817 25313 12851 25347
rect 12851 25313 12860 25347
rect 12808 25304 12860 25313
rect 13268 25347 13320 25356
rect 13268 25313 13277 25347
rect 13277 25313 13311 25347
rect 13311 25313 13320 25347
rect 13268 25304 13320 25313
rect 13728 25304 13780 25356
rect 14556 25347 14608 25356
rect 14556 25313 14565 25347
rect 14565 25313 14599 25347
rect 14599 25313 14608 25347
rect 14556 25304 14608 25313
rect 15384 25347 15436 25356
rect 15384 25313 15393 25347
rect 15393 25313 15427 25347
rect 15427 25313 15436 25347
rect 15384 25304 15436 25313
rect 15476 25304 15528 25356
rect 19248 25381 19257 25415
rect 19257 25381 19291 25415
rect 19291 25381 19300 25415
rect 19248 25372 19300 25381
rect 20076 25372 20128 25424
rect 18236 25304 18288 25356
rect 19156 25304 19208 25356
rect 19432 25347 19484 25356
rect 19432 25313 19441 25347
rect 19441 25313 19475 25347
rect 19475 25313 19484 25347
rect 19432 25304 19484 25313
rect 20812 25304 20864 25356
rect 8484 25236 8536 25288
rect 11336 25236 11388 25288
rect 12624 25279 12676 25288
rect 12624 25245 12633 25279
rect 12633 25245 12667 25279
rect 12667 25245 12676 25279
rect 12624 25236 12676 25245
rect 18512 25236 18564 25288
rect 20444 25236 20496 25288
rect 21732 25347 21784 25356
rect 21732 25313 21741 25347
rect 21741 25313 21775 25347
rect 21775 25313 21784 25347
rect 22284 25347 22336 25356
rect 21732 25304 21784 25313
rect 22284 25313 22293 25347
rect 22293 25313 22327 25347
rect 22327 25313 22336 25347
rect 22284 25304 22336 25313
rect 22008 25236 22060 25288
rect 24860 25304 24912 25356
rect 25136 25347 25188 25356
rect 25136 25313 25145 25347
rect 25145 25313 25179 25347
rect 25179 25313 25188 25347
rect 25136 25304 25188 25313
rect 26516 25372 26568 25424
rect 29276 25415 29328 25424
rect 26608 25347 26660 25356
rect 26608 25313 26617 25347
rect 26617 25313 26651 25347
rect 26651 25313 26660 25347
rect 26608 25304 26660 25313
rect 29276 25381 29285 25415
rect 29285 25381 29319 25415
rect 29319 25381 29328 25415
rect 29276 25372 29328 25381
rect 28908 25304 28960 25356
rect 29920 25347 29972 25356
rect 29920 25313 29929 25347
rect 29929 25313 29963 25347
rect 29963 25313 29972 25347
rect 29920 25304 29972 25313
rect 30012 25279 30064 25288
rect 30012 25245 30021 25279
rect 30021 25245 30055 25279
rect 30055 25245 30064 25279
rect 30012 25236 30064 25245
rect 30380 25279 30432 25288
rect 30380 25245 30389 25279
rect 30389 25245 30423 25279
rect 30423 25245 30432 25279
rect 30380 25236 30432 25245
rect 31024 25304 31076 25356
rect 32496 25347 32548 25356
rect 32496 25313 32505 25347
rect 32505 25313 32539 25347
rect 32539 25313 32548 25347
rect 32496 25304 32548 25313
rect 33600 25440 33652 25492
rect 34060 25440 34112 25492
rect 34612 25372 34664 25424
rect 35164 25372 35216 25424
rect 38200 25415 38252 25424
rect 38200 25381 38209 25415
rect 38209 25381 38243 25415
rect 38243 25381 38252 25415
rect 38200 25372 38252 25381
rect 33324 25347 33376 25356
rect 33324 25313 33333 25347
rect 33333 25313 33367 25347
rect 33367 25313 33376 25347
rect 33324 25304 33376 25313
rect 34336 25304 34388 25356
rect 34796 25304 34848 25356
rect 35440 25304 35492 25356
rect 35624 25304 35676 25356
rect 36544 25347 36596 25356
rect 36544 25313 36553 25347
rect 36553 25313 36587 25347
rect 36587 25313 36596 25347
rect 36544 25304 36596 25313
rect 36636 25304 36688 25356
rect 38292 25347 38344 25356
rect 38292 25313 38301 25347
rect 38301 25313 38335 25347
rect 38335 25313 38344 25347
rect 38292 25304 38344 25313
rect 33416 25236 33468 25288
rect 38752 25279 38804 25288
rect 38752 25245 38761 25279
rect 38761 25245 38795 25279
rect 38795 25245 38804 25279
rect 38752 25236 38804 25245
rect 3976 25168 4028 25220
rect 7196 25168 7248 25220
rect 8392 25168 8444 25220
rect 8576 25168 8628 25220
rect 30564 25168 30616 25220
rect 31116 25211 31168 25220
rect 31116 25177 31125 25211
rect 31125 25177 31159 25211
rect 31159 25177 31168 25211
rect 31116 25168 31168 25177
rect 36912 25211 36964 25220
rect 36912 25177 36921 25211
rect 36921 25177 36955 25211
rect 36955 25177 36964 25211
rect 36912 25168 36964 25177
rect 14372 25100 14424 25152
rect 23756 25100 23808 25152
rect 25320 25100 25372 25152
rect 29000 25100 29052 25152
rect 36544 25100 36596 25152
rect 4246 24998 4298 25050
rect 4310 24998 4362 25050
rect 4374 24998 4426 25050
rect 4438 24998 4490 25050
rect 34966 24998 35018 25050
rect 35030 24998 35082 25050
rect 35094 24998 35146 25050
rect 35158 24998 35210 25050
rect 2780 24828 2832 24880
rect 3424 24828 3476 24880
rect 5724 24896 5776 24948
rect 2872 24760 2924 24812
rect 8208 24828 8260 24880
rect 4988 24760 5040 24812
rect 7012 24760 7064 24812
rect 1584 24735 1636 24744
rect 1584 24701 1593 24735
rect 1593 24701 1627 24735
rect 1627 24701 1636 24735
rect 1584 24692 1636 24701
rect 2228 24735 2280 24744
rect 2228 24701 2237 24735
rect 2237 24701 2271 24735
rect 2271 24701 2280 24735
rect 2228 24692 2280 24701
rect 2688 24692 2740 24744
rect 2964 24735 3016 24744
rect 2964 24701 2973 24735
rect 2973 24701 3007 24735
rect 3007 24701 3016 24735
rect 2964 24692 3016 24701
rect 7380 24692 7432 24744
rect 6276 24624 6328 24676
rect 7564 24692 7616 24744
rect 7656 24692 7708 24744
rect 8116 24692 8168 24744
rect 8392 24692 8444 24744
rect 9864 24760 9916 24812
rect 11520 24828 11572 24880
rect 13820 24871 13872 24880
rect 13820 24837 13829 24871
rect 13829 24837 13863 24871
rect 13863 24837 13872 24871
rect 13820 24828 13872 24837
rect 11336 24760 11388 24812
rect 15384 24896 15436 24948
rect 18512 24939 18564 24948
rect 18512 24905 18521 24939
rect 18521 24905 18555 24939
rect 18555 24905 18564 24939
rect 18512 24896 18564 24905
rect 24400 24896 24452 24948
rect 25504 24896 25556 24948
rect 26516 24939 26568 24948
rect 26516 24905 26525 24939
rect 26525 24905 26559 24939
rect 26559 24905 26568 24939
rect 26516 24896 26568 24905
rect 16212 24828 16264 24880
rect 16764 24803 16816 24812
rect 9772 24735 9824 24744
rect 9772 24701 9781 24735
rect 9781 24701 9815 24735
rect 9815 24701 9824 24735
rect 9772 24692 9824 24701
rect 9956 24735 10008 24744
rect 9956 24701 9965 24735
rect 9965 24701 9999 24735
rect 9999 24701 10008 24735
rect 9956 24692 10008 24701
rect 11060 24735 11112 24744
rect 11060 24701 11069 24735
rect 11069 24701 11103 24735
rect 11103 24701 11112 24735
rect 11060 24692 11112 24701
rect 11428 24735 11480 24744
rect 2412 24556 2464 24608
rect 5816 24556 5868 24608
rect 10232 24624 10284 24676
rect 8116 24556 8168 24608
rect 10508 24556 10560 24608
rect 11428 24701 11437 24735
rect 11437 24701 11471 24735
rect 11471 24701 11480 24735
rect 11428 24692 11480 24701
rect 11520 24692 11572 24744
rect 11888 24624 11940 24676
rect 14556 24692 14608 24744
rect 15476 24624 15528 24676
rect 12440 24556 12492 24608
rect 15660 24556 15712 24608
rect 16396 24692 16448 24744
rect 16764 24769 16773 24803
rect 16773 24769 16807 24803
rect 16807 24769 16816 24803
rect 16764 24760 16816 24769
rect 18052 24803 18104 24812
rect 18052 24769 18061 24803
rect 18061 24769 18095 24803
rect 18095 24769 18104 24803
rect 18052 24760 18104 24769
rect 16672 24735 16724 24744
rect 16672 24701 16681 24735
rect 16681 24701 16715 24735
rect 16715 24701 16724 24735
rect 16672 24692 16724 24701
rect 17500 24692 17552 24744
rect 18144 24624 18196 24676
rect 18236 24667 18288 24676
rect 18236 24633 18245 24667
rect 18245 24633 18279 24667
rect 18279 24633 18288 24667
rect 18236 24624 18288 24633
rect 20812 24828 20864 24880
rect 21088 24760 21140 24812
rect 20812 24735 20864 24744
rect 20812 24701 20821 24735
rect 20821 24701 20855 24735
rect 20855 24701 20864 24735
rect 20812 24692 20864 24701
rect 22192 24828 22244 24880
rect 29920 24828 29972 24880
rect 23664 24760 23716 24812
rect 24216 24760 24268 24812
rect 25412 24803 25464 24812
rect 25412 24769 25421 24803
rect 25421 24769 25455 24803
rect 25455 24769 25464 24803
rect 25412 24760 25464 24769
rect 29184 24760 29236 24812
rect 22192 24735 22244 24744
rect 20720 24624 20772 24676
rect 19432 24556 19484 24608
rect 22192 24701 22201 24735
rect 22201 24701 22235 24735
rect 22235 24701 22244 24735
rect 22192 24692 22244 24701
rect 22928 24692 22980 24744
rect 23848 24692 23900 24744
rect 25136 24735 25188 24744
rect 25136 24701 25145 24735
rect 25145 24701 25179 24735
rect 25179 24701 25188 24735
rect 25136 24692 25188 24701
rect 28264 24735 28316 24744
rect 28264 24701 28273 24735
rect 28273 24701 28307 24735
rect 28307 24701 28316 24735
rect 28264 24692 28316 24701
rect 22284 24624 22336 24676
rect 26792 24624 26844 24676
rect 27620 24624 27672 24676
rect 28632 24692 28684 24744
rect 34612 24760 34664 24812
rect 34888 24760 34940 24812
rect 35440 24803 35492 24812
rect 35440 24769 35449 24803
rect 35449 24769 35483 24803
rect 35483 24769 35492 24803
rect 35440 24760 35492 24769
rect 37004 24760 37056 24812
rect 37464 24760 37516 24812
rect 38292 24760 38344 24812
rect 30656 24692 30708 24744
rect 30564 24624 30616 24676
rect 31024 24692 31076 24744
rect 31668 24735 31720 24744
rect 31668 24701 31677 24735
rect 31677 24701 31711 24735
rect 31711 24701 31720 24735
rect 31668 24692 31720 24701
rect 32220 24692 32272 24744
rect 32588 24735 32640 24744
rect 32588 24701 32597 24735
rect 32597 24701 32631 24735
rect 32631 24701 32640 24735
rect 32588 24692 32640 24701
rect 35256 24692 35308 24744
rect 35716 24692 35768 24744
rect 32404 24624 32456 24676
rect 33324 24624 33376 24676
rect 34520 24624 34572 24676
rect 35072 24624 35124 24676
rect 36360 24692 36412 24744
rect 37372 24692 37424 24744
rect 24308 24556 24360 24608
rect 30472 24556 30524 24608
rect 36360 24556 36412 24608
rect 36728 24599 36780 24608
rect 36728 24565 36737 24599
rect 36737 24565 36771 24599
rect 36771 24565 36780 24599
rect 36728 24556 36780 24565
rect 37924 24556 37976 24608
rect 19606 24454 19658 24506
rect 19670 24454 19722 24506
rect 19734 24454 19786 24506
rect 19798 24454 19850 24506
rect 15936 24395 15988 24404
rect 15936 24361 15945 24395
rect 15945 24361 15979 24395
rect 15979 24361 15988 24395
rect 15936 24352 15988 24361
rect 20720 24352 20772 24404
rect 22008 24352 22060 24404
rect 22100 24352 22152 24404
rect 1676 24284 1728 24336
rect 2412 24259 2464 24268
rect 2412 24225 2421 24259
rect 2421 24225 2455 24259
rect 2455 24225 2464 24259
rect 2412 24216 2464 24225
rect 2780 24216 2832 24268
rect 2964 24216 3016 24268
rect 4528 24216 4580 24268
rect 5540 24216 5592 24268
rect 6276 24259 6328 24268
rect 5816 24148 5868 24200
rect 6276 24225 6285 24259
rect 6285 24225 6319 24259
rect 6319 24225 6328 24259
rect 6276 24216 6328 24225
rect 7012 24259 7064 24268
rect 7012 24225 7021 24259
rect 7021 24225 7055 24259
rect 7055 24225 7064 24259
rect 7012 24216 7064 24225
rect 7748 24259 7800 24268
rect 6184 24191 6236 24200
rect 6184 24157 6193 24191
rect 6193 24157 6227 24191
rect 6227 24157 6236 24191
rect 6184 24148 6236 24157
rect 7472 24080 7524 24132
rect 3700 24012 3752 24064
rect 7748 24225 7757 24259
rect 7757 24225 7791 24259
rect 7791 24225 7800 24259
rect 7748 24216 7800 24225
rect 8208 24216 8260 24268
rect 12992 24284 13044 24336
rect 16212 24284 16264 24336
rect 8484 24216 8536 24268
rect 10324 24259 10376 24268
rect 9404 24148 9456 24200
rect 9864 24148 9916 24200
rect 10324 24225 10333 24259
rect 10333 24225 10367 24259
rect 10367 24225 10376 24259
rect 10324 24216 10376 24225
rect 10508 24259 10560 24268
rect 10508 24225 10517 24259
rect 10517 24225 10551 24259
rect 10551 24225 10560 24259
rect 10508 24216 10560 24225
rect 11152 24259 11204 24268
rect 11152 24225 11161 24259
rect 11161 24225 11195 24259
rect 11195 24225 11204 24259
rect 11152 24216 11204 24225
rect 11612 24216 11664 24268
rect 9956 24123 10008 24132
rect 9956 24089 9965 24123
rect 9965 24089 9999 24123
rect 9999 24089 10008 24123
rect 9956 24080 10008 24089
rect 10232 24148 10284 24200
rect 14372 24216 14424 24268
rect 14464 24216 14516 24268
rect 15476 24216 15528 24268
rect 16028 24216 16080 24268
rect 17132 24284 17184 24336
rect 17224 24216 17276 24268
rect 18236 24259 18288 24268
rect 18236 24225 18245 24259
rect 18245 24225 18279 24259
rect 18279 24225 18288 24259
rect 18236 24216 18288 24225
rect 18512 24284 18564 24336
rect 22744 24284 22796 24336
rect 23020 24327 23072 24336
rect 23020 24293 23029 24327
rect 23029 24293 23063 24327
rect 23063 24293 23072 24327
rect 23020 24284 23072 24293
rect 10968 24080 11020 24132
rect 12624 24080 12676 24132
rect 8392 24012 8444 24064
rect 8760 24055 8812 24064
rect 8760 24021 8769 24055
rect 8769 24021 8803 24055
rect 8803 24021 8812 24055
rect 8760 24012 8812 24021
rect 10324 24012 10376 24064
rect 14740 24191 14792 24200
rect 14740 24157 14749 24191
rect 14749 24157 14783 24191
rect 14783 24157 14792 24191
rect 14740 24148 14792 24157
rect 19892 24216 19944 24268
rect 20076 24259 20128 24268
rect 20076 24225 20085 24259
rect 20085 24225 20119 24259
rect 20119 24225 20128 24259
rect 20076 24216 20128 24225
rect 21640 24259 21692 24268
rect 21640 24225 21649 24259
rect 21649 24225 21683 24259
rect 21683 24225 21692 24259
rect 21640 24216 21692 24225
rect 21732 24216 21784 24268
rect 23296 24216 23348 24268
rect 23756 24259 23808 24268
rect 23756 24225 23765 24259
rect 23765 24225 23799 24259
rect 23799 24225 23808 24259
rect 24032 24259 24084 24268
rect 23756 24216 23808 24225
rect 24032 24225 24041 24259
rect 24041 24225 24075 24259
rect 24075 24225 24084 24259
rect 24032 24216 24084 24225
rect 25688 24352 25740 24404
rect 27344 24352 27396 24404
rect 28540 24352 28592 24404
rect 24860 24259 24912 24268
rect 24860 24225 24869 24259
rect 24869 24225 24903 24259
rect 24903 24225 24912 24259
rect 24860 24216 24912 24225
rect 25320 24216 25372 24268
rect 28908 24284 28960 24336
rect 25780 24259 25832 24268
rect 25780 24225 25789 24259
rect 25789 24225 25823 24259
rect 25823 24225 25832 24259
rect 25780 24216 25832 24225
rect 27344 24259 27396 24268
rect 27344 24225 27353 24259
rect 27353 24225 27387 24259
rect 27387 24225 27396 24259
rect 27344 24216 27396 24225
rect 27620 24259 27672 24268
rect 27620 24225 27629 24259
rect 27629 24225 27663 24259
rect 27663 24225 27672 24259
rect 27620 24216 27672 24225
rect 29184 24216 29236 24268
rect 30840 24352 30892 24404
rect 35900 24352 35952 24404
rect 37280 24352 37332 24404
rect 30012 24284 30064 24336
rect 29368 24191 29420 24200
rect 14464 24012 14516 24064
rect 14556 24012 14608 24064
rect 16672 24080 16724 24132
rect 18052 24123 18104 24132
rect 18052 24089 18061 24123
rect 18061 24089 18095 24123
rect 18095 24089 18104 24123
rect 18052 24080 18104 24089
rect 18144 24080 18196 24132
rect 19340 24080 19392 24132
rect 20628 24080 20680 24132
rect 21180 24123 21232 24132
rect 21180 24089 21189 24123
rect 21189 24089 21223 24123
rect 21223 24089 21232 24123
rect 21180 24080 21232 24089
rect 21640 24080 21692 24132
rect 25964 24080 26016 24132
rect 17316 24012 17368 24064
rect 17684 24012 17736 24064
rect 22836 24012 22888 24064
rect 23204 24012 23256 24064
rect 29368 24157 29377 24191
rect 29377 24157 29411 24191
rect 29411 24157 29420 24191
rect 29368 24148 29420 24157
rect 30472 24259 30524 24268
rect 29920 24148 29972 24200
rect 30472 24225 30481 24259
rect 30481 24225 30515 24259
rect 30515 24225 30524 24259
rect 30472 24216 30524 24225
rect 30656 24216 30708 24268
rect 32496 24259 32548 24268
rect 32496 24225 32505 24259
rect 32505 24225 32539 24259
rect 32539 24225 32548 24259
rect 32496 24216 32548 24225
rect 33324 24259 33376 24268
rect 32588 24191 32640 24200
rect 32588 24157 32597 24191
rect 32597 24157 32631 24191
rect 32631 24157 32640 24191
rect 32588 24148 32640 24157
rect 33324 24225 33333 24259
rect 33333 24225 33367 24259
rect 33367 24225 33376 24259
rect 33324 24216 33376 24225
rect 33600 24259 33652 24268
rect 33600 24225 33609 24259
rect 33609 24225 33643 24259
rect 33643 24225 33652 24259
rect 33600 24216 33652 24225
rect 34888 24284 34940 24336
rect 36084 24284 36136 24336
rect 38200 24284 38252 24336
rect 35072 24259 35124 24268
rect 35072 24225 35081 24259
rect 35081 24225 35115 24259
rect 35115 24225 35124 24259
rect 35072 24216 35124 24225
rect 35348 24216 35400 24268
rect 35532 24216 35584 24268
rect 37004 24216 37056 24268
rect 37832 24259 37884 24268
rect 37832 24225 37841 24259
rect 37841 24225 37875 24259
rect 37875 24225 37884 24259
rect 37832 24216 37884 24225
rect 38292 24259 38344 24268
rect 38292 24225 38301 24259
rect 38301 24225 38335 24259
rect 38335 24225 38344 24259
rect 38292 24216 38344 24225
rect 34520 24148 34572 24200
rect 33600 24080 33652 24132
rect 30840 24012 30892 24064
rect 31024 24012 31076 24064
rect 32220 24012 32272 24064
rect 34336 24012 34388 24064
rect 36360 24055 36412 24064
rect 36360 24021 36369 24055
rect 36369 24021 36403 24055
rect 36403 24021 36412 24055
rect 36360 24012 36412 24021
rect 4246 23910 4298 23962
rect 4310 23910 4362 23962
rect 4374 23910 4426 23962
rect 4438 23910 4490 23962
rect 34966 23910 35018 23962
rect 35030 23910 35082 23962
rect 35094 23910 35146 23962
rect 35158 23910 35210 23962
rect 5632 23783 5684 23792
rect 5632 23749 5641 23783
rect 5641 23749 5675 23783
rect 5675 23749 5684 23783
rect 5632 23740 5684 23749
rect 2780 23715 2832 23724
rect 2780 23681 2789 23715
rect 2789 23681 2823 23715
rect 2823 23681 2832 23715
rect 3424 23715 3476 23724
rect 2780 23672 2832 23681
rect 3424 23681 3433 23715
rect 3433 23681 3467 23715
rect 3467 23681 3476 23715
rect 3424 23672 3476 23681
rect 3700 23715 3752 23724
rect 3700 23681 3709 23715
rect 3709 23681 3743 23715
rect 3743 23681 3752 23715
rect 3700 23672 3752 23681
rect 8208 23808 8260 23860
rect 11244 23740 11296 23792
rect 11428 23740 11480 23792
rect 2044 23647 2096 23656
rect 2044 23613 2053 23647
rect 2053 23613 2087 23647
rect 2087 23613 2096 23647
rect 2044 23604 2096 23613
rect 2412 23647 2464 23656
rect 2412 23613 2421 23647
rect 2421 23613 2455 23647
rect 2455 23613 2464 23647
rect 2412 23604 2464 23613
rect 5724 23647 5776 23656
rect 5724 23613 5733 23647
rect 5733 23613 5767 23647
rect 5767 23613 5776 23647
rect 5724 23604 5776 23613
rect 6828 23604 6880 23656
rect 8392 23647 8444 23656
rect 4712 23468 4764 23520
rect 4988 23511 5040 23520
rect 4988 23477 4997 23511
rect 4997 23477 5031 23511
rect 5031 23477 5040 23511
rect 4988 23468 5040 23477
rect 8392 23613 8401 23647
rect 8401 23613 8435 23647
rect 8435 23613 8444 23647
rect 8392 23604 8444 23613
rect 10508 23672 10560 23724
rect 11796 23672 11848 23724
rect 14740 23808 14792 23860
rect 15660 23808 15712 23860
rect 17316 23808 17368 23860
rect 19340 23808 19392 23860
rect 22928 23851 22980 23860
rect 22928 23817 22937 23851
rect 22937 23817 22971 23851
rect 22971 23817 22980 23851
rect 22928 23808 22980 23817
rect 23572 23808 23624 23860
rect 18236 23740 18288 23792
rect 19984 23740 20036 23792
rect 21640 23740 21692 23792
rect 21824 23740 21876 23792
rect 25596 23740 25648 23792
rect 30656 23740 30708 23792
rect 8208 23536 8260 23588
rect 8484 23536 8536 23588
rect 9864 23647 9916 23656
rect 9864 23613 9873 23647
rect 9873 23613 9907 23647
rect 9907 23613 9916 23647
rect 9864 23604 9916 23613
rect 10324 23647 10376 23656
rect 10324 23613 10333 23647
rect 10333 23613 10367 23647
rect 10367 23613 10376 23647
rect 10324 23604 10376 23613
rect 10784 23604 10836 23656
rect 11704 23647 11756 23656
rect 11704 23613 11713 23647
rect 11713 23613 11747 23647
rect 11747 23613 11756 23647
rect 11704 23604 11756 23613
rect 12716 23647 12768 23656
rect 9772 23536 9824 23588
rect 12716 23613 12725 23647
rect 12725 23613 12759 23647
rect 12759 23613 12768 23647
rect 12716 23604 12768 23613
rect 14556 23647 14608 23656
rect 14556 23613 14565 23647
rect 14565 23613 14599 23647
rect 14599 23613 14608 23647
rect 14556 23604 14608 23613
rect 15292 23647 15344 23656
rect 15292 23613 15301 23647
rect 15301 23613 15335 23647
rect 15335 23613 15344 23647
rect 15292 23604 15344 23613
rect 16120 23647 16172 23656
rect 16120 23613 16129 23647
rect 16129 23613 16163 23647
rect 16163 23613 16172 23647
rect 16120 23604 16172 23613
rect 18052 23647 18104 23656
rect 18052 23613 18061 23647
rect 18061 23613 18095 23647
rect 18095 23613 18104 23647
rect 18052 23604 18104 23613
rect 18880 23647 18932 23656
rect 16580 23536 16632 23588
rect 17500 23536 17552 23588
rect 18880 23613 18889 23647
rect 18889 23613 18923 23647
rect 18923 23613 18932 23647
rect 18880 23604 18932 23613
rect 20076 23604 20128 23656
rect 20720 23604 20772 23656
rect 21088 23604 21140 23656
rect 23388 23672 23440 23724
rect 25320 23715 25372 23724
rect 25320 23681 25329 23715
rect 25329 23681 25363 23715
rect 25363 23681 25372 23715
rect 25320 23672 25372 23681
rect 21640 23604 21692 23656
rect 23020 23604 23072 23656
rect 23848 23647 23900 23656
rect 23848 23613 23857 23647
rect 23857 23613 23891 23647
rect 23891 23613 23900 23647
rect 23848 23604 23900 23613
rect 20996 23536 21048 23588
rect 24860 23604 24912 23656
rect 30564 23672 30616 23724
rect 25688 23647 25740 23656
rect 25688 23613 25697 23647
rect 25697 23613 25731 23647
rect 25731 23613 25740 23647
rect 25688 23604 25740 23613
rect 25964 23647 26016 23656
rect 25964 23613 25973 23647
rect 25973 23613 26007 23647
rect 26007 23613 26016 23647
rect 25964 23604 26016 23613
rect 26976 23647 27028 23656
rect 26516 23536 26568 23588
rect 10324 23468 10376 23520
rect 14464 23468 14516 23520
rect 18236 23468 18288 23520
rect 19984 23468 20036 23520
rect 20168 23468 20220 23520
rect 20720 23468 20772 23520
rect 21364 23468 21416 23520
rect 21732 23468 21784 23520
rect 25136 23468 25188 23520
rect 26976 23613 26985 23647
rect 26985 23613 27019 23647
rect 27019 23613 27028 23647
rect 26976 23604 27028 23613
rect 30472 23604 30524 23656
rect 28356 23579 28408 23588
rect 28356 23545 28365 23579
rect 28365 23545 28399 23579
rect 28399 23545 28408 23579
rect 28356 23536 28408 23545
rect 29644 23536 29696 23588
rect 32956 23604 33008 23656
rect 33324 23647 33376 23656
rect 33324 23613 33333 23647
rect 33333 23613 33367 23647
rect 33367 23613 33376 23647
rect 33324 23604 33376 23613
rect 33784 23647 33836 23656
rect 33784 23613 33793 23647
rect 33793 23613 33827 23647
rect 33827 23613 33836 23647
rect 33784 23604 33836 23613
rect 37372 23808 37424 23860
rect 34428 23740 34480 23792
rect 35164 23740 35216 23792
rect 37004 23715 37056 23724
rect 37004 23681 37013 23715
rect 37013 23681 37047 23715
rect 37047 23681 37056 23715
rect 37004 23672 37056 23681
rect 37280 23715 37332 23724
rect 37280 23681 37289 23715
rect 37289 23681 37323 23715
rect 37323 23681 37332 23715
rect 37280 23672 37332 23681
rect 34244 23579 34296 23588
rect 27620 23468 27672 23520
rect 34244 23545 34253 23579
rect 34253 23545 34287 23579
rect 34287 23545 34296 23579
rect 34244 23536 34296 23545
rect 35532 23604 35584 23656
rect 36084 23647 36136 23656
rect 36084 23613 36093 23647
rect 36093 23613 36127 23647
rect 36127 23613 36136 23647
rect 36084 23604 36136 23613
rect 36268 23604 36320 23656
rect 36728 23604 36780 23656
rect 34520 23536 34572 23588
rect 35624 23536 35676 23588
rect 31024 23468 31076 23520
rect 31392 23468 31444 23520
rect 33324 23468 33376 23520
rect 33416 23468 33468 23520
rect 35440 23468 35492 23520
rect 19606 23366 19658 23418
rect 19670 23366 19722 23418
rect 19734 23366 19786 23418
rect 19798 23366 19850 23418
rect 5540 23264 5592 23316
rect 4896 23171 4948 23180
rect 4896 23137 4905 23171
rect 4905 23137 4939 23171
rect 4939 23137 4948 23171
rect 4896 23128 4948 23137
rect 6000 23196 6052 23248
rect 6092 23171 6144 23180
rect 1400 23103 1452 23112
rect 1400 23069 1409 23103
rect 1409 23069 1443 23103
rect 1443 23069 1452 23103
rect 1400 23060 1452 23069
rect 1768 23060 1820 23112
rect 3332 23060 3384 23112
rect 6092 23137 6101 23171
rect 6101 23137 6135 23171
rect 6135 23137 6144 23171
rect 6092 23128 6144 23137
rect 6184 23128 6236 23180
rect 10784 23264 10836 23316
rect 14004 23264 14056 23316
rect 16120 23264 16172 23316
rect 20996 23264 21048 23316
rect 23020 23264 23072 23316
rect 23204 23264 23256 23316
rect 7840 23171 7892 23180
rect 7840 23137 7849 23171
rect 7849 23137 7883 23171
rect 7883 23137 7892 23171
rect 7840 23128 7892 23137
rect 12624 23196 12676 23248
rect 15292 23239 15344 23248
rect 15292 23205 15301 23239
rect 15301 23205 15335 23239
rect 15335 23205 15344 23239
rect 15292 23196 15344 23205
rect 7288 23060 7340 23112
rect 4712 23035 4764 23044
rect 4712 23001 4721 23035
rect 4721 23001 4755 23035
rect 4755 23001 4764 23035
rect 4712 22992 4764 23001
rect 4988 22992 5040 23044
rect 10140 23128 10192 23180
rect 10324 23171 10376 23180
rect 10324 23137 10333 23171
rect 10333 23137 10367 23171
rect 10367 23137 10376 23171
rect 10324 23128 10376 23137
rect 10876 23171 10928 23180
rect 10876 23137 10885 23171
rect 10885 23137 10919 23171
rect 10919 23137 10928 23171
rect 10876 23128 10928 23137
rect 11244 23171 11296 23180
rect 11244 23137 11253 23171
rect 11253 23137 11287 23171
rect 11287 23137 11296 23171
rect 11244 23128 11296 23137
rect 11796 23128 11848 23180
rect 12164 23171 12216 23180
rect 12164 23137 12173 23171
rect 12173 23137 12207 23171
rect 12207 23137 12216 23171
rect 12164 23128 12216 23137
rect 12348 23128 12400 23180
rect 11060 23103 11112 23112
rect 11060 23069 11069 23103
rect 11069 23069 11103 23103
rect 11103 23069 11112 23103
rect 11060 23060 11112 23069
rect 14556 23128 14608 23180
rect 15660 23128 15712 23180
rect 15844 23128 15896 23180
rect 16672 23196 16724 23248
rect 16396 23128 16448 23180
rect 14004 23060 14056 23112
rect 14372 23060 14424 23112
rect 2964 22967 3016 22976
rect 2964 22933 2973 22967
rect 2973 22933 3007 22967
rect 3007 22933 3016 22967
rect 2964 22924 3016 22933
rect 3516 22924 3568 22976
rect 7104 22924 7156 22976
rect 10876 22924 10928 22976
rect 19248 23196 19300 23248
rect 18696 23171 18748 23180
rect 18328 23060 18380 23112
rect 18696 23137 18705 23171
rect 18705 23137 18739 23171
rect 18739 23137 18748 23171
rect 18696 23128 18748 23137
rect 21640 23196 21692 23248
rect 22008 23196 22060 23248
rect 20996 23171 21048 23180
rect 17592 22992 17644 23044
rect 20352 23060 20404 23112
rect 20996 23137 21005 23171
rect 21005 23137 21039 23171
rect 21039 23137 21048 23171
rect 20996 23128 21048 23137
rect 22928 23171 22980 23180
rect 22928 23137 22937 23171
rect 22937 23137 22971 23171
rect 22971 23137 22980 23171
rect 22928 23128 22980 23137
rect 26976 23196 27028 23248
rect 23664 23128 23716 23180
rect 23940 23128 23992 23180
rect 25688 23128 25740 23180
rect 21916 23103 21968 23112
rect 20260 22992 20312 23044
rect 21916 23069 21925 23103
rect 21925 23069 21959 23103
rect 21959 23069 21968 23103
rect 21916 23060 21968 23069
rect 22008 23060 22060 23112
rect 21824 23035 21876 23044
rect 21824 23001 21833 23035
rect 21833 23001 21867 23035
rect 21867 23001 21876 23035
rect 21824 22992 21876 23001
rect 23296 22992 23348 23044
rect 25044 23060 25096 23112
rect 16028 22924 16080 22976
rect 16304 22924 16356 22976
rect 26792 23128 26844 23180
rect 26240 23060 26292 23112
rect 29368 23264 29420 23316
rect 27896 23196 27948 23248
rect 27804 23128 27856 23180
rect 28264 23128 28316 23180
rect 28540 23196 28592 23248
rect 28448 23128 28500 23180
rect 28908 23128 28960 23180
rect 29920 23128 29972 23180
rect 30656 23128 30708 23180
rect 30840 23171 30892 23180
rect 30840 23137 30849 23171
rect 30849 23137 30883 23171
rect 30883 23137 30892 23171
rect 30840 23128 30892 23137
rect 33784 23196 33836 23248
rect 34336 23239 34388 23248
rect 34336 23205 34345 23239
rect 34345 23205 34379 23239
rect 34379 23205 34388 23239
rect 34336 23196 34388 23205
rect 35256 23196 35308 23248
rect 32496 23171 32548 23180
rect 32496 23137 32505 23171
rect 32505 23137 32539 23171
rect 32539 23137 32548 23171
rect 32496 23128 32548 23137
rect 33048 23171 33100 23180
rect 33048 23137 33057 23171
rect 33057 23137 33091 23171
rect 33091 23137 33100 23171
rect 33048 23128 33100 23137
rect 34244 23171 34296 23180
rect 34244 23137 34253 23171
rect 34253 23137 34287 23171
rect 34287 23137 34296 23171
rect 34244 23128 34296 23137
rect 34612 23128 34664 23180
rect 35532 23171 35584 23180
rect 27620 23060 27672 23112
rect 29092 23103 29144 23112
rect 27712 22992 27764 23044
rect 29092 23069 29101 23103
rect 29101 23069 29135 23103
rect 29135 23069 29144 23103
rect 29092 23060 29144 23069
rect 29828 23060 29880 23112
rect 32956 23103 33008 23112
rect 32956 23069 32965 23103
rect 32965 23069 32999 23103
rect 32999 23069 33008 23103
rect 32956 23060 33008 23069
rect 35532 23137 35541 23171
rect 35541 23137 35575 23171
rect 35575 23137 35584 23171
rect 35532 23128 35584 23137
rect 36452 23171 36504 23180
rect 36452 23137 36461 23171
rect 36461 23137 36495 23171
rect 36495 23137 36504 23171
rect 36452 23128 36504 23137
rect 38660 23196 38712 23248
rect 38200 23171 38252 23180
rect 35440 23060 35492 23112
rect 36820 23103 36872 23112
rect 36820 23069 36829 23103
rect 36829 23069 36863 23103
rect 36863 23069 36872 23103
rect 36820 23060 36872 23069
rect 29276 22992 29328 23044
rect 29552 22992 29604 23044
rect 31024 23035 31076 23044
rect 29460 22924 29512 22976
rect 30012 22924 30064 22976
rect 31024 23001 31033 23035
rect 31033 23001 31067 23035
rect 31067 23001 31076 23035
rect 31024 22992 31076 23001
rect 31208 22992 31260 23044
rect 38200 23137 38209 23171
rect 38209 23137 38243 23171
rect 38243 23137 38252 23171
rect 38200 23128 38252 23137
rect 38384 23128 38436 23180
rect 38844 23060 38896 23112
rect 31484 22924 31536 22976
rect 34612 22924 34664 22976
rect 35348 22924 35400 22976
rect 35716 22924 35768 22976
rect 4246 22822 4298 22874
rect 4310 22822 4362 22874
rect 4374 22822 4426 22874
rect 4438 22822 4490 22874
rect 34966 22822 35018 22874
rect 35030 22822 35082 22874
rect 35094 22822 35146 22874
rect 35158 22822 35210 22874
rect 1768 22763 1820 22772
rect 1768 22729 1777 22763
rect 1777 22729 1811 22763
rect 1811 22729 1820 22763
rect 1768 22720 1820 22729
rect 7288 22720 7340 22772
rect 11888 22720 11940 22772
rect 12716 22720 12768 22772
rect 21180 22720 21232 22772
rect 26516 22763 26568 22772
rect 2044 22652 2096 22704
rect 3332 22652 3384 22704
rect 6000 22652 6052 22704
rect 6092 22652 6144 22704
rect 7012 22652 7064 22704
rect 2780 22584 2832 22636
rect 4620 22584 4672 22636
rect 6828 22627 6880 22636
rect 6828 22593 6837 22627
rect 6837 22593 6871 22627
rect 6871 22593 6880 22627
rect 6828 22584 6880 22593
rect 2964 22516 3016 22568
rect 3332 22559 3384 22568
rect 3332 22525 3341 22559
rect 3341 22525 3375 22559
rect 3375 22525 3384 22559
rect 3332 22516 3384 22525
rect 3516 22559 3568 22568
rect 3516 22525 3525 22559
rect 3525 22525 3559 22559
rect 3559 22525 3568 22559
rect 3516 22516 3568 22525
rect 3792 22559 3844 22568
rect 3792 22525 3801 22559
rect 3801 22525 3835 22559
rect 3835 22525 3844 22559
rect 3792 22516 3844 22525
rect 4712 22559 4764 22568
rect 4712 22525 4721 22559
rect 4721 22525 4755 22559
rect 4755 22525 4764 22559
rect 4712 22516 4764 22525
rect 5632 22516 5684 22568
rect 2780 22448 2832 22500
rect 3700 22448 3752 22500
rect 6184 22516 6236 22568
rect 7104 22491 7156 22500
rect 7104 22457 7113 22491
rect 7113 22457 7147 22491
rect 7147 22457 7156 22491
rect 7104 22448 7156 22457
rect 5356 22380 5408 22432
rect 6184 22380 6236 22432
rect 12900 22652 12952 22704
rect 7840 22584 7892 22636
rect 8484 22627 8536 22636
rect 8484 22593 8493 22627
rect 8493 22593 8527 22627
rect 8527 22593 8536 22627
rect 8484 22584 8536 22593
rect 10140 22584 10192 22636
rect 13912 22584 13964 22636
rect 14464 22584 14516 22636
rect 15292 22584 15344 22636
rect 15752 22627 15804 22636
rect 15752 22593 15761 22627
rect 15761 22593 15795 22627
rect 15795 22593 15804 22627
rect 15752 22584 15804 22593
rect 17224 22627 17276 22636
rect 17224 22593 17233 22627
rect 17233 22593 17267 22627
rect 17267 22593 17276 22627
rect 17224 22584 17276 22593
rect 18328 22584 18380 22636
rect 11796 22516 11848 22568
rect 12440 22559 12492 22568
rect 12440 22525 12449 22559
rect 12449 22525 12483 22559
rect 12483 22525 12492 22559
rect 13176 22559 13228 22568
rect 12440 22516 12492 22525
rect 13176 22525 13185 22559
rect 13185 22525 13219 22559
rect 13219 22525 13228 22559
rect 13176 22516 13228 22525
rect 13728 22559 13780 22568
rect 13728 22525 13737 22559
rect 13737 22525 13771 22559
rect 13771 22525 13780 22559
rect 13728 22516 13780 22525
rect 11612 22448 11664 22500
rect 14372 22448 14424 22500
rect 15108 22516 15160 22568
rect 16764 22559 16816 22568
rect 16764 22525 16773 22559
rect 16773 22525 16807 22559
rect 16807 22525 16816 22559
rect 16764 22516 16816 22525
rect 16856 22516 16908 22568
rect 18420 22559 18472 22568
rect 18420 22525 18429 22559
rect 18429 22525 18463 22559
rect 18463 22525 18472 22559
rect 18420 22516 18472 22525
rect 17960 22448 18012 22500
rect 18696 22448 18748 22500
rect 21088 22516 21140 22568
rect 21824 22652 21876 22704
rect 26516 22729 26525 22763
rect 26525 22729 26559 22763
rect 26559 22729 26568 22763
rect 26516 22720 26568 22729
rect 28724 22720 28776 22772
rect 29828 22720 29880 22772
rect 30564 22720 30616 22772
rect 36268 22720 36320 22772
rect 37188 22720 37240 22772
rect 38200 22720 38252 22772
rect 21364 22627 21416 22636
rect 21364 22593 21373 22627
rect 21373 22593 21407 22627
rect 21407 22593 21416 22627
rect 21364 22584 21416 22593
rect 21456 22516 21508 22568
rect 22836 22516 22888 22568
rect 23940 22584 23992 22636
rect 24032 22584 24084 22636
rect 24216 22627 24268 22636
rect 24216 22593 24225 22627
rect 24225 22593 24259 22627
rect 24259 22593 24268 22627
rect 24216 22584 24268 22593
rect 28356 22627 28408 22636
rect 28356 22593 28365 22627
rect 28365 22593 28399 22627
rect 28399 22593 28408 22627
rect 28356 22584 28408 22593
rect 31024 22652 31076 22704
rect 34520 22652 34572 22704
rect 23020 22516 23072 22568
rect 23756 22559 23808 22568
rect 23756 22525 23765 22559
rect 23765 22525 23799 22559
rect 23799 22525 23808 22559
rect 23756 22516 23808 22525
rect 23848 22516 23900 22568
rect 24676 22516 24728 22568
rect 25136 22559 25188 22568
rect 25136 22525 25145 22559
rect 25145 22525 25179 22559
rect 25179 22525 25188 22559
rect 25136 22516 25188 22525
rect 25412 22559 25464 22568
rect 25412 22525 25421 22559
rect 25421 22525 25455 22559
rect 25455 22525 25464 22559
rect 25412 22516 25464 22525
rect 25688 22516 25740 22568
rect 27896 22559 27948 22568
rect 23572 22448 23624 22500
rect 27896 22525 27905 22559
rect 27905 22525 27939 22559
rect 27939 22525 27948 22559
rect 27896 22516 27948 22525
rect 28632 22516 28684 22568
rect 29460 22559 29512 22568
rect 29460 22525 29469 22559
rect 29469 22525 29503 22559
rect 29503 22525 29512 22559
rect 29460 22516 29512 22525
rect 8208 22380 8260 22432
rect 9772 22380 9824 22432
rect 11152 22423 11204 22432
rect 11152 22389 11161 22423
rect 11161 22389 11195 22423
rect 11195 22389 11204 22423
rect 11152 22380 11204 22389
rect 11244 22423 11296 22432
rect 11244 22389 11253 22423
rect 11253 22389 11287 22423
rect 11287 22389 11296 22423
rect 11244 22380 11296 22389
rect 19156 22380 19208 22432
rect 23664 22380 23716 22432
rect 27988 22380 28040 22432
rect 29000 22448 29052 22500
rect 33692 22584 33744 22636
rect 31208 22559 31260 22568
rect 29828 22448 29880 22500
rect 31208 22525 31217 22559
rect 31217 22525 31251 22559
rect 31251 22525 31260 22559
rect 31208 22516 31260 22525
rect 31576 22516 31628 22568
rect 33324 22559 33376 22568
rect 33324 22525 33333 22559
rect 33333 22525 33367 22559
rect 33367 22525 33376 22559
rect 36360 22584 36412 22636
rect 37464 22627 37516 22636
rect 37464 22593 37473 22627
rect 37473 22593 37507 22627
rect 37507 22593 37516 22627
rect 37464 22584 37516 22593
rect 38752 22584 38804 22636
rect 33324 22516 33376 22525
rect 34612 22516 34664 22568
rect 35164 22559 35216 22568
rect 35164 22525 35173 22559
rect 35173 22525 35207 22559
rect 35207 22525 35216 22559
rect 35164 22516 35216 22525
rect 33508 22448 33560 22500
rect 29552 22380 29604 22432
rect 30012 22380 30064 22432
rect 30932 22380 30984 22432
rect 36452 22380 36504 22432
rect 38844 22380 38896 22432
rect 19606 22278 19658 22330
rect 19670 22278 19722 22330
rect 19734 22278 19786 22330
rect 19798 22278 19850 22330
rect 4896 22176 4948 22228
rect 7196 22176 7248 22228
rect 7380 22176 7432 22228
rect 1492 22083 1544 22092
rect 1492 22049 1501 22083
rect 1501 22049 1535 22083
rect 1535 22049 1544 22083
rect 1492 22040 1544 22049
rect 2964 22083 3016 22092
rect 2964 22049 2973 22083
rect 2973 22049 3007 22083
rect 3007 22049 3016 22083
rect 2964 22040 3016 22049
rect 3700 22040 3752 22092
rect 4068 22083 4120 22092
rect 4068 22049 4077 22083
rect 4077 22049 4111 22083
rect 4111 22049 4120 22083
rect 4068 22040 4120 22049
rect 4620 22083 4672 22092
rect 4620 22049 4629 22083
rect 4629 22049 4663 22083
rect 4663 22049 4672 22083
rect 4620 22040 4672 22049
rect 5356 22083 5408 22092
rect 5356 22049 5365 22083
rect 5365 22049 5399 22083
rect 5399 22049 5408 22083
rect 5356 22040 5408 22049
rect 5816 22083 5868 22092
rect 5816 22049 5825 22083
rect 5825 22049 5859 22083
rect 5859 22049 5868 22083
rect 5816 22040 5868 22049
rect 6276 22040 6328 22092
rect 6920 22083 6972 22092
rect 6920 22049 6929 22083
rect 6929 22049 6963 22083
rect 6963 22049 6972 22083
rect 6920 22040 6972 22049
rect 7104 22040 7156 22092
rect 7748 22083 7800 22092
rect 4896 21972 4948 22024
rect 7748 22049 7757 22083
rect 7757 22049 7791 22083
rect 7791 22049 7800 22083
rect 7748 22040 7800 22049
rect 8116 22040 8168 22092
rect 8576 22176 8628 22228
rect 11244 22176 11296 22228
rect 12348 22176 12400 22228
rect 13544 22176 13596 22228
rect 15752 22176 15804 22228
rect 16856 22219 16908 22228
rect 8760 22151 8812 22160
rect 8760 22117 8769 22151
rect 8769 22117 8803 22151
rect 8803 22117 8812 22151
rect 8760 22108 8812 22117
rect 9680 22108 9732 22160
rect 10968 22108 11020 22160
rect 8300 21972 8352 22024
rect 8484 21972 8536 22024
rect 2412 21904 2464 21956
rect 3792 21904 3844 21956
rect 10876 22040 10928 22092
rect 11704 22040 11756 22092
rect 12348 22083 12400 22092
rect 12348 22049 12357 22083
rect 12357 22049 12391 22083
rect 12391 22049 12400 22083
rect 12348 22040 12400 22049
rect 13176 22083 13228 22092
rect 13176 22049 13185 22083
rect 13185 22049 13219 22083
rect 13219 22049 13228 22083
rect 13176 22040 13228 22049
rect 14004 22040 14056 22092
rect 14832 22083 14884 22092
rect 14832 22049 14841 22083
rect 14841 22049 14875 22083
rect 14875 22049 14884 22083
rect 14832 22040 14884 22049
rect 9956 21972 10008 22024
rect 10232 22015 10284 22024
rect 10232 21981 10241 22015
rect 10241 21981 10275 22015
rect 10275 21981 10284 22015
rect 10232 21972 10284 21981
rect 11060 21972 11112 22024
rect 13912 22015 13964 22024
rect 10324 21904 10376 21956
rect 13912 21981 13921 22015
rect 13921 21981 13955 22015
rect 13955 21981 13964 22015
rect 13912 21972 13964 21981
rect 16396 22108 16448 22160
rect 16856 22185 16865 22219
rect 16865 22185 16899 22219
rect 16899 22185 16908 22219
rect 16856 22176 16908 22185
rect 23756 22176 23808 22228
rect 27712 22219 27764 22228
rect 27712 22185 27721 22219
rect 27721 22185 27755 22219
rect 27755 22185 27764 22219
rect 27712 22176 27764 22185
rect 27896 22176 27948 22228
rect 21088 22108 21140 22160
rect 1676 21836 1728 21888
rect 2872 21879 2924 21888
rect 2872 21845 2881 21879
rect 2881 21845 2915 21879
rect 2915 21845 2924 21879
rect 2872 21836 2924 21845
rect 3056 21836 3108 21888
rect 4988 21836 5040 21888
rect 13820 21836 13872 21888
rect 15752 22040 15804 22092
rect 16212 22040 16264 22092
rect 17960 22040 18012 22092
rect 19156 22040 19208 22092
rect 19340 22040 19392 22092
rect 19432 22083 19484 22092
rect 19432 22049 19441 22083
rect 19441 22049 19475 22083
rect 19475 22049 19484 22083
rect 19432 22040 19484 22049
rect 20260 22040 20312 22092
rect 16396 21972 16448 22024
rect 17868 21972 17920 22024
rect 20996 22040 21048 22092
rect 21548 22040 21600 22092
rect 22008 22108 22060 22160
rect 21824 22040 21876 22092
rect 22744 22083 22796 22092
rect 22744 22049 22753 22083
rect 22753 22049 22787 22083
rect 22787 22049 22796 22083
rect 22744 22040 22796 22049
rect 22836 22040 22888 22092
rect 23388 22083 23440 22092
rect 23388 22049 23397 22083
rect 23397 22049 23431 22083
rect 23431 22049 23440 22083
rect 23388 22040 23440 22049
rect 25136 22108 25188 22160
rect 25504 22108 25556 22160
rect 25228 22040 25280 22092
rect 25596 22040 25648 22092
rect 26516 22083 26568 22092
rect 26516 22049 26525 22083
rect 26525 22049 26559 22083
rect 26559 22049 26568 22083
rect 26516 22040 26568 22049
rect 27620 22083 27672 22092
rect 27620 22049 27629 22083
rect 27629 22049 27663 22083
rect 27663 22049 27672 22083
rect 27620 22040 27672 22049
rect 27804 22040 27856 22092
rect 29092 22108 29144 22160
rect 29644 22083 29696 22092
rect 25964 22015 26016 22024
rect 22652 21904 22704 21956
rect 25964 21981 25973 22015
rect 25973 21981 26007 22015
rect 26007 21981 26016 22015
rect 25964 21972 26016 21981
rect 29644 22049 29653 22083
rect 29653 22049 29687 22083
rect 29687 22049 29696 22083
rect 29644 22040 29696 22049
rect 28724 21972 28776 22024
rect 29092 21972 29144 22024
rect 30196 22176 30248 22228
rect 35900 22176 35952 22228
rect 33232 22108 33284 22160
rect 33692 22108 33744 22160
rect 30012 22040 30064 22092
rect 35072 22040 35124 22092
rect 35256 22083 35308 22092
rect 35256 22049 35265 22083
rect 35265 22049 35299 22083
rect 35299 22049 35308 22083
rect 35256 22040 35308 22049
rect 35440 22083 35492 22092
rect 35440 22049 35449 22083
rect 35449 22049 35483 22083
rect 35483 22049 35492 22083
rect 35440 22040 35492 22049
rect 37004 22108 37056 22160
rect 32128 22015 32180 22024
rect 32128 21981 32137 22015
rect 32137 21981 32171 22015
rect 32171 21981 32180 22015
rect 32128 21972 32180 21981
rect 32404 22015 32456 22024
rect 32404 21981 32413 22015
rect 32413 21981 32447 22015
rect 32447 21981 32456 22015
rect 32404 21972 32456 21981
rect 34612 21972 34664 22024
rect 35164 22015 35216 22024
rect 35164 21981 35173 22015
rect 35173 21981 35207 22015
rect 35207 21981 35216 22015
rect 35164 21972 35216 21981
rect 26240 21904 26292 21956
rect 33508 21904 33560 21956
rect 34888 21904 34940 21956
rect 15384 21879 15436 21888
rect 15384 21845 15393 21879
rect 15393 21845 15427 21879
rect 15427 21845 15436 21879
rect 15384 21836 15436 21845
rect 19432 21836 19484 21888
rect 20536 21836 20588 21888
rect 21364 21836 21416 21888
rect 21548 21836 21600 21888
rect 22928 21836 22980 21888
rect 24860 21836 24912 21888
rect 29092 21879 29144 21888
rect 29092 21845 29101 21879
rect 29101 21845 29135 21879
rect 29135 21845 29144 21879
rect 29092 21836 29144 21845
rect 33692 21879 33744 21888
rect 33692 21845 33701 21879
rect 33701 21845 33735 21879
rect 33735 21845 33744 21879
rect 33692 21836 33744 21845
rect 34796 21836 34848 21888
rect 37832 22083 37884 22092
rect 37832 22049 37841 22083
rect 37841 22049 37875 22083
rect 37875 22049 37884 22083
rect 37832 22040 37884 22049
rect 36820 21904 36872 21956
rect 36452 21836 36504 21888
rect 37556 21904 37608 21956
rect 4246 21734 4298 21786
rect 4310 21734 4362 21786
rect 4374 21734 4426 21786
rect 4438 21734 4490 21786
rect 34966 21734 35018 21786
rect 35030 21734 35082 21786
rect 35094 21734 35146 21786
rect 35158 21734 35210 21786
rect 4068 21632 4120 21684
rect 6828 21632 6880 21684
rect 9864 21632 9916 21684
rect 11060 21632 11112 21684
rect 11520 21675 11572 21684
rect 11520 21641 11529 21675
rect 11529 21641 11563 21675
rect 11563 21641 11572 21675
rect 11520 21632 11572 21641
rect 15476 21632 15528 21684
rect 19340 21632 19392 21684
rect 20076 21632 20128 21684
rect 1492 21564 1544 21616
rect 8392 21564 8444 21616
rect 9680 21564 9732 21616
rect 14280 21607 14332 21616
rect 2872 21496 2924 21548
rect 2596 21471 2648 21480
rect 2596 21437 2605 21471
rect 2605 21437 2639 21471
rect 2639 21437 2648 21471
rect 2596 21428 2648 21437
rect 2964 21471 3016 21480
rect 2964 21437 2973 21471
rect 2973 21437 3007 21471
rect 3007 21437 3016 21471
rect 2964 21428 3016 21437
rect 3240 21428 3292 21480
rect 4988 21471 5040 21480
rect 4988 21437 4997 21471
rect 4997 21437 5031 21471
rect 5031 21437 5040 21471
rect 4988 21428 5040 21437
rect 8944 21496 8996 21548
rect 10232 21496 10284 21548
rect 5448 21471 5500 21480
rect 5448 21437 5457 21471
rect 5457 21437 5491 21471
rect 5491 21437 5500 21471
rect 5448 21428 5500 21437
rect 7196 21428 7248 21480
rect 8024 21428 8076 21480
rect 8392 21428 8444 21480
rect 9864 21471 9916 21480
rect 3792 21360 3844 21412
rect 4804 21360 4856 21412
rect 9220 21360 9272 21412
rect 9864 21437 9873 21471
rect 9873 21437 9907 21471
rect 9907 21437 9916 21471
rect 9864 21428 9916 21437
rect 10324 21471 10376 21480
rect 10324 21437 10333 21471
rect 10333 21437 10367 21471
rect 10367 21437 10376 21471
rect 10324 21428 10376 21437
rect 14280 21573 14289 21607
rect 14289 21573 14323 21607
rect 14323 21573 14332 21607
rect 14280 21564 14332 21573
rect 12532 21496 12584 21548
rect 13176 21539 13228 21548
rect 11244 21471 11296 21480
rect 11244 21437 11253 21471
rect 11253 21437 11287 21471
rect 11287 21437 11296 21471
rect 11244 21428 11296 21437
rect 12624 21471 12676 21480
rect 10876 21360 10928 21412
rect 10968 21360 11020 21412
rect 12624 21437 12633 21471
rect 12633 21437 12667 21471
rect 12667 21437 12676 21471
rect 12624 21428 12676 21437
rect 13176 21505 13185 21539
rect 13185 21505 13219 21539
rect 13219 21505 13228 21539
rect 13176 21496 13228 21505
rect 16580 21607 16632 21616
rect 16580 21573 16589 21607
rect 16589 21573 16623 21607
rect 16623 21573 16632 21607
rect 16580 21564 16632 21573
rect 13820 21471 13872 21480
rect 13820 21437 13829 21471
rect 13829 21437 13863 21471
rect 13863 21437 13872 21471
rect 13820 21428 13872 21437
rect 17592 21496 17644 21548
rect 13084 21360 13136 21412
rect 15568 21428 15620 21480
rect 16580 21428 16632 21480
rect 16764 21428 16816 21480
rect 20720 21564 20772 21616
rect 19156 21496 19208 21548
rect 19248 21496 19300 21548
rect 18052 21471 18104 21480
rect 18052 21437 18061 21471
rect 18061 21437 18095 21471
rect 18095 21437 18104 21471
rect 18052 21428 18104 21437
rect 19432 21428 19484 21480
rect 15844 21360 15896 21412
rect 19248 21403 19300 21412
rect 19248 21369 19257 21403
rect 19257 21369 19291 21403
rect 19291 21369 19300 21403
rect 19248 21360 19300 21369
rect 19892 21360 19944 21412
rect 20168 21428 20220 21480
rect 21732 21564 21784 21616
rect 22008 21564 22060 21616
rect 23388 21632 23440 21684
rect 25228 21632 25280 21684
rect 29000 21632 29052 21684
rect 29092 21632 29144 21684
rect 33784 21632 33836 21684
rect 34796 21632 34848 21684
rect 38844 21675 38896 21684
rect 38844 21641 38853 21675
rect 38853 21641 38887 21675
rect 38887 21641 38896 21675
rect 38844 21632 38896 21641
rect 23572 21564 23624 21616
rect 25412 21564 25464 21616
rect 28632 21564 28684 21616
rect 21272 21496 21324 21548
rect 21916 21539 21968 21548
rect 21456 21471 21508 21480
rect 21456 21437 21465 21471
rect 21465 21437 21499 21471
rect 21499 21437 21508 21471
rect 21456 21428 21508 21437
rect 21548 21428 21600 21480
rect 21916 21505 21925 21539
rect 21925 21505 21959 21539
rect 21959 21505 21968 21539
rect 21916 21496 21968 21505
rect 23480 21496 23532 21548
rect 24860 21496 24912 21548
rect 25964 21496 26016 21548
rect 27712 21539 27764 21548
rect 27712 21505 27721 21539
rect 27721 21505 27755 21539
rect 27755 21505 27764 21539
rect 27712 21496 27764 21505
rect 23388 21428 23440 21480
rect 23940 21471 23992 21480
rect 23940 21437 23949 21471
rect 23949 21437 23983 21471
rect 23983 21437 23992 21471
rect 23940 21428 23992 21437
rect 26516 21471 26568 21480
rect 23204 21360 23256 21412
rect 12256 21292 12308 21344
rect 17132 21292 17184 21344
rect 19340 21292 19392 21344
rect 19432 21292 19484 21344
rect 22928 21292 22980 21344
rect 24676 21292 24728 21344
rect 26516 21437 26525 21471
rect 26525 21437 26559 21471
rect 26559 21437 26568 21471
rect 26516 21428 26568 21437
rect 27988 21471 28040 21480
rect 27988 21437 27997 21471
rect 27997 21437 28031 21471
rect 28031 21437 28040 21471
rect 27988 21428 28040 21437
rect 28632 21428 28684 21480
rect 29184 21428 29236 21480
rect 30288 21539 30340 21548
rect 30288 21505 30297 21539
rect 30297 21505 30331 21539
rect 30331 21505 30340 21539
rect 30288 21496 30340 21505
rect 36636 21496 36688 21548
rect 37556 21539 37608 21548
rect 37556 21505 37565 21539
rect 37565 21505 37599 21539
rect 37599 21505 37608 21539
rect 37556 21496 37608 21505
rect 30104 21471 30156 21480
rect 30104 21437 30113 21471
rect 30113 21437 30147 21471
rect 30147 21437 30156 21471
rect 30104 21428 30156 21437
rect 30564 21471 30616 21480
rect 30564 21437 30573 21471
rect 30573 21437 30607 21471
rect 30607 21437 30616 21471
rect 30564 21428 30616 21437
rect 31116 21428 31168 21480
rect 31852 21471 31904 21480
rect 31852 21437 31861 21471
rect 31861 21437 31895 21471
rect 31895 21437 31904 21471
rect 31852 21428 31904 21437
rect 32036 21471 32088 21480
rect 32036 21437 32045 21471
rect 32045 21437 32079 21471
rect 32079 21437 32088 21471
rect 32036 21428 32088 21437
rect 32312 21428 32364 21480
rect 33232 21471 33284 21480
rect 33232 21437 33241 21471
rect 33241 21437 33275 21471
rect 33275 21437 33284 21471
rect 33232 21428 33284 21437
rect 35716 21471 35768 21480
rect 29828 21360 29880 21412
rect 30012 21360 30064 21412
rect 35716 21437 35725 21471
rect 35725 21437 35759 21471
rect 35759 21437 35768 21471
rect 35716 21428 35768 21437
rect 35808 21428 35860 21480
rect 36084 21428 36136 21480
rect 36360 21471 36412 21480
rect 36360 21437 36369 21471
rect 36369 21437 36403 21471
rect 36403 21437 36412 21471
rect 36360 21428 36412 21437
rect 37280 21471 37332 21480
rect 37280 21437 37289 21471
rect 37289 21437 37323 21471
rect 37323 21437 37332 21471
rect 37280 21428 37332 21437
rect 35256 21360 35308 21412
rect 29276 21292 29328 21344
rect 31300 21335 31352 21344
rect 31300 21301 31309 21335
rect 31309 21301 31343 21335
rect 31343 21301 31352 21335
rect 31300 21292 31352 21301
rect 32404 21292 32456 21344
rect 34336 21292 34388 21344
rect 19606 21190 19658 21242
rect 19670 21190 19722 21242
rect 19734 21190 19786 21242
rect 19798 21190 19850 21242
rect 11152 21088 11204 21140
rect 2964 21020 3016 21072
rect 1400 20995 1452 21004
rect 1400 20961 1409 20995
rect 1409 20961 1443 20995
rect 1443 20961 1452 20995
rect 1400 20952 1452 20961
rect 1676 20995 1728 21004
rect 1676 20961 1685 20995
rect 1685 20961 1719 20995
rect 1719 20961 1728 20995
rect 1676 20952 1728 20961
rect 2596 20952 2648 21004
rect 4712 21020 4764 21072
rect 5448 21020 5500 21072
rect 4804 20995 4856 21004
rect 4804 20961 4813 20995
rect 4813 20961 4847 20995
rect 4847 20961 4856 20995
rect 4804 20952 4856 20961
rect 6276 20995 6328 21004
rect 6276 20961 6285 20995
rect 6285 20961 6319 20995
rect 6319 20961 6328 20995
rect 6276 20952 6328 20961
rect 6920 20952 6972 21004
rect 8024 21020 8076 21072
rect 7840 20995 7892 21004
rect 7840 20961 7849 20995
rect 7849 20961 7883 20995
rect 7883 20961 7892 20995
rect 7840 20952 7892 20961
rect 8392 20995 8444 21004
rect 8392 20961 8401 20995
rect 8401 20961 8435 20995
rect 8435 20961 8444 20995
rect 8392 20952 8444 20961
rect 5816 20927 5868 20936
rect 5816 20893 5825 20927
rect 5825 20893 5859 20927
rect 5859 20893 5868 20927
rect 5816 20884 5868 20893
rect 9772 20952 9824 21004
rect 9956 20995 10008 21004
rect 9956 20961 9965 20995
rect 9965 20961 9999 20995
rect 9999 20961 10008 20995
rect 9956 20952 10008 20961
rect 12532 21088 12584 21140
rect 16764 21131 16816 21140
rect 16764 21097 16773 21131
rect 16773 21097 16807 21131
rect 16807 21097 16816 21131
rect 16764 21088 16816 21097
rect 18052 21088 18104 21140
rect 15752 21020 15804 21072
rect 12532 20995 12584 21004
rect 12532 20961 12541 20995
rect 12541 20961 12575 20995
rect 12575 20961 12584 20995
rect 13084 20995 13136 21004
rect 12532 20952 12584 20961
rect 13084 20961 13093 20995
rect 13093 20961 13127 20995
rect 13127 20961 13136 20995
rect 13084 20952 13136 20961
rect 14648 20952 14700 21004
rect 16948 21020 17000 21072
rect 19340 21020 19392 21072
rect 16764 20952 16816 21004
rect 5356 20816 5408 20868
rect 15108 20884 15160 20936
rect 17868 20952 17920 21004
rect 19892 21020 19944 21072
rect 21456 21088 21508 21140
rect 17960 20884 18012 20936
rect 19156 20884 19208 20936
rect 20168 20952 20220 21004
rect 21088 20995 21140 21004
rect 21088 20961 21097 20995
rect 21097 20961 21131 20995
rect 21131 20961 21140 20995
rect 21088 20952 21140 20961
rect 20260 20884 20312 20936
rect 21548 20884 21600 20936
rect 10876 20816 10928 20868
rect 22100 21088 22152 21140
rect 22928 21088 22980 21140
rect 23112 21131 23164 21140
rect 23112 21097 23121 21131
rect 23121 21097 23155 21131
rect 23155 21097 23164 21131
rect 23112 21088 23164 21097
rect 23204 21088 23256 21140
rect 21824 20995 21876 21004
rect 21824 20961 21833 20995
rect 21833 20961 21867 20995
rect 21867 20961 21876 20995
rect 21824 20952 21876 20961
rect 22284 20952 22336 21004
rect 22836 20952 22888 21004
rect 23572 21020 23624 21072
rect 24124 21020 24176 21072
rect 24952 21063 25004 21072
rect 24952 21029 24961 21063
rect 24961 21029 24995 21063
rect 24995 21029 25004 21063
rect 24952 21020 25004 21029
rect 25136 21088 25188 21140
rect 28632 21131 28684 21140
rect 28632 21097 28641 21131
rect 28641 21097 28675 21131
rect 28675 21097 28684 21131
rect 28632 21088 28684 21097
rect 35716 21088 35768 21140
rect 36452 21088 36504 21140
rect 29092 21020 29144 21072
rect 22560 20927 22612 20936
rect 22560 20893 22569 20927
rect 22569 20893 22603 20927
rect 22603 20893 22612 20927
rect 22560 20884 22612 20893
rect 7472 20748 7524 20800
rect 8208 20748 8260 20800
rect 8944 20791 8996 20800
rect 8944 20757 8953 20791
rect 8953 20757 8987 20791
rect 8987 20757 8996 20791
rect 8944 20748 8996 20757
rect 13084 20748 13136 20800
rect 16212 20748 16264 20800
rect 22008 20816 22060 20868
rect 24400 20995 24452 21004
rect 24400 20961 24409 20995
rect 24409 20961 24443 20995
rect 24443 20961 24452 20995
rect 24400 20952 24452 20961
rect 24676 20952 24728 21004
rect 27620 20995 27672 21004
rect 24216 20927 24268 20936
rect 24216 20893 24225 20927
rect 24225 20893 24259 20927
rect 24259 20893 24268 20927
rect 24216 20884 24268 20893
rect 27620 20961 27629 20995
rect 27629 20961 27663 20995
rect 27663 20961 27672 20995
rect 27620 20952 27672 20961
rect 27712 20952 27764 21004
rect 28356 20995 28408 21004
rect 28356 20961 28365 20995
rect 28365 20961 28399 20995
rect 28399 20961 28408 20995
rect 28356 20952 28408 20961
rect 29276 20995 29328 21004
rect 29276 20961 29285 20995
rect 29285 20961 29319 20995
rect 29319 20961 29328 20995
rect 29276 20952 29328 20961
rect 29828 20995 29880 21004
rect 29828 20961 29837 20995
rect 29837 20961 29871 20995
rect 29871 20961 29880 20995
rect 29828 20952 29880 20961
rect 30288 20995 30340 21004
rect 30288 20961 30297 20995
rect 30297 20961 30331 20995
rect 30331 20961 30340 20995
rect 30288 20952 30340 20961
rect 32036 21020 32088 21072
rect 32680 20952 32732 21004
rect 33508 21020 33560 21072
rect 33784 21020 33836 21072
rect 32864 20995 32916 21004
rect 32864 20961 32873 20995
rect 32873 20961 32907 20995
rect 32907 20961 32916 20995
rect 33416 20995 33468 21004
rect 32864 20952 32916 20961
rect 33416 20961 33425 20995
rect 33425 20961 33459 20995
rect 33459 20961 33468 20995
rect 33416 20952 33468 20961
rect 34336 20995 34388 21004
rect 34336 20961 34345 20995
rect 34345 20961 34379 20995
rect 34379 20961 34388 20995
rect 34336 20952 34388 20961
rect 34980 20952 35032 21004
rect 33048 20927 33100 20936
rect 19892 20748 19944 20800
rect 20076 20748 20128 20800
rect 21456 20748 21508 20800
rect 22744 20748 22796 20800
rect 22836 20748 22888 20800
rect 33048 20893 33057 20927
rect 33057 20893 33091 20927
rect 33091 20893 33100 20927
rect 33048 20884 33100 20893
rect 34520 20927 34572 20936
rect 34520 20893 34529 20927
rect 34529 20893 34563 20927
rect 34563 20893 34572 20927
rect 34520 20884 34572 20893
rect 35348 20952 35400 21004
rect 38660 21020 38712 21072
rect 37832 20995 37884 21004
rect 37832 20961 37841 20995
rect 37841 20961 37875 20995
rect 37875 20961 37884 20995
rect 37832 20952 37884 20961
rect 38568 20995 38620 21004
rect 38568 20961 38577 20995
rect 38577 20961 38611 20995
rect 38611 20961 38620 20995
rect 38568 20952 38620 20961
rect 35440 20884 35492 20936
rect 35900 20884 35952 20936
rect 38476 20884 38528 20936
rect 27620 20816 27672 20868
rect 31576 20816 31628 20868
rect 37188 20816 37240 20868
rect 37740 20816 37792 20868
rect 38108 20748 38160 20800
rect 4246 20646 4298 20698
rect 4310 20646 4362 20698
rect 4374 20646 4426 20698
rect 4438 20646 4490 20698
rect 34966 20646 35018 20698
rect 35030 20646 35082 20698
rect 35094 20646 35146 20698
rect 35158 20646 35210 20698
rect 2964 20408 3016 20460
rect 2780 20340 2832 20392
rect 3240 20383 3292 20392
rect 3240 20349 3249 20383
rect 3249 20349 3283 20383
rect 3283 20349 3292 20383
rect 3240 20340 3292 20349
rect 6460 20544 6512 20596
rect 4620 20476 4672 20528
rect 5448 20408 5500 20460
rect 5356 20340 5408 20392
rect 6828 20476 6880 20528
rect 5908 20340 5960 20392
rect 6828 20383 6880 20392
rect 6828 20349 6837 20383
rect 6837 20349 6871 20383
rect 6871 20349 6880 20383
rect 6828 20340 6880 20349
rect 8116 20544 8168 20596
rect 16396 20544 16448 20596
rect 20260 20544 20312 20596
rect 8392 20476 8444 20528
rect 8024 20408 8076 20460
rect 9864 20383 9916 20392
rect 9864 20349 9873 20383
rect 9873 20349 9907 20383
rect 9907 20349 9916 20383
rect 9864 20340 9916 20349
rect 11336 20340 11388 20392
rect 12900 20476 12952 20528
rect 15292 20519 15344 20528
rect 15292 20485 15301 20519
rect 15301 20485 15335 20519
rect 15335 20485 15344 20519
rect 15292 20476 15344 20485
rect 13084 20408 13136 20460
rect 14740 20408 14792 20460
rect 14924 20408 14976 20460
rect 15108 20408 15160 20460
rect 11704 20383 11756 20392
rect 11704 20349 11713 20383
rect 11713 20349 11747 20383
rect 11747 20349 11756 20383
rect 11704 20340 11756 20349
rect 12716 20340 12768 20392
rect 12992 20383 13044 20392
rect 12992 20349 13001 20383
rect 13001 20349 13035 20383
rect 13035 20349 13044 20383
rect 12992 20340 13044 20349
rect 13912 20340 13964 20392
rect 15200 20340 15252 20392
rect 16304 20383 16356 20392
rect 16304 20349 16313 20383
rect 16313 20349 16347 20383
rect 16347 20349 16356 20383
rect 16304 20340 16356 20349
rect 16672 20340 16724 20392
rect 18236 20476 18288 20528
rect 21088 20476 21140 20528
rect 22008 20476 22060 20528
rect 17500 20451 17552 20460
rect 17500 20417 17509 20451
rect 17509 20417 17543 20451
rect 17543 20417 17552 20451
rect 17500 20408 17552 20417
rect 17408 20340 17460 20392
rect 17776 20340 17828 20392
rect 21548 20451 21600 20460
rect 21548 20417 21557 20451
rect 21557 20417 21591 20451
rect 21591 20417 21600 20451
rect 25596 20544 25648 20596
rect 26700 20544 26752 20596
rect 31116 20544 31168 20596
rect 28172 20476 28224 20528
rect 21548 20408 21600 20417
rect 21272 20383 21324 20392
rect 21272 20349 21281 20383
rect 21281 20349 21315 20383
rect 21315 20349 21324 20383
rect 21272 20340 21324 20349
rect 21364 20340 21416 20392
rect 8392 20247 8444 20256
rect 8392 20213 8401 20247
rect 8401 20213 8435 20247
rect 8435 20213 8444 20247
rect 8392 20204 8444 20213
rect 13544 20272 13596 20324
rect 18420 20315 18472 20324
rect 18420 20281 18429 20315
rect 18429 20281 18463 20315
rect 18463 20281 18472 20315
rect 18420 20272 18472 20281
rect 22560 20408 22612 20460
rect 22836 20383 22888 20392
rect 22836 20349 22845 20383
rect 22845 20349 22879 20383
rect 22879 20349 22888 20383
rect 22836 20340 22888 20349
rect 22928 20340 22980 20392
rect 23480 20340 23532 20392
rect 24400 20340 24452 20392
rect 25964 20383 26016 20392
rect 25964 20349 25973 20383
rect 25973 20349 26007 20383
rect 26007 20349 26016 20383
rect 25964 20340 26016 20349
rect 27620 20408 27672 20460
rect 27528 20340 27580 20392
rect 28448 20383 28500 20392
rect 28448 20349 28457 20383
rect 28457 20349 28491 20383
rect 28491 20349 28500 20383
rect 28448 20340 28500 20349
rect 28540 20383 28592 20392
rect 28540 20349 28549 20383
rect 28549 20349 28583 20383
rect 28583 20349 28592 20383
rect 28540 20340 28592 20349
rect 30288 20340 30340 20392
rect 31300 20408 31352 20460
rect 33048 20544 33100 20596
rect 35348 20476 35400 20528
rect 34520 20408 34572 20460
rect 35900 20408 35952 20460
rect 25504 20315 25556 20324
rect 25504 20281 25513 20315
rect 25513 20281 25547 20315
rect 25547 20281 25556 20315
rect 25504 20272 25556 20281
rect 34060 20340 34112 20392
rect 35256 20383 35308 20392
rect 35256 20349 35265 20383
rect 35265 20349 35299 20383
rect 35299 20349 35308 20383
rect 35256 20340 35308 20349
rect 36084 20340 36136 20392
rect 36268 20340 36320 20392
rect 37740 20451 37792 20460
rect 37740 20417 37749 20451
rect 37749 20417 37783 20451
rect 37783 20417 37792 20451
rect 37740 20408 37792 20417
rect 34520 20272 34572 20324
rect 37280 20340 37332 20392
rect 13820 20204 13872 20256
rect 16120 20247 16172 20256
rect 16120 20213 16129 20247
rect 16129 20213 16163 20247
rect 16163 20213 16172 20247
rect 16120 20204 16172 20213
rect 16212 20204 16264 20256
rect 19432 20204 19484 20256
rect 22192 20204 22244 20256
rect 23848 20247 23900 20256
rect 23848 20213 23857 20247
rect 23857 20213 23891 20247
rect 23891 20213 23900 20247
rect 23848 20204 23900 20213
rect 24308 20204 24360 20256
rect 25136 20204 25188 20256
rect 26332 20204 26384 20256
rect 29736 20204 29788 20256
rect 32496 20204 32548 20256
rect 32680 20247 32732 20256
rect 32680 20213 32689 20247
rect 32689 20213 32723 20247
rect 32723 20213 32732 20247
rect 32680 20204 32732 20213
rect 33048 20204 33100 20256
rect 33784 20204 33836 20256
rect 38108 20204 38160 20256
rect 19606 20102 19658 20154
rect 19670 20102 19722 20154
rect 19734 20102 19786 20154
rect 19798 20102 19850 20154
rect 3240 19932 3292 19984
rect 1400 19907 1452 19916
rect 1400 19873 1409 19907
rect 1409 19873 1443 19907
rect 1443 19873 1452 19907
rect 1400 19864 1452 19873
rect 3884 19864 3936 19916
rect 11336 20000 11388 20052
rect 11704 20000 11756 20052
rect 12808 20043 12860 20052
rect 12808 20009 12817 20043
rect 12817 20009 12851 20043
rect 12851 20009 12860 20043
rect 12808 20000 12860 20009
rect 12992 20000 13044 20052
rect 13360 20000 13412 20052
rect 16212 20000 16264 20052
rect 17408 20043 17460 20052
rect 17408 20009 17417 20043
rect 17417 20009 17451 20043
rect 17451 20009 17460 20043
rect 17408 20000 17460 20009
rect 17500 20000 17552 20052
rect 19156 20000 19208 20052
rect 5816 19932 5868 19984
rect 5540 19907 5592 19916
rect 5540 19873 5549 19907
rect 5549 19873 5583 19907
rect 5583 19873 5592 19907
rect 5540 19864 5592 19873
rect 5632 19864 5684 19916
rect 1676 19839 1728 19848
rect 1676 19805 1685 19839
rect 1685 19805 1719 19839
rect 1719 19805 1728 19839
rect 1676 19796 1728 19805
rect 5356 19839 5408 19848
rect 5356 19805 5365 19839
rect 5365 19805 5399 19839
rect 5399 19805 5408 19839
rect 5356 19796 5408 19805
rect 3424 19660 3476 19712
rect 6920 19864 6972 19916
rect 6828 19796 6880 19848
rect 7472 19839 7524 19848
rect 7472 19805 7481 19839
rect 7481 19805 7515 19839
rect 7515 19805 7524 19839
rect 7472 19796 7524 19805
rect 8944 19864 8996 19916
rect 9128 19907 9180 19916
rect 9128 19873 9137 19907
rect 9137 19873 9171 19907
rect 9171 19873 9180 19907
rect 9128 19864 9180 19873
rect 11520 19864 11572 19916
rect 12900 19907 12952 19916
rect 12900 19873 12909 19907
rect 12909 19873 12943 19907
rect 12943 19873 12952 19907
rect 12900 19864 12952 19873
rect 13544 19907 13596 19916
rect 8208 19796 8260 19848
rect 9036 19796 9088 19848
rect 9312 19796 9364 19848
rect 10416 19796 10468 19848
rect 10600 19839 10652 19848
rect 10600 19805 10609 19839
rect 10609 19805 10643 19839
rect 10643 19805 10652 19839
rect 10600 19796 10652 19805
rect 13544 19873 13553 19907
rect 13553 19873 13587 19907
rect 13587 19873 13596 19907
rect 13544 19864 13596 19873
rect 14464 19907 14516 19916
rect 14464 19873 14473 19907
rect 14473 19873 14507 19907
rect 14507 19873 14516 19907
rect 14464 19864 14516 19873
rect 13452 19796 13504 19848
rect 14648 19864 14700 19916
rect 15108 19864 15160 19916
rect 16948 19907 17000 19916
rect 16948 19873 16957 19907
rect 16957 19873 16991 19907
rect 16991 19873 17000 19907
rect 16948 19864 17000 19873
rect 17500 19864 17552 19916
rect 17592 19864 17644 19916
rect 19248 19932 19300 19984
rect 19340 19907 19392 19916
rect 17776 19796 17828 19848
rect 19340 19873 19349 19907
rect 19349 19873 19383 19907
rect 19383 19873 19392 19907
rect 19340 19864 19392 19873
rect 20260 19907 20312 19916
rect 20260 19873 20269 19907
rect 20269 19873 20303 19907
rect 20303 19873 20312 19907
rect 20260 19864 20312 19873
rect 22008 20000 22060 20052
rect 25964 20000 26016 20052
rect 26516 20000 26568 20052
rect 27436 20000 27488 20052
rect 30012 20000 30064 20052
rect 21640 19864 21692 19916
rect 21824 19864 21876 19916
rect 25136 19907 25188 19916
rect 8116 19660 8168 19712
rect 9864 19660 9916 19712
rect 16028 19728 16080 19780
rect 19432 19728 19484 19780
rect 23848 19728 23900 19780
rect 24676 19728 24728 19780
rect 25136 19873 25145 19907
rect 25145 19873 25179 19907
rect 25179 19873 25188 19907
rect 25136 19864 25188 19873
rect 25412 19907 25464 19916
rect 25412 19873 25421 19907
rect 25421 19873 25455 19907
rect 25455 19873 25464 19907
rect 25412 19864 25464 19873
rect 25504 19864 25556 19916
rect 26608 19864 26660 19916
rect 27436 19864 27488 19916
rect 28540 19907 28592 19916
rect 28540 19873 28549 19907
rect 28549 19873 28583 19907
rect 28583 19873 28592 19907
rect 28540 19864 28592 19873
rect 29000 19907 29052 19916
rect 29000 19873 29009 19907
rect 29009 19873 29043 19907
rect 29043 19873 29052 19907
rect 29000 19864 29052 19873
rect 32036 19864 32088 19916
rect 34336 19932 34388 19984
rect 35624 20000 35676 20052
rect 27620 19796 27672 19848
rect 29092 19839 29144 19848
rect 29092 19805 29101 19839
rect 29101 19805 29135 19839
rect 29135 19805 29144 19839
rect 29092 19796 29144 19805
rect 14648 19703 14700 19712
rect 14648 19669 14657 19703
rect 14657 19669 14691 19703
rect 14691 19669 14700 19703
rect 14648 19660 14700 19669
rect 14832 19660 14884 19712
rect 16120 19660 16172 19712
rect 18696 19660 18748 19712
rect 22560 19660 22612 19712
rect 22928 19660 22980 19712
rect 25964 19660 26016 19712
rect 27068 19660 27120 19712
rect 27712 19703 27764 19712
rect 27712 19669 27721 19703
rect 27721 19669 27755 19703
rect 27755 19669 27764 19703
rect 27712 19660 27764 19669
rect 29644 19660 29696 19712
rect 29828 19703 29880 19712
rect 29828 19669 29837 19703
rect 29837 19669 29871 19703
rect 29871 19669 29880 19703
rect 29828 19660 29880 19669
rect 30656 19660 30708 19712
rect 32036 19660 32088 19712
rect 33508 19907 33560 19916
rect 33508 19873 33517 19907
rect 33517 19873 33551 19907
rect 33551 19873 33560 19907
rect 33508 19864 33560 19873
rect 33968 19907 34020 19916
rect 33968 19873 33977 19907
rect 33977 19873 34011 19907
rect 34011 19873 34020 19907
rect 33968 19864 34020 19873
rect 35440 19907 35492 19916
rect 35440 19873 35449 19907
rect 35449 19873 35483 19907
rect 35483 19873 35492 19907
rect 35440 19864 35492 19873
rect 35532 19796 35584 19848
rect 33968 19728 34020 19780
rect 35348 19660 35400 19712
rect 35992 19864 36044 19916
rect 38108 19907 38160 19916
rect 38108 19873 38117 19907
rect 38117 19873 38151 19907
rect 38151 19873 38160 19907
rect 38108 19864 38160 19873
rect 38476 19907 38528 19916
rect 38476 19873 38485 19907
rect 38485 19873 38519 19907
rect 38519 19873 38528 19907
rect 38476 19864 38528 19873
rect 38660 19907 38712 19916
rect 38660 19873 38669 19907
rect 38669 19873 38703 19907
rect 38703 19873 38712 19907
rect 38660 19864 38712 19873
rect 37004 19660 37056 19712
rect 4246 19558 4298 19610
rect 4310 19558 4362 19610
rect 4374 19558 4426 19610
rect 4438 19558 4490 19610
rect 34966 19558 35018 19610
rect 35030 19558 35082 19610
rect 35094 19558 35146 19610
rect 35158 19558 35210 19610
rect 1676 19456 1728 19508
rect 4068 19456 4120 19508
rect 9772 19456 9824 19508
rect 11336 19456 11388 19508
rect 15200 19456 15252 19508
rect 16672 19456 16724 19508
rect 18052 19456 18104 19508
rect 27068 19456 27120 19508
rect 3056 19388 3108 19440
rect 7288 19388 7340 19440
rect 9312 19388 9364 19440
rect 24032 19431 24084 19440
rect 24032 19397 24041 19431
rect 24041 19397 24075 19431
rect 24075 19397 24084 19431
rect 24032 19388 24084 19397
rect 28540 19456 28592 19508
rect 34796 19456 34848 19508
rect 35532 19456 35584 19508
rect 7840 19363 7892 19372
rect 7840 19329 7849 19363
rect 7849 19329 7883 19363
rect 7883 19329 7892 19363
rect 7840 19320 7892 19329
rect 3240 19252 3292 19304
rect 3332 19295 3384 19304
rect 3332 19261 3341 19295
rect 3341 19261 3375 19295
rect 3375 19261 3384 19295
rect 3700 19295 3752 19304
rect 3332 19252 3384 19261
rect 3700 19261 3709 19295
rect 3709 19261 3743 19295
rect 3743 19261 3752 19295
rect 3700 19252 3752 19261
rect 4252 19295 4304 19304
rect 4252 19261 4261 19295
rect 4261 19261 4295 19295
rect 4295 19261 4304 19295
rect 4252 19252 4304 19261
rect 4896 19252 4948 19304
rect 5540 19252 5592 19304
rect 5816 19295 5868 19304
rect 5816 19261 5825 19295
rect 5825 19261 5859 19295
rect 5859 19261 5868 19295
rect 5816 19252 5868 19261
rect 7104 19295 7156 19304
rect 7104 19261 7113 19295
rect 7113 19261 7147 19295
rect 7147 19261 7156 19295
rect 7104 19252 7156 19261
rect 2780 19184 2832 19236
rect 6000 19227 6052 19236
rect 6000 19193 6009 19227
rect 6009 19193 6043 19227
rect 6043 19193 6052 19227
rect 6000 19184 6052 19193
rect 7748 19295 7800 19304
rect 7748 19261 7757 19295
rect 7757 19261 7791 19295
rect 7791 19261 7800 19295
rect 7748 19252 7800 19261
rect 8300 19252 8352 19304
rect 9128 19252 9180 19304
rect 9588 19295 9640 19304
rect 9588 19261 9597 19295
rect 9597 19261 9631 19295
rect 9631 19261 9640 19295
rect 9588 19252 9640 19261
rect 10600 19320 10652 19372
rect 13728 19363 13780 19372
rect 9956 19252 10008 19304
rect 10968 19295 11020 19304
rect 10968 19261 10977 19295
rect 10977 19261 11011 19295
rect 11011 19261 11020 19295
rect 10968 19252 11020 19261
rect 3056 19116 3108 19168
rect 3976 19116 4028 19168
rect 7564 19116 7616 19168
rect 7748 19116 7800 19168
rect 8392 19116 8444 19168
rect 13728 19329 13737 19363
rect 13737 19329 13771 19363
rect 13771 19329 13780 19363
rect 13728 19320 13780 19329
rect 12256 19295 12308 19304
rect 12256 19261 12265 19295
rect 12265 19261 12299 19295
rect 12299 19261 12308 19295
rect 12256 19252 12308 19261
rect 12808 19295 12860 19304
rect 12808 19261 12817 19295
rect 12817 19261 12851 19295
rect 12851 19261 12860 19295
rect 12808 19252 12860 19261
rect 13176 19295 13228 19304
rect 13176 19261 13185 19295
rect 13185 19261 13219 19295
rect 13219 19261 13228 19295
rect 13176 19252 13228 19261
rect 14832 19320 14884 19372
rect 12440 19184 12492 19236
rect 16212 19252 16264 19304
rect 16488 19252 16540 19304
rect 16672 19252 16724 19304
rect 15200 19184 15252 19236
rect 18144 19252 18196 19304
rect 18696 19295 18748 19304
rect 18696 19261 18705 19295
rect 18705 19261 18739 19295
rect 18739 19261 18748 19295
rect 18696 19252 18748 19261
rect 18972 19295 19024 19304
rect 18972 19261 18981 19295
rect 18981 19261 19015 19295
rect 19015 19261 19024 19295
rect 18972 19252 19024 19261
rect 19064 19252 19116 19304
rect 21272 19320 21324 19372
rect 21548 19320 21600 19372
rect 28448 19320 28500 19372
rect 20904 19252 20956 19304
rect 21088 19252 21140 19304
rect 23848 19252 23900 19304
rect 24676 19295 24728 19304
rect 24676 19261 24685 19295
rect 24685 19261 24719 19295
rect 24719 19261 24728 19295
rect 24676 19252 24728 19261
rect 25136 19295 25188 19304
rect 25136 19261 25145 19295
rect 25145 19261 25179 19295
rect 25179 19261 25188 19295
rect 25136 19252 25188 19261
rect 25412 19295 25464 19304
rect 25412 19261 25421 19295
rect 25421 19261 25455 19295
rect 25455 19261 25464 19295
rect 25412 19252 25464 19261
rect 25504 19252 25556 19304
rect 26332 19295 26384 19304
rect 26332 19261 26341 19295
rect 26341 19261 26375 19295
rect 26375 19261 26384 19295
rect 26332 19252 26384 19261
rect 27068 19295 27120 19304
rect 27068 19261 27077 19295
rect 27077 19261 27111 19295
rect 27111 19261 27120 19295
rect 27068 19252 27120 19261
rect 27160 19252 27212 19304
rect 29000 19252 29052 19304
rect 29460 19320 29512 19372
rect 32496 19320 32548 19372
rect 33968 19320 34020 19372
rect 30012 19252 30064 19304
rect 31852 19252 31904 19304
rect 32036 19295 32088 19304
rect 32036 19261 32045 19295
rect 32045 19261 32079 19295
rect 32079 19261 32088 19295
rect 32036 19252 32088 19261
rect 32956 19252 33008 19304
rect 34520 19320 34572 19372
rect 36084 19320 36136 19372
rect 23204 19227 23256 19236
rect 18420 19116 18472 19168
rect 23204 19193 23213 19227
rect 23213 19193 23247 19227
rect 23247 19193 23256 19227
rect 23204 19184 23256 19193
rect 26056 19184 26108 19236
rect 33140 19184 33192 19236
rect 36268 19252 36320 19304
rect 37280 19320 37332 19372
rect 37188 19295 37240 19304
rect 37188 19261 37197 19295
rect 37197 19261 37231 19295
rect 37231 19261 37240 19295
rect 37188 19252 37240 19261
rect 38384 19252 38436 19304
rect 19248 19116 19300 19168
rect 19340 19116 19392 19168
rect 21824 19116 21876 19168
rect 22928 19116 22980 19168
rect 27620 19116 27672 19168
rect 28080 19116 28132 19168
rect 29644 19116 29696 19168
rect 35808 19116 35860 19168
rect 38936 19116 38988 19168
rect 19606 19014 19658 19066
rect 19670 19014 19722 19066
rect 19734 19014 19786 19066
rect 19798 19014 19850 19066
rect 3240 18912 3292 18964
rect 2780 18844 2832 18896
rect 3424 18844 3476 18896
rect 5632 18912 5684 18964
rect 9772 18912 9824 18964
rect 9864 18912 9916 18964
rect 2872 18819 2924 18828
rect 2872 18785 2881 18819
rect 2881 18785 2915 18819
rect 2915 18785 2924 18819
rect 2872 18776 2924 18785
rect 2964 18776 3016 18828
rect 3332 18776 3384 18828
rect 3516 18819 3568 18828
rect 3516 18785 3525 18819
rect 3525 18785 3559 18819
rect 3559 18785 3568 18819
rect 3516 18776 3568 18785
rect 5724 18819 5776 18828
rect 4252 18708 4304 18760
rect 5356 18640 5408 18692
rect 5724 18785 5733 18819
rect 5733 18785 5767 18819
rect 5767 18785 5776 18819
rect 5724 18776 5776 18785
rect 6000 18776 6052 18828
rect 7748 18819 7800 18828
rect 7748 18785 7757 18819
rect 7757 18785 7791 18819
rect 7791 18785 7800 18819
rect 7748 18776 7800 18785
rect 8300 18776 8352 18828
rect 5908 18751 5960 18760
rect 5908 18717 5917 18751
rect 5917 18717 5951 18751
rect 5951 18717 5960 18751
rect 5908 18708 5960 18717
rect 8576 18708 8628 18760
rect 9588 18844 9640 18896
rect 9680 18844 9732 18896
rect 10048 18912 10100 18964
rect 14740 18912 14792 18964
rect 15568 18955 15620 18964
rect 15568 18921 15577 18955
rect 15577 18921 15611 18955
rect 15611 18921 15620 18955
rect 15568 18912 15620 18921
rect 16212 18912 16264 18964
rect 23204 18912 23256 18964
rect 26700 18955 26752 18964
rect 26700 18921 26709 18955
rect 26709 18921 26743 18955
rect 26743 18921 26752 18955
rect 26700 18912 26752 18921
rect 27896 18912 27948 18964
rect 34152 18912 34204 18964
rect 12808 18844 12860 18896
rect 14096 18844 14148 18896
rect 14648 18844 14700 18896
rect 18972 18844 19024 18896
rect 13360 18776 13412 18828
rect 13820 18819 13872 18828
rect 13820 18785 13829 18819
rect 13829 18785 13863 18819
rect 13863 18785 13872 18819
rect 13820 18776 13872 18785
rect 14464 18819 14516 18828
rect 14464 18785 14473 18819
rect 14473 18785 14507 18819
rect 14507 18785 14516 18819
rect 14464 18776 14516 18785
rect 2228 18572 2280 18624
rect 3884 18572 3936 18624
rect 5724 18572 5776 18624
rect 6092 18572 6144 18624
rect 10048 18708 10100 18760
rect 11060 18751 11112 18760
rect 9864 18640 9916 18692
rect 10600 18640 10652 18692
rect 11060 18717 11069 18751
rect 11069 18717 11103 18751
rect 11103 18717 11112 18751
rect 11060 18708 11112 18717
rect 12716 18708 12768 18760
rect 13084 18708 13136 18760
rect 13912 18708 13964 18760
rect 15936 18776 15988 18828
rect 19064 18776 19116 18828
rect 19340 18819 19392 18828
rect 19340 18785 19349 18819
rect 19349 18785 19383 18819
rect 19383 18785 19392 18819
rect 19340 18776 19392 18785
rect 19524 18776 19576 18828
rect 19708 18776 19760 18828
rect 17960 18708 18012 18760
rect 18328 18708 18380 18760
rect 19248 18708 19300 18760
rect 18052 18640 18104 18692
rect 19984 18751 20036 18760
rect 19984 18717 19993 18751
rect 19993 18717 20027 18751
rect 20027 18717 20036 18751
rect 21088 18844 21140 18896
rect 21364 18844 21416 18896
rect 21824 18844 21876 18896
rect 22008 18887 22060 18896
rect 22008 18853 22017 18887
rect 22017 18853 22051 18887
rect 22051 18853 22060 18887
rect 22008 18844 22060 18853
rect 23848 18844 23900 18896
rect 19984 18708 20036 18717
rect 22468 18776 22520 18828
rect 22100 18708 22152 18760
rect 22284 18708 22336 18760
rect 21180 18640 21232 18692
rect 22836 18776 22888 18828
rect 23204 18776 23256 18828
rect 24860 18844 24912 18896
rect 24400 18776 24452 18828
rect 25228 18819 25280 18828
rect 25228 18785 25237 18819
rect 25237 18785 25271 18819
rect 25271 18785 25280 18819
rect 25228 18776 25280 18785
rect 26240 18776 26292 18828
rect 24308 18708 24360 18760
rect 24860 18751 24912 18760
rect 24860 18717 24869 18751
rect 24869 18717 24903 18751
rect 24903 18717 24912 18751
rect 24860 18708 24912 18717
rect 26148 18708 26200 18760
rect 28080 18776 28132 18828
rect 28540 18776 28592 18828
rect 29736 18776 29788 18828
rect 30196 18819 30248 18828
rect 30196 18785 30205 18819
rect 30205 18785 30239 18819
rect 30239 18785 30248 18819
rect 30196 18776 30248 18785
rect 30656 18819 30708 18828
rect 29092 18708 29144 18760
rect 29552 18751 29604 18760
rect 29552 18717 29561 18751
rect 29561 18717 29595 18751
rect 29595 18717 29604 18751
rect 29552 18708 29604 18717
rect 30656 18785 30665 18819
rect 30665 18785 30699 18819
rect 30699 18785 30708 18819
rect 30656 18776 30708 18785
rect 31852 18776 31904 18828
rect 32036 18776 32088 18828
rect 32496 18819 32548 18828
rect 32496 18785 32505 18819
rect 32505 18785 32539 18819
rect 32539 18785 32548 18819
rect 32496 18776 32548 18785
rect 32956 18819 33008 18828
rect 32956 18785 32965 18819
rect 32965 18785 32999 18819
rect 32999 18785 33008 18819
rect 32956 18776 33008 18785
rect 33048 18776 33100 18828
rect 34796 18844 34848 18896
rect 34520 18819 34572 18828
rect 34520 18785 34529 18819
rect 34529 18785 34563 18819
rect 34563 18785 34572 18819
rect 34520 18776 34572 18785
rect 34704 18776 34756 18828
rect 35900 18776 35952 18828
rect 36912 18887 36964 18896
rect 36912 18853 36921 18887
rect 36921 18853 36955 18887
rect 36955 18853 36964 18887
rect 36912 18844 36964 18853
rect 38384 18844 38436 18896
rect 34612 18751 34664 18760
rect 34612 18717 34621 18751
rect 34621 18717 34655 18751
rect 34655 18717 34664 18751
rect 34612 18708 34664 18717
rect 38108 18776 38160 18828
rect 38476 18776 38528 18828
rect 38200 18708 38252 18760
rect 23204 18640 23256 18692
rect 23848 18640 23900 18692
rect 25504 18683 25556 18692
rect 25504 18649 25513 18683
rect 25513 18649 25547 18683
rect 25547 18649 25556 18683
rect 25504 18640 25556 18649
rect 29368 18640 29420 18692
rect 33048 18640 33100 18692
rect 38660 18640 38712 18692
rect 9772 18572 9824 18624
rect 17868 18572 17920 18624
rect 18420 18572 18472 18624
rect 19984 18572 20036 18624
rect 21640 18572 21692 18624
rect 27344 18615 27396 18624
rect 27344 18581 27353 18615
rect 27353 18581 27387 18615
rect 27387 18581 27396 18615
rect 27344 18572 27396 18581
rect 27436 18572 27488 18624
rect 31944 18572 31996 18624
rect 35900 18572 35952 18624
rect 4246 18470 4298 18522
rect 4310 18470 4362 18522
rect 4374 18470 4426 18522
rect 4438 18470 4490 18522
rect 34966 18470 35018 18522
rect 35030 18470 35082 18522
rect 35094 18470 35146 18522
rect 35158 18470 35210 18522
rect 9772 18368 9824 18420
rect 9956 18368 10008 18420
rect 12348 18368 12400 18420
rect 4620 18300 4672 18352
rect 6828 18300 6880 18352
rect 7840 18300 7892 18352
rect 10324 18300 10376 18352
rect 13912 18300 13964 18352
rect 2872 18232 2924 18284
rect 2780 18207 2832 18216
rect 2780 18173 2789 18207
rect 2789 18173 2823 18207
rect 2823 18173 2832 18207
rect 3516 18207 3568 18216
rect 2780 18164 2832 18173
rect 3516 18173 3525 18207
rect 3525 18173 3559 18207
rect 3559 18173 3568 18207
rect 3516 18164 3568 18173
rect 5448 18232 5500 18284
rect 5632 18207 5684 18216
rect 3516 18028 3568 18080
rect 4712 18096 4764 18148
rect 5632 18173 5641 18207
rect 5641 18173 5675 18207
rect 5675 18173 5684 18207
rect 5632 18164 5684 18173
rect 5816 18096 5868 18148
rect 7196 18207 7248 18216
rect 6920 18096 6972 18148
rect 7196 18173 7205 18207
rect 7205 18173 7239 18207
rect 7239 18173 7248 18207
rect 7196 18164 7248 18173
rect 14832 18232 14884 18284
rect 15200 18275 15252 18284
rect 15200 18241 15209 18275
rect 15209 18241 15243 18275
rect 15243 18241 15252 18275
rect 15200 18232 15252 18241
rect 8392 18207 8444 18216
rect 8392 18173 8401 18207
rect 8401 18173 8435 18207
rect 8435 18173 8444 18207
rect 8392 18164 8444 18173
rect 8116 18096 8168 18148
rect 8300 18096 8352 18148
rect 10232 18164 10284 18216
rect 12624 18207 12676 18216
rect 12624 18173 12633 18207
rect 12633 18173 12667 18207
rect 12667 18173 12676 18207
rect 12624 18164 12676 18173
rect 10416 18028 10468 18080
rect 12256 18096 12308 18148
rect 14096 18164 14148 18216
rect 14188 18096 14240 18148
rect 15292 18164 15344 18216
rect 15936 18164 15988 18216
rect 17868 18368 17920 18420
rect 19524 18368 19576 18420
rect 19708 18368 19760 18420
rect 22284 18368 22336 18420
rect 22836 18368 22888 18420
rect 29276 18368 29328 18420
rect 35716 18368 35768 18420
rect 36636 18368 36688 18420
rect 39028 18368 39080 18420
rect 21180 18300 21232 18352
rect 22192 18300 22244 18352
rect 23940 18343 23992 18352
rect 23940 18309 23949 18343
rect 23949 18309 23983 18343
rect 23983 18309 23992 18343
rect 23940 18300 23992 18309
rect 29460 18343 29512 18352
rect 29460 18309 29469 18343
rect 29469 18309 29503 18343
rect 29503 18309 29512 18343
rect 29460 18300 29512 18309
rect 32956 18343 33008 18352
rect 32956 18309 32965 18343
rect 32965 18309 32999 18343
rect 32999 18309 33008 18343
rect 32956 18300 33008 18309
rect 34336 18300 34388 18352
rect 18696 18232 18748 18284
rect 23848 18275 23900 18284
rect 18144 18164 18196 18216
rect 18328 18207 18380 18216
rect 18328 18173 18337 18207
rect 18337 18173 18371 18207
rect 18371 18173 18380 18207
rect 18328 18164 18380 18173
rect 20444 18207 20496 18216
rect 20444 18173 20453 18207
rect 20453 18173 20487 18207
rect 20487 18173 20496 18207
rect 20444 18164 20496 18173
rect 12440 18028 12492 18080
rect 14924 18028 14976 18080
rect 16120 18028 16172 18080
rect 16304 18071 16356 18080
rect 16304 18037 16313 18071
rect 16313 18037 16347 18071
rect 16347 18037 16356 18071
rect 16304 18028 16356 18037
rect 17408 18071 17460 18080
rect 17408 18037 17417 18071
rect 17417 18037 17451 18071
rect 17451 18037 17460 18071
rect 17408 18028 17460 18037
rect 19340 18028 19392 18080
rect 23848 18241 23857 18275
rect 23857 18241 23891 18275
rect 23891 18241 23900 18275
rect 23848 18232 23900 18241
rect 27160 18275 27212 18284
rect 27160 18241 27169 18275
rect 27169 18241 27203 18275
rect 27203 18241 27212 18275
rect 27160 18232 27212 18241
rect 22560 18207 22612 18216
rect 22560 18173 22569 18207
rect 22569 18173 22603 18207
rect 22603 18173 22612 18207
rect 22560 18164 22612 18173
rect 22744 18164 22796 18216
rect 24676 18164 24728 18216
rect 25136 18164 25188 18216
rect 25320 18207 25372 18216
rect 25320 18173 25329 18207
rect 25329 18173 25363 18207
rect 25363 18173 25372 18207
rect 25320 18164 25372 18173
rect 25504 18207 25556 18216
rect 25504 18173 25513 18207
rect 25513 18173 25547 18207
rect 25547 18173 25556 18207
rect 25504 18164 25556 18173
rect 26516 18207 26568 18216
rect 26516 18173 26525 18207
rect 26525 18173 26559 18207
rect 26559 18173 26568 18207
rect 26516 18164 26568 18173
rect 27344 18164 27396 18216
rect 30196 18232 30248 18284
rect 33600 18275 33652 18284
rect 28632 18207 28684 18216
rect 22008 18096 22060 18148
rect 23204 18096 23256 18148
rect 28632 18173 28641 18207
rect 28641 18173 28675 18207
rect 28675 18173 28684 18207
rect 28632 18164 28684 18173
rect 29276 18207 29328 18216
rect 29276 18173 29285 18207
rect 29285 18173 29319 18207
rect 29319 18173 29328 18207
rect 29276 18164 29328 18173
rect 29552 18164 29604 18216
rect 30840 18164 30892 18216
rect 33140 18207 33192 18216
rect 22100 18028 22152 18080
rect 27988 18028 28040 18080
rect 29092 18096 29144 18148
rect 28724 18028 28776 18080
rect 30288 18028 30340 18080
rect 33140 18173 33149 18207
rect 33149 18173 33183 18207
rect 33183 18173 33192 18207
rect 33140 18164 33192 18173
rect 33600 18241 33609 18275
rect 33609 18241 33643 18275
rect 33643 18241 33652 18275
rect 33600 18232 33652 18241
rect 34428 18232 34480 18284
rect 36084 18232 36136 18284
rect 38568 18275 38620 18284
rect 38568 18241 38577 18275
rect 38577 18241 38611 18275
rect 38611 18241 38620 18275
rect 38568 18232 38620 18241
rect 33508 18207 33560 18216
rect 33508 18173 33517 18207
rect 33517 18173 33551 18207
rect 33551 18173 33560 18207
rect 33508 18164 33560 18173
rect 33692 18164 33744 18216
rect 34796 18164 34848 18216
rect 35992 18207 36044 18216
rect 35992 18173 36001 18207
rect 36001 18173 36035 18207
rect 36035 18173 36044 18207
rect 35992 18164 36044 18173
rect 38200 18207 38252 18216
rect 38200 18173 38209 18207
rect 38209 18173 38243 18207
rect 38243 18173 38252 18207
rect 38200 18164 38252 18173
rect 38384 18207 38436 18216
rect 38384 18173 38393 18207
rect 38393 18173 38427 18207
rect 38427 18173 38436 18207
rect 38384 18164 38436 18173
rect 38660 18207 38712 18216
rect 38660 18173 38669 18207
rect 38669 18173 38703 18207
rect 38703 18173 38712 18207
rect 38660 18164 38712 18173
rect 34520 18096 34572 18148
rect 32864 18028 32916 18080
rect 38568 18096 38620 18148
rect 19606 17926 19658 17978
rect 19670 17926 19722 17978
rect 19734 17926 19786 17978
rect 19798 17926 19850 17978
rect 5448 17824 5500 17876
rect 3884 17756 3936 17808
rect 10324 17824 10376 17876
rect 13084 17824 13136 17876
rect 24032 17824 24084 17876
rect 25780 17824 25832 17876
rect 32404 17867 32456 17876
rect 32404 17833 32413 17867
rect 32413 17833 32447 17867
rect 32447 17833 32456 17867
rect 32404 17824 32456 17833
rect 35348 17824 35400 17876
rect 1400 17688 1452 17740
rect 3976 17688 4028 17740
rect 4896 17731 4948 17740
rect 4896 17697 4905 17731
rect 4905 17697 4939 17731
rect 4939 17697 4948 17731
rect 4896 17688 4948 17697
rect 5356 17731 5408 17740
rect 5356 17697 5365 17731
rect 5365 17697 5399 17731
rect 5399 17697 5408 17731
rect 5356 17688 5408 17697
rect 5908 17688 5960 17740
rect 6092 17731 6144 17740
rect 6092 17697 6101 17731
rect 6101 17697 6135 17731
rect 6135 17697 6144 17731
rect 6092 17688 6144 17697
rect 7104 17731 7156 17740
rect 1768 17663 1820 17672
rect 1768 17629 1777 17663
rect 1777 17629 1811 17663
rect 1811 17629 1820 17663
rect 1768 17620 1820 17629
rect 7104 17697 7113 17731
rect 7113 17697 7147 17731
rect 7147 17697 7156 17731
rect 7104 17688 7156 17697
rect 7656 17731 7708 17740
rect 7656 17697 7665 17731
rect 7665 17697 7699 17731
rect 7699 17697 7708 17731
rect 7656 17688 7708 17697
rect 9220 17756 9272 17808
rect 8576 17731 8628 17740
rect 8576 17697 8585 17731
rect 8585 17697 8619 17731
rect 8619 17697 8628 17731
rect 8576 17688 8628 17697
rect 11060 17756 11112 17808
rect 17960 17756 18012 17808
rect 10416 17731 10468 17740
rect 10416 17697 10425 17731
rect 10425 17697 10459 17731
rect 10459 17697 10468 17731
rect 10416 17688 10468 17697
rect 13912 17731 13964 17740
rect 13912 17697 13921 17731
rect 13921 17697 13955 17731
rect 13955 17697 13964 17731
rect 13912 17688 13964 17697
rect 14188 17688 14240 17740
rect 15292 17731 15344 17740
rect 15292 17697 15301 17731
rect 15301 17697 15335 17731
rect 15335 17697 15344 17731
rect 15292 17688 15344 17697
rect 17592 17731 17644 17740
rect 17592 17697 17601 17731
rect 17601 17697 17635 17731
rect 17635 17697 17644 17731
rect 17592 17688 17644 17697
rect 17776 17688 17828 17740
rect 18880 17688 18932 17740
rect 20076 17688 20128 17740
rect 11244 17620 11296 17672
rect 11612 17663 11664 17672
rect 8300 17552 8352 17604
rect 9772 17552 9824 17604
rect 11612 17629 11621 17663
rect 11621 17629 11655 17663
rect 11655 17629 11664 17663
rect 11612 17620 11664 17629
rect 13636 17663 13688 17672
rect 13636 17629 13645 17663
rect 13645 17629 13679 17663
rect 13679 17629 13688 17663
rect 13636 17620 13688 17629
rect 15568 17663 15620 17672
rect 15568 17629 15577 17663
rect 15577 17629 15611 17663
rect 15611 17629 15620 17663
rect 15568 17620 15620 17629
rect 18604 17663 18656 17672
rect 18604 17629 18613 17663
rect 18613 17629 18647 17663
rect 18647 17629 18656 17663
rect 18604 17620 18656 17629
rect 14004 17552 14056 17604
rect 17408 17552 17460 17604
rect 21088 17620 21140 17672
rect 19156 17552 19208 17604
rect 21732 17688 21784 17740
rect 3976 17484 4028 17536
rect 8116 17484 8168 17536
rect 12900 17527 12952 17536
rect 12900 17493 12909 17527
rect 12909 17493 12943 17527
rect 12943 17493 12952 17527
rect 12900 17484 12952 17493
rect 16672 17527 16724 17536
rect 16672 17493 16681 17527
rect 16681 17493 16715 17527
rect 16715 17493 16724 17527
rect 16672 17484 16724 17493
rect 17868 17527 17920 17536
rect 17868 17493 17877 17527
rect 17877 17493 17911 17527
rect 17911 17493 17920 17527
rect 17868 17484 17920 17493
rect 18328 17484 18380 17536
rect 22100 17484 22152 17536
rect 22744 17756 22796 17808
rect 24216 17756 24268 17808
rect 22928 17688 22980 17740
rect 23848 17731 23900 17740
rect 23848 17697 23857 17731
rect 23857 17697 23891 17731
rect 23891 17697 23900 17731
rect 23848 17688 23900 17697
rect 24676 17688 24728 17740
rect 25136 17688 25188 17740
rect 25320 17731 25372 17740
rect 25320 17697 25329 17731
rect 25329 17697 25363 17731
rect 25363 17697 25372 17731
rect 25320 17688 25372 17697
rect 25504 17731 25556 17740
rect 25504 17697 25513 17731
rect 25513 17697 25547 17731
rect 25547 17697 25556 17731
rect 25504 17688 25556 17697
rect 26792 17731 26844 17740
rect 26792 17697 26801 17731
rect 26801 17697 26835 17731
rect 26835 17697 26844 17731
rect 26792 17688 26844 17697
rect 26976 17688 27028 17740
rect 23756 17552 23808 17604
rect 26424 17620 26476 17672
rect 26608 17595 26660 17604
rect 26608 17561 26617 17595
rect 26617 17561 26651 17595
rect 26651 17561 26660 17595
rect 26608 17552 26660 17561
rect 27068 17552 27120 17604
rect 27712 17552 27764 17604
rect 24124 17484 24176 17536
rect 24308 17484 24360 17536
rect 25228 17484 25280 17536
rect 28632 17688 28684 17740
rect 28816 17688 28868 17740
rect 30196 17756 30248 17808
rect 31116 17731 31168 17740
rect 29092 17663 29144 17672
rect 29092 17629 29101 17663
rect 29101 17629 29135 17663
rect 29135 17629 29144 17663
rect 29092 17620 29144 17629
rect 31116 17697 31125 17731
rect 31125 17697 31159 17731
rect 31159 17697 31168 17731
rect 31116 17688 31168 17697
rect 34520 17756 34572 17808
rect 32312 17731 32364 17740
rect 32312 17697 32321 17731
rect 32321 17697 32355 17731
rect 32355 17697 32364 17731
rect 32312 17688 32364 17697
rect 32680 17731 32732 17740
rect 32680 17697 32689 17731
rect 32689 17697 32723 17731
rect 32723 17697 32732 17731
rect 32680 17688 32732 17697
rect 33600 17688 33652 17740
rect 33692 17688 33744 17740
rect 34612 17731 34664 17740
rect 34612 17697 34621 17731
rect 34621 17697 34655 17731
rect 34655 17697 34664 17731
rect 34612 17688 34664 17697
rect 34796 17731 34848 17740
rect 34796 17697 34805 17731
rect 34805 17697 34839 17731
rect 34839 17697 34848 17731
rect 34796 17688 34848 17697
rect 36452 17756 36504 17808
rect 30012 17620 30064 17672
rect 30196 17620 30248 17672
rect 36360 17688 36412 17740
rect 38568 17731 38620 17740
rect 35808 17620 35860 17672
rect 38568 17697 38577 17731
rect 38577 17697 38611 17731
rect 38611 17697 38620 17731
rect 38568 17688 38620 17697
rect 38844 17620 38896 17672
rect 32496 17484 32548 17536
rect 34796 17484 34848 17536
rect 35532 17484 35584 17536
rect 35716 17527 35768 17536
rect 35716 17493 35725 17527
rect 35725 17493 35759 17527
rect 35759 17493 35768 17527
rect 35716 17484 35768 17493
rect 36268 17484 36320 17536
rect 36544 17552 36596 17604
rect 37556 17484 37608 17536
rect 4246 17382 4298 17434
rect 4310 17382 4362 17434
rect 4374 17382 4426 17434
rect 4438 17382 4490 17434
rect 34966 17382 35018 17434
rect 35030 17382 35082 17434
rect 35094 17382 35146 17434
rect 35158 17382 35210 17434
rect 2780 17280 2832 17332
rect 4712 17280 4764 17332
rect 6920 17323 6972 17332
rect 6920 17289 6929 17323
rect 6929 17289 6963 17323
rect 6963 17289 6972 17323
rect 6920 17280 6972 17289
rect 9220 17323 9272 17332
rect 9220 17289 9229 17323
rect 9229 17289 9263 17323
rect 9263 17289 9272 17323
rect 9220 17280 9272 17289
rect 10232 17323 10284 17332
rect 10232 17289 10241 17323
rect 10241 17289 10275 17323
rect 10275 17289 10284 17323
rect 10232 17280 10284 17289
rect 11612 17323 11664 17332
rect 11612 17289 11621 17323
rect 11621 17289 11655 17323
rect 11655 17289 11664 17323
rect 11612 17280 11664 17289
rect 14740 17280 14792 17332
rect 10048 17212 10100 17264
rect 3056 17187 3108 17196
rect 3056 17153 3065 17187
rect 3065 17153 3099 17187
rect 3099 17153 3108 17187
rect 3056 17144 3108 17153
rect 1952 17076 2004 17128
rect 2228 17119 2280 17128
rect 2228 17085 2237 17119
rect 2237 17085 2271 17119
rect 2271 17085 2280 17119
rect 2228 17076 2280 17085
rect 2780 17076 2832 17128
rect 4620 17144 4672 17196
rect 4712 17144 4764 17196
rect 6184 17187 6236 17196
rect 3424 17119 3476 17128
rect 3424 17085 3433 17119
rect 3433 17085 3467 17119
rect 3467 17085 3476 17119
rect 3424 17076 3476 17085
rect 3976 17119 4028 17128
rect 3976 17085 3985 17119
rect 3985 17085 4019 17119
rect 4019 17085 4028 17119
rect 3976 17076 4028 17085
rect 4896 17119 4948 17128
rect 4896 17085 4905 17119
rect 4905 17085 4939 17119
rect 4939 17085 4948 17119
rect 4896 17076 4948 17085
rect 5448 17119 5500 17128
rect 5448 17085 5457 17119
rect 5457 17085 5491 17119
rect 5491 17085 5500 17119
rect 5448 17076 5500 17085
rect 6184 17153 6193 17187
rect 6193 17153 6227 17187
rect 6227 17153 6236 17187
rect 6184 17144 6236 17153
rect 11244 17144 11296 17196
rect 6276 17119 6328 17128
rect 6276 17085 6285 17119
rect 6285 17085 6319 17119
rect 6319 17085 6328 17119
rect 6276 17076 6328 17085
rect 7840 17119 7892 17128
rect 7840 17085 7849 17119
rect 7849 17085 7883 17119
rect 7883 17085 7892 17119
rect 7840 17076 7892 17085
rect 8576 17076 8628 17128
rect 10692 17076 10744 17128
rect 11428 17119 11480 17128
rect 11428 17085 11437 17119
rect 11437 17085 11471 17119
rect 11471 17085 11480 17119
rect 12716 17119 12768 17128
rect 11428 17076 11480 17085
rect 12716 17085 12725 17119
rect 12725 17085 12759 17119
rect 12759 17085 12768 17119
rect 12716 17076 12768 17085
rect 12900 17119 12952 17128
rect 12900 17085 12909 17119
rect 12909 17085 12943 17119
rect 12943 17085 12952 17119
rect 12900 17076 12952 17085
rect 13820 17212 13872 17264
rect 15844 17255 15896 17264
rect 13636 17187 13688 17196
rect 13636 17153 13645 17187
rect 13645 17153 13679 17187
rect 13679 17153 13688 17187
rect 13636 17144 13688 17153
rect 15292 17144 15344 17196
rect 14924 17119 14976 17128
rect 14924 17085 14933 17119
rect 14933 17085 14967 17119
rect 14967 17085 14976 17119
rect 14924 17076 14976 17085
rect 15200 17076 15252 17128
rect 15844 17221 15853 17255
rect 15853 17221 15887 17255
rect 15887 17221 15896 17255
rect 15844 17212 15896 17221
rect 16120 17280 16172 17332
rect 18604 17212 18656 17264
rect 18696 17144 18748 17196
rect 19156 17187 19208 17196
rect 19156 17153 19165 17187
rect 19165 17153 19199 17187
rect 19199 17153 19208 17187
rect 19156 17144 19208 17153
rect 16672 17119 16724 17128
rect 16672 17085 16681 17119
rect 16681 17085 16715 17119
rect 16715 17085 16724 17119
rect 16672 17076 16724 17085
rect 17224 17119 17276 17128
rect 17224 17085 17233 17119
rect 17233 17085 17267 17119
rect 17267 17085 17276 17119
rect 17224 17076 17276 17085
rect 18144 17076 18196 17128
rect 23480 17280 23532 17332
rect 26516 17280 26568 17332
rect 27528 17280 27580 17332
rect 28356 17280 28408 17332
rect 22652 17255 22704 17264
rect 22652 17221 22661 17255
rect 22661 17221 22695 17255
rect 22695 17221 22704 17255
rect 22652 17212 22704 17221
rect 24032 17212 24084 17264
rect 25688 17212 25740 17264
rect 33140 17280 33192 17332
rect 34612 17280 34664 17332
rect 38108 17280 38160 17332
rect 38568 17280 38620 17332
rect 21364 17144 21416 17196
rect 21640 17076 21692 17128
rect 22744 17144 22796 17196
rect 24492 17144 24544 17196
rect 22008 17076 22060 17128
rect 22192 17076 22244 17128
rect 23572 17076 23624 17128
rect 24400 17076 24452 17128
rect 26148 17119 26200 17128
rect 6552 17008 6604 17060
rect 1768 16940 1820 16992
rect 11244 16940 11296 16992
rect 15476 17008 15528 17060
rect 17408 17008 17460 17060
rect 20168 17008 20220 17060
rect 26148 17085 26157 17119
rect 26157 17085 26191 17119
rect 26191 17085 26200 17119
rect 26148 17076 26200 17085
rect 26240 17119 26292 17128
rect 26240 17085 26249 17119
rect 26249 17085 26283 17119
rect 26283 17085 26292 17119
rect 26792 17144 26844 17196
rect 28816 17144 28868 17196
rect 34336 17212 34388 17264
rect 32404 17187 32456 17196
rect 26240 17076 26292 17085
rect 27528 17076 27580 17128
rect 27988 17119 28040 17128
rect 27988 17085 27997 17119
rect 27997 17085 28031 17119
rect 28031 17085 28040 17119
rect 27988 17076 28040 17085
rect 28080 17119 28132 17128
rect 28080 17085 28089 17119
rect 28089 17085 28123 17119
rect 28123 17085 28132 17119
rect 28080 17076 28132 17085
rect 27436 17008 27488 17060
rect 27712 17008 27764 17060
rect 28448 17119 28500 17128
rect 28448 17085 28457 17119
rect 28457 17085 28491 17119
rect 28491 17085 28500 17119
rect 29552 17119 29604 17128
rect 28448 17076 28500 17085
rect 29552 17085 29561 17119
rect 29561 17085 29595 17119
rect 29595 17085 29604 17119
rect 29552 17076 29604 17085
rect 30012 17119 30064 17128
rect 30012 17085 30021 17119
rect 30021 17085 30055 17119
rect 30055 17085 30064 17119
rect 30012 17076 30064 17085
rect 30288 17119 30340 17128
rect 30288 17085 30297 17119
rect 30297 17085 30331 17119
rect 30331 17085 30340 17119
rect 30288 17076 30340 17085
rect 31944 17076 31996 17128
rect 32128 17119 32180 17128
rect 32128 17085 32137 17119
rect 32137 17085 32171 17119
rect 32171 17085 32180 17119
rect 32128 17076 32180 17085
rect 32404 17153 32413 17187
rect 32413 17153 32447 17187
rect 32447 17153 32456 17187
rect 32404 17144 32456 17153
rect 32772 17076 32824 17128
rect 35808 17144 35860 17196
rect 36360 17144 36412 17196
rect 34520 17076 34572 17128
rect 35348 17119 35400 17128
rect 35348 17085 35357 17119
rect 35357 17085 35391 17119
rect 35391 17085 35400 17119
rect 35348 17076 35400 17085
rect 35716 17119 35768 17128
rect 35716 17085 35725 17119
rect 35725 17085 35759 17119
rect 35759 17085 35768 17119
rect 35716 17076 35768 17085
rect 36084 17076 36136 17128
rect 37188 17144 37240 17196
rect 37832 17076 37884 17128
rect 38660 17119 38712 17128
rect 38660 17085 38669 17119
rect 38669 17085 38703 17119
rect 38703 17085 38712 17119
rect 38660 17076 38712 17085
rect 13544 16940 13596 16992
rect 17500 16940 17552 16992
rect 20628 16940 20680 16992
rect 24308 16983 24360 16992
rect 24308 16949 24317 16983
rect 24317 16949 24351 16983
rect 24351 16949 24360 16983
rect 24308 16940 24360 16949
rect 24768 16940 24820 16992
rect 24952 16983 25004 16992
rect 24952 16949 24961 16983
rect 24961 16949 24995 16983
rect 24995 16949 25004 16983
rect 24952 16940 25004 16949
rect 25688 16940 25740 16992
rect 27528 16940 27580 16992
rect 30380 16940 30432 16992
rect 33968 16940 34020 16992
rect 34612 16940 34664 16992
rect 36452 16940 36504 16992
rect 19606 16838 19658 16890
rect 19670 16838 19722 16890
rect 19734 16838 19786 16890
rect 19798 16838 19850 16890
rect 4804 16736 4856 16788
rect 5356 16736 5408 16788
rect 8208 16736 8260 16788
rect 11428 16736 11480 16788
rect 12716 16736 12768 16788
rect 3056 16600 3108 16652
rect 3332 16643 3384 16652
rect 3332 16609 3341 16643
rect 3341 16609 3375 16643
rect 3375 16609 3384 16643
rect 3332 16600 3384 16609
rect 8576 16711 8628 16720
rect 8576 16677 8585 16711
rect 8585 16677 8619 16711
rect 8619 16677 8628 16711
rect 8576 16668 8628 16677
rect 14004 16736 14056 16788
rect 19984 16736 20036 16788
rect 20720 16736 20772 16788
rect 22008 16736 22060 16788
rect 6184 16643 6236 16652
rect 6184 16609 6193 16643
rect 6193 16609 6227 16643
rect 6227 16609 6236 16643
rect 6184 16600 6236 16609
rect 6552 16643 6604 16652
rect 6552 16609 6561 16643
rect 6561 16609 6595 16643
rect 6595 16609 6604 16643
rect 6552 16600 6604 16609
rect 7196 16643 7248 16652
rect 7196 16609 7205 16643
rect 7205 16609 7239 16643
rect 7239 16609 7248 16643
rect 7196 16600 7248 16609
rect 8116 16643 8168 16652
rect 3516 16532 3568 16584
rect 3976 16464 4028 16516
rect 4436 16532 4488 16584
rect 8116 16609 8125 16643
rect 8125 16609 8159 16643
rect 8159 16609 8168 16643
rect 8116 16600 8168 16609
rect 8392 16600 8444 16652
rect 9956 16600 10008 16652
rect 17868 16668 17920 16720
rect 29000 16736 29052 16788
rect 15476 16643 15528 16652
rect 15476 16609 15485 16643
rect 15485 16609 15519 16643
rect 15519 16609 15528 16643
rect 15476 16600 15528 16609
rect 16304 16600 16356 16652
rect 17500 16600 17552 16652
rect 17684 16643 17736 16652
rect 17684 16609 17693 16643
rect 17693 16609 17727 16643
rect 17727 16609 17736 16643
rect 17684 16600 17736 16609
rect 18420 16643 18472 16652
rect 18420 16609 18429 16643
rect 18429 16609 18463 16643
rect 18463 16609 18472 16643
rect 18420 16600 18472 16609
rect 18512 16600 18564 16652
rect 20168 16643 20220 16652
rect 20168 16609 20177 16643
rect 20177 16609 20211 16643
rect 20211 16609 20220 16643
rect 20168 16600 20220 16609
rect 21640 16600 21692 16652
rect 22008 16643 22060 16652
rect 22008 16609 22017 16643
rect 22017 16609 22051 16643
rect 22051 16609 22060 16643
rect 22008 16600 22060 16609
rect 12532 16532 12584 16584
rect 13084 16575 13136 16584
rect 13084 16541 13093 16575
rect 13093 16541 13127 16575
rect 13127 16541 13136 16575
rect 13084 16532 13136 16541
rect 15292 16532 15344 16584
rect 17040 16532 17092 16584
rect 18328 16532 18380 16584
rect 19340 16575 19392 16584
rect 19340 16541 19349 16575
rect 19349 16541 19383 16575
rect 19383 16541 19392 16575
rect 19340 16532 19392 16541
rect 20720 16532 20772 16584
rect 24032 16668 24084 16720
rect 24952 16668 25004 16720
rect 22744 16643 22796 16652
rect 22744 16609 22753 16643
rect 22753 16609 22787 16643
rect 22787 16609 22796 16643
rect 22744 16600 22796 16609
rect 23756 16643 23808 16652
rect 23756 16609 23765 16643
rect 23765 16609 23799 16643
rect 23799 16609 23808 16643
rect 23756 16600 23808 16609
rect 24400 16600 24452 16652
rect 24860 16643 24912 16652
rect 24860 16609 24869 16643
rect 24869 16609 24903 16643
rect 24903 16609 24912 16643
rect 24860 16600 24912 16609
rect 25320 16643 25372 16652
rect 25320 16609 25329 16643
rect 25329 16609 25363 16643
rect 25363 16609 25372 16643
rect 25320 16600 25372 16609
rect 25780 16643 25832 16652
rect 25780 16609 25789 16643
rect 25789 16609 25823 16643
rect 25823 16609 25832 16643
rect 25780 16600 25832 16609
rect 26792 16600 26844 16652
rect 27068 16643 27120 16652
rect 27068 16609 27077 16643
rect 27077 16609 27111 16643
rect 27111 16609 27120 16643
rect 27068 16600 27120 16609
rect 27436 16643 27488 16652
rect 1492 16396 1544 16448
rect 4068 16396 4120 16448
rect 10048 16396 10100 16448
rect 10784 16396 10836 16448
rect 21456 16464 21508 16516
rect 22560 16464 22612 16516
rect 23572 16464 23624 16516
rect 24492 16532 24544 16584
rect 24676 16532 24728 16584
rect 25044 16532 25096 16584
rect 26608 16532 26660 16584
rect 27436 16609 27445 16643
rect 27445 16609 27479 16643
rect 27479 16609 27488 16643
rect 27436 16600 27488 16609
rect 27620 16600 27672 16652
rect 28172 16600 28224 16652
rect 28356 16600 28408 16652
rect 28816 16643 28868 16652
rect 28816 16609 28825 16643
rect 28825 16609 28859 16643
rect 28859 16609 28868 16643
rect 28816 16600 28868 16609
rect 27160 16464 27212 16516
rect 29092 16600 29144 16652
rect 29368 16643 29420 16652
rect 29368 16609 29377 16643
rect 29377 16609 29411 16643
rect 29411 16609 29420 16643
rect 29368 16600 29420 16609
rect 29736 16532 29788 16584
rect 30380 16643 30432 16652
rect 30380 16609 30389 16643
rect 30389 16609 30423 16643
rect 30423 16609 30432 16643
rect 32220 16668 32272 16720
rect 33692 16736 33744 16788
rect 34980 16779 35032 16788
rect 34980 16745 34989 16779
rect 34989 16745 35023 16779
rect 35023 16745 35032 16779
rect 34980 16736 35032 16745
rect 35992 16736 36044 16788
rect 38844 16736 38896 16788
rect 30380 16600 30432 16609
rect 31116 16600 31168 16652
rect 30472 16532 30524 16584
rect 34060 16668 34112 16720
rect 33232 16600 33284 16652
rect 34612 16600 34664 16652
rect 35624 16643 35676 16652
rect 35624 16609 35633 16643
rect 35633 16609 35667 16643
rect 35667 16609 35676 16643
rect 35624 16600 35676 16609
rect 36268 16643 36320 16652
rect 36268 16609 36277 16643
rect 36277 16609 36311 16643
rect 36311 16609 36320 16643
rect 36268 16600 36320 16609
rect 36544 16643 36596 16652
rect 36544 16609 36553 16643
rect 36553 16609 36587 16643
rect 36587 16609 36596 16643
rect 36544 16600 36596 16609
rect 38568 16643 38620 16652
rect 33508 16532 33560 16584
rect 36084 16532 36136 16584
rect 37556 16532 37608 16584
rect 38568 16609 38577 16643
rect 38577 16609 38611 16643
rect 38611 16609 38620 16643
rect 38568 16600 38620 16609
rect 30012 16464 30064 16516
rect 30840 16507 30892 16516
rect 30840 16473 30849 16507
rect 30849 16473 30883 16507
rect 30883 16473 30892 16507
rect 30840 16464 30892 16473
rect 15568 16396 15620 16448
rect 19340 16396 19392 16448
rect 21180 16396 21232 16448
rect 24216 16396 24268 16448
rect 24676 16396 24728 16448
rect 28172 16439 28224 16448
rect 28172 16405 28181 16439
rect 28181 16405 28215 16439
rect 28215 16405 28224 16439
rect 28172 16396 28224 16405
rect 28908 16396 28960 16448
rect 36636 16464 36688 16516
rect 33508 16396 33560 16448
rect 36360 16396 36412 16448
rect 4246 16294 4298 16346
rect 4310 16294 4362 16346
rect 4374 16294 4426 16346
rect 4438 16294 4490 16346
rect 34966 16294 35018 16346
rect 35030 16294 35082 16346
rect 35094 16294 35146 16346
rect 35158 16294 35210 16346
rect 3148 16192 3200 16244
rect 3976 16192 4028 16244
rect 3424 16056 3476 16108
rect 6276 16192 6328 16244
rect 13728 16192 13780 16244
rect 13084 16124 13136 16176
rect 4804 16056 4856 16108
rect 6552 16056 6604 16108
rect 7840 16056 7892 16108
rect 1492 15988 1544 16040
rect 1676 16031 1728 16040
rect 1676 15997 1685 16031
rect 1685 15997 1719 16031
rect 1719 15997 1728 16031
rect 1676 15988 1728 15997
rect 3700 16031 3752 16040
rect 3700 15997 3709 16031
rect 3709 15997 3743 16031
rect 3743 15997 3752 16031
rect 3700 15988 3752 15997
rect 5172 15988 5224 16040
rect 7012 15988 7064 16040
rect 8668 16031 8720 16040
rect 8668 15997 8677 16031
rect 8677 15997 8711 16031
rect 8711 15997 8720 16031
rect 8668 15988 8720 15997
rect 10784 16056 10836 16108
rect 18328 16099 18380 16108
rect 3792 15852 3844 15904
rect 11520 16031 11572 16040
rect 11520 15997 11529 16031
rect 11529 15997 11563 16031
rect 11563 15997 11572 16031
rect 11520 15988 11572 15997
rect 12900 16031 12952 16040
rect 12900 15997 12909 16031
rect 12909 15997 12943 16031
rect 12943 15997 12952 16031
rect 12900 15988 12952 15997
rect 13084 15988 13136 16040
rect 13544 15988 13596 16040
rect 13820 15988 13872 16040
rect 14832 16031 14884 16040
rect 12532 15920 12584 15972
rect 14832 15997 14841 16031
rect 14841 15997 14875 16031
rect 14875 15997 14884 16031
rect 14832 15988 14884 15997
rect 15476 15988 15528 16040
rect 11612 15895 11664 15904
rect 11612 15861 11621 15895
rect 11621 15861 11655 15895
rect 11655 15861 11664 15895
rect 11612 15852 11664 15861
rect 15936 15895 15988 15904
rect 15936 15861 15945 15895
rect 15945 15861 15979 15895
rect 15979 15861 15988 15895
rect 15936 15852 15988 15861
rect 16672 15852 16724 15904
rect 18328 16065 18337 16099
rect 18337 16065 18371 16099
rect 18371 16065 18380 16099
rect 18328 16056 18380 16065
rect 26516 16192 26568 16244
rect 29000 16192 29052 16244
rect 30196 16192 30248 16244
rect 35532 16192 35584 16244
rect 38200 16192 38252 16244
rect 26424 16167 26476 16176
rect 18696 15988 18748 16040
rect 20720 16031 20772 16040
rect 19892 15920 19944 15972
rect 19432 15895 19484 15904
rect 19432 15861 19441 15895
rect 19441 15861 19475 15895
rect 19475 15861 19484 15895
rect 20720 15997 20729 16031
rect 20729 15997 20763 16031
rect 20763 15997 20772 16031
rect 20720 15988 20772 15997
rect 21272 16056 21324 16108
rect 22100 16031 22152 16040
rect 22100 15997 22109 16031
rect 22109 15997 22143 16031
rect 22143 15997 22152 16031
rect 22100 15988 22152 15997
rect 22284 16031 22336 16040
rect 22284 15997 22293 16031
rect 22293 15997 22327 16031
rect 22327 15997 22336 16031
rect 22284 15988 22336 15997
rect 22652 15988 22704 16040
rect 22928 15988 22980 16040
rect 23480 15988 23532 16040
rect 23848 15988 23900 16040
rect 24124 16031 24176 16040
rect 24124 15997 24133 16031
rect 24133 15997 24167 16031
rect 24167 15997 24176 16031
rect 24124 15988 24176 15997
rect 24400 16031 24452 16040
rect 24400 15997 24409 16031
rect 24409 15997 24443 16031
rect 24443 15997 24452 16031
rect 24400 15988 24452 15997
rect 24492 16031 24544 16040
rect 24492 15997 24501 16031
rect 24501 15997 24535 16031
rect 24535 15997 24544 16031
rect 24676 16031 24728 16040
rect 24492 15988 24544 15997
rect 24676 15997 24685 16031
rect 24685 15997 24719 16031
rect 24719 15997 24728 16031
rect 24676 15988 24728 15997
rect 24952 16031 25004 16040
rect 24952 15997 24961 16031
rect 24961 15997 24995 16031
rect 24995 15997 25004 16031
rect 24952 15988 25004 15997
rect 20812 15920 20864 15972
rect 19432 15852 19484 15861
rect 22100 15852 22152 15904
rect 23020 15852 23072 15904
rect 25136 15920 25188 15972
rect 24400 15852 24452 15904
rect 26424 16133 26433 16167
rect 26433 16133 26467 16167
rect 26467 16133 26476 16167
rect 26424 16124 26476 16133
rect 27344 16099 27396 16108
rect 27344 16065 27353 16099
rect 27353 16065 27387 16099
rect 27387 16065 27396 16099
rect 27344 16056 27396 16065
rect 26148 16031 26200 16040
rect 26148 15997 26157 16031
rect 26157 15997 26191 16031
rect 26191 15997 26200 16031
rect 26148 15988 26200 15997
rect 26332 15988 26384 16040
rect 28356 16056 28408 16108
rect 29276 16056 29328 16108
rect 30472 16099 30524 16108
rect 30472 16065 30481 16099
rect 30481 16065 30515 16099
rect 30515 16065 30524 16099
rect 30472 16056 30524 16065
rect 31116 16056 31168 16108
rect 26056 15920 26108 15972
rect 27804 15988 27856 16040
rect 27252 15920 27304 15972
rect 29184 15988 29236 16040
rect 30288 15988 30340 16040
rect 31024 16031 31076 16040
rect 31024 15997 31033 16031
rect 31033 15997 31067 16031
rect 31067 15997 31076 16031
rect 31024 15988 31076 15997
rect 32220 15988 32272 16040
rect 35624 16124 35676 16176
rect 34336 16056 34388 16108
rect 32956 15988 33008 16040
rect 33692 16031 33744 16040
rect 33692 15997 33701 16031
rect 33701 15997 33735 16031
rect 33735 15997 33744 16031
rect 33692 15988 33744 15997
rect 35440 15988 35492 16040
rect 35808 16031 35860 16040
rect 35808 15997 35817 16031
rect 35817 15997 35851 16031
rect 35851 15997 35860 16031
rect 35808 15988 35860 15997
rect 36084 16056 36136 16108
rect 36360 15988 36412 16040
rect 37188 16056 37240 16108
rect 38752 15988 38804 16040
rect 36544 15920 36596 15972
rect 32036 15852 32088 15904
rect 33784 15852 33836 15904
rect 19606 15750 19658 15802
rect 19670 15750 19722 15802
rect 19734 15750 19786 15802
rect 19798 15750 19850 15802
rect 3700 15648 3752 15700
rect 9680 15648 9732 15700
rect 1676 15580 1728 15632
rect 12624 15648 12676 15700
rect 13636 15648 13688 15700
rect 14464 15648 14516 15700
rect 20812 15648 20864 15700
rect 25228 15648 25280 15700
rect 26608 15691 26660 15700
rect 26608 15657 26617 15691
rect 26617 15657 26651 15691
rect 26651 15657 26660 15691
rect 26608 15648 26660 15657
rect 29276 15691 29328 15700
rect 29276 15657 29285 15691
rect 29285 15657 29319 15691
rect 29319 15657 29328 15691
rect 29276 15648 29328 15657
rect 29644 15648 29696 15700
rect 29920 15648 29972 15700
rect 30012 15648 30064 15700
rect 32312 15648 32364 15700
rect 37832 15691 37884 15700
rect 2780 15512 2832 15564
rect 3884 15555 3936 15564
rect 3884 15521 3893 15555
rect 3893 15521 3927 15555
rect 3927 15521 3936 15555
rect 3884 15512 3936 15521
rect 2688 15444 2740 15496
rect 3792 15444 3844 15496
rect 4068 15487 4120 15496
rect 4068 15453 4077 15487
rect 4077 15453 4111 15487
rect 4111 15453 4120 15487
rect 4068 15444 4120 15453
rect 4804 15444 4856 15496
rect 6920 15444 6972 15496
rect 3516 15376 3568 15428
rect 8484 15512 8536 15564
rect 10416 15555 10468 15564
rect 8852 15444 8904 15496
rect 10416 15521 10425 15555
rect 10425 15521 10459 15555
rect 10459 15521 10468 15555
rect 11612 15580 11664 15632
rect 10416 15512 10468 15521
rect 9772 15444 9824 15496
rect 10508 15487 10560 15496
rect 10508 15453 10517 15487
rect 10517 15453 10551 15487
rect 10551 15453 10560 15487
rect 10508 15444 10560 15453
rect 11060 15555 11112 15564
rect 11060 15521 11069 15555
rect 11069 15521 11103 15555
rect 11103 15521 11112 15555
rect 11060 15512 11112 15521
rect 11704 15555 11756 15564
rect 11704 15521 11713 15555
rect 11713 15521 11747 15555
rect 11747 15521 11756 15555
rect 11704 15512 11756 15521
rect 12808 15580 12860 15632
rect 12532 15512 12584 15564
rect 12992 15555 13044 15564
rect 12992 15521 13001 15555
rect 13001 15521 13035 15555
rect 13035 15521 13044 15555
rect 12992 15512 13044 15521
rect 13084 15512 13136 15564
rect 16396 15555 16448 15564
rect 14464 15444 14516 15496
rect 16396 15521 16405 15555
rect 16405 15521 16439 15555
rect 16439 15521 16448 15555
rect 16396 15512 16448 15521
rect 16488 15512 16540 15564
rect 10232 15376 10284 15428
rect 3240 15308 3292 15360
rect 9036 15308 9088 15360
rect 10140 15308 10192 15360
rect 15292 15308 15344 15360
rect 16672 15444 16724 15496
rect 16948 15308 17000 15360
rect 17592 15580 17644 15632
rect 18512 15580 18564 15632
rect 17960 15555 18012 15564
rect 17960 15521 17969 15555
rect 17969 15521 18003 15555
rect 18003 15521 18012 15555
rect 17960 15512 18012 15521
rect 18696 15555 18748 15564
rect 18696 15521 18705 15555
rect 18705 15521 18739 15555
rect 18739 15521 18748 15555
rect 18696 15512 18748 15521
rect 17684 15487 17736 15496
rect 17684 15453 17693 15487
rect 17693 15453 17727 15487
rect 17727 15453 17736 15487
rect 17684 15444 17736 15453
rect 18144 15444 18196 15496
rect 20536 15512 20588 15564
rect 22192 15580 22244 15632
rect 24400 15580 24452 15632
rect 22100 15555 22152 15564
rect 22100 15521 22109 15555
rect 22109 15521 22143 15555
rect 22143 15521 22152 15555
rect 22284 15555 22336 15564
rect 22100 15512 22152 15521
rect 22284 15521 22293 15555
rect 22293 15521 22327 15555
rect 22327 15521 22336 15555
rect 22284 15512 22336 15521
rect 22560 15555 22612 15564
rect 22560 15521 22569 15555
rect 22569 15521 22603 15555
rect 22603 15521 22612 15555
rect 22560 15512 22612 15521
rect 22652 15555 22704 15564
rect 22652 15521 22661 15555
rect 22661 15521 22695 15555
rect 22695 15521 22704 15555
rect 22652 15512 22704 15521
rect 23296 15512 23348 15564
rect 24124 15555 24176 15564
rect 24124 15521 24133 15555
rect 24133 15521 24167 15555
rect 24167 15521 24176 15555
rect 24124 15512 24176 15521
rect 24952 15555 25004 15564
rect 18972 15487 19024 15496
rect 18972 15453 18981 15487
rect 18981 15453 19015 15487
rect 19015 15453 19024 15487
rect 18972 15444 19024 15453
rect 20812 15444 20864 15496
rect 20720 15376 20772 15428
rect 24032 15444 24084 15496
rect 24400 15444 24452 15496
rect 24952 15521 24961 15555
rect 24961 15521 24995 15555
rect 24995 15521 25004 15555
rect 24952 15512 25004 15521
rect 26884 15512 26936 15564
rect 27160 15555 27212 15564
rect 27160 15521 27169 15555
rect 27169 15521 27203 15555
rect 27203 15521 27212 15555
rect 27160 15512 27212 15521
rect 27896 15555 27948 15564
rect 27896 15521 27905 15555
rect 27905 15521 27939 15555
rect 27939 15521 27948 15555
rect 27896 15512 27948 15521
rect 29368 15580 29420 15632
rect 29736 15580 29788 15632
rect 29828 15555 29880 15564
rect 29828 15521 29837 15555
rect 29837 15521 29871 15555
rect 29871 15521 29880 15555
rect 29828 15512 29880 15521
rect 30196 15555 30248 15564
rect 30196 15521 30205 15555
rect 30205 15521 30239 15555
rect 30239 15521 30248 15555
rect 30196 15512 30248 15521
rect 33508 15580 33560 15632
rect 32956 15512 33008 15564
rect 33140 15512 33192 15564
rect 33784 15555 33836 15564
rect 33784 15521 33793 15555
rect 33793 15521 33827 15555
rect 33827 15521 33836 15555
rect 33784 15512 33836 15521
rect 36268 15580 36320 15632
rect 37832 15657 37841 15691
rect 37841 15657 37875 15691
rect 37875 15657 37884 15691
rect 37832 15648 37884 15657
rect 39028 15691 39080 15700
rect 39028 15657 39037 15691
rect 39037 15657 39071 15691
rect 39071 15657 39080 15691
rect 39028 15648 39080 15657
rect 36176 15555 36228 15564
rect 36176 15521 36185 15555
rect 36185 15521 36219 15555
rect 36219 15521 36228 15555
rect 36176 15512 36228 15521
rect 36452 15555 36504 15564
rect 36452 15521 36461 15555
rect 36461 15521 36495 15555
rect 36495 15521 36504 15555
rect 36452 15512 36504 15521
rect 36544 15512 36596 15564
rect 38936 15555 38988 15564
rect 26148 15444 26200 15496
rect 27988 15487 28040 15496
rect 27988 15453 27997 15487
rect 27997 15453 28031 15487
rect 28031 15453 28040 15487
rect 27988 15444 28040 15453
rect 32128 15444 32180 15496
rect 34244 15444 34296 15496
rect 34428 15444 34480 15496
rect 38936 15521 38945 15555
rect 38945 15521 38979 15555
rect 38979 15521 38988 15555
rect 38936 15512 38988 15521
rect 24676 15376 24728 15428
rect 27436 15419 27488 15428
rect 27436 15385 27445 15419
rect 27445 15385 27479 15419
rect 27479 15385 27488 15419
rect 27436 15376 27488 15385
rect 27804 15376 27856 15428
rect 30932 15376 30984 15428
rect 32036 15376 32088 15428
rect 20536 15308 20588 15360
rect 22928 15308 22980 15360
rect 23388 15308 23440 15360
rect 24492 15308 24544 15360
rect 25688 15351 25740 15360
rect 25688 15317 25697 15351
rect 25697 15317 25731 15351
rect 25731 15317 25740 15351
rect 25688 15308 25740 15317
rect 30564 15308 30616 15360
rect 35348 15308 35400 15360
rect 4246 15206 4298 15258
rect 4310 15206 4362 15258
rect 4374 15206 4426 15258
rect 4438 15206 4490 15258
rect 34966 15206 35018 15258
rect 35030 15206 35082 15258
rect 35094 15206 35146 15258
rect 35158 15206 35210 15258
rect 2780 15147 2832 15156
rect 2780 15113 2789 15147
rect 2789 15113 2823 15147
rect 2823 15113 2832 15147
rect 2780 15104 2832 15113
rect 7012 15104 7064 15156
rect 9220 15104 9272 15156
rect 11060 15104 11112 15156
rect 11796 15104 11848 15156
rect 6920 15036 6972 15088
rect 1492 14900 1544 14952
rect 4068 14943 4120 14952
rect 4068 14909 4077 14943
rect 4077 14909 4111 14943
rect 4111 14909 4120 14943
rect 4068 14900 4120 14909
rect 4620 14900 4672 14952
rect 7104 14764 7156 14816
rect 9496 14968 9548 15020
rect 11704 15036 11756 15088
rect 13360 15079 13412 15088
rect 13360 15045 13369 15079
rect 13369 15045 13403 15079
rect 13403 15045 13412 15079
rect 13360 15036 13412 15045
rect 16028 15104 16080 15156
rect 15660 15036 15712 15088
rect 19432 15104 19484 15156
rect 20444 15104 20496 15156
rect 38752 15147 38804 15156
rect 17224 15036 17276 15088
rect 17868 15036 17920 15088
rect 13820 15011 13872 15020
rect 9036 14943 9088 14952
rect 8116 14764 8168 14816
rect 8208 14764 8260 14816
rect 9036 14909 9045 14943
rect 9045 14909 9079 14943
rect 9079 14909 9088 14943
rect 9036 14900 9088 14909
rect 9220 14943 9272 14952
rect 9220 14909 9229 14943
rect 9229 14909 9263 14943
rect 9263 14909 9272 14943
rect 9220 14900 9272 14909
rect 9588 14943 9640 14952
rect 9588 14909 9597 14943
rect 9597 14909 9631 14943
rect 9631 14909 9640 14943
rect 9588 14900 9640 14909
rect 10600 14900 10652 14952
rect 10784 14943 10836 14952
rect 10784 14909 10793 14943
rect 10793 14909 10827 14943
rect 10827 14909 10836 14943
rect 10784 14900 10836 14909
rect 11428 14900 11480 14952
rect 12624 14900 12676 14952
rect 13820 14977 13829 15011
rect 13829 14977 13863 15011
rect 13863 14977 13872 15011
rect 13820 14968 13872 14977
rect 13636 14943 13688 14952
rect 13636 14909 13645 14943
rect 13645 14909 13679 14943
rect 13679 14909 13688 14943
rect 15292 14968 15344 15020
rect 16396 15011 16448 15020
rect 13636 14900 13688 14909
rect 15384 14900 15436 14952
rect 15568 14900 15620 14952
rect 16396 14977 16405 15011
rect 16405 14977 16439 15011
rect 16439 14977 16448 15011
rect 16396 14968 16448 14977
rect 18512 14968 18564 15020
rect 18972 15011 19024 15020
rect 18972 14977 18981 15011
rect 18981 14977 19015 15011
rect 19015 14977 19024 15011
rect 18972 14968 19024 14977
rect 19340 15036 19392 15088
rect 22744 15036 22796 15088
rect 23020 15036 23072 15088
rect 17960 14900 18012 14952
rect 19340 14943 19392 14952
rect 8944 14832 8996 14884
rect 17684 14832 17736 14884
rect 10416 14764 10468 14816
rect 10968 14807 11020 14816
rect 10968 14773 10977 14807
rect 10977 14773 11011 14807
rect 11011 14773 11020 14807
rect 10968 14764 11020 14773
rect 11704 14807 11756 14816
rect 11704 14773 11713 14807
rect 11713 14773 11747 14807
rect 11747 14773 11756 14807
rect 11704 14764 11756 14773
rect 11796 14764 11848 14816
rect 15108 14764 15160 14816
rect 15384 14764 15436 14816
rect 17960 14764 18012 14816
rect 18420 14764 18472 14816
rect 19340 14909 19349 14943
rect 19349 14909 19383 14943
rect 19383 14909 19392 14943
rect 19340 14900 19392 14909
rect 19984 14943 20036 14952
rect 19984 14909 19993 14943
rect 19993 14909 20027 14943
rect 20027 14909 20036 14943
rect 19984 14900 20036 14909
rect 20720 14943 20772 14952
rect 20720 14909 20729 14943
rect 20729 14909 20763 14943
rect 20763 14909 20772 14943
rect 20720 14900 20772 14909
rect 21180 14943 21232 14952
rect 21180 14909 21189 14943
rect 21189 14909 21223 14943
rect 21223 14909 21232 14943
rect 21180 14900 21232 14909
rect 21456 14900 21508 14952
rect 20904 14832 20956 14884
rect 21272 14832 21324 14884
rect 23112 14900 23164 14952
rect 24952 15036 25004 15088
rect 27896 15036 27948 15088
rect 24492 14900 24544 14952
rect 25596 14943 25648 14952
rect 25596 14909 25605 14943
rect 25605 14909 25639 14943
rect 25639 14909 25648 14943
rect 25596 14900 25648 14909
rect 26424 14900 26476 14952
rect 26608 14943 26660 14952
rect 26608 14909 26617 14943
rect 26617 14909 26651 14943
rect 26651 14909 26660 14943
rect 26608 14900 26660 14909
rect 26884 14900 26936 14952
rect 27528 14900 27580 14952
rect 22560 14875 22612 14884
rect 22560 14841 22569 14875
rect 22569 14841 22603 14875
rect 22603 14841 22612 14875
rect 22560 14832 22612 14841
rect 20812 14764 20864 14816
rect 23664 14764 23716 14816
rect 23940 14807 23992 14816
rect 23940 14773 23949 14807
rect 23949 14773 23983 14807
rect 23983 14773 23992 14807
rect 23940 14764 23992 14773
rect 24124 14832 24176 14884
rect 28172 14900 28224 14952
rect 38752 15113 38761 15147
rect 38761 15113 38795 15147
rect 38795 15113 38804 15147
rect 38752 15104 38804 15113
rect 33140 15079 33192 15088
rect 33140 15045 33149 15079
rect 33149 15045 33183 15079
rect 33183 15045 33192 15079
rect 33140 15036 33192 15045
rect 29552 14968 29604 15020
rect 36176 15011 36228 15020
rect 29736 14943 29788 14952
rect 29736 14909 29745 14943
rect 29745 14909 29779 14943
rect 29779 14909 29788 14943
rect 29736 14900 29788 14909
rect 29828 14900 29880 14952
rect 30288 14943 30340 14952
rect 30288 14909 30297 14943
rect 30297 14909 30331 14943
rect 30331 14909 30340 14943
rect 30288 14900 30340 14909
rect 31484 14900 31536 14952
rect 36176 14977 36185 15011
rect 36185 14977 36219 15011
rect 36219 14977 36228 15011
rect 36176 14968 36228 14977
rect 36636 14968 36688 15020
rect 33140 14943 33192 14952
rect 33140 14909 33149 14943
rect 33149 14909 33183 14943
rect 33183 14909 33192 14943
rect 33140 14900 33192 14909
rect 34428 14900 34480 14952
rect 35256 14943 35308 14952
rect 35256 14909 35265 14943
rect 35265 14909 35299 14943
rect 35299 14909 35308 14943
rect 35256 14900 35308 14909
rect 35716 14943 35768 14952
rect 35716 14909 35725 14943
rect 35725 14909 35759 14943
rect 35759 14909 35768 14943
rect 35716 14900 35768 14909
rect 36360 14900 36412 14952
rect 25412 14764 25464 14816
rect 26056 14764 26108 14816
rect 28724 14832 28776 14884
rect 30288 14764 30340 14816
rect 30564 14832 30616 14884
rect 31116 14832 31168 14884
rect 31392 14875 31444 14884
rect 31392 14841 31401 14875
rect 31401 14841 31435 14875
rect 31435 14841 31444 14875
rect 31392 14832 31444 14841
rect 32220 14832 32272 14884
rect 33968 14832 34020 14884
rect 36544 14900 36596 14952
rect 37740 14943 37792 14952
rect 37740 14909 37749 14943
rect 37749 14909 37783 14943
rect 37783 14909 37792 14943
rect 37740 14900 37792 14909
rect 38568 14943 38620 14952
rect 38568 14909 38577 14943
rect 38577 14909 38611 14943
rect 38611 14909 38620 14943
rect 38568 14900 38620 14909
rect 34336 14764 34388 14816
rect 37832 14764 37884 14816
rect 19606 14662 19658 14714
rect 19670 14662 19722 14714
rect 19734 14662 19786 14714
rect 19798 14662 19850 14714
rect 1860 14560 1912 14612
rect 3976 14560 4028 14612
rect 4804 14535 4856 14544
rect 4804 14501 4813 14535
rect 4813 14501 4847 14535
rect 4847 14501 4856 14535
rect 4804 14492 4856 14501
rect 8116 14492 8168 14544
rect 1952 14424 2004 14476
rect 2504 14467 2556 14476
rect 2504 14433 2513 14467
rect 2513 14433 2547 14467
rect 2547 14433 2556 14467
rect 2504 14424 2556 14433
rect 3240 14467 3292 14476
rect 3240 14433 3249 14467
rect 3249 14433 3283 14467
rect 3283 14433 3292 14467
rect 3240 14424 3292 14433
rect 4068 14356 4120 14408
rect 5448 14424 5500 14476
rect 10324 14492 10376 14544
rect 11520 14560 11572 14612
rect 11888 14560 11940 14612
rect 15660 14560 15712 14612
rect 15844 14560 15896 14612
rect 18512 14560 18564 14612
rect 13360 14492 13412 14544
rect 18880 14492 18932 14544
rect 22008 14560 22060 14612
rect 23664 14560 23716 14612
rect 24216 14560 24268 14612
rect 26608 14603 26660 14612
rect 26608 14569 26617 14603
rect 26617 14569 26651 14603
rect 26651 14569 26660 14603
rect 26608 14560 26660 14569
rect 28816 14560 28868 14612
rect 30564 14603 30616 14612
rect 30564 14569 30573 14603
rect 30573 14569 30607 14603
rect 30607 14569 30616 14603
rect 30564 14560 30616 14569
rect 38568 14560 38620 14612
rect 23388 14492 23440 14544
rect 26424 14492 26476 14544
rect 30748 14492 30800 14544
rect 32864 14492 32916 14544
rect 33324 14492 33376 14544
rect 34336 14492 34388 14544
rect 9036 14424 9088 14476
rect 10232 14467 10284 14476
rect 10232 14433 10241 14467
rect 10241 14433 10275 14467
rect 10275 14433 10284 14467
rect 10232 14424 10284 14433
rect 10508 14467 10560 14476
rect 10508 14433 10517 14467
rect 10517 14433 10551 14467
rect 10551 14433 10560 14467
rect 10508 14424 10560 14433
rect 10600 14424 10652 14476
rect 5080 14356 5132 14408
rect 6184 14399 6236 14408
rect 3424 14263 3476 14272
rect 3424 14229 3433 14263
rect 3433 14229 3467 14263
rect 3467 14229 3476 14263
rect 3424 14220 3476 14229
rect 6184 14365 6193 14399
rect 6193 14365 6227 14399
rect 6227 14365 6236 14399
rect 6184 14356 6236 14365
rect 8668 14399 8720 14408
rect 8668 14365 8677 14399
rect 8677 14365 8711 14399
rect 8711 14365 8720 14399
rect 8668 14356 8720 14365
rect 13544 14424 13596 14476
rect 13820 14467 13872 14476
rect 13820 14433 13829 14467
rect 13829 14433 13863 14467
rect 13863 14433 13872 14467
rect 13820 14424 13872 14433
rect 14464 14467 14516 14476
rect 14464 14433 14473 14467
rect 14473 14433 14507 14467
rect 14507 14433 14516 14467
rect 14464 14424 14516 14433
rect 16488 14424 16540 14476
rect 9956 14288 10008 14340
rect 12532 14288 12584 14340
rect 12992 14288 13044 14340
rect 13268 14288 13320 14340
rect 18052 14399 18104 14408
rect 18052 14365 18061 14399
rect 18061 14365 18095 14399
rect 18095 14365 18104 14399
rect 18052 14356 18104 14365
rect 19708 14424 19760 14476
rect 23020 14467 23072 14476
rect 23020 14433 23029 14467
rect 23029 14433 23063 14467
rect 23063 14433 23072 14467
rect 23020 14424 23072 14433
rect 23112 14424 23164 14476
rect 18696 14356 18748 14408
rect 21180 14399 21232 14408
rect 21180 14365 21189 14399
rect 21189 14365 21223 14399
rect 21223 14365 21232 14399
rect 21180 14356 21232 14365
rect 22744 14356 22796 14408
rect 24952 14424 25004 14476
rect 24492 14399 24544 14408
rect 24492 14365 24501 14399
rect 24501 14365 24535 14399
rect 24535 14365 24544 14399
rect 24492 14356 24544 14365
rect 25504 14424 25556 14476
rect 26700 14467 26752 14476
rect 26700 14433 26709 14467
rect 26709 14433 26743 14467
rect 26743 14433 26752 14467
rect 26700 14424 26752 14433
rect 7564 14220 7616 14272
rect 15200 14220 15252 14272
rect 20168 14288 20220 14340
rect 25596 14288 25648 14340
rect 25964 14356 26016 14408
rect 27896 14424 27948 14476
rect 29276 14467 29328 14476
rect 29276 14433 29285 14467
rect 29285 14433 29319 14467
rect 29319 14433 29328 14467
rect 29276 14424 29328 14433
rect 29828 14467 29880 14476
rect 29828 14433 29837 14467
rect 29837 14433 29871 14467
rect 29871 14433 29880 14467
rect 29828 14424 29880 14433
rect 29920 14424 29972 14476
rect 32588 14467 32640 14476
rect 27620 14356 27672 14408
rect 28448 14356 28500 14408
rect 29736 14356 29788 14408
rect 30196 14356 30248 14408
rect 32588 14433 32597 14467
rect 32597 14433 32631 14467
rect 32631 14433 32640 14467
rect 32588 14424 32640 14433
rect 33968 14424 34020 14476
rect 33232 14356 33284 14408
rect 33600 14399 33652 14408
rect 33600 14365 33609 14399
rect 33609 14365 33643 14399
rect 33643 14365 33652 14399
rect 33600 14356 33652 14365
rect 27068 14288 27120 14340
rect 33692 14288 33744 14340
rect 19432 14220 19484 14272
rect 21364 14220 21416 14272
rect 23296 14220 23348 14272
rect 23572 14220 23624 14272
rect 29276 14220 29328 14272
rect 34612 14467 34664 14476
rect 34612 14433 34621 14467
rect 34621 14433 34655 14467
rect 34655 14433 34664 14467
rect 34612 14424 34664 14433
rect 34796 14424 34848 14476
rect 36176 14424 36228 14476
rect 37740 14492 37792 14544
rect 38660 14492 38712 14544
rect 37924 14467 37976 14476
rect 37924 14433 37933 14467
rect 37933 14433 37967 14467
rect 37967 14433 37976 14467
rect 37924 14424 37976 14433
rect 38016 14467 38068 14476
rect 38016 14433 38025 14467
rect 38025 14433 38059 14467
rect 38059 14433 38068 14467
rect 38936 14467 38988 14476
rect 38016 14424 38068 14433
rect 38936 14433 38945 14467
rect 38945 14433 38979 14467
rect 38979 14433 38988 14467
rect 38936 14424 38988 14433
rect 34336 14356 34388 14408
rect 36912 14356 36964 14408
rect 37740 14399 37792 14408
rect 37740 14365 37749 14399
rect 37749 14365 37783 14399
rect 37783 14365 37792 14399
rect 37740 14356 37792 14365
rect 35440 14220 35492 14272
rect 35532 14220 35584 14272
rect 4246 14118 4298 14170
rect 4310 14118 4362 14170
rect 4374 14118 4426 14170
rect 4438 14118 4490 14170
rect 34966 14118 35018 14170
rect 35030 14118 35082 14170
rect 35094 14118 35146 14170
rect 35158 14118 35210 14170
rect 3884 13948 3936 14000
rect 1492 13880 1544 13932
rect 1860 13923 1912 13932
rect 1860 13889 1869 13923
rect 1869 13889 1903 13923
rect 1903 13889 1912 13923
rect 1860 13880 1912 13889
rect 4620 13923 4672 13932
rect 4620 13889 4629 13923
rect 4629 13889 4663 13923
rect 4663 13889 4672 13923
rect 4620 13880 4672 13889
rect 3976 13855 4028 13864
rect 3976 13821 3985 13855
rect 3985 13821 4019 13855
rect 4019 13821 4028 13855
rect 3976 13812 4028 13821
rect 4160 13855 4212 13864
rect 4160 13821 4169 13855
rect 4169 13821 4203 13855
rect 4203 13821 4212 13855
rect 4160 13812 4212 13821
rect 6184 13948 6236 14000
rect 8944 14016 8996 14068
rect 9312 14016 9364 14068
rect 11428 14016 11480 14068
rect 13820 14016 13872 14068
rect 19248 14016 19300 14068
rect 20904 14016 20956 14068
rect 24860 14016 24912 14068
rect 27528 14016 27580 14068
rect 12440 13948 12492 14000
rect 16488 13991 16540 14000
rect 16488 13957 16497 13991
rect 16497 13957 16531 13991
rect 16531 13957 16540 13991
rect 16488 13948 16540 13957
rect 5264 13923 5316 13932
rect 5264 13889 5273 13923
rect 5273 13889 5307 13923
rect 5307 13889 5316 13923
rect 5264 13880 5316 13889
rect 10048 13880 10100 13932
rect 15568 13880 15620 13932
rect 17960 13948 18012 14000
rect 18052 13948 18104 14000
rect 19616 13948 19668 14000
rect 19984 13948 20036 14000
rect 30380 14016 30432 14068
rect 31484 14016 31536 14068
rect 34336 14016 34388 14068
rect 35532 14016 35584 14068
rect 5356 13855 5408 13864
rect 5356 13821 5365 13855
rect 5365 13821 5399 13855
rect 5399 13821 5408 13855
rect 5356 13812 5408 13821
rect 5816 13855 5868 13864
rect 5816 13821 5825 13855
rect 5825 13821 5859 13855
rect 5859 13821 5868 13855
rect 5816 13812 5868 13821
rect 7380 13855 7432 13864
rect 2964 13719 3016 13728
rect 2964 13685 2973 13719
rect 2973 13685 3007 13719
rect 3007 13685 3016 13719
rect 2964 13676 3016 13685
rect 7380 13821 7389 13855
rect 7389 13821 7423 13855
rect 7423 13821 7432 13855
rect 7380 13812 7432 13821
rect 7564 13855 7616 13864
rect 7564 13821 7573 13855
rect 7573 13821 7607 13855
rect 7607 13821 7616 13855
rect 7564 13812 7616 13821
rect 8208 13855 8260 13864
rect 8208 13821 8217 13855
rect 8217 13821 8251 13855
rect 8251 13821 8260 13855
rect 8208 13812 8260 13821
rect 7656 13744 7708 13796
rect 9220 13855 9272 13864
rect 9220 13821 9229 13855
rect 9229 13821 9263 13855
rect 9263 13821 9272 13855
rect 9220 13812 9272 13821
rect 9588 13855 9640 13864
rect 9588 13821 9597 13855
rect 9597 13821 9631 13855
rect 9631 13821 9640 13855
rect 9588 13812 9640 13821
rect 10140 13855 10192 13864
rect 10140 13821 10149 13855
rect 10149 13821 10183 13855
rect 10183 13821 10192 13855
rect 10140 13812 10192 13821
rect 11520 13855 11572 13864
rect 9864 13744 9916 13796
rect 10968 13744 11020 13796
rect 11520 13821 11529 13855
rect 11529 13821 11563 13855
rect 11563 13821 11572 13855
rect 11520 13812 11572 13821
rect 11888 13855 11940 13864
rect 11888 13821 11897 13855
rect 11897 13821 11931 13855
rect 11931 13821 11940 13855
rect 11888 13812 11940 13821
rect 12532 13855 12584 13864
rect 12532 13821 12541 13855
rect 12541 13821 12575 13855
rect 12575 13821 12584 13855
rect 12532 13812 12584 13821
rect 13268 13812 13320 13864
rect 13636 13812 13688 13864
rect 15292 13855 15344 13864
rect 15292 13821 15301 13855
rect 15301 13821 15335 13855
rect 15335 13821 15344 13855
rect 15292 13812 15344 13821
rect 21180 13923 21232 13932
rect 16672 13812 16724 13864
rect 17684 13812 17736 13864
rect 18420 13855 18472 13864
rect 16764 13744 16816 13796
rect 18420 13821 18429 13855
rect 18429 13821 18463 13855
rect 18463 13821 18472 13855
rect 18420 13812 18472 13821
rect 18880 13812 18932 13864
rect 8300 13676 8352 13728
rect 9588 13676 9640 13728
rect 14740 13676 14792 13728
rect 21180 13889 21189 13923
rect 21189 13889 21223 13923
rect 21223 13889 21232 13923
rect 21180 13880 21232 13889
rect 19248 13855 19300 13864
rect 19248 13821 19257 13855
rect 19257 13821 19291 13855
rect 19291 13821 19300 13855
rect 19248 13812 19300 13821
rect 19616 13855 19668 13864
rect 19616 13821 19625 13855
rect 19625 13821 19659 13855
rect 19659 13821 19668 13855
rect 19616 13812 19668 13821
rect 20168 13812 20220 13864
rect 20812 13855 20864 13864
rect 20812 13821 20821 13855
rect 20821 13821 20855 13855
rect 20855 13821 20864 13855
rect 20812 13812 20864 13821
rect 21272 13855 21324 13864
rect 21272 13821 21281 13855
rect 21281 13821 21315 13855
rect 21315 13821 21324 13855
rect 21272 13812 21324 13821
rect 22560 13880 22612 13932
rect 26056 13923 26108 13932
rect 26056 13889 26065 13923
rect 26065 13889 26099 13923
rect 26099 13889 26108 13923
rect 26056 13880 26108 13889
rect 26148 13880 26200 13932
rect 29828 13923 29880 13932
rect 29828 13889 29837 13923
rect 29837 13889 29871 13923
rect 29871 13889 29880 13923
rect 29828 13880 29880 13889
rect 19156 13744 19208 13796
rect 19984 13676 20036 13728
rect 20904 13744 20956 13796
rect 22192 13812 22244 13864
rect 23664 13855 23716 13864
rect 23664 13821 23673 13855
rect 23673 13821 23707 13855
rect 23707 13821 23716 13855
rect 23664 13812 23716 13821
rect 25596 13812 25648 13864
rect 28448 13855 28500 13864
rect 28448 13821 28457 13855
rect 28457 13821 28491 13855
rect 28491 13821 28500 13855
rect 28448 13812 28500 13821
rect 29644 13855 29696 13864
rect 29644 13821 29653 13855
rect 29653 13821 29687 13855
rect 29687 13821 29696 13855
rect 29644 13812 29696 13821
rect 29736 13812 29788 13864
rect 30564 13855 30616 13864
rect 21456 13676 21508 13728
rect 22468 13744 22520 13796
rect 30564 13821 30573 13855
rect 30573 13821 30607 13855
rect 30607 13821 30616 13855
rect 30564 13812 30616 13821
rect 31116 13948 31168 14000
rect 32588 13948 32640 14000
rect 33140 13923 33192 13932
rect 33140 13889 33149 13923
rect 33149 13889 33183 13923
rect 33183 13889 33192 13923
rect 33140 13880 33192 13889
rect 31392 13855 31444 13864
rect 31392 13821 31401 13855
rect 31401 13821 31435 13855
rect 31435 13821 31444 13855
rect 31392 13812 31444 13821
rect 31944 13812 31996 13864
rect 32496 13855 32548 13864
rect 32496 13821 32505 13855
rect 32505 13821 32539 13855
rect 32539 13821 32548 13855
rect 32496 13812 32548 13821
rect 33324 13812 33376 13864
rect 33508 13855 33560 13864
rect 33508 13821 33517 13855
rect 33517 13821 33551 13855
rect 33551 13821 33560 13855
rect 33508 13812 33560 13821
rect 35440 13923 35492 13932
rect 35440 13889 35449 13923
rect 35449 13889 35483 13923
rect 35483 13889 35492 13923
rect 35440 13880 35492 13889
rect 33876 13812 33928 13864
rect 35624 13855 35676 13864
rect 35624 13821 35633 13855
rect 35633 13821 35667 13855
rect 35667 13821 35676 13855
rect 37832 14016 37884 14068
rect 38108 13948 38160 14000
rect 38568 13880 38620 13932
rect 35624 13812 35676 13821
rect 36084 13812 36136 13864
rect 37372 13855 37424 13864
rect 37372 13821 37381 13855
rect 37381 13821 37415 13855
rect 37415 13821 37424 13855
rect 37372 13812 37424 13821
rect 37556 13855 37608 13864
rect 37556 13821 37565 13855
rect 37565 13821 37599 13855
rect 37599 13821 37608 13855
rect 37556 13812 37608 13821
rect 37832 13812 37884 13864
rect 34796 13744 34848 13796
rect 36544 13744 36596 13796
rect 37280 13744 37332 13796
rect 37740 13744 37792 13796
rect 22192 13676 22244 13728
rect 24768 13676 24820 13728
rect 27528 13676 27580 13728
rect 32956 13676 33008 13728
rect 33140 13676 33192 13728
rect 33784 13676 33836 13728
rect 34336 13676 34388 13728
rect 34612 13676 34664 13728
rect 19606 13574 19658 13626
rect 19670 13574 19722 13626
rect 19734 13574 19786 13626
rect 19798 13574 19850 13626
rect 1676 13472 1728 13524
rect 2964 13404 3016 13456
rect 5080 13404 5132 13456
rect 11244 13404 11296 13456
rect 15844 13472 15896 13524
rect 16856 13472 16908 13524
rect 18236 13515 18288 13524
rect 18236 13481 18245 13515
rect 18245 13481 18279 13515
rect 18279 13481 18288 13515
rect 18236 13472 18288 13481
rect 18328 13472 18380 13524
rect 19156 13472 19208 13524
rect 21272 13472 21324 13524
rect 23756 13472 23808 13524
rect 2780 13379 2832 13388
rect 2780 13345 2789 13379
rect 2789 13345 2823 13379
rect 2823 13345 2832 13379
rect 2780 13336 2832 13345
rect 3332 13336 3384 13388
rect 4804 13336 4856 13388
rect 7104 13379 7156 13388
rect 7104 13345 7113 13379
rect 7113 13345 7147 13379
rect 7147 13345 7156 13379
rect 7104 13336 7156 13345
rect 7196 13336 7248 13388
rect 7656 13379 7708 13388
rect 7656 13345 7665 13379
rect 7665 13345 7699 13379
rect 7699 13345 7708 13379
rect 7656 13336 7708 13345
rect 8300 13379 8352 13388
rect 8300 13345 8309 13379
rect 8309 13345 8343 13379
rect 8343 13345 8352 13379
rect 8300 13336 8352 13345
rect 8852 13379 8904 13388
rect 8852 13345 8861 13379
rect 8861 13345 8895 13379
rect 8895 13345 8904 13379
rect 8852 13336 8904 13345
rect 9864 13379 9916 13388
rect 9864 13345 9873 13379
rect 9873 13345 9907 13379
rect 9907 13345 9916 13379
rect 9864 13336 9916 13345
rect 10048 13336 10100 13388
rect 11520 13379 11572 13388
rect 11520 13345 11529 13379
rect 11529 13345 11563 13379
rect 11563 13345 11572 13379
rect 11520 13336 11572 13345
rect 12532 13404 12584 13456
rect 11980 13379 12032 13388
rect 11980 13345 11989 13379
rect 11989 13345 12023 13379
rect 12023 13345 12032 13379
rect 11980 13336 12032 13345
rect 2688 13311 2740 13320
rect 2688 13277 2697 13311
rect 2697 13277 2731 13311
rect 2731 13277 2740 13311
rect 2688 13268 2740 13277
rect 3424 13200 3476 13252
rect 5172 13268 5224 13320
rect 9312 13268 9364 13320
rect 10968 13268 11020 13320
rect 13636 13379 13688 13388
rect 13636 13345 13645 13379
rect 13645 13345 13679 13379
rect 13679 13345 13688 13379
rect 13636 13336 13688 13345
rect 13728 13336 13780 13388
rect 15292 13379 15344 13388
rect 15292 13345 15301 13379
rect 15301 13345 15335 13379
rect 15335 13345 15344 13379
rect 15292 13336 15344 13345
rect 15936 13336 15988 13388
rect 16764 13379 16816 13388
rect 12256 13311 12308 13320
rect 12256 13277 12265 13311
rect 12265 13277 12299 13311
rect 12299 13277 12308 13311
rect 12256 13268 12308 13277
rect 9220 13200 9272 13252
rect 15476 13243 15528 13252
rect 15476 13209 15485 13243
rect 15485 13209 15519 13243
rect 15519 13209 15528 13243
rect 15476 13200 15528 13209
rect 1952 13175 2004 13184
rect 1952 13141 1961 13175
rect 1961 13141 1995 13175
rect 1995 13141 2004 13175
rect 1952 13132 2004 13141
rect 6828 13132 6880 13184
rect 7656 13132 7708 13184
rect 9680 13132 9732 13184
rect 10968 13132 11020 13184
rect 13636 13132 13688 13184
rect 14556 13132 14608 13184
rect 15016 13132 15068 13184
rect 16764 13345 16773 13379
rect 16773 13345 16807 13379
rect 16807 13345 16816 13379
rect 16764 13336 16816 13345
rect 17132 13379 17184 13388
rect 17132 13345 17141 13379
rect 17141 13345 17175 13379
rect 17175 13345 17184 13379
rect 17132 13336 17184 13345
rect 17868 13336 17920 13388
rect 18236 13336 18288 13388
rect 21364 13379 21416 13388
rect 21364 13345 21373 13379
rect 21373 13345 21407 13379
rect 21407 13345 21416 13379
rect 21364 13336 21416 13345
rect 21456 13336 21508 13388
rect 22560 13379 22612 13388
rect 22560 13345 22569 13379
rect 22569 13345 22603 13379
rect 22603 13345 22612 13379
rect 22560 13336 22612 13345
rect 24768 13404 24820 13456
rect 28448 13472 28500 13524
rect 33692 13515 33744 13524
rect 24952 13404 25004 13456
rect 18328 13268 18380 13320
rect 19432 13268 19484 13320
rect 23940 13268 23992 13320
rect 20536 13200 20588 13252
rect 26240 13336 26292 13388
rect 27436 13379 27488 13388
rect 27436 13345 27445 13379
rect 27445 13345 27479 13379
rect 27479 13345 27488 13379
rect 27436 13336 27488 13345
rect 26608 13268 26660 13320
rect 29092 13336 29144 13388
rect 29644 13379 29696 13388
rect 29644 13345 29653 13379
rect 29653 13345 29687 13379
rect 29687 13345 29696 13379
rect 29644 13336 29696 13345
rect 30840 13404 30892 13456
rect 32128 13404 32180 13456
rect 29736 13268 29788 13320
rect 30196 13268 30248 13320
rect 30288 13268 30340 13320
rect 31116 13336 31168 13388
rect 32128 13268 32180 13320
rect 33692 13481 33701 13515
rect 33701 13481 33735 13515
rect 33735 13481 33744 13515
rect 33692 13472 33744 13481
rect 33876 13472 33928 13524
rect 34612 13472 34664 13524
rect 36176 13472 36228 13524
rect 32864 13404 32916 13456
rect 32956 13336 33008 13388
rect 33508 13404 33560 13456
rect 33968 13404 34020 13456
rect 33784 13336 33836 13388
rect 34888 13336 34940 13388
rect 35440 13379 35492 13388
rect 35440 13345 35449 13379
rect 35449 13345 35483 13379
rect 35483 13345 35492 13379
rect 35440 13336 35492 13345
rect 37372 13472 37424 13524
rect 36544 13404 36596 13456
rect 21548 13132 21600 13184
rect 22008 13132 22060 13184
rect 28080 13132 28132 13184
rect 30472 13132 30524 13184
rect 32956 13243 33008 13252
rect 32956 13209 32965 13243
rect 32965 13209 32999 13243
rect 32999 13209 33008 13243
rect 32956 13200 33008 13209
rect 34612 13268 34664 13320
rect 35256 13268 35308 13320
rect 36176 13268 36228 13320
rect 37556 13404 37608 13456
rect 37372 13336 37424 13388
rect 38108 13379 38160 13388
rect 38108 13345 38117 13379
rect 38117 13345 38151 13379
rect 38151 13345 38160 13379
rect 38108 13336 38160 13345
rect 38568 13379 38620 13388
rect 38568 13345 38577 13379
rect 38577 13345 38611 13379
rect 38611 13345 38620 13379
rect 38568 13336 38620 13345
rect 37188 13311 37240 13320
rect 37188 13277 37197 13311
rect 37197 13277 37231 13311
rect 37231 13277 37240 13311
rect 37188 13268 37240 13277
rect 36084 13200 36136 13252
rect 38476 13200 38528 13252
rect 35624 13132 35676 13184
rect 4246 13030 4298 13082
rect 4310 13030 4362 13082
rect 4374 13030 4426 13082
rect 4438 13030 4490 13082
rect 34966 13030 35018 13082
rect 35030 13030 35082 13082
rect 35094 13030 35146 13082
rect 35158 13030 35210 13082
rect 2780 12971 2832 12980
rect 2780 12937 2789 12971
rect 2789 12937 2823 12971
rect 2823 12937 2832 12971
rect 2780 12928 2832 12937
rect 5356 12928 5408 12980
rect 8300 12860 8352 12912
rect 9312 12860 9364 12912
rect 1676 12835 1728 12844
rect 1676 12801 1685 12835
rect 1685 12801 1719 12835
rect 1719 12801 1728 12835
rect 1676 12792 1728 12801
rect 2872 12792 2924 12844
rect 5264 12792 5316 12844
rect 9588 12792 9640 12844
rect 3516 12767 3568 12776
rect 3516 12733 3525 12767
rect 3525 12733 3559 12767
rect 3559 12733 3568 12767
rect 3516 12724 3568 12733
rect 3792 12767 3844 12776
rect 3792 12733 3801 12767
rect 3801 12733 3835 12767
rect 3835 12733 3844 12767
rect 3792 12724 3844 12733
rect 5724 12767 5776 12776
rect 5724 12733 5733 12767
rect 5733 12733 5767 12767
rect 5767 12733 5776 12767
rect 6828 12767 6880 12776
rect 5724 12724 5776 12733
rect 6828 12733 6837 12767
rect 6837 12733 6871 12767
rect 6871 12733 6880 12767
rect 6828 12724 6880 12733
rect 7656 12767 7708 12776
rect 7656 12733 7665 12767
rect 7665 12733 7699 12767
rect 7699 12733 7708 12767
rect 7656 12724 7708 12733
rect 7932 12767 7984 12776
rect 7932 12733 7941 12767
rect 7941 12733 7975 12767
rect 7975 12733 7984 12767
rect 7932 12724 7984 12733
rect 8208 12767 8260 12776
rect 8208 12733 8217 12767
rect 8217 12733 8251 12767
rect 8251 12733 8260 12767
rect 8208 12724 8260 12733
rect 8392 12724 8444 12776
rect 9220 12724 9272 12776
rect 10968 12767 11020 12776
rect 10968 12733 10977 12767
rect 10977 12733 11011 12767
rect 11011 12733 11020 12767
rect 10968 12724 11020 12733
rect 11244 12767 11296 12776
rect 11244 12733 11253 12767
rect 11253 12733 11287 12767
rect 11287 12733 11296 12767
rect 11244 12724 11296 12733
rect 11428 12767 11480 12776
rect 11428 12733 11437 12767
rect 11437 12733 11471 12767
rect 11471 12733 11480 12767
rect 11428 12724 11480 12733
rect 12348 12724 12400 12776
rect 12532 12724 12584 12776
rect 12900 12767 12952 12776
rect 12900 12733 12909 12767
rect 12909 12733 12943 12767
rect 12943 12733 12952 12767
rect 12900 12724 12952 12733
rect 15200 12792 15252 12844
rect 15844 12928 15896 12980
rect 18328 12971 18380 12980
rect 18328 12937 18337 12971
rect 18337 12937 18371 12971
rect 18371 12937 18380 12971
rect 18328 12928 18380 12937
rect 19340 12928 19392 12980
rect 19984 12928 20036 12980
rect 20720 12928 20772 12980
rect 26056 12928 26108 12980
rect 30196 12928 30248 12980
rect 31392 12928 31444 12980
rect 32128 12928 32180 12980
rect 33784 12928 33836 12980
rect 36360 12971 36412 12980
rect 36360 12937 36369 12971
rect 36369 12937 36403 12971
rect 36403 12937 36412 12971
rect 36360 12928 36412 12937
rect 36912 12928 36964 12980
rect 16212 12860 16264 12912
rect 17316 12792 17368 12844
rect 19064 12792 19116 12844
rect 14740 12767 14792 12776
rect 14740 12733 14749 12767
rect 14749 12733 14783 12767
rect 14783 12733 14792 12767
rect 14740 12724 14792 12733
rect 15108 12767 15160 12776
rect 15108 12733 15117 12767
rect 15117 12733 15151 12767
rect 15151 12733 15160 12767
rect 15108 12724 15160 12733
rect 16212 12767 16264 12776
rect 16212 12733 16221 12767
rect 16221 12733 16255 12767
rect 16255 12733 16264 12767
rect 16212 12724 16264 12733
rect 18880 12767 18932 12776
rect 16764 12656 16816 12708
rect 14004 12588 14056 12640
rect 18880 12733 18889 12767
rect 18889 12733 18923 12767
rect 18923 12733 18932 12767
rect 18880 12724 18932 12733
rect 19432 12724 19484 12776
rect 19984 12767 20036 12776
rect 19984 12733 19993 12767
rect 19993 12733 20027 12767
rect 20027 12733 20036 12767
rect 19984 12724 20036 12733
rect 19892 12656 19944 12708
rect 19432 12588 19484 12640
rect 25504 12860 25556 12912
rect 25872 12903 25924 12912
rect 25872 12869 25881 12903
rect 25881 12869 25915 12903
rect 25915 12869 25924 12903
rect 25872 12860 25924 12869
rect 27988 12860 28040 12912
rect 30748 12860 30800 12912
rect 33968 12860 34020 12912
rect 23940 12835 23992 12844
rect 21272 12767 21324 12776
rect 21272 12733 21281 12767
rect 21281 12733 21315 12767
rect 21315 12733 21324 12767
rect 21272 12724 21324 12733
rect 21548 12767 21600 12776
rect 21548 12733 21557 12767
rect 21557 12733 21591 12767
rect 21591 12733 21600 12767
rect 21548 12724 21600 12733
rect 23296 12656 23348 12708
rect 22652 12631 22704 12640
rect 22652 12597 22661 12631
rect 22661 12597 22695 12631
rect 22695 12597 22704 12631
rect 22652 12588 22704 12597
rect 23388 12588 23440 12640
rect 23940 12801 23949 12835
rect 23949 12801 23983 12835
rect 23983 12801 23992 12835
rect 23940 12792 23992 12801
rect 27620 12792 27672 12844
rect 30288 12792 30340 12844
rect 30840 12835 30892 12844
rect 30840 12801 30849 12835
rect 30849 12801 30883 12835
rect 30883 12801 30892 12835
rect 30840 12792 30892 12801
rect 33324 12792 33376 12844
rect 33508 12792 33560 12844
rect 23664 12767 23716 12776
rect 23664 12733 23673 12767
rect 23673 12733 23707 12767
rect 23707 12733 23716 12767
rect 23664 12724 23716 12733
rect 24216 12724 24268 12776
rect 25872 12724 25924 12776
rect 26516 12724 26568 12776
rect 26700 12724 26752 12776
rect 28448 12724 28500 12776
rect 28632 12656 28684 12708
rect 29920 12724 29972 12776
rect 31116 12767 31168 12776
rect 31116 12733 31125 12767
rect 31125 12733 31159 12767
rect 31159 12733 31168 12767
rect 31116 12724 31168 12733
rect 31392 12724 31444 12776
rect 32220 12767 32272 12776
rect 32220 12733 32229 12767
rect 32229 12733 32263 12767
rect 32263 12733 32272 12767
rect 32220 12724 32272 12733
rect 33140 12767 33192 12776
rect 33140 12733 33149 12767
rect 33149 12733 33183 12767
rect 33183 12733 33192 12767
rect 33140 12724 33192 12733
rect 34520 12792 34572 12844
rect 34796 12792 34848 12844
rect 35256 12767 35308 12776
rect 31668 12656 31720 12708
rect 24032 12588 24084 12640
rect 25044 12631 25096 12640
rect 25044 12597 25053 12631
rect 25053 12597 25087 12631
rect 25087 12597 25096 12631
rect 25044 12588 25096 12597
rect 25320 12588 25372 12640
rect 27528 12588 27580 12640
rect 30564 12588 30616 12640
rect 32128 12588 32180 12640
rect 32404 12631 32456 12640
rect 32404 12597 32413 12631
rect 32413 12597 32447 12631
rect 32447 12597 32456 12631
rect 32404 12588 32456 12597
rect 33140 12588 33192 12640
rect 33784 12656 33836 12708
rect 33968 12699 34020 12708
rect 33968 12665 33977 12699
rect 33977 12665 34011 12699
rect 34011 12665 34020 12699
rect 33968 12656 34020 12665
rect 35256 12733 35265 12767
rect 35265 12733 35299 12767
rect 35299 12733 35308 12767
rect 35256 12724 35308 12733
rect 35440 12767 35492 12776
rect 35440 12733 35449 12767
rect 35449 12733 35483 12767
rect 35483 12733 35492 12767
rect 35440 12724 35492 12733
rect 33508 12631 33560 12640
rect 33508 12597 33517 12631
rect 33517 12597 33551 12631
rect 33551 12597 33560 12631
rect 33508 12588 33560 12597
rect 34428 12588 34480 12640
rect 38568 12860 38620 12912
rect 36636 12792 36688 12844
rect 37188 12792 37240 12844
rect 37004 12767 37056 12776
rect 37004 12733 37013 12767
rect 37013 12733 37047 12767
rect 37047 12733 37056 12767
rect 37924 12767 37976 12776
rect 37004 12724 37056 12733
rect 37924 12733 37933 12767
rect 37933 12733 37967 12767
rect 37967 12733 37976 12767
rect 37924 12724 37976 12733
rect 38844 12767 38896 12776
rect 38844 12733 38853 12767
rect 38853 12733 38887 12767
rect 38887 12733 38896 12767
rect 38844 12724 38896 12733
rect 19606 12486 19658 12538
rect 19670 12486 19722 12538
rect 19734 12486 19786 12538
rect 19798 12486 19850 12538
rect 3792 12316 3844 12368
rect 2044 12291 2096 12300
rect 2044 12257 2053 12291
rect 2053 12257 2087 12291
rect 2087 12257 2096 12291
rect 2044 12248 2096 12257
rect 2320 12248 2372 12300
rect 6184 12248 6236 12300
rect 7380 12291 7432 12300
rect 7380 12257 7389 12291
rect 7389 12257 7423 12291
rect 7423 12257 7432 12291
rect 7380 12248 7432 12257
rect 7932 12291 7984 12300
rect 7932 12257 7941 12291
rect 7941 12257 7975 12291
rect 7975 12257 7984 12291
rect 7932 12248 7984 12257
rect 8024 12248 8076 12300
rect 10140 12291 10192 12300
rect 10140 12257 10149 12291
rect 10149 12257 10183 12291
rect 10183 12257 10192 12291
rect 10140 12248 10192 12257
rect 10324 12291 10376 12300
rect 10324 12257 10333 12291
rect 10333 12257 10367 12291
rect 10367 12257 10376 12291
rect 10324 12248 10376 12257
rect 10508 12291 10560 12300
rect 10508 12257 10517 12291
rect 10517 12257 10551 12291
rect 10551 12257 10560 12291
rect 10508 12248 10560 12257
rect 5172 12223 5224 12232
rect 5172 12189 5181 12223
rect 5181 12189 5215 12223
rect 5215 12189 5224 12223
rect 5172 12180 5224 12189
rect 5448 12223 5500 12232
rect 5448 12189 5457 12223
rect 5457 12189 5491 12223
rect 5491 12189 5500 12223
rect 5448 12180 5500 12189
rect 12900 12384 12952 12436
rect 12256 12316 12308 12368
rect 15108 12316 15160 12368
rect 12900 12248 12952 12300
rect 13728 12248 13780 12300
rect 15200 12248 15252 12300
rect 16764 12316 16816 12368
rect 19064 12384 19116 12436
rect 16948 12248 17000 12300
rect 9956 12155 10008 12164
rect 9956 12121 9965 12155
rect 9965 12121 9999 12155
rect 9999 12121 10008 12155
rect 9956 12112 10008 12121
rect 2320 12044 2372 12096
rect 6920 12044 6972 12096
rect 12900 12112 12952 12164
rect 16672 12112 16724 12164
rect 14464 12087 14516 12096
rect 14464 12053 14473 12087
rect 14473 12053 14507 12087
rect 14507 12053 14516 12087
rect 14464 12044 14516 12053
rect 14648 12044 14700 12096
rect 18144 12316 18196 12368
rect 19340 12316 19392 12368
rect 18420 12291 18472 12300
rect 18420 12257 18429 12291
rect 18429 12257 18463 12291
rect 18463 12257 18472 12291
rect 18420 12248 18472 12257
rect 19248 12248 19300 12300
rect 19892 12223 19944 12232
rect 19892 12189 19901 12223
rect 19901 12189 19935 12223
rect 19935 12189 19944 12223
rect 19892 12180 19944 12189
rect 21364 12316 21416 12368
rect 20720 12248 20772 12300
rect 20812 12248 20864 12300
rect 22560 12384 22612 12436
rect 22468 12316 22520 12368
rect 25320 12384 25372 12436
rect 26056 12384 26108 12436
rect 28724 12427 28776 12436
rect 28724 12393 28733 12427
rect 28733 12393 28767 12427
rect 28767 12393 28776 12427
rect 28724 12384 28776 12393
rect 29736 12384 29788 12436
rect 31392 12384 31444 12436
rect 33784 12384 33836 12436
rect 34336 12384 34388 12436
rect 34428 12384 34480 12436
rect 38936 12384 38988 12436
rect 22284 12291 22336 12300
rect 22284 12257 22293 12291
rect 22293 12257 22327 12291
rect 22327 12257 22336 12291
rect 22284 12248 22336 12257
rect 23388 12248 23440 12300
rect 24952 12316 25004 12368
rect 30104 12316 30156 12368
rect 25044 12248 25096 12300
rect 26056 12248 26108 12300
rect 26516 12291 26568 12300
rect 26516 12257 26525 12291
rect 26525 12257 26559 12291
rect 26559 12257 26568 12291
rect 26516 12248 26568 12257
rect 27160 12291 27212 12300
rect 27160 12257 27169 12291
rect 27169 12257 27203 12291
rect 27203 12257 27212 12291
rect 27160 12248 27212 12257
rect 27528 12248 27580 12300
rect 30564 12316 30616 12368
rect 30932 12316 30984 12368
rect 32680 12316 32732 12368
rect 30656 12291 30708 12300
rect 30656 12257 30665 12291
rect 30665 12257 30699 12291
rect 30699 12257 30708 12291
rect 30656 12248 30708 12257
rect 30748 12248 30800 12300
rect 31668 12248 31720 12300
rect 32496 12248 32548 12300
rect 33968 12248 34020 12300
rect 34612 12291 34664 12300
rect 34612 12257 34621 12291
rect 34621 12257 34655 12291
rect 34655 12257 34664 12291
rect 34612 12248 34664 12257
rect 37280 12316 37332 12368
rect 36084 12291 36136 12300
rect 36084 12257 36093 12291
rect 36093 12257 36127 12291
rect 36127 12257 36136 12291
rect 36084 12248 36136 12257
rect 20628 12112 20680 12164
rect 21364 12112 21416 12164
rect 21548 12155 21600 12164
rect 21548 12121 21557 12155
rect 21557 12121 21591 12155
rect 21591 12121 21600 12155
rect 21548 12112 21600 12121
rect 23480 12112 23532 12164
rect 30748 12155 30800 12164
rect 17684 12044 17736 12096
rect 17776 12044 17828 12096
rect 21640 12044 21692 12096
rect 23388 12044 23440 12096
rect 24952 12044 25004 12096
rect 30748 12121 30757 12155
rect 30757 12121 30791 12155
rect 30791 12121 30800 12155
rect 30748 12112 30800 12121
rect 31392 12223 31444 12232
rect 31392 12189 31401 12223
rect 31401 12189 31435 12223
rect 31435 12189 31444 12223
rect 31392 12180 31444 12189
rect 31668 12112 31720 12164
rect 33784 12112 33836 12164
rect 29092 12044 29144 12096
rect 30196 12044 30248 12096
rect 33508 12044 33560 12096
rect 34428 12180 34480 12232
rect 34796 12180 34848 12232
rect 35992 12180 36044 12232
rect 36452 12180 36504 12232
rect 33968 12112 34020 12164
rect 34520 12044 34572 12096
rect 35348 12044 35400 12096
rect 37832 12248 37884 12300
rect 38200 12248 38252 12300
rect 38568 12291 38620 12300
rect 38568 12257 38577 12291
rect 38577 12257 38611 12291
rect 38611 12257 38620 12291
rect 38568 12248 38620 12257
rect 38752 12223 38804 12232
rect 38752 12189 38761 12223
rect 38761 12189 38795 12223
rect 38795 12189 38804 12223
rect 38752 12180 38804 12189
rect 37740 12112 37792 12164
rect 4246 11942 4298 11994
rect 4310 11942 4362 11994
rect 4374 11942 4426 11994
rect 4438 11942 4490 11994
rect 34966 11942 35018 11994
rect 35030 11942 35082 11994
rect 35094 11942 35146 11994
rect 35158 11942 35210 11994
rect 5724 11840 5776 11892
rect 6184 11883 6236 11892
rect 6184 11849 6193 11883
rect 6193 11849 6227 11883
rect 6227 11849 6236 11883
rect 6184 11840 6236 11849
rect 7196 11883 7248 11892
rect 7196 11849 7205 11883
rect 7205 11849 7239 11883
rect 7239 11849 7248 11883
rect 7196 11840 7248 11849
rect 12348 11840 12400 11892
rect 14464 11840 14516 11892
rect 15568 11840 15620 11892
rect 10140 11772 10192 11824
rect 12716 11815 12768 11824
rect 3516 11704 3568 11756
rect 3332 11679 3384 11688
rect 3332 11645 3341 11679
rect 3341 11645 3375 11679
rect 3375 11645 3384 11679
rect 3332 11636 3384 11645
rect 6920 11636 6972 11688
rect 7564 11636 7616 11688
rect 8300 11704 8352 11756
rect 10324 11704 10376 11756
rect 10508 11747 10560 11756
rect 10508 11713 10517 11747
rect 10517 11713 10551 11747
rect 10551 11713 10560 11747
rect 10508 11704 10560 11713
rect 11428 11747 11480 11756
rect 11428 11713 11437 11747
rect 11437 11713 11471 11747
rect 11471 11713 11480 11747
rect 11428 11704 11480 11713
rect 12716 11781 12725 11815
rect 12725 11781 12759 11815
rect 12759 11781 12768 11815
rect 12716 11772 12768 11781
rect 14372 11772 14424 11824
rect 8484 11679 8536 11688
rect 7932 11568 7984 11620
rect 8484 11645 8493 11679
rect 8493 11645 8527 11679
rect 8527 11645 8536 11679
rect 8484 11636 8536 11645
rect 9680 11636 9732 11688
rect 9680 11500 9732 11552
rect 10048 11636 10100 11688
rect 11336 11679 11388 11688
rect 11336 11645 11345 11679
rect 11345 11645 11379 11679
rect 11379 11645 11388 11679
rect 11336 11636 11388 11645
rect 11704 11679 11756 11688
rect 11704 11645 11713 11679
rect 11713 11645 11747 11679
rect 11747 11645 11756 11679
rect 11704 11636 11756 11645
rect 13544 11704 13596 11756
rect 17776 11772 17828 11824
rect 18236 11840 18288 11892
rect 19892 11840 19944 11892
rect 21640 11840 21692 11892
rect 23480 11840 23532 11892
rect 23756 11883 23808 11892
rect 23756 11849 23765 11883
rect 23765 11849 23799 11883
rect 23799 11849 23808 11883
rect 23756 11840 23808 11849
rect 23940 11840 23992 11892
rect 24216 11840 24268 11892
rect 13084 11679 13136 11688
rect 13084 11645 13093 11679
rect 13093 11645 13127 11679
rect 13127 11645 13136 11679
rect 13084 11636 13136 11645
rect 13268 11679 13320 11688
rect 13268 11645 13277 11679
rect 13277 11645 13311 11679
rect 13311 11645 13320 11679
rect 13268 11636 13320 11645
rect 17868 11704 17920 11756
rect 13636 11568 13688 11620
rect 9956 11500 10008 11552
rect 11244 11500 11296 11552
rect 14096 11500 14148 11552
rect 15108 11679 15160 11688
rect 15108 11645 15117 11679
rect 15117 11645 15151 11679
rect 15151 11645 15160 11679
rect 15108 11636 15160 11645
rect 16212 11679 16264 11688
rect 16212 11645 16221 11679
rect 16221 11645 16255 11679
rect 16255 11645 16264 11679
rect 16212 11636 16264 11645
rect 16580 11679 16632 11688
rect 16580 11645 16589 11679
rect 16589 11645 16623 11679
rect 16623 11645 16632 11679
rect 16580 11636 16632 11645
rect 17132 11679 17184 11688
rect 17132 11645 17141 11679
rect 17141 11645 17175 11679
rect 17175 11645 17184 11679
rect 17132 11636 17184 11645
rect 18512 11679 18564 11688
rect 18512 11645 18521 11679
rect 18521 11645 18555 11679
rect 18555 11645 18564 11679
rect 18512 11636 18564 11645
rect 23388 11772 23440 11824
rect 19248 11747 19300 11756
rect 19248 11713 19257 11747
rect 19257 11713 19291 11747
rect 19291 11713 19300 11747
rect 19248 11704 19300 11713
rect 19892 11704 19944 11756
rect 20352 11679 20404 11688
rect 20352 11645 20361 11679
rect 20361 11645 20395 11679
rect 20395 11645 20404 11679
rect 20352 11636 20404 11645
rect 22652 11704 22704 11756
rect 26332 11840 26384 11892
rect 27160 11840 27212 11892
rect 30472 11840 30524 11892
rect 38936 11883 38988 11892
rect 30748 11772 30800 11824
rect 32496 11815 32548 11824
rect 28908 11704 28960 11756
rect 32496 11781 32505 11815
rect 32505 11781 32539 11815
rect 32539 11781 32548 11815
rect 32496 11772 32548 11781
rect 33324 11772 33376 11824
rect 20996 11636 21048 11688
rect 21364 11679 21416 11688
rect 21364 11645 21373 11679
rect 21373 11645 21407 11679
rect 21407 11645 21416 11679
rect 21364 11636 21416 11645
rect 23296 11636 23348 11688
rect 24216 11636 24268 11688
rect 24492 11679 24544 11688
rect 24492 11645 24501 11679
rect 24501 11645 24535 11679
rect 24535 11645 24544 11679
rect 24492 11636 24544 11645
rect 24952 11679 25004 11688
rect 24952 11645 24961 11679
rect 24961 11645 24995 11679
rect 24995 11645 25004 11679
rect 24952 11636 25004 11645
rect 25136 11636 25188 11688
rect 16488 11568 16540 11620
rect 20168 11568 20220 11620
rect 22008 11500 22060 11552
rect 22284 11500 22336 11552
rect 23388 11500 23440 11552
rect 24768 11568 24820 11620
rect 25320 11568 25372 11620
rect 25596 11568 25648 11620
rect 27620 11636 27672 11688
rect 28540 11679 28592 11688
rect 28540 11645 28549 11679
rect 28549 11645 28583 11679
rect 28583 11645 28592 11679
rect 28540 11636 28592 11645
rect 30196 11636 30248 11688
rect 30564 11636 30616 11688
rect 31484 11636 31536 11688
rect 33600 11679 33652 11688
rect 26700 11500 26752 11552
rect 30748 11568 30800 11620
rect 33232 11568 33284 11620
rect 33600 11645 33609 11679
rect 33609 11645 33643 11679
rect 33643 11645 33652 11679
rect 33600 11636 33652 11645
rect 33876 11772 33928 11824
rect 38936 11849 38945 11883
rect 38945 11849 38979 11883
rect 38979 11849 38988 11883
rect 38936 11840 38988 11849
rect 34428 11772 34480 11824
rect 35348 11679 35400 11688
rect 35348 11645 35357 11679
rect 35357 11645 35391 11679
rect 35391 11645 35400 11679
rect 35348 11636 35400 11645
rect 35532 11679 35584 11688
rect 35532 11645 35541 11679
rect 35541 11645 35575 11679
rect 35575 11645 35584 11679
rect 35532 11636 35584 11645
rect 35808 11636 35860 11688
rect 35992 11679 36044 11688
rect 35992 11645 36001 11679
rect 36001 11645 36035 11679
rect 36035 11645 36044 11679
rect 36820 11679 36872 11688
rect 35992 11636 36044 11645
rect 36820 11645 36829 11679
rect 36829 11645 36863 11679
rect 36863 11645 36872 11679
rect 36820 11636 36872 11645
rect 37372 11679 37424 11688
rect 37372 11645 37381 11679
rect 37381 11645 37415 11679
rect 37415 11645 37424 11679
rect 37372 11636 37424 11645
rect 37188 11568 37240 11620
rect 37832 11636 37884 11688
rect 38384 11568 38436 11620
rect 29920 11500 29972 11552
rect 32496 11500 32548 11552
rect 36176 11500 36228 11552
rect 19606 11398 19658 11450
rect 19670 11398 19722 11450
rect 19734 11398 19786 11450
rect 19798 11398 19850 11450
rect 2320 11160 2372 11212
rect 3240 11203 3292 11212
rect 3240 11169 3249 11203
rect 3249 11169 3283 11203
rect 3283 11169 3292 11203
rect 3240 11160 3292 11169
rect 3884 11160 3936 11212
rect 5356 11203 5408 11212
rect 5356 11169 5365 11203
rect 5365 11169 5399 11203
rect 5399 11169 5408 11203
rect 5356 11160 5408 11169
rect 6184 11228 6236 11280
rect 10324 11296 10376 11348
rect 13728 11296 13780 11348
rect 3332 11135 3384 11144
rect 3332 11101 3341 11135
rect 3341 11101 3375 11135
rect 3375 11101 3384 11135
rect 3332 11092 3384 11101
rect 5448 11135 5500 11144
rect 5448 11101 5457 11135
rect 5457 11101 5491 11135
rect 5491 11101 5500 11135
rect 5448 11092 5500 11101
rect 7104 11228 7156 11280
rect 7012 11160 7064 11212
rect 8024 11203 8076 11212
rect 8024 11169 8033 11203
rect 8033 11169 8067 11203
rect 8067 11169 8076 11203
rect 8024 11160 8076 11169
rect 9036 11228 9088 11280
rect 9772 11203 9824 11212
rect 9772 11169 9781 11203
rect 9781 11169 9815 11203
rect 9815 11169 9824 11203
rect 9772 11160 9824 11169
rect 10048 11203 10100 11212
rect 10048 11169 10057 11203
rect 10057 11169 10091 11203
rect 10091 11169 10100 11203
rect 10048 11160 10100 11169
rect 11704 11228 11756 11280
rect 13084 11228 13136 11280
rect 18880 11296 18932 11348
rect 20628 11296 20680 11348
rect 30196 11296 30248 11348
rect 31208 11296 31260 11348
rect 31576 11296 31628 11348
rect 35532 11296 35584 11348
rect 35900 11296 35952 11348
rect 20352 11271 20404 11280
rect 10784 11160 10836 11212
rect 11612 11203 11664 11212
rect 11612 11169 11621 11203
rect 11621 11169 11655 11203
rect 11655 11169 11664 11203
rect 11612 11160 11664 11169
rect 12072 11203 12124 11212
rect 12072 11169 12081 11203
rect 12081 11169 12115 11203
rect 12115 11169 12124 11203
rect 12072 11160 12124 11169
rect 12164 11160 12216 11212
rect 20352 11237 20361 11271
rect 20361 11237 20395 11271
rect 20395 11237 20404 11271
rect 20352 11228 20404 11237
rect 22468 11228 22520 11280
rect 13544 11203 13596 11212
rect 13544 11169 13553 11203
rect 13553 11169 13587 11203
rect 13587 11169 13596 11203
rect 13544 11160 13596 11169
rect 13912 11203 13964 11212
rect 13912 11169 13921 11203
rect 13921 11169 13955 11203
rect 13955 11169 13964 11203
rect 13912 11160 13964 11169
rect 14464 11160 14516 11212
rect 14648 11203 14700 11212
rect 14648 11169 14657 11203
rect 14657 11169 14691 11203
rect 14691 11169 14700 11203
rect 15292 11203 15344 11212
rect 14648 11160 14700 11169
rect 15292 11169 15301 11203
rect 15301 11169 15335 11203
rect 15335 11169 15344 11203
rect 15292 11160 15344 11169
rect 16948 11160 17000 11212
rect 18512 11203 18564 11212
rect 18512 11169 18521 11203
rect 18521 11169 18555 11203
rect 18555 11169 18564 11203
rect 18512 11160 18564 11169
rect 16120 11092 16172 11144
rect 16488 11135 16540 11144
rect 16488 11101 16497 11135
rect 16497 11101 16531 11135
rect 16531 11101 16540 11135
rect 16488 11092 16540 11101
rect 10968 11067 11020 11076
rect 4620 10956 4672 11008
rect 10968 11033 10977 11067
rect 10977 11033 11011 11067
rect 11011 11033 11020 11067
rect 10968 11024 11020 11033
rect 13452 11024 13504 11076
rect 15568 11024 15620 11076
rect 16212 11024 16264 11076
rect 19340 11160 19392 11212
rect 19984 11160 20036 11212
rect 20168 11203 20220 11212
rect 20168 11169 20177 11203
rect 20177 11169 20211 11203
rect 20211 11169 20220 11203
rect 20168 11160 20220 11169
rect 21548 11203 21600 11212
rect 21548 11169 21557 11203
rect 21557 11169 21591 11203
rect 21591 11169 21600 11203
rect 21548 11160 21600 11169
rect 21916 11160 21968 11212
rect 22836 11203 22888 11212
rect 22836 11169 22845 11203
rect 22845 11169 22879 11203
rect 22879 11169 22888 11203
rect 22836 11160 22888 11169
rect 23296 11203 23348 11212
rect 23296 11169 23305 11203
rect 23305 11169 23339 11203
rect 23339 11169 23348 11203
rect 23296 11160 23348 11169
rect 21640 11092 21692 11144
rect 24768 11203 24820 11212
rect 24768 11169 24777 11203
rect 24777 11169 24811 11203
rect 24811 11169 24820 11203
rect 24768 11160 24820 11169
rect 25320 11203 25372 11212
rect 25320 11169 25329 11203
rect 25329 11169 25363 11203
rect 25363 11169 25372 11203
rect 25320 11160 25372 11169
rect 26700 11228 26752 11280
rect 31392 11228 31444 11280
rect 26608 11203 26660 11212
rect 26608 11169 26617 11203
rect 26617 11169 26651 11203
rect 26651 11169 26660 11203
rect 26608 11160 26660 11169
rect 27344 11160 27396 11212
rect 29920 11203 29972 11212
rect 29920 11169 29929 11203
rect 29929 11169 29963 11203
rect 29963 11169 29972 11203
rect 29920 11160 29972 11169
rect 30840 11160 30892 11212
rect 31116 11160 31168 11212
rect 33140 11160 33192 11212
rect 33324 11203 33376 11212
rect 33324 11169 33333 11203
rect 33333 11169 33367 11203
rect 33367 11169 33376 11203
rect 33324 11160 33376 11169
rect 33784 11228 33836 11280
rect 22008 11024 22060 11076
rect 23112 11024 23164 11076
rect 7472 10956 7524 11008
rect 14096 10956 14148 11008
rect 16580 10956 16632 11008
rect 25136 11024 25188 11076
rect 25688 10956 25740 11008
rect 28540 11024 28592 11076
rect 31484 11092 31536 11144
rect 34520 11160 34572 11212
rect 34796 11203 34848 11212
rect 34796 11169 34805 11203
rect 34805 11169 34839 11203
rect 34839 11169 34848 11203
rect 34796 11160 34848 11169
rect 35808 11228 35860 11280
rect 36176 11271 36228 11280
rect 36176 11237 36185 11271
rect 36185 11237 36219 11271
rect 36219 11237 36228 11271
rect 36176 11228 36228 11237
rect 35992 11160 36044 11212
rect 36452 11203 36504 11212
rect 36452 11169 36461 11203
rect 36461 11169 36495 11203
rect 36495 11169 36504 11203
rect 36452 11160 36504 11169
rect 27252 10956 27304 11008
rect 27712 10956 27764 11008
rect 27896 10956 27948 11008
rect 28080 10956 28132 11008
rect 31668 11024 31720 11076
rect 38200 11228 38252 11280
rect 35900 10956 35952 11008
rect 36360 10956 36412 11008
rect 38568 11203 38620 11212
rect 38568 11169 38577 11203
rect 38577 11169 38611 11203
rect 38611 11169 38620 11203
rect 38568 11160 38620 11169
rect 37832 11135 37884 11144
rect 37832 11101 37841 11135
rect 37841 11101 37875 11135
rect 37875 11101 37884 11135
rect 37832 11092 37884 11101
rect 4246 10854 4298 10906
rect 4310 10854 4362 10906
rect 4374 10854 4426 10906
rect 4438 10854 4490 10906
rect 34966 10854 35018 10906
rect 35030 10854 35082 10906
rect 35094 10854 35146 10906
rect 35158 10854 35210 10906
rect 2504 10795 2556 10804
rect 2504 10761 2513 10795
rect 2513 10761 2547 10795
rect 2547 10761 2556 10795
rect 2504 10752 2556 10761
rect 3240 10752 3292 10804
rect 3884 10752 3936 10804
rect 7104 10752 7156 10804
rect 7564 10752 7616 10804
rect 9036 10795 9088 10804
rect 9036 10761 9045 10795
rect 9045 10761 9079 10795
rect 9079 10761 9088 10795
rect 9036 10752 9088 10761
rect 10692 10752 10744 10804
rect 28080 10752 28132 10804
rect 31208 10752 31260 10804
rect 2872 10616 2924 10668
rect 2964 10548 3016 10600
rect 4620 10616 4672 10668
rect 4344 10548 4396 10600
rect 6184 10548 6236 10600
rect 12624 10684 12676 10736
rect 13268 10727 13320 10736
rect 13268 10693 13277 10727
rect 13277 10693 13311 10727
rect 13311 10693 13320 10727
rect 13268 10684 13320 10693
rect 16120 10684 16172 10736
rect 8484 10616 8536 10668
rect 7656 10591 7708 10600
rect 7656 10557 7665 10591
rect 7665 10557 7699 10591
rect 7699 10557 7708 10591
rect 7656 10548 7708 10557
rect 9036 10616 9088 10668
rect 8852 10591 8904 10600
rect 8852 10557 8861 10591
rect 8861 10557 8895 10591
rect 8895 10557 8904 10591
rect 10968 10616 11020 10668
rect 11980 10616 12032 10668
rect 12072 10616 12124 10668
rect 13912 10616 13964 10668
rect 17132 10659 17184 10668
rect 17132 10625 17141 10659
rect 17141 10625 17175 10659
rect 17175 10625 17184 10659
rect 17132 10616 17184 10625
rect 17868 10616 17920 10668
rect 9864 10591 9916 10600
rect 8852 10548 8904 10557
rect 9864 10557 9873 10591
rect 9873 10557 9907 10591
rect 9907 10557 9916 10591
rect 9864 10548 9916 10557
rect 11428 10591 11480 10600
rect 3608 10480 3660 10532
rect 1400 10412 1452 10464
rect 3516 10412 3568 10464
rect 8668 10480 8720 10532
rect 11428 10557 11437 10591
rect 11437 10557 11471 10591
rect 11471 10557 11480 10591
rect 11428 10548 11480 10557
rect 11704 10591 11756 10600
rect 11704 10557 11713 10591
rect 11713 10557 11747 10591
rect 11747 10557 11756 10591
rect 11704 10548 11756 10557
rect 12440 10591 12492 10600
rect 12440 10557 12449 10591
rect 12449 10557 12483 10591
rect 12483 10557 12492 10591
rect 12992 10591 13044 10600
rect 12440 10548 12492 10557
rect 12992 10557 13001 10591
rect 13001 10557 13035 10591
rect 13035 10557 13044 10591
rect 12992 10548 13044 10557
rect 13360 10591 13412 10600
rect 13360 10557 13369 10591
rect 13369 10557 13403 10591
rect 13403 10557 13412 10591
rect 13360 10548 13412 10557
rect 13636 10548 13688 10600
rect 14464 10591 14516 10600
rect 14464 10557 14473 10591
rect 14473 10557 14507 10591
rect 14507 10557 14516 10591
rect 14464 10548 14516 10557
rect 12348 10480 12400 10532
rect 12716 10480 12768 10532
rect 15292 10548 15344 10600
rect 15384 10548 15436 10600
rect 16580 10548 16632 10600
rect 17224 10548 17276 10600
rect 18420 10548 18472 10600
rect 19432 10548 19484 10600
rect 20536 10616 20588 10668
rect 21456 10616 21508 10668
rect 17960 10480 18012 10532
rect 20168 10548 20220 10600
rect 21640 10591 21692 10600
rect 21640 10557 21649 10591
rect 21649 10557 21683 10591
rect 21683 10557 21692 10591
rect 21640 10548 21692 10557
rect 22836 10616 22888 10668
rect 24584 10616 24636 10668
rect 25596 10616 25648 10668
rect 29460 10684 29512 10736
rect 38752 10752 38804 10804
rect 28080 10616 28132 10668
rect 22652 10591 22704 10600
rect 19984 10480 20036 10532
rect 21548 10480 21600 10532
rect 22652 10557 22661 10591
rect 22661 10557 22695 10591
rect 22695 10557 22704 10591
rect 22652 10548 22704 10557
rect 23204 10548 23256 10600
rect 24952 10591 25004 10600
rect 24952 10557 24961 10591
rect 24961 10557 24995 10591
rect 24995 10557 25004 10591
rect 24952 10548 25004 10557
rect 27068 10591 27120 10600
rect 27068 10557 27077 10591
rect 27077 10557 27111 10591
rect 27111 10557 27120 10591
rect 27068 10548 27120 10557
rect 27160 10591 27212 10600
rect 27160 10557 27169 10591
rect 27169 10557 27203 10591
rect 27203 10557 27212 10591
rect 27528 10591 27580 10600
rect 27160 10548 27212 10557
rect 27528 10557 27537 10591
rect 27537 10557 27571 10591
rect 27571 10557 27580 10591
rect 27528 10548 27580 10557
rect 27988 10548 28040 10600
rect 23296 10480 23348 10532
rect 26056 10480 26108 10532
rect 28080 10480 28132 10532
rect 28448 10480 28500 10532
rect 28632 10548 28684 10600
rect 29460 10591 29512 10600
rect 29460 10557 29469 10591
rect 29469 10557 29503 10591
rect 29503 10557 29512 10591
rect 29460 10548 29512 10557
rect 31392 10548 31444 10600
rect 35624 10616 35676 10668
rect 37280 10684 37332 10736
rect 36360 10616 36412 10668
rect 37740 10659 37792 10668
rect 37740 10625 37749 10659
rect 37749 10625 37783 10659
rect 37783 10625 37792 10659
rect 37740 10616 37792 10625
rect 37832 10616 37884 10668
rect 31760 10548 31812 10600
rect 32220 10548 32272 10600
rect 33232 10591 33284 10600
rect 12624 10412 12676 10464
rect 13084 10412 13136 10464
rect 13728 10412 13780 10464
rect 14188 10412 14240 10464
rect 15476 10412 15528 10464
rect 16396 10412 16448 10464
rect 19340 10412 19392 10464
rect 22008 10412 22060 10464
rect 22284 10412 22336 10464
rect 26148 10412 26200 10464
rect 27344 10412 27396 10464
rect 27712 10412 27764 10464
rect 31484 10480 31536 10532
rect 33232 10557 33241 10591
rect 33241 10557 33275 10591
rect 33275 10557 33284 10591
rect 33232 10548 33284 10557
rect 33508 10591 33560 10600
rect 33508 10557 33517 10591
rect 33517 10557 33551 10591
rect 33551 10557 33560 10591
rect 33508 10548 33560 10557
rect 33692 10548 33744 10600
rect 36728 10591 36780 10600
rect 36728 10557 36737 10591
rect 36737 10557 36771 10591
rect 36771 10557 36780 10591
rect 36728 10548 36780 10557
rect 37464 10591 37516 10600
rect 37464 10557 37473 10591
rect 37473 10557 37507 10591
rect 37507 10557 37516 10591
rect 37464 10548 37516 10557
rect 36084 10480 36136 10532
rect 36360 10480 36412 10532
rect 37556 10480 37608 10532
rect 30472 10455 30524 10464
rect 30472 10421 30481 10455
rect 30481 10421 30515 10455
rect 30515 10421 30524 10455
rect 30472 10412 30524 10421
rect 33140 10412 33192 10464
rect 33232 10412 33284 10464
rect 34336 10412 34388 10464
rect 34796 10412 34848 10464
rect 38936 10412 38988 10464
rect 19606 10310 19658 10362
rect 19670 10310 19722 10362
rect 19734 10310 19786 10362
rect 19798 10310 19850 10362
rect 4344 10208 4396 10260
rect 7656 10208 7708 10260
rect 5356 10140 5408 10192
rect 13084 10208 13136 10260
rect 13176 10208 13228 10260
rect 13728 10208 13780 10260
rect 12716 10140 12768 10192
rect 15292 10183 15344 10192
rect 2504 10072 2556 10124
rect 4988 10072 5040 10124
rect 5172 10072 5224 10124
rect 6184 10115 6236 10124
rect 6184 10081 6193 10115
rect 6193 10081 6227 10115
rect 6227 10081 6236 10115
rect 6184 10072 6236 10081
rect 6920 10072 6972 10124
rect 8852 10115 8904 10124
rect 8852 10081 8867 10115
rect 8867 10081 8901 10115
rect 8901 10081 8904 10115
rect 10508 10115 10560 10124
rect 8852 10072 8904 10081
rect 10508 10081 10517 10115
rect 10517 10081 10551 10115
rect 10551 10081 10560 10115
rect 10508 10072 10560 10081
rect 10784 10115 10836 10124
rect 10784 10081 10793 10115
rect 10793 10081 10827 10115
rect 10827 10081 10836 10115
rect 10784 10072 10836 10081
rect 12532 10115 12584 10124
rect 1400 10047 1452 10056
rect 1400 10013 1409 10047
rect 1409 10013 1443 10047
rect 1443 10013 1452 10047
rect 1400 10004 1452 10013
rect 2780 10047 2832 10056
rect 2780 10013 2789 10047
rect 2789 10013 2823 10047
rect 2823 10013 2832 10047
rect 2780 10004 2832 10013
rect 4712 10004 4764 10056
rect 8208 10004 8260 10056
rect 8576 10004 8628 10056
rect 9588 10004 9640 10056
rect 12532 10081 12541 10115
rect 12541 10081 12575 10115
rect 12575 10081 12584 10115
rect 12532 10072 12584 10081
rect 13544 10072 13596 10124
rect 13912 10115 13964 10124
rect 13912 10081 13921 10115
rect 13921 10081 13955 10115
rect 13955 10081 13964 10115
rect 13912 10072 13964 10081
rect 15292 10149 15301 10183
rect 15301 10149 15335 10183
rect 15335 10149 15344 10183
rect 15292 10140 15344 10149
rect 16580 10072 16632 10124
rect 14188 10004 14240 10056
rect 9680 9936 9732 9988
rect 12808 9936 12860 9988
rect 15752 10004 15804 10056
rect 16396 10047 16448 10056
rect 16396 10013 16405 10047
rect 16405 10013 16439 10047
rect 16439 10013 16448 10047
rect 16396 10004 16448 10013
rect 17224 10072 17276 10124
rect 17960 10115 18012 10124
rect 17960 10081 17969 10115
rect 17969 10081 18003 10115
rect 18003 10081 18012 10115
rect 17960 10072 18012 10081
rect 19156 10072 19208 10124
rect 19340 10115 19392 10124
rect 19340 10081 19349 10115
rect 19349 10081 19383 10115
rect 19383 10081 19392 10115
rect 19340 10072 19392 10081
rect 19892 10115 19944 10124
rect 19892 10081 19901 10115
rect 19901 10081 19935 10115
rect 19935 10081 19944 10115
rect 19892 10072 19944 10081
rect 18328 10004 18380 10056
rect 5448 9868 5500 9920
rect 10508 9868 10560 9920
rect 12072 9868 12124 9920
rect 12716 9868 12768 9920
rect 17224 9868 17276 9920
rect 18420 9868 18472 9920
rect 19984 9868 20036 9920
rect 22836 10208 22888 10260
rect 24216 10208 24268 10260
rect 27160 10208 27212 10260
rect 27620 10251 27672 10260
rect 27620 10217 27629 10251
rect 27629 10217 27663 10251
rect 27663 10217 27672 10251
rect 27620 10208 27672 10217
rect 23756 10140 23808 10192
rect 25320 10140 25372 10192
rect 21548 10115 21600 10124
rect 21548 10081 21557 10115
rect 21557 10081 21591 10115
rect 21591 10081 21600 10115
rect 21548 10072 21600 10081
rect 21916 10115 21968 10124
rect 21916 10081 21925 10115
rect 21925 10081 21959 10115
rect 21959 10081 21968 10115
rect 21916 10072 21968 10081
rect 23388 10072 23440 10124
rect 21456 10047 21508 10056
rect 21456 10013 21465 10047
rect 21465 10013 21499 10047
rect 21499 10013 21508 10047
rect 21456 10004 21508 10013
rect 22008 10047 22060 10056
rect 22008 10013 22017 10047
rect 22017 10013 22051 10047
rect 22051 10013 22060 10047
rect 22008 10004 22060 10013
rect 22744 10047 22796 10056
rect 22744 10013 22753 10047
rect 22753 10013 22787 10047
rect 22787 10013 22796 10047
rect 22744 10004 22796 10013
rect 24860 10072 24912 10124
rect 25688 10115 25740 10124
rect 25688 10081 25697 10115
rect 25697 10081 25731 10115
rect 25731 10081 25740 10115
rect 25688 10072 25740 10081
rect 27252 10140 27304 10192
rect 30380 10208 30432 10260
rect 31300 10208 31352 10260
rect 33508 10208 33560 10260
rect 37280 10208 37332 10260
rect 37372 10208 37424 10260
rect 28448 10115 28500 10124
rect 21272 9936 21324 9988
rect 27160 10004 27212 10056
rect 27896 10004 27948 10056
rect 27988 10004 28040 10056
rect 28448 10081 28457 10115
rect 28457 10081 28491 10115
rect 28491 10081 28500 10115
rect 28448 10072 28500 10081
rect 30564 10115 30616 10124
rect 30564 10081 30573 10115
rect 30573 10081 30607 10115
rect 30607 10081 30616 10115
rect 30564 10072 30616 10081
rect 30840 10072 30892 10124
rect 31116 10072 31168 10124
rect 30656 10004 30708 10056
rect 32312 10115 32364 10124
rect 32312 10081 32321 10115
rect 32321 10081 32355 10115
rect 32355 10081 32364 10115
rect 32680 10115 32732 10124
rect 32312 10072 32364 10081
rect 32680 10081 32689 10115
rect 32689 10081 32723 10115
rect 32723 10081 32732 10115
rect 32680 10072 32732 10081
rect 32772 10072 32824 10124
rect 33784 10072 33836 10124
rect 35624 10115 35676 10124
rect 35624 10081 35633 10115
rect 35633 10081 35667 10115
rect 35667 10081 35676 10115
rect 35624 10072 35676 10081
rect 35808 10115 35860 10124
rect 35808 10081 35817 10115
rect 35817 10081 35851 10115
rect 35851 10081 35860 10115
rect 35808 10072 35860 10081
rect 38016 10115 38068 10124
rect 38016 10081 38025 10115
rect 38025 10081 38059 10115
rect 38059 10081 38068 10115
rect 38016 10072 38068 10081
rect 38936 10115 38988 10124
rect 38936 10081 38945 10115
rect 38945 10081 38979 10115
rect 38979 10081 38988 10115
rect 38936 10072 38988 10081
rect 36452 10004 36504 10056
rect 27528 9936 27580 9988
rect 28080 9936 28132 9988
rect 29368 9936 29420 9988
rect 24676 9868 24728 9920
rect 28172 9868 28224 9920
rect 28632 9868 28684 9920
rect 30104 9868 30156 9920
rect 30564 9936 30616 9988
rect 31392 9936 31444 9988
rect 32312 9936 32364 9988
rect 35808 9936 35860 9988
rect 4246 9766 4298 9818
rect 4310 9766 4362 9818
rect 4374 9766 4426 9818
rect 4438 9766 4490 9818
rect 34966 9766 35018 9818
rect 35030 9766 35082 9818
rect 35094 9766 35146 9818
rect 35158 9766 35210 9818
rect 20168 9664 20220 9716
rect 22744 9664 22796 9716
rect 24584 9664 24636 9716
rect 4068 9596 4120 9648
rect 4620 9596 4672 9648
rect 10784 9596 10836 9648
rect 12808 9639 12860 9648
rect 12808 9605 12817 9639
rect 12817 9605 12851 9639
rect 12851 9605 12860 9639
rect 12808 9596 12860 9605
rect 13636 9639 13688 9648
rect 13636 9605 13645 9639
rect 13645 9605 13679 9639
rect 13679 9605 13688 9639
rect 13636 9596 13688 9605
rect 14464 9596 14516 9648
rect 4712 9528 4764 9580
rect 2320 9503 2372 9512
rect 2320 9469 2329 9503
rect 2329 9469 2363 9503
rect 2363 9469 2372 9503
rect 2320 9460 2372 9469
rect 3884 9503 3936 9512
rect 1676 9324 1728 9376
rect 3884 9469 3893 9503
rect 3893 9469 3927 9503
rect 3927 9469 3936 9503
rect 3884 9460 3936 9469
rect 4436 9392 4488 9444
rect 5172 9392 5224 9444
rect 6092 9392 6144 9444
rect 4160 9324 4212 9376
rect 4896 9324 4948 9376
rect 6184 9324 6236 9376
rect 7288 9503 7340 9512
rect 6460 9392 6512 9444
rect 7288 9469 7297 9503
rect 7297 9469 7331 9503
rect 7331 9469 7340 9503
rect 7288 9460 7340 9469
rect 7748 9528 7800 9580
rect 12532 9528 12584 9580
rect 9956 9503 10008 9512
rect 9956 9469 9965 9503
rect 9965 9469 9999 9503
rect 9999 9469 10008 9503
rect 9956 9460 10008 9469
rect 8760 9392 8812 9444
rect 10600 9324 10652 9376
rect 10784 9503 10836 9512
rect 10784 9469 10793 9503
rect 10793 9469 10827 9503
rect 10827 9469 10836 9503
rect 10784 9460 10836 9469
rect 10968 9460 11020 9512
rect 12256 9460 12308 9512
rect 13268 9460 13320 9512
rect 13544 9503 13596 9512
rect 13544 9469 13553 9503
rect 13553 9469 13587 9503
rect 13587 9469 13596 9503
rect 13544 9460 13596 9469
rect 17408 9596 17460 9648
rect 18604 9596 18656 9648
rect 17316 9571 17368 9580
rect 17316 9537 17325 9571
rect 17325 9537 17359 9571
rect 17359 9537 17368 9571
rect 17316 9528 17368 9537
rect 19984 9528 20036 9580
rect 21456 9528 21508 9580
rect 22008 9596 22060 9648
rect 23296 9596 23348 9648
rect 24952 9596 25004 9648
rect 27436 9664 27488 9716
rect 30196 9664 30248 9716
rect 30380 9664 30432 9716
rect 31852 9664 31904 9716
rect 32680 9664 32732 9716
rect 33784 9664 33836 9716
rect 35716 9664 35768 9716
rect 38016 9664 38068 9716
rect 26240 9596 26292 9648
rect 27068 9596 27120 9648
rect 13728 9392 13780 9444
rect 15568 9503 15620 9512
rect 15568 9469 15577 9503
rect 15577 9469 15611 9503
rect 15611 9469 15620 9503
rect 15568 9460 15620 9469
rect 15660 9460 15712 9512
rect 16672 9460 16724 9512
rect 17224 9503 17276 9512
rect 17224 9469 17233 9503
rect 17233 9469 17267 9503
rect 17267 9469 17276 9503
rect 17224 9460 17276 9469
rect 18420 9503 18472 9512
rect 18420 9469 18429 9503
rect 18429 9469 18463 9503
rect 18463 9469 18472 9503
rect 18420 9460 18472 9469
rect 18788 9503 18840 9512
rect 18788 9469 18797 9503
rect 18797 9469 18831 9503
rect 18831 9469 18840 9503
rect 18788 9460 18840 9469
rect 19064 9460 19116 9512
rect 21640 9503 21692 9512
rect 21640 9469 21649 9503
rect 21649 9469 21683 9503
rect 21683 9469 21692 9503
rect 21640 9460 21692 9469
rect 21824 9460 21876 9512
rect 22836 9503 22888 9512
rect 22836 9469 22845 9503
rect 22845 9469 22879 9503
rect 22879 9469 22888 9503
rect 22836 9460 22888 9469
rect 23112 9460 23164 9512
rect 23664 9460 23716 9512
rect 12440 9324 12492 9376
rect 12808 9324 12860 9376
rect 15752 9324 15804 9376
rect 16028 9324 16080 9376
rect 20996 9324 21048 9376
rect 21824 9324 21876 9376
rect 24032 9324 24084 9376
rect 29000 9596 29052 9648
rect 30656 9639 30708 9648
rect 30656 9605 30665 9639
rect 30665 9605 30699 9639
rect 30699 9605 30708 9639
rect 30656 9596 30708 9605
rect 34060 9596 34112 9648
rect 34336 9596 34388 9648
rect 25320 9460 25372 9512
rect 27068 9503 27120 9512
rect 25044 9392 25096 9444
rect 24768 9324 24820 9376
rect 27068 9469 27077 9503
rect 27077 9469 27111 9503
rect 27111 9469 27120 9503
rect 27068 9460 27120 9469
rect 26332 9392 26384 9444
rect 27620 9503 27672 9512
rect 27620 9469 27629 9503
rect 27629 9469 27663 9503
rect 27663 9469 27672 9503
rect 27620 9460 27672 9469
rect 30472 9528 30524 9580
rect 31668 9528 31720 9580
rect 29092 9503 29144 9512
rect 29092 9469 29101 9503
rect 29101 9469 29135 9503
rect 29135 9469 29144 9503
rect 29092 9460 29144 9469
rect 29184 9460 29236 9512
rect 29368 9460 29420 9512
rect 31392 9503 31444 9512
rect 31392 9469 31401 9503
rect 31401 9469 31435 9503
rect 31435 9469 31444 9503
rect 31392 9460 31444 9469
rect 34520 9528 34572 9580
rect 35808 9571 35860 9580
rect 35808 9537 35817 9571
rect 35817 9537 35851 9571
rect 35851 9537 35860 9571
rect 35808 9528 35860 9537
rect 37372 9528 37424 9580
rect 32220 9503 32272 9512
rect 32220 9469 32229 9503
rect 32229 9469 32263 9503
rect 32263 9469 32272 9503
rect 32220 9460 32272 9469
rect 33968 9503 34020 9512
rect 28264 9392 28316 9444
rect 33968 9469 33977 9503
rect 33977 9469 34011 9503
rect 34011 9469 34020 9503
rect 33968 9460 34020 9469
rect 34060 9503 34112 9512
rect 34060 9469 34069 9503
rect 34069 9469 34103 9503
rect 34103 9469 34112 9503
rect 34060 9460 34112 9469
rect 35072 9460 35124 9512
rect 35716 9503 35768 9512
rect 35716 9469 35725 9503
rect 35725 9469 35759 9503
rect 35759 9469 35768 9503
rect 35716 9460 35768 9469
rect 37188 9503 37240 9512
rect 37188 9469 37197 9503
rect 37197 9469 37231 9503
rect 37231 9469 37240 9503
rect 37188 9460 37240 9469
rect 26516 9324 26568 9376
rect 29184 9324 29236 9376
rect 30840 9324 30892 9376
rect 31484 9367 31536 9376
rect 31484 9333 31493 9367
rect 31493 9333 31527 9367
rect 31527 9333 31536 9367
rect 31484 9324 31536 9333
rect 35256 9324 35308 9376
rect 19606 9222 19658 9274
rect 19670 9222 19722 9274
rect 19734 9222 19786 9274
rect 19798 9222 19850 9274
rect 2964 9163 3016 9172
rect 2964 9129 2973 9163
rect 2973 9129 3007 9163
rect 3007 9129 3016 9163
rect 2964 9120 3016 9129
rect 13360 9120 13412 9172
rect 15476 9120 15528 9172
rect 18328 9163 18380 9172
rect 18328 9129 18337 9163
rect 18337 9129 18371 9163
rect 18371 9129 18380 9163
rect 18328 9120 18380 9129
rect 21364 9120 21416 9172
rect 23388 9120 23440 9172
rect 1676 9027 1728 9036
rect 1676 8993 1685 9027
rect 1685 8993 1719 9027
rect 1719 8993 1728 9027
rect 1676 8984 1728 8993
rect 4068 8984 4120 9036
rect 4436 9027 4488 9036
rect 4436 8993 4445 9027
rect 4445 8993 4479 9027
rect 4479 8993 4488 9027
rect 4436 8984 4488 8993
rect 4896 9027 4948 9036
rect 4896 8993 4905 9027
rect 4905 8993 4939 9027
rect 4939 8993 4948 9027
rect 4896 8984 4948 8993
rect 5172 8984 5224 9036
rect 5448 9027 5500 9036
rect 5448 8993 5457 9027
rect 5457 8993 5491 9027
rect 5491 8993 5500 9027
rect 5448 8984 5500 8993
rect 6092 9027 6144 9036
rect 6092 8993 6101 9027
rect 6101 8993 6135 9027
rect 6135 8993 6144 9027
rect 6092 8984 6144 8993
rect 7104 8984 7156 9036
rect 7748 9027 7800 9036
rect 7748 8993 7757 9027
rect 7757 8993 7791 9027
rect 7791 8993 7800 9027
rect 7748 8984 7800 8993
rect 8116 9027 8168 9036
rect 8116 8993 8125 9027
rect 8125 8993 8159 9027
rect 8159 8993 8168 9027
rect 8116 8984 8168 8993
rect 9036 9027 9088 9036
rect 9036 8993 9045 9027
rect 9045 8993 9079 9027
rect 9079 8993 9088 9027
rect 9036 8984 9088 8993
rect 10140 8984 10192 9036
rect 12348 9027 12400 9036
rect 12348 8993 12357 9027
rect 12357 8993 12391 9027
rect 12391 8993 12400 9027
rect 12348 8984 12400 8993
rect 12716 9027 12768 9036
rect 12716 8993 12725 9027
rect 12725 8993 12759 9027
rect 12759 8993 12768 9027
rect 12716 8984 12768 8993
rect 13268 8984 13320 9036
rect 13728 8984 13780 9036
rect 15752 8984 15804 9036
rect 16304 9027 16356 9036
rect 16304 8993 16313 9027
rect 16313 8993 16347 9027
rect 16347 8993 16356 9027
rect 16304 8984 16356 8993
rect 1400 8959 1452 8968
rect 1400 8925 1409 8959
rect 1409 8925 1443 8959
rect 1443 8925 1452 8959
rect 1400 8916 1452 8925
rect 4804 8959 4856 8968
rect 4804 8925 4813 8959
rect 4813 8925 4847 8959
rect 4847 8925 4856 8959
rect 4804 8916 4856 8925
rect 7288 8959 7340 8968
rect 7288 8925 7297 8959
rect 7297 8925 7331 8959
rect 7331 8925 7340 8959
rect 7288 8916 7340 8925
rect 11152 8959 11204 8968
rect 11152 8925 11161 8959
rect 11161 8925 11195 8959
rect 11195 8925 11204 8959
rect 11152 8916 11204 8925
rect 12256 8959 12308 8968
rect 12256 8925 12265 8959
rect 12265 8925 12299 8959
rect 12299 8925 12308 8959
rect 12256 8916 12308 8925
rect 3700 8823 3752 8832
rect 3700 8789 3709 8823
rect 3709 8789 3743 8823
rect 3743 8789 3752 8823
rect 3700 8780 3752 8789
rect 14188 8916 14240 8968
rect 14372 8959 14424 8968
rect 14372 8925 14381 8959
rect 14381 8925 14415 8959
rect 14415 8925 14424 8959
rect 14372 8916 14424 8925
rect 15844 8959 15896 8968
rect 15844 8925 15853 8959
rect 15853 8925 15887 8959
rect 15887 8925 15896 8959
rect 15844 8916 15896 8925
rect 16212 8916 16264 8968
rect 16948 8959 17000 8968
rect 16948 8925 16957 8959
rect 16957 8925 16991 8959
rect 16991 8925 17000 8959
rect 16948 8916 17000 8925
rect 19064 9052 19116 9104
rect 19340 9052 19392 9104
rect 17316 8984 17368 9036
rect 19800 9027 19852 9036
rect 19800 8993 19809 9027
rect 19809 8993 19843 9027
rect 19843 8993 19852 9027
rect 19800 8984 19852 8993
rect 19892 9027 19944 9036
rect 19892 8993 19901 9027
rect 19901 8993 19935 9027
rect 19935 8993 19944 9027
rect 20168 9027 20220 9036
rect 19892 8984 19944 8993
rect 20168 8993 20177 9027
rect 20177 8993 20211 9027
rect 20211 8993 20220 9027
rect 20168 8984 20220 8993
rect 22192 9027 22244 9036
rect 13084 8848 13136 8900
rect 15660 8848 15712 8900
rect 13912 8780 13964 8832
rect 18052 8780 18104 8832
rect 19432 8916 19484 8968
rect 21364 8959 21416 8968
rect 21364 8925 21373 8959
rect 21373 8925 21407 8959
rect 21407 8925 21416 8959
rect 21364 8916 21416 8925
rect 21456 8916 21508 8968
rect 22192 8993 22201 9027
rect 22201 8993 22235 9027
rect 22235 8993 22244 9027
rect 22192 8984 22244 8993
rect 23756 9052 23808 9104
rect 24768 9120 24820 9172
rect 23480 8984 23532 9036
rect 23848 9027 23900 9036
rect 23388 8916 23440 8968
rect 23848 8993 23857 9027
rect 23857 8993 23891 9027
rect 23891 8993 23900 9027
rect 23848 8984 23900 8993
rect 24032 8916 24084 8968
rect 22100 8891 22152 8900
rect 22100 8857 22109 8891
rect 22109 8857 22143 8891
rect 22143 8857 22152 8891
rect 22100 8848 22152 8857
rect 26240 9120 26292 9172
rect 26884 9120 26936 9172
rect 30196 9163 30248 9172
rect 30196 9129 30205 9163
rect 30205 9129 30239 9163
rect 30239 9129 30248 9163
rect 30196 9120 30248 9129
rect 31484 9120 31536 9172
rect 36360 9163 36412 9172
rect 31208 9052 31260 9104
rect 31944 9052 31996 9104
rect 34244 9052 34296 9104
rect 35072 9052 35124 9104
rect 36360 9129 36369 9163
rect 36369 9129 36403 9163
rect 36403 9129 36412 9163
rect 36360 9120 36412 9129
rect 37188 9120 37240 9172
rect 25228 9027 25280 9036
rect 25228 8993 25237 9027
rect 25237 8993 25271 9027
rect 25271 8993 25280 9027
rect 25228 8984 25280 8993
rect 24860 8916 24912 8968
rect 26240 8984 26292 9036
rect 27436 8916 27488 8968
rect 27988 8959 28040 8968
rect 27988 8925 27997 8959
rect 27997 8925 28031 8959
rect 28031 8925 28040 8959
rect 27988 8916 28040 8925
rect 28356 8984 28408 9036
rect 30104 9027 30156 9036
rect 30104 8993 30113 9027
rect 30113 8993 30147 9027
rect 30147 8993 30156 9027
rect 30104 8984 30156 8993
rect 31024 8984 31076 9036
rect 33140 9027 33192 9036
rect 33140 8993 33149 9027
rect 33149 8993 33183 9027
rect 33183 8993 33192 9027
rect 33140 8984 33192 8993
rect 35256 9027 35308 9036
rect 35256 8993 35265 9027
rect 35265 8993 35299 9027
rect 35299 8993 35308 9027
rect 35256 8984 35308 8993
rect 37556 8984 37608 9036
rect 38476 9027 38528 9036
rect 38476 8993 38485 9027
rect 38485 8993 38519 9027
rect 38519 8993 38528 9027
rect 38476 8984 38528 8993
rect 31300 8916 31352 8968
rect 33508 8916 33560 8968
rect 34336 8916 34388 8968
rect 24952 8848 25004 8900
rect 29000 8848 29052 8900
rect 29828 8848 29880 8900
rect 31668 8848 31720 8900
rect 24860 8780 24912 8832
rect 25872 8780 25924 8832
rect 29276 8780 29328 8832
rect 31852 8780 31904 8832
rect 34428 8823 34480 8832
rect 34428 8789 34437 8823
rect 34437 8789 34471 8823
rect 34471 8789 34480 8823
rect 34428 8780 34480 8789
rect 4246 8678 4298 8730
rect 4310 8678 4362 8730
rect 4374 8678 4426 8730
rect 4438 8678 4490 8730
rect 34966 8678 35018 8730
rect 35030 8678 35082 8730
rect 35094 8678 35146 8730
rect 35158 8678 35210 8730
rect 4068 8619 4120 8628
rect 4068 8585 4077 8619
rect 4077 8585 4111 8619
rect 4111 8585 4120 8619
rect 4068 8576 4120 8585
rect 6184 8619 6236 8628
rect 6184 8585 6193 8619
rect 6193 8585 6227 8619
rect 6227 8585 6236 8619
rect 6184 8576 6236 8585
rect 12256 8576 12308 8628
rect 6460 8508 6512 8560
rect 12348 8508 12400 8560
rect 12900 8508 12952 8560
rect 13084 8551 13136 8560
rect 13084 8517 13093 8551
rect 13093 8517 13127 8551
rect 13127 8517 13136 8551
rect 13084 8508 13136 8517
rect 2780 8483 2832 8492
rect 2780 8449 2789 8483
rect 2789 8449 2823 8483
rect 2823 8449 2832 8483
rect 2780 8440 2832 8449
rect 4804 8440 4856 8492
rect 7196 8483 7248 8492
rect 7196 8449 7205 8483
rect 7205 8449 7239 8483
rect 7239 8449 7248 8483
rect 7196 8440 7248 8449
rect 1400 8415 1452 8424
rect 1400 8381 1409 8415
rect 1409 8381 1443 8415
rect 1443 8381 1452 8415
rect 1400 8372 1452 8381
rect 1676 8415 1728 8424
rect 1676 8381 1685 8415
rect 1685 8381 1719 8415
rect 1719 8381 1728 8415
rect 1676 8372 1728 8381
rect 4988 8372 5040 8424
rect 5172 8372 5224 8424
rect 6460 8372 6512 8424
rect 7104 8415 7156 8424
rect 7104 8381 7113 8415
rect 7113 8381 7147 8415
rect 7147 8381 7156 8415
rect 7104 8372 7156 8381
rect 8668 8440 8720 8492
rect 13268 8440 13320 8492
rect 8116 8415 8168 8424
rect 8116 8381 8125 8415
rect 8125 8381 8159 8415
rect 8159 8381 8168 8415
rect 8116 8372 8168 8381
rect 9036 8415 9088 8424
rect 5908 8304 5960 8356
rect 9036 8381 9045 8415
rect 9045 8381 9079 8415
rect 9079 8381 9088 8415
rect 9036 8372 9088 8381
rect 9680 8372 9732 8424
rect 9864 8372 9916 8424
rect 10600 8415 10652 8424
rect 10600 8381 10609 8415
rect 10609 8381 10643 8415
rect 10643 8381 10652 8415
rect 10600 8372 10652 8381
rect 11244 8372 11296 8424
rect 12072 8372 12124 8424
rect 12532 8372 12584 8424
rect 21456 8576 21508 8628
rect 23848 8576 23900 8628
rect 24400 8576 24452 8628
rect 26240 8619 26292 8628
rect 26240 8585 26249 8619
rect 26249 8585 26283 8619
rect 26283 8585 26292 8619
rect 26240 8576 26292 8585
rect 31024 8576 31076 8628
rect 14188 8508 14240 8560
rect 16212 8508 16264 8560
rect 16028 8483 16080 8492
rect 16028 8449 16037 8483
rect 16037 8449 16071 8483
rect 16071 8449 16080 8483
rect 16028 8440 16080 8449
rect 16396 8440 16448 8492
rect 16120 8415 16172 8424
rect 16120 8381 16129 8415
rect 16129 8381 16163 8415
rect 16163 8381 16172 8415
rect 16120 8372 16172 8381
rect 17132 8372 17184 8424
rect 23296 8508 23348 8560
rect 34060 8576 34112 8628
rect 38292 8576 38344 8628
rect 33232 8551 33284 8560
rect 33232 8517 33241 8551
rect 33241 8517 33275 8551
rect 33275 8517 33284 8551
rect 33232 8508 33284 8517
rect 18788 8440 18840 8492
rect 19800 8440 19852 8492
rect 21548 8440 21600 8492
rect 22192 8483 22244 8492
rect 22192 8449 22201 8483
rect 22201 8449 22235 8483
rect 22235 8449 22244 8483
rect 22192 8440 22244 8449
rect 17408 8415 17460 8424
rect 17408 8381 17417 8415
rect 17417 8381 17451 8415
rect 17451 8381 17460 8415
rect 18052 8415 18104 8424
rect 17408 8372 17460 8381
rect 18052 8381 18061 8415
rect 18061 8381 18095 8415
rect 18095 8381 18104 8415
rect 18052 8372 18104 8381
rect 15384 8304 15436 8356
rect 19064 8372 19116 8424
rect 20996 8415 21048 8424
rect 20996 8381 21005 8415
rect 21005 8381 21039 8415
rect 21039 8381 21048 8415
rect 20996 8372 21048 8381
rect 21916 8415 21968 8424
rect 21456 8304 21508 8356
rect 21916 8381 21925 8415
rect 21925 8381 21959 8415
rect 21959 8381 21968 8415
rect 21916 8372 21968 8381
rect 22468 8415 22520 8424
rect 22468 8381 22477 8415
rect 22477 8381 22511 8415
rect 22511 8381 22520 8415
rect 22468 8372 22520 8381
rect 22652 8415 22704 8424
rect 22652 8381 22661 8415
rect 22661 8381 22695 8415
rect 22695 8381 22704 8415
rect 22652 8372 22704 8381
rect 24584 8440 24636 8492
rect 24952 8483 25004 8492
rect 24952 8449 24961 8483
rect 24961 8449 24995 8483
rect 24995 8449 25004 8483
rect 24952 8440 25004 8449
rect 27988 8440 28040 8492
rect 28356 8440 28408 8492
rect 26332 8372 26384 8424
rect 27712 8372 27764 8424
rect 29092 8372 29144 8424
rect 29552 8415 29604 8424
rect 29552 8381 29561 8415
rect 29561 8381 29595 8415
rect 29595 8381 29604 8415
rect 29552 8372 29604 8381
rect 31392 8415 31444 8424
rect 31392 8381 31401 8415
rect 31401 8381 31435 8415
rect 31435 8381 31444 8415
rect 31392 8372 31444 8381
rect 31944 8372 31996 8424
rect 32220 8415 32272 8424
rect 32220 8381 32229 8415
rect 32229 8381 32263 8415
rect 32263 8381 32272 8415
rect 32220 8372 32272 8381
rect 33784 8415 33836 8424
rect 33784 8381 33793 8415
rect 33793 8381 33827 8415
rect 33827 8381 33836 8415
rect 33784 8372 33836 8381
rect 33876 8415 33928 8424
rect 33876 8381 33885 8415
rect 33885 8381 33919 8415
rect 33919 8381 33928 8415
rect 33876 8372 33928 8381
rect 34336 8372 34388 8424
rect 34520 8372 34572 8424
rect 37832 8372 37884 8424
rect 38384 8415 38436 8424
rect 38384 8381 38393 8415
rect 38393 8381 38427 8415
rect 38427 8381 38436 8415
rect 38384 8372 38436 8381
rect 4988 8236 5040 8288
rect 12532 8236 12584 8288
rect 13452 8236 13504 8288
rect 18788 8236 18840 8288
rect 34244 8304 34296 8356
rect 36820 8304 36872 8356
rect 25872 8236 25924 8288
rect 33324 8236 33376 8288
rect 19606 8134 19658 8186
rect 19670 8134 19722 8186
rect 19734 8134 19786 8186
rect 19798 8134 19850 8186
rect 8668 8075 8720 8084
rect 8668 8041 8677 8075
rect 8677 8041 8711 8075
rect 8711 8041 8720 8075
rect 8668 8032 8720 8041
rect 16672 8075 16724 8084
rect 4620 7964 4672 8016
rect 7840 7964 7892 8016
rect 15568 7964 15620 8016
rect 4160 7896 4212 7948
rect 4804 7939 4856 7948
rect 4804 7905 4813 7939
rect 4813 7905 4847 7939
rect 4847 7905 4856 7939
rect 4804 7896 4856 7905
rect 5356 7896 5408 7948
rect 5908 7896 5960 7948
rect 6092 7896 6144 7948
rect 6460 7939 6512 7948
rect 6460 7905 6469 7939
rect 6469 7905 6503 7939
rect 6503 7905 6512 7939
rect 6460 7896 6512 7905
rect 7196 7896 7248 7948
rect 10048 7896 10100 7948
rect 12072 7896 12124 7948
rect 12440 7939 12492 7948
rect 12440 7905 12449 7939
rect 12449 7905 12483 7939
rect 12483 7905 12492 7939
rect 12440 7896 12492 7905
rect 12992 7896 13044 7948
rect 14188 7939 14240 7948
rect 14188 7905 14197 7939
rect 14197 7905 14231 7939
rect 14231 7905 14240 7939
rect 14188 7896 14240 7905
rect 15476 7939 15528 7948
rect 15476 7905 15485 7939
rect 15485 7905 15519 7939
rect 15519 7905 15528 7939
rect 15476 7896 15528 7905
rect 16672 8041 16681 8075
rect 16681 8041 16715 8075
rect 16715 8041 16724 8075
rect 16672 8032 16724 8041
rect 16948 8032 17000 8084
rect 18880 8032 18932 8084
rect 22008 8032 22060 8084
rect 25872 8075 25924 8084
rect 16120 7964 16172 8016
rect 15936 7896 15988 7948
rect 19156 7964 19208 8016
rect 24768 7964 24820 8016
rect 25872 8041 25881 8075
rect 25881 8041 25915 8075
rect 25915 8041 25924 8075
rect 25872 8032 25924 8041
rect 27528 8032 27580 8084
rect 27712 8075 27764 8084
rect 27712 8041 27721 8075
rect 27721 8041 27755 8075
rect 27755 8041 27764 8075
rect 27712 8032 27764 8041
rect 29368 8075 29420 8084
rect 29368 8041 29377 8075
rect 29377 8041 29411 8075
rect 29411 8041 29420 8075
rect 29368 8032 29420 8041
rect 31300 8075 31352 8084
rect 31300 8041 31309 8075
rect 31309 8041 31343 8075
rect 31343 8041 31352 8075
rect 31300 8032 31352 8041
rect 33876 8032 33928 8084
rect 1400 7871 1452 7880
rect 1400 7837 1409 7871
rect 1409 7837 1443 7871
rect 1443 7837 1452 7871
rect 1400 7828 1452 7837
rect 2504 7828 2556 7880
rect 9956 7871 10008 7880
rect 9956 7837 9965 7871
rect 9965 7837 9999 7871
rect 9999 7837 10008 7871
rect 9956 7828 10008 7837
rect 3516 7760 3568 7812
rect 2964 7735 3016 7744
rect 2964 7701 2973 7735
rect 2973 7701 3007 7735
rect 3007 7701 3016 7735
rect 2964 7692 3016 7701
rect 4988 7692 5040 7744
rect 15292 7828 15344 7880
rect 15384 7828 15436 7880
rect 16488 7828 16540 7880
rect 17224 7896 17276 7948
rect 17500 7896 17552 7948
rect 18788 7939 18840 7948
rect 18788 7905 18797 7939
rect 18797 7905 18831 7939
rect 18831 7905 18840 7939
rect 18788 7896 18840 7905
rect 18880 7896 18932 7948
rect 19800 7896 19852 7948
rect 19984 7939 20036 7948
rect 19984 7905 19993 7939
rect 19993 7905 20027 7939
rect 20027 7905 20036 7939
rect 19984 7896 20036 7905
rect 22100 7896 22152 7948
rect 23296 7939 23348 7948
rect 23296 7905 23305 7939
rect 23305 7905 23339 7939
rect 23339 7905 23348 7939
rect 23296 7896 23348 7905
rect 24032 7896 24084 7948
rect 24676 7896 24728 7948
rect 25412 7896 25464 7948
rect 11060 7760 11112 7812
rect 11980 7760 12032 7812
rect 21272 7828 21324 7880
rect 21456 7828 21508 7880
rect 27068 7896 27120 7948
rect 34336 7964 34388 8016
rect 34428 7964 34480 8016
rect 27436 7896 27488 7948
rect 28356 7939 28408 7948
rect 28356 7905 28365 7939
rect 28365 7905 28399 7939
rect 28399 7905 28408 7939
rect 28356 7896 28408 7905
rect 29276 7939 29328 7948
rect 29276 7905 29285 7939
rect 29285 7905 29319 7939
rect 29319 7905 29328 7939
rect 29276 7896 29328 7905
rect 33508 7896 33560 7948
rect 35348 7896 35400 7948
rect 11520 7692 11572 7744
rect 17040 7735 17092 7744
rect 17040 7701 17049 7735
rect 17049 7701 17083 7735
rect 17083 7701 17092 7735
rect 17040 7692 17092 7701
rect 17592 7692 17644 7744
rect 17868 7692 17920 7744
rect 19064 7692 19116 7744
rect 19248 7760 19300 7812
rect 23388 7803 23440 7812
rect 23388 7769 23397 7803
rect 23397 7769 23431 7803
rect 23431 7769 23440 7803
rect 23388 7760 23440 7769
rect 29092 7828 29144 7880
rect 30564 7828 30616 7880
rect 32404 7871 32456 7880
rect 32404 7837 32413 7871
rect 32413 7837 32447 7871
rect 32447 7837 32456 7871
rect 32404 7828 32456 7837
rect 33692 7828 33744 7880
rect 34796 7871 34848 7880
rect 34796 7837 34805 7871
rect 34805 7837 34839 7871
rect 34839 7837 34848 7871
rect 34796 7828 34848 7837
rect 36084 7828 36136 7880
rect 28172 7760 28224 7812
rect 21824 7692 21876 7744
rect 22468 7692 22520 7744
rect 25320 7692 25372 7744
rect 29460 7692 29512 7744
rect 36268 7692 36320 7744
rect 4246 7590 4298 7642
rect 4310 7590 4362 7642
rect 4374 7590 4426 7642
rect 4438 7590 4490 7642
rect 34966 7590 35018 7642
rect 35030 7590 35082 7642
rect 35094 7590 35146 7642
rect 35158 7590 35210 7642
rect 2320 7327 2372 7336
rect 2320 7293 2329 7327
rect 2329 7293 2363 7327
rect 2363 7293 2372 7327
rect 2320 7284 2372 7293
rect 4896 7488 4948 7540
rect 6092 7488 6144 7540
rect 6552 7488 6604 7540
rect 7104 7488 7156 7540
rect 4620 7420 4672 7472
rect 7840 7463 7892 7472
rect 7840 7429 7849 7463
rect 7849 7429 7883 7463
rect 7883 7429 7892 7463
rect 7840 7420 7892 7429
rect 3516 7395 3568 7404
rect 3516 7361 3525 7395
rect 3525 7361 3559 7395
rect 3559 7361 3568 7395
rect 3516 7352 3568 7361
rect 4988 7352 5040 7404
rect 5172 7284 5224 7336
rect 5264 7284 5316 7336
rect 7472 7284 7524 7336
rect 8300 7284 8352 7336
rect 8392 7327 8444 7336
rect 8392 7293 8401 7327
rect 8401 7293 8435 7327
rect 8435 7293 8444 7327
rect 11244 7488 11296 7540
rect 15936 7488 15988 7540
rect 16488 7488 16540 7540
rect 14188 7463 14240 7472
rect 14188 7429 14197 7463
rect 14197 7429 14231 7463
rect 14231 7429 14240 7463
rect 14188 7420 14240 7429
rect 9956 7395 10008 7404
rect 9956 7361 9965 7395
rect 9965 7361 9999 7395
rect 9999 7361 10008 7395
rect 9956 7352 10008 7361
rect 8392 7284 8444 7293
rect 9864 7327 9916 7336
rect 9864 7293 9873 7327
rect 9873 7293 9907 7327
rect 9907 7293 9916 7327
rect 11980 7352 12032 7404
rect 12072 7352 12124 7404
rect 9864 7284 9916 7293
rect 10784 7327 10836 7336
rect 10784 7293 10793 7327
rect 10793 7293 10827 7327
rect 10827 7293 10836 7327
rect 10784 7284 10836 7293
rect 11520 7327 11572 7336
rect 11520 7293 11529 7327
rect 11529 7293 11563 7327
rect 11563 7293 11572 7327
rect 11520 7284 11572 7293
rect 13728 7352 13780 7404
rect 10600 7216 10652 7268
rect 13820 7284 13872 7336
rect 14004 7327 14056 7336
rect 14004 7293 14013 7327
rect 14013 7293 14047 7327
rect 14047 7293 14056 7327
rect 14004 7284 14056 7293
rect 18144 7352 18196 7404
rect 14280 7216 14332 7268
rect 1676 7148 1728 7200
rect 16856 7284 16908 7336
rect 24768 7488 24820 7540
rect 25320 7488 25372 7540
rect 33416 7488 33468 7540
rect 22376 7463 22428 7472
rect 18880 7352 18932 7404
rect 19248 7395 19300 7404
rect 19248 7361 19257 7395
rect 19257 7361 19291 7395
rect 19291 7361 19300 7395
rect 19248 7352 19300 7361
rect 19064 7284 19116 7336
rect 21548 7327 21600 7336
rect 21548 7293 21557 7327
rect 21557 7293 21591 7327
rect 21591 7293 21600 7327
rect 21548 7284 21600 7293
rect 21824 7284 21876 7336
rect 22376 7429 22385 7463
rect 22385 7429 22419 7463
rect 22419 7429 22428 7463
rect 22376 7420 22428 7429
rect 23848 7420 23900 7472
rect 24860 7420 24912 7472
rect 28172 7420 28224 7472
rect 30840 7420 30892 7472
rect 22468 7327 22520 7336
rect 22468 7293 22477 7327
rect 22477 7293 22511 7327
rect 22511 7293 22520 7327
rect 22468 7284 22520 7293
rect 20260 7216 20312 7268
rect 29552 7352 29604 7404
rect 31024 7352 31076 7404
rect 31576 7395 31628 7404
rect 31576 7361 31585 7395
rect 31585 7361 31619 7395
rect 31619 7361 31628 7395
rect 31576 7352 31628 7361
rect 23848 7327 23900 7336
rect 23848 7293 23857 7327
rect 23857 7293 23891 7327
rect 23891 7293 23900 7327
rect 23848 7284 23900 7293
rect 24032 7327 24084 7336
rect 24032 7293 24041 7327
rect 24041 7293 24075 7327
rect 24075 7293 24084 7327
rect 24032 7284 24084 7293
rect 24400 7327 24452 7336
rect 24400 7293 24409 7327
rect 24409 7293 24443 7327
rect 24443 7293 24452 7327
rect 24400 7284 24452 7293
rect 25228 7284 25280 7336
rect 25780 7327 25832 7336
rect 25780 7293 25789 7327
rect 25789 7293 25823 7327
rect 25823 7293 25832 7327
rect 25780 7284 25832 7293
rect 26332 7327 26384 7336
rect 26332 7293 26341 7327
rect 26341 7293 26375 7327
rect 26375 7293 26384 7327
rect 26332 7284 26384 7293
rect 27804 7284 27856 7336
rect 29000 7284 29052 7336
rect 31852 7327 31904 7336
rect 16672 7148 16724 7200
rect 17224 7148 17276 7200
rect 19248 7148 19300 7200
rect 21732 7148 21784 7200
rect 22008 7148 22060 7200
rect 22652 7148 22704 7200
rect 23940 7148 23992 7200
rect 29552 7216 29604 7268
rect 31852 7293 31861 7327
rect 31861 7293 31895 7327
rect 31895 7293 31904 7327
rect 31852 7284 31904 7293
rect 32036 7327 32088 7336
rect 32036 7293 32045 7327
rect 32045 7293 32079 7327
rect 32079 7293 32088 7327
rect 32036 7284 32088 7293
rect 35440 7352 35492 7404
rect 36728 7395 36780 7404
rect 36728 7361 36737 7395
rect 36737 7361 36771 7395
rect 36771 7361 36780 7395
rect 36728 7352 36780 7361
rect 37372 7395 37424 7404
rect 37372 7361 37381 7395
rect 37381 7361 37415 7395
rect 37415 7361 37424 7395
rect 37372 7352 37424 7361
rect 37648 7395 37700 7404
rect 37648 7361 37657 7395
rect 37657 7361 37691 7395
rect 37691 7361 37700 7395
rect 37648 7352 37700 7361
rect 33324 7327 33376 7336
rect 30288 7216 30340 7268
rect 31116 7216 31168 7268
rect 32772 7216 32824 7268
rect 27988 7148 28040 7200
rect 30932 7148 30984 7200
rect 31576 7148 31628 7200
rect 32680 7148 32732 7200
rect 33324 7293 33333 7327
rect 33333 7293 33367 7327
rect 33367 7293 33376 7327
rect 33324 7284 33376 7293
rect 35072 7327 35124 7336
rect 35072 7293 35081 7327
rect 35081 7293 35115 7327
rect 35115 7293 35124 7327
rect 35072 7284 35124 7293
rect 33600 7148 33652 7200
rect 19606 7046 19658 7098
rect 19670 7046 19722 7098
rect 19734 7046 19786 7098
rect 19798 7046 19850 7098
rect 8300 6944 8352 6996
rect 10324 6944 10376 6996
rect 20260 6944 20312 6996
rect 22652 6944 22704 6996
rect 24676 6944 24728 6996
rect 29460 6944 29512 6996
rect 29552 6944 29604 6996
rect 35072 6944 35124 6996
rect 4988 6876 5040 6928
rect 2780 6808 2832 6860
rect 2872 6740 2924 6792
rect 4620 6808 4672 6860
rect 15292 6876 15344 6928
rect 15660 6876 15712 6928
rect 16856 6919 16908 6928
rect 16856 6885 16865 6919
rect 16865 6885 16899 6919
rect 16899 6885 16908 6919
rect 16856 6876 16908 6885
rect 17500 6876 17552 6928
rect 18420 6919 18472 6928
rect 6276 6851 6328 6860
rect 6276 6817 6285 6851
rect 6285 6817 6319 6851
rect 6319 6817 6328 6851
rect 6276 6808 6328 6817
rect 6552 6851 6604 6860
rect 6552 6817 6561 6851
rect 6561 6817 6595 6851
rect 6595 6817 6604 6851
rect 6552 6808 6604 6817
rect 10508 6808 10560 6860
rect 11060 6851 11112 6860
rect 11060 6817 11069 6851
rect 11069 6817 11103 6851
rect 11103 6817 11112 6851
rect 11060 6808 11112 6817
rect 12440 6808 12492 6860
rect 13544 6808 13596 6860
rect 4896 6672 4948 6724
rect 6184 6740 6236 6792
rect 6828 6740 6880 6792
rect 7472 6740 7524 6792
rect 11152 6783 11204 6792
rect 7012 6672 7064 6724
rect 11152 6749 11161 6783
rect 11161 6749 11195 6783
rect 11195 6749 11204 6783
rect 11152 6740 11204 6749
rect 12072 6783 12124 6792
rect 12072 6749 12081 6783
rect 12081 6749 12115 6783
rect 12115 6749 12124 6783
rect 12072 6740 12124 6749
rect 16580 6808 16632 6860
rect 17040 6808 17092 6860
rect 17132 6808 17184 6860
rect 17592 6851 17644 6860
rect 17592 6817 17601 6851
rect 17601 6817 17635 6851
rect 17635 6817 17644 6851
rect 17592 6808 17644 6817
rect 18420 6885 18429 6919
rect 18429 6885 18463 6919
rect 18463 6885 18472 6919
rect 18420 6876 18472 6885
rect 19432 6876 19484 6928
rect 21088 6876 21140 6928
rect 11796 6672 11848 6724
rect 13636 6672 13688 6724
rect 2504 6647 2556 6656
rect 2504 6613 2513 6647
rect 2513 6613 2547 6647
rect 2547 6613 2556 6647
rect 2504 6604 2556 6613
rect 4620 6604 4672 6656
rect 7564 6604 7616 6656
rect 13360 6604 13412 6656
rect 14188 6604 14240 6656
rect 16764 6740 16816 6792
rect 17224 6740 17276 6792
rect 18144 6808 18196 6860
rect 19248 6808 19300 6860
rect 19892 6808 19944 6860
rect 19984 6783 20036 6792
rect 19984 6749 19993 6783
rect 19993 6749 20027 6783
rect 20027 6749 20036 6783
rect 19984 6740 20036 6749
rect 20168 6808 20220 6860
rect 20628 6808 20680 6860
rect 21916 6851 21968 6860
rect 20260 6740 20312 6792
rect 21456 6783 21508 6792
rect 21456 6749 21465 6783
rect 21465 6749 21499 6783
rect 21499 6749 21508 6783
rect 21456 6740 21508 6749
rect 21916 6817 21925 6851
rect 21925 6817 21959 6851
rect 21959 6817 21968 6851
rect 21916 6808 21968 6817
rect 22008 6808 22060 6860
rect 23112 6851 23164 6860
rect 23112 6817 23121 6851
rect 23121 6817 23155 6851
rect 23155 6817 23164 6851
rect 23112 6808 23164 6817
rect 25780 6876 25832 6928
rect 29000 6919 29052 6928
rect 29000 6885 29009 6919
rect 29009 6885 29043 6919
rect 29043 6885 29052 6919
rect 29000 6876 29052 6885
rect 24676 6808 24728 6860
rect 25136 6851 25188 6860
rect 22560 6740 22612 6792
rect 15844 6672 15896 6724
rect 20352 6604 20404 6656
rect 21916 6604 21968 6656
rect 22192 6604 22244 6656
rect 25136 6817 25145 6851
rect 25145 6817 25179 6851
rect 25179 6817 25188 6851
rect 25136 6808 25188 6817
rect 26332 6808 26384 6860
rect 24952 6783 25004 6792
rect 24952 6749 24961 6783
rect 24961 6749 24995 6783
rect 24995 6749 25004 6783
rect 24952 6740 25004 6749
rect 25872 6740 25924 6792
rect 28172 6808 28224 6860
rect 29828 6851 29880 6860
rect 27620 6740 27672 6792
rect 28632 6740 28684 6792
rect 29828 6817 29837 6851
rect 29837 6817 29871 6851
rect 29871 6817 29880 6851
rect 29828 6808 29880 6817
rect 30564 6851 30616 6860
rect 30564 6817 30573 6851
rect 30573 6817 30607 6851
rect 30607 6817 30616 6851
rect 30564 6808 30616 6817
rect 31116 6851 31168 6860
rect 31116 6817 31125 6851
rect 31125 6817 31159 6851
rect 31159 6817 31168 6851
rect 31116 6808 31168 6817
rect 29920 6740 29972 6792
rect 32036 6808 32088 6860
rect 33692 6851 33744 6860
rect 31760 6740 31812 6792
rect 33416 6783 33468 6792
rect 33416 6749 33425 6783
rect 33425 6749 33459 6783
rect 33459 6749 33468 6783
rect 33416 6740 33468 6749
rect 33692 6817 33701 6851
rect 33701 6817 33735 6851
rect 33735 6817 33744 6851
rect 33692 6808 33744 6817
rect 36912 6808 36964 6860
rect 33600 6740 33652 6792
rect 34428 6740 34480 6792
rect 26056 6604 26108 6656
rect 26332 6604 26384 6656
rect 27528 6604 27580 6656
rect 31484 6604 31536 6656
rect 34704 6604 34756 6656
rect 36912 6647 36964 6656
rect 36912 6613 36921 6647
rect 36921 6613 36955 6647
rect 36955 6613 36964 6647
rect 36912 6604 36964 6613
rect 4246 6502 4298 6554
rect 4310 6502 4362 6554
rect 4374 6502 4426 6554
rect 4438 6502 4490 6554
rect 34966 6502 35018 6554
rect 35030 6502 35082 6554
rect 35094 6502 35146 6554
rect 35158 6502 35210 6554
rect 8116 6400 8168 6452
rect 9864 6443 9916 6452
rect 9864 6409 9873 6443
rect 9873 6409 9907 6443
rect 9907 6409 9916 6443
rect 9864 6400 9916 6409
rect 4712 6332 4764 6384
rect 6276 6332 6328 6384
rect 4344 6307 4396 6316
rect 4344 6273 4353 6307
rect 4353 6273 4387 6307
rect 4387 6273 4396 6307
rect 4344 6264 4396 6273
rect 4988 6196 5040 6248
rect 5540 6196 5592 6248
rect 6552 6264 6604 6316
rect 7472 6307 7524 6316
rect 7472 6273 7481 6307
rect 7481 6273 7515 6307
rect 7515 6273 7524 6307
rect 7472 6264 7524 6273
rect 6092 6239 6144 6248
rect 6092 6205 6101 6239
rect 6101 6205 6135 6239
rect 6135 6205 6144 6239
rect 6092 6196 6144 6205
rect 7104 6239 7156 6248
rect 7104 6205 7113 6239
rect 7113 6205 7147 6239
rect 7147 6205 7156 6239
rect 7104 6196 7156 6205
rect 7840 6196 7892 6248
rect 8116 6239 8168 6248
rect 8116 6205 8125 6239
rect 8125 6205 8159 6239
rect 8159 6205 8168 6239
rect 8116 6196 8168 6205
rect 9680 6332 9732 6384
rect 10784 6332 10836 6384
rect 12072 6332 12124 6384
rect 8300 6239 8352 6248
rect 8300 6205 8309 6239
rect 8309 6205 8343 6239
rect 8343 6205 8352 6239
rect 8300 6196 8352 6205
rect 9864 6196 9916 6248
rect 4620 6128 4672 6180
rect 6184 6171 6236 6180
rect 6184 6137 6193 6171
rect 6193 6137 6227 6171
rect 6227 6137 6236 6171
rect 10600 6196 10652 6248
rect 11152 6239 11204 6248
rect 11152 6205 11161 6239
rect 11161 6205 11195 6239
rect 11195 6205 11204 6239
rect 11152 6196 11204 6205
rect 6184 6128 6236 6137
rect 10876 6128 10928 6180
rect 13176 6196 13228 6248
rect 11704 6171 11756 6180
rect 11704 6137 11713 6171
rect 11713 6137 11747 6171
rect 11747 6137 11756 6171
rect 11704 6128 11756 6137
rect 13360 6239 13412 6248
rect 13360 6205 13369 6239
rect 13369 6205 13403 6239
rect 13403 6205 13412 6239
rect 14004 6239 14056 6248
rect 13360 6196 13412 6205
rect 14004 6205 14013 6239
rect 14013 6205 14047 6239
rect 14047 6205 14056 6239
rect 14004 6196 14056 6205
rect 14096 6196 14148 6248
rect 15476 6196 15528 6248
rect 15752 6307 15804 6316
rect 15752 6273 15761 6307
rect 15761 6273 15795 6307
rect 15795 6273 15804 6307
rect 15752 6264 15804 6273
rect 14188 6128 14240 6180
rect 16120 6332 16172 6384
rect 19432 6332 19484 6384
rect 20628 6400 20680 6452
rect 20812 6332 20864 6384
rect 16396 6264 16448 6316
rect 24308 6400 24360 6452
rect 26056 6443 26108 6452
rect 26056 6409 26065 6443
rect 26065 6409 26099 6443
rect 26099 6409 26108 6443
rect 26056 6400 26108 6409
rect 27528 6400 27580 6452
rect 28172 6443 28224 6452
rect 28172 6409 28181 6443
rect 28181 6409 28215 6443
rect 28215 6409 28224 6443
rect 28172 6400 28224 6409
rect 29460 6443 29512 6452
rect 29460 6409 29469 6443
rect 29469 6409 29503 6443
rect 29503 6409 29512 6443
rect 29460 6400 29512 6409
rect 29920 6400 29972 6452
rect 34612 6400 34664 6452
rect 16580 6239 16632 6248
rect 16580 6205 16589 6239
rect 16589 6205 16623 6239
rect 16623 6205 16632 6239
rect 16580 6196 16632 6205
rect 16672 6196 16724 6248
rect 18420 6196 18472 6248
rect 19064 6196 19116 6248
rect 19156 6196 19208 6248
rect 8300 6060 8352 6112
rect 17960 6128 18012 6180
rect 20720 6196 20772 6248
rect 20812 6196 20864 6248
rect 34888 6332 34940 6384
rect 37096 6332 37148 6384
rect 22100 6264 22152 6316
rect 22468 6307 22520 6316
rect 21640 6196 21692 6248
rect 22468 6273 22477 6307
rect 22477 6273 22511 6307
rect 22511 6273 22520 6307
rect 22468 6264 22520 6273
rect 23940 6239 23992 6248
rect 23940 6205 23949 6239
rect 23949 6205 23983 6239
rect 23983 6205 23992 6239
rect 23940 6196 23992 6205
rect 24032 6239 24084 6248
rect 24032 6205 24041 6239
rect 24041 6205 24075 6239
rect 24075 6205 24084 6239
rect 24676 6239 24728 6248
rect 24032 6196 24084 6205
rect 24676 6205 24685 6239
rect 24685 6205 24719 6239
rect 24719 6205 24728 6239
rect 24676 6196 24728 6205
rect 26424 6264 26476 6316
rect 26976 6264 27028 6316
rect 27896 6264 27948 6316
rect 30104 6264 30156 6316
rect 30932 6264 30984 6316
rect 31484 6307 31536 6316
rect 31484 6273 31493 6307
rect 31493 6273 31527 6307
rect 31527 6273 31536 6307
rect 31484 6264 31536 6273
rect 32404 6264 32456 6316
rect 32772 6307 32824 6316
rect 32772 6273 32781 6307
rect 32781 6273 32815 6307
rect 32815 6273 32824 6307
rect 32772 6264 32824 6273
rect 26884 6239 26936 6248
rect 22468 6128 22520 6180
rect 17776 6060 17828 6112
rect 19064 6103 19116 6112
rect 19064 6069 19073 6103
rect 19073 6069 19107 6103
rect 19107 6069 19116 6103
rect 19064 6060 19116 6069
rect 26884 6205 26893 6239
rect 26893 6205 26927 6239
rect 26927 6205 26936 6239
rect 26884 6196 26936 6205
rect 29276 6239 29328 6248
rect 29276 6205 29285 6239
rect 29285 6205 29319 6239
rect 29319 6205 29328 6239
rect 29276 6196 29328 6205
rect 31944 6196 31996 6248
rect 36084 6264 36136 6316
rect 30932 6128 30984 6180
rect 31760 6128 31812 6180
rect 33600 6196 33652 6248
rect 29092 6060 29144 6112
rect 33508 6060 33560 6112
rect 34428 6060 34480 6112
rect 37096 6196 37148 6248
rect 36728 6128 36780 6180
rect 19606 5958 19658 6010
rect 19670 5958 19722 6010
rect 19734 5958 19786 6010
rect 19798 5958 19850 6010
rect 5540 5856 5592 5908
rect 11520 5856 11572 5908
rect 12164 5856 12216 5908
rect 8208 5788 8260 5840
rect 8392 5788 8444 5840
rect 4344 5763 4396 5772
rect 4344 5729 4353 5763
rect 4353 5729 4387 5763
rect 4387 5729 4396 5763
rect 4344 5720 4396 5729
rect 6920 5720 6972 5772
rect 7104 5720 7156 5772
rect 8116 5763 8168 5772
rect 4068 5695 4120 5704
rect 4068 5661 4077 5695
rect 4077 5661 4111 5695
rect 4111 5661 4120 5695
rect 4068 5652 4120 5661
rect 6552 5652 6604 5704
rect 8116 5729 8125 5763
rect 8125 5729 8159 5763
rect 8159 5729 8168 5763
rect 8116 5720 8168 5729
rect 8760 5720 8812 5772
rect 9588 5720 9640 5772
rect 9772 5720 9824 5772
rect 7012 5584 7064 5636
rect 7288 5627 7340 5636
rect 7288 5593 7297 5627
rect 7297 5593 7331 5627
rect 7331 5593 7340 5627
rect 7288 5584 7340 5593
rect 10140 5516 10192 5568
rect 11060 5720 11112 5772
rect 11520 5763 11572 5772
rect 10508 5695 10560 5704
rect 10508 5661 10517 5695
rect 10517 5661 10551 5695
rect 10551 5661 10560 5695
rect 10508 5652 10560 5661
rect 10416 5584 10468 5636
rect 11520 5729 11529 5763
rect 11529 5729 11563 5763
rect 11563 5729 11572 5763
rect 11520 5720 11572 5729
rect 12256 5763 12308 5772
rect 12256 5729 12265 5763
rect 12265 5729 12299 5763
rect 12299 5729 12308 5763
rect 12256 5720 12308 5729
rect 13820 5856 13872 5908
rect 14280 5899 14332 5908
rect 14280 5865 14289 5899
rect 14289 5865 14323 5899
rect 14323 5865 14332 5899
rect 14280 5856 14332 5865
rect 13728 5788 13780 5840
rect 13544 5763 13596 5772
rect 13544 5729 13553 5763
rect 13553 5729 13587 5763
rect 13587 5729 13596 5763
rect 13544 5720 13596 5729
rect 13820 5720 13872 5772
rect 16120 5856 16172 5908
rect 17592 5856 17644 5908
rect 20260 5856 20312 5908
rect 21640 5856 21692 5908
rect 25872 5856 25924 5908
rect 14556 5720 14608 5772
rect 17776 5788 17828 5840
rect 15200 5720 15252 5772
rect 15936 5763 15988 5772
rect 15936 5729 15945 5763
rect 15945 5729 15979 5763
rect 15979 5729 15988 5763
rect 15936 5720 15988 5729
rect 16028 5763 16080 5772
rect 16028 5729 16037 5763
rect 16037 5729 16071 5763
rect 16071 5729 16080 5763
rect 16028 5720 16080 5729
rect 13636 5584 13688 5636
rect 14740 5584 14792 5636
rect 16580 5720 16632 5772
rect 17960 5763 18012 5772
rect 17960 5729 17969 5763
rect 17969 5729 18003 5763
rect 18003 5729 18012 5763
rect 17960 5720 18012 5729
rect 21732 5763 21784 5772
rect 21732 5729 21741 5763
rect 21741 5729 21775 5763
rect 21775 5729 21784 5763
rect 21732 5720 21784 5729
rect 16948 5584 17000 5636
rect 12808 5516 12860 5568
rect 13452 5516 13504 5568
rect 13544 5516 13596 5568
rect 15936 5516 15988 5568
rect 17592 5516 17644 5568
rect 21640 5652 21692 5704
rect 21824 5695 21876 5704
rect 21824 5661 21833 5695
rect 21833 5661 21867 5695
rect 21867 5661 21876 5695
rect 21824 5652 21876 5661
rect 26884 5788 26936 5840
rect 22376 5720 22428 5772
rect 24216 5720 24268 5772
rect 25136 5763 25188 5772
rect 24124 5652 24176 5704
rect 24860 5627 24912 5636
rect 24860 5593 24869 5627
rect 24869 5593 24903 5627
rect 24903 5593 24912 5627
rect 24860 5584 24912 5593
rect 17960 5516 18012 5568
rect 19064 5516 19116 5568
rect 19984 5516 20036 5568
rect 21640 5516 21692 5568
rect 25136 5729 25145 5763
rect 25145 5729 25179 5763
rect 25179 5729 25188 5763
rect 25136 5720 25188 5729
rect 26332 5720 26384 5772
rect 27620 5763 27672 5772
rect 27620 5729 27629 5763
rect 27629 5729 27663 5763
rect 27663 5729 27672 5763
rect 27620 5720 27672 5729
rect 27896 5763 27948 5772
rect 27896 5729 27905 5763
rect 27905 5729 27939 5763
rect 27939 5729 27948 5763
rect 27896 5720 27948 5729
rect 28172 5856 28224 5908
rect 29920 5856 29972 5908
rect 31024 5856 31076 5908
rect 28632 5788 28684 5840
rect 35348 5856 35400 5908
rect 36728 5856 36780 5908
rect 29276 5720 29328 5772
rect 29920 5763 29972 5772
rect 29920 5729 29929 5763
rect 29929 5729 29963 5763
rect 29963 5729 29972 5763
rect 29920 5720 29972 5729
rect 30104 5720 30156 5772
rect 34796 5788 34848 5840
rect 31760 5720 31812 5772
rect 32680 5763 32732 5772
rect 32680 5729 32689 5763
rect 32689 5729 32723 5763
rect 32723 5729 32732 5763
rect 32680 5720 32732 5729
rect 29368 5695 29420 5704
rect 29368 5661 29377 5695
rect 29377 5661 29411 5695
rect 29411 5661 29420 5695
rect 29368 5652 29420 5661
rect 32588 5652 32640 5704
rect 29000 5584 29052 5636
rect 28908 5516 28960 5568
rect 33232 5720 33284 5772
rect 33600 5720 33652 5772
rect 34520 5763 34572 5772
rect 34520 5729 34529 5763
rect 34529 5729 34563 5763
rect 34563 5729 34572 5763
rect 34520 5720 34572 5729
rect 34704 5763 34756 5772
rect 34704 5729 34713 5763
rect 34713 5729 34747 5763
rect 34747 5729 34756 5763
rect 34704 5720 34756 5729
rect 34888 5720 34940 5772
rect 35624 5720 35676 5772
rect 36544 5720 36596 5772
rect 36912 5720 36964 5772
rect 33692 5695 33744 5704
rect 33692 5661 33701 5695
rect 33701 5661 33735 5695
rect 33735 5661 33744 5695
rect 33692 5652 33744 5661
rect 34612 5652 34664 5704
rect 4246 5414 4298 5466
rect 4310 5414 4362 5466
rect 4374 5414 4426 5466
rect 4438 5414 4490 5466
rect 34966 5414 35018 5466
rect 35030 5414 35082 5466
rect 35094 5414 35146 5466
rect 35158 5414 35210 5466
rect 6092 5312 6144 5364
rect 9772 5312 9824 5364
rect 11060 5312 11112 5364
rect 11520 5312 11572 5364
rect 13452 5312 13504 5364
rect 13728 5312 13780 5364
rect 17592 5312 17644 5364
rect 26424 5355 26476 5364
rect 12256 5244 12308 5296
rect 4068 5176 4120 5228
rect 4896 5219 4948 5228
rect 2320 5108 2372 5160
rect 4528 5108 4580 5160
rect 4896 5185 4905 5219
rect 4905 5185 4939 5219
rect 4939 5185 4948 5219
rect 4896 5176 4948 5185
rect 7288 5219 7340 5228
rect 7288 5185 7297 5219
rect 7297 5185 7331 5219
rect 7331 5185 7340 5219
rect 7288 5176 7340 5185
rect 8484 5176 8536 5228
rect 9864 5176 9916 5228
rect 6828 5108 6880 5160
rect 8116 5108 8168 5160
rect 8392 5108 8444 5160
rect 9680 5151 9732 5160
rect 9680 5117 9689 5151
rect 9689 5117 9723 5151
rect 9723 5117 9732 5151
rect 10416 5176 10468 5228
rect 10600 5176 10652 5228
rect 12716 5219 12768 5228
rect 9680 5108 9732 5117
rect 10324 5151 10376 5160
rect 10324 5117 10333 5151
rect 10333 5117 10367 5151
rect 10367 5117 10376 5151
rect 10324 5108 10376 5117
rect 12716 5185 12725 5219
rect 12725 5185 12759 5219
rect 12759 5185 12768 5219
rect 12716 5176 12768 5185
rect 11428 5108 11480 5160
rect 12808 5151 12860 5160
rect 12808 5117 12817 5151
rect 12817 5117 12851 5151
rect 12851 5117 12860 5151
rect 12808 5108 12860 5117
rect 13636 5151 13688 5160
rect 4068 5083 4120 5092
rect 4068 5049 4077 5083
rect 4077 5049 4111 5083
rect 4111 5049 4120 5083
rect 4068 5040 4120 5049
rect 13636 5117 13645 5151
rect 13645 5117 13679 5151
rect 13679 5117 13688 5151
rect 13636 5108 13688 5117
rect 14004 5151 14056 5160
rect 14004 5117 14013 5151
rect 14013 5117 14047 5151
rect 14047 5117 14056 5151
rect 14004 5108 14056 5117
rect 16396 5244 16448 5296
rect 16212 5219 16264 5228
rect 16212 5185 16221 5219
rect 16221 5185 16255 5219
rect 16255 5185 16264 5219
rect 16212 5176 16264 5185
rect 16304 5176 16356 5228
rect 26424 5321 26433 5355
rect 26433 5321 26467 5355
rect 26467 5321 26476 5355
rect 26424 5312 26476 5321
rect 33232 5312 33284 5364
rect 36728 5312 36780 5364
rect 15200 5108 15252 5160
rect 15660 5108 15712 5160
rect 16028 5151 16080 5160
rect 13452 5040 13504 5092
rect 16028 5117 16037 5151
rect 16037 5117 16071 5151
rect 16071 5117 16080 5151
rect 16028 5108 16080 5117
rect 16488 5040 16540 5092
rect 16764 5108 16816 5160
rect 17776 5108 17828 5160
rect 18696 5151 18748 5160
rect 18696 5117 18705 5151
rect 18705 5117 18739 5151
rect 18739 5117 18748 5151
rect 18696 5108 18748 5117
rect 21732 5176 21784 5228
rect 28172 5219 28224 5228
rect 28172 5185 28181 5219
rect 28181 5185 28215 5219
rect 28215 5185 28224 5219
rect 28172 5176 28224 5185
rect 28632 5219 28684 5228
rect 28632 5185 28641 5219
rect 28641 5185 28675 5219
rect 28675 5185 28684 5219
rect 28632 5176 28684 5185
rect 16856 5040 16908 5092
rect 18052 4972 18104 5024
rect 22100 5151 22152 5160
rect 22100 5117 22109 5151
rect 22109 5117 22143 5151
rect 22143 5117 22152 5151
rect 22100 5108 22152 5117
rect 23940 5108 23992 5160
rect 24308 5108 24360 5160
rect 24860 5151 24912 5160
rect 24860 5117 24869 5151
rect 24869 5117 24903 5151
rect 24903 5117 24912 5151
rect 24860 5108 24912 5117
rect 27528 5108 27580 5160
rect 28264 5108 28316 5160
rect 29092 5108 29144 5160
rect 37096 5176 37148 5228
rect 29552 5151 29604 5160
rect 29552 5117 29561 5151
rect 29561 5117 29595 5151
rect 29595 5117 29604 5151
rect 29552 5108 29604 5117
rect 32128 5108 32180 5160
rect 34520 5108 34572 5160
rect 35624 5151 35676 5160
rect 35624 5117 35633 5151
rect 35633 5117 35667 5151
rect 35667 5117 35676 5151
rect 35624 5108 35676 5117
rect 36084 5151 36136 5160
rect 22192 5040 22244 5092
rect 22836 5040 22888 5092
rect 27620 5083 27672 5092
rect 27620 5049 27629 5083
rect 27629 5049 27663 5083
rect 27663 5049 27672 5083
rect 27620 5040 27672 5049
rect 24216 5015 24268 5024
rect 24216 4981 24225 5015
rect 24225 4981 24259 5015
rect 24259 4981 24268 5015
rect 36084 5117 36093 5151
rect 36093 5117 36127 5151
rect 36127 5117 36136 5151
rect 36084 5108 36136 5117
rect 36544 5151 36596 5160
rect 36544 5117 36553 5151
rect 36553 5117 36587 5151
rect 36587 5117 36596 5151
rect 36544 5108 36596 5117
rect 35992 5040 36044 5092
rect 24216 4972 24268 4981
rect 30012 4972 30064 5024
rect 34428 4972 34480 5024
rect 19606 4870 19658 4922
rect 19670 4870 19722 4922
rect 19734 4870 19786 4922
rect 19798 4870 19850 4922
rect 2872 4768 2924 4820
rect 5172 4768 5224 4820
rect 6920 4768 6972 4820
rect 8116 4811 8168 4820
rect 8116 4777 8125 4811
rect 8125 4777 8159 4811
rect 8159 4777 8168 4811
rect 8116 4768 8168 4777
rect 4804 4632 4856 4684
rect 6368 4632 6420 4684
rect 11244 4768 11296 4820
rect 11428 4768 11480 4820
rect 11796 4768 11848 4820
rect 8668 4675 8720 4684
rect 8668 4641 8677 4675
rect 8677 4641 8711 4675
rect 8711 4641 8720 4675
rect 8668 4632 8720 4641
rect 9680 4632 9732 4684
rect 10324 4632 10376 4684
rect 10508 4675 10560 4684
rect 10508 4641 10517 4675
rect 10517 4641 10551 4675
rect 10551 4641 10560 4675
rect 10508 4632 10560 4641
rect 12716 4632 12768 4684
rect 14372 4632 14424 4684
rect 15200 4632 15252 4684
rect 19064 4768 19116 4820
rect 24308 4811 24360 4820
rect 24308 4777 24317 4811
rect 24317 4777 24351 4811
rect 24351 4777 24360 4811
rect 24308 4768 24360 4777
rect 25044 4768 25096 4820
rect 36636 4811 36688 4820
rect 36636 4777 36645 4811
rect 36645 4777 36679 4811
rect 36679 4777 36688 4811
rect 36636 4768 36688 4777
rect 16120 4632 16172 4684
rect 16856 4675 16908 4684
rect 16856 4641 16865 4675
rect 16865 4641 16899 4675
rect 16899 4641 16908 4675
rect 16856 4632 16908 4641
rect 17408 4700 17460 4752
rect 29552 4700 29604 4752
rect 32128 4743 32180 4752
rect 32128 4709 32137 4743
rect 32137 4709 32171 4743
rect 32171 4709 32180 4743
rect 32128 4700 32180 4709
rect 3700 4564 3752 4616
rect 6920 4564 6972 4616
rect 9128 4607 9180 4616
rect 9128 4573 9137 4607
rect 9137 4573 9171 4607
rect 9171 4573 9180 4607
rect 9128 4564 9180 4573
rect 20812 4632 20864 4684
rect 21456 4632 21508 4684
rect 21824 4632 21876 4684
rect 24860 4632 24912 4684
rect 26148 4632 26200 4684
rect 27620 4675 27672 4684
rect 27620 4641 27629 4675
rect 27629 4641 27663 4675
rect 27663 4641 27672 4675
rect 27620 4632 27672 4641
rect 27804 4632 27856 4684
rect 29368 4632 29420 4684
rect 31392 4632 31444 4684
rect 32588 4632 32640 4684
rect 34336 4632 34388 4684
rect 34428 4675 34480 4684
rect 34428 4641 34437 4675
rect 34437 4641 34471 4675
rect 34471 4641 34480 4675
rect 34428 4632 34480 4641
rect 17960 4607 18012 4616
rect 8116 4496 8168 4548
rect 10048 4496 10100 4548
rect 17960 4573 17969 4607
rect 17969 4573 18003 4607
rect 18003 4573 18012 4607
rect 17960 4564 18012 4573
rect 21548 4564 21600 4616
rect 29000 4564 29052 4616
rect 31024 4564 31076 4616
rect 31760 4564 31812 4616
rect 33600 4607 33652 4616
rect 33600 4573 33609 4607
rect 33609 4573 33643 4607
rect 33643 4573 33652 4607
rect 33600 4564 33652 4573
rect 34520 4564 34572 4616
rect 35348 4607 35400 4616
rect 13452 4496 13504 4548
rect 20720 4496 20772 4548
rect 26884 4496 26936 4548
rect 35348 4573 35357 4607
rect 35357 4573 35391 4607
rect 35391 4573 35400 4607
rect 35348 4564 35400 4573
rect 7012 4428 7064 4480
rect 4246 4326 4298 4378
rect 4310 4326 4362 4378
rect 4374 4326 4426 4378
rect 4438 4326 4490 4378
rect 34966 4326 35018 4378
rect 35030 4326 35082 4378
rect 35094 4326 35146 4378
rect 35158 4326 35210 4378
rect 5816 4224 5868 4276
rect 35900 4224 35952 4276
rect 3700 4131 3752 4140
rect 3700 4097 3709 4131
rect 3709 4097 3743 4131
rect 3743 4097 3752 4131
rect 3700 4088 3752 4097
rect 4068 4088 4120 4140
rect 6368 4088 6420 4140
rect 6000 4063 6052 4072
rect 6000 4029 6009 4063
rect 6009 4029 6043 4063
rect 6043 4029 6052 4063
rect 6000 4020 6052 4029
rect 7104 4063 7156 4072
rect 7104 4029 7113 4063
rect 7113 4029 7147 4063
rect 7147 4029 7156 4063
rect 7104 4020 7156 4029
rect 8576 4156 8628 4208
rect 8116 4088 8168 4140
rect 8484 4020 8536 4072
rect 9220 4088 9272 4140
rect 12900 4088 12952 4140
rect 14740 4131 14792 4140
rect 14740 4097 14749 4131
rect 14749 4097 14783 4131
rect 14783 4097 14792 4131
rect 14740 4088 14792 4097
rect 15384 4088 15436 4140
rect 16304 4088 16356 4140
rect 17776 4088 17828 4140
rect 9312 4020 9364 4072
rect 5264 3927 5316 3936
rect 5264 3893 5273 3927
rect 5273 3893 5307 3927
rect 5307 3893 5316 3927
rect 5264 3884 5316 3893
rect 6920 3927 6972 3936
rect 6920 3893 6929 3927
rect 6929 3893 6963 3927
rect 6963 3893 6972 3927
rect 6920 3884 6972 3893
rect 10048 3884 10100 3936
rect 11244 4020 11296 4072
rect 11520 4063 11572 4072
rect 10324 3952 10376 4004
rect 11520 4029 11529 4063
rect 11529 4029 11563 4063
rect 11563 4029 11572 4063
rect 11520 4020 11572 4029
rect 13268 4063 13320 4072
rect 13268 4029 13277 4063
rect 13277 4029 13311 4063
rect 13311 4029 13320 4063
rect 13268 4020 13320 4029
rect 13452 4063 13504 4072
rect 13452 4029 13461 4063
rect 13461 4029 13495 4063
rect 13495 4029 13504 4063
rect 13452 4020 13504 4029
rect 14464 4063 14516 4072
rect 14464 4029 14473 4063
rect 14473 4029 14507 4063
rect 14507 4029 14516 4063
rect 14464 4020 14516 4029
rect 11888 3952 11940 4004
rect 13820 3952 13872 4004
rect 17224 4063 17276 4072
rect 17224 4029 17233 4063
rect 17233 4029 17267 4063
rect 17267 4029 17276 4063
rect 17224 4020 17276 4029
rect 18144 3952 18196 4004
rect 18696 4020 18748 4072
rect 19064 4063 19116 4072
rect 19064 4029 19073 4063
rect 19073 4029 19107 4063
rect 19107 4029 19116 4063
rect 19064 4020 19116 4029
rect 22100 4156 22152 4208
rect 19248 4088 19300 4140
rect 20444 4088 20496 4140
rect 26424 4088 26476 4140
rect 26700 4088 26752 4140
rect 29460 4199 29512 4208
rect 29460 4165 29469 4199
rect 29469 4165 29503 4199
rect 29503 4165 29512 4199
rect 29460 4156 29512 4165
rect 30932 4131 30984 4140
rect 19984 4063 20036 4072
rect 19340 3995 19392 4004
rect 19340 3961 19349 3995
rect 19349 3961 19383 3995
rect 19383 3961 19392 3995
rect 19340 3952 19392 3961
rect 19984 4029 19993 4063
rect 19993 4029 20027 4063
rect 20027 4029 20036 4063
rect 19984 4020 20036 4029
rect 21732 4020 21784 4072
rect 22192 4063 22244 4072
rect 22192 4029 22201 4063
rect 22201 4029 22235 4063
rect 22235 4029 22244 4063
rect 22192 4020 22244 4029
rect 25872 4063 25924 4072
rect 20996 3952 21048 4004
rect 24492 3952 24544 4004
rect 25872 4029 25881 4063
rect 25881 4029 25915 4063
rect 25915 4029 25924 4063
rect 25872 4020 25924 4029
rect 26056 4063 26108 4072
rect 26056 4029 26065 4063
rect 26065 4029 26099 4063
rect 26099 4029 26108 4063
rect 26056 4020 26108 4029
rect 26332 4020 26384 4072
rect 27068 4020 27120 4072
rect 29276 4063 29328 4072
rect 29276 4029 29285 4063
rect 29285 4029 29319 4063
rect 29319 4029 29328 4063
rect 29276 4020 29328 4029
rect 17868 3884 17920 3936
rect 18420 3884 18472 3936
rect 18972 3884 19024 3936
rect 23756 3884 23808 3936
rect 27528 3952 27580 4004
rect 26424 3884 26476 3936
rect 26516 3884 26568 3936
rect 27896 3927 27948 3936
rect 27896 3893 27905 3927
rect 27905 3893 27939 3927
rect 27939 3893 27948 3927
rect 27896 3884 27948 3893
rect 30932 4097 30941 4131
rect 30941 4097 30975 4131
rect 30975 4097 30984 4131
rect 30932 4088 30984 4097
rect 33968 4156 34020 4208
rect 31944 4088 31996 4140
rect 31760 4020 31812 4072
rect 32128 4020 32180 4072
rect 32772 4088 32824 4140
rect 33048 4088 33100 4140
rect 34428 4156 34480 4208
rect 32864 4063 32916 4072
rect 32864 4029 32873 4063
rect 32873 4029 32907 4063
rect 32907 4029 32916 4063
rect 32864 4020 32916 4029
rect 33876 4063 33928 4072
rect 33876 4029 33885 4063
rect 33885 4029 33919 4063
rect 33919 4029 33928 4063
rect 33876 4020 33928 4029
rect 33968 4020 34020 4072
rect 34612 4088 34664 4140
rect 34428 4020 34480 4072
rect 35440 4063 35492 4072
rect 35440 4029 35449 4063
rect 35449 4029 35483 4063
rect 35483 4029 35492 4063
rect 35440 4020 35492 4029
rect 35992 4088 36044 4140
rect 31852 3995 31904 4004
rect 31852 3961 31861 3995
rect 31861 3961 31895 3995
rect 31895 3961 31904 3995
rect 31852 3952 31904 3961
rect 32036 3952 32088 4004
rect 35348 3884 35400 3936
rect 19606 3782 19658 3834
rect 19670 3782 19722 3834
rect 19734 3782 19786 3834
rect 19798 3782 19850 3834
rect 7380 3680 7432 3732
rect 7472 3680 7524 3732
rect 6000 3612 6052 3664
rect 5264 3587 5316 3596
rect 5264 3553 5273 3587
rect 5273 3553 5307 3587
rect 5307 3553 5316 3587
rect 5264 3544 5316 3553
rect 6368 3587 6420 3596
rect 6368 3553 6377 3587
rect 6377 3553 6411 3587
rect 6411 3553 6420 3587
rect 6368 3544 6420 3553
rect 7104 3587 7156 3596
rect 7104 3553 7113 3587
rect 7113 3553 7147 3587
rect 7147 3553 7156 3587
rect 7104 3544 7156 3553
rect 8576 3544 8628 3596
rect 8760 3612 8812 3664
rect 20996 3680 21048 3732
rect 8944 3544 8996 3596
rect 10324 3612 10376 3664
rect 10416 3612 10468 3664
rect 27068 3680 27120 3732
rect 10140 3587 10192 3596
rect 5172 3519 5224 3528
rect 5172 3485 5181 3519
rect 5181 3485 5215 3519
rect 5215 3485 5224 3519
rect 5172 3476 5224 3485
rect 5724 3519 5776 3528
rect 5724 3485 5733 3519
rect 5733 3485 5767 3519
rect 5767 3485 5776 3519
rect 5724 3476 5776 3485
rect 6092 3408 6144 3460
rect 6828 3408 6880 3460
rect 8668 3408 8720 3460
rect 10140 3553 10149 3587
rect 10149 3553 10183 3587
rect 10183 3553 10192 3587
rect 10140 3544 10192 3553
rect 11244 3544 11296 3596
rect 11888 3587 11940 3596
rect 11888 3553 11897 3587
rect 11897 3553 11931 3587
rect 11931 3553 11940 3587
rect 11888 3544 11940 3553
rect 13268 3544 13320 3596
rect 14188 3587 14240 3596
rect 14188 3553 14197 3587
rect 14197 3553 14231 3587
rect 14231 3553 14240 3587
rect 14188 3544 14240 3553
rect 14464 3544 14516 3596
rect 16212 3587 16264 3596
rect 10416 3476 10468 3528
rect 13544 3476 13596 3528
rect 14280 3519 14332 3528
rect 14280 3485 14289 3519
rect 14289 3485 14323 3519
rect 14323 3485 14332 3519
rect 14280 3476 14332 3485
rect 16212 3553 16221 3587
rect 16221 3553 16255 3587
rect 16255 3553 16264 3587
rect 16212 3544 16264 3553
rect 16304 3544 16356 3596
rect 18052 3587 18104 3596
rect 18052 3553 18061 3587
rect 18061 3553 18095 3587
rect 18095 3553 18104 3587
rect 18052 3544 18104 3553
rect 21364 3587 21416 3596
rect 17960 3476 18012 3528
rect 18236 3476 18288 3528
rect 18420 3476 18472 3528
rect 19892 3476 19944 3528
rect 21364 3553 21373 3587
rect 21373 3553 21407 3587
rect 21407 3553 21416 3587
rect 21364 3544 21416 3553
rect 22652 3544 22704 3596
rect 22836 3587 22888 3596
rect 22836 3553 22845 3587
rect 22845 3553 22879 3587
rect 22879 3553 22888 3587
rect 22836 3544 22888 3553
rect 25872 3544 25924 3596
rect 27896 3612 27948 3664
rect 30104 3680 30156 3732
rect 30288 3680 30340 3732
rect 30656 3680 30708 3732
rect 31392 3680 31444 3732
rect 32864 3680 32916 3732
rect 34336 3680 34388 3732
rect 27988 3587 28040 3596
rect 27988 3553 27997 3587
rect 27997 3553 28031 3587
rect 28031 3553 28040 3587
rect 27988 3544 28040 3553
rect 28264 3587 28316 3596
rect 28264 3553 28273 3587
rect 28273 3553 28307 3587
rect 28307 3553 28316 3587
rect 28264 3544 28316 3553
rect 31944 3612 31996 3664
rect 32128 3655 32180 3664
rect 32128 3621 32137 3655
rect 32137 3621 32171 3655
rect 32171 3621 32180 3655
rect 32128 3612 32180 3621
rect 31852 3544 31904 3596
rect 21732 3476 21784 3528
rect 22100 3476 22152 3528
rect 27804 3476 27856 3528
rect 10048 3408 10100 3460
rect 11152 3408 11204 3460
rect 19064 3408 19116 3460
rect 22284 3408 22336 3460
rect 23848 3408 23900 3460
rect 26700 3408 26752 3460
rect 27068 3408 27120 3460
rect 29092 3476 29144 3528
rect 29552 3476 29604 3528
rect 30564 3476 30616 3528
rect 33416 3544 33468 3596
rect 33692 3544 33744 3596
rect 35992 3544 36044 3596
rect 32680 3519 32732 3528
rect 32680 3485 32689 3519
rect 32689 3485 32723 3519
rect 32723 3485 32732 3519
rect 32680 3476 32732 3485
rect 6552 3383 6604 3392
rect 6552 3349 6561 3383
rect 6561 3349 6595 3383
rect 6595 3349 6604 3383
rect 6552 3340 6604 3349
rect 16580 3340 16632 3392
rect 18328 3340 18380 3392
rect 21548 3340 21600 3392
rect 24124 3383 24176 3392
rect 24124 3349 24133 3383
rect 24133 3349 24167 3383
rect 24167 3349 24176 3383
rect 24124 3340 24176 3349
rect 24768 3340 24820 3392
rect 26884 3340 26936 3392
rect 28264 3340 28316 3392
rect 30564 3340 30616 3392
rect 30656 3340 30708 3392
rect 33508 3476 33560 3528
rect 33416 3340 33468 3392
rect 35716 3340 35768 3392
rect 4246 3238 4298 3290
rect 4310 3238 4362 3290
rect 4374 3238 4426 3290
rect 4438 3238 4490 3290
rect 34966 3238 35018 3290
rect 35030 3238 35082 3290
rect 35094 3238 35146 3290
rect 35158 3238 35210 3290
rect 6552 3136 6604 3188
rect 10876 3179 10928 3188
rect 1400 3000 1452 3052
rect 7104 3000 7156 3052
rect 7472 3043 7524 3052
rect 7472 3009 7481 3043
rect 7481 3009 7515 3043
rect 7515 3009 7524 3043
rect 7472 3000 7524 3009
rect 9128 3000 9180 3052
rect 10876 3145 10885 3179
rect 10885 3145 10919 3179
rect 10919 3145 10928 3179
rect 10876 3136 10928 3145
rect 11060 3136 11112 3188
rect 11704 3068 11756 3120
rect 18236 3136 18288 3188
rect 13544 3043 13596 3052
rect 1952 2932 2004 2984
rect 5816 2975 5868 2984
rect 5816 2941 5825 2975
rect 5825 2941 5859 2975
rect 5859 2941 5868 2975
rect 5816 2932 5868 2941
rect 6092 2975 6144 2984
rect 6092 2941 6101 2975
rect 6101 2941 6135 2975
rect 6135 2941 6144 2975
rect 6092 2932 6144 2941
rect 6920 2932 6972 2984
rect 10416 2932 10468 2984
rect 11152 2932 11204 2984
rect 12348 2932 12400 2984
rect 13544 3009 13553 3043
rect 13553 3009 13587 3043
rect 13587 3009 13596 3043
rect 13544 3000 13596 3009
rect 13820 3043 13872 3052
rect 13820 3009 13829 3043
rect 13829 3009 13863 3043
rect 13863 3009 13872 3043
rect 13820 3000 13872 3009
rect 16120 3068 16172 3120
rect 23848 3136 23900 3188
rect 26056 3136 26108 3188
rect 27712 3136 27764 3188
rect 27804 3136 27856 3188
rect 28724 3136 28776 3188
rect 31392 3179 31444 3188
rect 31392 3145 31401 3179
rect 31401 3145 31435 3179
rect 31435 3145 31444 3179
rect 31392 3136 31444 3145
rect 33968 3136 34020 3188
rect 2596 2796 2648 2848
rect 12440 2796 12492 2848
rect 16580 3000 16632 3052
rect 15200 2864 15252 2916
rect 18144 2975 18196 2984
rect 18144 2941 18153 2975
rect 18153 2941 18187 2975
rect 18187 2941 18196 2975
rect 18144 2932 18196 2941
rect 18604 2975 18656 2984
rect 18604 2941 18613 2975
rect 18613 2941 18647 2975
rect 18647 2941 18656 2975
rect 18604 2932 18656 2941
rect 17224 2907 17276 2916
rect 17224 2873 17233 2907
rect 17233 2873 17267 2907
rect 17267 2873 17276 2907
rect 17224 2864 17276 2873
rect 18880 2907 18932 2916
rect 18880 2873 18889 2907
rect 18889 2873 18923 2907
rect 18923 2873 18932 2907
rect 18880 2864 18932 2873
rect 19340 3000 19392 3052
rect 19432 2932 19484 2984
rect 21824 2932 21876 2984
rect 24124 3000 24176 3052
rect 24032 2932 24084 2984
rect 24768 2932 24820 2984
rect 24308 2864 24360 2916
rect 26332 2932 26384 2984
rect 27068 2975 27120 2984
rect 27068 2941 27077 2975
rect 27077 2941 27111 2975
rect 27111 2941 27120 2975
rect 27068 2932 27120 2941
rect 26424 2864 26476 2916
rect 27712 2932 27764 2984
rect 29092 2932 29144 2984
rect 32036 2932 32088 2984
rect 33600 3000 33652 3052
rect 34520 3000 34572 3052
rect 35440 3043 35492 3052
rect 35440 3009 35449 3043
rect 35449 3009 35483 3043
rect 35483 3009 35492 3043
rect 35440 3000 35492 3009
rect 30104 2864 30156 2916
rect 27988 2796 28040 2848
rect 30288 2796 30340 2848
rect 32036 2796 32088 2848
rect 33140 2932 33192 2984
rect 35716 2975 35768 2984
rect 35716 2941 35725 2975
rect 35725 2941 35759 2975
rect 35759 2941 35768 2975
rect 35716 2932 35768 2941
rect 36360 2864 36412 2916
rect 33508 2796 33560 2848
rect 19606 2694 19658 2746
rect 19670 2694 19722 2746
rect 19734 2694 19786 2746
rect 19798 2694 19850 2746
rect 8576 2592 8628 2644
rect 16488 2592 16540 2644
rect 18604 2592 18656 2644
rect 19984 2592 20036 2644
rect 24032 2592 24084 2644
rect 30288 2592 30340 2644
rect 15200 2524 15252 2576
rect 3700 2456 3752 2508
rect 4988 2456 5040 2508
rect 6920 2499 6972 2508
rect 6920 2465 6929 2499
rect 6929 2465 6963 2499
rect 6963 2465 6972 2499
rect 6920 2456 6972 2465
rect 8852 2456 8904 2508
rect 10416 2499 10468 2508
rect 10416 2465 10425 2499
rect 10425 2465 10459 2499
rect 10459 2465 10468 2499
rect 10416 2456 10468 2465
rect 11060 2456 11112 2508
rect 14280 2456 14332 2508
rect 17224 2456 17276 2508
rect 18328 2499 18380 2508
rect 18328 2465 18337 2499
rect 18337 2465 18371 2499
rect 18371 2465 18380 2499
rect 18328 2456 18380 2465
rect 18880 2456 18932 2508
rect 19524 2456 19576 2508
rect 21364 2524 21416 2576
rect 22100 2499 22152 2508
rect 22100 2465 22109 2499
rect 22109 2465 22143 2499
rect 22143 2465 22152 2499
rect 26608 2524 26660 2576
rect 22100 2456 22152 2465
rect 24308 2499 24360 2508
rect 24308 2465 24317 2499
rect 24317 2465 24351 2499
rect 24351 2465 24360 2499
rect 24308 2456 24360 2465
rect 26884 2499 26936 2508
rect 26884 2465 26893 2499
rect 26893 2465 26927 2499
rect 26927 2465 26936 2499
rect 26884 2456 26936 2465
rect 29460 2524 29512 2576
rect 5724 2388 5776 2440
rect 18052 2388 18104 2440
rect 22560 2388 22612 2440
rect 26700 2388 26752 2440
rect 30012 2456 30064 2508
rect 33876 2524 33928 2576
rect 30564 2499 30616 2508
rect 30564 2465 30573 2499
rect 30573 2465 30607 2499
rect 30607 2465 30616 2499
rect 30564 2456 30616 2465
rect 31392 2456 31444 2508
rect 33416 2499 33468 2508
rect 33140 2431 33192 2440
rect 4712 2252 4764 2304
rect 28724 2320 28776 2372
rect 33140 2397 33149 2431
rect 33149 2397 33183 2431
rect 33183 2397 33192 2431
rect 33140 2388 33192 2397
rect 33416 2465 33425 2499
rect 33425 2465 33459 2499
rect 33459 2465 33468 2499
rect 33416 2456 33468 2465
rect 11060 2252 11112 2304
rect 13084 2252 13136 2304
rect 17316 2252 17368 2304
rect 23388 2295 23440 2304
rect 23388 2261 23397 2295
rect 23397 2261 23431 2295
rect 23431 2261 23440 2295
rect 23388 2252 23440 2261
rect 25596 2295 25648 2304
rect 25596 2261 25605 2295
rect 25605 2261 25639 2295
rect 25639 2261 25648 2295
rect 25596 2252 25648 2261
rect 38476 2295 38528 2304
rect 38476 2261 38485 2295
rect 38485 2261 38519 2295
rect 38519 2261 38528 2295
rect 38476 2252 38528 2261
rect 4246 2150 4298 2202
rect 4310 2150 4362 2202
rect 4374 2150 4426 2202
rect 4438 2150 4490 2202
rect 34966 2150 35018 2202
rect 35030 2150 35082 2202
rect 35094 2150 35146 2202
rect 35158 2150 35210 2202
rect 19524 2048 19576 2100
rect 20076 2048 20128 2100
rect 23388 2048 23440 2100
rect 34244 2048 34296 2100
rect 25596 1980 25648 2032
rect 36452 1980 36504 2032
rect 19892 1912 19944 1964
rect 25780 1912 25832 1964
rect 572 1776 624 1828
rect 8760 1776 8812 1828
<< metal2 >>
rect 1306 40200 1362 41000
rect 3330 40200 3386 41000
rect 5538 40200 5594 41000
rect 7562 40200 7618 41000
rect 9770 40200 9826 41000
rect 11794 40200 11850 41000
rect 14002 40200 14058 41000
rect 16026 40200 16082 41000
rect 18234 40200 18290 41000
rect 20258 40200 20314 41000
rect 22466 40200 22522 41000
rect 24490 40200 24546 41000
rect 26698 40200 26754 41000
rect 28722 40200 28778 41000
rect 30930 40200 30986 41000
rect 32954 40200 33010 41000
rect 35162 40200 35218 41000
rect 37186 40200 37242 41000
rect 39394 40200 39450 41000
rect 1320 38418 1348 40200
rect 1308 38412 1360 38418
rect 1308 38354 1360 38360
rect 1858 38176 1914 38185
rect 1858 38111 1914 38120
rect 1872 37330 1900 38111
rect 3344 37874 3372 40200
rect 5552 38196 5580 40200
rect 7576 38554 7604 40200
rect 7564 38548 7616 38554
rect 7564 38490 7616 38496
rect 9680 38480 9732 38486
rect 9678 38448 9680 38457
rect 9732 38448 9734 38457
rect 9036 38412 9088 38418
rect 9678 38383 9734 38392
rect 9036 38354 9088 38360
rect 6092 38344 6144 38350
rect 6092 38286 6144 38292
rect 7932 38344 7984 38350
rect 7932 38286 7984 38292
rect 5552 38168 5672 38196
rect 4220 38108 4516 38128
rect 4276 38106 4300 38108
rect 4356 38106 4380 38108
rect 4436 38106 4460 38108
rect 4298 38054 4300 38106
rect 4362 38054 4374 38106
rect 4436 38054 4438 38106
rect 4276 38052 4300 38054
rect 4356 38052 4380 38054
rect 4436 38052 4460 38054
rect 4220 38032 4516 38052
rect 3332 37868 3384 37874
rect 3332 37810 3384 37816
rect 5172 37800 5224 37806
rect 5172 37742 5224 37748
rect 1860 37324 1912 37330
rect 1860 37266 1912 37272
rect 4220 37020 4516 37040
rect 4276 37018 4300 37020
rect 4356 37018 4380 37020
rect 4436 37018 4460 37020
rect 4298 36966 4300 37018
rect 4362 36966 4374 37018
rect 4436 36966 4438 37018
rect 4276 36964 4300 36966
rect 4356 36964 4380 36966
rect 4436 36964 4460 36966
rect 4220 36944 4516 36964
rect 4988 36100 5040 36106
rect 4988 36042 5040 36048
rect 4220 35932 4516 35952
rect 4276 35930 4300 35932
rect 4356 35930 4380 35932
rect 4436 35930 4460 35932
rect 4298 35878 4300 35930
rect 4362 35878 4374 35930
rect 4436 35878 4438 35930
rect 4276 35876 4300 35878
rect 4356 35876 4380 35878
rect 4436 35876 4460 35878
rect 4220 35856 4516 35876
rect 3792 35624 3844 35630
rect 3792 35566 3844 35572
rect 4160 35624 4212 35630
rect 4160 35566 4212 35572
rect 2872 35488 2924 35494
rect 2872 35430 2924 35436
rect 1952 35148 2004 35154
rect 1952 35090 2004 35096
rect 1964 34542 1992 35090
rect 2136 35080 2188 35086
rect 2136 35022 2188 35028
rect 2688 35080 2740 35086
rect 2688 35022 2740 35028
rect 2148 34746 2176 35022
rect 2136 34740 2188 34746
rect 2136 34682 2188 34688
rect 2700 34610 2728 35022
rect 2780 34944 2832 34950
rect 2780 34886 2832 34892
rect 2688 34604 2740 34610
rect 2688 34546 2740 34552
rect 1768 34536 1820 34542
rect 1768 34478 1820 34484
rect 1952 34536 2004 34542
rect 1952 34478 2004 34484
rect 1780 34134 1808 34478
rect 1768 34128 1820 34134
rect 1768 34070 1820 34076
rect 2700 32978 2728 34546
rect 2792 34134 2820 34886
rect 2780 34128 2832 34134
rect 2780 34070 2832 34076
rect 2792 33454 2820 34070
rect 2780 33448 2832 33454
rect 2780 33390 2832 33396
rect 2688 32972 2740 32978
rect 2688 32914 2740 32920
rect 1676 32904 1728 32910
rect 1676 32846 1728 32852
rect 1688 32026 1716 32846
rect 1676 32020 1728 32026
rect 1676 31962 1728 31968
rect 2504 31884 2556 31890
rect 2504 31826 2556 31832
rect 1676 31272 1728 31278
rect 1676 31214 1728 31220
rect 1688 30938 1716 31214
rect 1676 30932 1728 30938
rect 1676 30874 1728 30880
rect 2516 30818 2544 31826
rect 2700 31346 2728 32914
rect 2884 31929 2912 35430
rect 3606 35184 3662 35193
rect 3606 35119 3662 35128
rect 3056 34128 3108 34134
rect 3056 34070 3108 34076
rect 2964 33992 3016 33998
rect 2964 33934 3016 33940
rect 2976 32434 3004 33934
rect 3068 32502 3096 34070
rect 3148 34060 3200 34066
rect 3148 34002 3200 34008
rect 3332 34060 3384 34066
rect 3332 34002 3384 34008
rect 3160 33658 3188 34002
rect 3148 33652 3200 33658
rect 3148 33594 3200 33600
rect 3056 32496 3108 32502
rect 3056 32438 3108 32444
rect 2964 32428 3016 32434
rect 2964 32370 3016 32376
rect 2870 31920 2926 31929
rect 2870 31855 2926 31864
rect 2872 31476 2924 31482
rect 2872 31418 2924 31424
rect 2688 31340 2740 31346
rect 2688 31282 2740 31288
rect 2884 30870 2912 31418
rect 2872 30864 2924 30870
rect 2516 30802 2728 30818
rect 2872 30806 2924 30812
rect 2516 30796 2740 30802
rect 2516 30790 2688 30796
rect 2688 30738 2740 30744
rect 2412 30184 2464 30190
rect 2412 30126 2464 30132
rect 1400 29640 1452 29646
rect 1400 29582 1452 29588
rect 1860 29640 1912 29646
rect 1860 29582 1912 29588
rect 1412 27538 1440 29582
rect 1872 29306 1900 29582
rect 1860 29300 1912 29306
rect 1860 29242 1912 29248
rect 2424 29102 2452 30126
rect 2412 29096 2464 29102
rect 2412 29038 2464 29044
rect 2320 28620 2372 28626
rect 2320 28562 2372 28568
rect 1952 28416 2004 28422
rect 1952 28358 2004 28364
rect 1400 27532 1452 27538
rect 1400 27474 1452 27480
rect 1964 26518 1992 28358
rect 2332 28014 2360 28562
rect 2412 28416 2464 28422
rect 2412 28358 2464 28364
rect 2320 28008 2372 28014
rect 2320 27950 2372 27956
rect 2332 27130 2360 27950
rect 2424 27538 2452 28358
rect 2700 27606 2728 30738
rect 2780 30592 2832 30598
rect 2780 30534 2832 30540
rect 2792 30190 2820 30534
rect 2780 30184 2832 30190
rect 2780 30126 2832 30132
rect 2976 29238 3004 32370
rect 3056 32292 3108 32298
rect 3056 32234 3108 32240
rect 3068 31890 3096 32234
rect 3160 32230 3188 33594
rect 3344 33454 3372 34002
rect 3332 33448 3384 33454
rect 3332 33390 3384 33396
rect 3344 33046 3372 33390
rect 3332 33040 3384 33046
rect 3332 32982 3384 32988
rect 3240 32496 3292 32502
rect 3240 32438 3292 32444
rect 3148 32224 3200 32230
rect 3148 32166 3200 32172
rect 3252 31890 3280 32438
rect 3344 32366 3372 32982
rect 3332 32360 3384 32366
rect 3332 32302 3384 32308
rect 3056 31884 3108 31890
rect 3056 31826 3108 31832
rect 3240 31884 3292 31890
rect 3240 31826 3292 31832
rect 3240 31136 3292 31142
rect 3240 31078 3292 31084
rect 3252 30802 3280 31078
rect 3240 30796 3292 30802
rect 3240 30738 3292 30744
rect 3056 30184 3108 30190
rect 3056 30126 3108 30132
rect 3240 30184 3292 30190
rect 3240 30126 3292 30132
rect 2964 29232 3016 29238
rect 2964 29174 3016 29180
rect 3068 29102 3096 30126
rect 3148 30048 3200 30054
rect 3148 29990 3200 29996
rect 3160 29510 3188 29990
rect 3148 29504 3200 29510
rect 3148 29446 3200 29452
rect 3056 29096 3108 29102
rect 3056 29038 3108 29044
rect 3054 28928 3110 28937
rect 3054 28863 3110 28872
rect 3068 28234 3096 28863
rect 3160 28626 3188 29446
rect 3252 29102 3280 30126
rect 3240 29096 3292 29102
rect 3240 29038 3292 29044
rect 3148 28620 3200 28626
rect 3148 28562 3200 28568
rect 3068 28206 3188 28234
rect 2964 28008 3016 28014
rect 2964 27950 3016 27956
rect 2976 27674 3004 27950
rect 2964 27668 3016 27674
rect 2964 27610 3016 27616
rect 2688 27600 2740 27606
rect 2688 27542 2740 27548
rect 2412 27532 2464 27538
rect 2412 27474 2464 27480
rect 2320 27124 2372 27130
rect 2320 27066 2372 27072
rect 2412 26920 2464 26926
rect 2412 26862 2464 26868
rect 1952 26512 2004 26518
rect 1952 26454 2004 26460
rect 2424 26450 2452 26862
rect 2412 26444 2464 26450
rect 2412 26386 2464 26392
rect 1676 25288 1728 25294
rect 1676 25230 1728 25236
rect 1584 24744 1636 24750
rect 1584 24686 1636 24692
rect 1400 23112 1452 23118
rect 1400 23054 1452 23060
rect 1412 21010 1440 23054
rect 1596 22681 1624 24686
rect 1688 24342 1716 25230
rect 2700 24750 2728 27542
rect 2780 27464 2832 27470
rect 2780 27406 2832 27412
rect 2792 25906 2820 27406
rect 2976 27062 3004 27610
rect 2964 27056 3016 27062
rect 2964 26998 3016 27004
rect 2872 26920 2924 26926
rect 2872 26862 2924 26868
rect 3056 26920 3108 26926
rect 3056 26862 3108 26868
rect 2884 26450 2912 26862
rect 2872 26444 2924 26450
rect 2872 26386 2924 26392
rect 2780 25900 2832 25906
rect 2780 25842 2832 25848
rect 2792 25362 2820 25842
rect 2884 25498 2912 26386
rect 2964 26376 3016 26382
rect 3068 26330 3096 26862
rect 3016 26324 3096 26330
rect 2964 26318 3096 26324
rect 2976 26302 3096 26318
rect 2872 25492 2924 25498
rect 2872 25434 2924 25440
rect 2780 25356 2832 25362
rect 2780 25298 2832 25304
rect 2792 24886 2820 25298
rect 2780 24880 2832 24886
rect 2780 24822 2832 24828
rect 2884 24818 2912 25434
rect 2976 25362 3004 26302
rect 2964 25356 3016 25362
rect 2964 25298 3016 25304
rect 2872 24812 2924 24818
rect 2872 24754 2924 24760
rect 2228 24744 2280 24750
rect 2228 24686 2280 24692
rect 2688 24744 2740 24750
rect 2688 24686 2740 24692
rect 1676 24336 1728 24342
rect 1676 24278 1728 24284
rect 2044 23656 2096 23662
rect 2044 23598 2096 23604
rect 1768 23112 1820 23118
rect 1768 23054 1820 23060
rect 1780 22778 1808 23054
rect 1768 22772 1820 22778
rect 1768 22714 1820 22720
rect 2056 22710 2084 23598
rect 2044 22704 2096 22710
rect 1582 22672 1638 22681
rect 2044 22646 2096 22652
rect 1582 22607 1638 22616
rect 1492 22092 1544 22098
rect 2240 22080 2268 24686
rect 2412 24608 2464 24614
rect 2412 24550 2464 24556
rect 2424 24274 2452 24550
rect 2412 24268 2464 24274
rect 2412 24210 2464 24216
rect 2780 24268 2832 24274
rect 2884 24256 2912 24754
rect 2976 24750 3004 25298
rect 2964 24744 3016 24750
rect 2964 24686 3016 24692
rect 2976 24274 3004 24686
rect 2832 24228 2912 24256
rect 2964 24268 3016 24274
rect 2780 24210 2832 24216
rect 2964 24210 3016 24216
rect 2780 23724 2832 23730
rect 2780 23666 2832 23672
rect 2412 23656 2464 23662
rect 2412 23598 2464 23604
rect 1492 22034 1544 22040
rect 2056 22052 2268 22080
rect 1504 21622 1532 22034
rect 1676 21888 1728 21894
rect 1676 21830 1728 21836
rect 1492 21616 1544 21622
rect 1492 21558 1544 21564
rect 1688 21010 1716 21830
rect 1400 21004 1452 21010
rect 1400 20946 1452 20952
rect 1676 21004 1728 21010
rect 1676 20946 1728 20952
rect 1412 19922 1440 20946
rect 1400 19916 1452 19922
rect 1400 19858 1452 19864
rect 1412 17746 1440 19858
rect 1676 19848 1728 19854
rect 1676 19790 1728 19796
rect 1688 19514 1716 19790
rect 1676 19508 1728 19514
rect 1676 19450 1728 19456
rect 1400 17740 1452 17746
rect 1452 17700 1532 17728
rect 1400 17682 1452 17688
rect 1504 16454 1532 17700
rect 1768 17672 1820 17678
rect 1768 17614 1820 17620
rect 1780 16998 1808 17614
rect 1952 17128 2004 17134
rect 1952 17070 2004 17076
rect 1768 16992 1820 16998
rect 1768 16934 1820 16940
rect 1492 16448 1544 16454
rect 1492 16390 1544 16396
rect 1504 16046 1532 16390
rect 1492 16040 1544 16046
rect 1492 15982 1544 15988
rect 1676 16040 1728 16046
rect 1676 15982 1728 15988
rect 1504 14958 1532 15982
rect 1688 15638 1716 15982
rect 1676 15632 1728 15638
rect 1676 15574 1728 15580
rect 1492 14952 1544 14958
rect 1492 14894 1544 14900
rect 1504 13938 1532 14894
rect 1860 14612 1912 14618
rect 1860 14554 1912 14560
rect 1872 13938 1900 14554
rect 1964 14482 1992 17070
rect 1952 14476 2004 14482
rect 1952 14418 2004 14424
rect 1492 13932 1544 13938
rect 1492 13874 1544 13880
rect 1860 13932 1912 13938
rect 1860 13874 1912 13880
rect 1676 13524 1728 13530
rect 1676 13466 1728 13472
rect 1688 12850 1716 13466
rect 1952 13184 2004 13190
rect 1952 13126 2004 13132
rect 1676 12844 1728 12850
rect 1676 12786 1728 12792
rect 1400 10464 1452 10470
rect 1400 10406 1452 10412
rect 1412 10062 1440 10406
rect 1400 10056 1452 10062
rect 1400 9998 1452 10004
rect 1412 8974 1440 9998
rect 1676 9376 1728 9382
rect 1676 9318 1728 9324
rect 1688 9042 1716 9318
rect 1676 9036 1728 9042
rect 1676 8978 1728 8984
rect 1400 8968 1452 8974
rect 1400 8910 1452 8916
rect 1412 8430 1440 8910
rect 1400 8424 1452 8430
rect 1400 8366 1452 8372
rect 1676 8424 1728 8430
rect 1676 8366 1728 8372
rect 1412 7886 1440 8366
rect 1400 7880 1452 7886
rect 1400 7822 1452 7828
rect 1412 3058 1440 7822
rect 1688 7206 1716 8366
rect 1676 7200 1728 7206
rect 1676 7142 1728 7148
rect 1400 3052 1452 3058
rect 1400 2994 1452 3000
rect 1964 2990 1992 13126
rect 2056 12306 2084 22052
rect 2424 21962 2452 23598
rect 2792 22642 2820 23666
rect 2964 22976 3016 22982
rect 2964 22918 3016 22924
rect 2780 22636 2832 22642
rect 2780 22578 2832 22584
rect 2976 22574 3004 22918
rect 2964 22568 3016 22574
rect 2964 22510 3016 22516
rect 2780 22500 2832 22506
rect 2780 22442 2832 22448
rect 2792 21978 2820 22442
rect 2964 22092 3016 22098
rect 2964 22034 3016 22040
rect 2976 21978 3004 22034
rect 2412 21956 2464 21962
rect 2792 21950 3004 21978
rect 2412 21898 2464 21904
rect 2872 21888 2924 21894
rect 2872 21830 2924 21836
rect 3056 21888 3108 21894
rect 3056 21830 3108 21836
rect 2884 21554 2912 21830
rect 2872 21548 2924 21554
rect 2872 21490 2924 21496
rect 2596 21480 2648 21486
rect 2596 21422 2648 21428
rect 2608 21010 2636 21422
rect 2596 21004 2648 21010
rect 2596 20946 2648 20952
rect 2780 20392 2832 20398
rect 2780 20334 2832 20340
rect 2792 19281 2820 20334
rect 2884 19394 2912 21490
rect 2964 21480 3016 21486
rect 2964 21422 3016 21428
rect 2976 21078 3004 21422
rect 2964 21072 3016 21078
rect 2964 21014 3016 21020
rect 2976 20466 3004 21014
rect 2964 20460 3016 20466
rect 2964 20402 3016 20408
rect 3068 19446 3096 21830
rect 3056 19440 3108 19446
rect 2884 19366 3004 19394
rect 3056 19382 3108 19388
rect 2778 19272 2834 19281
rect 2778 19207 2780 19216
rect 2832 19207 2834 19216
rect 2780 19178 2832 19184
rect 2792 19147 2820 19178
rect 2780 18896 2832 18902
rect 2780 18838 2832 18844
rect 2228 18624 2280 18630
rect 2228 18566 2280 18572
rect 2240 17134 2268 18566
rect 2792 18222 2820 18838
rect 2976 18834 3004 19366
rect 3056 19168 3108 19174
rect 3056 19110 3108 19116
rect 2872 18828 2924 18834
rect 2872 18770 2924 18776
rect 2964 18828 3016 18834
rect 2964 18770 3016 18776
rect 2884 18714 2912 18770
rect 3068 18714 3096 19110
rect 2884 18686 3096 18714
rect 2884 18290 2912 18686
rect 2872 18284 2924 18290
rect 2872 18226 2924 18232
rect 2780 18216 2832 18222
rect 2780 18158 2832 18164
rect 2780 17332 2832 17338
rect 2780 17274 2832 17280
rect 2792 17134 2820 17274
rect 3056 17196 3108 17202
rect 3056 17138 3108 17144
rect 2228 17128 2280 17134
rect 2228 17070 2280 17076
rect 2780 17128 2832 17134
rect 2780 17070 2832 17076
rect 3068 16658 3096 17138
rect 3056 16652 3108 16658
rect 3056 16594 3108 16600
rect 3160 16250 3188 28206
rect 3252 28082 3280 29038
rect 3240 28076 3292 28082
rect 3240 28018 3292 28024
rect 3332 28008 3384 28014
rect 3332 27950 3384 27956
rect 3344 26994 3372 27950
rect 3332 26988 3384 26994
rect 3332 26930 3384 26936
rect 3424 24880 3476 24886
rect 3424 24822 3476 24828
rect 3436 23730 3464 24822
rect 3424 23724 3476 23730
rect 3424 23666 3476 23672
rect 3332 23112 3384 23118
rect 3332 23054 3384 23060
rect 3344 22710 3372 23054
rect 3516 22976 3568 22982
rect 3516 22918 3568 22924
rect 3332 22704 3384 22710
rect 3332 22646 3384 22652
rect 3344 22574 3372 22646
rect 3528 22574 3556 22918
rect 3332 22568 3384 22574
rect 3332 22510 3384 22516
rect 3516 22568 3568 22574
rect 3516 22510 3568 22516
rect 3240 21480 3292 21486
rect 3240 21422 3292 21428
rect 3252 20398 3280 21422
rect 3240 20392 3292 20398
rect 3240 20334 3292 20340
rect 3252 19990 3280 20334
rect 3240 19984 3292 19990
rect 3240 19926 3292 19932
rect 3424 19712 3476 19718
rect 3424 19654 3476 19660
rect 3240 19304 3292 19310
rect 3240 19246 3292 19252
rect 3332 19304 3384 19310
rect 3332 19246 3384 19252
rect 3252 18970 3280 19246
rect 3240 18964 3292 18970
rect 3240 18906 3292 18912
rect 3344 18834 3372 19246
rect 3436 18902 3464 19654
rect 3424 18896 3476 18902
rect 3424 18838 3476 18844
rect 3332 18828 3384 18834
rect 3332 18770 3384 18776
rect 3516 18828 3568 18834
rect 3516 18770 3568 18776
rect 3528 18222 3556 18770
rect 3516 18216 3568 18222
rect 3516 18158 3568 18164
rect 3516 18080 3568 18086
rect 3516 18022 3568 18028
rect 3424 17128 3476 17134
rect 3424 17070 3476 17076
rect 3330 16688 3386 16697
rect 3330 16623 3332 16632
rect 3384 16623 3386 16632
rect 3332 16594 3384 16600
rect 3148 16244 3200 16250
rect 3148 16186 3200 16192
rect 3436 16114 3464 17070
rect 3528 16590 3556 18022
rect 3516 16584 3568 16590
rect 3516 16526 3568 16532
rect 3424 16108 3476 16114
rect 3424 16050 3476 16056
rect 2780 15564 2832 15570
rect 2780 15506 2832 15512
rect 2688 15496 2740 15502
rect 2688 15438 2740 15444
rect 2502 14784 2558 14793
rect 2502 14719 2558 14728
rect 2516 14482 2544 14719
rect 2504 14476 2556 14482
rect 2504 14418 2556 14424
rect 2700 13326 2728 15438
rect 2792 15162 2820 15506
rect 3240 15360 3292 15366
rect 3240 15302 3292 15308
rect 2780 15156 2832 15162
rect 2780 15098 2832 15104
rect 3252 14482 3280 15302
rect 3240 14476 3292 14482
rect 3240 14418 3292 14424
rect 2964 13728 3016 13734
rect 2964 13670 3016 13676
rect 2976 13462 3004 13670
rect 2964 13456 3016 13462
rect 2964 13398 3016 13404
rect 2780 13388 2832 13394
rect 3252 13376 3280 14418
rect 3436 14278 3464 16050
rect 3528 15434 3556 16526
rect 3516 15428 3568 15434
rect 3516 15370 3568 15376
rect 3424 14272 3476 14278
rect 3424 14214 3476 14220
rect 3332 13388 3384 13394
rect 3252 13348 3332 13376
rect 2780 13330 2832 13336
rect 3332 13330 3384 13336
rect 2688 13320 2740 13326
rect 2688 13262 2740 13268
rect 2792 12986 2820 13330
rect 3436 13258 3464 14214
rect 3424 13252 3476 13258
rect 3424 13194 3476 13200
rect 2780 12980 2832 12986
rect 2780 12922 2832 12928
rect 2872 12844 2924 12850
rect 2872 12786 2924 12792
rect 2044 12300 2096 12306
rect 2044 12242 2096 12248
rect 2320 12300 2372 12306
rect 2320 12242 2372 12248
rect 2332 12102 2360 12242
rect 2320 12096 2372 12102
rect 2320 12038 2372 12044
rect 2332 11218 2360 12038
rect 2320 11212 2372 11218
rect 2320 11154 2372 11160
rect 2332 9518 2360 11154
rect 2504 10804 2556 10810
rect 2504 10746 2556 10752
rect 2516 10130 2544 10746
rect 2884 10674 2912 12786
rect 3516 12776 3568 12782
rect 3516 12718 3568 12724
rect 3528 11762 3556 12718
rect 3516 11756 3568 11762
rect 3516 11698 3568 11704
rect 3332 11688 3384 11694
rect 3332 11630 3384 11636
rect 3240 11212 3292 11218
rect 3240 11154 3292 11160
rect 3252 10810 3280 11154
rect 3344 11150 3372 11630
rect 3332 11144 3384 11150
rect 3332 11086 3384 11092
rect 3240 10804 3292 10810
rect 3240 10746 3292 10752
rect 2872 10668 2924 10674
rect 2872 10610 2924 10616
rect 2778 10160 2834 10169
rect 2504 10124 2556 10130
rect 2778 10095 2834 10104
rect 2504 10066 2556 10072
rect 2792 10062 2820 10095
rect 2780 10056 2832 10062
rect 2780 9998 2832 10004
rect 2320 9512 2372 9518
rect 2320 9454 2372 9460
rect 2332 7342 2360 9454
rect 2780 8492 2832 8498
rect 2780 8434 2832 8440
rect 2504 7880 2556 7886
rect 2504 7822 2556 7828
rect 2320 7336 2372 7342
rect 2320 7278 2372 7284
rect 2332 5166 2360 7278
rect 2516 6662 2544 7822
rect 2792 6866 2820 8434
rect 2780 6860 2832 6866
rect 2780 6802 2832 6808
rect 2884 6798 2912 10610
rect 2964 10600 3016 10606
rect 2964 10542 3016 10548
rect 2976 9178 3004 10542
rect 3528 10470 3556 11698
rect 3620 10538 3648 35119
rect 3804 34746 3832 35566
rect 4172 35494 4200 35566
rect 4160 35488 4212 35494
rect 4160 35430 4212 35436
rect 4172 35154 4200 35430
rect 5000 35154 5028 36042
rect 4160 35148 4212 35154
rect 4160 35090 4212 35096
rect 4988 35148 5040 35154
rect 4988 35090 5040 35096
rect 4220 34844 4516 34864
rect 4276 34842 4300 34844
rect 4356 34842 4380 34844
rect 4436 34842 4460 34844
rect 4298 34790 4300 34842
rect 4362 34790 4374 34842
rect 4436 34790 4438 34842
rect 4276 34788 4300 34790
rect 4356 34788 4380 34790
rect 4436 34788 4460 34790
rect 4220 34768 4516 34788
rect 3792 34740 3844 34746
rect 3792 34682 3844 34688
rect 3700 34060 3752 34066
rect 3700 34002 3752 34008
rect 3712 33454 3740 34002
rect 3804 33522 3832 34682
rect 4160 34536 4212 34542
rect 4160 34478 4212 34484
rect 4172 34134 4200 34478
rect 4712 34468 4764 34474
rect 4712 34410 4764 34416
rect 4160 34128 4212 34134
rect 4160 34070 4212 34076
rect 4620 33992 4672 33998
rect 4620 33934 4672 33940
rect 4220 33756 4516 33776
rect 4276 33754 4300 33756
rect 4356 33754 4380 33756
rect 4436 33754 4460 33756
rect 4298 33702 4300 33754
rect 4362 33702 4374 33754
rect 4436 33702 4438 33754
rect 4276 33700 4300 33702
rect 4356 33700 4380 33702
rect 4436 33700 4460 33702
rect 4220 33680 4516 33700
rect 3792 33516 3844 33522
rect 3792 33458 3844 33464
rect 3700 33448 3752 33454
rect 3700 33390 3752 33396
rect 3712 30802 3740 33390
rect 4632 33046 4660 33934
rect 4724 33454 4752 34410
rect 5080 33992 5132 33998
rect 5080 33934 5132 33940
rect 5092 33658 5120 33934
rect 5080 33652 5132 33658
rect 5080 33594 5132 33600
rect 4712 33448 4764 33454
rect 4712 33390 4764 33396
rect 5092 33046 5120 33594
rect 4620 33040 4672 33046
rect 4620 32982 4672 32988
rect 5080 33040 5132 33046
rect 5080 32982 5132 32988
rect 4712 32972 4764 32978
rect 4712 32914 4764 32920
rect 4988 32972 5040 32978
rect 4988 32914 5040 32920
rect 4068 32904 4120 32910
rect 4068 32846 4120 32852
rect 4080 32434 4108 32846
rect 4220 32668 4516 32688
rect 4276 32666 4300 32668
rect 4356 32666 4380 32668
rect 4436 32666 4460 32668
rect 4298 32614 4300 32666
rect 4362 32614 4374 32666
rect 4436 32614 4438 32666
rect 4276 32612 4300 32614
rect 4356 32612 4380 32614
rect 4436 32612 4460 32614
rect 4220 32592 4516 32612
rect 4160 32496 4212 32502
rect 4160 32438 4212 32444
rect 4620 32496 4672 32502
rect 4620 32438 4672 32444
rect 4068 32428 4120 32434
rect 4068 32370 4120 32376
rect 4080 32042 4108 32370
rect 4172 32366 4200 32438
rect 4160 32360 4212 32366
rect 4160 32302 4212 32308
rect 3988 32026 4108 32042
rect 3988 32020 4120 32026
rect 3988 32014 4068 32020
rect 3988 31278 4016 32014
rect 4068 31962 4120 31968
rect 4068 31884 4120 31890
rect 4068 31826 4120 31832
rect 4080 31482 4108 31826
rect 4220 31580 4516 31600
rect 4276 31578 4300 31580
rect 4356 31578 4380 31580
rect 4436 31578 4460 31580
rect 4298 31526 4300 31578
rect 4362 31526 4374 31578
rect 4436 31526 4438 31578
rect 4276 31524 4300 31526
rect 4356 31524 4380 31526
rect 4436 31524 4460 31526
rect 4220 31504 4516 31524
rect 4068 31476 4120 31482
rect 4068 31418 4120 31424
rect 4632 31346 4660 32438
rect 4724 32298 4752 32914
rect 5000 32502 5028 32914
rect 4988 32496 5040 32502
rect 4988 32438 5040 32444
rect 5092 32366 5120 32982
rect 5080 32360 5132 32366
rect 5080 32302 5132 32308
rect 4712 32292 4764 32298
rect 4712 32234 4764 32240
rect 4620 31340 4672 31346
rect 4620 31282 4672 31288
rect 3976 31272 4028 31278
rect 3976 31214 4028 31220
rect 3700 30796 3752 30802
rect 3700 30738 3752 30744
rect 4068 30796 4120 30802
rect 4068 30738 4120 30744
rect 3712 30326 3740 30738
rect 3700 30320 3752 30326
rect 3700 30262 3752 30268
rect 4080 30190 4108 30738
rect 4220 30492 4516 30512
rect 4276 30490 4300 30492
rect 4356 30490 4380 30492
rect 4436 30490 4460 30492
rect 4298 30438 4300 30490
rect 4362 30438 4374 30490
rect 4436 30438 4438 30490
rect 4276 30436 4300 30438
rect 4356 30436 4380 30438
rect 4436 30436 4460 30438
rect 4220 30416 4516 30436
rect 4632 30258 4660 31282
rect 4724 31278 4752 32234
rect 4712 31272 4764 31278
rect 4712 31214 4764 31220
rect 4896 31272 4948 31278
rect 4896 31214 4948 31220
rect 4712 30592 4764 30598
rect 4712 30534 4764 30540
rect 4620 30252 4672 30258
rect 4620 30194 4672 30200
rect 4068 30184 4120 30190
rect 4068 30126 4120 30132
rect 4528 30184 4580 30190
rect 4528 30126 4580 30132
rect 4540 29782 4568 30126
rect 4528 29776 4580 29782
rect 4528 29718 4580 29724
rect 4632 29714 4660 30194
rect 4724 30190 4752 30534
rect 4712 30184 4764 30190
rect 4712 30126 4764 30132
rect 4620 29708 4672 29714
rect 4620 29650 4672 29656
rect 3976 29504 4028 29510
rect 3976 29446 4028 29452
rect 3884 27872 3936 27878
rect 3884 27814 3936 27820
rect 3896 26926 3924 27814
rect 3884 26920 3936 26926
rect 3884 26862 3936 26868
rect 3988 26450 4016 29446
rect 4220 29404 4516 29424
rect 4276 29402 4300 29404
rect 4356 29402 4380 29404
rect 4436 29402 4460 29404
rect 4298 29350 4300 29402
rect 4362 29350 4374 29402
rect 4436 29350 4438 29402
rect 4276 29348 4300 29350
rect 4356 29348 4380 29350
rect 4436 29348 4460 29350
rect 4220 29328 4516 29348
rect 4632 29102 4660 29650
rect 4908 29646 4936 31214
rect 5080 30728 5132 30734
rect 5080 30670 5132 30676
rect 4896 29640 4948 29646
rect 4896 29582 4948 29588
rect 4804 29572 4856 29578
rect 4804 29514 4856 29520
rect 4816 29102 4844 29514
rect 4160 29096 4212 29102
rect 4160 29038 4212 29044
rect 4620 29096 4672 29102
rect 4620 29038 4672 29044
rect 4804 29096 4856 29102
rect 4804 29038 4856 29044
rect 4172 28762 4200 29038
rect 4908 29034 4936 29582
rect 5092 29306 5120 30670
rect 5080 29300 5132 29306
rect 5080 29242 5132 29248
rect 4896 29028 4948 29034
rect 4896 28970 4948 28976
rect 4160 28756 4212 28762
rect 4160 28698 4212 28704
rect 5092 28558 5120 29242
rect 4712 28552 4764 28558
rect 4712 28494 4764 28500
rect 5080 28552 5132 28558
rect 5080 28494 5132 28500
rect 4620 28416 4672 28422
rect 4620 28358 4672 28364
rect 4220 28316 4516 28336
rect 4276 28314 4300 28316
rect 4356 28314 4380 28316
rect 4436 28314 4460 28316
rect 4298 28262 4300 28314
rect 4362 28262 4374 28314
rect 4436 28262 4438 28314
rect 4276 28260 4300 28262
rect 4356 28260 4380 28262
rect 4436 28260 4460 28262
rect 4220 28240 4516 28260
rect 4068 28144 4120 28150
rect 4068 28086 4120 28092
rect 4080 27334 4108 28086
rect 4436 28008 4488 28014
rect 4488 27968 4568 27996
rect 4436 27950 4488 27956
rect 4540 27418 4568 27968
rect 4632 27538 4660 28358
rect 4620 27532 4672 27538
rect 4620 27474 4672 27480
rect 4540 27390 4660 27418
rect 4068 27328 4120 27334
rect 4068 27270 4120 27276
rect 4080 26926 4108 27270
rect 4220 27228 4516 27248
rect 4276 27226 4300 27228
rect 4356 27226 4380 27228
rect 4436 27226 4460 27228
rect 4298 27174 4300 27226
rect 4362 27174 4374 27226
rect 4436 27174 4438 27226
rect 4276 27172 4300 27174
rect 4356 27172 4380 27174
rect 4436 27172 4460 27174
rect 4220 27152 4516 27172
rect 4068 26920 4120 26926
rect 4068 26862 4120 26868
rect 3976 26444 4028 26450
rect 3976 26386 4028 26392
rect 4220 26140 4516 26160
rect 4276 26138 4300 26140
rect 4356 26138 4380 26140
rect 4436 26138 4460 26140
rect 4298 26086 4300 26138
rect 4362 26086 4374 26138
rect 4436 26086 4438 26138
rect 4276 26084 4300 26086
rect 4356 26084 4380 26086
rect 4436 26084 4460 26086
rect 4220 26064 4516 26084
rect 4632 26042 4660 27390
rect 4724 26994 4752 28494
rect 5092 27470 5120 28494
rect 5080 27464 5132 27470
rect 5080 27406 5132 27412
rect 4804 27056 4856 27062
rect 4804 26998 4856 27004
rect 4712 26988 4764 26994
rect 4712 26930 4764 26936
rect 4816 26450 4844 26998
rect 4988 26784 5040 26790
rect 4988 26726 5040 26732
rect 4804 26444 4856 26450
rect 4804 26386 4856 26392
rect 4620 26036 4672 26042
rect 4620 25978 4672 25984
rect 4632 25838 4660 25978
rect 4160 25832 4212 25838
rect 4160 25774 4212 25780
rect 4620 25832 4672 25838
rect 4620 25774 4672 25780
rect 4068 25696 4120 25702
rect 3974 25664 4030 25673
rect 4068 25638 4120 25644
rect 3974 25599 4030 25608
rect 3988 25226 4016 25599
rect 4080 25430 4108 25638
rect 4172 25498 4200 25774
rect 4160 25492 4212 25498
rect 4160 25434 4212 25440
rect 4068 25424 4120 25430
rect 4068 25366 4120 25372
rect 3976 25220 4028 25226
rect 3976 25162 4028 25168
rect 4220 25052 4516 25072
rect 4276 25050 4300 25052
rect 4356 25050 4380 25052
rect 4436 25050 4460 25052
rect 4298 24998 4300 25050
rect 4362 24998 4374 25050
rect 4436 24998 4438 25050
rect 4276 24996 4300 24998
rect 4356 24996 4380 24998
rect 4436 24996 4460 24998
rect 4220 24976 4516 24996
rect 5000 24818 5028 26726
rect 5092 26382 5120 27406
rect 5080 26376 5132 26382
rect 5080 26318 5132 26324
rect 5080 26240 5132 26246
rect 5080 26182 5132 26188
rect 5092 25294 5120 26182
rect 5080 25288 5132 25294
rect 5080 25230 5132 25236
rect 4988 24812 5040 24818
rect 4988 24754 5040 24760
rect 4528 24268 4580 24274
rect 4580 24228 4660 24256
rect 4528 24210 4580 24216
rect 3700 24064 3752 24070
rect 3700 24006 3752 24012
rect 3712 23730 3740 24006
rect 4220 23964 4516 23984
rect 4276 23962 4300 23964
rect 4356 23962 4380 23964
rect 4436 23962 4460 23964
rect 4298 23910 4300 23962
rect 4362 23910 4374 23962
rect 4436 23910 4438 23962
rect 4276 23908 4300 23910
rect 4356 23908 4380 23910
rect 4436 23908 4460 23910
rect 4220 23888 4516 23908
rect 3700 23724 3752 23730
rect 3700 23666 3752 23672
rect 4220 22876 4516 22896
rect 4276 22874 4300 22876
rect 4356 22874 4380 22876
rect 4436 22874 4460 22876
rect 4298 22822 4300 22874
rect 4362 22822 4374 22874
rect 4436 22822 4438 22874
rect 4276 22820 4300 22822
rect 4356 22820 4380 22822
rect 4436 22820 4460 22822
rect 4220 22800 4516 22820
rect 4632 22642 4660 24228
rect 4712 23520 4764 23526
rect 4712 23462 4764 23468
rect 4988 23520 5040 23526
rect 4988 23462 5040 23468
rect 4724 23050 4752 23462
rect 4896 23180 4948 23186
rect 4896 23122 4948 23128
rect 4712 23044 4764 23050
rect 4712 22986 4764 22992
rect 4620 22636 4672 22642
rect 4620 22578 4672 22584
rect 3792 22568 3844 22574
rect 3792 22510 3844 22516
rect 4712 22568 4764 22574
rect 4712 22510 4764 22516
rect 3700 22500 3752 22506
rect 3700 22442 3752 22448
rect 3712 22098 3740 22442
rect 3700 22092 3752 22098
rect 3700 22034 3752 22040
rect 3804 21962 3832 22510
rect 4068 22092 4120 22098
rect 4068 22034 4120 22040
rect 4620 22092 4672 22098
rect 4620 22034 4672 22040
rect 3792 21956 3844 21962
rect 3792 21898 3844 21904
rect 3804 21418 3832 21898
rect 4080 21690 4108 22034
rect 4220 21788 4516 21808
rect 4276 21786 4300 21788
rect 4356 21786 4380 21788
rect 4436 21786 4460 21788
rect 4298 21734 4300 21786
rect 4362 21734 4374 21786
rect 4436 21734 4438 21786
rect 4276 21732 4300 21734
rect 4356 21732 4380 21734
rect 4436 21732 4460 21734
rect 4220 21712 4516 21732
rect 4068 21684 4120 21690
rect 4068 21626 4120 21632
rect 3792 21412 3844 21418
rect 3792 21354 3844 21360
rect 4220 20700 4516 20720
rect 4276 20698 4300 20700
rect 4356 20698 4380 20700
rect 4436 20698 4460 20700
rect 4298 20646 4300 20698
rect 4362 20646 4374 20698
rect 4436 20646 4438 20698
rect 4276 20644 4300 20646
rect 4356 20644 4380 20646
rect 4436 20644 4460 20646
rect 4220 20624 4516 20644
rect 4632 20534 4660 22034
rect 4724 21078 4752 22510
rect 4908 22234 4936 23122
rect 5000 23050 5028 23462
rect 4988 23044 5040 23050
rect 4988 22986 5040 22992
rect 4896 22228 4948 22234
rect 4896 22170 4948 22176
rect 4896 22024 4948 22030
rect 4896 21966 4948 21972
rect 4804 21412 4856 21418
rect 4804 21354 4856 21360
rect 4712 21072 4764 21078
rect 4712 21014 4764 21020
rect 4816 21010 4844 21354
rect 4804 21004 4856 21010
rect 4804 20946 4856 20952
rect 4620 20528 4672 20534
rect 4620 20470 4672 20476
rect 3884 19916 3936 19922
rect 3884 19858 3936 19864
rect 3700 19304 3752 19310
rect 3698 19272 3700 19281
rect 3752 19272 3754 19281
rect 3698 19207 3754 19216
rect 3896 18630 3924 19858
rect 4220 19612 4516 19632
rect 4276 19610 4300 19612
rect 4356 19610 4380 19612
rect 4436 19610 4460 19612
rect 4298 19558 4300 19610
rect 4362 19558 4374 19610
rect 4436 19558 4438 19610
rect 4276 19556 4300 19558
rect 4356 19556 4380 19558
rect 4436 19556 4460 19558
rect 4220 19536 4516 19556
rect 4068 19508 4120 19514
rect 4068 19450 4120 19456
rect 4080 19417 4108 19450
rect 4066 19408 4122 19417
rect 4066 19343 4122 19352
rect 4908 19310 4936 21966
rect 4988 21888 5040 21894
rect 4988 21830 5040 21836
rect 5000 21486 5028 21830
rect 4988 21480 5040 21486
rect 4988 21422 5040 21428
rect 4252 19304 4304 19310
rect 4252 19246 4304 19252
rect 4896 19304 4948 19310
rect 4896 19246 4948 19252
rect 3976 19168 4028 19174
rect 3976 19110 4028 19116
rect 3884 18624 3936 18630
rect 3884 18566 3936 18572
rect 3896 17814 3924 18566
rect 3884 17808 3936 17814
rect 3884 17750 3936 17756
rect 3988 17746 4016 19110
rect 4264 18766 4292 19246
rect 4252 18760 4304 18766
rect 4252 18702 4304 18708
rect 4220 18524 4516 18544
rect 4276 18522 4300 18524
rect 4356 18522 4380 18524
rect 4436 18522 4460 18524
rect 4298 18470 4300 18522
rect 4362 18470 4374 18522
rect 4436 18470 4438 18522
rect 4276 18468 4300 18470
rect 4356 18468 4380 18470
rect 4436 18468 4460 18470
rect 4220 18448 4516 18468
rect 4620 18352 4672 18358
rect 4620 18294 4672 18300
rect 3976 17740 4028 17746
rect 3976 17682 4028 17688
rect 3976 17536 4028 17542
rect 3976 17478 4028 17484
rect 3988 17134 4016 17478
rect 4220 17436 4516 17456
rect 4276 17434 4300 17436
rect 4356 17434 4380 17436
rect 4436 17434 4460 17436
rect 4298 17382 4300 17434
rect 4362 17382 4374 17434
rect 4436 17382 4438 17434
rect 4276 17380 4300 17382
rect 4356 17380 4380 17382
rect 4436 17380 4460 17382
rect 4220 17360 4516 17380
rect 4632 17202 4660 18294
rect 4712 18148 4764 18154
rect 4712 18090 4764 18096
rect 4724 17338 4752 18090
rect 4896 17740 4948 17746
rect 4896 17682 4948 17688
rect 4712 17332 4764 17338
rect 4712 17274 4764 17280
rect 4724 17202 4752 17274
rect 4620 17196 4672 17202
rect 4620 17138 4672 17144
rect 4712 17196 4764 17202
rect 4712 17138 4764 17144
rect 4908 17134 4936 17682
rect 3976 17128 4028 17134
rect 3976 17070 4028 17076
rect 4896 17128 4948 17134
rect 4896 17070 4948 17076
rect 4804 16788 4856 16794
rect 4804 16730 4856 16736
rect 4434 16688 4490 16697
rect 4434 16623 4490 16632
rect 4448 16590 4476 16623
rect 4436 16584 4488 16590
rect 4436 16526 4488 16532
rect 3976 16516 4028 16522
rect 3976 16458 4028 16464
rect 3988 16250 4016 16458
rect 4068 16448 4120 16454
rect 4066 16416 4068 16425
rect 4120 16416 4122 16425
rect 4066 16351 4122 16360
rect 4220 16348 4516 16368
rect 4276 16346 4300 16348
rect 4356 16346 4380 16348
rect 4436 16346 4460 16348
rect 4298 16294 4300 16346
rect 4362 16294 4374 16346
rect 4436 16294 4438 16346
rect 4276 16292 4300 16294
rect 4356 16292 4380 16294
rect 4436 16292 4460 16294
rect 4220 16272 4516 16292
rect 3976 16244 4028 16250
rect 3976 16186 4028 16192
rect 4816 16114 4844 16730
rect 4804 16108 4856 16114
rect 4804 16050 4856 16056
rect 3700 16040 3752 16046
rect 3700 15982 3752 15988
rect 3712 15706 3740 15982
rect 3792 15904 3844 15910
rect 3792 15846 3844 15852
rect 3700 15700 3752 15706
rect 3700 15642 3752 15648
rect 3804 15502 3832 15846
rect 3884 15564 3936 15570
rect 3884 15506 3936 15512
rect 3792 15496 3844 15502
rect 3792 15438 3844 15444
rect 3896 14006 3924 15506
rect 4068 15496 4120 15502
rect 4068 15438 4120 15444
rect 4804 15496 4856 15502
rect 4804 15438 4856 15444
rect 4080 14958 4108 15438
rect 4220 15260 4516 15280
rect 4276 15258 4300 15260
rect 4356 15258 4380 15260
rect 4436 15258 4460 15260
rect 4298 15206 4300 15258
rect 4362 15206 4374 15258
rect 4436 15206 4438 15258
rect 4276 15204 4300 15206
rect 4356 15204 4380 15206
rect 4436 15204 4460 15206
rect 4220 15184 4516 15204
rect 4068 14952 4120 14958
rect 4068 14894 4120 14900
rect 4620 14952 4672 14958
rect 4620 14894 4672 14900
rect 3976 14612 4028 14618
rect 3976 14554 4028 14560
rect 3884 14000 3936 14006
rect 3884 13942 3936 13948
rect 3792 12776 3844 12782
rect 3792 12718 3844 12724
rect 3804 12374 3832 12718
rect 3792 12368 3844 12374
rect 3792 12310 3844 12316
rect 3896 11218 3924 13942
rect 3988 13870 4016 14554
rect 4068 14408 4120 14414
rect 4068 14350 4120 14356
rect 3976 13864 4028 13870
rect 4080 13852 4108 14350
rect 4220 14172 4516 14192
rect 4276 14170 4300 14172
rect 4356 14170 4380 14172
rect 4436 14170 4460 14172
rect 4298 14118 4300 14170
rect 4362 14118 4374 14170
rect 4436 14118 4438 14170
rect 4276 14116 4300 14118
rect 4356 14116 4380 14118
rect 4436 14116 4460 14118
rect 4220 14096 4516 14116
rect 4632 13938 4660 14894
rect 4816 14550 4844 15438
rect 4804 14544 4856 14550
rect 4804 14486 4856 14492
rect 5092 14414 5120 25230
rect 5184 16046 5212 37742
rect 5540 37392 5592 37398
rect 5540 37334 5592 37340
rect 5552 36786 5580 37334
rect 5644 36854 5672 38168
rect 6104 37670 6132 38286
rect 7472 37800 7524 37806
rect 7472 37742 7524 37748
rect 7748 37800 7800 37806
rect 7748 37742 7800 37748
rect 6092 37664 6144 37670
rect 6092 37606 6144 37612
rect 6920 37664 6972 37670
rect 6920 37606 6972 37612
rect 6104 37262 6132 37606
rect 6092 37256 6144 37262
rect 6092 37198 6144 37204
rect 5632 36848 5684 36854
rect 5632 36790 5684 36796
rect 5540 36780 5592 36786
rect 5540 36722 5592 36728
rect 5816 36644 5868 36650
rect 5816 36586 5868 36592
rect 5724 36304 5776 36310
rect 5724 36246 5776 36252
rect 5540 36236 5592 36242
rect 5540 36178 5592 36184
rect 5356 36100 5408 36106
rect 5356 36042 5408 36048
rect 5368 35630 5396 36042
rect 5552 35698 5580 36178
rect 5540 35692 5592 35698
rect 5540 35634 5592 35640
rect 5356 35624 5408 35630
rect 5356 35566 5408 35572
rect 5368 34542 5396 35566
rect 5632 34944 5684 34950
rect 5632 34886 5684 34892
rect 5356 34536 5408 34542
rect 5356 34478 5408 34484
rect 5644 34134 5672 34886
rect 5736 34678 5764 36246
rect 5828 35766 5856 36586
rect 5816 35760 5868 35766
rect 5816 35702 5868 35708
rect 6104 35086 6132 37198
rect 6932 36718 6960 37606
rect 7196 37120 7248 37126
rect 7196 37062 7248 37068
rect 7208 36718 7236 37062
rect 6920 36712 6972 36718
rect 6920 36654 6972 36660
rect 7196 36712 7248 36718
rect 7196 36654 7248 36660
rect 7208 36310 7236 36654
rect 7484 36378 7512 37742
rect 7472 36372 7524 36378
rect 7472 36314 7524 36320
rect 7196 36304 7248 36310
rect 7196 36246 7248 36252
rect 6736 36236 6788 36242
rect 6736 36178 6788 36184
rect 7380 36236 7432 36242
rect 7380 36178 7432 36184
rect 6748 35494 6776 36178
rect 6828 35624 6880 35630
rect 6828 35566 6880 35572
rect 6736 35488 6788 35494
rect 6736 35430 6788 35436
rect 6644 35216 6696 35222
rect 6644 35158 6696 35164
rect 6092 35080 6144 35086
rect 6092 35022 6144 35028
rect 5908 34944 5960 34950
rect 5908 34886 5960 34892
rect 5724 34672 5776 34678
rect 5724 34614 5776 34620
rect 5920 34542 5948 34886
rect 5908 34536 5960 34542
rect 5908 34478 5960 34484
rect 5724 34400 5776 34406
rect 5724 34342 5776 34348
rect 5632 34128 5684 34134
rect 5632 34070 5684 34076
rect 5736 33862 5764 34342
rect 5908 33992 5960 33998
rect 5908 33934 5960 33940
rect 5724 33856 5776 33862
rect 5724 33798 5776 33804
rect 5736 32366 5764 33798
rect 5920 32570 5948 33934
rect 6104 33930 6132 35022
rect 6656 34066 6684 35158
rect 6748 34542 6776 35430
rect 6840 35154 6868 35566
rect 6828 35148 6880 35154
rect 6828 35090 6880 35096
rect 7392 35018 7420 36178
rect 7472 36168 7524 36174
rect 7472 36110 7524 36116
rect 7484 35698 7512 36110
rect 7760 35698 7788 37742
rect 7840 36372 7892 36378
rect 7840 36314 7892 36320
rect 7472 35692 7524 35698
rect 7472 35634 7524 35640
rect 7748 35692 7800 35698
rect 7748 35634 7800 35640
rect 7484 35154 7512 35634
rect 7472 35148 7524 35154
rect 7472 35090 7524 35096
rect 7380 35012 7432 35018
rect 7380 34954 7432 34960
rect 7392 34542 7420 34954
rect 6736 34536 6788 34542
rect 6736 34478 6788 34484
rect 7380 34536 7432 34542
rect 7380 34478 7432 34484
rect 6644 34060 6696 34066
rect 6644 34002 6696 34008
rect 6920 34060 6972 34066
rect 6920 34002 6972 34008
rect 7196 34060 7248 34066
rect 7196 34002 7248 34008
rect 6092 33924 6144 33930
rect 6092 33866 6144 33872
rect 6000 33108 6052 33114
rect 6000 33050 6052 33056
rect 5908 32564 5960 32570
rect 5908 32506 5960 32512
rect 5724 32360 5776 32366
rect 5724 32302 5776 32308
rect 6012 31754 6040 33050
rect 6104 32910 6132 33866
rect 6932 33674 6960 34002
rect 7104 33992 7156 33998
rect 7104 33934 7156 33940
rect 6748 33646 6960 33674
rect 6748 33522 6776 33646
rect 6736 33516 6788 33522
rect 6736 33458 6788 33464
rect 6920 33516 6972 33522
rect 6920 33458 6972 33464
rect 6092 32904 6144 32910
rect 6092 32846 6144 32852
rect 6460 32904 6512 32910
rect 6460 32846 6512 32852
rect 6736 32904 6788 32910
rect 6736 32846 6788 32852
rect 6000 31748 6052 31754
rect 6000 31690 6052 31696
rect 5632 31680 5684 31686
rect 5632 31622 5684 31628
rect 5644 30802 5672 31622
rect 5816 31136 5868 31142
rect 5816 31078 5868 31084
rect 5632 30796 5684 30802
rect 5632 30738 5684 30744
rect 5828 30190 5856 31078
rect 5816 30184 5868 30190
rect 5816 30126 5868 30132
rect 5448 30116 5500 30122
rect 5448 30058 5500 30064
rect 5460 29714 5488 30058
rect 5540 29844 5592 29850
rect 5540 29786 5592 29792
rect 5448 29708 5500 29714
rect 5448 29650 5500 29656
rect 5356 28620 5408 28626
rect 5460 28608 5488 29650
rect 5552 28694 5580 29786
rect 5828 29646 5856 30126
rect 5816 29640 5868 29646
rect 5816 29582 5868 29588
rect 5632 29572 5684 29578
rect 5632 29514 5684 29520
rect 5540 28688 5592 28694
rect 5540 28630 5592 28636
rect 5408 28580 5488 28608
rect 5356 28562 5408 28568
rect 5460 27946 5488 28580
rect 5644 28014 5672 29514
rect 5724 28552 5776 28558
rect 5724 28494 5776 28500
rect 5736 28150 5764 28494
rect 5724 28144 5776 28150
rect 5724 28086 5776 28092
rect 5828 28014 5856 29582
rect 5632 28008 5684 28014
rect 5632 27950 5684 27956
rect 5816 28008 5868 28014
rect 5816 27950 5868 27956
rect 5448 27940 5500 27946
rect 5448 27882 5500 27888
rect 6012 27334 6040 31690
rect 6092 31680 6144 31686
rect 6092 31622 6144 31628
rect 6104 31278 6132 31622
rect 6472 31278 6500 32846
rect 6748 32434 6776 32846
rect 6736 32428 6788 32434
rect 6736 32370 6788 32376
rect 6932 32366 6960 33458
rect 7116 33454 7144 33934
rect 7208 33658 7236 34002
rect 7852 33998 7880 36314
rect 7840 33992 7892 33998
rect 7840 33934 7892 33940
rect 7196 33652 7248 33658
rect 7196 33594 7248 33600
rect 7104 33448 7156 33454
rect 7104 33390 7156 33396
rect 7116 32774 7144 33390
rect 7208 33318 7236 33594
rect 7380 33380 7432 33386
rect 7380 33322 7432 33328
rect 7196 33312 7248 33318
rect 7196 33254 7248 33260
rect 7104 32768 7156 32774
rect 7104 32710 7156 32716
rect 7392 32434 7420 33322
rect 7380 32428 7432 32434
rect 7380 32370 7432 32376
rect 6920 32360 6972 32366
rect 6920 32302 6972 32308
rect 6552 32292 6604 32298
rect 6552 32234 6604 32240
rect 7288 32292 7340 32298
rect 7288 32234 7340 32240
rect 6092 31272 6144 31278
rect 6092 31214 6144 31220
rect 6460 31272 6512 31278
rect 6460 31214 6512 31220
rect 6564 29850 6592 32234
rect 7196 31952 7248 31958
rect 7196 31894 7248 31900
rect 7208 30870 7236 31894
rect 7300 31890 7328 32234
rect 7288 31884 7340 31890
rect 7288 31826 7340 31832
rect 7380 31204 7432 31210
rect 7380 31146 7432 31152
rect 7196 30864 7248 30870
rect 7196 30806 7248 30812
rect 7012 30728 7064 30734
rect 7012 30670 7064 30676
rect 7024 30190 7052 30670
rect 7104 30660 7156 30666
rect 7104 30602 7156 30608
rect 7012 30184 7064 30190
rect 7012 30126 7064 30132
rect 6552 29844 6604 29850
rect 6552 29786 6604 29792
rect 7024 29714 7052 30126
rect 7012 29708 7064 29714
rect 7012 29650 7064 29656
rect 7012 29232 7064 29238
rect 7012 29174 7064 29180
rect 7024 29102 7052 29174
rect 7012 29096 7064 29102
rect 7012 29038 7064 29044
rect 6920 29028 6972 29034
rect 6920 28970 6972 28976
rect 6932 28762 6960 28970
rect 6920 28756 6972 28762
rect 6920 28698 6972 28704
rect 7116 28150 7144 30602
rect 7392 29646 7420 31146
rect 7656 30796 7708 30802
rect 7656 30738 7708 30744
rect 7840 30796 7892 30802
rect 7840 30738 7892 30744
rect 7668 30326 7696 30738
rect 7656 30320 7708 30326
rect 7656 30262 7708 30268
rect 7852 30258 7880 30738
rect 7840 30252 7892 30258
rect 7840 30194 7892 30200
rect 7380 29640 7432 29646
rect 7380 29582 7432 29588
rect 7392 28694 7420 29582
rect 7748 29504 7800 29510
rect 7748 29446 7800 29452
rect 7564 29096 7616 29102
rect 7564 29038 7616 29044
rect 7380 28688 7432 28694
rect 7380 28630 7432 28636
rect 7104 28144 7156 28150
rect 7104 28086 7156 28092
rect 6828 28008 6880 28014
rect 6828 27950 6880 27956
rect 6840 27470 6868 27950
rect 7116 27674 7144 28086
rect 7104 27668 7156 27674
rect 7104 27610 7156 27616
rect 7576 27538 7604 29038
rect 7760 28966 7788 29446
rect 7748 28960 7800 28966
rect 7748 28902 7800 28908
rect 7564 27532 7616 27538
rect 7564 27474 7616 27480
rect 6828 27464 6880 27470
rect 6828 27406 6880 27412
rect 7380 27464 7432 27470
rect 7380 27406 7432 27412
rect 6000 27328 6052 27334
rect 6000 27270 6052 27276
rect 6460 27328 6512 27334
rect 6460 27270 6512 27276
rect 5540 26920 5592 26926
rect 5540 26862 5592 26868
rect 5552 25294 5580 26862
rect 6184 26852 6236 26858
rect 6184 26794 6236 26800
rect 5724 25832 5776 25838
rect 5724 25774 5776 25780
rect 5540 25288 5592 25294
rect 5540 25230 5592 25236
rect 5736 24954 5764 25774
rect 5816 25696 5868 25702
rect 5816 25638 5868 25644
rect 5828 25362 5856 25638
rect 5816 25356 5868 25362
rect 6092 25356 6144 25362
rect 5816 25298 5868 25304
rect 6012 25316 6092 25344
rect 5724 24948 5776 24954
rect 5724 24890 5776 24896
rect 5540 24268 5592 24274
rect 5540 24210 5592 24216
rect 5552 23322 5580 24210
rect 5632 23792 5684 23798
rect 5632 23734 5684 23740
rect 5540 23316 5592 23322
rect 5540 23258 5592 23264
rect 5644 22574 5672 23734
rect 5736 23662 5764 24890
rect 5828 24614 5856 25298
rect 5816 24608 5868 24614
rect 5816 24550 5868 24556
rect 5828 24206 5856 24550
rect 5816 24200 5868 24206
rect 5816 24142 5868 24148
rect 5724 23656 5776 23662
rect 5724 23598 5776 23604
rect 6012 23254 6040 25316
rect 6092 25298 6144 25304
rect 6196 24206 6224 26794
rect 6276 24676 6328 24682
rect 6276 24618 6328 24624
rect 6288 24274 6316 24618
rect 6276 24268 6328 24274
rect 6276 24210 6328 24216
rect 6184 24200 6236 24206
rect 6184 24142 6236 24148
rect 6000 23248 6052 23254
rect 6000 23190 6052 23196
rect 6012 22710 6040 23190
rect 6092 23180 6144 23186
rect 6092 23122 6144 23128
rect 6184 23180 6236 23186
rect 6184 23122 6236 23128
rect 6104 22710 6132 23122
rect 6000 22704 6052 22710
rect 6000 22646 6052 22652
rect 6092 22704 6144 22710
rect 6092 22646 6144 22652
rect 6196 22574 6224 23122
rect 5632 22568 5684 22574
rect 5632 22510 5684 22516
rect 6184 22568 6236 22574
rect 6184 22510 6236 22516
rect 6196 22438 6224 22510
rect 5356 22432 5408 22438
rect 5356 22374 5408 22380
rect 6184 22432 6236 22438
rect 6184 22374 6236 22380
rect 5368 22098 5396 22374
rect 5356 22092 5408 22098
rect 5356 22034 5408 22040
rect 5816 22092 5868 22098
rect 6196 22080 6224 22374
rect 6276 22092 6328 22098
rect 6196 22052 6276 22080
rect 5816 22034 5868 22040
rect 6276 22034 6328 22040
rect 5368 20874 5396 22034
rect 5448 21480 5500 21486
rect 5448 21422 5500 21428
rect 5460 21078 5488 21422
rect 5448 21072 5500 21078
rect 5448 21014 5500 21020
rect 5356 20868 5408 20874
rect 5356 20810 5408 20816
rect 5460 20466 5488 21014
rect 5828 20942 5856 22034
rect 6288 21010 6316 22034
rect 6276 21004 6328 21010
rect 6276 20946 6328 20952
rect 5816 20936 5868 20942
rect 5816 20878 5868 20884
rect 5448 20460 5500 20466
rect 5448 20402 5500 20408
rect 5356 20392 5408 20398
rect 5356 20334 5408 20340
rect 5368 19854 5396 20334
rect 5828 19990 5856 20878
rect 6472 20602 6500 27270
rect 6828 26240 6880 26246
rect 6828 26182 6880 26188
rect 6840 25362 6868 26182
rect 7104 25832 7156 25838
rect 7104 25774 7156 25780
rect 7012 25492 7064 25498
rect 7012 25434 7064 25440
rect 6828 25356 6880 25362
rect 6828 25298 6880 25304
rect 6840 23662 6868 25298
rect 7024 24818 7052 25434
rect 7116 25294 7144 25774
rect 7104 25288 7156 25294
rect 7104 25230 7156 25236
rect 7196 25220 7248 25226
rect 7196 25162 7248 25168
rect 7012 24812 7064 24818
rect 7012 24754 7064 24760
rect 7024 24274 7052 24754
rect 7012 24268 7064 24274
rect 7012 24210 7064 24216
rect 6828 23656 6880 23662
rect 6828 23598 6880 23604
rect 7024 22710 7052 24210
rect 7104 22976 7156 22982
rect 7104 22918 7156 22924
rect 7012 22704 7064 22710
rect 7012 22646 7064 22652
rect 6828 22636 6880 22642
rect 6828 22578 6880 22584
rect 6840 21690 6868 22578
rect 7116 22506 7144 22918
rect 7208 22658 7236 25162
rect 7392 24750 7420 27406
rect 7840 26920 7892 26926
rect 7840 26862 7892 26868
rect 7748 26580 7800 26586
rect 7748 26522 7800 26528
rect 7472 25764 7524 25770
rect 7472 25706 7524 25712
rect 7380 24744 7432 24750
rect 7380 24686 7432 24692
rect 7288 23112 7340 23118
rect 7288 23054 7340 23060
rect 7300 22778 7328 23054
rect 7288 22772 7340 22778
rect 7288 22714 7340 22720
rect 7208 22630 7328 22658
rect 7104 22500 7156 22506
rect 7104 22442 7156 22448
rect 7116 22098 7144 22442
rect 7196 22228 7248 22234
rect 7196 22170 7248 22176
rect 6920 22092 6972 22098
rect 6920 22034 6972 22040
rect 7104 22092 7156 22098
rect 7104 22034 7156 22040
rect 6828 21684 6880 21690
rect 6828 21626 6880 21632
rect 6932 21010 6960 22034
rect 7208 21486 7236 22170
rect 7196 21480 7248 21486
rect 7196 21422 7248 21428
rect 6920 21004 6972 21010
rect 6920 20946 6972 20952
rect 6460 20596 6512 20602
rect 6460 20538 6512 20544
rect 6828 20528 6880 20534
rect 6880 20476 6960 20482
rect 6828 20470 6960 20476
rect 6840 20454 6960 20470
rect 5908 20392 5960 20398
rect 5906 20360 5908 20369
rect 6828 20392 6880 20398
rect 5960 20360 5962 20369
rect 6828 20334 6880 20340
rect 5906 20295 5962 20304
rect 5816 19984 5868 19990
rect 5816 19926 5868 19932
rect 5540 19916 5592 19922
rect 5540 19858 5592 19864
rect 5632 19916 5684 19922
rect 5632 19858 5684 19864
rect 5356 19848 5408 19854
rect 5356 19790 5408 19796
rect 5552 19310 5580 19858
rect 5540 19304 5592 19310
rect 5540 19246 5592 19252
rect 5356 18692 5408 18698
rect 5356 18634 5408 18640
rect 5368 17746 5396 18634
rect 5552 18306 5580 19246
rect 5644 18970 5672 19858
rect 5828 19310 5856 19926
rect 5816 19304 5868 19310
rect 5816 19246 5868 19252
rect 5632 18964 5684 18970
rect 5632 18906 5684 18912
rect 5460 18290 5580 18306
rect 5448 18284 5580 18290
rect 5500 18278 5580 18284
rect 5448 18226 5500 18232
rect 5644 18222 5672 18906
rect 5724 18828 5776 18834
rect 5724 18770 5776 18776
rect 5736 18630 5764 18770
rect 5724 18624 5776 18630
rect 5724 18566 5776 18572
rect 5632 18216 5684 18222
rect 5632 18158 5684 18164
rect 5828 18154 5856 19246
rect 5920 18766 5948 20295
rect 6840 19854 6868 20334
rect 6932 19922 6960 20454
rect 6920 19916 6972 19922
rect 6920 19858 6972 19864
rect 6828 19848 6880 19854
rect 6828 19790 6880 19796
rect 6000 19236 6052 19242
rect 6000 19178 6052 19184
rect 6012 18834 6040 19178
rect 6000 18828 6052 18834
rect 6000 18770 6052 18776
rect 5908 18760 5960 18766
rect 5908 18702 5960 18708
rect 5816 18148 5868 18154
rect 5816 18090 5868 18096
rect 5448 17876 5500 17882
rect 5448 17818 5500 17824
rect 5356 17740 5408 17746
rect 5356 17682 5408 17688
rect 5368 16794 5396 17682
rect 5460 17134 5488 17818
rect 6012 17762 6040 18770
rect 6092 18624 6144 18630
rect 6092 18566 6144 18572
rect 6104 17785 6132 18566
rect 6840 18358 6868 19790
rect 7300 19446 7328 22630
rect 7392 22234 7420 24686
rect 7484 24138 7512 25706
rect 7656 25696 7708 25702
rect 7656 25638 7708 25644
rect 7564 25356 7616 25362
rect 7564 25298 7616 25304
rect 7576 24750 7604 25298
rect 7668 24750 7696 25638
rect 7760 25294 7788 26522
rect 7852 26246 7880 26862
rect 7840 26240 7892 26246
rect 7840 26182 7892 26188
rect 7748 25288 7800 25294
rect 7748 25230 7800 25236
rect 7564 24744 7616 24750
rect 7564 24686 7616 24692
rect 7656 24744 7708 24750
rect 7656 24686 7708 24692
rect 7760 24274 7788 25230
rect 7748 24268 7800 24274
rect 7748 24210 7800 24216
rect 7472 24132 7524 24138
rect 7472 24074 7524 24080
rect 7380 22228 7432 22234
rect 7380 22170 7432 22176
rect 7760 22098 7788 24210
rect 7840 23180 7892 23186
rect 7840 23122 7892 23128
rect 7852 22642 7880 23122
rect 7840 22636 7892 22642
rect 7840 22578 7892 22584
rect 7748 22092 7800 22098
rect 7748 22034 7800 22040
rect 7840 21004 7892 21010
rect 7840 20946 7892 20952
rect 7472 20800 7524 20806
rect 7472 20742 7524 20748
rect 7484 19854 7512 20742
rect 7472 19848 7524 19854
rect 7472 19790 7524 19796
rect 7288 19440 7340 19446
rect 7288 19382 7340 19388
rect 7104 19304 7156 19310
rect 7104 19246 7156 19252
rect 6828 18352 6880 18358
rect 6828 18294 6880 18300
rect 6920 18148 6972 18154
rect 6920 18090 6972 18096
rect 5920 17746 6040 17762
rect 5908 17740 6040 17746
rect 5960 17734 6040 17740
rect 6090 17776 6146 17785
rect 6090 17711 6092 17720
rect 5908 17682 5960 17688
rect 6144 17711 6146 17720
rect 6092 17682 6144 17688
rect 6104 17651 6132 17682
rect 6932 17338 6960 18090
rect 7116 17785 7144 19246
rect 7196 18216 7248 18222
rect 7196 18158 7248 18164
rect 7102 17776 7158 17785
rect 7102 17711 7104 17720
rect 7156 17711 7158 17720
rect 7104 17682 7156 17688
rect 6920 17332 6972 17338
rect 6920 17274 6972 17280
rect 6184 17196 6236 17202
rect 6184 17138 6236 17144
rect 5448 17128 5500 17134
rect 5448 17070 5500 17076
rect 5356 16788 5408 16794
rect 5356 16730 5408 16736
rect 6196 16658 6224 17138
rect 6276 17128 6328 17134
rect 6276 17070 6328 17076
rect 6184 16652 6236 16658
rect 6184 16594 6236 16600
rect 6288 16250 6316 17070
rect 6552 17060 6604 17066
rect 6552 17002 6604 17008
rect 6564 16658 6592 17002
rect 7208 16658 7236 18158
rect 6552 16652 6604 16658
rect 6552 16594 6604 16600
rect 7196 16652 7248 16658
rect 7196 16594 7248 16600
rect 6276 16244 6328 16250
rect 6276 16186 6328 16192
rect 6564 16114 6592 16594
rect 6552 16108 6604 16114
rect 6552 16050 6604 16056
rect 5172 16040 5224 16046
rect 5172 15982 5224 15988
rect 7012 16040 7064 16046
rect 7012 15982 7064 15988
rect 6920 15496 6972 15502
rect 6920 15438 6972 15444
rect 6932 15094 6960 15438
rect 7024 15162 7052 15982
rect 7012 15156 7064 15162
rect 7012 15098 7064 15104
rect 6920 15088 6972 15094
rect 6920 15030 6972 15036
rect 7104 14816 7156 14822
rect 7104 14758 7156 14764
rect 5446 14512 5502 14521
rect 5446 14447 5448 14456
rect 5500 14447 5502 14456
rect 5448 14418 5500 14424
rect 5080 14408 5132 14414
rect 5080 14350 5132 14356
rect 6184 14408 6236 14414
rect 6184 14350 6236 14356
rect 6196 14006 6224 14350
rect 6184 14000 6236 14006
rect 6184 13942 6236 13948
rect 4620 13932 4672 13938
rect 4620 13874 4672 13880
rect 5264 13932 5316 13938
rect 5264 13874 5316 13880
rect 4160 13864 4212 13870
rect 4080 13824 4160 13852
rect 3976 13806 4028 13812
rect 4160 13806 4212 13812
rect 5080 13456 5132 13462
rect 5080 13398 5132 13404
rect 4804 13388 4856 13394
rect 4804 13330 4856 13336
rect 4220 13084 4516 13104
rect 4276 13082 4300 13084
rect 4356 13082 4380 13084
rect 4436 13082 4460 13084
rect 4298 13030 4300 13082
rect 4362 13030 4374 13082
rect 4436 13030 4438 13082
rect 4276 13028 4300 13030
rect 4356 13028 4380 13030
rect 4436 13028 4460 13030
rect 4220 13008 4516 13028
rect 4220 11996 4516 12016
rect 4276 11994 4300 11996
rect 4356 11994 4380 11996
rect 4436 11994 4460 11996
rect 4298 11942 4300 11994
rect 4362 11942 4374 11994
rect 4436 11942 4438 11994
rect 4276 11940 4300 11942
rect 4356 11940 4380 11942
rect 4436 11940 4460 11942
rect 4220 11920 4516 11940
rect 3884 11212 3936 11218
rect 3884 11154 3936 11160
rect 4620 11008 4672 11014
rect 4620 10950 4672 10956
rect 4220 10908 4516 10928
rect 4276 10906 4300 10908
rect 4356 10906 4380 10908
rect 4436 10906 4460 10908
rect 4298 10854 4300 10906
rect 4362 10854 4374 10906
rect 4436 10854 4438 10906
rect 4276 10852 4300 10854
rect 4356 10852 4380 10854
rect 4436 10852 4460 10854
rect 4220 10832 4516 10852
rect 3884 10804 3936 10810
rect 3884 10746 3936 10752
rect 3608 10532 3660 10538
rect 3608 10474 3660 10480
rect 3516 10464 3568 10470
rect 3516 10406 3568 10412
rect 3896 9518 3924 10746
rect 4632 10674 4660 10950
rect 4620 10668 4672 10674
rect 4620 10610 4672 10616
rect 4344 10600 4396 10606
rect 4344 10542 4396 10548
rect 4356 10266 4384 10542
rect 4344 10260 4396 10266
rect 4344 10202 4396 10208
rect 4220 9820 4516 9840
rect 4276 9818 4300 9820
rect 4356 9818 4380 9820
rect 4436 9818 4460 9820
rect 4298 9766 4300 9818
rect 4362 9766 4374 9818
rect 4436 9766 4438 9818
rect 4276 9764 4300 9766
rect 4356 9764 4380 9766
rect 4436 9764 4460 9766
rect 4220 9744 4516 9764
rect 4632 9654 4660 10610
rect 4712 10056 4764 10062
rect 4712 9998 4764 10004
rect 4068 9648 4120 9654
rect 4068 9590 4120 9596
rect 4620 9648 4672 9654
rect 4620 9590 4672 9596
rect 3884 9512 3936 9518
rect 3884 9454 3936 9460
rect 2964 9172 3016 9178
rect 2964 9114 3016 9120
rect 4080 9042 4108 9590
rect 4724 9586 4752 9998
rect 4712 9580 4764 9586
rect 4712 9522 4764 9528
rect 4436 9444 4488 9450
rect 4436 9386 4488 9392
rect 4160 9376 4212 9382
rect 4160 9318 4212 9324
rect 4068 9036 4120 9042
rect 4068 8978 4120 8984
rect 4172 8922 4200 9318
rect 4448 9042 4476 9386
rect 4816 9058 4844 13330
rect 4988 10124 5040 10130
rect 4988 10066 5040 10072
rect 4896 9376 4948 9382
rect 4896 9318 4948 9324
rect 4436 9036 4488 9042
rect 4724 9030 4844 9058
rect 4908 9042 4936 9318
rect 4896 9036 4948 9042
rect 4488 8996 4568 9024
rect 4436 8978 4488 8984
rect 4080 8894 4200 8922
rect 4540 8922 4568 8996
rect 4540 8894 4660 8922
rect 3700 8832 3752 8838
rect 3700 8774 3752 8780
rect 3516 7812 3568 7818
rect 3516 7754 3568 7760
rect 2964 7744 3016 7750
rect 2964 7686 3016 7692
rect 2872 6792 2924 6798
rect 2872 6734 2924 6740
rect 2504 6656 2556 6662
rect 2504 6598 2556 6604
rect 2320 5160 2372 5166
rect 2320 5102 2372 5108
rect 2884 4826 2912 6734
rect 2976 6633 3004 7686
rect 3528 7410 3556 7754
rect 3516 7404 3568 7410
rect 3516 7346 3568 7352
rect 2962 6624 3018 6633
rect 2962 6559 3018 6568
rect 2872 4820 2924 4826
rect 2872 4762 2924 4768
rect 3712 4622 3740 8774
rect 4080 8634 4108 8894
rect 4220 8732 4516 8752
rect 4276 8730 4300 8732
rect 4356 8730 4380 8732
rect 4436 8730 4460 8732
rect 4298 8678 4300 8730
rect 4362 8678 4374 8730
rect 4436 8678 4438 8730
rect 4276 8676 4300 8678
rect 4356 8676 4380 8678
rect 4436 8676 4460 8678
rect 4220 8656 4516 8676
rect 4068 8628 4120 8634
rect 4068 8570 4120 8576
rect 4080 8514 4108 8570
rect 4080 8486 4200 8514
rect 4172 7954 4200 8486
rect 4632 8022 4660 8894
rect 4620 8016 4672 8022
rect 4620 7958 4672 7964
rect 4160 7948 4212 7954
rect 4160 7890 4212 7896
rect 4220 7644 4516 7664
rect 4276 7642 4300 7644
rect 4356 7642 4380 7644
rect 4436 7642 4460 7644
rect 4298 7590 4300 7642
rect 4362 7590 4374 7642
rect 4436 7590 4438 7642
rect 4276 7588 4300 7590
rect 4356 7588 4380 7590
rect 4436 7588 4460 7590
rect 4220 7568 4516 7588
rect 4632 7478 4660 7958
rect 4620 7472 4672 7478
rect 4620 7414 4672 7420
rect 4632 6866 4660 7414
rect 4724 6916 4752 9030
rect 4896 8978 4948 8984
rect 4804 8968 4856 8974
rect 4804 8910 4856 8916
rect 4816 8498 4844 8910
rect 4804 8492 4856 8498
rect 4804 8434 4856 8440
rect 4804 7948 4856 7954
rect 4804 7890 4856 7896
rect 4816 7426 4844 7890
rect 4908 7546 4936 8978
rect 5000 8430 5028 10066
rect 4988 8424 5040 8430
rect 4988 8366 5040 8372
rect 4988 8288 5040 8294
rect 4988 8230 5040 8236
rect 5000 7750 5028 8230
rect 4988 7744 5040 7750
rect 4988 7686 5040 7692
rect 4896 7540 4948 7546
rect 4896 7482 4948 7488
rect 4816 7398 4936 7426
rect 5000 7410 5028 7686
rect 4908 6916 4936 7398
rect 4988 7404 5040 7410
rect 4988 7346 5040 7352
rect 4988 6928 5040 6934
rect 4724 6888 4844 6916
rect 4908 6888 4988 6916
rect 4620 6860 4672 6866
rect 4672 6820 4752 6848
rect 4620 6802 4672 6808
rect 4620 6656 4672 6662
rect 4620 6598 4672 6604
rect 4220 6556 4516 6576
rect 4276 6554 4300 6556
rect 4356 6554 4380 6556
rect 4436 6554 4460 6556
rect 4298 6502 4300 6554
rect 4362 6502 4374 6554
rect 4436 6502 4438 6554
rect 4276 6500 4300 6502
rect 4356 6500 4380 6502
rect 4436 6500 4460 6502
rect 4220 6480 4516 6500
rect 4344 6316 4396 6322
rect 4344 6258 4396 6264
rect 4356 5778 4384 6258
rect 4632 6186 4660 6598
rect 4724 6390 4752 6820
rect 4712 6384 4764 6390
rect 4712 6326 4764 6332
rect 4620 6180 4672 6186
rect 4620 6122 4672 6128
rect 4344 5772 4396 5778
rect 4344 5714 4396 5720
rect 4068 5704 4120 5710
rect 4068 5646 4120 5652
rect 4080 5234 4108 5646
rect 4220 5468 4516 5488
rect 4276 5466 4300 5468
rect 4356 5466 4380 5468
rect 4436 5466 4460 5468
rect 4298 5414 4300 5466
rect 4362 5414 4374 5466
rect 4436 5414 4438 5466
rect 4276 5412 4300 5414
rect 4356 5412 4380 5414
rect 4436 5412 4460 5414
rect 4220 5392 4516 5412
rect 4068 5228 4120 5234
rect 4068 5170 4120 5176
rect 4528 5160 4580 5166
rect 4632 5148 4660 6122
rect 4580 5120 4660 5148
rect 4528 5102 4580 5108
rect 4068 5092 4120 5098
rect 4068 5034 4120 5040
rect 3700 4616 3752 4622
rect 3700 4558 3752 4564
rect 3712 4146 3740 4558
rect 4080 4146 4108 5034
rect 4816 4690 4844 6888
rect 4988 6870 5040 6876
rect 4896 6724 4948 6730
rect 4896 6666 4948 6672
rect 4908 5234 4936 6666
rect 5000 6254 5028 6870
rect 4988 6248 5040 6254
rect 4988 6190 5040 6196
rect 5092 6066 5120 13398
rect 5172 13320 5224 13326
rect 5172 13262 5224 13268
rect 5184 12238 5212 13262
rect 5276 12850 5304 13874
rect 5356 13864 5408 13870
rect 5816 13864 5868 13870
rect 5356 13806 5408 13812
rect 5814 13832 5816 13841
rect 5868 13832 5870 13841
rect 5368 12986 5396 13806
rect 5814 13767 5870 13776
rect 7116 13394 7144 14758
rect 7104 13388 7156 13394
rect 7104 13330 7156 13336
rect 7196 13388 7248 13394
rect 7196 13330 7248 13336
rect 6828 13184 6880 13190
rect 6828 13126 6880 13132
rect 5356 12980 5408 12986
rect 5356 12922 5408 12928
rect 5264 12844 5316 12850
rect 5264 12786 5316 12792
rect 6840 12782 6868 13126
rect 5724 12776 5776 12782
rect 5724 12718 5776 12724
rect 6828 12776 6880 12782
rect 6828 12718 6880 12724
rect 5172 12232 5224 12238
rect 5172 12174 5224 12180
rect 5448 12232 5500 12238
rect 5448 12174 5500 12180
rect 5184 10130 5212 12174
rect 5356 11212 5408 11218
rect 5356 11154 5408 11160
rect 5368 10198 5396 11154
rect 5460 11150 5488 12174
rect 5736 11898 5764 12718
rect 6184 12300 6236 12306
rect 6184 12242 6236 12248
rect 6196 11898 6224 12242
rect 6920 12096 6972 12102
rect 6920 12038 6972 12044
rect 5724 11892 5776 11898
rect 5724 11834 5776 11840
rect 6184 11892 6236 11898
rect 6184 11834 6236 11840
rect 6196 11286 6224 11834
rect 6932 11694 6960 12038
rect 7208 11898 7236 13330
rect 7196 11892 7248 11898
rect 7196 11834 7248 11840
rect 6920 11688 6972 11694
rect 6920 11630 6972 11636
rect 6184 11280 6236 11286
rect 6184 11222 6236 11228
rect 5448 11144 5500 11150
rect 5448 11086 5500 11092
rect 6184 10600 6236 10606
rect 6184 10542 6236 10548
rect 5356 10192 5408 10198
rect 5276 10152 5356 10180
rect 5172 10124 5224 10130
rect 5172 10066 5224 10072
rect 5172 9444 5224 9450
rect 5172 9386 5224 9392
rect 5184 9042 5212 9386
rect 5172 9036 5224 9042
rect 5172 8978 5224 8984
rect 5172 8424 5224 8430
rect 5172 8366 5224 8372
rect 5184 7342 5212 8366
rect 5276 7342 5304 10152
rect 5356 10134 5408 10140
rect 6196 10130 6224 10542
rect 6932 10130 6960 11630
rect 7104 11280 7156 11286
rect 7104 11222 7156 11228
rect 7012 11212 7064 11218
rect 7012 11154 7064 11160
rect 6184 10124 6236 10130
rect 6184 10066 6236 10072
rect 6920 10124 6972 10130
rect 6920 10066 6972 10072
rect 5448 9920 5500 9926
rect 5448 9862 5500 9868
rect 5460 9042 5488 9862
rect 6092 9444 6144 9450
rect 6092 9386 6144 9392
rect 6460 9444 6512 9450
rect 6460 9386 6512 9392
rect 6104 9042 6132 9386
rect 6184 9376 6236 9382
rect 6184 9318 6236 9324
rect 5448 9036 5500 9042
rect 5448 8978 5500 8984
rect 6092 9036 6144 9042
rect 6092 8978 6144 8984
rect 5356 7948 5408 7954
rect 5460 7936 5488 8978
rect 5908 8356 5960 8362
rect 5908 8298 5960 8304
rect 5920 7954 5948 8298
rect 6104 7954 6132 8978
rect 6196 8634 6224 9318
rect 6184 8628 6236 8634
rect 6184 8570 6236 8576
rect 6472 8566 6500 9386
rect 6460 8560 6512 8566
rect 6460 8502 6512 8508
rect 6472 8430 6500 8502
rect 6460 8424 6512 8430
rect 6460 8366 6512 8372
rect 6472 7954 6500 8366
rect 5408 7908 5488 7936
rect 5908 7948 5960 7954
rect 5356 7890 5408 7896
rect 5908 7890 5960 7896
rect 6092 7948 6144 7954
rect 6092 7890 6144 7896
rect 6460 7948 6512 7954
rect 6460 7890 6512 7896
rect 6104 7546 6132 7890
rect 6092 7540 6144 7546
rect 6092 7482 6144 7488
rect 6552 7540 6604 7546
rect 6552 7482 6604 7488
rect 5172 7336 5224 7342
rect 5172 7278 5224 7284
rect 5264 7336 5316 7342
rect 5264 7278 5316 7284
rect 6564 6866 6592 7482
rect 6276 6860 6328 6866
rect 6276 6802 6328 6808
rect 6552 6860 6604 6866
rect 6552 6802 6604 6808
rect 6184 6792 6236 6798
rect 6184 6734 6236 6740
rect 5540 6248 5592 6254
rect 5540 6190 5592 6196
rect 6092 6248 6144 6254
rect 6092 6190 6144 6196
rect 5000 6038 5120 6066
rect 4896 5228 4948 5234
rect 4896 5170 4948 5176
rect 4804 4684 4856 4690
rect 4804 4626 4856 4632
rect 4220 4380 4516 4400
rect 4276 4378 4300 4380
rect 4356 4378 4380 4380
rect 4436 4378 4460 4380
rect 4298 4326 4300 4378
rect 4362 4326 4374 4378
rect 4436 4326 4438 4378
rect 4276 4324 4300 4326
rect 4356 4324 4380 4326
rect 4436 4324 4460 4326
rect 4220 4304 4516 4324
rect 3700 4140 3752 4146
rect 3700 4082 3752 4088
rect 4068 4140 4120 4146
rect 4068 4082 4120 4088
rect 1952 2984 2004 2990
rect 1952 2926 2004 2932
rect 2596 2848 2648 2854
rect 2596 2790 2648 2796
rect 572 1828 624 1834
rect 572 1770 624 1776
rect 584 800 612 1770
rect 2608 800 2636 2790
rect 3712 2514 3740 4082
rect 4220 3292 4516 3312
rect 4276 3290 4300 3292
rect 4356 3290 4380 3292
rect 4436 3290 4460 3292
rect 4298 3238 4300 3290
rect 4362 3238 4374 3290
rect 4436 3238 4438 3290
rect 4276 3236 4300 3238
rect 4356 3236 4380 3238
rect 4436 3236 4460 3238
rect 4220 3216 4516 3236
rect 5000 2514 5028 6038
rect 5552 5914 5580 6190
rect 5540 5908 5592 5914
rect 5540 5850 5592 5856
rect 6104 5370 6132 6190
rect 6196 6186 6224 6734
rect 6288 6390 6316 6802
rect 6276 6384 6328 6390
rect 6276 6326 6328 6332
rect 6564 6322 6592 6802
rect 6828 6792 6880 6798
rect 6828 6734 6880 6740
rect 6552 6316 6604 6322
rect 6552 6258 6604 6264
rect 6184 6180 6236 6186
rect 6184 6122 6236 6128
rect 6552 5704 6604 5710
rect 6552 5646 6604 5652
rect 6092 5364 6144 5370
rect 6092 5306 6144 5312
rect 5172 4820 5224 4826
rect 5172 4762 5224 4768
rect 5184 3534 5212 4762
rect 6368 4684 6420 4690
rect 6368 4626 6420 4632
rect 5816 4276 5868 4282
rect 5816 4218 5868 4224
rect 5264 3936 5316 3942
rect 5264 3878 5316 3884
rect 5276 3602 5304 3878
rect 5264 3596 5316 3602
rect 5264 3538 5316 3544
rect 5172 3528 5224 3534
rect 5172 3470 5224 3476
rect 5724 3528 5776 3534
rect 5724 3470 5776 3476
rect 3700 2508 3752 2514
rect 3700 2450 3752 2456
rect 4988 2508 5040 2514
rect 4988 2450 5040 2456
rect 5736 2446 5764 3470
rect 5828 2990 5856 4218
rect 6380 4146 6408 4626
rect 6368 4140 6420 4146
rect 6368 4082 6420 4088
rect 6000 4072 6052 4078
rect 6000 4014 6052 4020
rect 6012 3670 6040 4014
rect 6000 3664 6052 3670
rect 6000 3606 6052 3612
rect 6380 3602 6408 4082
rect 6368 3596 6420 3602
rect 6368 3538 6420 3544
rect 6092 3460 6144 3466
rect 6092 3402 6144 3408
rect 6104 2990 6132 3402
rect 6564 3398 6592 5646
rect 6840 5166 6868 6734
rect 7024 6730 7052 11154
rect 7116 10810 7144 11222
rect 7104 10804 7156 10810
rect 7104 10746 7156 10752
rect 7300 9602 7328 19382
rect 7852 19378 7880 20946
rect 7840 19372 7892 19378
rect 7840 19314 7892 19320
rect 7748 19304 7800 19310
rect 7668 19252 7748 19258
rect 7668 19246 7800 19252
rect 7668 19230 7788 19246
rect 7564 19168 7616 19174
rect 7668 19122 7696 19230
rect 7616 19116 7696 19122
rect 7564 19110 7696 19116
rect 7748 19168 7800 19174
rect 7748 19110 7800 19116
rect 7576 19094 7696 19110
rect 7668 17746 7696 19094
rect 7760 18834 7788 19110
rect 7748 18828 7800 18834
rect 7748 18770 7800 18776
rect 7840 18352 7892 18358
rect 7840 18294 7892 18300
rect 7656 17740 7708 17746
rect 7656 17682 7708 17688
rect 7852 17134 7880 18294
rect 7840 17128 7892 17134
rect 7840 17070 7892 17076
rect 7852 16114 7880 17070
rect 7840 16108 7892 16114
rect 7840 16050 7892 16056
rect 7944 14396 7972 38286
rect 8116 38208 8168 38214
rect 8116 38150 8168 38156
rect 8128 37874 8156 38150
rect 8116 37868 8168 37874
rect 8116 37810 8168 37816
rect 8208 37868 8260 37874
rect 8208 37810 8260 37816
rect 8220 37330 8248 37810
rect 9048 37398 9076 38354
rect 9784 38010 9812 40200
rect 10968 38412 11020 38418
rect 10968 38354 11020 38360
rect 11336 38412 11388 38418
rect 11336 38354 11388 38360
rect 11428 38412 11480 38418
rect 11428 38354 11480 38360
rect 10784 38208 10836 38214
rect 10784 38150 10836 38156
rect 9772 38004 9824 38010
rect 9772 37946 9824 37952
rect 9680 37800 9732 37806
rect 9680 37742 9732 37748
rect 9036 37392 9088 37398
rect 9036 37334 9088 37340
rect 9692 37330 9720 37742
rect 8208 37324 8260 37330
rect 8208 37266 8260 37272
rect 8668 37324 8720 37330
rect 8668 37266 8720 37272
rect 9680 37324 9732 37330
rect 9680 37266 9732 37272
rect 8484 37256 8536 37262
rect 8484 37198 8536 37204
rect 8496 36786 8524 37198
rect 8680 36922 8708 37266
rect 9220 37256 9272 37262
rect 9220 37198 9272 37204
rect 9864 37256 9916 37262
rect 9864 37198 9916 37204
rect 8668 36916 8720 36922
rect 8668 36858 8720 36864
rect 9232 36854 9260 37198
rect 9680 37120 9732 37126
rect 9680 37062 9732 37068
rect 9220 36848 9272 36854
rect 9220 36790 9272 36796
rect 8484 36780 8536 36786
rect 8484 36722 8536 36728
rect 8576 36712 8628 36718
rect 8576 36654 8628 36660
rect 8116 36644 8168 36650
rect 8116 36586 8168 36592
rect 8024 36576 8076 36582
rect 8024 36518 8076 36524
rect 8036 35154 8064 36518
rect 8024 35148 8076 35154
rect 8024 35090 8076 35096
rect 8128 34746 8156 36586
rect 8588 36242 8616 36654
rect 8576 36236 8628 36242
rect 8576 36178 8628 36184
rect 9036 36032 9088 36038
rect 9036 35974 9088 35980
rect 8300 35624 8352 35630
rect 8300 35566 8352 35572
rect 8208 35148 8260 35154
rect 8208 35090 8260 35096
rect 8220 35018 8248 35090
rect 8208 35012 8260 35018
rect 8208 34954 8260 34960
rect 8116 34740 8168 34746
rect 8116 34682 8168 34688
rect 8128 34134 8156 34682
rect 8312 34202 8340 35566
rect 8484 35012 8536 35018
rect 8484 34954 8536 34960
rect 8392 34468 8444 34474
rect 8392 34410 8444 34416
rect 8300 34196 8352 34202
rect 8300 34138 8352 34144
rect 8116 34128 8168 34134
rect 8116 34070 8168 34076
rect 8128 33454 8156 34070
rect 8208 34060 8260 34066
rect 8208 34002 8260 34008
rect 8220 33590 8248 34002
rect 8404 33930 8432 34410
rect 8496 34066 8524 34954
rect 8760 34672 8812 34678
rect 8760 34614 8812 34620
rect 8576 34128 8628 34134
rect 8576 34070 8628 34076
rect 8484 34060 8536 34066
rect 8484 34002 8536 34008
rect 8392 33924 8444 33930
rect 8392 33866 8444 33872
rect 8300 33856 8352 33862
rect 8300 33798 8352 33804
rect 8208 33584 8260 33590
rect 8208 33526 8260 33532
rect 8312 33454 8340 33798
rect 8116 33448 8168 33454
rect 8116 33390 8168 33396
rect 8300 33448 8352 33454
rect 8300 33390 8352 33396
rect 8128 32842 8156 33390
rect 8404 33114 8432 33866
rect 8588 33658 8616 34070
rect 8576 33652 8628 33658
rect 8576 33594 8628 33600
rect 8392 33108 8444 33114
rect 8392 33050 8444 33056
rect 8588 32978 8616 33594
rect 8772 33318 8800 34614
rect 8944 34536 8996 34542
rect 8944 34478 8996 34484
rect 8852 34400 8904 34406
rect 8852 34342 8904 34348
rect 8864 34066 8892 34342
rect 8852 34060 8904 34066
rect 8852 34002 8904 34008
rect 8956 33402 8984 34478
rect 9048 34134 9076 35974
rect 9036 34128 9088 34134
rect 9036 34070 9088 34076
rect 8864 33386 8984 33402
rect 8852 33380 8984 33386
rect 8904 33374 8984 33380
rect 8852 33322 8904 33328
rect 8760 33312 8812 33318
rect 8760 33254 8812 33260
rect 8576 32972 8628 32978
rect 8576 32914 8628 32920
rect 8116 32836 8168 32842
rect 8116 32778 8168 32784
rect 8772 32774 8800 33254
rect 8956 33046 8984 33374
rect 8944 33040 8996 33046
rect 8944 32982 8996 32988
rect 9128 32972 9180 32978
rect 9128 32914 9180 32920
rect 8208 32768 8260 32774
rect 8208 32710 8260 32716
rect 8760 32768 8812 32774
rect 8760 32710 8812 32716
rect 8220 31890 8248 32710
rect 8300 32360 8352 32366
rect 8300 32302 8352 32308
rect 8760 32360 8812 32366
rect 8760 32302 8812 32308
rect 8208 31884 8260 31890
rect 8208 31826 8260 31832
rect 8220 31346 8248 31826
rect 8208 31340 8260 31346
rect 8208 31282 8260 31288
rect 8312 30258 8340 32302
rect 8772 31958 8800 32302
rect 8760 31952 8812 31958
rect 8760 31894 8812 31900
rect 8772 31278 8800 31894
rect 8760 31272 8812 31278
rect 8760 31214 8812 31220
rect 8392 30796 8444 30802
rect 8392 30738 8444 30744
rect 8300 30252 8352 30258
rect 8300 30194 8352 30200
rect 8404 30190 8432 30738
rect 8944 30592 8996 30598
rect 8944 30534 8996 30540
rect 8484 30252 8536 30258
rect 8484 30194 8536 30200
rect 8392 30184 8444 30190
rect 8392 30126 8444 30132
rect 8300 30116 8352 30122
rect 8300 30058 8352 30064
rect 8116 29708 8168 29714
rect 8116 29650 8168 29656
rect 8128 29170 8156 29650
rect 8312 29170 8340 30058
rect 8404 29510 8432 30126
rect 8392 29504 8444 29510
rect 8392 29446 8444 29452
rect 8404 29238 8432 29446
rect 8496 29306 8524 30194
rect 8760 30048 8812 30054
rect 8760 29990 8812 29996
rect 8484 29300 8536 29306
rect 8484 29242 8536 29248
rect 8392 29232 8444 29238
rect 8392 29174 8444 29180
rect 8116 29164 8168 29170
rect 8116 29106 8168 29112
rect 8300 29164 8352 29170
rect 8300 29106 8352 29112
rect 8128 27334 8156 29106
rect 8208 28552 8260 28558
rect 8208 28494 8260 28500
rect 8220 27674 8248 28494
rect 8208 27668 8260 27674
rect 8208 27610 8260 27616
rect 8116 27328 8168 27334
rect 8116 27270 8168 27276
rect 8116 26852 8168 26858
rect 8116 26794 8168 26800
rect 8024 25696 8076 25702
rect 8024 25638 8076 25644
rect 8036 21486 8064 25638
rect 8128 25430 8156 26794
rect 8220 26450 8248 27610
rect 8668 27532 8720 27538
rect 8668 27474 8720 27480
rect 8392 27328 8444 27334
rect 8392 27270 8444 27276
rect 8208 26444 8260 26450
rect 8208 26386 8260 26392
rect 8220 25838 8248 26386
rect 8208 25832 8260 25838
rect 8208 25774 8260 25780
rect 8116 25424 8168 25430
rect 8116 25366 8168 25372
rect 8404 25226 8432 27270
rect 8680 27130 8708 27474
rect 8668 27124 8720 27130
rect 8668 27066 8720 27072
rect 8576 27056 8628 27062
rect 8576 26998 8628 27004
rect 8588 25770 8616 26998
rect 8772 26586 8800 29990
rect 8852 29096 8904 29102
rect 8852 29038 8904 29044
rect 8864 26790 8892 29038
rect 8956 27946 8984 30534
rect 9140 30054 9168 32914
rect 9232 30598 9260 36790
rect 9692 36786 9720 37062
rect 9680 36780 9732 36786
rect 9680 36722 9732 36728
rect 9404 36236 9456 36242
rect 9404 36178 9456 36184
rect 9416 35834 9444 36178
rect 9404 35828 9456 35834
rect 9404 35770 9456 35776
rect 9876 35698 9904 37198
rect 10796 36718 10824 38150
rect 10980 37806 11008 38354
rect 11060 38208 11112 38214
rect 11060 38150 11112 38156
rect 10968 37800 11020 37806
rect 10968 37742 11020 37748
rect 10048 36712 10100 36718
rect 10048 36654 10100 36660
rect 10784 36712 10836 36718
rect 10784 36654 10836 36660
rect 10060 36106 10088 36654
rect 10324 36236 10376 36242
rect 10324 36178 10376 36184
rect 10784 36236 10836 36242
rect 10784 36178 10836 36184
rect 10048 36100 10100 36106
rect 10048 36042 10100 36048
rect 9864 35692 9916 35698
rect 9864 35634 9916 35640
rect 9588 35012 9640 35018
rect 9588 34954 9640 34960
rect 9600 34610 9628 34954
rect 9772 34944 9824 34950
rect 9772 34886 9824 34892
rect 9588 34604 9640 34610
rect 9588 34546 9640 34552
rect 9588 34128 9640 34134
rect 9588 34070 9640 34076
rect 9600 33386 9628 34070
rect 9588 33380 9640 33386
rect 9588 33322 9640 33328
rect 9680 32904 9732 32910
rect 9680 32846 9732 32852
rect 9588 32768 9640 32774
rect 9588 32710 9640 32716
rect 9600 32298 9628 32710
rect 9496 32292 9548 32298
rect 9496 32234 9548 32240
rect 9588 32292 9640 32298
rect 9588 32234 9640 32240
rect 9508 31482 9536 32234
rect 9600 31890 9628 32234
rect 9692 31890 9720 32846
rect 9588 31884 9640 31890
rect 9588 31826 9640 31832
rect 9680 31884 9732 31890
rect 9680 31826 9732 31832
rect 9496 31476 9548 31482
rect 9496 31418 9548 31424
rect 9784 30682 9812 34886
rect 9876 34406 9904 35634
rect 10336 35154 10364 36178
rect 10796 35630 10824 36178
rect 10980 35766 11008 37742
rect 11072 37330 11100 38150
rect 11060 37324 11112 37330
rect 11060 37266 11112 37272
rect 11348 36786 11376 38354
rect 11440 37806 11468 38354
rect 11428 37800 11480 37806
rect 11428 37742 11480 37748
rect 11808 37346 11836 40200
rect 13728 38412 13780 38418
rect 13728 38354 13780 38360
rect 12716 38208 12768 38214
rect 12716 38150 12768 38156
rect 12440 37800 12492 37806
rect 12440 37742 12492 37748
rect 11808 37318 12204 37346
rect 11888 37188 11940 37194
rect 11888 37130 11940 37136
rect 11336 36780 11388 36786
rect 11336 36722 11388 36728
rect 11900 36718 11928 37130
rect 11888 36712 11940 36718
rect 11888 36654 11940 36660
rect 11796 36576 11848 36582
rect 11796 36518 11848 36524
rect 11808 36242 11836 36518
rect 11796 36236 11848 36242
rect 11796 36178 11848 36184
rect 11244 36168 11296 36174
rect 11244 36110 11296 36116
rect 10968 35760 11020 35766
rect 10968 35702 11020 35708
rect 11256 35698 11284 36110
rect 11244 35692 11296 35698
rect 11244 35634 11296 35640
rect 10784 35624 10836 35630
rect 10784 35566 10836 35572
rect 11612 35624 11664 35630
rect 11612 35566 11664 35572
rect 10324 35148 10376 35154
rect 10324 35090 10376 35096
rect 10232 34536 10284 34542
rect 10232 34478 10284 34484
rect 9864 34400 9916 34406
rect 9864 34342 9916 34348
rect 9876 33930 9904 34342
rect 10244 34134 10272 34478
rect 10232 34128 10284 34134
rect 10232 34070 10284 34076
rect 9864 33924 9916 33930
rect 9864 33866 9916 33872
rect 10048 33924 10100 33930
rect 10048 33866 10100 33872
rect 9864 32360 9916 32366
rect 9864 32302 9916 32308
rect 9876 31686 9904 32302
rect 10060 31822 10088 33866
rect 10336 33454 10364 35090
rect 10796 35086 10824 35566
rect 11624 35154 11652 35566
rect 11612 35148 11664 35154
rect 11612 35090 11664 35096
rect 10784 35080 10836 35086
rect 10784 35022 10836 35028
rect 11624 34746 11652 35090
rect 11612 34740 11664 34746
rect 11612 34682 11664 34688
rect 11060 34536 11112 34542
rect 11060 34478 11112 34484
rect 10508 34400 10560 34406
rect 10508 34342 10560 34348
rect 10520 33454 10548 34342
rect 11072 34202 11100 34478
rect 11520 34468 11572 34474
rect 11520 34410 11572 34416
rect 11060 34196 11112 34202
rect 11060 34138 11112 34144
rect 10968 34128 11020 34134
rect 10968 34070 11020 34076
rect 10600 33992 10652 33998
rect 10600 33934 10652 33940
rect 10612 33454 10640 33934
rect 10324 33448 10376 33454
rect 10324 33390 10376 33396
rect 10508 33448 10560 33454
rect 10508 33390 10560 33396
rect 10600 33448 10652 33454
rect 10600 33390 10652 33396
rect 10232 32904 10284 32910
rect 10232 32846 10284 32852
rect 10244 32434 10272 32846
rect 10232 32428 10284 32434
rect 10232 32370 10284 32376
rect 10612 32366 10640 33390
rect 10980 33386 11008 34070
rect 11072 33454 11100 34138
rect 11532 34066 11560 34410
rect 11520 34060 11572 34066
rect 11520 34002 11572 34008
rect 11244 33992 11296 33998
rect 11244 33934 11296 33940
rect 11256 33658 11284 33934
rect 11244 33652 11296 33658
rect 11244 33594 11296 33600
rect 11060 33448 11112 33454
rect 11060 33390 11112 33396
rect 10968 33380 11020 33386
rect 10968 33322 11020 33328
rect 10980 33114 11008 33322
rect 10968 33108 11020 33114
rect 10968 33050 11020 33056
rect 10980 32502 11008 33050
rect 11072 32910 11100 33390
rect 11336 32972 11388 32978
rect 11336 32914 11388 32920
rect 11428 32972 11480 32978
rect 11428 32914 11480 32920
rect 11060 32904 11112 32910
rect 11060 32846 11112 32852
rect 10968 32496 11020 32502
rect 10968 32438 11020 32444
rect 11072 32366 11100 32846
rect 11348 32842 11376 32914
rect 11336 32836 11388 32842
rect 11336 32778 11388 32784
rect 10600 32360 10652 32366
rect 10600 32302 10652 32308
rect 11060 32360 11112 32366
rect 11060 32302 11112 32308
rect 10612 32026 10640 32302
rect 11072 32026 11100 32302
rect 11440 32298 11468 32914
rect 11428 32292 11480 32298
rect 11428 32234 11480 32240
rect 10600 32020 10652 32026
rect 10600 31962 10652 31968
rect 11060 32020 11112 32026
rect 11060 31962 11112 31968
rect 10048 31816 10100 31822
rect 10048 31758 10100 31764
rect 11336 31816 11388 31822
rect 11336 31758 11388 31764
rect 9864 31680 9916 31686
rect 9864 31622 9916 31628
rect 9876 31414 9904 31622
rect 9864 31408 9916 31414
rect 9864 31350 9916 31356
rect 10876 31204 10928 31210
rect 10876 31146 10928 31152
rect 10888 30802 10916 31146
rect 10416 30796 10468 30802
rect 10416 30738 10468 30744
rect 10876 30796 10928 30802
rect 10876 30738 10928 30744
rect 9784 30654 9904 30682
rect 9876 30598 9904 30654
rect 9220 30592 9272 30598
rect 9220 30534 9272 30540
rect 9864 30592 9916 30598
rect 9864 30534 9916 30540
rect 10140 30592 10192 30598
rect 10140 30534 10192 30540
rect 9876 30394 9904 30534
rect 9864 30388 9916 30394
rect 9864 30330 9916 30336
rect 9588 30252 9640 30258
rect 9588 30194 9640 30200
rect 9312 30184 9364 30190
rect 9600 30161 9628 30194
rect 9312 30126 9364 30132
rect 9586 30152 9642 30161
rect 9128 30048 9180 30054
rect 9128 29990 9180 29996
rect 9220 30048 9272 30054
rect 9220 29990 9272 29996
rect 9140 28694 9168 29990
rect 9232 29102 9260 29990
rect 9324 29850 9352 30126
rect 9586 30087 9642 30096
rect 9876 29866 9904 30330
rect 9956 30320 10008 30326
rect 9956 30262 10008 30268
rect 9312 29844 9364 29850
rect 9312 29786 9364 29792
rect 9692 29838 9904 29866
rect 9588 29776 9640 29782
rect 9588 29718 9640 29724
rect 9220 29096 9272 29102
rect 9220 29038 9272 29044
rect 9600 28966 9628 29718
rect 9692 29578 9720 29838
rect 9772 29776 9824 29782
rect 9772 29718 9824 29724
rect 9680 29572 9732 29578
rect 9680 29514 9732 29520
rect 9784 29238 9812 29718
rect 9772 29232 9824 29238
rect 9772 29174 9824 29180
rect 9588 28960 9640 28966
rect 9588 28902 9640 28908
rect 9128 28688 9180 28694
rect 9128 28630 9180 28636
rect 9128 28552 9180 28558
rect 9128 28494 9180 28500
rect 9140 28014 9168 28494
rect 9680 28076 9732 28082
rect 9680 28018 9732 28024
rect 9128 28008 9180 28014
rect 9128 27950 9180 27956
rect 8944 27940 8996 27946
rect 8944 27882 8996 27888
rect 8852 26784 8904 26790
rect 8852 26726 8904 26732
rect 8760 26580 8812 26586
rect 8760 26522 8812 26528
rect 8668 26444 8720 26450
rect 8668 26386 8720 26392
rect 8680 25838 8708 26386
rect 8668 25832 8720 25838
rect 8668 25774 8720 25780
rect 8576 25764 8628 25770
rect 8576 25706 8628 25712
rect 8588 25362 8616 25706
rect 8576 25356 8628 25362
rect 8576 25298 8628 25304
rect 8484 25288 8536 25294
rect 8484 25230 8536 25236
rect 8392 25220 8444 25226
rect 8392 25162 8444 25168
rect 8208 24880 8260 24886
rect 8208 24822 8260 24828
rect 8116 24744 8168 24750
rect 8116 24686 8168 24692
rect 8128 24614 8156 24686
rect 8116 24608 8168 24614
rect 8116 24550 8168 24556
rect 8128 22098 8156 24550
rect 8220 24274 8248 24822
rect 8392 24744 8444 24750
rect 8392 24686 8444 24692
rect 8208 24268 8260 24274
rect 8208 24210 8260 24216
rect 8404 24070 8432 24686
rect 8496 24274 8524 25230
rect 8576 25220 8628 25226
rect 8576 25162 8628 25168
rect 8484 24268 8536 24274
rect 8484 24210 8536 24216
rect 8392 24064 8444 24070
rect 8392 24006 8444 24012
rect 8496 23882 8524 24210
rect 8208 23860 8260 23866
rect 8208 23802 8260 23808
rect 8312 23854 8524 23882
rect 8220 23594 8248 23802
rect 8208 23588 8260 23594
rect 8208 23530 8260 23536
rect 8208 22432 8260 22438
rect 8208 22374 8260 22380
rect 8116 22092 8168 22098
rect 8116 22034 8168 22040
rect 8024 21480 8076 21486
rect 8024 21422 8076 21428
rect 8036 21078 8064 21422
rect 8024 21072 8076 21078
rect 8024 21014 8076 21020
rect 8220 20806 8248 22374
rect 8312 22030 8340 23854
rect 8392 23656 8444 23662
rect 8392 23598 8444 23604
rect 8300 22024 8352 22030
rect 8300 21966 8352 21972
rect 8404 21622 8432 23598
rect 8484 23588 8536 23594
rect 8484 23530 8536 23536
rect 8496 22642 8524 23530
rect 8484 22636 8536 22642
rect 8484 22578 8536 22584
rect 8588 22234 8616 25162
rect 8760 24064 8812 24070
rect 8760 24006 8812 24012
rect 8576 22228 8628 22234
rect 8576 22170 8628 22176
rect 8772 22166 8800 24006
rect 8760 22160 8812 22166
rect 8760 22102 8812 22108
rect 8484 22024 8536 22030
rect 8484 21966 8536 21972
rect 8392 21616 8444 21622
rect 8392 21558 8444 21564
rect 8404 21486 8432 21558
rect 8392 21480 8444 21486
rect 8392 21422 8444 21428
rect 8392 21004 8444 21010
rect 8392 20946 8444 20952
rect 8208 20800 8260 20806
rect 8208 20742 8260 20748
rect 8116 20596 8168 20602
rect 8116 20538 8168 20544
rect 8024 20460 8076 20466
rect 8024 20402 8076 20408
rect 8036 20369 8064 20402
rect 8022 20360 8078 20369
rect 8022 20295 8078 20304
rect 8128 19718 8156 20538
rect 8404 20534 8432 20946
rect 8392 20528 8444 20534
rect 8392 20470 8444 20476
rect 8392 20256 8444 20262
rect 8392 20198 8444 20204
rect 8208 19848 8260 19854
rect 8208 19790 8260 19796
rect 8116 19712 8168 19718
rect 8116 19654 8168 19660
rect 8116 18148 8168 18154
rect 8116 18090 8168 18096
rect 8128 17542 8156 18090
rect 8116 17536 8168 17542
rect 8116 17478 8168 17484
rect 8128 16658 8156 17478
rect 8220 16794 8248 19790
rect 8300 19304 8352 19310
rect 8300 19246 8352 19252
rect 8312 18834 8340 19246
rect 8404 19174 8432 20198
rect 8392 19168 8444 19174
rect 8392 19110 8444 19116
rect 8300 18828 8352 18834
rect 8300 18770 8352 18776
rect 8392 18216 8444 18222
rect 8392 18158 8444 18164
rect 8300 18148 8352 18154
rect 8300 18090 8352 18096
rect 8312 17610 8340 18090
rect 8300 17604 8352 17610
rect 8300 17546 8352 17552
rect 8208 16788 8260 16794
rect 8208 16730 8260 16736
rect 8404 16658 8432 18158
rect 8116 16652 8168 16658
rect 8116 16594 8168 16600
rect 8392 16652 8444 16658
rect 8392 16594 8444 16600
rect 8496 15570 8524 21966
rect 8956 21554 8984 27882
rect 9312 27872 9364 27878
rect 9312 27814 9364 27820
rect 9128 27532 9180 27538
rect 9128 27474 9180 27480
rect 9036 26580 9088 26586
rect 9036 26522 9088 26528
rect 8944 21548 8996 21554
rect 8944 21490 8996 21496
rect 8944 20800 8996 20806
rect 8944 20742 8996 20748
rect 8956 19922 8984 20742
rect 8944 19916 8996 19922
rect 8944 19858 8996 19864
rect 9048 19854 9076 26522
rect 9140 26518 9168 27474
rect 9324 26994 9352 27814
rect 9692 27470 9720 28018
rect 9680 27464 9732 27470
rect 9680 27406 9732 27412
rect 9312 26988 9364 26994
rect 9312 26930 9364 26936
rect 9128 26512 9180 26518
rect 9128 26454 9180 26460
rect 9772 26308 9824 26314
rect 9772 26250 9824 26256
rect 9404 25832 9456 25838
rect 9404 25774 9456 25780
rect 9416 24206 9444 25774
rect 9784 24750 9812 26250
rect 9876 24818 9904 29838
rect 9968 29102 9996 30262
rect 10152 30190 10180 30534
rect 10428 30394 10456 30738
rect 11152 30728 11204 30734
rect 11152 30670 11204 30676
rect 10600 30592 10652 30598
rect 10600 30534 10652 30540
rect 10232 30388 10284 30394
rect 10232 30330 10284 30336
rect 10416 30388 10468 30394
rect 10416 30330 10468 30336
rect 10244 30190 10272 30330
rect 10612 30326 10640 30534
rect 10968 30388 11020 30394
rect 10968 30330 11020 30336
rect 10600 30320 10652 30326
rect 10600 30262 10652 30268
rect 10140 30184 10192 30190
rect 10140 30126 10192 30132
rect 10232 30184 10284 30190
rect 10232 30126 10284 30132
rect 9956 29096 10008 29102
rect 9956 29038 10008 29044
rect 10152 28626 10180 30126
rect 10784 29504 10836 29510
rect 10784 29446 10836 29452
rect 10876 29504 10928 29510
rect 10876 29446 10928 29452
rect 10796 29102 10824 29446
rect 10888 29238 10916 29446
rect 10876 29232 10928 29238
rect 10876 29174 10928 29180
rect 10600 29096 10652 29102
rect 10600 29038 10652 29044
rect 10784 29096 10836 29102
rect 10784 29038 10836 29044
rect 10416 29028 10468 29034
rect 10416 28970 10468 28976
rect 10140 28620 10192 28626
rect 10140 28562 10192 28568
rect 10428 27538 10456 28970
rect 10612 28626 10640 29038
rect 10600 28620 10652 28626
rect 10600 28562 10652 28568
rect 10876 28620 10928 28626
rect 10876 28562 10928 28568
rect 10416 27532 10468 27538
rect 10416 27474 10468 27480
rect 10888 27470 10916 28562
rect 10876 27464 10928 27470
rect 10876 27406 10928 27412
rect 10508 26920 10560 26926
rect 10508 26862 10560 26868
rect 9864 24812 9916 24818
rect 9864 24754 9916 24760
rect 9772 24744 9824 24750
rect 9772 24686 9824 24692
rect 9956 24744 10008 24750
rect 9956 24686 10008 24692
rect 9404 24200 9456 24206
rect 9404 24142 9456 24148
rect 9864 24200 9916 24206
rect 9864 24142 9916 24148
rect 9876 23662 9904 24142
rect 9968 24138 9996 24686
rect 10232 24676 10284 24682
rect 10232 24618 10284 24624
rect 10244 24206 10272 24618
rect 10520 24614 10548 26862
rect 10784 26784 10836 26790
rect 10784 26726 10836 26732
rect 10796 26382 10824 26726
rect 10784 26376 10836 26382
rect 10784 26318 10836 26324
rect 10508 24608 10560 24614
rect 10508 24550 10560 24556
rect 10520 24274 10548 24550
rect 10324 24268 10376 24274
rect 10324 24210 10376 24216
rect 10508 24268 10560 24274
rect 10508 24210 10560 24216
rect 10232 24200 10284 24206
rect 10232 24142 10284 24148
rect 9956 24132 10008 24138
rect 9956 24074 10008 24080
rect 10336 24070 10364 24210
rect 10324 24064 10376 24070
rect 10324 24006 10376 24012
rect 10336 23662 10364 24006
rect 10520 23730 10548 24210
rect 10508 23724 10560 23730
rect 10508 23666 10560 23672
rect 10796 23662 10824 26318
rect 10888 25838 10916 27406
rect 10980 25974 11008 30330
rect 11164 29646 11192 30670
rect 11348 30190 11376 31758
rect 11704 30592 11756 30598
rect 11704 30534 11756 30540
rect 11716 30394 11744 30534
rect 11704 30388 11756 30394
rect 11704 30330 11756 30336
rect 11336 30184 11388 30190
rect 11336 30126 11388 30132
rect 11152 29640 11204 29646
rect 11152 29582 11204 29588
rect 11164 28422 11192 29582
rect 11348 29238 11376 30126
rect 11336 29232 11388 29238
rect 11336 29174 11388 29180
rect 11704 28960 11756 28966
rect 11704 28902 11756 28908
rect 11336 28688 11388 28694
rect 11336 28630 11388 28636
rect 11244 28484 11296 28490
rect 11244 28426 11296 28432
rect 11152 28416 11204 28422
rect 11152 28358 11204 28364
rect 11164 28150 11192 28358
rect 11152 28144 11204 28150
rect 11152 28086 11204 28092
rect 11164 27538 11192 28086
rect 11152 27532 11204 27538
rect 11152 27474 11204 27480
rect 11060 26444 11112 26450
rect 11060 26386 11112 26392
rect 11072 25974 11100 26386
rect 10968 25968 11020 25974
rect 10968 25910 11020 25916
rect 11060 25968 11112 25974
rect 11060 25910 11112 25916
rect 10876 25832 10928 25838
rect 10876 25774 10928 25780
rect 10980 25702 11008 25910
rect 11164 25820 11192 27474
rect 11256 26450 11284 28426
rect 11348 28150 11376 28630
rect 11612 28484 11664 28490
rect 11612 28426 11664 28432
rect 11336 28144 11388 28150
rect 11336 28086 11388 28092
rect 11348 27130 11376 28086
rect 11624 28014 11652 28426
rect 11716 28422 11744 28902
rect 11704 28416 11756 28422
rect 11704 28358 11756 28364
rect 12176 28150 12204 37318
rect 12452 37262 12480 37742
rect 12440 37256 12492 37262
rect 12440 37198 12492 37204
rect 12728 36310 12756 38150
rect 13544 37800 13596 37806
rect 13544 37742 13596 37748
rect 13176 37120 13228 37126
rect 13176 37062 13228 37068
rect 13188 36650 13216 37062
rect 13176 36644 13228 36650
rect 13176 36586 13228 36592
rect 12900 36576 12952 36582
rect 12900 36518 12952 36524
rect 12912 36378 12940 36518
rect 12900 36372 12952 36378
rect 12900 36314 12952 36320
rect 12716 36304 12768 36310
rect 12716 36246 12768 36252
rect 12532 36236 12584 36242
rect 12532 36178 12584 36184
rect 12544 35698 12572 36178
rect 12532 35692 12584 35698
rect 12532 35634 12584 35640
rect 12440 35624 12492 35630
rect 12440 35566 12492 35572
rect 12452 35222 12480 35566
rect 12544 35290 12572 35634
rect 12912 35630 12940 36314
rect 12900 35624 12952 35630
rect 12900 35566 12952 35572
rect 13084 35488 13136 35494
rect 13084 35430 13136 35436
rect 12532 35284 12584 35290
rect 12532 35226 12584 35232
rect 12440 35216 12492 35222
rect 12440 35158 12492 35164
rect 13096 35154 13124 35430
rect 13084 35148 13136 35154
rect 13084 35090 13136 35096
rect 13176 35080 13228 35086
rect 13176 35022 13228 35028
rect 12624 34536 12676 34542
rect 12624 34478 12676 34484
rect 12636 34406 12664 34478
rect 12624 34400 12676 34406
rect 12624 34342 12676 34348
rect 12636 34134 12664 34342
rect 12624 34128 12676 34134
rect 12624 34070 12676 34076
rect 13188 33862 13216 35022
rect 13360 34060 13412 34066
rect 13360 34002 13412 34008
rect 13176 33856 13228 33862
rect 13176 33798 13228 33804
rect 13188 32434 13216 33798
rect 13372 33590 13400 34002
rect 13360 33584 13412 33590
rect 13360 33526 13412 33532
rect 13372 33046 13400 33526
rect 13452 33380 13504 33386
rect 13452 33322 13504 33328
rect 13360 33040 13412 33046
rect 13360 32982 13412 32988
rect 13464 32434 13492 33322
rect 13176 32428 13228 32434
rect 13176 32370 13228 32376
rect 13452 32428 13504 32434
rect 13452 32370 13504 32376
rect 12256 31884 12308 31890
rect 12256 31826 12308 31832
rect 12992 31884 13044 31890
rect 12992 31826 13044 31832
rect 12268 29578 12296 31826
rect 12900 31272 12952 31278
rect 12900 31214 12952 31220
rect 12440 30320 12492 30326
rect 12440 30262 12492 30268
rect 12256 29572 12308 29578
rect 12256 29514 12308 29520
rect 12164 28144 12216 28150
rect 12164 28086 12216 28092
rect 11612 28008 11664 28014
rect 11612 27950 11664 27956
rect 11612 27872 11664 27878
rect 11612 27814 11664 27820
rect 11624 27538 11652 27814
rect 11612 27532 11664 27538
rect 11612 27474 11664 27480
rect 11428 27464 11480 27470
rect 11428 27406 11480 27412
rect 11336 27124 11388 27130
rect 11336 27066 11388 27072
rect 11440 26858 11468 27406
rect 12268 27334 12296 29514
rect 12256 27328 12308 27334
rect 12256 27270 12308 27276
rect 11428 26852 11480 26858
rect 11428 26794 11480 26800
rect 11440 26450 11468 26794
rect 12268 26518 12296 27270
rect 12452 26926 12480 30262
rect 12532 30184 12584 30190
rect 12532 30126 12584 30132
rect 12544 29646 12572 30126
rect 12532 29640 12584 29646
rect 12532 29582 12584 29588
rect 12912 29578 12940 31214
rect 13004 30394 13032 31826
rect 13360 31136 13412 31142
rect 13360 31078 13412 31084
rect 12992 30388 13044 30394
rect 12992 30330 13044 30336
rect 13372 29714 13400 31078
rect 13360 29708 13412 29714
rect 13360 29650 13412 29656
rect 12900 29572 12952 29578
rect 12900 29514 12952 29520
rect 12716 29096 12768 29102
rect 12716 29038 12768 29044
rect 12624 28484 12676 28490
rect 12624 28426 12676 28432
rect 12636 27010 12664 28426
rect 12728 27130 12756 29038
rect 12716 27124 12768 27130
rect 12716 27066 12768 27072
rect 13556 27010 13584 37742
rect 13740 37330 13768 38354
rect 14016 38010 14044 40200
rect 14004 38004 14056 38010
rect 14004 37946 14056 37952
rect 15292 37868 15344 37874
rect 15292 37810 15344 37816
rect 14004 37664 14056 37670
rect 14004 37606 14056 37612
rect 14016 37398 14044 37606
rect 14004 37392 14056 37398
rect 14004 37334 14056 37340
rect 13728 37324 13780 37330
rect 13728 37266 13780 37272
rect 13740 37126 13768 37266
rect 13912 37256 13964 37262
rect 13912 37198 13964 37204
rect 13728 37120 13780 37126
rect 13728 37062 13780 37068
rect 13728 36712 13780 36718
rect 13728 36654 13780 36660
rect 13740 36242 13768 36654
rect 13924 36242 13952 37198
rect 14016 36718 14044 37334
rect 14096 37324 14148 37330
rect 14096 37266 14148 37272
rect 14372 37324 14424 37330
rect 14372 37266 14424 37272
rect 14004 36712 14056 36718
rect 14004 36654 14056 36660
rect 14108 36310 14136 37266
rect 14384 37194 14412 37266
rect 15304 37244 15332 37810
rect 15844 37800 15896 37806
rect 15844 37742 15896 37748
rect 15752 37324 15804 37330
rect 15752 37266 15804 37272
rect 15384 37256 15436 37262
rect 15304 37216 15384 37244
rect 14372 37188 14424 37194
rect 14424 37148 14504 37176
rect 14372 37130 14424 37136
rect 14384 37065 14412 37130
rect 14372 36916 14424 36922
rect 14372 36858 14424 36864
rect 14280 36712 14332 36718
rect 14280 36654 14332 36660
rect 14096 36304 14148 36310
rect 14096 36246 14148 36252
rect 14292 36242 14320 36654
rect 13728 36236 13780 36242
rect 13728 36178 13780 36184
rect 13912 36236 13964 36242
rect 13912 36178 13964 36184
rect 14280 36236 14332 36242
rect 14280 36178 14332 36184
rect 13820 36100 13872 36106
rect 13820 36042 13872 36048
rect 13832 33998 13860 36042
rect 13924 35766 13952 36178
rect 13912 35760 13964 35766
rect 13912 35702 13964 35708
rect 14292 34950 14320 36178
rect 14384 35630 14412 36858
rect 14476 36718 14504 37148
rect 15016 37120 15068 37126
rect 15016 37062 15068 37068
rect 15200 37120 15252 37126
rect 15200 37062 15252 37068
rect 15028 36718 15056 37062
rect 15212 36786 15240 37062
rect 15200 36780 15252 36786
rect 15200 36722 15252 36728
rect 14464 36712 14516 36718
rect 14464 36654 14516 36660
rect 15016 36712 15068 36718
rect 15016 36654 15068 36660
rect 14372 35624 14424 35630
rect 14372 35566 14424 35572
rect 14004 34944 14056 34950
rect 14004 34886 14056 34892
rect 14280 34944 14332 34950
rect 14280 34886 14332 34892
rect 13912 34604 13964 34610
rect 13912 34546 13964 34552
rect 13924 34066 13952 34546
rect 14016 34542 14044 34886
rect 14476 34542 14504 36654
rect 14924 35692 14976 35698
rect 14924 35634 14976 35640
rect 14832 35556 14884 35562
rect 14832 35498 14884 35504
rect 14844 35154 14872 35498
rect 14832 35148 14884 35154
rect 14832 35090 14884 35096
rect 14004 34536 14056 34542
rect 14004 34478 14056 34484
rect 14464 34536 14516 34542
rect 14464 34478 14516 34484
rect 13912 34060 13964 34066
rect 13912 34002 13964 34008
rect 13820 33992 13872 33998
rect 13820 33934 13872 33940
rect 13636 33448 13688 33454
rect 13636 33390 13688 33396
rect 13912 33448 13964 33454
rect 13912 33390 13964 33396
rect 14004 33448 14056 33454
rect 14004 33390 14056 33396
rect 13648 32026 13676 33390
rect 13636 32020 13688 32026
rect 13636 31962 13688 31968
rect 13924 31958 13952 33390
rect 13912 31952 13964 31958
rect 13912 31894 13964 31900
rect 14016 31890 14044 33390
rect 14464 32972 14516 32978
rect 14464 32914 14516 32920
rect 14476 32026 14504 32914
rect 14556 32428 14608 32434
rect 14556 32370 14608 32376
rect 14464 32020 14516 32026
rect 14464 31962 14516 31968
rect 13636 31884 13688 31890
rect 13636 31826 13688 31832
rect 14004 31884 14056 31890
rect 14004 31826 14056 31832
rect 13648 31278 13676 31826
rect 14016 31278 14044 31826
rect 13636 31272 13688 31278
rect 13636 31214 13688 31220
rect 14004 31272 14056 31278
rect 14004 31214 14056 31220
rect 14280 30796 14332 30802
rect 14280 30738 14332 30744
rect 14188 30728 14240 30734
rect 14188 30670 14240 30676
rect 13912 30184 13964 30190
rect 13912 30126 13964 30132
rect 13820 30048 13872 30054
rect 13820 29990 13872 29996
rect 13636 29844 13688 29850
rect 13636 29786 13688 29792
rect 13648 29238 13676 29786
rect 13832 29306 13860 29990
rect 13924 29782 13952 30126
rect 14004 29844 14056 29850
rect 14004 29786 14056 29792
rect 13912 29776 13964 29782
rect 13912 29718 13964 29724
rect 13924 29306 13952 29718
rect 14016 29510 14044 29786
rect 14096 29708 14148 29714
rect 14096 29650 14148 29656
rect 14004 29504 14056 29510
rect 14004 29446 14056 29452
rect 13820 29300 13872 29306
rect 13820 29242 13872 29248
rect 13912 29300 13964 29306
rect 13912 29242 13964 29248
rect 13636 29232 13688 29238
rect 13636 29174 13688 29180
rect 14108 29170 14136 29650
rect 14096 29164 14148 29170
rect 14096 29106 14148 29112
rect 14108 29034 14136 29106
rect 14200 29102 14228 30670
rect 14292 29714 14320 30738
rect 14464 30184 14516 30190
rect 14568 30172 14596 32370
rect 14832 32292 14884 32298
rect 14832 32234 14884 32240
rect 14648 31680 14700 31686
rect 14648 31622 14700 31628
rect 14660 31278 14688 31622
rect 14648 31272 14700 31278
rect 14648 31214 14700 31220
rect 14660 31142 14688 31214
rect 14648 31136 14700 31142
rect 14648 31078 14700 31084
rect 14516 30144 14596 30172
rect 14464 30126 14516 30132
rect 14280 29708 14332 29714
rect 14280 29650 14332 29656
rect 14476 29170 14504 30126
rect 14660 30122 14688 31078
rect 14844 30802 14872 32234
rect 14832 30796 14884 30802
rect 14832 30738 14884 30744
rect 14844 30258 14872 30738
rect 14832 30252 14884 30258
rect 14832 30194 14884 30200
rect 14648 30116 14700 30122
rect 14648 30058 14700 30064
rect 14464 29164 14516 29170
rect 14464 29106 14516 29112
rect 14660 29102 14688 30058
rect 14188 29096 14240 29102
rect 14188 29038 14240 29044
rect 14648 29096 14700 29102
rect 14648 29038 14700 29044
rect 14096 29028 14148 29034
rect 14096 28970 14148 28976
rect 14108 28626 14136 28970
rect 13636 28620 13688 28626
rect 13636 28562 13688 28568
rect 14096 28620 14148 28626
rect 14096 28562 14148 28568
rect 13648 28014 13676 28562
rect 14004 28552 14056 28558
rect 14004 28494 14056 28500
rect 14016 28014 14044 28494
rect 13636 28008 13688 28014
rect 13636 27950 13688 27956
rect 14004 28008 14056 28014
rect 14004 27950 14056 27956
rect 13648 27538 13676 27950
rect 14016 27606 14044 27950
rect 14556 27872 14608 27878
rect 14556 27814 14608 27820
rect 14004 27600 14056 27606
rect 14004 27542 14056 27548
rect 13636 27532 13688 27538
rect 13636 27474 13688 27480
rect 13912 27396 13964 27402
rect 13912 27338 13964 27344
rect 12636 26982 12940 27010
rect 13556 26982 13676 27010
rect 12440 26920 12492 26926
rect 12440 26862 12492 26868
rect 12256 26512 12308 26518
rect 12256 26454 12308 26460
rect 11244 26444 11296 26450
rect 11244 26386 11296 26392
rect 11428 26444 11480 26450
rect 11428 26386 11480 26392
rect 11520 26444 11572 26450
rect 11520 26386 11572 26392
rect 11428 26240 11480 26246
rect 11428 26182 11480 26188
rect 11244 25968 11296 25974
rect 11244 25910 11296 25916
rect 11072 25792 11192 25820
rect 10968 25696 11020 25702
rect 10968 25638 11020 25644
rect 11072 25362 11100 25792
rect 11152 25424 11204 25430
rect 11152 25366 11204 25372
rect 11060 25356 11112 25362
rect 11060 25298 11112 25304
rect 11060 24744 11112 24750
rect 11060 24686 11112 24692
rect 10968 24132 11020 24138
rect 10968 24074 11020 24080
rect 9864 23656 9916 23662
rect 9864 23598 9916 23604
rect 10324 23656 10376 23662
rect 10324 23598 10376 23604
rect 10784 23656 10836 23662
rect 10784 23598 10836 23604
rect 9772 23588 9824 23594
rect 9772 23530 9824 23536
rect 9784 22438 9812 23530
rect 10324 23520 10376 23526
rect 10324 23462 10376 23468
rect 10336 23186 10364 23462
rect 10796 23322 10824 23598
rect 10784 23316 10836 23322
rect 10784 23258 10836 23264
rect 10140 23180 10192 23186
rect 10140 23122 10192 23128
rect 10324 23180 10376 23186
rect 10324 23122 10376 23128
rect 10876 23180 10928 23186
rect 10876 23122 10928 23128
rect 10152 22642 10180 23122
rect 10140 22636 10192 22642
rect 10140 22578 10192 22584
rect 9772 22432 9824 22438
rect 9772 22374 9824 22380
rect 9680 22160 9732 22166
rect 9680 22102 9732 22108
rect 9692 21622 9720 22102
rect 9680 21616 9732 21622
rect 9680 21558 9732 21564
rect 9220 21412 9272 21418
rect 9220 21354 9272 21360
rect 9128 19916 9180 19922
rect 9128 19858 9180 19864
rect 9036 19848 9088 19854
rect 9036 19790 9088 19796
rect 9140 19310 9168 19858
rect 9128 19304 9180 19310
rect 9128 19246 9180 19252
rect 8576 18760 8628 18766
rect 8576 18702 8628 18708
rect 8588 17746 8616 18702
rect 9232 17898 9260 21354
rect 9784 21010 9812 22374
rect 9956 22024 10008 22030
rect 9956 21966 10008 21972
rect 10232 22024 10284 22030
rect 10232 21966 10284 21972
rect 9864 21684 9916 21690
rect 9864 21626 9916 21632
rect 9876 21486 9904 21626
rect 9864 21480 9916 21486
rect 9864 21422 9916 21428
rect 9968 21010 9996 21966
rect 10244 21554 10272 21966
rect 10336 21962 10364 23122
rect 10888 22982 10916 23122
rect 10876 22976 10928 22982
rect 10876 22918 10928 22924
rect 10888 22098 10916 22918
rect 10980 22166 11008 24074
rect 11072 23118 11100 24686
rect 11164 24274 11192 25366
rect 11152 24268 11204 24274
rect 11152 24210 11204 24216
rect 11256 23798 11284 25910
rect 11440 25770 11468 26182
rect 11428 25764 11480 25770
rect 11428 25706 11480 25712
rect 11532 25430 11560 26386
rect 11980 26308 12032 26314
rect 11980 26250 12032 26256
rect 11992 25906 12020 26250
rect 11980 25900 12032 25906
rect 11980 25842 12032 25848
rect 11992 25430 12020 25842
rect 12532 25832 12584 25838
rect 12532 25774 12584 25780
rect 11520 25424 11572 25430
rect 11520 25366 11572 25372
rect 11980 25424 12032 25430
rect 11980 25366 12032 25372
rect 11336 25288 11388 25294
rect 11336 25230 11388 25236
rect 11348 24818 11376 25230
rect 11520 24880 11572 24886
rect 11520 24822 11572 24828
rect 11336 24812 11388 24818
rect 11336 24754 11388 24760
rect 11532 24750 11560 24822
rect 11428 24744 11480 24750
rect 11428 24686 11480 24692
rect 11520 24744 11572 24750
rect 11520 24686 11572 24692
rect 11440 23798 11468 24686
rect 11888 24676 11940 24682
rect 11888 24618 11940 24624
rect 11612 24268 11664 24274
rect 11612 24210 11664 24216
rect 11244 23792 11296 23798
rect 11244 23734 11296 23740
rect 11428 23792 11480 23798
rect 11428 23734 11480 23740
rect 11256 23186 11284 23734
rect 11244 23180 11296 23186
rect 11244 23122 11296 23128
rect 11060 23112 11112 23118
rect 11060 23054 11112 23060
rect 11624 22506 11652 24210
rect 11796 23724 11848 23730
rect 11796 23666 11848 23672
rect 11704 23656 11756 23662
rect 11704 23598 11756 23604
rect 11612 22500 11664 22506
rect 11612 22442 11664 22448
rect 11152 22432 11204 22438
rect 11152 22374 11204 22380
rect 11244 22432 11296 22438
rect 11244 22374 11296 22380
rect 10968 22160 11020 22166
rect 10968 22102 11020 22108
rect 10876 22092 10928 22098
rect 10876 22034 10928 22040
rect 10324 21956 10376 21962
rect 10324 21898 10376 21904
rect 10232 21548 10284 21554
rect 10232 21490 10284 21496
rect 10336 21486 10364 21898
rect 10324 21480 10376 21486
rect 10324 21422 10376 21428
rect 10888 21418 10916 22034
rect 11060 22024 11112 22030
rect 11060 21966 11112 21972
rect 11072 21690 11100 21966
rect 11060 21684 11112 21690
rect 11060 21626 11112 21632
rect 10876 21412 10928 21418
rect 10876 21354 10928 21360
rect 10968 21412 11020 21418
rect 10968 21354 11020 21360
rect 9772 21004 9824 21010
rect 9772 20946 9824 20952
rect 9956 21004 10008 21010
rect 9956 20946 10008 20952
rect 10888 20874 10916 21354
rect 10876 20868 10928 20874
rect 10876 20810 10928 20816
rect 9864 20392 9916 20398
rect 9864 20334 9916 20340
rect 9312 19848 9364 19854
rect 9312 19790 9364 19796
rect 9324 19446 9352 19790
rect 9876 19718 9904 20334
rect 10414 19952 10470 19961
rect 10414 19887 10470 19896
rect 10428 19854 10456 19887
rect 10416 19848 10468 19854
rect 10416 19790 10468 19796
rect 10600 19848 10652 19854
rect 10600 19790 10652 19796
rect 9864 19712 9916 19718
rect 9864 19654 9916 19660
rect 9772 19508 9824 19514
rect 9772 19450 9824 19456
rect 9312 19440 9364 19446
rect 9312 19382 9364 19388
rect 9588 19304 9640 19310
rect 9588 19246 9640 19252
rect 9600 18902 9628 19246
rect 9784 18970 9812 19450
rect 10612 19378 10640 19790
rect 10600 19372 10652 19378
rect 10600 19314 10652 19320
rect 9956 19304 10008 19310
rect 9956 19246 10008 19252
rect 9772 18964 9824 18970
rect 9772 18906 9824 18912
rect 9864 18964 9916 18970
rect 9864 18906 9916 18912
rect 9588 18896 9640 18902
rect 9588 18838 9640 18844
rect 9680 18896 9732 18902
rect 9876 18850 9904 18906
rect 9732 18844 9904 18850
rect 9680 18838 9904 18844
rect 9692 18822 9904 18838
rect 9770 18728 9826 18737
rect 9770 18663 9826 18672
rect 9864 18692 9916 18698
rect 9784 18630 9812 18663
rect 9864 18634 9916 18640
rect 9772 18624 9824 18630
rect 9772 18566 9824 18572
rect 9772 18420 9824 18426
rect 9876 18408 9904 18634
rect 9968 18426 9996 19246
rect 10048 18964 10100 18970
rect 10048 18906 10100 18912
rect 10060 18766 10088 18906
rect 10048 18760 10100 18766
rect 10048 18702 10100 18708
rect 9824 18380 9904 18408
rect 9956 18420 10008 18426
rect 9772 18362 9824 18368
rect 9956 18362 10008 18368
rect 9232 17870 9352 17898
rect 9220 17808 9272 17814
rect 9220 17750 9272 17756
rect 8576 17740 8628 17746
rect 8576 17682 8628 17688
rect 9232 17338 9260 17750
rect 9220 17332 9272 17338
rect 9220 17274 9272 17280
rect 8576 17128 8628 17134
rect 8576 17070 8628 17076
rect 8588 16726 8616 17070
rect 8576 16720 8628 16726
rect 8576 16662 8628 16668
rect 8668 16040 8720 16046
rect 8668 15982 8720 15988
rect 8484 15564 8536 15570
rect 8484 15506 8536 15512
rect 8116 14816 8168 14822
rect 8116 14758 8168 14764
rect 8208 14816 8260 14822
rect 8208 14758 8260 14764
rect 8128 14550 8156 14758
rect 8116 14544 8168 14550
rect 8116 14486 8168 14492
rect 7944 14368 8156 14396
rect 7564 14272 7616 14278
rect 7564 14214 7616 14220
rect 7576 13870 7604 14214
rect 7380 13864 7432 13870
rect 7380 13806 7432 13812
rect 7564 13864 7616 13870
rect 7564 13806 7616 13812
rect 7392 12306 7420 13806
rect 7380 12300 7432 12306
rect 7380 12242 7432 12248
rect 7576 11694 7604 13806
rect 7656 13796 7708 13802
rect 7656 13738 7708 13744
rect 7668 13394 7696 13738
rect 7656 13388 7708 13394
rect 7656 13330 7708 13336
rect 7656 13184 7708 13190
rect 7656 13126 7708 13132
rect 7668 12782 7696 13126
rect 7656 12776 7708 12782
rect 7656 12718 7708 12724
rect 7932 12776 7984 12782
rect 7932 12718 7984 12724
rect 7944 12306 7972 12718
rect 7932 12300 7984 12306
rect 7932 12242 7984 12248
rect 8024 12300 8076 12306
rect 8024 12242 8076 12248
rect 7564 11688 7616 11694
rect 7564 11630 7616 11636
rect 7944 11626 7972 12242
rect 7932 11620 7984 11626
rect 7932 11562 7984 11568
rect 8036 11218 8064 12242
rect 8024 11212 8076 11218
rect 8024 11154 8076 11160
rect 7472 11008 7524 11014
rect 7472 10950 7524 10956
rect 7300 9574 7420 9602
rect 7288 9512 7340 9518
rect 7288 9454 7340 9460
rect 7104 9036 7156 9042
rect 7104 8978 7156 8984
rect 7116 8430 7144 8978
rect 7300 8974 7328 9454
rect 7288 8968 7340 8974
rect 7288 8910 7340 8916
rect 7196 8492 7248 8498
rect 7196 8434 7248 8440
rect 7104 8424 7156 8430
rect 7104 8366 7156 8372
rect 7116 7546 7144 8366
rect 7208 7954 7236 8434
rect 7196 7948 7248 7954
rect 7196 7890 7248 7896
rect 7104 7540 7156 7546
rect 7104 7482 7156 7488
rect 7012 6724 7064 6730
rect 7012 6666 7064 6672
rect 6920 5772 6972 5778
rect 6920 5714 6972 5720
rect 6828 5160 6880 5166
rect 6828 5102 6880 5108
rect 6932 4826 6960 5714
rect 7024 5642 7052 6666
rect 7116 6254 7144 7482
rect 7104 6248 7156 6254
rect 7104 6190 7156 6196
rect 7116 5778 7144 6190
rect 7104 5772 7156 5778
rect 7104 5714 7156 5720
rect 7012 5636 7064 5642
rect 7012 5578 7064 5584
rect 7288 5636 7340 5642
rect 7288 5578 7340 5584
rect 7300 5234 7328 5578
rect 7288 5228 7340 5234
rect 7288 5170 7340 5176
rect 6920 4820 6972 4826
rect 6920 4762 6972 4768
rect 6920 4616 6972 4622
rect 6920 4558 6972 4564
rect 6932 3942 6960 4558
rect 7012 4480 7064 4486
rect 7012 4422 7064 4428
rect 6920 3936 6972 3942
rect 6920 3878 6972 3884
rect 7024 3754 7052 4422
rect 7104 4072 7156 4078
rect 7102 4040 7104 4049
rect 7156 4040 7158 4049
rect 7102 3975 7158 3984
rect 6932 3726 7052 3754
rect 7392 3738 7420 9574
rect 7484 7342 7512 10950
rect 7564 10804 7616 10810
rect 7564 10746 7616 10752
rect 7472 7336 7524 7342
rect 7472 7278 7524 7284
rect 7472 6792 7524 6798
rect 7472 6734 7524 6740
rect 7484 6322 7512 6734
rect 7576 6662 7604 10746
rect 7656 10600 7708 10606
rect 7656 10542 7708 10548
rect 7668 10266 7696 10542
rect 7656 10260 7708 10266
rect 7656 10202 7708 10208
rect 8128 9908 8156 14368
rect 8220 13870 8248 14758
rect 8680 14414 8708 15982
rect 8852 15496 8904 15502
rect 8852 15438 8904 15444
rect 8668 14408 8720 14414
rect 8668 14350 8720 14356
rect 8208 13864 8260 13870
rect 8208 13806 8260 13812
rect 8300 13728 8352 13734
rect 8300 13670 8352 13676
rect 8312 13394 8340 13670
rect 8864 13394 8892 15438
rect 9036 15360 9088 15366
rect 9036 15302 9088 15308
rect 9048 14958 9076 15302
rect 9220 15156 9272 15162
rect 9220 15098 9272 15104
rect 9232 14958 9260 15098
rect 9036 14952 9088 14958
rect 9036 14894 9088 14900
rect 9220 14952 9272 14958
rect 9220 14894 9272 14900
rect 8944 14884 8996 14890
rect 8944 14826 8996 14832
rect 8956 14793 8984 14826
rect 8942 14784 8998 14793
rect 8942 14719 8998 14728
rect 9048 14482 9076 14894
rect 9036 14476 9088 14482
rect 9036 14418 9088 14424
rect 8944 14068 8996 14074
rect 8944 14010 8996 14016
rect 8300 13388 8352 13394
rect 8852 13388 8904 13394
rect 8352 13348 8432 13376
rect 8300 13330 8352 13336
rect 8300 12912 8352 12918
rect 8300 12854 8352 12860
rect 8208 12776 8260 12782
rect 8208 12718 8260 12724
rect 8220 10062 8248 12718
rect 8312 11762 8340 12854
rect 8404 12782 8432 13348
rect 8852 13330 8904 13336
rect 8392 12776 8444 12782
rect 8392 12718 8444 12724
rect 8300 11756 8352 11762
rect 8300 11698 8352 11704
rect 8484 11688 8536 11694
rect 8484 11630 8536 11636
rect 8496 10674 8524 11630
rect 8484 10668 8536 10674
rect 8484 10610 8536 10616
rect 8852 10600 8904 10606
rect 8852 10542 8904 10548
rect 8668 10532 8720 10538
rect 8668 10474 8720 10480
rect 8208 10056 8260 10062
rect 8208 9998 8260 10004
rect 8576 10056 8628 10062
rect 8576 9998 8628 10004
rect 8128 9880 8248 9908
rect 7748 9580 7800 9586
rect 7748 9522 7800 9528
rect 7760 9042 7788 9522
rect 7748 9036 7800 9042
rect 7748 8978 7800 8984
rect 8116 9036 8168 9042
rect 8116 8978 8168 8984
rect 8128 8430 8156 8978
rect 8116 8424 8168 8430
rect 8116 8366 8168 8372
rect 7840 8016 7892 8022
rect 7840 7958 7892 7964
rect 7852 7478 7880 7958
rect 7840 7472 7892 7478
rect 7840 7414 7892 7420
rect 7564 6656 7616 6662
rect 7564 6598 7616 6604
rect 7472 6316 7524 6322
rect 7472 6258 7524 6264
rect 7852 6254 7880 7414
rect 8128 6458 8156 8366
rect 8116 6452 8168 6458
rect 8116 6394 8168 6400
rect 8128 6254 8156 6394
rect 7840 6248 7892 6254
rect 7840 6190 7892 6196
rect 8116 6248 8168 6254
rect 8116 6190 8168 6196
rect 8128 5778 8156 6190
rect 8220 5846 8248 9880
rect 8300 7336 8352 7342
rect 8300 7278 8352 7284
rect 8392 7336 8444 7342
rect 8392 7278 8444 7284
rect 8312 7002 8340 7278
rect 8300 6996 8352 7002
rect 8300 6938 8352 6944
rect 8300 6248 8352 6254
rect 8300 6190 8352 6196
rect 8312 6118 8340 6190
rect 8300 6112 8352 6118
rect 8300 6054 8352 6060
rect 8404 5846 8432 7278
rect 8208 5840 8260 5846
rect 8208 5782 8260 5788
rect 8392 5840 8444 5846
rect 8392 5782 8444 5788
rect 8116 5772 8168 5778
rect 8116 5714 8168 5720
rect 8404 5166 8432 5782
rect 8484 5228 8536 5234
rect 8484 5170 8536 5176
rect 8116 5160 8168 5166
rect 8116 5102 8168 5108
rect 8392 5160 8444 5166
rect 8392 5102 8444 5108
rect 8128 4826 8156 5102
rect 8116 4820 8168 4826
rect 8116 4762 8168 4768
rect 8128 4554 8156 4762
rect 8116 4548 8168 4554
rect 8116 4490 8168 4496
rect 8128 4146 8156 4490
rect 8116 4140 8168 4146
rect 8116 4082 8168 4088
rect 8496 4078 8524 5170
rect 8588 4214 8616 9998
rect 8680 8498 8708 10474
rect 8864 10130 8892 10542
rect 8852 10124 8904 10130
rect 8852 10066 8904 10072
rect 8760 9444 8812 9450
rect 8760 9386 8812 9392
rect 8668 8492 8720 8498
rect 8668 8434 8720 8440
rect 8680 8090 8708 8434
rect 8668 8084 8720 8090
rect 8668 8026 8720 8032
rect 8772 5817 8800 9386
rect 8758 5808 8814 5817
rect 8758 5743 8760 5752
rect 8812 5743 8814 5752
rect 8760 5714 8812 5720
rect 8772 5683 8800 5714
rect 8668 4684 8720 4690
rect 8668 4626 8720 4632
rect 8576 4208 8628 4214
rect 8576 4150 8628 4156
rect 8484 4072 8536 4078
rect 8484 4014 8536 4020
rect 7380 3732 7432 3738
rect 6828 3460 6880 3466
rect 6828 3402 6880 3408
rect 6552 3392 6604 3398
rect 6552 3334 6604 3340
rect 6564 3194 6592 3334
rect 6552 3188 6604 3194
rect 6552 3130 6604 3136
rect 5816 2984 5868 2990
rect 5816 2926 5868 2932
rect 6092 2984 6144 2990
rect 6092 2926 6144 2932
rect 5724 2440 5776 2446
rect 5724 2382 5776 2388
rect 4712 2304 4764 2310
rect 4712 2246 4764 2252
rect 4220 2204 4516 2224
rect 4276 2202 4300 2204
rect 4356 2202 4380 2204
rect 4436 2202 4460 2204
rect 4298 2150 4300 2202
rect 4362 2150 4374 2202
rect 4436 2150 4438 2202
rect 4276 2148 4300 2150
rect 4356 2148 4380 2150
rect 4436 2148 4460 2150
rect 4220 2128 4516 2148
rect 4724 1170 4752 2246
rect 4632 1142 4752 1170
rect 4632 800 4660 1142
rect 6840 800 6868 3402
rect 6932 2990 6960 3726
rect 7380 3674 7432 3680
rect 7472 3732 7524 3738
rect 7472 3674 7524 3680
rect 7104 3596 7156 3602
rect 7104 3538 7156 3544
rect 7116 3058 7144 3538
rect 7484 3058 7512 3674
rect 8576 3596 8628 3602
rect 8576 3538 8628 3544
rect 7104 3052 7156 3058
rect 7104 2994 7156 3000
rect 7472 3052 7524 3058
rect 7472 2994 7524 3000
rect 6920 2984 6972 2990
rect 6920 2926 6972 2932
rect 6932 2514 6960 2926
rect 8588 2650 8616 3538
rect 8680 3466 8708 4626
rect 8760 3664 8812 3670
rect 8760 3606 8812 3612
rect 8668 3460 8720 3466
rect 8668 3402 8720 3408
rect 8576 2644 8628 2650
rect 8576 2586 8628 2592
rect 6920 2508 6972 2514
rect 6920 2450 6972 2456
rect 8772 1834 8800 3606
rect 8956 3602 8984 14010
rect 9232 13870 9260 14894
rect 9324 14074 9352 17870
rect 9784 17610 9812 18362
rect 9772 17604 9824 17610
rect 9772 17546 9824 17552
rect 9680 15700 9732 15706
rect 9680 15642 9732 15648
rect 9692 15042 9720 15642
rect 9784 15502 9812 17546
rect 9968 16658 9996 18362
rect 10060 17270 10088 18702
rect 10612 18698 10640 19314
rect 10980 19310 11008 21354
rect 11164 21146 11192 22374
rect 11256 22234 11284 22374
rect 11244 22228 11296 22234
rect 11244 22170 11296 22176
rect 11716 22098 11744 23598
rect 11808 23186 11836 23666
rect 11796 23180 11848 23186
rect 11796 23122 11848 23128
rect 11808 22574 11836 23122
rect 11900 22778 11928 24618
rect 12440 24608 12492 24614
rect 12440 24550 12492 24556
rect 12162 23352 12218 23361
rect 12162 23287 12218 23296
rect 12176 23186 12204 23287
rect 12164 23180 12216 23186
rect 12164 23122 12216 23128
rect 12348 23180 12400 23186
rect 12348 23122 12400 23128
rect 11888 22772 11940 22778
rect 11888 22714 11940 22720
rect 11796 22568 11848 22574
rect 11796 22510 11848 22516
rect 12360 22234 12388 23122
rect 12452 22574 12480 24550
rect 12440 22568 12492 22574
rect 12440 22510 12492 22516
rect 12348 22228 12400 22234
rect 12348 22170 12400 22176
rect 12360 22098 12388 22170
rect 11704 22092 11756 22098
rect 11704 22034 11756 22040
rect 12348 22092 12400 22098
rect 12348 22034 12400 22040
rect 11520 21684 11572 21690
rect 11520 21626 11572 21632
rect 11244 21480 11296 21486
rect 11244 21422 11296 21428
rect 11152 21140 11204 21146
rect 11152 21082 11204 21088
rect 10968 19304 11020 19310
rect 10968 19246 11020 19252
rect 11060 18760 11112 18766
rect 11060 18702 11112 18708
rect 10600 18692 10652 18698
rect 10600 18634 10652 18640
rect 10324 18352 10376 18358
rect 10324 18294 10376 18300
rect 10232 18216 10284 18222
rect 10232 18158 10284 18164
rect 10244 17338 10272 18158
rect 10336 17882 10364 18294
rect 10416 18080 10468 18086
rect 10416 18022 10468 18028
rect 10324 17876 10376 17882
rect 10324 17818 10376 17824
rect 10428 17746 10456 18022
rect 11072 17814 11100 18702
rect 11060 17808 11112 17814
rect 11060 17750 11112 17756
rect 10416 17740 10468 17746
rect 10416 17682 10468 17688
rect 11256 17678 11284 21422
rect 11336 20392 11388 20398
rect 11336 20334 11388 20340
rect 11348 20058 11376 20334
rect 11336 20052 11388 20058
rect 11336 19994 11388 20000
rect 11348 19514 11376 19994
rect 11532 19922 11560 21626
rect 12544 21554 12572 25774
rect 12808 25356 12860 25362
rect 12808 25298 12860 25304
rect 12624 25288 12676 25294
rect 12624 25230 12676 25236
rect 12636 24138 12664 25230
rect 12624 24132 12676 24138
rect 12624 24074 12676 24080
rect 12716 23656 12768 23662
rect 12716 23598 12768 23604
rect 12624 23248 12676 23254
rect 12624 23190 12676 23196
rect 12532 21548 12584 21554
rect 12532 21490 12584 21496
rect 12256 21344 12308 21350
rect 12256 21286 12308 21292
rect 11704 20392 11756 20398
rect 11704 20334 11756 20340
rect 11716 20058 11744 20334
rect 11704 20052 11756 20058
rect 11704 19994 11756 20000
rect 11520 19916 11572 19922
rect 11520 19858 11572 19864
rect 11336 19508 11388 19514
rect 11336 19450 11388 19456
rect 12268 19310 12296 21286
rect 12544 21146 12572 21490
rect 12636 21486 12664 23190
rect 12728 22778 12756 23598
rect 12716 22772 12768 22778
rect 12716 22714 12768 22720
rect 12624 21480 12676 21486
rect 12624 21422 12676 21428
rect 12532 21140 12584 21146
rect 12532 21082 12584 21088
rect 12544 21010 12572 21082
rect 12532 21004 12584 21010
rect 12532 20946 12584 20952
rect 12716 20392 12768 20398
rect 12716 20334 12768 20340
rect 12256 19304 12308 19310
rect 12256 19246 12308 19252
rect 12268 18154 12296 19246
rect 12440 19236 12492 19242
rect 12440 19178 12492 19184
rect 12452 18442 12480 19178
rect 12728 18766 12756 20334
rect 12820 20058 12848 25298
rect 12912 22710 12940 26982
rect 13544 26920 13596 26926
rect 13544 26862 13596 26868
rect 13268 26308 13320 26314
rect 13268 26250 13320 26256
rect 13084 25900 13136 25906
rect 13084 25842 13136 25848
rect 12992 24336 13044 24342
rect 12990 24304 12992 24313
rect 13044 24304 13046 24313
rect 12990 24239 13046 24248
rect 12900 22704 12952 22710
rect 12900 22646 12952 22652
rect 13096 21418 13124 25842
rect 13176 25764 13228 25770
rect 13176 25706 13228 25712
rect 13188 22574 13216 25706
rect 13280 25362 13308 26250
rect 13268 25356 13320 25362
rect 13268 25298 13320 25304
rect 13176 22568 13228 22574
rect 13176 22510 13228 22516
rect 13556 22234 13584 26862
rect 13544 22228 13596 22234
rect 13544 22170 13596 22176
rect 13176 22092 13228 22098
rect 13176 22034 13228 22040
rect 13188 21554 13216 22034
rect 13176 21548 13228 21554
rect 13176 21490 13228 21496
rect 13084 21412 13136 21418
rect 13084 21354 13136 21360
rect 13096 21010 13124 21354
rect 13084 21004 13136 21010
rect 13084 20946 13136 20952
rect 13096 20806 13124 20946
rect 13084 20800 13136 20806
rect 13084 20742 13136 20748
rect 12900 20528 12952 20534
rect 12900 20470 12952 20476
rect 12808 20052 12860 20058
rect 12808 19994 12860 20000
rect 12912 19922 12940 20470
rect 13084 20460 13136 20466
rect 13084 20402 13136 20408
rect 12992 20392 13044 20398
rect 12992 20334 13044 20340
rect 13004 20058 13032 20334
rect 12992 20052 13044 20058
rect 12992 19994 13044 20000
rect 12900 19916 12952 19922
rect 12900 19858 12952 19864
rect 12808 19304 12860 19310
rect 12808 19246 12860 19252
rect 12820 18902 12848 19246
rect 12808 18896 12860 18902
rect 12808 18838 12860 18844
rect 13096 18766 13124 20402
rect 13544 20324 13596 20330
rect 13544 20266 13596 20272
rect 13360 20052 13412 20058
rect 13360 19994 13412 20000
rect 13176 19304 13228 19310
rect 13176 19246 13228 19252
rect 12716 18760 12768 18766
rect 12716 18702 12768 18708
rect 13084 18760 13136 18766
rect 13084 18702 13136 18708
rect 12360 18426 12572 18442
rect 12348 18420 12572 18426
rect 12400 18414 12572 18420
rect 12348 18362 12400 18368
rect 12256 18148 12308 18154
rect 12256 18090 12308 18096
rect 12440 18080 12492 18086
rect 12440 18022 12492 18028
rect 11244 17672 11296 17678
rect 11244 17614 11296 17620
rect 11612 17672 11664 17678
rect 11612 17614 11664 17620
rect 10232 17332 10284 17338
rect 10232 17274 10284 17280
rect 10048 17264 10100 17270
rect 10048 17206 10100 17212
rect 11256 17202 11284 17614
rect 11624 17338 11652 17614
rect 11612 17332 11664 17338
rect 11612 17274 11664 17280
rect 11244 17196 11296 17202
rect 11244 17138 11296 17144
rect 10692 17128 10744 17134
rect 10692 17070 10744 17076
rect 9956 16652 10008 16658
rect 9956 16594 10008 16600
rect 9772 15496 9824 15502
rect 9772 15438 9824 15444
rect 9508 15026 9720 15042
rect 9496 15020 9720 15026
rect 9548 15014 9720 15020
rect 9496 14962 9548 14968
rect 9588 14952 9640 14958
rect 9588 14894 9640 14900
rect 9312 14068 9364 14074
rect 9312 14010 9364 14016
rect 9600 13870 9628 14894
rect 9968 14346 9996 16594
rect 10048 16448 10100 16454
rect 10048 16390 10100 16396
rect 9956 14340 10008 14346
rect 9956 14282 10008 14288
rect 10060 13938 10088 16390
rect 10416 15564 10468 15570
rect 10416 15506 10468 15512
rect 10232 15428 10284 15434
rect 10232 15370 10284 15376
rect 10140 15360 10192 15366
rect 10140 15302 10192 15308
rect 10048 13932 10100 13938
rect 10048 13874 10100 13880
rect 9220 13864 9272 13870
rect 9220 13806 9272 13812
rect 9588 13864 9640 13870
rect 9588 13806 9640 13812
rect 9864 13796 9916 13802
rect 9864 13738 9916 13744
rect 9588 13728 9640 13734
rect 9588 13670 9640 13676
rect 9312 13320 9364 13326
rect 9312 13262 9364 13268
rect 9220 13252 9272 13258
rect 9220 13194 9272 13200
rect 9232 12782 9260 13194
rect 9324 12918 9352 13262
rect 9312 12912 9364 12918
rect 9312 12854 9364 12860
rect 9600 12850 9628 13670
rect 9876 13394 9904 13738
rect 10060 13394 10088 13874
rect 10152 13870 10180 15302
rect 10244 14482 10272 15370
rect 10428 14822 10456 15506
rect 10508 15496 10560 15502
rect 10508 15438 10560 15444
rect 10416 14816 10468 14822
rect 10322 14784 10378 14793
rect 10416 14758 10468 14764
rect 10322 14719 10378 14728
rect 10336 14550 10364 14719
rect 10324 14544 10376 14550
rect 10324 14486 10376 14492
rect 10520 14482 10548 15438
rect 10600 14952 10652 14958
rect 10600 14894 10652 14900
rect 10612 14482 10640 14894
rect 10232 14476 10284 14482
rect 10232 14418 10284 14424
rect 10508 14476 10560 14482
rect 10508 14418 10560 14424
rect 10600 14476 10652 14482
rect 10600 14418 10652 14424
rect 10140 13864 10192 13870
rect 10140 13806 10192 13812
rect 9864 13388 9916 13394
rect 9864 13330 9916 13336
rect 10048 13388 10100 13394
rect 10048 13330 10100 13336
rect 9680 13184 9732 13190
rect 9680 13126 9732 13132
rect 9588 12844 9640 12850
rect 9588 12786 9640 12792
rect 9220 12776 9272 12782
rect 9220 12718 9272 12724
rect 9036 11280 9088 11286
rect 9036 11222 9088 11228
rect 9048 10810 9076 11222
rect 9036 10804 9088 10810
rect 9036 10746 9088 10752
rect 9048 10674 9076 10746
rect 9036 10668 9088 10674
rect 9036 10610 9088 10616
rect 9600 10062 9628 12786
rect 9692 11694 9720 13126
rect 9680 11688 9732 11694
rect 9680 11630 9732 11636
rect 9680 11552 9732 11558
rect 9680 11494 9732 11500
rect 9588 10056 9640 10062
rect 9588 9998 9640 10004
rect 9692 9994 9720 11494
rect 9772 11212 9824 11218
rect 9772 11154 9824 11160
rect 9680 9988 9732 9994
rect 9680 9930 9732 9936
rect 9036 9036 9088 9042
rect 9036 8978 9088 8984
rect 9048 8430 9076 8978
rect 9036 8424 9088 8430
rect 9036 8366 9088 8372
rect 9680 8424 9732 8430
rect 9680 8366 9732 8372
rect 9692 6390 9720 8366
rect 9680 6384 9732 6390
rect 9680 6326 9732 6332
rect 9692 5794 9720 6326
rect 9600 5778 9720 5794
rect 9784 5778 9812 11154
rect 9876 10606 9904 13330
rect 9954 13288 10010 13297
rect 9954 13223 10010 13232
rect 9968 12170 9996 13223
rect 10140 12300 10192 12306
rect 10140 12242 10192 12248
rect 10324 12300 10376 12306
rect 10324 12242 10376 12248
rect 10508 12300 10560 12306
rect 10508 12242 10560 12248
rect 9956 12164 10008 12170
rect 9956 12106 10008 12112
rect 10152 11830 10180 12242
rect 10140 11824 10192 11830
rect 10140 11766 10192 11772
rect 10048 11688 10100 11694
rect 10048 11630 10100 11636
rect 9956 11552 10008 11558
rect 9956 11494 10008 11500
rect 9864 10600 9916 10606
rect 9864 10542 9916 10548
rect 9876 8430 9904 10542
rect 9968 9518 9996 11494
rect 10060 11218 10088 11630
rect 10048 11212 10100 11218
rect 10048 11154 10100 11160
rect 9956 9512 10008 9518
rect 9956 9454 10008 9460
rect 10152 9042 10180 11766
rect 10336 11762 10364 12242
rect 10520 11762 10548 12242
rect 10324 11756 10376 11762
rect 10324 11698 10376 11704
rect 10508 11756 10560 11762
rect 10508 11698 10560 11704
rect 10324 11348 10376 11354
rect 10324 11290 10376 11296
rect 10140 9036 10192 9042
rect 10140 8978 10192 8984
rect 9864 8424 9916 8430
rect 9864 8366 9916 8372
rect 10048 7948 10100 7954
rect 10048 7890 10100 7896
rect 9956 7880 10008 7886
rect 9956 7822 10008 7828
rect 9968 7410 9996 7822
rect 9956 7404 10008 7410
rect 9956 7346 10008 7352
rect 9864 7336 9916 7342
rect 9864 7278 9916 7284
rect 9876 6458 9904 7278
rect 9864 6452 9916 6458
rect 9864 6394 9916 6400
rect 9864 6248 9916 6254
rect 9864 6190 9916 6196
rect 9588 5772 9720 5778
rect 9640 5766 9720 5772
rect 9772 5772 9824 5778
rect 9588 5714 9640 5720
rect 9772 5714 9824 5720
rect 9784 5370 9812 5714
rect 9772 5364 9824 5370
rect 9772 5306 9824 5312
rect 9876 5234 9904 6190
rect 9864 5228 9916 5234
rect 9864 5170 9916 5176
rect 9680 5160 9732 5166
rect 9680 5102 9732 5108
rect 9692 4690 9720 5102
rect 9680 4684 9732 4690
rect 9680 4626 9732 4632
rect 9128 4616 9180 4622
rect 9128 4558 9180 4564
rect 8944 3596 8996 3602
rect 8944 3538 8996 3544
rect 9140 3058 9168 4558
rect 10060 4554 10088 7890
rect 10336 7002 10364 11290
rect 10704 10810 10732 17070
rect 11256 16998 11284 17138
rect 11428 17128 11480 17134
rect 11428 17070 11480 17076
rect 11244 16992 11296 16998
rect 11244 16934 11296 16940
rect 11440 16794 11468 17070
rect 11428 16788 11480 16794
rect 11428 16730 11480 16736
rect 10784 16448 10836 16454
rect 10784 16390 10836 16396
rect 10796 16114 10824 16390
rect 10784 16108 10836 16114
rect 10784 16050 10836 16056
rect 11520 16040 11572 16046
rect 11520 15982 11572 15988
rect 11060 15564 11112 15570
rect 11060 15506 11112 15512
rect 11072 15162 11100 15506
rect 11060 15156 11112 15162
rect 11060 15098 11112 15104
rect 10784 14952 10836 14958
rect 10784 14894 10836 14900
rect 11428 14952 11480 14958
rect 11428 14894 11480 14900
rect 10796 11218 10824 14894
rect 10968 14816 11020 14822
rect 10968 14758 11020 14764
rect 10980 13802 11008 14758
rect 11440 14074 11468 14894
rect 11532 14618 11560 15982
rect 11612 15904 11664 15910
rect 11612 15846 11664 15852
rect 11624 15638 11652 15846
rect 11612 15632 11664 15638
rect 11612 15574 11664 15580
rect 11520 14612 11572 14618
rect 11520 14554 11572 14560
rect 11428 14068 11480 14074
rect 11428 14010 11480 14016
rect 11520 13864 11572 13870
rect 11520 13806 11572 13812
rect 10968 13796 11020 13802
rect 10968 13738 11020 13744
rect 10980 13326 11008 13738
rect 11244 13456 11296 13462
rect 11244 13398 11296 13404
rect 10968 13320 11020 13326
rect 10968 13262 11020 13268
rect 10968 13184 11020 13190
rect 10968 13126 11020 13132
rect 10980 12782 11008 13126
rect 11256 12782 11284 13398
rect 11532 13394 11560 13806
rect 11520 13388 11572 13394
rect 11520 13330 11572 13336
rect 10968 12776 11020 12782
rect 10968 12718 11020 12724
rect 11244 12776 11296 12782
rect 11244 12718 11296 12724
rect 11428 12776 11480 12782
rect 11428 12718 11480 12724
rect 11256 11558 11284 12718
rect 11440 11762 11468 12718
rect 11428 11756 11480 11762
rect 11428 11698 11480 11704
rect 11336 11688 11388 11694
rect 11336 11630 11388 11636
rect 11244 11552 11296 11558
rect 11244 11494 11296 11500
rect 10784 11212 10836 11218
rect 10784 11154 10836 11160
rect 10968 11076 11020 11082
rect 10968 11018 11020 11024
rect 10692 10804 10744 10810
rect 10692 10746 10744 10752
rect 10980 10674 11008 11018
rect 10968 10668 11020 10674
rect 10968 10610 11020 10616
rect 10508 10124 10560 10130
rect 10508 10066 10560 10072
rect 10784 10124 10836 10130
rect 10784 10066 10836 10072
rect 10520 9926 10548 10066
rect 10508 9920 10560 9926
rect 10508 9862 10560 9868
rect 10324 6996 10376 7002
rect 10324 6938 10376 6944
rect 10140 5568 10192 5574
rect 10140 5510 10192 5516
rect 10048 4548 10100 4554
rect 10048 4490 10100 4496
rect 9220 4140 9272 4146
rect 9220 4082 9272 4088
rect 9232 3913 9260 4082
rect 9312 4072 9364 4078
rect 9310 4040 9312 4049
rect 9364 4040 9366 4049
rect 9310 3975 9366 3984
rect 10048 3936 10100 3942
rect 9218 3904 9274 3913
rect 10048 3878 10100 3884
rect 9218 3839 9274 3848
rect 10060 3466 10088 3878
rect 10152 3602 10180 5510
rect 10336 5166 10364 6938
rect 10520 6866 10548 9862
rect 10796 9654 10824 10066
rect 10784 9648 10836 9654
rect 10784 9590 10836 9596
rect 10980 9518 11008 10610
rect 10784 9512 10836 9518
rect 10612 9472 10784 9500
rect 10612 9382 10640 9472
rect 10784 9454 10836 9460
rect 10968 9512 11020 9518
rect 10968 9454 11020 9460
rect 10600 9376 10652 9382
rect 10600 9318 10652 9324
rect 11152 8968 11204 8974
rect 11152 8910 11204 8916
rect 10600 8424 10652 8430
rect 10600 8366 10652 8372
rect 10612 7274 10640 8366
rect 11060 7812 11112 7818
rect 11060 7754 11112 7760
rect 10784 7336 10836 7342
rect 10784 7278 10836 7284
rect 10600 7268 10652 7274
rect 10600 7210 10652 7216
rect 10508 6860 10560 6866
rect 10508 6802 10560 6808
rect 10796 6390 10824 7278
rect 11072 6866 11100 7754
rect 11060 6860 11112 6866
rect 11060 6802 11112 6808
rect 11164 6798 11192 8910
rect 11244 8424 11296 8430
rect 11244 8366 11296 8372
rect 11256 7546 11284 8366
rect 11244 7540 11296 7546
rect 11244 7482 11296 7488
rect 11152 6792 11204 6798
rect 11152 6734 11204 6740
rect 10784 6384 10836 6390
rect 10784 6326 10836 6332
rect 10600 6248 10652 6254
rect 10600 6190 10652 6196
rect 11152 6248 11204 6254
rect 11152 6190 11204 6196
rect 10508 5704 10560 5710
rect 10508 5646 10560 5652
rect 10416 5636 10468 5642
rect 10416 5578 10468 5584
rect 10428 5234 10456 5578
rect 10416 5228 10468 5234
rect 10416 5170 10468 5176
rect 10324 5160 10376 5166
rect 10324 5102 10376 5108
rect 10520 4690 10548 5646
rect 10612 5234 10640 6190
rect 10876 6180 10928 6186
rect 10876 6122 10928 6128
rect 10600 5228 10652 5234
rect 10600 5170 10652 5176
rect 10324 4684 10376 4690
rect 10508 4684 10560 4690
rect 10376 4644 10456 4672
rect 10324 4626 10376 4632
rect 10324 4004 10376 4010
rect 10324 3946 10376 3952
rect 10336 3670 10364 3946
rect 10428 3670 10456 4644
rect 10508 4626 10560 4632
rect 10324 3664 10376 3670
rect 10324 3606 10376 3612
rect 10416 3664 10468 3670
rect 10416 3606 10468 3612
rect 10140 3596 10192 3602
rect 10140 3538 10192 3544
rect 10416 3528 10468 3534
rect 10416 3470 10468 3476
rect 10048 3460 10100 3466
rect 10048 3402 10100 3408
rect 9128 3052 9180 3058
rect 9128 2994 9180 3000
rect 10428 2990 10456 3470
rect 10888 3194 10916 6122
rect 11060 5772 11112 5778
rect 11060 5714 11112 5720
rect 11072 5370 11100 5714
rect 11060 5364 11112 5370
rect 11060 5306 11112 5312
rect 11164 3466 11192 6190
rect 11256 4826 11284 7482
rect 11244 4820 11296 4826
rect 11244 4762 11296 4768
rect 11348 4298 11376 11630
rect 11624 11218 11652 15574
rect 11704 15564 11756 15570
rect 11704 15506 11756 15512
rect 11716 15473 11744 15506
rect 11702 15464 11758 15473
rect 11702 15399 11758 15408
rect 11716 15094 11744 15399
rect 11796 15156 11848 15162
rect 11796 15098 11848 15104
rect 11704 15088 11756 15094
rect 11704 15030 11756 15036
rect 11808 14822 11836 15098
rect 11704 14816 11756 14822
rect 11702 14784 11704 14793
rect 11796 14816 11848 14822
rect 11756 14784 11758 14793
rect 11796 14758 11848 14764
rect 11702 14719 11758 14728
rect 11888 14612 11940 14618
rect 11888 14554 11940 14560
rect 11900 13870 11928 14554
rect 12452 14006 12480 18022
rect 12544 16590 12572 18414
rect 12624 18216 12676 18222
rect 12624 18158 12676 18164
rect 12532 16584 12584 16590
rect 12532 16526 12584 16532
rect 12544 15978 12572 16526
rect 12532 15972 12584 15978
rect 12532 15914 12584 15920
rect 12544 15570 12572 15914
rect 12636 15706 12664 18158
rect 12728 17134 12756 18702
rect 13084 17876 13136 17882
rect 13084 17818 13136 17824
rect 12900 17536 12952 17542
rect 12900 17478 12952 17484
rect 12912 17134 12940 17478
rect 12716 17128 12768 17134
rect 12716 17070 12768 17076
rect 12900 17128 12952 17134
rect 12900 17070 12952 17076
rect 12728 16794 12756 17070
rect 12716 16788 12768 16794
rect 12716 16730 12768 16736
rect 13096 16590 13124 17818
rect 13084 16584 13136 16590
rect 13084 16526 13136 16532
rect 13084 16176 13136 16182
rect 13004 16136 13084 16164
rect 12900 16040 12952 16046
rect 12900 15982 12952 15988
rect 12624 15700 12676 15706
rect 12624 15642 12676 15648
rect 12808 15632 12860 15638
rect 12912 15620 12940 15982
rect 12860 15592 12940 15620
rect 12808 15574 12860 15580
rect 13004 15570 13032 16136
rect 13084 16118 13136 16124
rect 13084 16040 13136 16046
rect 13084 15982 13136 15988
rect 13096 15570 13124 15982
rect 12532 15564 12584 15570
rect 12532 15506 12584 15512
rect 12992 15564 13044 15570
rect 12992 15506 13044 15512
rect 13084 15564 13136 15570
rect 13084 15506 13136 15512
rect 12622 15056 12678 15065
rect 12622 14991 12678 15000
rect 12636 14958 12664 14991
rect 12624 14952 12676 14958
rect 12624 14894 12676 14900
rect 12532 14340 12584 14346
rect 12532 14282 12584 14288
rect 12440 14000 12492 14006
rect 12440 13942 12492 13948
rect 11888 13864 11940 13870
rect 11888 13806 11940 13812
rect 11980 13388 12032 13394
rect 11980 13330 12032 13336
rect 11704 11688 11756 11694
rect 11704 11630 11756 11636
rect 11716 11286 11744 11630
rect 11704 11280 11756 11286
rect 11704 11222 11756 11228
rect 11612 11212 11664 11218
rect 11612 11154 11664 11160
rect 11716 10606 11744 11222
rect 11992 10674 12020 13330
rect 12256 13320 12308 13326
rect 12256 13262 12308 13268
rect 12268 12374 12296 13262
rect 12348 12776 12400 12782
rect 12348 12718 12400 12724
rect 12256 12368 12308 12374
rect 12256 12310 12308 12316
rect 12360 11898 12388 12718
rect 12348 11892 12400 11898
rect 12348 11834 12400 11840
rect 12072 11212 12124 11218
rect 12072 11154 12124 11160
rect 12164 11212 12216 11218
rect 12164 11154 12216 11160
rect 12084 10674 12112 11154
rect 11980 10668 12032 10674
rect 11980 10610 12032 10616
rect 12072 10668 12124 10674
rect 12072 10610 12124 10616
rect 11428 10600 11480 10606
rect 11428 10542 11480 10548
rect 11704 10600 11756 10606
rect 11704 10542 11756 10548
rect 11440 5166 11468 10542
rect 12084 9926 12112 10610
rect 12072 9920 12124 9926
rect 12072 9862 12124 9868
rect 12072 8424 12124 8430
rect 12072 8366 12124 8372
rect 12084 7954 12112 8366
rect 12072 7948 12124 7954
rect 12072 7890 12124 7896
rect 11980 7812 12032 7818
rect 11980 7754 12032 7760
rect 11520 7744 11572 7750
rect 11520 7686 11572 7692
rect 11532 7342 11560 7686
rect 11992 7410 12020 7754
rect 12084 7410 12112 7890
rect 11980 7404 12032 7410
rect 11980 7346 12032 7352
rect 12072 7404 12124 7410
rect 12072 7346 12124 7352
rect 11520 7336 11572 7342
rect 11520 7278 11572 7284
rect 12072 6792 12124 6798
rect 12072 6734 12124 6740
rect 11796 6724 11848 6730
rect 11796 6666 11848 6672
rect 11704 6180 11756 6186
rect 11704 6122 11756 6128
rect 11520 5908 11572 5914
rect 11520 5850 11572 5856
rect 11532 5778 11560 5850
rect 11520 5772 11572 5778
rect 11520 5714 11572 5720
rect 11532 5681 11560 5714
rect 11518 5672 11574 5681
rect 11518 5607 11574 5616
rect 11520 5364 11572 5370
rect 11520 5306 11572 5312
rect 11428 5160 11480 5166
rect 11428 5102 11480 5108
rect 11440 4826 11468 5102
rect 11428 4820 11480 4826
rect 11428 4762 11480 4768
rect 11256 4270 11376 4298
rect 11256 4078 11284 4270
rect 11532 4078 11560 5306
rect 11244 4072 11296 4078
rect 11244 4014 11296 4020
rect 11520 4072 11572 4078
rect 11520 4014 11572 4020
rect 11256 3602 11284 4014
rect 11244 3596 11296 3602
rect 11244 3538 11296 3544
rect 11152 3460 11204 3466
rect 11152 3402 11204 3408
rect 10876 3188 10928 3194
rect 10876 3130 10928 3136
rect 11060 3188 11112 3194
rect 11060 3130 11112 3136
rect 10416 2984 10468 2990
rect 10416 2926 10468 2932
rect 10428 2514 10456 2926
rect 11072 2514 11100 3130
rect 11164 2990 11192 3402
rect 11716 3126 11744 6122
rect 11808 4826 11836 6666
rect 12084 6390 12112 6734
rect 12072 6384 12124 6390
rect 12072 6326 12124 6332
rect 12176 5914 12204 11154
rect 12452 10606 12480 13942
rect 12544 13870 12572 14282
rect 12532 13864 12584 13870
rect 12532 13806 12584 13812
rect 12532 13456 12584 13462
rect 12532 13398 12584 13404
rect 12544 12782 12572 13398
rect 12532 12776 12584 12782
rect 12532 12718 12584 12724
rect 12636 10742 12664 14894
rect 12992 14340 13044 14346
rect 12992 14282 13044 14288
rect 12900 12776 12952 12782
rect 12900 12718 12952 12724
rect 12912 12442 12940 12718
rect 12900 12436 12952 12442
rect 12900 12378 12952 12384
rect 12912 12306 12940 12378
rect 12900 12300 12952 12306
rect 12900 12242 12952 12248
rect 13004 12186 13032 14282
rect 12912 12170 13032 12186
rect 12900 12164 13032 12170
rect 12952 12158 13032 12164
rect 12900 12106 12952 12112
rect 12716 11824 12768 11830
rect 12714 11792 12716 11801
rect 12768 11792 12770 11801
rect 12714 11727 12770 11736
rect 12624 10736 12676 10742
rect 12624 10678 12676 10684
rect 12440 10600 12492 10606
rect 12440 10542 12492 10548
rect 12348 10532 12400 10538
rect 12348 10474 12400 10480
rect 12716 10532 12768 10538
rect 12716 10474 12768 10480
rect 12256 9512 12308 9518
rect 12256 9454 12308 9460
rect 12268 8974 12296 9454
rect 12360 9042 12388 10474
rect 12624 10464 12676 10470
rect 12624 10406 12676 10412
rect 12532 10124 12584 10130
rect 12532 10066 12584 10072
rect 12544 9586 12572 10066
rect 12636 9908 12664 10406
rect 12728 10198 12756 10474
rect 12716 10192 12768 10198
rect 12716 10134 12768 10140
rect 12808 9988 12860 9994
rect 12808 9930 12860 9936
rect 12716 9920 12768 9926
rect 12636 9880 12716 9908
rect 12716 9862 12768 9868
rect 12532 9580 12584 9586
rect 12532 9522 12584 9528
rect 12440 9376 12492 9382
rect 12440 9318 12492 9324
rect 12348 9036 12400 9042
rect 12348 8978 12400 8984
rect 12256 8968 12308 8974
rect 12256 8910 12308 8916
rect 12268 8634 12296 8910
rect 12256 8628 12308 8634
rect 12256 8570 12308 8576
rect 12348 8560 12400 8566
rect 12348 8502 12400 8508
rect 12360 7834 12388 8502
rect 12452 7954 12480 9318
rect 12728 9042 12756 9862
rect 12820 9654 12848 9930
rect 12808 9648 12860 9654
rect 12808 9590 12860 9596
rect 12820 9382 12848 9590
rect 12808 9376 12860 9382
rect 12808 9318 12860 9324
rect 12716 9036 12768 9042
rect 12716 8978 12768 8984
rect 12912 8566 12940 12106
rect 13084 11688 13136 11694
rect 13084 11630 13136 11636
rect 13096 11286 13124 11630
rect 13084 11280 13136 11286
rect 13084 11222 13136 11228
rect 12992 10600 13044 10606
rect 12992 10542 13044 10548
rect 12900 8560 12952 8566
rect 12900 8502 12952 8508
rect 12532 8424 12584 8430
rect 12532 8366 12584 8372
rect 12544 8294 12572 8366
rect 12532 8288 12584 8294
rect 12532 8230 12584 8236
rect 13004 7954 13032 10542
rect 13084 10464 13136 10470
rect 13084 10406 13136 10412
rect 13096 10266 13124 10406
rect 13188 10266 13216 19246
rect 13372 18834 13400 19994
rect 13556 19922 13584 20266
rect 13544 19916 13596 19922
rect 13544 19858 13596 19864
rect 13452 19848 13504 19854
rect 13452 19790 13504 19796
rect 13360 18828 13412 18834
rect 13360 18770 13412 18776
rect 13360 15088 13412 15094
rect 13360 15030 13412 15036
rect 13372 14550 13400 15030
rect 13360 14544 13412 14550
rect 13360 14486 13412 14492
rect 13268 14340 13320 14346
rect 13268 14282 13320 14288
rect 13280 13870 13308 14282
rect 13268 13864 13320 13870
rect 13268 13806 13320 13812
rect 13268 11688 13320 11694
rect 13268 11630 13320 11636
rect 13280 10742 13308 11630
rect 13268 10736 13320 10742
rect 13268 10678 13320 10684
rect 13372 10690 13400 14486
rect 13464 11082 13492 19790
rect 13648 17762 13676 26982
rect 13924 26926 13952 27338
rect 14016 27062 14044 27542
rect 14004 27056 14056 27062
rect 14004 26998 14056 27004
rect 13912 26920 13964 26926
rect 13912 26862 13964 26868
rect 13820 26852 13872 26858
rect 13820 26794 13872 26800
rect 13832 26586 13860 26794
rect 14016 26586 14044 26998
rect 13820 26580 13872 26586
rect 13820 26522 13872 26528
rect 14004 26580 14056 26586
rect 14004 26522 14056 26528
rect 14568 25838 14596 27814
rect 13820 25832 13872 25838
rect 13820 25774 13872 25780
rect 14280 25832 14332 25838
rect 14280 25774 14332 25780
rect 14556 25832 14608 25838
rect 14556 25774 14608 25780
rect 13728 25696 13780 25702
rect 13728 25638 13780 25644
rect 13740 25362 13768 25638
rect 13728 25356 13780 25362
rect 13728 25298 13780 25304
rect 13832 24886 13860 25774
rect 13820 24880 13872 24886
rect 13820 24822 13872 24828
rect 14004 23316 14056 23322
rect 14004 23258 14056 23264
rect 14016 23118 14044 23258
rect 14004 23112 14056 23118
rect 14004 23054 14056 23060
rect 13912 22636 13964 22642
rect 13912 22578 13964 22584
rect 13728 22568 13780 22574
rect 13728 22510 13780 22516
rect 13740 19378 13768 22510
rect 13924 22030 13952 22578
rect 14004 22092 14056 22098
rect 14004 22034 14056 22040
rect 13912 22024 13964 22030
rect 13912 21966 13964 21972
rect 13820 21888 13872 21894
rect 13820 21830 13872 21836
rect 13832 21486 13860 21830
rect 13820 21480 13872 21486
rect 13820 21422 13872 21428
rect 13924 20398 13952 21966
rect 13912 20392 13964 20398
rect 13912 20334 13964 20340
rect 13820 20256 13872 20262
rect 13818 20224 13820 20233
rect 13872 20224 13874 20233
rect 13818 20159 13874 20168
rect 13728 19372 13780 19378
rect 13728 19314 13780 19320
rect 13820 18828 13872 18834
rect 13820 18770 13872 18776
rect 13648 17734 13768 17762
rect 13636 17672 13688 17678
rect 13636 17614 13688 17620
rect 13648 17202 13676 17614
rect 13636 17196 13688 17202
rect 13636 17138 13688 17144
rect 13544 16992 13596 16998
rect 13544 16934 13596 16940
rect 13556 16046 13584 16934
rect 13740 16250 13768 17734
rect 13832 17270 13860 18770
rect 13912 18760 13964 18766
rect 13912 18702 13964 18708
rect 13924 18358 13952 18702
rect 13912 18352 13964 18358
rect 13912 18294 13964 18300
rect 13912 17740 13964 17746
rect 13912 17682 13964 17688
rect 13820 17264 13872 17270
rect 13820 17206 13872 17212
rect 13728 16244 13780 16250
rect 13728 16186 13780 16192
rect 13544 16040 13596 16046
rect 13544 15982 13596 15988
rect 13820 16040 13872 16046
rect 13820 15982 13872 15988
rect 13556 14482 13584 15982
rect 13636 15700 13688 15706
rect 13636 15642 13688 15648
rect 13648 14958 13676 15642
rect 13832 15026 13860 15982
rect 13820 15020 13872 15026
rect 13820 14962 13872 14968
rect 13636 14952 13688 14958
rect 13636 14894 13688 14900
rect 13544 14476 13596 14482
rect 13544 14418 13596 14424
rect 13820 14476 13872 14482
rect 13820 14418 13872 14424
rect 13832 14074 13860 14418
rect 13820 14068 13872 14074
rect 13820 14010 13872 14016
rect 13636 13864 13688 13870
rect 13636 13806 13688 13812
rect 13648 13394 13676 13806
rect 13924 13716 13952 17682
rect 14016 17610 14044 22034
rect 14292 21622 14320 25774
rect 14556 25356 14608 25362
rect 14556 25298 14608 25304
rect 14372 25152 14424 25158
rect 14372 25094 14424 25100
rect 14384 24274 14412 25094
rect 14568 24750 14596 25298
rect 14556 24744 14608 24750
rect 14556 24686 14608 24692
rect 14372 24268 14424 24274
rect 14372 24210 14424 24216
rect 14464 24268 14516 24274
rect 14464 24210 14516 24216
rect 14384 23118 14412 24210
rect 14476 24070 14504 24210
rect 14740 24200 14792 24206
rect 14740 24142 14792 24148
rect 14464 24064 14516 24070
rect 14464 24006 14516 24012
rect 14556 24064 14608 24070
rect 14556 24006 14608 24012
rect 14476 23526 14504 24006
rect 14568 23662 14596 24006
rect 14752 23866 14780 24142
rect 14740 23860 14792 23866
rect 14740 23802 14792 23808
rect 14556 23656 14608 23662
rect 14556 23598 14608 23604
rect 14464 23520 14516 23526
rect 14464 23462 14516 23468
rect 14372 23112 14424 23118
rect 14372 23054 14424 23060
rect 14476 22642 14504 23462
rect 14568 23186 14596 23598
rect 14556 23180 14608 23186
rect 14556 23122 14608 23128
rect 14464 22636 14516 22642
rect 14464 22578 14516 22584
rect 14372 22500 14424 22506
rect 14372 22442 14424 22448
rect 14280 21616 14332 21622
rect 14280 21558 14332 21564
rect 14096 18896 14148 18902
rect 14096 18838 14148 18844
rect 14108 18222 14136 18838
rect 14096 18216 14148 18222
rect 14096 18158 14148 18164
rect 14188 18148 14240 18154
rect 14188 18090 14240 18096
rect 14200 17746 14228 18090
rect 14188 17740 14240 17746
rect 14188 17682 14240 17688
rect 14004 17604 14056 17610
rect 14004 17546 14056 17552
rect 14004 16788 14056 16794
rect 14004 16730 14056 16736
rect 13832 13688 13952 13716
rect 13636 13388 13688 13394
rect 13636 13330 13688 13336
rect 13728 13388 13780 13394
rect 13728 13330 13780 13336
rect 13636 13184 13688 13190
rect 13636 13126 13688 13132
rect 13544 11756 13596 11762
rect 13544 11698 13596 11704
rect 13556 11218 13584 11698
rect 13648 11626 13676 13126
rect 13740 12306 13768 13330
rect 13728 12300 13780 12306
rect 13728 12242 13780 12248
rect 13636 11620 13688 11626
rect 13636 11562 13688 11568
rect 13544 11212 13596 11218
rect 13544 11154 13596 11160
rect 13452 11076 13504 11082
rect 13452 11018 13504 11024
rect 13372 10662 13492 10690
rect 13360 10600 13412 10606
rect 13360 10542 13412 10548
rect 13084 10260 13136 10266
rect 13084 10202 13136 10208
rect 13176 10260 13228 10266
rect 13176 10202 13228 10208
rect 13096 9738 13124 10202
rect 13096 9710 13216 9738
rect 13084 8900 13136 8906
rect 13084 8842 13136 8848
rect 13096 8566 13124 8842
rect 13084 8560 13136 8566
rect 13084 8502 13136 8508
rect 12440 7948 12492 7954
rect 12440 7890 12492 7896
rect 12992 7948 13044 7954
rect 12992 7890 13044 7896
rect 12360 7806 12480 7834
rect 12452 6866 12480 7806
rect 12440 6860 12492 6866
rect 12440 6802 12492 6808
rect 13188 6254 13216 9710
rect 13268 9512 13320 9518
rect 13268 9454 13320 9460
rect 13280 9042 13308 9454
rect 13372 9178 13400 10542
rect 13360 9172 13412 9178
rect 13360 9114 13412 9120
rect 13268 9036 13320 9042
rect 13268 8978 13320 8984
rect 13280 8498 13308 8978
rect 13268 8492 13320 8498
rect 13268 8434 13320 8440
rect 13464 8294 13492 10662
rect 13556 10130 13584 11154
rect 13648 10606 13676 11562
rect 13740 11354 13768 12242
rect 13728 11348 13780 11354
rect 13728 11290 13780 11296
rect 13636 10600 13688 10606
rect 13636 10542 13688 10548
rect 13728 10464 13780 10470
rect 13728 10406 13780 10412
rect 13740 10266 13768 10406
rect 13728 10260 13780 10266
rect 13728 10202 13780 10208
rect 13544 10124 13596 10130
rect 13544 10066 13596 10072
rect 13556 9518 13584 10066
rect 13636 9648 13688 9654
rect 13832 9602 13860 13688
rect 14016 12646 14044 16730
rect 14004 12640 14056 12646
rect 14004 12582 14056 12588
rect 13912 11212 13964 11218
rect 13912 11154 13964 11160
rect 13924 10674 13952 11154
rect 13912 10668 13964 10674
rect 13912 10610 13964 10616
rect 13912 10124 13964 10130
rect 13912 10066 13964 10072
rect 13688 9596 13860 9602
rect 13636 9590 13860 9596
rect 13648 9574 13860 9590
rect 13544 9512 13596 9518
rect 13544 9454 13596 9460
rect 13728 9444 13780 9450
rect 13728 9386 13780 9392
rect 13740 9042 13768 9386
rect 13728 9036 13780 9042
rect 13728 8978 13780 8984
rect 13452 8288 13504 8294
rect 13452 8230 13504 8236
rect 13740 7410 13768 8978
rect 13924 8838 13952 10066
rect 13912 8832 13964 8838
rect 13912 8774 13964 8780
rect 13728 7404 13780 7410
rect 13728 7346 13780 7352
rect 13544 6860 13596 6866
rect 13544 6802 13596 6808
rect 13360 6656 13412 6662
rect 13360 6598 13412 6604
rect 13372 6254 13400 6598
rect 13176 6248 13228 6254
rect 13176 6190 13228 6196
rect 13360 6248 13412 6254
rect 13360 6190 13412 6196
rect 13372 5953 13400 6190
rect 13358 5944 13414 5953
rect 12164 5908 12216 5914
rect 13358 5879 13414 5888
rect 12164 5850 12216 5856
rect 13556 5778 13584 6802
rect 13636 6724 13688 6730
rect 13636 6666 13688 6672
rect 12256 5772 12308 5778
rect 12256 5714 12308 5720
rect 13544 5772 13596 5778
rect 13544 5714 13596 5720
rect 12268 5302 12296 5714
rect 13648 5642 13676 6666
rect 13740 5846 13768 7346
rect 14016 7342 14044 12582
rect 14384 11830 14412 22442
rect 14832 22092 14884 22098
rect 14832 22034 14884 22040
rect 14648 21004 14700 21010
rect 14648 20946 14700 20952
rect 14660 19922 14688 20946
rect 14740 20460 14792 20466
rect 14740 20402 14792 20408
rect 14464 19916 14516 19922
rect 14464 19858 14516 19864
rect 14648 19916 14700 19922
rect 14648 19858 14700 19864
rect 14476 18834 14504 19858
rect 14660 19718 14688 19858
rect 14648 19712 14700 19718
rect 14648 19654 14700 19660
rect 14660 18902 14688 19654
rect 14752 18970 14780 20402
rect 14844 19802 14872 22034
rect 14936 20466 14964 35634
rect 15028 34746 15056 36654
rect 15304 36106 15332 37216
rect 15384 37198 15436 37204
rect 15764 36582 15792 37266
rect 15856 36922 15884 37742
rect 16040 37482 16068 40200
rect 17224 37868 17276 37874
rect 17224 37810 17276 37816
rect 16040 37454 16528 37482
rect 17236 37466 17264 37810
rect 17960 37800 18012 37806
rect 17960 37742 18012 37748
rect 17972 37466 18000 37742
rect 16028 37324 16080 37330
rect 16028 37266 16080 37272
rect 15844 36916 15896 36922
rect 15844 36858 15896 36864
rect 15936 36644 15988 36650
rect 15936 36586 15988 36592
rect 15752 36576 15804 36582
rect 15752 36518 15804 36524
rect 15292 36100 15344 36106
rect 15292 36042 15344 36048
rect 15304 35630 15332 36042
rect 15764 35834 15792 36518
rect 15752 35828 15804 35834
rect 15752 35770 15804 35776
rect 15292 35624 15344 35630
rect 15292 35566 15344 35572
rect 15016 34740 15068 34746
rect 15016 34682 15068 34688
rect 15304 34610 15332 35566
rect 15752 35080 15804 35086
rect 15752 35022 15804 35028
rect 15292 34604 15344 34610
rect 15292 34546 15344 34552
rect 15108 34536 15160 34542
rect 15108 34478 15160 34484
rect 15120 34202 15148 34478
rect 15108 34196 15160 34202
rect 15108 34138 15160 34144
rect 15764 33980 15792 35022
rect 15948 34218 15976 36586
rect 16040 35698 16068 37266
rect 16028 35692 16080 35698
rect 16028 35634 16080 35640
rect 15948 34190 16068 34218
rect 15936 33992 15988 33998
rect 15764 33952 15936 33980
rect 15936 33934 15988 33940
rect 15108 33448 15160 33454
rect 15108 33390 15160 33396
rect 15120 33114 15148 33390
rect 15844 33312 15896 33318
rect 15844 33254 15896 33260
rect 15108 33108 15160 33114
rect 15108 33050 15160 33056
rect 15660 32972 15712 32978
rect 15660 32914 15712 32920
rect 15672 32570 15700 32914
rect 15660 32564 15712 32570
rect 15660 32506 15712 32512
rect 15856 32366 15884 33254
rect 15108 32360 15160 32366
rect 15108 32302 15160 32308
rect 15844 32360 15896 32366
rect 15844 32302 15896 32308
rect 15120 31822 15148 32302
rect 15856 31890 15884 32302
rect 15200 31884 15252 31890
rect 15200 31826 15252 31832
rect 15844 31884 15896 31890
rect 15844 31826 15896 31832
rect 15108 31816 15160 31822
rect 15108 31758 15160 31764
rect 15120 31482 15148 31758
rect 15108 31476 15160 31482
rect 15108 31418 15160 31424
rect 15212 30666 15240 31826
rect 15856 31754 15884 31826
rect 15844 31748 15896 31754
rect 15844 31690 15896 31696
rect 15384 31272 15436 31278
rect 15384 31214 15436 31220
rect 15568 31272 15620 31278
rect 15568 31214 15620 31220
rect 15660 31272 15712 31278
rect 15660 31214 15712 31220
rect 15292 31204 15344 31210
rect 15292 31146 15344 31152
rect 15200 30660 15252 30666
rect 15200 30602 15252 30608
rect 15200 29708 15252 29714
rect 15200 29650 15252 29656
rect 15212 29578 15240 29650
rect 15304 29578 15332 31146
rect 15200 29572 15252 29578
rect 15200 29514 15252 29520
rect 15292 29572 15344 29578
rect 15292 29514 15344 29520
rect 15292 28960 15344 28966
rect 15292 28902 15344 28908
rect 15304 28626 15332 28902
rect 15292 28620 15344 28626
rect 15292 28562 15344 28568
rect 15396 28014 15424 31214
rect 15476 30728 15528 30734
rect 15476 30670 15528 30676
rect 15488 29782 15516 30670
rect 15580 30258 15608 31214
rect 15672 30598 15700 31214
rect 15856 30802 15884 31690
rect 15844 30796 15896 30802
rect 15844 30738 15896 30744
rect 15660 30592 15712 30598
rect 15660 30534 15712 30540
rect 15568 30252 15620 30258
rect 15568 30194 15620 30200
rect 15476 29776 15528 29782
rect 15476 29718 15528 29724
rect 15672 29034 15700 30534
rect 15844 30184 15896 30190
rect 15842 30152 15844 30161
rect 15896 30152 15898 30161
rect 15842 30087 15898 30096
rect 15844 29708 15896 29714
rect 15844 29650 15896 29656
rect 15856 29034 15884 29650
rect 15660 29028 15712 29034
rect 15660 28970 15712 28976
rect 15844 29028 15896 29034
rect 15844 28970 15896 28976
rect 15568 28756 15620 28762
rect 15568 28698 15620 28704
rect 15476 28552 15528 28558
rect 15476 28494 15528 28500
rect 15488 28218 15516 28494
rect 15476 28212 15528 28218
rect 15476 28154 15528 28160
rect 15384 28008 15436 28014
rect 15384 27950 15436 27956
rect 15580 27946 15608 28698
rect 15752 28552 15804 28558
rect 15752 28494 15804 28500
rect 15568 27940 15620 27946
rect 15568 27882 15620 27888
rect 15476 26920 15528 26926
rect 15476 26862 15528 26868
rect 15384 26512 15436 26518
rect 15384 26454 15436 26460
rect 15292 26376 15344 26382
rect 15292 26318 15344 26324
rect 15304 25838 15332 26318
rect 15292 25832 15344 25838
rect 15292 25774 15344 25780
rect 15396 25362 15424 26454
rect 15488 26314 15516 26862
rect 15580 26790 15608 27882
rect 15764 27470 15792 28494
rect 15752 27464 15804 27470
rect 15752 27406 15804 27412
rect 15568 26784 15620 26790
rect 15568 26726 15620 26732
rect 15476 26308 15528 26314
rect 15476 26250 15528 26256
rect 15752 25832 15804 25838
rect 15752 25774 15804 25780
rect 15384 25356 15436 25362
rect 15384 25298 15436 25304
rect 15476 25356 15528 25362
rect 15476 25298 15528 25304
rect 15396 24954 15424 25298
rect 15384 24948 15436 24954
rect 15384 24890 15436 24896
rect 15488 24682 15516 25298
rect 15476 24676 15528 24682
rect 15476 24618 15528 24624
rect 15488 24274 15516 24618
rect 15660 24608 15712 24614
rect 15660 24550 15712 24556
rect 15476 24268 15528 24274
rect 15476 24210 15528 24216
rect 15292 23656 15344 23662
rect 15292 23598 15344 23604
rect 15304 23254 15332 23598
rect 15292 23248 15344 23254
rect 15292 23190 15344 23196
rect 15292 22636 15344 22642
rect 15292 22578 15344 22584
rect 15108 22568 15160 22574
rect 15108 22510 15160 22516
rect 15120 20942 15148 22510
rect 15108 20936 15160 20942
rect 15108 20878 15160 20884
rect 15304 20534 15332 22578
rect 15384 21888 15436 21894
rect 15384 21830 15436 21836
rect 15292 20528 15344 20534
rect 15292 20470 15344 20476
rect 14924 20460 14976 20466
rect 14924 20402 14976 20408
rect 15108 20460 15160 20466
rect 15108 20402 15160 20408
rect 15120 19922 15148 20402
rect 15200 20392 15252 20398
rect 15200 20334 15252 20340
rect 15108 19916 15160 19922
rect 15108 19858 15160 19864
rect 14844 19774 15056 19802
rect 14832 19712 14884 19718
rect 14832 19654 14884 19660
rect 14844 19378 14872 19654
rect 14832 19372 14884 19378
rect 14832 19314 14884 19320
rect 14740 18964 14792 18970
rect 14740 18906 14792 18912
rect 14648 18896 14700 18902
rect 14648 18838 14700 18844
rect 14464 18828 14516 18834
rect 14464 18770 14516 18776
rect 14752 17338 14780 18906
rect 14832 18284 14884 18290
rect 14832 18226 14884 18232
rect 14740 17332 14792 17338
rect 14740 17274 14792 17280
rect 14844 16046 14872 18226
rect 14924 18080 14976 18086
rect 14924 18022 14976 18028
rect 14936 17134 14964 18022
rect 14924 17128 14976 17134
rect 14924 17070 14976 17076
rect 14832 16040 14884 16046
rect 14832 15982 14884 15988
rect 14464 15700 14516 15706
rect 14464 15642 14516 15648
rect 14476 15502 14504 15642
rect 14464 15496 14516 15502
rect 14464 15438 14516 15444
rect 14476 14482 14504 15438
rect 14464 14476 14516 14482
rect 14464 14418 14516 14424
rect 14740 13728 14792 13734
rect 14740 13670 14792 13676
rect 14556 13184 14608 13190
rect 14556 13126 14608 13132
rect 14464 12096 14516 12102
rect 14464 12038 14516 12044
rect 14476 11898 14504 12038
rect 14464 11892 14516 11898
rect 14464 11834 14516 11840
rect 14372 11824 14424 11830
rect 14372 11766 14424 11772
rect 14096 11552 14148 11558
rect 14096 11494 14148 11500
rect 14108 11014 14136 11494
rect 14476 11218 14504 11834
rect 14464 11212 14516 11218
rect 14464 11154 14516 11160
rect 14096 11008 14148 11014
rect 14096 10950 14148 10956
rect 13820 7336 13872 7342
rect 13820 7278 13872 7284
rect 14004 7336 14056 7342
rect 14004 7278 14056 7284
rect 13832 5914 13860 7278
rect 14002 6352 14058 6361
rect 14002 6287 14058 6296
rect 14016 6254 14044 6287
rect 14108 6254 14136 10950
rect 14464 10600 14516 10606
rect 14464 10542 14516 10548
rect 14188 10464 14240 10470
rect 14188 10406 14240 10412
rect 14200 10062 14228 10406
rect 14188 10056 14240 10062
rect 14188 9998 14240 10004
rect 14476 9654 14504 10542
rect 14464 9648 14516 9654
rect 14464 9590 14516 9596
rect 14188 8968 14240 8974
rect 14188 8910 14240 8916
rect 14372 8968 14424 8974
rect 14372 8910 14424 8916
rect 14200 8566 14228 8910
rect 14188 8560 14240 8566
rect 14188 8502 14240 8508
rect 14188 7948 14240 7954
rect 14188 7890 14240 7896
rect 14200 7478 14228 7890
rect 14188 7472 14240 7478
rect 14188 7414 14240 7420
rect 14280 7268 14332 7274
rect 14280 7210 14332 7216
rect 14188 6656 14240 6662
rect 14188 6598 14240 6604
rect 14004 6248 14056 6254
rect 14004 6190 14056 6196
rect 14096 6248 14148 6254
rect 14096 6190 14148 6196
rect 13820 5908 13872 5914
rect 13820 5850 13872 5856
rect 13728 5840 13780 5846
rect 13728 5782 13780 5788
rect 13820 5772 13872 5778
rect 13820 5714 13872 5720
rect 13832 5658 13860 5714
rect 13636 5636 13688 5642
rect 13636 5578 13688 5584
rect 13740 5630 13860 5658
rect 12808 5568 12860 5574
rect 12808 5510 12860 5516
rect 13452 5568 13504 5574
rect 13452 5510 13504 5516
rect 13544 5568 13596 5574
rect 13544 5510 13596 5516
rect 12256 5296 12308 5302
rect 12256 5238 12308 5244
rect 12716 5228 12768 5234
rect 12716 5170 12768 5176
rect 11796 4820 11848 4826
rect 11796 4762 11848 4768
rect 12728 4690 12756 5170
rect 12820 5166 12848 5510
rect 13464 5370 13492 5510
rect 13452 5364 13504 5370
rect 13452 5306 13504 5312
rect 12808 5160 12860 5166
rect 12808 5102 12860 5108
rect 13452 5092 13504 5098
rect 13452 5034 13504 5040
rect 12716 4684 12768 4690
rect 12716 4626 12768 4632
rect 13464 4554 13492 5034
rect 13452 4548 13504 4554
rect 13452 4490 13504 4496
rect 12900 4140 12952 4146
rect 12900 4082 12952 4088
rect 11888 4004 11940 4010
rect 11888 3946 11940 3952
rect 11900 3602 11928 3946
rect 12912 3777 12940 4082
rect 13464 4078 13492 4490
rect 13268 4072 13320 4078
rect 13268 4014 13320 4020
rect 13452 4072 13504 4078
rect 13452 4014 13504 4020
rect 12898 3768 12954 3777
rect 12898 3703 12954 3712
rect 13280 3602 13308 4014
rect 11888 3596 11940 3602
rect 11888 3538 11940 3544
rect 13268 3596 13320 3602
rect 13268 3538 13320 3544
rect 13556 3534 13584 5510
rect 13648 5166 13676 5578
rect 13740 5370 13768 5630
rect 13728 5364 13780 5370
rect 13728 5306 13780 5312
rect 14016 5166 14044 6190
rect 14200 6186 14228 6598
rect 14188 6180 14240 6186
rect 14188 6122 14240 6128
rect 13636 5160 13688 5166
rect 13636 5102 13688 5108
rect 14004 5160 14056 5166
rect 14004 5102 14056 5108
rect 13820 4004 13872 4010
rect 13820 3946 13872 3952
rect 13544 3528 13596 3534
rect 13544 3470 13596 3476
rect 11704 3120 11756 3126
rect 11704 3062 11756 3068
rect 13556 3058 13584 3470
rect 13832 3058 13860 3946
rect 14200 3602 14228 6122
rect 14292 5914 14320 7210
rect 14280 5908 14332 5914
rect 14280 5850 14332 5856
rect 14384 4690 14412 8910
rect 14568 5778 14596 13126
rect 14752 12782 14780 13670
rect 15028 13190 15056 19774
rect 15212 19514 15240 20334
rect 15200 19508 15252 19514
rect 15200 19450 15252 19456
rect 15200 19236 15252 19242
rect 15200 19178 15252 19184
rect 15212 18290 15240 19178
rect 15200 18284 15252 18290
rect 15200 18226 15252 18232
rect 15292 18216 15344 18222
rect 15292 18158 15344 18164
rect 15304 17746 15332 18158
rect 15292 17740 15344 17746
rect 15292 17682 15344 17688
rect 15292 17196 15344 17202
rect 15396 17184 15424 21830
rect 15488 21690 15516 24210
rect 15672 23866 15700 24550
rect 15660 23860 15712 23866
rect 15660 23802 15712 23808
rect 15672 23186 15700 23802
rect 15660 23180 15712 23186
rect 15660 23122 15712 23128
rect 15764 22642 15792 25774
rect 15856 23186 15884 28970
rect 15948 24410 15976 33934
rect 16040 26858 16068 34190
rect 16212 33516 16264 33522
rect 16212 33458 16264 33464
rect 16224 32978 16252 33458
rect 16120 32972 16172 32978
rect 16120 32914 16172 32920
rect 16212 32972 16264 32978
rect 16212 32914 16264 32920
rect 16132 31958 16160 32914
rect 16224 32570 16252 32914
rect 16396 32904 16448 32910
rect 16396 32846 16448 32852
rect 16212 32564 16264 32570
rect 16212 32506 16264 32512
rect 16212 32224 16264 32230
rect 16212 32166 16264 32172
rect 16120 31952 16172 31958
rect 16120 31894 16172 31900
rect 16224 31890 16252 32166
rect 16408 31890 16436 32846
rect 16212 31884 16264 31890
rect 16212 31826 16264 31832
rect 16396 31884 16448 31890
rect 16396 31826 16448 31832
rect 16212 30796 16264 30802
rect 16212 30738 16264 30744
rect 16120 30592 16172 30598
rect 16120 30534 16172 30540
rect 16132 29714 16160 30534
rect 16120 29708 16172 29714
rect 16120 29650 16172 29656
rect 16120 29300 16172 29306
rect 16120 29242 16172 29248
rect 16132 29034 16160 29242
rect 16120 29028 16172 29034
rect 16120 28970 16172 28976
rect 16132 28218 16160 28970
rect 16120 28212 16172 28218
rect 16120 28154 16172 28160
rect 16120 27532 16172 27538
rect 16120 27474 16172 27480
rect 16132 26926 16160 27474
rect 16120 26920 16172 26926
rect 16120 26862 16172 26868
rect 16028 26852 16080 26858
rect 16028 26794 16080 26800
rect 16040 26382 16068 26794
rect 16224 26586 16252 30738
rect 16396 30184 16448 30190
rect 16396 30126 16448 30132
rect 16304 29844 16356 29850
rect 16304 29786 16356 29792
rect 16316 29714 16344 29786
rect 16304 29708 16356 29714
rect 16304 29650 16356 29656
rect 16316 29102 16344 29650
rect 16408 29170 16436 30126
rect 16396 29164 16448 29170
rect 16396 29106 16448 29112
rect 16304 29096 16356 29102
rect 16356 29044 16436 29050
rect 16304 29038 16436 29044
rect 16316 29022 16436 29038
rect 16408 28014 16436 29022
rect 16304 28008 16356 28014
rect 16304 27950 16356 27956
rect 16396 28008 16448 28014
rect 16396 27950 16448 27956
rect 16212 26580 16264 26586
rect 16212 26522 16264 26528
rect 16028 26376 16080 26382
rect 16028 26318 16080 26324
rect 16120 25832 16172 25838
rect 16120 25774 16172 25780
rect 16132 25498 16160 25774
rect 16120 25492 16172 25498
rect 16120 25434 16172 25440
rect 16212 24880 16264 24886
rect 16212 24822 16264 24828
rect 15936 24404 15988 24410
rect 15936 24346 15988 24352
rect 15844 23180 15896 23186
rect 15844 23122 15896 23128
rect 15752 22636 15804 22642
rect 15752 22578 15804 22584
rect 15752 22228 15804 22234
rect 15752 22170 15804 22176
rect 15764 22098 15792 22170
rect 15752 22092 15804 22098
rect 15752 22034 15804 22040
rect 15476 21684 15528 21690
rect 15476 21626 15528 21632
rect 15568 21480 15620 21486
rect 15568 21422 15620 21428
rect 15580 18970 15608 21422
rect 15764 21078 15792 22034
rect 15844 21412 15896 21418
rect 15844 21354 15896 21360
rect 15752 21072 15804 21078
rect 15752 21014 15804 21020
rect 15568 18964 15620 18970
rect 15568 18906 15620 18912
rect 15568 17672 15620 17678
rect 15568 17614 15620 17620
rect 15344 17156 15424 17184
rect 15292 17138 15344 17144
rect 15200 17128 15252 17134
rect 15200 17070 15252 17076
rect 15108 14816 15160 14822
rect 15108 14758 15160 14764
rect 15016 13184 15068 13190
rect 15016 13126 15068 13132
rect 15120 12782 15148 14758
rect 15212 14385 15240 17070
rect 15292 16584 15344 16590
rect 15292 16526 15344 16532
rect 15304 15366 15332 16526
rect 15396 16028 15424 17156
rect 15476 17060 15528 17066
rect 15476 17002 15528 17008
rect 15488 16658 15516 17002
rect 15476 16652 15528 16658
rect 15476 16594 15528 16600
rect 15580 16454 15608 17614
rect 15856 17270 15884 21354
rect 15948 18834 15976 24346
rect 16224 24342 16252 24822
rect 16212 24336 16264 24342
rect 16212 24278 16264 24284
rect 16028 24268 16080 24274
rect 16028 24210 16080 24216
rect 16040 22982 16068 24210
rect 16120 23656 16172 23662
rect 16120 23598 16172 23604
rect 16132 23322 16160 23598
rect 16120 23316 16172 23322
rect 16120 23258 16172 23264
rect 16316 23168 16344 27950
rect 16396 27464 16448 27470
rect 16396 27406 16448 27412
rect 16408 27130 16436 27406
rect 16396 27124 16448 27130
rect 16396 27066 16448 27072
rect 16396 26308 16448 26314
rect 16396 26250 16448 26256
rect 16408 24750 16436 26250
rect 16396 24744 16448 24750
rect 16396 24686 16448 24692
rect 16132 23140 16344 23168
rect 16396 23180 16448 23186
rect 16028 22976 16080 22982
rect 16028 22918 16080 22924
rect 16132 22386 16160 23140
rect 16396 23122 16448 23128
rect 16304 22976 16356 22982
rect 16304 22918 16356 22924
rect 16040 22358 16160 22386
rect 16040 19786 16068 22358
rect 16212 22092 16264 22098
rect 16212 22034 16264 22040
rect 16224 20806 16252 22034
rect 16212 20800 16264 20806
rect 16212 20742 16264 20748
rect 16316 20398 16344 22918
rect 16408 22166 16436 23122
rect 16396 22160 16448 22166
rect 16396 22102 16448 22108
rect 16396 22024 16448 22030
rect 16396 21966 16448 21972
rect 16408 20602 16436 21966
rect 16396 20596 16448 20602
rect 16396 20538 16448 20544
rect 16304 20392 16356 20398
rect 16304 20334 16356 20340
rect 16120 20256 16172 20262
rect 16120 20198 16172 20204
rect 16212 20256 16264 20262
rect 16212 20198 16264 20204
rect 16028 19780 16080 19786
rect 16028 19722 16080 19728
rect 15936 18828 15988 18834
rect 15936 18770 15988 18776
rect 15948 18222 15976 18770
rect 15936 18216 15988 18222
rect 15936 18158 15988 18164
rect 15844 17264 15896 17270
rect 15844 17206 15896 17212
rect 15568 16448 15620 16454
rect 15568 16390 15620 16396
rect 15476 16040 15528 16046
rect 15396 16000 15476 16028
rect 15292 15360 15344 15366
rect 15292 15302 15344 15308
rect 15292 15020 15344 15026
rect 15292 14962 15344 14968
rect 15198 14376 15254 14385
rect 15198 14311 15254 14320
rect 15200 14272 15252 14278
rect 15200 14214 15252 14220
rect 15212 12850 15240 14214
rect 15304 13870 15332 14962
rect 15396 14958 15424 16000
rect 15476 15982 15528 15988
rect 15936 15904 15988 15910
rect 15936 15846 15988 15852
rect 15660 15088 15712 15094
rect 15660 15030 15712 15036
rect 15384 14952 15436 14958
rect 15384 14894 15436 14900
rect 15568 14952 15620 14958
rect 15568 14894 15620 14900
rect 15396 14822 15424 14894
rect 15384 14816 15436 14822
rect 15384 14758 15436 14764
rect 15580 14498 15608 14894
rect 15672 14618 15700 15030
rect 15660 14612 15712 14618
rect 15660 14554 15712 14560
rect 15844 14612 15896 14618
rect 15844 14554 15896 14560
rect 15856 14498 15884 14554
rect 15580 14470 15884 14498
rect 15580 13938 15608 14470
rect 15568 13932 15620 13938
rect 15568 13874 15620 13880
rect 15292 13864 15344 13870
rect 15292 13806 15344 13812
rect 15844 13524 15896 13530
rect 15844 13466 15896 13472
rect 15292 13388 15344 13394
rect 15292 13330 15344 13336
rect 15200 12844 15252 12850
rect 15200 12786 15252 12792
rect 14740 12776 14792 12782
rect 14740 12718 14792 12724
rect 15108 12776 15160 12782
rect 15108 12718 15160 12724
rect 15120 12374 15148 12718
rect 15108 12368 15160 12374
rect 15108 12310 15160 12316
rect 15212 12306 15240 12786
rect 15200 12300 15252 12306
rect 15200 12242 15252 12248
rect 14648 12096 14700 12102
rect 14648 12038 14700 12044
rect 14660 11218 14688 12038
rect 15106 11792 15162 11801
rect 15106 11727 15162 11736
rect 15120 11694 15148 11727
rect 15108 11688 15160 11694
rect 15108 11630 15160 11636
rect 14648 11212 14700 11218
rect 14648 11154 14700 11160
rect 15212 5778 15240 12242
rect 15304 11218 15332 13330
rect 15476 13252 15528 13258
rect 15476 13194 15528 13200
rect 15488 12617 15516 13194
rect 15856 12986 15884 13466
rect 15948 13394 15976 15846
rect 16040 15162 16068 19722
rect 16132 19718 16160 20198
rect 16224 20058 16252 20198
rect 16212 20052 16264 20058
rect 16212 19994 16264 20000
rect 16120 19712 16172 19718
rect 16120 19654 16172 19660
rect 16500 19310 16528 37454
rect 17224 37460 17276 37466
rect 17224 37402 17276 37408
rect 17960 37460 18012 37466
rect 17960 37402 18012 37408
rect 17500 37324 17552 37330
rect 17500 37266 17552 37272
rect 16672 36168 16724 36174
rect 16672 36110 16724 36116
rect 16684 35834 16712 36110
rect 16672 35828 16724 35834
rect 16672 35770 16724 35776
rect 17040 34944 17092 34950
rect 17040 34886 17092 34892
rect 17052 34542 17080 34886
rect 17224 34740 17276 34746
rect 17224 34682 17276 34688
rect 17040 34536 17092 34542
rect 17040 34478 17092 34484
rect 17236 34066 17264 34682
rect 17224 34060 17276 34066
rect 17224 34002 17276 34008
rect 16580 33448 16632 33454
rect 16580 33390 16632 33396
rect 16592 33046 16620 33390
rect 17132 33312 17184 33318
rect 17132 33254 17184 33260
rect 16672 33108 16724 33114
rect 16672 33050 16724 33056
rect 16580 33040 16632 33046
rect 16580 32982 16632 32988
rect 16684 32434 16712 33050
rect 17144 32978 17172 33254
rect 17512 33130 17540 37266
rect 17972 36786 18000 37402
rect 17960 36780 18012 36786
rect 17960 36722 18012 36728
rect 17972 36242 18000 36722
rect 18144 36712 18196 36718
rect 18144 36654 18196 36660
rect 17960 36236 18012 36242
rect 17960 36178 18012 36184
rect 18156 36038 18184 36654
rect 18248 36038 18276 40200
rect 19580 38652 19876 38672
rect 19636 38650 19660 38652
rect 19716 38650 19740 38652
rect 19796 38650 19820 38652
rect 19658 38598 19660 38650
rect 19722 38598 19734 38650
rect 19796 38598 19798 38650
rect 19636 38596 19660 38598
rect 19716 38596 19740 38598
rect 19796 38596 19820 38598
rect 19580 38576 19876 38596
rect 19168 38554 19288 38570
rect 19168 38548 19300 38554
rect 19168 38542 19248 38548
rect 19168 38457 19196 38542
rect 19248 38490 19300 38496
rect 19154 38448 19210 38457
rect 19154 38383 19210 38392
rect 18788 37664 18840 37670
rect 18788 37606 18840 37612
rect 18696 36236 18748 36242
rect 18696 36178 18748 36184
rect 18144 36032 18196 36038
rect 18144 35974 18196 35980
rect 18236 36032 18288 36038
rect 18236 35974 18288 35980
rect 18052 35828 18104 35834
rect 18052 35770 18104 35776
rect 18064 35154 18092 35770
rect 18052 35148 18104 35154
rect 18052 35090 18104 35096
rect 17960 33312 18012 33318
rect 17960 33254 18012 33260
rect 17420 33102 17540 33130
rect 17132 32972 17184 32978
rect 17132 32914 17184 32920
rect 16672 32428 16724 32434
rect 16672 32370 16724 32376
rect 16684 29306 16712 32370
rect 17224 31816 17276 31822
rect 17224 31758 17276 31764
rect 17132 30796 17184 30802
rect 17132 30738 17184 30744
rect 16764 30184 16816 30190
rect 16764 30126 16816 30132
rect 16776 29782 16804 30126
rect 16764 29776 16816 29782
rect 16764 29718 16816 29724
rect 16672 29300 16724 29306
rect 16672 29242 16724 29248
rect 16776 28422 16804 29718
rect 16580 28416 16632 28422
rect 16580 28358 16632 28364
rect 16764 28416 16816 28422
rect 16764 28358 16816 28364
rect 16592 28218 16620 28358
rect 16580 28212 16632 28218
rect 16580 28154 16632 28160
rect 16672 28144 16724 28150
rect 16672 28086 16724 28092
rect 16684 26926 16712 28086
rect 16672 26920 16724 26926
rect 16672 26862 16724 26868
rect 16776 24818 16804 28358
rect 17040 28008 17092 28014
rect 17040 27950 17092 27956
rect 17052 26790 17080 27950
rect 17040 26784 17092 26790
rect 17040 26726 17092 26732
rect 16948 26444 17000 26450
rect 16948 26386 17000 26392
rect 16960 25838 16988 26386
rect 16948 25832 17000 25838
rect 16948 25774 17000 25780
rect 16764 24812 16816 24818
rect 16764 24754 16816 24760
rect 16672 24744 16724 24750
rect 16672 24686 16724 24692
rect 16684 24138 16712 24686
rect 17144 24342 17172 30738
rect 17236 30258 17264 31758
rect 17316 31204 17368 31210
rect 17316 31146 17368 31152
rect 17328 30802 17356 31146
rect 17316 30796 17368 30802
rect 17316 30738 17368 30744
rect 17224 30252 17276 30258
rect 17224 30194 17276 30200
rect 17316 29572 17368 29578
rect 17316 29514 17368 29520
rect 17328 29102 17356 29514
rect 17316 29096 17368 29102
rect 17316 29038 17368 29044
rect 17224 28008 17276 28014
rect 17224 27950 17276 27956
rect 17236 27538 17264 27950
rect 17224 27532 17276 27538
rect 17224 27474 17276 27480
rect 17132 24336 17184 24342
rect 17132 24278 17184 24284
rect 17224 24268 17276 24274
rect 17224 24210 17276 24216
rect 16672 24132 16724 24138
rect 16672 24074 16724 24080
rect 16580 23588 16632 23594
rect 16580 23530 16632 23536
rect 16592 21622 16620 23530
rect 16684 23254 16712 24074
rect 16672 23248 16724 23254
rect 16672 23190 16724 23196
rect 17236 22642 17264 24210
rect 17316 24064 17368 24070
rect 17316 24006 17368 24012
rect 17328 23866 17356 24006
rect 17316 23860 17368 23866
rect 17316 23802 17368 23808
rect 17420 23746 17448 33102
rect 17868 32768 17920 32774
rect 17868 32710 17920 32716
rect 17500 32360 17552 32366
rect 17500 32302 17552 32308
rect 17512 31822 17540 32302
rect 17776 32292 17828 32298
rect 17776 32234 17828 32240
rect 17500 31816 17552 31822
rect 17500 31758 17552 31764
rect 17512 30870 17540 31758
rect 17788 31278 17816 32234
rect 17880 31890 17908 32710
rect 17972 32366 18000 33254
rect 17960 32360 18012 32366
rect 17960 32302 18012 32308
rect 17868 31884 17920 31890
rect 17868 31826 17920 31832
rect 17776 31272 17828 31278
rect 17776 31214 17828 31220
rect 17788 30938 17816 31214
rect 18052 31136 18104 31142
rect 18052 31078 18104 31084
rect 17776 30932 17828 30938
rect 17776 30874 17828 30880
rect 17500 30864 17552 30870
rect 17500 30806 17552 30812
rect 17960 30796 18012 30802
rect 17960 30738 18012 30744
rect 17972 30326 18000 30738
rect 18064 30326 18092 31078
rect 17960 30320 18012 30326
rect 17960 30262 18012 30268
rect 18052 30320 18104 30326
rect 18052 30262 18104 30268
rect 17868 30184 17920 30190
rect 18156 30138 18184 35974
rect 18708 35834 18736 36178
rect 18696 35828 18748 35834
rect 18696 35770 18748 35776
rect 18420 33856 18472 33862
rect 18420 33798 18472 33804
rect 18328 32904 18380 32910
rect 18328 32846 18380 32852
rect 18340 32570 18368 32846
rect 18328 32564 18380 32570
rect 18328 32506 18380 32512
rect 18340 32450 18368 32506
rect 18248 32422 18368 32450
rect 18248 30734 18276 32422
rect 18328 31816 18380 31822
rect 18328 31758 18380 31764
rect 18340 31346 18368 31758
rect 18328 31340 18380 31346
rect 18328 31282 18380 31288
rect 18340 31142 18368 31282
rect 18328 31136 18380 31142
rect 18328 31078 18380 31084
rect 18236 30728 18288 30734
rect 18236 30670 18288 30676
rect 17868 30126 17920 30132
rect 17880 29866 17908 30126
rect 17972 30110 18184 30138
rect 17972 30054 18000 30110
rect 17960 30048 18012 30054
rect 17960 29990 18012 29996
rect 18248 29866 18276 30670
rect 18328 30184 18380 30190
rect 18328 30126 18380 30132
rect 17880 29838 18276 29866
rect 17972 28558 18000 29838
rect 18340 29306 18368 30126
rect 18328 29300 18380 29306
rect 18328 29242 18380 29248
rect 18052 28620 18104 28626
rect 18052 28562 18104 28568
rect 17960 28552 18012 28558
rect 17960 28494 18012 28500
rect 17500 26784 17552 26790
rect 17500 26726 17552 26732
rect 17512 26382 17540 26726
rect 17684 26444 17736 26450
rect 17684 26386 17736 26392
rect 17500 26376 17552 26382
rect 17500 26318 17552 26324
rect 17512 24750 17540 26318
rect 17696 25838 17724 26386
rect 18064 26382 18092 28562
rect 18236 28552 18288 28558
rect 18236 28494 18288 28500
rect 18248 28150 18276 28494
rect 18236 28144 18288 28150
rect 18236 28086 18288 28092
rect 18144 27600 18196 27606
rect 18144 27542 18196 27548
rect 18156 27062 18184 27542
rect 18144 27056 18196 27062
rect 18144 26998 18196 27004
rect 18052 26376 18104 26382
rect 18052 26318 18104 26324
rect 17684 25832 17736 25838
rect 17684 25774 17736 25780
rect 17500 24744 17552 24750
rect 17500 24686 17552 24692
rect 17696 24070 17724 25774
rect 18052 25764 18104 25770
rect 18052 25706 18104 25712
rect 18064 24818 18092 25706
rect 18248 25362 18276 28086
rect 18328 27668 18380 27674
rect 18328 27610 18380 27616
rect 18340 26450 18368 27610
rect 18328 26444 18380 26450
rect 18328 26386 18380 26392
rect 18328 26308 18380 26314
rect 18328 26250 18380 26256
rect 18236 25356 18288 25362
rect 18236 25298 18288 25304
rect 18340 25242 18368 26250
rect 18248 25214 18368 25242
rect 18052 24812 18104 24818
rect 18052 24754 18104 24760
rect 18248 24682 18276 25214
rect 18144 24676 18196 24682
rect 18144 24618 18196 24624
rect 18236 24676 18288 24682
rect 18236 24618 18288 24624
rect 18156 24138 18184 24618
rect 18236 24268 18288 24274
rect 18236 24210 18288 24216
rect 18052 24132 18104 24138
rect 18052 24074 18104 24080
rect 18144 24132 18196 24138
rect 18144 24074 18196 24080
rect 17684 24064 17736 24070
rect 17684 24006 17736 24012
rect 17328 23718 17448 23746
rect 17224 22636 17276 22642
rect 17224 22578 17276 22584
rect 16764 22568 16816 22574
rect 16764 22510 16816 22516
rect 16856 22568 16908 22574
rect 16856 22510 16908 22516
rect 16580 21616 16632 21622
rect 16580 21558 16632 21564
rect 16776 21570 16804 22510
rect 16868 22234 16896 22510
rect 16856 22228 16908 22234
rect 16856 22170 16908 22176
rect 16776 21542 16896 21570
rect 16580 21480 16632 21486
rect 16580 21422 16632 21428
rect 16764 21480 16816 21486
rect 16764 21422 16816 21428
rect 16212 19304 16264 19310
rect 16212 19246 16264 19252
rect 16488 19304 16540 19310
rect 16488 19246 16540 19252
rect 16224 18970 16252 19246
rect 16212 18964 16264 18970
rect 16212 18906 16264 18912
rect 16120 18080 16172 18086
rect 16120 18022 16172 18028
rect 16304 18080 16356 18086
rect 16304 18022 16356 18028
rect 16132 17338 16160 18022
rect 16120 17332 16172 17338
rect 16120 17274 16172 17280
rect 16316 16658 16344 18022
rect 16304 16652 16356 16658
rect 16304 16594 16356 16600
rect 16396 15564 16448 15570
rect 16396 15506 16448 15512
rect 16488 15564 16540 15570
rect 16488 15506 16540 15512
rect 16028 15156 16080 15162
rect 16028 15098 16080 15104
rect 16408 15026 16436 15506
rect 16396 15020 16448 15026
rect 16396 14962 16448 14968
rect 16500 14482 16528 15506
rect 16488 14476 16540 14482
rect 16488 14418 16540 14424
rect 16592 14090 16620 21422
rect 16776 21146 16804 21422
rect 16764 21140 16816 21146
rect 16764 21082 16816 21088
rect 16764 21004 16816 21010
rect 16764 20946 16816 20952
rect 16672 20392 16724 20398
rect 16672 20334 16724 20340
rect 16684 19514 16712 20334
rect 16672 19508 16724 19514
rect 16672 19450 16724 19456
rect 16672 19304 16724 19310
rect 16670 19272 16672 19281
rect 16724 19272 16726 19281
rect 16670 19207 16726 19216
rect 16776 18737 16804 20946
rect 16762 18728 16818 18737
rect 16762 18663 16818 18672
rect 16672 17536 16724 17542
rect 16672 17478 16724 17484
rect 16684 17134 16712 17478
rect 16672 17128 16724 17134
rect 16672 17070 16724 17076
rect 16672 15904 16724 15910
rect 16672 15846 16724 15852
rect 16684 15502 16712 15846
rect 16672 15496 16724 15502
rect 16672 15438 16724 15444
rect 16500 14062 16620 14090
rect 16500 14006 16528 14062
rect 16488 14000 16540 14006
rect 16684 13954 16712 15438
rect 16488 13942 16540 13948
rect 16592 13926 16712 13954
rect 15936 13388 15988 13394
rect 15936 13330 15988 13336
rect 15844 12980 15896 12986
rect 15844 12922 15896 12928
rect 15474 12608 15530 12617
rect 15474 12543 15530 12552
rect 15568 11892 15620 11898
rect 15568 11834 15620 11840
rect 15292 11212 15344 11218
rect 15344 11172 15424 11200
rect 15292 11154 15344 11160
rect 15396 10606 15424 11172
rect 15580 11082 15608 11834
rect 15568 11076 15620 11082
rect 15568 11018 15620 11024
rect 15292 10600 15344 10606
rect 15292 10542 15344 10548
rect 15384 10600 15436 10606
rect 15384 10542 15436 10548
rect 15304 10198 15332 10542
rect 15476 10464 15528 10470
rect 15476 10406 15528 10412
rect 15292 10192 15344 10198
rect 15292 10134 15344 10140
rect 15488 9178 15516 10406
rect 15752 10056 15804 10062
rect 15752 9998 15804 10004
rect 15568 9512 15620 9518
rect 15568 9454 15620 9460
rect 15660 9512 15712 9518
rect 15660 9454 15712 9460
rect 15476 9172 15528 9178
rect 15476 9114 15528 9120
rect 15384 8356 15436 8362
rect 15384 8298 15436 8304
rect 15396 7886 15424 8298
rect 15488 7954 15516 9114
rect 15580 8022 15608 9454
rect 15672 8906 15700 9454
rect 15764 9382 15792 9998
rect 15752 9376 15804 9382
rect 15752 9318 15804 9324
rect 15752 9036 15804 9042
rect 15752 8978 15804 8984
rect 15660 8900 15712 8906
rect 15660 8842 15712 8848
rect 15568 8016 15620 8022
rect 15568 7958 15620 7964
rect 15476 7948 15528 7954
rect 15476 7890 15528 7896
rect 15292 7880 15344 7886
rect 15292 7822 15344 7828
rect 15384 7880 15436 7886
rect 15384 7822 15436 7828
rect 15304 6934 15332 7822
rect 15292 6928 15344 6934
rect 15292 6870 15344 6876
rect 15488 6254 15516 7890
rect 15660 6928 15712 6934
rect 15660 6870 15712 6876
rect 15476 6248 15528 6254
rect 15476 6190 15528 6196
rect 14556 5772 14608 5778
rect 14556 5714 14608 5720
rect 15200 5772 15252 5778
rect 15200 5714 15252 5720
rect 14740 5636 14792 5642
rect 14740 5578 14792 5584
rect 14372 4684 14424 4690
rect 14372 4626 14424 4632
rect 14752 4146 14780 5578
rect 15212 5166 15240 5714
rect 15672 5166 15700 6870
rect 15764 6322 15792 8978
rect 15856 8974 15884 12922
rect 16212 12912 16264 12918
rect 16212 12854 16264 12860
rect 16224 12782 16252 12854
rect 16212 12776 16264 12782
rect 16212 12718 16264 12724
rect 16224 11694 16252 12718
rect 16592 11694 16620 13926
rect 16672 13864 16724 13870
rect 16672 13806 16724 13812
rect 16684 12170 16712 13806
rect 16764 13796 16816 13802
rect 16764 13738 16816 13744
rect 16776 13394 16804 13738
rect 16868 13530 16896 21542
rect 17132 21344 17184 21350
rect 17132 21286 17184 21292
rect 16948 21072 17000 21078
rect 16948 21014 17000 21020
rect 16960 19922 16988 21014
rect 16948 19916 17000 19922
rect 16948 19858 17000 19864
rect 17040 16584 17092 16590
rect 17040 16526 17092 16532
rect 16948 15360 17000 15366
rect 16948 15302 17000 15308
rect 16856 13524 16908 13530
rect 16856 13466 16908 13472
rect 16764 13388 16816 13394
rect 16764 13330 16816 13336
rect 16764 12708 16816 12714
rect 16764 12650 16816 12656
rect 16776 12374 16804 12650
rect 16764 12368 16816 12374
rect 16764 12310 16816 12316
rect 16672 12164 16724 12170
rect 16672 12106 16724 12112
rect 16212 11688 16264 11694
rect 16212 11630 16264 11636
rect 16580 11688 16632 11694
rect 16580 11630 16632 11636
rect 16488 11620 16540 11626
rect 16488 11562 16540 11568
rect 16500 11150 16528 11562
rect 16120 11144 16172 11150
rect 16120 11086 16172 11092
rect 16488 11144 16540 11150
rect 16488 11086 16540 11092
rect 16592 11098 16620 11630
rect 16132 10742 16160 11086
rect 16212 11076 16264 11082
rect 16592 11070 16712 11098
rect 16212 11018 16264 11024
rect 16120 10736 16172 10742
rect 16120 10678 16172 10684
rect 16028 9376 16080 9382
rect 16028 9318 16080 9324
rect 15844 8968 15896 8974
rect 15844 8910 15896 8916
rect 16040 8498 16068 9318
rect 16224 8974 16252 11018
rect 16580 11008 16632 11014
rect 16580 10950 16632 10956
rect 16592 10606 16620 10950
rect 16580 10600 16632 10606
rect 16580 10542 16632 10548
rect 16396 10464 16448 10470
rect 16396 10406 16448 10412
rect 16408 10062 16436 10406
rect 16592 10130 16620 10542
rect 16580 10124 16632 10130
rect 16580 10066 16632 10072
rect 16396 10056 16448 10062
rect 16396 9998 16448 10004
rect 16304 9036 16356 9042
rect 16304 8978 16356 8984
rect 16212 8968 16264 8974
rect 16212 8910 16264 8916
rect 16224 8566 16252 8910
rect 16212 8560 16264 8566
rect 16212 8502 16264 8508
rect 16028 8492 16080 8498
rect 16028 8434 16080 8440
rect 16120 8424 16172 8430
rect 16120 8366 16172 8372
rect 16132 8022 16160 8366
rect 16120 8016 16172 8022
rect 16120 7958 16172 7964
rect 15936 7948 15988 7954
rect 15936 7890 15988 7896
rect 15948 7546 15976 7890
rect 15936 7540 15988 7546
rect 15936 7482 15988 7488
rect 15844 6724 15896 6730
rect 15844 6666 15896 6672
rect 15856 6361 15884 6666
rect 16120 6384 16172 6390
rect 15842 6352 15898 6361
rect 15752 6316 15804 6322
rect 16120 6326 16172 6332
rect 15842 6287 15898 6296
rect 15752 6258 15804 6264
rect 16026 5944 16082 5953
rect 16132 5914 16160 6326
rect 16026 5879 16082 5888
rect 16120 5908 16172 5914
rect 16040 5778 16068 5879
rect 16120 5850 16172 5856
rect 15936 5772 15988 5778
rect 15936 5714 15988 5720
rect 16028 5772 16080 5778
rect 16028 5714 16080 5720
rect 15948 5574 15976 5714
rect 15936 5568 15988 5574
rect 15936 5510 15988 5516
rect 16040 5166 16068 5714
rect 16316 5234 16344 8978
rect 16408 8498 16436 9998
rect 16684 9518 16712 11070
rect 16672 9512 16724 9518
rect 16592 9472 16672 9500
rect 16396 8492 16448 8498
rect 16396 8434 16448 8440
rect 16488 7880 16540 7886
rect 16488 7822 16540 7828
rect 16500 7546 16528 7822
rect 16488 7540 16540 7546
rect 16488 7482 16540 7488
rect 16592 6866 16620 9472
rect 16672 9454 16724 9460
rect 16672 8084 16724 8090
rect 16672 8026 16724 8032
rect 16684 7206 16712 8026
rect 16776 7426 16804 12310
rect 16960 12306 16988 15302
rect 17052 13977 17080 16526
rect 17144 15065 17172 21286
rect 17224 17128 17276 17134
rect 17224 17070 17276 17076
rect 17236 15094 17264 17070
rect 17224 15088 17276 15094
rect 17130 15056 17186 15065
rect 17224 15030 17276 15036
rect 17130 14991 17186 15000
rect 17038 13968 17094 13977
rect 17038 13903 17094 13912
rect 17132 13388 17184 13394
rect 17132 13330 17184 13336
rect 17144 13297 17172 13330
rect 17130 13288 17186 13297
rect 17130 13223 17186 13232
rect 17328 12850 17356 23718
rect 17500 23588 17552 23594
rect 17500 23530 17552 23536
rect 17512 20466 17540 23530
rect 17592 23044 17644 23050
rect 17592 22986 17644 22992
rect 17604 21554 17632 22986
rect 17592 21548 17644 21554
rect 17592 21490 17644 21496
rect 17500 20460 17552 20466
rect 17500 20402 17552 20408
rect 17408 20392 17460 20398
rect 17408 20334 17460 20340
rect 17420 20058 17448 20334
rect 17590 20224 17646 20233
rect 17590 20159 17646 20168
rect 17408 20052 17460 20058
rect 17408 19994 17460 20000
rect 17500 20052 17552 20058
rect 17500 19994 17552 20000
rect 17512 19922 17540 19994
rect 17604 19922 17632 20159
rect 17500 19916 17552 19922
rect 17500 19858 17552 19864
rect 17592 19916 17644 19922
rect 17592 19858 17644 19864
rect 17590 19272 17646 19281
rect 17590 19207 17646 19216
rect 17408 18080 17460 18086
rect 17408 18022 17460 18028
rect 17420 17610 17448 18022
rect 17604 17746 17632 19207
rect 17592 17740 17644 17746
rect 17592 17682 17644 17688
rect 17408 17604 17460 17610
rect 17408 17546 17460 17552
rect 17420 17066 17448 17546
rect 17408 17060 17460 17066
rect 17408 17002 17460 17008
rect 17500 16992 17552 16998
rect 17500 16934 17552 16940
rect 17512 16658 17540 16934
rect 17696 16810 17724 24006
rect 18064 23662 18092 24074
rect 18248 23798 18276 24210
rect 18236 23792 18288 23798
rect 18236 23734 18288 23740
rect 18052 23656 18104 23662
rect 18052 23598 18104 23604
rect 18248 23526 18276 23734
rect 18236 23520 18288 23526
rect 18236 23462 18288 23468
rect 18328 23112 18380 23118
rect 18328 23054 18380 23060
rect 18340 22642 18368 23054
rect 18328 22636 18380 22642
rect 18328 22578 18380 22584
rect 17960 22500 18012 22506
rect 17960 22442 18012 22448
rect 17972 22098 18000 22442
rect 17960 22092 18012 22098
rect 17960 22034 18012 22040
rect 17868 22024 17920 22030
rect 17868 21966 17920 21972
rect 17880 21010 17908 21966
rect 17868 21004 17920 21010
rect 17868 20946 17920 20952
rect 17972 20942 18000 22034
rect 18052 21480 18104 21486
rect 18052 21422 18104 21428
rect 18064 21146 18092 21422
rect 18052 21140 18104 21146
rect 18052 21082 18104 21088
rect 17960 20936 18012 20942
rect 17960 20878 18012 20884
rect 17776 20392 17828 20398
rect 17776 20334 17828 20340
rect 17788 19854 17816 20334
rect 17776 19848 17828 19854
rect 17776 19790 17828 19796
rect 17972 18850 18000 20878
rect 18236 20528 18288 20534
rect 18236 20470 18288 20476
rect 18052 19508 18104 19514
rect 18052 19450 18104 19456
rect 17880 18822 18000 18850
rect 17880 18630 17908 18822
rect 17960 18760 18012 18766
rect 17960 18702 18012 18708
rect 17868 18624 17920 18630
rect 17868 18566 17920 18572
rect 17880 18426 17908 18566
rect 17868 18420 17920 18426
rect 17868 18362 17920 18368
rect 17972 17814 18000 18702
rect 18064 18698 18092 19450
rect 18144 19304 18196 19310
rect 18144 19246 18196 19252
rect 18052 18692 18104 18698
rect 18052 18634 18104 18640
rect 18156 18222 18184 19246
rect 18144 18216 18196 18222
rect 18144 18158 18196 18164
rect 17960 17808 18012 17814
rect 17960 17750 18012 17756
rect 17776 17740 17828 17746
rect 17776 17682 17828 17688
rect 17604 16782 17724 16810
rect 17500 16652 17552 16658
rect 17500 16594 17552 16600
rect 17316 12844 17368 12850
rect 17316 12786 17368 12792
rect 16948 12300 17000 12306
rect 16948 12242 17000 12248
rect 17132 11688 17184 11694
rect 17132 11630 17184 11636
rect 16948 11212 17000 11218
rect 16948 11154 17000 11160
rect 16960 8974 16988 11154
rect 17144 10674 17172 11630
rect 17132 10668 17184 10674
rect 17132 10610 17184 10616
rect 17224 10600 17276 10606
rect 17224 10542 17276 10548
rect 17236 10130 17264 10542
rect 17224 10124 17276 10130
rect 17224 10066 17276 10072
rect 17236 10010 17264 10066
rect 17144 9982 17264 10010
rect 16948 8968 17000 8974
rect 16948 8910 17000 8916
rect 16960 8090 16988 8910
rect 17144 8616 17172 9982
rect 17224 9920 17276 9926
rect 17224 9862 17276 9868
rect 17236 9518 17264 9862
rect 17408 9648 17460 9654
rect 17408 9590 17460 9596
rect 17316 9580 17368 9586
rect 17316 9522 17368 9528
rect 17224 9512 17276 9518
rect 17224 9454 17276 9460
rect 17328 9042 17356 9522
rect 17316 9036 17368 9042
rect 17316 8978 17368 8984
rect 17144 8588 17264 8616
rect 17132 8424 17184 8430
rect 17132 8366 17184 8372
rect 16948 8084 17000 8090
rect 16948 8026 17000 8032
rect 17040 7744 17092 7750
rect 17040 7686 17092 7692
rect 16776 7398 16988 7426
rect 16856 7336 16908 7342
rect 16856 7278 16908 7284
rect 16672 7200 16724 7206
rect 16672 7142 16724 7148
rect 16868 6934 16896 7278
rect 16856 6928 16908 6934
rect 16856 6870 16908 6876
rect 16580 6860 16632 6866
rect 16580 6802 16632 6808
rect 16592 6338 16620 6802
rect 16764 6792 16816 6798
rect 16762 6760 16764 6769
rect 16816 6760 16818 6769
rect 16762 6695 16818 6704
rect 16396 6316 16448 6322
rect 16592 6310 16712 6338
rect 16396 6258 16448 6264
rect 16408 5302 16436 6258
rect 16684 6254 16712 6310
rect 16580 6248 16632 6254
rect 16580 6190 16632 6196
rect 16672 6248 16724 6254
rect 16672 6190 16724 6196
rect 16592 5778 16620 6190
rect 16580 5772 16632 5778
rect 16580 5714 16632 5720
rect 16396 5296 16448 5302
rect 16396 5238 16448 5244
rect 16212 5228 16264 5234
rect 16212 5170 16264 5176
rect 16304 5228 16356 5234
rect 16304 5170 16356 5176
rect 15200 5160 15252 5166
rect 15200 5102 15252 5108
rect 15660 5160 15712 5166
rect 15660 5102 15712 5108
rect 16028 5160 16080 5166
rect 16080 5120 16160 5148
rect 16028 5102 16080 5108
rect 15212 4690 15240 5102
rect 16132 4690 16160 5120
rect 15200 4684 15252 4690
rect 15200 4626 15252 4632
rect 16120 4684 16172 4690
rect 16120 4626 16172 4632
rect 14740 4140 14792 4146
rect 14740 4082 14792 4088
rect 15384 4140 15436 4146
rect 15384 4082 15436 4088
rect 14464 4072 14516 4078
rect 14464 4014 14516 4020
rect 14476 3602 14504 4014
rect 14188 3596 14240 3602
rect 14188 3538 14240 3544
rect 14464 3596 14516 3602
rect 14464 3538 14516 3544
rect 14280 3528 14332 3534
rect 14280 3470 14332 3476
rect 13544 3052 13596 3058
rect 13544 2994 13596 3000
rect 13820 3052 13872 3058
rect 13820 2994 13872 3000
rect 11152 2984 11204 2990
rect 11152 2926 11204 2932
rect 12348 2984 12400 2990
rect 12348 2926 12400 2932
rect 12360 2836 12388 2926
rect 12440 2848 12492 2854
rect 12360 2808 12440 2836
rect 12440 2790 12492 2796
rect 14292 2514 14320 3470
rect 15200 2916 15252 2922
rect 15200 2858 15252 2864
rect 15212 2582 15240 2858
rect 15200 2576 15252 2582
rect 15200 2518 15252 2524
rect 8852 2508 8904 2514
rect 8852 2450 8904 2456
rect 10416 2508 10468 2514
rect 10416 2450 10468 2456
rect 11060 2508 11112 2514
rect 11060 2450 11112 2456
rect 14280 2508 14332 2514
rect 14280 2450 14332 2456
rect 8760 1828 8812 1834
rect 8760 1770 8812 1776
rect 8864 800 8892 2450
rect 11060 2304 11112 2310
rect 11060 2246 11112 2252
rect 13084 2304 13136 2310
rect 13084 2246 13136 2252
rect 11072 800 11100 2246
rect 13096 800 13124 2246
rect 15396 2088 15424 4082
rect 16224 3602 16252 5170
rect 16316 4146 16344 5170
rect 16776 5166 16804 6695
rect 16960 5642 16988 7398
rect 17052 6866 17080 7686
rect 17144 6866 17172 8366
rect 17236 7954 17264 8588
rect 17420 8430 17448 9590
rect 17408 8424 17460 8430
rect 17408 8366 17460 8372
rect 17224 7948 17276 7954
rect 17224 7890 17276 7896
rect 17236 7206 17264 7890
rect 17224 7200 17276 7206
rect 17224 7142 17276 7148
rect 17040 6860 17092 6866
rect 17040 6802 17092 6808
rect 17132 6860 17184 6866
rect 17132 6802 17184 6808
rect 17236 6798 17264 7142
rect 17224 6792 17276 6798
rect 17224 6734 17276 6740
rect 16948 5636 17000 5642
rect 16948 5578 17000 5584
rect 16764 5160 16816 5166
rect 16764 5102 16816 5108
rect 16488 5092 16540 5098
rect 16488 5034 16540 5040
rect 16856 5092 16908 5098
rect 16960 5080 16988 5578
rect 16908 5052 16988 5080
rect 16856 5034 16908 5040
rect 16304 4140 16356 4146
rect 16304 4082 16356 4088
rect 16212 3596 16264 3602
rect 16212 3538 16264 3544
rect 16304 3596 16356 3602
rect 16304 3538 16356 3544
rect 16316 3482 16344 3538
rect 16132 3454 16344 3482
rect 16132 3126 16160 3454
rect 16120 3120 16172 3126
rect 16120 3062 16172 3068
rect 16500 2650 16528 5034
rect 16868 4690 16896 5034
rect 17420 4758 17448 8366
rect 17512 7954 17540 16594
rect 17604 15638 17632 16782
rect 17684 16652 17736 16658
rect 17684 16594 17736 16600
rect 17592 15632 17644 15638
rect 17592 15574 17644 15580
rect 17696 15502 17724 16594
rect 17684 15496 17736 15502
rect 17684 15438 17736 15444
rect 17684 14884 17736 14890
rect 17684 14826 17736 14832
rect 17696 13870 17724 14826
rect 17684 13864 17736 13870
rect 17684 13806 17736 13812
rect 17788 12186 17816 17682
rect 17868 17536 17920 17542
rect 17868 17478 17920 17484
rect 17880 16726 17908 17478
rect 18156 17134 18184 18158
rect 18144 17128 18196 17134
rect 18144 17070 18196 17076
rect 17868 16720 17920 16726
rect 17868 16662 17920 16668
rect 17960 15564 18012 15570
rect 17960 15506 18012 15512
rect 17868 15088 17920 15094
rect 17868 15030 17920 15036
rect 17880 13394 17908 15030
rect 17972 14958 18000 15506
rect 18144 15496 18196 15502
rect 18142 15464 18144 15473
rect 18196 15464 18198 15473
rect 18142 15399 18198 15408
rect 17960 14952 18012 14958
rect 17960 14894 18012 14900
rect 17972 14822 18000 14894
rect 17960 14816 18012 14822
rect 17960 14758 18012 14764
rect 17972 14006 18000 14758
rect 18052 14408 18104 14414
rect 18052 14350 18104 14356
rect 18064 14006 18092 14350
rect 17960 14000 18012 14006
rect 17960 13942 18012 13948
rect 18052 14000 18104 14006
rect 18052 13942 18104 13948
rect 17868 13388 17920 13394
rect 17868 13330 17920 13336
rect 17604 12158 17816 12186
rect 17500 7948 17552 7954
rect 17500 7890 17552 7896
rect 17512 6934 17540 7890
rect 17604 7750 17632 12158
rect 17684 12096 17736 12102
rect 17684 12038 17736 12044
rect 17776 12096 17828 12102
rect 17776 12038 17828 12044
rect 17592 7744 17644 7750
rect 17592 7686 17644 7692
rect 17500 6928 17552 6934
rect 17500 6870 17552 6876
rect 17592 6860 17644 6866
rect 17592 6802 17644 6808
rect 17604 5914 17632 6802
rect 17592 5908 17644 5914
rect 17592 5850 17644 5856
rect 17592 5568 17644 5574
rect 17592 5510 17644 5516
rect 17604 5370 17632 5510
rect 17592 5364 17644 5370
rect 17592 5306 17644 5312
rect 17408 4752 17460 4758
rect 17408 4694 17460 4700
rect 16856 4684 16908 4690
rect 16856 4626 16908 4632
rect 17224 4072 17276 4078
rect 17696 4060 17724 12038
rect 17788 11830 17816 12038
rect 17776 11824 17828 11830
rect 17776 11766 17828 11772
rect 17868 11756 17920 11762
rect 17868 11698 17920 11704
rect 17880 10674 17908 11698
rect 17868 10668 17920 10674
rect 17868 10610 17920 10616
rect 17972 10538 18000 13942
rect 18156 12374 18184 15399
rect 18248 13530 18276 20470
rect 18340 18766 18368 22578
rect 18432 22574 18460 33798
rect 18512 32360 18564 32366
rect 18512 32302 18564 32308
rect 18524 32230 18552 32302
rect 18512 32224 18564 32230
rect 18512 32166 18564 32172
rect 18524 31482 18552 32166
rect 18604 31884 18656 31890
rect 18604 31826 18656 31832
rect 18512 31476 18564 31482
rect 18512 31418 18564 31424
rect 18616 31210 18644 31826
rect 18604 31204 18656 31210
rect 18604 31146 18656 31152
rect 18616 29073 18644 31146
rect 18602 29064 18658 29073
rect 18602 28999 18658 29008
rect 18800 28966 18828 37606
rect 19580 37564 19876 37584
rect 19636 37562 19660 37564
rect 19716 37562 19740 37564
rect 19796 37562 19820 37564
rect 19658 37510 19660 37562
rect 19722 37510 19734 37562
rect 19796 37510 19798 37562
rect 19636 37508 19660 37510
rect 19716 37508 19740 37510
rect 19796 37508 19820 37510
rect 19580 37488 19876 37508
rect 20168 37256 20220 37262
rect 20168 37198 20220 37204
rect 20180 36786 20208 37198
rect 20272 36938 20300 40200
rect 21456 37800 21508 37806
rect 21456 37742 21508 37748
rect 21824 37800 21876 37806
rect 21824 37742 21876 37748
rect 21468 37670 21496 37742
rect 21456 37664 21508 37670
rect 21456 37606 21508 37612
rect 21180 37256 21232 37262
rect 21180 37198 21232 37204
rect 20272 36922 20392 36938
rect 20272 36916 20404 36922
rect 20272 36910 20352 36916
rect 20352 36858 20404 36864
rect 20168 36780 20220 36786
rect 20168 36722 20220 36728
rect 20444 36712 20496 36718
rect 20444 36654 20496 36660
rect 20536 36712 20588 36718
rect 20536 36654 20588 36660
rect 20076 36644 20128 36650
rect 20076 36586 20128 36592
rect 19580 36476 19876 36496
rect 19636 36474 19660 36476
rect 19716 36474 19740 36476
rect 19796 36474 19820 36476
rect 19658 36422 19660 36474
rect 19722 36422 19734 36474
rect 19796 36422 19798 36474
rect 19636 36420 19660 36422
rect 19716 36420 19740 36422
rect 19796 36420 19820 36422
rect 19580 36400 19876 36420
rect 20088 36174 20116 36586
rect 20456 36310 20484 36654
rect 20444 36304 20496 36310
rect 20444 36246 20496 36252
rect 20076 36168 20128 36174
rect 20076 36110 20128 36116
rect 20088 35630 20116 36110
rect 20456 35698 20484 36246
rect 20444 35692 20496 35698
rect 20444 35634 20496 35640
rect 19248 35624 19300 35630
rect 19248 35566 19300 35572
rect 20076 35624 20128 35630
rect 20076 35566 20128 35572
rect 18972 34944 19024 34950
rect 18972 34886 19024 34892
rect 18984 34542 19012 34886
rect 18972 34536 19024 34542
rect 18972 34478 19024 34484
rect 19260 33318 19288 35566
rect 19580 35388 19876 35408
rect 19636 35386 19660 35388
rect 19716 35386 19740 35388
rect 19796 35386 19820 35388
rect 19658 35334 19660 35386
rect 19722 35334 19734 35386
rect 19796 35334 19798 35386
rect 19636 35332 19660 35334
rect 19716 35332 19740 35334
rect 19796 35332 19820 35334
rect 19580 35312 19876 35332
rect 20352 34604 20404 34610
rect 20352 34546 20404 34552
rect 19892 34536 19944 34542
rect 19892 34478 19944 34484
rect 20168 34536 20220 34542
rect 20168 34478 20220 34484
rect 19432 34468 19484 34474
rect 19432 34410 19484 34416
rect 19444 34066 19472 34410
rect 19580 34300 19876 34320
rect 19636 34298 19660 34300
rect 19716 34298 19740 34300
rect 19796 34298 19820 34300
rect 19658 34246 19660 34298
rect 19722 34246 19734 34298
rect 19796 34246 19798 34298
rect 19636 34244 19660 34246
rect 19716 34244 19740 34246
rect 19796 34244 19820 34246
rect 19580 34224 19876 34244
rect 19432 34060 19484 34066
rect 19432 34002 19484 34008
rect 19904 33998 19932 34478
rect 19892 33992 19944 33998
rect 19892 33934 19944 33940
rect 19248 33312 19300 33318
rect 19248 33254 19300 33260
rect 19580 33212 19876 33232
rect 19636 33210 19660 33212
rect 19716 33210 19740 33212
rect 19796 33210 19820 33212
rect 19658 33158 19660 33210
rect 19722 33158 19734 33210
rect 19796 33158 19798 33210
rect 19636 33156 19660 33158
rect 19716 33156 19740 33158
rect 19796 33156 19820 33158
rect 19580 33136 19876 33156
rect 19904 32978 19932 33934
rect 20180 33658 20208 34478
rect 20260 33856 20312 33862
rect 20260 33798 20312 33804
rect 20168 33652 20220 33658
rect 20168 33594 20220 33600
rect 19892 32972 19944 32978
rect 19892 32914 19944 32920
rect 18972 32904 19024 32910
rect 18972 32846 19024 32852
rect 18984 32502 19012 32846
rect 19156 32768 19208 32774
rect 19156 32710 19208 32716
rect 18972 32496 19024 32502
rect 18972 32438 19024 32444
rect 18880 32360 18932 32366
rect 18880 32302 18932 32308
rect 18892 32026 18920 32302
rect 18880 32020 18932 32026
rect 18880 31962 18932 31968
rect 19168 31890 19196 32710
rect 19580 32124 19876 32144
rect 19636 32122 19660 32124
rect 19716 32122 19740 32124
rect 19796 32122 19820 32124
rect 19658 32070 19660 32122
rect 19722 32070 19734 32122
rect 19796 32070 19798 32122
rect 19636 32068 19660 32070
rect 19716 32068 19740 32070
rect 19796 32068 19820 32070
rect 19580 32048 19876 32068
rect 19156 31884 19208 31890
rect 19208 31844 19288 31872
rect 19156 31826 19208 31832
rect 19156 31272 19208 31278
rect 19156 31214 19208 31220
rect 19168 30802 19196 31214
rect 19156 30796 19208 30802
rect 19156 30738 19208 30744
rect 19168 30122 19196 30738
rect 19260 30258 19288 31844
rect 19432 31340 19484 31346
rect 19432 31282 19484 31288
rect 19444 30802 19472 31282
rect 19892 31272 19944 31278
rect 19892 31214 19944 31220
rect 19580 31036 19876 31056
rect 19636 31034 19660 31036
rect 19716 31034 19740 31036
rect 19796 31034 19820 31036
rect 19658 30982 19660 31034
rect 19722 30982 19734 31034
rect 19796 30982 19798 31034
rect 19636 30980 19660 30982
rect 19716 30980 19740 30982
rect 19796 30980 19820 30982
rect 19580 30960 19876 30980
rect 19904 30802 19932 31214
rect 19432 30796 19484 30802
rect 19432 30738 19484 30744
rect 19892 30796 19944 30802
rect 19892 30738 19944 30744
rect 19340 30388 19392 30394
rect 19340 30330 19392 30336
rect 19248 30252 19300 30258
rect 19248 30194 19300 30200
rect 19156 30116 19208 30122
rect 19156 30058 19208 30064
rect 19064 29708 19116 29714
rect 19064 29650 19116 29656
rect 19076 29102 19104 29650
rect 19168 29510 19196 30058
rect 19156 29504 19208 29510
rect 19156 29446 19208 29452
rect 18972 29096 19024 29102
rect 18972 29038 19024 29044
rect 19064 29096 19116 29102
rect 19064 29038 19116 29044
rect 18512 28960 18564 28966
rect 18512 28902 18564 28908
rect 18788 28960 18840 28966
rect 18880 28960 18932 28966
rect 18788 28902 18840 28908
rect 18878 28928 18880 28937
rect 18932 28928 18934 28937
rect 18524 28626 18552 28902
rect 18878 28863 18934 28872
rect 18512 28620 18564 28626
rect 18512 28562 18564 28568
rect 18510 28520 18566 28529
rect 18510 28455 18566 28464
rect 18524 26790 18552 28455
rect 18984 26994 19012 29038
rect 19076 27674 19104 29038
rect 19064 27668 19116 27674
rect 19064 27610 19116 27616
rect 19168 27538 19196 29446
rect 19260 28558 19288 30194
rect 19352 29646 19380 30330
rect 19904 30258 19932 30738
rect 19892 30252 19944 30258
rect 19892 30194 19944 30200
rect 19580 29948 19876 29968
rect 19636 29946 19660 29948
rect 19716 29946 19740 29948
rect 19796 29946 19820 29948
rect 19658 29894 19660 29946
rect 19722 29894 19734 29946
rect 19796 29894 19798 29946
rect 19636 29892 19660 29894
rect 19716 29892 19740 29894
rect 19796 29892 19820 29894
rect 19580 29872 19876 29892
rect 19340 29640 19392 29646
rect 19340 29582 19392 29588
rect 19248 28552 19300 28558
rect 19248 28494 19300 28500
rect 19248 28416 19300 28422
rect 19248 28358 19300 28364
rect 19156 27532 19208 27538
rect 19156 27474 19208 27480
rect 18972 26988 19024 26994
rect 18972 26930 19024 26936
rect 19064 26920 19116 26926
rect 19064 26862 19116 26868
rect 18512 26784 18564 26790
rect 18512 26726 18564 26732
rect 19076 26450 19104 26862
rect 18604 26444 18656 26450
rect 18604 26386 18656 26392
rect 19064 26444 19116 26450
rect 19064 26386 19116 26392
rect 18616 26246 18644 26386
rect 18604 26240 18656 26246
rect 18604 26182 18656 26188
rect 18616 25820 18644 26182
rect 18696 25832 18748 25838
rect 18616 25792 18696 25820
rect 18696 25774 18748 25780
rect 19156 25832 19208 25838
rect 19156 25774 19208 25780
rect 19168 25362 19196 25774
rect 19260 25430 19288 28358
rect 19352 27538 19380 29582
rect 19432 29028 19484 29034
rect 19432 28970 19484 28976
rect 19444 27946 19472 28970
rect 19580 28860 19876 28880
rect 19636 28858 19660 28860
rect 19716 28858 19740 28860
rect 19796 28858 19820 28860
rect 19658 28806 19660 28858
rect 19722 28806 19734 28858
rect 19796 28806 19798 28858
rect 19636 28804 19660 28806
rect 19716 28804 19740 28806
rect 19796 28804 19820 28806
rect 19580 28784 19876 28804
rect 19432 27940 19484 27946
rect 19432 27882 19484 27888
rect 19580 27772 19876 27792
rect 19636 27770 19660 27772
rect 19716 27770 19740 27772
rect 19796 27770 19820 27772
rect 19658 27718 19660 27770
rect 19722 27718 19734 27770
rect 19796 27718 19798 27770
rect 19636 27716 19660 27718
rect 19716 27716 19740 27718
rect 19796 27716 19820 27718
rect 19580 27696 19876 27716
rect 19340 27532 19392 27538
rect 19340 27474 19392 27480
rect 19904 27470 19932 30194
rect 20168 30184 20220 30190
rect 20168 30126 20220 30132
rect 19984 29708 20036 29714
rect 19984 29650 20036 29656
rect 19996 28422 20024 29650
rect 20180 29238 20208 30126
rect 20168 29232 20220 29238
rect 20168 29174 20220 29180
rect 20180 28966 20208 29174
rect 20168 28960 20220 28966
rect 20168 28902 20220 28908
rect 20076 28688 20128 28694
rect 20076 28630 20128 28636
rect 19984 28416 20036 28422
rect 19984 28358 20036 28364
rect 19892 27464 19944 27470
rect 19892 27406 19944 27412
rect 19432 26920 19484 26926
rect 19432 26862 19484 26868
rect 19444 26500 19472 26862
rect 19580 26684 19876 26704
rect 19636 26682 19660 26684
rect 19716 26682 19740 26684
rect 19796 26682 19820 26684
rect 19658 26630 19660 26682
rect 19722 26630 19734 26682
rect 19796 26630 19798 26682
rect 19636 26628 19660 26630
rect 19716 26628 19740 26630
rect 19796 26628 19820 26630
rect 19580 26608 19876 26628
rect 19444 26472 19564 26500
rect 19432 26240 19484 26246
rect 19432 26182 19484 26188
rect 19536 26194 19564 26472
rect 19904 26450 19932 27406
rect 19996 26858 20024 28358
rect 20088 27010 20116 28630
rect 20088 26982 20208 27010
rect 20076 26920 20128 26926
rect 20076 26862 20128 26868
rect 19984 26852 20036 26858
rect 19984 26794 20036 26800
rect 19892 26444 19944 26450
rect 19720 26404 19892 26432
rect 19340 25900 19392 25906
rect 19340 25842 19392 25848
rect 19352 25498 19380 25842
rect 19444 25498 19472 26182
rect 19536 26166 19656 26194
rect 19628 25838 19656 26166
rect 19616 25832 19668 25838
rect 19616 25774 19668 25780
rect 19720 25770 19748 26404
rect 19892 26386 19944 26392
rect 19984 26444 20036 26450
rect 19984 26386 20036 26392
rect 19996 25906 20024 26386
rect 20088 26314 20116 26862
rect 20076 26308 20128 26314
rect 20076 26250 20128 26256
rect 19984 25900 20036 25906
rect 19984 25842 20036 25848
rect 19892 25832 19944 25838
rect 19892 25774 19944 25780
rect 19708 25764 19760 25770
rect 19708 25706 19760 25712
rect 19580 25596 19876 25616
rect 19636 25594 19660 25596
rect 19716 25594 19740 25596
rect 19796 25594 19820 25596
rect 19658 25542 19660 25594
rect 19722 25542 19734 25594
rect 19796 25542 19798 25594
rect 19636 25540 19660 25542
rect 19716 25540 19740 25542
rect 19796 25540 19820 25542
rect 19580 25520 19876 25540
rect 19340 25492 19392 25498
rect 19340 25434 19392 25440
rect 19432 25492 19484 25498
rect 19432 25434 19484 25440
rect 19248 25424 19300 25430
rect 19248 25366 19300 25372
rect 19156 25356 19208 25362
rect 19156 25298 19208 25304
rect 19432 25356 19484 25362
rect 19432 25298 19484 25304
rect 18512 25288 18564 25294
rect 18512 25230 18564 25236
rect 18524 24954 18552 25230
rect 18512 24948 18564 24954
rect 18512 24890 18564 24896
rect 19444 24614 19472 25298
rect 19432 24608 19484 24614
rect 19432 24550 19484 24556
rect 19580 24508 19876 24528
rect 19636 24506 19660 24508
rect 19716 24506 19740 24508
rect 19796 24506 19820 24508
rect 19658 24454 19660 24506
rect 19722 24454 19734 24506
rect 19796 24454 19798 24506
rect 19636 24452 19660 24454
rect 19716 24452 19740 24454
rect 19796 24452 19820 24454
rect 19580 24432 19876 24452
rect 18512 24336 18564 24342
rect 18510 24304 18512 24313
rect 18564 24304 18566 24313
rect 19904 24274 19932 25774
rect 19984 25764 20036 25770
rect 19984 25706 20036 25712
rect 18510 24239 18566 24248
rect 19892 24268 19944 24274
rect 19892 24210 19944 24216
rect 19340 24132 19392 24138
rect 19340 24074 19392 24080
rect 19352 23866 19380 24074
rect 19340 23860 19392 23866
rect 19340 23802 19392 23808
rect 18880 23656 18932 23662
rect 18880 23598 18932 23604
rect 18892 23361 18920 23598
rect 19580 23420 19876 23440
rect 19636 23418 19660 23420
rect 19716 23418 19740 23420
rect 19796 23418 19820 23420
rect 19658 23366 19660 23418
rect 19722 23366 19734 23418
rect 19796 23366 19798 23418
rect 19636 23364 19660 23366
rect 19716 23364 19740 23366
rect 19796 23364 19820 23366
rect 18878 23352 18934 23361
rect 19580 23344 19876 23364
rect 18878 23287 18934 23296
rect 19248 23248 19300 23254
rect 18878 23216 18934 23225
rect 18696 23180 18748 23186
rect 19248 23190 19300 23196
rect 18878 23151 18934 23160
rect 18696 23122 18748 23128
rect 18420 22568 18472 22574
rect 18420 22510 18472 22516
rect 18708 22506 18736 23122
rect 18696 22500 18748 22506
rect 18696 22442 18748 22448
rect 18420 20324 18472 20330
rect 18420 20266 18472 20272
rect 18432 19961 18460 20266
rect 18418 19952 18474 19961
rect 18418 19887 18474 19896
rect 18696 19712 18748 19718
rect 18696 19654 18748 19660
rect 18708 19310 18736 19654
rect 18696 19304 18748 19310
rect 18696 19246 18748 19252
rect 18420 19168 18472 19174
rect 18420 19110 18472 19116
rect 18328 18760 18380 18766
rect 18328 18702 18380 18708
rect 18340 18306 18368 18702
rect 18432 18630 18460 19110
rect 18420 18624 18472 18630
rect 18420 18566 18472 18572
rect 18340 18278 18460 18306
rect 18708 18290 18736 19246
rect 18328 18216 18380 18222
rect 18328 18158 18380 18164
rect 18340 17542 18368 18158
rect 18328 17536 18380 17542
rect 18328 17478 18380 17484
rect 18432 16658 18460 18278
rect 18696 18284 18748 18290
rect 18696 18226 18748 18232
rect 18604 17672 18656 17678
rect 18604 17614 18656 17620
rect 18616 17270 18644 17614
rect 18604 17264 18656 17270
rect 18604 17206 18656 17212
rect 18708 17202 18736 18226
rect 18892 17864 18920 23151
rect 19156 22432 19208 22438
rect 19156 22374 19208 22380
rect 19168 22098 19196 22374
rect 19156 22092 19208 22098
rect 19156 22034 19208 22040
rect 19168 21554 19196 22034
rect 19260 21554 19288 23190
rect 19580 22332 19876 22352
rect 19636 22330 19660 22332
rect 19716 22330 19740 22332
rect 19796 22330 19820 22332
rect 19658 22278 19660 22330
rect 19722 22278 19734 22330
rect 19796 22278 19798 22330
rect 19636 22276 19660 22278
rect 19716 22276 19740 22278
rect 19796 22276 19820 22278
rect 19580 22256 19876 22276
rect 19340 22092 19392 22098
rect 19340 22034 19392 22040
rect 19432 22092 19484 22098
rect 19432 22034 19484 22040
rect 19352 21690 19380 22034
rect 19444 21894 19472 22034
rect 19432 21888 19484 21894
rect 19432 21830 19484 21836
rect 19340 21684 19392 21690
rect 19340 21626 19392 21632
rect 19904 21593 19932 24210
rect 19996 23798 20024 25706
rect 20088 25430 20116 26250
rect 20076 25424 20128 25430
rect 20076 25366 20128 25372
rect 20076 24268 20128 24274
rect 20076 24210 20128 24216
rect 19984 23792 20036 23798
rect 19984 23734 20036 23740
rect 20088 23662 20116 24210
rect 20076 23656 20128 23662
rect 20076 23598 20128 23604
rect 19984 23520 20036 23526
rect 19984 23462 20036 23468
rect 19890 21584 19946 21593
rect 19156 21548 19208 21554
rect 19156 21490 19208 21496
rect 19248 21548 19300 21554
rect 19890 21519 19946 21528
rect 19248 21490 19300 21496
rect 19168 20942 19196 21490
rect 19432 21480 19484 21486
rect 19432 21422 19484 21428
rect 19248 21412 19300 21418
rect 19248 21354 19300 21360
rect 19156 20936 19208 20942
rect 19156 20878 19208 20884
rect 19168 20058 19196 20878
rect 19156 20052 19208 20058
rect 19156 19994 19208 20000
rect 19260 19990 19288 21354
rect 19444 21350 19472 21422
rect 19892 21412 19944 21418
rect 19892 21354 19944 21360
rect 19340 21344 19392 21350
rect 19340 21286 19392 21292
rect 19432 21344 19484 21350
rect 19432 21286 19484 21292
rect 19352 21078 19380 21286
rect 19580 21244 19876 21264
rect 19636 21242 19660 21244
rect 19716 21242 19740 21244
rect 19796 21242 19820 21244
rect 19658 21190 19660 21242
rect 19722 21190 19734 21242
rect 19796 21190 19798 21242
rect 19636 21188 19660 21190
rect 19716 21188 19740 21190
rect 19796 21188 19820 21190
rect 19580 21168 19876 21188
rect 19904 21078 19932 21354
rect 19340 21072 19392 21078
rect 19340 21014 19392 21020
rect 19892 21072 19944 21078
rect 19892 21014 19944 21020
rect 19248 19984 19300 19990
rect 19248 19926 19300 19932
rect 19352 19922 19380 21014
rect 19892 20800 19944 20806
rect 19892 20742 19944 20748
rect 19432 20256 19484 20262
rect 19432 20198 19484 20204
rect 19340 19916 19392 19922
rect 19340 19858 19392 19864
rect 19444 19786 19472 20198
rect 19580 20156 19876 20176
rect 19636 20154 19660 20156
rect 19716 20154 19740 20156
rect 19796 20154 19820 20156
rect 19658 20102 19660 20154
rect 19722 20102 19734 20154
rect 19796 20102 19798 20154
rect 19636 20100 19660 20102
rect 19716 20100 19740 20102
rect 19796 20100 19820 20102
rect 19580 20080 19876 20100
rect 19432 19780 19484 19786
rect 19432 19722 19484 19728
rect 18972 19304 19024 19310
rect 18972 19246 19024 19252
rect 19064 19304 19116 19310
rect 19064 19246 19116 19252
rect 18984 18902 19012 19246
rect 18972 18896 19024 18902
rect 18972 18838 19024 18844
rect 19076 18834 19104 19246
rect 19248 19168 19300 19174
rect 19248 19110 19300 19116
rect 19340 19168 19392 19174
rect 19340 19110 19392 19116
rect 19064 18828 19116 18834
rect 19064 18770 19116 18776
rect 19260 18766 19288 19110
rect 19352 18834 19380 19110
rect 19580 19068 19876 19088
rect 19636 19066 19660 19068
rect 19716 19066 19740 19068
rect 19796 19066 19820 19068
rect 19658 19014 19660 19066
rect 19722 19014 19734 19066
rect 19796 19014 19798 19066
rect 19636 19012 19660 19014
rect 19716 19012 19740 19014
rect 19796 19012 19820 19014
rect 19580 18992 19876 19012
rect 19340 18828 19392 18834
rect 19340 18770 19392 18776
rect 19524 18828 19576 18834
rect 19524 18770 19576 18776
rect 19708 18828 19760 18834
rect 19708 18770 19760 18776
rect 19248 18760 19300 18766
rect 19248 18702 19300 18708
rect 19536 18426 19564 18770
rect 19720 18426 19748 18770
rect 19524 18420 19576 18426
rect 19524 18362 19576 18368
rect 19708 18420 19760 18426
rect 19708 18362 19760 18368
rect 19340 18080 19392 18086
rect 19340 18022 19392 18028
rect 18800 17836 18920 17864
rect 18696 17196 18748 17202
rect 18696 17138 18748 17144
rect 18420 16652 18472 16658
rect 18420 16594 18472 16600
rect 18512 16652 18564 16658
rect 18512 16594 18564 16600
rect 18328 16584 18380 16590
rect 18328 16526 18380 16532
rect 18340 16114 18368 16526
rect 18328 16108 18380 16114
rect 18328 16050 18380 16056
rect 18432 14906 18460 16594
rect 18524 15638 18552 16594
rect 18708 16046 18736 17138
rect 18696 16040 18748 16046
rect 18696 15982 18748 15988
rect 18512 15632 18564 15638
rect 18512 15574 18564 15580
rect 18524 15026 18552 15574
rect 18708 15570 18736 15982
rect 18696 15564 18748 15570
rect 18696 15506 18748 15512
rect 18512 15020 18564 15026
rect 18512 14962 18564 14968
rect 18340 14878 18460 14906
rect 18340 13530 18368 14878
rect 18420 14816 18472 14822
rect 18420 14758 18472 14764
rect 18432 13870 18460 14758
rect 18524 14618 18552 14962
rect 18512 14612 18564 14618
rect 18512 14554 18564 14560
rect 18708 14414 18736 15506
rect 18696 14408 18748 14414
rect 18602 14376 18658 14385
rect 18696 14350 18748 14356
rect 18602 14311 18658 14320
rect 18420 13864 18472 13870
rect 18420 13806 18472 13812
rect 18236 13524 18288 13530
rect 18236 13466 18288 13472
rect 18328 13524 18380 13530
rect 18328 13466 18380 13472
rect 18236 13388 18288 13394
rect 18236 13330 18288 13336
rect 18144 12368 18196 12374
rect 18144 12310 18196 12316
rect 18248 11898 18276 13330
rect 18328 13320 18380 13326
rect 18328 13262 18380 13268
rect 18340 12986 18368 13262
rect 18328 12980 18380 12986
rect 18328 12922 18380 12928
rect 18418 12608 18474 12617
rect 18418 12543 18474 12552
rect 18432 12306 18460 12543
rect 18420 12300 18472 12306
rect 18420 12242 18472 12248
rect 18236 11892 18288 11898
rect 18236 11834 18288 11840
rect 18432 10606 18460 12242
rect 18512 11688 18564 11694
rect 18512 11630 18564 11636
rect 18524 11218 18552 11630
rect 18512 11212 18564 11218
rect 18512 11154 18564 11160
rect 18420 10600 18472 10606
rect 18420 10542 18472 10548
rect 17960 10532 18012 10538
rect 17960 10474 18012 10480
rect 17972 10130 18000 10474
rect 17960 10124 18012 10130
rect 17960 10066 18012 10072
rect 18328 10056 18380 10062
rect 18328 9998 18380 10004
rect 18340 9178 18368 9998
rect 18420 9920 18472 9926
rect 18420 9862 18472 9868
rect 18432 9518 18460 9862
rect 18616 9654 18644 14311
rect 18800 13841 18828 17836
rect 18880 17740 18932 17746
rect 18880 17682 18932 17688
rect 18892 14906 18920 17682
rect 19156 17604 19208 17610
rect 19156 17546 19208 17552
rect 19168 17202 19196 17546
rect 19156 17196 19208 17202
rect 19156 17138 19208 17144
rect 19352 16590 19380 18022
rect 19580 17980 19876 18000
rect 19636 17978 19660 17980
rect 19716 17978 19740 17980
rect 19796 17978 19820 17980
rect 19658 17926 19660 17978
rect 19722 17926 19734 17978
rect 19796 17926 19798 17978
rect 19636 17924 19660 17926
rect 19716 17924 19740 17926
rect 19796 17924 19820 17926
rect 19580 17904 19876 17924
rect 19580 16892 19876 16912
rect 19636 16890 19660 16892
rect 19716 16890 19740 16892
rect 19796 16890 19820 16892
rect 19658 16838 19660 16890
rect 19722 16838 19734 16890
rect 19796 16838 19798 16890
rect 19636 16836 19660 16838
rect 19716 16836 19740 16838
rect 19796 16836 19820 16838
rect 19580 16816 19876 16836
rect 19340 16584 19392 16590
rect 19340 16526 19392 16532
rect 19352 16454 19380 16526
rect 19340 16448 19392 16454
rect 19340 16390 19392 16396
rect 19904 15978 19932 20742
rect 19996 18766 20024 23462
rect 20088 21690 20116 23598
rect 20180 23526 20208 26982
rect 20168 23520 20220 23526
rect 20168 23462 20220 23468
rect 20272 23050 20300 33798
rect 20364 33522 20392 34546
rect 20352 33516 20404 33522
rect 20352 33458 20404 33464
rect 20364 28694 20392 33458
rect 20548 33454 20576 36654
rect 21192 36582 21220 37198
rect 20904 36576 20956 36582
rect 20904 36518 20956 36524
rect 21180 36576 21232 36582
rect 21180 36518 21232 36524
rect 20916 36242 20944 36518
rect 20904 36236 20956 36242
rect 20904 36178 20956 36184
rect 20812 36032 20864 36038
rect 20812 35974 20864 35980
rect 20996 36032 21048 36038
rect 20996 35974 21048 35980
rect 20824 33454 20852 35974
rect 21008 35630 21036 35974
rect 21468 35698 21496 37606
rect 21836 37466 21864 37742
rect 21824 37460 21876 37466
rect 21824 37402 21876 37408
rect 22480 36854 22508 40200
rect 24216 37800 24268 37806
rect 24216 37742 24268 37748
rect 23296 37732 23348 37738
rect 23296 37674 23348 37680
rect 23020 37664 23072 37670
rect 23020 37606 23072 37612
rect 23032 37262 23060 37606
rect 23308 37330 23336 37674
rect 24228 37466 24256 37742
rect 24216 37460 24268 37466
rect 24216 37402 24268 37408
rect 23296 37324 23348 37330
rect 23296 37266 23348 37272
rect 23020 37256 23072 37262
rect 23020 37198 23072 37204
rect 22468 36848 22520 36854
rect 22468 36790 22520 36796
rect 24216 36848 24268 36854
rect 24216 36790 24268 36796
rect 22468 36712 22520 36718
rect 22468 36654 22520 36660
rect 22836 36712 22888 36718
rect 22836 36654 22888 36660
rect 22376 36576 22428 36582
rect 22376 36518 22428 36524
rect 22388 35698 22416 36518
rect 22480 35834 22508 36654
rect 22652 36236 22704 36242
rect 22652 36178 22704 36184
rect 22664 35834 22692 36178
rect 22848 36106 22876 36654
rect 23112 36236 23164 36242
rect 23112 36178 23164 36184
rect 22836 36100 22888 36106
rect 22836 36042 22888 36048
rect 22468 35828 22520 35834
rect 22468 35770 22520 35776
rect 22652 35828 22704 35834
rect 22652 35770 22704 35776
rect 21456 35692 21508 35698
rect 21456 35634 21508 35640
rect 22376 35692 22428 35698
rect 22376 35634 22428 35640
rect 20996 35624 21048 35630
rect 20996 35566 21048 35572
rect 22664 35154 22692 35770
rect 23124 35154 23152 36178
rect 24124 36168 24176 36174
rect 24124 36110 24176 36116
rect 23940 35624 23992 35630
rect 23940 35566 23992 35572
rect 23952 35154 23980 35566
rect 24136 35494 24164 36110
rect 24124 35488 24176 35494
rect 24124 35430 24176 35436
rect 22652 35148 22704 35154
rect 22652 35090 22704 35096
rect 23112 35148 23164 35154
rect 23112 35090 23164 35096
rect 23388 35148 23440 35154
rect 23388 35090 23440 35096
rect 23940 35148 23992 35154
rect 23940 35090 23992 35096
rect 20904 35080 20956 35086
rect 20904 35022 20956 35028
rect 22100 35080 22152 35086
rect 22100 35022 22152 35028
rect 20536 33448 20588 33454
rect 20536 33390 20588 33396
rect 20812 33448 20864 33454
rect 20812 33390 20864 33396
rect 20444 32972 20496 32978
rect 20444 32914 20496 32920
rect 20456 32434 20484 32914
rect 20444 32428 20496 32434
rect 20444 32370 20496 32376
rect 20456 31754 20484 32370
rect 20720 32360 20772 32366
rect 20720 32302 20772 32308
rect 20444 31748 20496 31754
rect 20444 31690 20496 31696
rect 20732 31686 20760 32302
rect 20720 31680 20772 31686
rect 20720 31622 20772 31628
rect 20444 31272 20496 31278
rect 20444 31214 20496 31220
rect 20456 30394 20484 31214
rect 20444 30388 20496 30394
rect 20444 30330 20496 30336
rect 20444 29096 20496 29102
rect 20444 29038 20496 29044
rect 20352 28688 20404 28694
rect 20352 28630 20404 28636
rect 20352 28008 20404 28014
rect 20352 27950 20404 27956
rect 20364 26518 20392 27950
rect 20456 27062 20484 29038
rect 20628 28960 20680 28966
rect 20628 28902 20680 28908
rect 20536 28144 20588 28150
rect 20536 28086 20588 28092
rect 20444 27056 20496 27062
rect 20444 26998 20496 27004
rect 20548 26994 20576 28086
rect 20640 27674 20668 28902
rect 20628 27668 20680 27674
rect 20628 27610 20680 27616
rect 20628 27056 20680 27062
rect 20628 26998 20680 27004
rect 20536 26988 20588 26994
rect 20536 26930 20588 26936
rect 20444 26920 20496 26926
rect 20444 26862 20496 26868
rect 20456 26586 20484 26862
rect 20444 26580 20496 26586
rect 20444 26522 20496 26528
rect 20352 26512 20404 26518
rect 20352 26454 20404 26460
rect 20444 25832 20496 25838
rect 20444 25774 20496 25780
rect 20456 25294 20484 25774
rect 20444 25288 20496 25294
rect 20444 25230 20496 25236
rect 20640 24138 20668 26998
rect 20812 26920 20864 26926
rect 20812 26862 20864 26868
rect 20824 26518 20852 26862
rect 20812 26512 20864 26518
rect 20812 26454 20864 26460
rect 20824 25362 20852 26454
rect 20812 25356 20864 25362
rect 20812 25298 20864 25304
rect 20824 24886 20852 25298
rect 20812 24880 20864 24886
rect 20812 24822 20864 24828
rect 20812 24744 20864 24750
rect 20812 24686 20864 24692
rect 20720 24676 20772 24682
rect 20720 24618 20772 24624
rect 20732 24410 20760 24618
rect 20720 24404 20772 24410
rect 20720 24346 20772 24352
rect 20628 24132 20680 24138
rect 20824 24120 20852 24686
rect 20628 24074 20680 24080
rect 20732 24092 20852 24120
rect 20732 23662 20760 24092
rect 20720 23656 20772 23662
rect 20720 23598 20772 23604
rect 20732 23526 20760 23598
rect 20720 23520 20772 23526
rect 20720 23462 20772 23468
rect 20352 23112 20404 23118
rect 20352 23054 20404 23060
rect 20260 23044 20312 23050
rect 20260 22986 20312 22992
rect 20260 22092 20312 22098
rect 20260 22034 20312 22040
rect 20076 21684 20128 21690
rect 20076 21626 20128 21632
rect 20074 21584 20130 21593
rect 20074 21519 20130 21528
rect 20088 20806 20116 21519
rect 20168 21480 20220 21486
rect 20168 21422 20220 21428
rect 20180 21010 20208 21422
rect 20168 21004 20220 21010
rect 20168 20946 20220 20952
rect 20272 20942 20300 22034
rect 20260 20936 20312 20942
rect 20260 20878 20312 20884
rect 20076 20800 20128 20806
rect 20076 20742 20128 20748
rect 20260 20596 20312 20602
rect 20260 20538 20312 20544
rect 20272 19922 20300 20538
rect 20260 19916 20312 19922
rect 20260 19858 20312 19864
rect 19984 18760 20036 18766
rect 19984 18702 20036 18708
rect 19996 18630 20024 18702
rect 19984 18624 20036 18630
rect 19984 18566 20036 18572
rect 20076 17740 20128 17746
rect 20076 17682 20128 17688
rect 19984 16788 20036 16794
rect 19984 16730 20036 16736
rect 19996 16017 20024 16730
rect 19982 16008 20038 16017
rect 19892 15972 19944 15978
rect 19982 15943 20038 15952
rect 19892 15914 19944 15920
rect 19432 15904 19484 15910
rect 19432 15846 19484 15852
rect 18972 15496 19024 15502
rect 18972 15438 19024 15444
rect 18984 15026 19012 15438
rect 19444 15162 19472 15846
rect 19580 15804 19876 15824
rect 19636 15802 19660 15804
rect 19716 15802 19740 15804
rect 19796 15802 19820 15804
rect 19658 15750 19660 15802
rect 19722 15750 19734 15802
rect 19796 15750 19798 15802
rect 19636 15748 19660 15750
rect 19716 15748 19740 15750
rect 19796 15748 19820 15750
rect 19580 15728 19876 15748
rect 19432 15156 19484 15162
rect 19432 15098 19484 15104
rect 19340 15088 19392 15094
rect 19340 15030 19392 15036
rect 18972 15020 19024 15026
rect 18972 14962 19024 14968
rect 19352 14958 19380 15030
rect 19340 14952 19392 14958
rect 18892 14878 19012 14906
rect 19340 14894 19392 14900
rect 19984 14952 20036 14958
rect 19984 14894 20036 14900
rect 18880 14544 18932 14550
rect 18880 14486 18932 14492
rect 18892 13870 18920 14486
rect 18880 13864 18932 13870
rect 18786 13832 18842 13841
rect 18880 13806 18932 13812
rect 18786 13767 18842 13776
rect 18880 12776 18932 12782
rect 18880 12718 18932 12724
rect 18892 11354 18920 12718
rect 18880 11348 18932 11354
rect 18880 11290 18932 11296
rect 18604 9648 18656 9654
rect 18604 9590 18656 9596
rect 18420 9512 18472 9518
rect 18420 9454 18472 9460
rect 18788 9512 18840 9518
rect 18788 9454 18840 9460
rect 18328 9172 18380 9178
rect 18328 9114 18380 9120
rect 18052 8832 18104 8838
rect 18052 8774 18104 8780
rect 18064 8430 18092 8774
rect 18800 8498 18828 9454
rect 18788 8492 18840 8498
rect 18788 8434 18840 8440
rect 18052 8424 18104 8430
rect 18052 8366 18104 8372
rect 18788 8288 18840 8294
rect 18788 8230 18840 8236
rect 18800 7954 18828 8230
rect 18880 8084 18932 8090
rect 18880 8026 18932 8032
rect 18892 7954 18920 8026
rect 18788 7948 18840 7954
rect 18788 7890 18840 7896
rect 18880 7948 18932 7954
rect 18880 7890 18932 7896
rect 17868 7744 17920 7750
rect 17868 7686 17920 7692
rect 17776 6112 17828 6118
rect 17776 6054 17828 6060
rect 17788 5846 17816 6054
rect 17776 5840 17828 5846
rect 17776 5782 17828 5788
rect 17788 5166 17816 5782
rect 17776 5160 17828 5166
rect 17776 5102 17828 5108
rect 17774 4176 17830 4185
rect 17774 4111 17776 4120
rect 17828 4111 17830 4120
rect 17776 4082 17828 4088
rect 17276 4032 17724 4060
rect 17224 4014 17276 4020
rect 17880 3942 17908 7686
rect 18892 7410 18920 7890
rect 18144 7404 18196 7410
rect 18144 7346 18196 7352
rect 18880 7404 18932 7410
rect 18880 7346 18932 7352
rect 18156 6866 18184 7346
rect 18420 6928 18472 6934
rect 18420 6870 18472 6876
rect 18144 6860 18196 6866
rect 18144 6802 18196 6808
rect 18432 6254 18460 6870
rect 18420 6248 18472 6254
rect 18420 6190 18472 6196
rect 17960 6180 18012 6186
rect 17960 6122 18012 6128
rect 17972 5778 18000 6122
rect 17960 5772 18012 5778
rect 17960 5714 18012 5720
rect 17960 5568 18012 5574
rect 17960 5510 18012 5516
rect 17972 4622 18000 5510
rect 18696 5160 18748 5166
rect 18696 5102 18748 5108
rect 18052 5024 18104 5030
rect 18052 4966 18104 4972
rect 17960 4616 18012 4622
rect 17960 4558 18012 4564
rect 17868 3936 17920 3942
rect 17868 3878 17920 3884
rect 17972 3534 18000 4558
rect 18064 3602 18092 4966
rect 18708 4078 18736 5102
rect 18696 4072 18748 4078
rect 18696 4014 18748 4020
rect 18144 4004 18196 4010
rect 18144 3946 18196 3952
rect 18052 3596 18104 3602
rect 18052 3538 18104 3544
rect 17960 3528 18012 3534
rect 17960 3470 18012 3476
rect 16580 3392 16632 3398
rect 16580 3334 16632 3340
rect 16592 3058 16620 3334
rect 16580 3052 16632 3058
rect 16580 2994 16632 3000
rect 17224 2916 17276 2922
rect 17224 2858 17276 2864
rect 16488 2644 16540 2650
rect 16488 2586 16540 2592
rect 17236 2514 17264 2858
rect 17224 2508 17276 2514
rect 17224 2450 17276 2456
rect 18064 2446 18092 3538
rect 18156 2990 18184 3946
rect 18984 3942 19012 14878
rect 19154 14784 19210 14793
rect 19154 14719 19210 14728
rect 19168 13802 19196 14719
rect 19352 14521 19380 14894
rect 19580 14716 19876 14736
rect 19636 14714 19660 14716
rect 19716 14714 19740 14716
rect 19796 14714 19820 14716
rect 19658 14662 19660 14714
rect 19722 14662 19734 14714
rect 19796 14662 19798 14714
rect 19636 14660 19660 14662
rect 19716 14660 19740 14662
rect 19796 14660 19820 14662
rect 19580 14640 19876 14660
rect 19338 14512 19394 14521
rect 19338 14447 19394 14456
rect 19706 14512 19762 14521
rect 19706 14447 19708 14456
rect 19760 14447 19762 14456
rect 19708 14418 19760 14424
rect 19432 14272 19484 14278
rect 19432 14214 19484 14220
rect 19248 14068 19300 14074
rect 19248 14010 19300 14016
rect 19260 13870 19288 14010
rect 19248 13864 19300 13870
rect 19248 13806 19300 13812
rect 19156 13796 19208 13802
rect 19156 13738 19208 13744
rect 19156 13524 19208 13530
rect 19156 13466 19208 13472
rect 19064 12844 19116 12850
rect 19064 12786 19116 12792
rect 19076 12442 19104 12786
rect 19064 12436 19116 12442
rect 19064 12378 19116 12384
rect 19168 10130 19196 13466
rect 19444 13326 19472 14214
rect 19996 14006 20024 14894
rect 19616 14000 19668 14006
rect 19616 13942 19668 13948
rect 19984 14000 20036 14006
rect 19984 13942 20036 13948
rect 19628 13870 19656 13942
rect 19616 13864 19668 13870
rect 19616 13806 19668 13812
rect 19984 13728 20036 13734
rect 19984 13670 20036 13676
rect 19580 13628 19876 13648
rect 19636 13626 19660 13628
rect 19716 13626 19740 13628
rect 19796 13626 19820 13628
rect 19658 13574 19660 13626
rect 19722 13574 19734 13626
rect 19796 13574 19798 13626
rect 19636 13572 19660 13574
rect 19716 13572 19740 13574
rect 19796 13572 19820 13574
rect 19580 13552 19876 13572
rect 19432 13320 19484 13326
rect 19432 13262 19484 13268
rect 19340 12980 19392 12986
rect 19340 12922 19392 12928
rect 19352 12374 19380 12922
rect 19444 12782 19472 13262
rect 19996 12986 20024 13670
rect 19984 12980 20036 12986
rect 19984 12922 20036 12928
rect 19432 12776 19484 12782
rect 19432 12718 19484 12724
rect 19984 12776 20036 12782
rect 19984 12718 20036 12724
rect 19892 12708 19944 12714
rect 19892 12650 19944 12656
rect 19432 12640 19484 12646
rect 19432 12582 19484 12588
rect 19340 12368 19392 12374
rect 19340 12310 19392 12316
rect 19248 12300 19300 12306
rect 19248 12242 19300 12248
rect 19260 11762 19288 12242
rect 19248 11756 19300 11762
rect 19248 11698 19300 11704
rect 19340 11212 19392 11218
rect 19340 11154 19392 11160
rect 19352 10470 19380 11154
rect 19444 10606 19472 12582
rect 19580 12540 19876 12560
rect 19636 12538 19660 12540
rect 19716 12538 19740 12540
rect 19796 12538 19820 12540
rect 19658 12486 19660 12538
rect 19722 12486 19734 12538
rect 19796 12486 19798 12538
rect 19636 12484 19660 12486
rect 19716 12484 19740 12486
rect 19796 12484 19820 12486
rect 19580 12464 19876 12484
rect 19904 12238 19932 12650
rect 19892 12232 19944 12238
rect 19892 12174 19944 12180
rect 19904 11898 19932 12174
rect 19892 11892 19944 11898
rect 19892 11834 19944 11840
rect 19904 11762 19932 11834
rect 19892 11756 19944 11762
rect 19892 11698 19944 11704
rect 19580 11452 19876 11472
rect 19636 11450 19660 11452
rect 19716 11450 19740 11452
rect 19796 11450 19820 11452
rect 19658 11398 19660 11450
rect 19722 11398 19734 11450
rect 19796 11398 19798 11450
rect 19636 11396 19660 11398
rect 19716 11396 19740 11398
rect 19796 11396 19820 11398
rect 19580 11376 19876 11396
rect 19432 10600 19484 10606
rect 19432 10542 19484 10548
rect 19340 10464 19392 10470
rect 19392 10424 19472 10452
rect 19340 10406 19392 10412
rect 19156 10124 19208 10130
rect 19156 10066 19208 10072
rect 19340 10124 19392 10130
rect 19340 10066 19392 10072
rect 19064 9512 19116 9518
rect 19064 9454 19116 9460
rect 19076 9110 19104 9454
rect 19352 9110 19380 10066
rect 19064 9104 19116 9110
rect 19064 9046 19116 9052
rect 19340 9104 19392 9110
rect 19340 9046 19392 9052
rect 19076 8430 19104 9046
rect 19444 8974 19472 10424
rect 19580 10364 19876 10384
rect 19636 10362 19660 10364
rect 19716 10362 19740 10364
rect 19796 10362 19820 10364
rect 19658 10310 19660 10362
rect 19722 10310 19734 10362
rect 19796 10310 19798 10362
rect 19636 10308 19660 10310
rect 19716 10308 19740 10310
rect 19796 10308 19820 10310
rect 19580 10288 19876 10308
rect 19904 10130 19932 11698
rect 19996 11218 20024 12718
rect 19984 11212 20036 11218
rect 19984 11154 20036 11160
rect 19984 10532 20036 10538
rect 19984 10474 20036 10480
rect 19892 10124 19944 10130
rect 19892 10066 19944 10072
rect 19580 9276 19876 9296
rect 19636 9274 19660 9276
rect 19716 9274 19740 9276
rect 19796 9274 19820 9276
rect 19658 9222 19660 9274
rect 19722 9222 19734 9274
rect 19796 9222 19798 9274
rect 19636 9220 19660 9222
rect 19716 9220 19740 9222
rect 19796 9220 19820 9222
rect 19580 9200 19876 9220
rect 19904 9042 19932 10066
rect 19996 9926 20024 10474
rect 19984 9920 20036 9926
rect 19984 9862 20036 9868
rect 19996 9586 20024 9862
rect 19984 9580 20036 9586
rect 19984 9522 20036 9528
rect 19800 9036 19852 9042
rect 19800 8978 19852 8984
rect 19892 9036 19944 9042
rect 19892 8978 19944 8984
rect 19432 8968 19484 8974
rect 19432 8910 19484 8916
rect 19812 8498 19840 8978
rect 19800 8492 19852 8498
rect 19800 8434 19852 8440
rect 19064 8424 19116 8430
rect 19064 8366 19116 8372
rect 19580 8188 19876 8208
rect 19636 8186 19660 8188
rect 19716 8186 19740 8188
rect 19796 8186 19820 8188
rect 19658 8134 19660 8186
rect 19722 8134 19734 8186
rect 19796 8134 19798 8186
rect 19636 8132 19660 8134
rect 19716 8132 19740 8134
rect 19796 8132 19820 8134
rect 19580 8112 19876 8132
rect 19156 8016 19208 8022
rect 19156 7958 19208 7964
rect 19064 7744 19116 7750
rect 19064 7686 19116 7692
rect 19076 7342 19104 7686
rect 19064 7336 19116 7342
rect 19064 7278 19116 7284
rect 19076 6254 19104 7278
rect 19168 6254 19196 7958
rect 19800 7948 19852 7954
rect 19984 7948 20036 7954
rect 19852 7908 19932 7936
rect 19800 7890 19852 7896
rect 19248 7812 19300 7818
rect 19248 7754 19300 7760
rect 19260 7410 19288 7754
rect 19248 7404 19300 7410
rect 19248 7346 19300 7352
rect 19248 7200 19300 7206
rect 19248 7142 19300 7148
rect 19260 6866 19288 7142
rect 19580 7100 19876 7120
rect 19636 7098 19660 7100
rect 19716 7098 19740 7100
rect 19796 7098 19820 7100
rect 19658 7046 19660 7098
rect 19722 7046 19734 7098
rect 19796 7046 19798 7098
rect 19636 7044 19660 7046
rect 19716 7044 19740 7046
rect 19796 7044 19820 7046
rect 19580 7024 19876 7044
rect 19432 6928 19484 6934
rect 19432 6870 19484 6876
rect 19248 6860 19300 6866
rect 19248 6802 19300 6808
rect 19444 6390 19472 6870
rect 19904 6866 19932 7908
rect 19984 7890 20036 7896
rect 19892 6860 19944 6866
rect 19892 6802 19944 6808
rect 19996 6798 20024 7890
rect 19984 6792 20036 6798
rect 19984 6734 20036 6740
rect 19432 6384 19484 6390
rect 19432 6326 19484 6332
rect 19064 6248 19116 6254
rect 19064 6190 19116 6196
rect 19156 6248 19208 6254
rect 19156 6190 19208 6196
rect 19064 6112 19116 6118
rect 19064 6054 19116 6060
rect 19076 5574 19104 6054
rect 19580 6012 19876 6032
rect 19636 6010 19660 6012
rect 19716 6010 19740 6012
rect 19796 6010 19820 6012
rect 19658 5958 19660 6010
rect 19722 5958 19734 6010
rect 19796 5958 19798 6010
rect 19636 5956 19660 5958
rect 19716 5956 19740 5958
rect 19796 5956 19820 5958
rect 19580 5936 19876 5956
rect 19064 5568 19116 5574
rect 19064 5510 19116 5516
rect 19984 5568 20036 5574
rect 19984 5510 20036 5516
rect 19580 4924 19876 4944
rect 19636 4922 19660 4924
rect 19716 4922 19740 4924
rect 19796 4922 19820 4924
rect 19658 4870 19660 4922
rect 19722 4870 19734 4922
rect 19796 4870 19798 4922
rect 19636 4868 19660 4870
rect 19716 4868 19740 4870
rect 19796 4868 19820 4870
rect 19580 4848 19876 4868
rect 19064 4820 19116 4826
rect 19064 4762 19116 4768
rect 19076 4078 19104 4762
rect 19246 4176 19302 4185
rect 19246 4111 19248 4120
rect 19300 4111 19302 4120
rect 19248 4082 19300 4088
rect 19996 4078 20024 5510
rect 19064 4072 19116 4078
rect 19064 4014 19116 4020
rect 19984 4072 20036 4078
rect 19984 4014 20036 4020
rect 19340 4004 19392 4010
rect 19340 3946 19392 3952
rect 18420 3936 18472 3942
rect 18420 3878 18472 3884
rect 18972 3936 19024 3942
rect 18972 3878 19024 3884
rect 18432 3534 18460 3878
rect 19062 3768 19118 3777
rect 19062 3703 19118 3712
rect 18236 3528 18288 3534
rect 18236 3470 18288 3476
rect 18420 3528 18472 3534
rect 18420 3470 18472 3476
rect 18248 3194 18276 3470
rect 19076 3466 19104 3703
rect 19064 3460 19116 3466
rect 19064 3402 19116 3408
rect 18328 3392 18380 3398
rect 18328 3334 18380 3340
rect 18236 3188 18288 3194
rect 18236 3130 18288 3136
rect 18144 2984 18196 2990
rect 18144 2926 18196 2932
rect 18340 2514 18368 3334
rect 19352 3058 19380 3946
rect 19580 3836 19876 3856
rect 19636 3834 19660 3836
rect 19716 3834 19740 3836
rect 19796 3834 19820 3836
rect 19658 3782 19660 3834
rect 19722 3782 19734 3834
rect 19796 3782 19798 3834
rect 19636 3780 19660 3782
rect 19716 3780 19740 3782
rect 19796 3780 19820 3782
rect 19580 3760 19876 3780
rect 19892 3528 19944 3534
rect 19892 3470 19944 3476
rect 19340 3052 19392 3058
rect 19340 2994 19392 3000
rect 18604 2984 18656 2990
rect 18604 2926 18656 2932
rect 19432 2984 19484 2990
rect 19432 2926 19484 2932
rect 18616 2650 18644 2926
rect 18880 2916 18932 2922
rect 18880 2858 18932 2864
rect 18604 2644 18656 2650
rect 18604 2586 18656 2592
rect 18892 2514 18920 2858
rect 18328 2508 18380 2514
rect 18328 2450 18380 2456
rect 18880 2508 18932 2514
rect 19444 2496 19472 2926
rect 19580 2748 19876 2768
rect 19636 2746 19660 2748
rect 19716 2746 19740 2748
rect 19796 2746 19820 2748
rect 19658 2694 19660 2746
rect 19722 2694 19734 2746
rect 19796 2694 19798 2746
rect 19636 2692 19660 2694
rect 19716 2692 19740 2694
rect 19796 2692 19820 2694
rect 19580 2672 19876 2692
rect 19524 2508 19576 2514
rect 19444 2468 19524 2496
rect 18880 2450 18932 2456
rect 19524 2450 19576 2456
rect 18052 2440 18104 2446
rect 18052 2382 18104 2388
rect 17316 2304 17368 2310
rect 17316 2246 17368 2252
rect 15304 2060 15424 2088
rect 15304 800 15332 2060
rect 17328 800 17356 2246
rect 19524 2100 19576 2106
rect 19524 2042 19576 2048
rect 19536 800 19564 2042
rect 19904 1970 19932 3470
rect 19996 2650 20024 4014
rect 19984 2644 20036 2650
rect 19984 2586 20036 2592
rect 20088 2106 20116 17682
rect 20168 17060 20220 17066
rect 20168 17002 20220 17008
rect 20180 16658 20208 17002
rect 20168 16652 20220 16658
rect 20168 16594 20220 16600
rect 20168 14340 20220 14346
rect 20168 14282 20220 14288
rect 20180 13870 20208 14282
rect 20168 13864 20220 13870
rect 20166 13832 20168 13841
rect 20220 13832 20222 13841
rect 20166 13767 20222 13776
rect 20168 11620 20220 11626
rect 20168 11562 20220 11568
rect 20180 11218 20208 11562
rect 20168 11212 20220 11218
rect 20168 11154 20220 11160
rect 20168 10600 20220 10606
rect 20168 10542 20220 10548
rect 20180 9722 20208 10542
rect 20168 9716 20220 9722
rect 20168 9658 20220 9664
rect 20168 9036 20220 9042
rect 20168 8978 20220 8984
rect 20180 6866 20208 8978
rect 20272 7426 20300 19858
rect 20364 14498 20392 23054
rect 20536 21888 20588 21894
rect 20536 21830 20588 21836
rect 20444 18216 20496 18222
rect 20444 18158 20496 18164
rect 20456 15162 20484 18158
rect 20548 15570 20576 21830
rect 20720 21616 20772 21622
rect 20720 21558 20772 21564
rect 20628 16992 20680 16998
rect 20628 16934 20680 16940
rect 20536 15564 20588 15570
rect 20536 15506 20588 15512
rect 20536 15360 20588 15366
rect 20536 15302 20588 15308
rect 20444 15156 20496 15162
rect 20444 15098 20496 15104
rect 20364 14470 20484 14498
rect 20352 11688 20404 11694
rect 20352 11630 20404 11636
rect 20364 11286 20392 11630
rect 20352 11280 20404 11286
rect 20352 11222 20404 11228
rect 20272 7398 20392 7426
rect 20260 7268 20312 7274
rect 20260 7210 20312 7216
rect 20272 7002 20300 7210
rect 20260 6996 20312 7002
rect 20260 6938 20312 6944
rect 20168 6860 20220 6866
rect 20168 6802 20220 6808
rect 20260 6792 20312 6798
rect 20260 6734 20312 6740
rect 20272 5914 20300 6734
rect 20364 6662 20392 7398
rect 20352 6656 20404 6662
rect 20352 6598 20404 6604
rect 20260 5908 20312 5914
rect 20260 5850 20312 5856
rect 20456 4146 20484 14470
rect 20548 13258 20576 15302
rect 20536 13252 20588 13258
rect 20536 13194 20588 13200
rect 20548 10674 20576 13194
rect 20640 12170 20668 16934
rect 20732 16794 20760 21558
rect 20916 19310 20944 35022
rect 22112 34746 22140 35022
rect 22284 35012 22336 35018
rect 22284 34954 22336 34960
rect 22100 34740 22152 34746
rect 22100 34682 22152 34688
rect 21640 34604 21692 34610
rect 21640 34546 21692 34552
rect 20996 34060 21048 34066
rect 20996 34002 21048 34008
rect 21008 29306 21036 34002
rect 21652 33862 21680 34546
rect 22296 34542 22324 34954
rect 23400 34678 23428 35090
rect 23388 34672 23440 34678
rect 23388 34614 23440 34620
rect 24136 34542 24164 35430
rect 22284 34536 22336 34542
rect 22284 34478 22336 34484
rect 22744 34536 22796 34542
rect 22744 34478 22796 34484
rect 24124 34536 24176 34542
rect 24124 34478 24176 34484
rect 21824 34468 21876 34474
rect 21824 34410 21876 34416
rect 21640 33856 21692 33862
rect 21640 33798 21692 33804
rect 21652 33590 21680 33798
rect 21640 33584 21692 33590
rect 21640 33526 21692 33532
rect 21088 33516 21140 33522
rect 21088 33458 21140 33464
rect 21100 32434 21128 33458
rect 21836 33454 21864 34410
rect 22284 33992 22336 33998
rect 22284 33934 22336 33940
rect 22296 33522 22324 33934
rect 22284 33516 22336 33522
rect 22284 33458 22336 33464
rect 21824 33448 21876 33454
rect 21824 33390 21876 33396
rect 21180 33380 21232 33386
rect 21180 33322 21232 33328
rect 21192 32978 21220 33322
rect 21180 32972 21232 32978
rect 21180 32914 21232 32920
rect 22652 32564 22704 32570
rect 22652 32506 22704 32512
rect 21088 32428 21140 32434
rect 21088 32370 21140 32376
rect 21100 31822 21128 32370
rect 22664 31890 22692 32506
rect 21456 31884 21508 31890
rect 21456 31826 21508 31832
rect 22652 31884 22704 31890
rect 22652 31826 22704 31832
rect 21088 31816 21140 31822
rect 21088 31758 21140 31764
rect 21272 30116 21324 30122
rect 21272 30058 21324 30064
rect 21284 29714 21312 30058
rect 21272 29708 21324 29714
rect 21272 29650 21324 29656
rect 20996 29300 21048 29306
rect 20996 29242 21048 29248
rect 21364 29300 21416 29306
rect 21364 29242 21416 29248
rect 21088 29164 21140 29170
rect 21088 29106 21140 29112
rect 20996 28620 21048 28626
rect 20996 28562 21048 28568
rect 21008 27946 21036 28562
rect 20996 27940 21048 27946
rect 20996 27882 21048 27888
rect 21008 27674 21036 27882
rect 20996 27668 21048 27674
rect 20996 27610 21048 27616
rect 21100 27130 21128 29106
rect 21088 27124 21140 27130
rect 21088 27066 21140 27072
rect 21376 25906 21404 29242
rect 21468 28132 21496 31826
rect 21640 31272 21692 31278
rect 21640 31214 21692 31220
rect 21548 31136 21600 31142
rect 21548 31078 21600 31084
rect 21560 30802 21588 31078
rect 21548 30796 21600 30802
rect 21548 30738 21600 30744
rect 21652 30258 21680 31214
rect 22560 31204 22612 31210
rect 22560 31146 22612 31152
rect 22376 31136 22428 31142
rect 22376 31078 22428 31084
rect 22572 31090 22600 31146
rect 21640 30252 21692 30258
rect 21640 30194 21692 30200
rect 22008 30184 22060 30190
rect 22008 30126 22060 30132
rect 21732 30048 21784 30054
rect 21732 29990 21784 29996
rect 21744 29714 21772 29990
rect 22020 29782 22048 30126
rect 22008 29776 22060 29782
rect 22008 29718 22060 29724
rect 21732 29708 21784 29714
rect 21732 29650 21784 29656
rect 21548 29096 21600 29102
rect 21548 29038 21600 29044
rect 22100 29096 22152 29102
rect 22100 29038 22152 29044
rect 21560 28626 21588 29038
rect 22112 28626 22140 29038
rect 21548 28620 21600 28626
rect 21548 28562 21600 28568
rect 22100 28620 22152 28626
rect 22100 28562 22152 28568
rect 22284 28484 22336 28490
rect 22284 28426 22336 28432
rect 21468 28104 21588 28132
rect 21364 25900 21416 25906
rect 21364 25842 21416 25848
rect 21180 25832 21232 25838
rect 21180 25774 21232 25780
rect 21088 24812 21140 24818
rect 21088 24754 21140 24760
rect 21100 23662 21128 24754
rect 21192 24138 21220 25774
rect 21180 24132 21232 24138
rect 21180 24074 21232 24080
rect 21088 23656 21140 23662
rect 21088 23598 21140 23604
rect 20996 23588 21048 23594
rect 20996 23530 21048 23536
rect 21008 23322 21036 23530
rect 21364 23520 21416 23526
rect 21364 23462 21416 23468
rect 20996 23316 21048 23322
rect 20996 23258 21048 23264
rect 21008 23186 21036 23258
rect 20996 23180 21048 23186
rect 20996 23122 21048 23128
rect 21180 22772 21232 22778
rect 21180 22714 21232 22720
rect 21088 22568 21140 22574
rect 21088 22510 21140 22516
rect 21100 22166 21128 22510
rect 21088 22160 21140 22166
rect 21088 22102 21140 22108
rect 20996 22092 21048 22098
rect 20996 22034 21048 22040
rect 20904 19304 20956 19310
rect 20904 19246 20956 19252
rect 20720 16788 20772 16794
rect 20720 16730 20772 16736
rect 20720 16584 20772 16590
rect 20720 16526 20772 16532
rect 20732 16046 20760 16526
rect 20720 16040 20772 16046
rect 20720 15982 20772 15988
rect 20812 15972 20864 15978
rect 20812 15914 20864 15920
rect 20824 15706 20852 15914
rect 20812 15700 20864 15706
rect 20812 15642 20864 15648
rect 20812 15496 20864 15502
rect 20812 15438 20864 15444
rect 20720 15428 20772 15434
rect 20720 15370 20772 15376
rect 20732 14958 20760 15370
rect 20720 14952 20772 14958
rect 20720 14894 20772 14900
rect 20732 12986 20760 14894
rect 20824 14822 20852 15438
rect 20904 14884 20956 14890
rect 20904 14826 20956 14832
rect 20812 14816 20864 14822
rect 20812 14758 20864 14764
rect 20824 13870 20852 14758
rect 20916 14074 20944 14826
rect 20904 14068 20956 14074
rect 20904 14010 20956 14016
rect 20812 13864 20864 13870
rect 20812 13806 20864 13812
rect 20720 12980 20772 12986
rect 20720 12922 20772 12928
rect 20824 12306 20852 13806
rect 20916 13802 20944 14010
rect 20904 13796 20956 13802
rect 20904 13738 20956 13744
rect 21008 13297 21036 22034
rect 21088 21004 21140 21010
rect 21088 20946 21140 20952
rect 21100 20534 21128 20946
rect 21088 20528 21140 20534
rect 21088 20470 21140 20476
rect 21088 19304 21140 19310
rect 21088 19246 21140 19252
rect 21100 18902 21128 19246
rect 21088 18896 21140 18902
rect 21088 18838 21140 18844
rect 21192 18816 21220 22714
rect 21376 22642 21404 23462
rect 21364 22636 21416 22642
rect 21364 22578 21416 22584
rect 21456 22568 21508 22574
rect 21456 22510 21508 22516
rect 21364 21888 21416 21894
rect 21364 21830 21416 21836
rect 21272 21548 21324 21554
rect 21272 21490 21324 21496
rect 21284 20398 21312 21490
rect 21376 20398 21404 21830
rect 21468 21486 21496 22510
rect 21560 22098 21588 28104
rect 22296 27538 22324 28426
rect 21640 27532 21692 27538
rect 21640 27474 21692 27480
rect 22284 27532 22336 27538
rect 22284 27474 22336 27480
rect 21652 24274 21680 27474
rect 21916 26920 21968 26926
rect 21916 26862 21968 26868
rect 22284 26920 22336 26926
rect 22284 26862 22336 26868
rect 21928 26450 21956 26862
rect 21916 26444 21968 26450
rect 21916 26386 21968 26392
rect 22100 26376 22152 26382
rect 22100 26318 22152 26324
rect 22112 25906 22140 26318
rect 22100 25900 22152 25906
rect 22100 25842 22152 25848
rect 22296 25362 22324 26862
rect 21732 25356 21784 25362
rect 21732 25298 21784 25304
rect 22284 25356 22336 25362
rect 22284 25298 22336 25304
rect 21744 24274 21772 25298
rect 22008 25288 22060 25294
rect 22008 25230 22060 25236
rect 22020 24410 22048 25230
rect 22192 24880 22244 24886
rect 22296 24868 22324 25298
rect 22244 24840 22324 24868
rect 22192 24822 22244 24828
rect 22192 24744 22244 24750
rect 22192 24686 22244 24692
rect 22008 24404 22060 24410
rect 22008 24346 22060 24352
rect 22100 24404 22152 24410
rect 22100 24346 22152 24352
rect 21640 24268 21692 24274
rect 21640 24210 21692 24216
rect 21732 24268 21784 24274
rect 21732 24210 21784 24216
rect 21652 24138 21680 24210
rect 21640 24132 21692 24138
rect 21640 24074 21692 24080
rect 21652 23798 21680 24074
rect 21640 23792 21692 23798
rect 21640 23734 21692 23740
rect 21640 23656 21692 23662
rect 21640 23598 21692 23604
rect 21652 23254 21680 23598
rect 21744 23526 21772 24210
rect 21824 23792 21876 23798
rect 21824 23734 21876 23740
rect 21732 23520 21784 23526
rect 21732 23462 21784 23468
rect 21640 23248 21692 23254
rect 21640 23190 21692 23196
rect 21836 23050 21864 23734
rect 22020 23254 22048 24346
rect 22008 23248 22060 23254
rect 22008 23190 22060 23196
rect 21916 23112 21968 23118
rect 21916 23054 21968 23060
rect 22008 23112 22060 23118
rect 22008 23054 22060 23060
rect 21824 23044 21876 23050
rect 21824 22986 21876 22992
rect 21824 22704 21876 22710
rect 21824 22646 21876 22652
rect 21836 22098 21864 22646
rect 21548 22092 21600 22098
rect 21548 22034 21600 22040
rect 21824 22092 21876 22098
rect 21824 22034 21876 22040
rect 21548 21888 21600 21894
rect 21548 21830 21600 21836
rect 21560 21486 21588 21830
rect 21732 21616 21784 21622
rect 21732 21558 21784 21564
rect 21456 21480 21508 21486
rect 21456 21422 21508 21428
rect 21548 21480 21600 21486
rect 21548 21422 21600 21428
rect 21468 21146 21496 21422
rect 21456 21140 21508 21146
rect 21456 21082 21508 21088
rect 21468 20806 21496 21082
rect 21548 20936 21600 20942
rect 21548 20878 21600 20884
rect 21456 20800 21508 20806
rect 21456 20742 21508 20748
rect 21560 20466 21588 20878
rect 21548 20460 21600 20466
rect 21548 20402 21600 20408
rect 21272 20392 21324 20398
rect 21272 20334 21324 20340
rect 21364 20392 21416 20398
rect 21364 20334 21416 20340
rect 21284 19378 21312 20334
rect 21272 19372 21324 19378
rect 21272 19314 21324 19320
rect 21376 18902 21404 20334
rect 21640 19916 21692 19922
rect 21640 19858 21692 19864
rect 21548 19372 21600 19378
rect 21548 19314 21600 19320
rect 21364 18896 21416 18902
rect 21364 18838 21416 18844
rect 21192 18788 21312 18816
rect 21180 18692 21232 18698
rect 21180 18634 21232 18640
rect 21192 18358 21220 18634
rect 21180 18352 21232 18358
rect 21180 18294 21232 18300
rect 21088 17672 21140 17678
rect 21088 17614 21140 17620
rect 20994 13288 21050 13297
rect 20994 13223 21050 13232
rect 20720 12300 20772 12306
rect 20720 12242 20772 12248
rect 20812 12300 20864 12306
rect 20812 12242 20864 12248
rect 20732 12186 20760 12242
rect 20628 12164 20680 12170
rect 20732 12158 21036 12186
rect 20628 12106 20680 12112
rect 20640 11354 20668 12106
rect 21008 11694 21036 12158
rect 20996 11688 21048 11694
rect 20996 11630 21048 11636
rect 20628 11348 20680 11354
rect 20628 11290 20680 11296
rect 20536 10668 20588 10674
rect 20536 10610 20588 10616
rect 21008 9382 21036 11630
rect 20996 9376 21048 9382
rect 20996 9318 21048 9324
rect 21008 8430 21036 9318
rect 20996 8424 21048 8430
rect 20996 8366 21048 8372
rect 21100 6934 21128 17614
rect 21180 16448 21232 16454
rect 21180 16390 21232 16396
rect 21192 14958 21220 16390
rect 21284 16114 21312 18788
rect 21376 17202 21404 18838
rect 21364 17196 21416 17202
rect 21364 17138 21416 17144
rect 21454 16552 21510 16561
rect 21454 16487 21456 16496
rect 21508 16487 21510 16496
rect 21456 16458 21508 16464
rect 21272 16108 21324 16114
rect 21272 16050 21324 16056
rect 21180 14952 21232 14958
rect 21180 14894 21232 14900
rect 21456 14952 21508 14958
rect 21456 14894 21508 14900
rect 21272 14884 21324 14890
rect 21272 14826 21324 14832
rect 21180 14408 21232 14414
rect 21180 14350 21232 14356
rect 21192 13938 21220 14350
rect 21180 13932 21232 13938
rect 21180 13874 21232 13880
rect 21284 13870 21312 14826
rect 21364 14272 21416 14278
rect 21364 14214 21416 14220
rect 21272 13864 21324 13870
rect 21272 13806 21324 13812
rect 21284 13530 21312 13806
rect 21272 13524 21324 13530
rect 21272 13466 21324 13472
rect 21376 13394 21404 14214
rect 21468 13734 21496 14894
rect 21456 13728 21508 13734
rect 21456 13670 21508 13676
rect 21468 13394 21496 13670
rect 21364 13388 21416 13394
rect 21364 13330 21416 13336
rect 21456 13388 21508 13394
rect 21456 13330 21508 13336
rect 21272 12776 21324 12782
rect 21272 12718 21324 12724
rect 21284 9994 21312 12718
rect 21376 12374 21404 13330
rect 21560 13190 21588 19314
rect 21652 18630 21680 19858
rect 21640 18624 21692 18630
rect 21640 18566 21692 18572
rect 21744 17746 21772 21558
rect 21836 21010 21864 22034
rect 21928 21554 21956 23054
rect 22020 22166 22048 23054
rect 22008 22160 22060 22166
rect 22008 22102 22060 22108
rect 22020 21622 22048 22102
rect 22008 21616 22060 21622
rect 22008 21558 22060 21564
rect 21916 21548 21968 21554
rect 21916 21490 21968 21496
rect 22112 21146 22140 24346
rect 22100 21140 22152 21146
rect 22100 21082 22152 21088
rect 21824 21004 21876 21010
rect 21824 20946 21876 20952
rect 21836 19922 21864 20946
rect 22008 20868 22060 20874
rect 22008 20810 22060 20816
rect 22020 20534 22048 20810
rect 22008 20528 22060 20534
rect 22008 20470 22060 20476
rect 22020 20058 22048 20470
rect 22204 20262 22232 24686
rect 22296 24682 22324 24840
rect 22284 24676 22336 24682
rect 22284 24618 22336 24624
rect 22284 21004 22336 21010
rect 22284 20946 22336 20952
rect 22192 20256 22244 20262
rect 22192 20198 22244 20204
rect 22008 20052 22060 20058
rect 22008 19994 22060 20000
rect 21824 19916 21876 19922
rect 21824 19858 21876 19864
rect 21824 19168 21876 19174
rect 21824 19110 21876 19116
rect 21836 18902 21864 19110
rect 21824 18896 21876 18902
rect 21824 18838 21876 18844
rect 22008 18896 22060 18902
rect 22008 18838 22060 18844
rect 22020 18154 22048 18838
rect 22296 18766 22324 20946
rect 22100 18760 22152 18766
rect 22100 18702 22152 18708
rect 22284 18760 22336 18766
rect 22284 18702 22336 18708
rect 22008 18148 22060 18154
rect 22008 18090 22060 18096
rect 22112 18086 22140 18702
rect 22284 18420 22336 18426
rect 22284 18362 22336 18368
rect 22192 18352 22244 18358
rect 22192 18294 22244 18300
rect 22100 18080 22152 18086
rect 22100 18022 22152 18028
rect 21732 17740 21784 17746
rect 21732 17682 21784 17688
rect 21640 17128 21692 17134
rect 21744 17116 21772 17682
rect 22100 17536 22152 17542
rect 22100 17478 22152 17484
rect 21692 17088 21772 17116
rect 22008 17128 22060 17134
rect 21640 17070 21692 17076
rect 22008 17070 22060 17076
rect 21652 16658 21680 17070
rect 22020 16794 22048 17070
rect 22008 16788 22060 16794
rect 22008 16730 22060 16736
rect 22020 16658 22048 16730
rect 21640 16652 21692 16658
rect 21640 16594 21692 16600
rect 22008 16652 22060 16658
rect 22008 16594 22060 16600
rect 22112 16046 22140 17478
rect 22204 17134 22232 18294
rect 22192 17128 22244 17134
rect 22192 17070 22244 17076
rect 22100 16040 22152 16046
rect 22100 15982 22152 15988
rect 22100 15904 22152 15910
rect 22100 15846 22152 15852
rect 22112 15570 22140 15846
rect 22204 15638 22232 17070
rect 22296 16046 22324 18362
rect 22284 16040 22336 16046
rect 22284 15982 22336 15988
rect 22192 15632 22244 15638
rect 22192 15574 22244 15580
rect 22296 15570 22324 15982
rect 22100 15564 22152 15570
rect 22100 15506 22152 15512
rect 22284 15564 22336 15570
rect 22284 15506 22336 15512
rect 22008 14612 22060 14618
rect 22008 14554 22060 14560
rect 22020 13190 22048 14554
rect 22190 13968 22246 13977
rect 22190 13903 22246 13912
rect 22204 13870 22232 13903
rect 22192 13864 22244 13870
rect 22192 13806 22244 13812
rect 22192 13728 22244 13734
rect 22192 13670 22244 13676
rect 21548 13184 21600 13190
rect 21548 13126 21600 13132
rect 22008 13184 22060 13190
rect 22008 13126 22060 13132
rect 21548 12776 21600 12782
rect 21548 12718 21600 12724
rect 21364 12368 21416 12374
rect 21364 12310 21416 12316
rect 21560 12170 21588 12718
rect 21364 12164 21416 12170
rect 21364 12106 21416 12112
rect 21548 12164 21600 12170
rect 21548 12106 21600 12112
rect 21376 11694 21404 12106
rect 21640 12096 21692 12102
rect 21640 12038 21692 12044
rect 21652 11898 21680 12038
rect 21640 11892 21692 11898
rect 21640 11834 21692 11840
rect 21364 11688 21416 11694
rect 21364 11630 21416 11636
rect 22008 11552 22060 11558
rect 22008 11494 22060 11500
rect 21548 11212 21600 11218
rect 21548 11154 21600 11160
rect 21916 11212 21968 11218
rect 21916 11154 21968 11160
rect 21456 10668 21508 10674
rect 21456 10610 21508 10616
rect 21468 10062 21496 10610
rect 21560 10538 21588 11154
rect 21640 11144 21692 11150
rect 21640 11086 21692 11092
rect 21652 10606 21680 11086
rect 21928 10713 21956 11154
rect 22020 11082 22048 11494
rect 22008 11076 22060 11082
rect 22008 11018 22060 11024
rect 21914 10704 21970 10713
rect 21914 10639 21970 10648
rect 21640 10600 21692 10606
rect 21640 10542 21692 10548
rect 21548 10532 21600 10538
rect 21548 10474 21600 10480
rect 22008 10464 22060 10470
rect 22204 10452 22232 13670
rect 22284 12300 22336 12306
rect 22284 12242 22336 12248
rect 22296 11558 22324 12242
rect 22284 11552 22336 11558
rect 22284 11494 22336 11500
rect 22284 10464 22336 10470
rect 22204 10424 22284 10452
rect 22008 10406 22060 10412
rect 22284 10406 22336 10412
rect 21548 10124 21600 10130
rect 21548 10066 21600 10072
rect 21916 10124 21968 10130
rect 21916 10066 21968 10072
rect 21456 10056 21508 10062
rect 21456 9998 21508 10004
rect 21272 9988 21324 9994
rect 21272 9930 21324 9936
rect 21284 7886 21312 9930
rect 21468 9586 21496 9998
rect 21456 9580 21508 9586
rect 21456 9522 21508 9528
rect 21364 9172 21416 9178
rect 21364 9114 21416 9120
rect 21376 8974 21404 9114
rect 21364 8968 21416 8974
rect 21364 8910 21416 8916
rect 21456 8968 21508 8974
rect 21456 8910 21508 8916
rect 21272 7880 21324 7886
rect 21272 7822 21324 7828
rect 21376 7562 21404 8910
rect 21468 8634 21496 8910
rect 21456 8628 21508 8634
rect 21456 8570 21508 8576
rect 21560 8498 21588 10066
rect 21640 9512 21692 9518
rect 21640 9454 21692 9460
rect 21824 9512 21876 9518
rect 21824 9454 21876 9460
rect 21548 8492 21600 8498
rect 21548 8434 21600 8440
rect 21456 8356 21508 8362
rect 21456 8298 21508 8304
rect 21468 7886 21496 8298
rect 21456 7880 21508 7886
rect 21456 7822 21508 7828
rect 21376 7534 21588 7562
rect 21560 7342 21588 7534
rect 21548 7336 21600 7342
rect 21548 7278 21600 7284
rect 21088 6928 21140 6934
rect 21088 6870 21140 6876
rect 20628 6860 20680 6866
rect 20628 6802 20680 6808
rect 20640 6458 20668 6802
rect 21456 6792 21508 6798
rect 21456 6734 21508 6740
rect 20628 6452 20680 6458
rect 20628 6394 20680 6400
rect 20812 6384 20864 6390
rect 20812 6326 20864 6332
rect 20824 6254 20852 6326
rect 20720 6248 20772 6254
rect 20720 6190 20772 6196
rect 20812 6248 20864 6254
rect 20812 6190 20864 6196
rect 20732 4554 20760 6190
rect 20824 4690 20852 6190
rect 21468 4690 21496 6734
rect 20812 4684 20864 4690
rect 20812 4626 20864 4632
rect 21456 4684 21508 4690
rect 21456 4626 21508 4632
rect 21560 4622 21588 7278
rect 21652 6254 21680 9454
rect 21836 9382 21864 9454
rect 21824 9376 21876 9382
rect 21824 9318 21876 9324
rect 21928 8430 21956 10066
rect 22020 10062 22048 10406
rect 22008 10056 22060 10062
rect 22008 9998 22060 10004
rect 22020 9654 22048 9998
rect 22008 9648 22060 9654
rect 22008 9590 22060 9596
rect 22192 9036 22244 9042
rect 22192 8978 22244 8984
rect 22100 8900 22152 8906
rect 22100 8842 22152 8848
rect 21916 8424 21968 8430
rect 21968 8384 22048 8412
rect 21916 8366 21968 8372
rect 22020 8090 22048 8384
rect 22008 8084 22060 8090
rect 22008 8026 22060 8032
rect 22112 7954 22140 8842
rect 22204 8498 22232 8978
rect 22192 8492 22244 8498
rect 22192 8434 22244 8440
rect 22100 7948 22152 7954
rect 22100 7890 22152 7896
rect 21824 7744 21876 7750
rect 22296 7698 22324 10406
rect 21824 7686 21876 7692
rect 21836 7342 21864 7686
rect 22204 7670 22324 7698
rect 21824 7336 21876 7342
rect 21824 7278 21876 7284
rect 21732 7200 21784 7206
rect 21732 7142 21784 7148
rect 22008 7200 22060 7206
rect 22008 7142 22060 7148
rect 21640 6248 21692 6254
rect 21640 6190 21692 6196
rect 21652 5914 21680 6190
rect 21640 5908 21692 5914
rect 21640 5850 21692 5856
rect 21744 5778 21772 7142
rect 22020 6866 22048 7142
rect 21916 6860 21968 6866
rect 21916 6802 21968 6808
rect 22008 6860 22060 6866
rect 22008 6802 22060 6808
rect 21928 6662 21956 6802
rect 22204 6662 22232 7670
rect 22388 7562 22416 31078
rect 22572 31062 22692 31090
rect 22664 30598 22692 31062
rect 22652 30592 22704 30598
rect 22652 30534 22704 30540
rect 22664 30190 22692 30534
rect 22652 30184 22704 30190
rect 22652 30126 22704 30132
rect 22664 29646 22692 30126
rect 22652 29640 22704 29646
rect 22652 29582 22704 29588
rect 22560 28008 22612 28014
rect 22560 27950 22612 27956
rect 22468 27532 22520 27538
rect 22468 27474 22520 27480
rect 22480 26042 22508 27474
rect 22468 26036 22520 26042
rect 22468 25978 22520 25984
rect 22572 25702 22600 27950
rect 22560 25696 22612 25702
rect 22560 25638 22612 25644
rect 22756 24342 22784 34478
rect 24228 34066 24256 36790
rect 24504 36786 24532 40200
rect 25504 38276 25556 38282
rect 25504 38218 25556 38224
rect 25516 37874 25544 38218
rect 26712 37874 26740 40200
rect 26792 38208 26844 38214
rect 26792 38150 26844 38156
rect 26804 38010 26832 38150
rect 26792 38004 26844 38010
rect 26792 37946 26844 37952
rect 25504 37868 25556 37874
rect 25504 37810 25556 37816
rect 26700 37868 26752 37874
rect 26700 37810 26752 37816
rect 26424 37800 26476 37806
rect 26424 37742 26476 37748
rect 24584 37664 24636 37670
rect 24584 37606 24636 37612
rect 24596 36854 24624 37606
rect 25320 37460 25372 37466
rect 25320 37402 25372 37408
rect 24584 36848 24636 36854
rect 24584 36790 24636 36796
rect 24492 36780 24544 36786
rect 24492 36722 24544 36728
rect 25332 36718 25360 37402
rect 26436 37330 26464 37742
rect 26792 37664 26844 37670
rect 26792 37606 26844 37612
rect 26804 37330 26832 37606
rect 28736 37466 28764 40200
rect 29828 38548 29880 38554
rect 29828 38490 29880 38496
rect 29840 37806 29868 38490
rect 30472 38344 30524 38350
rect 30472 38286 30524 38292
rect 30484 37806 30512 38286
rect 30656 38276 30708 38282
rect 30656 38218 30708 38224
rect 29828 37800 29880 37806
rect 29828 37742 29880 37748
rect 30472 37800 30524 37806
rect 30472 37742 30524 37748
rect 28724 37460 28776 37466
rect 28724 37402 28776 37408
rect 25504 37324 25556 37330
rect 25504 37266 25556 37272
rect 26240 37324 26292 37330
rect 26240 37266 26292 37272
rect 26424 37324 26476 37330
rect 26424 37266 26476 37272
rect 26792 37324 26844 37330
rect 26792 37266 26844 37272
rect 25516 36786 25544 37266
rect 25504 36780 25556 36786
rect 25504 36722 25556 36728
rect 24676 36712 24728 36718
rect 24676 36654 24728 36660
rect 25320 36712 25372 36718
rect 25320 36654 25372 36660
rect 24400 36168 24452 36174
rect 24400 36110 24452 36116
rect 24412 35766 24440 36110
rect 24400 35760 24452 35766
rect 24400 35702 24452 35708
rect 24688 35290 24716 36654
rect 25228 36576 25280 36582
rect 25228 36518 25280 36524
rect 25136 35760 25188 35766
rect 25136 35702 25188 35708
rect 24768 35692 24820 35698
rect 24768 35634 24820 35640
rect 24676 35284 24728 35290
rect 24676 35226 24728 35232
rect 24492 34944 24544 34950
rect 24492 34886 24544 34892
rect 24504 34610 24532 34886
rect 24688 34746 24716 35226
rect 24780 35154 24808 35634
rect 25148 35562 25176 35702
rect 25240 35630 25268 36518
rect 25516 36378 25544 36722
rect 25504 36372 25556 36378
rect 25504 36314 25556 36320
rect 25516 35630 25544 36314
rect 26252 35630 26280 37266
rect 26436 36786 26464 37266
rect 28908 37256 28960 37262
rect 28908 37198 28960 37204
rect 27712 37120 27764 37126
rect 27712 37062 27764 37068
rect 27724 36786 27752 37062
rect 28920 36786 28948 37198
rect 30012 37120 30064 37126
rect 30012 37062 30064 37068
rect 30024 36786 30052 37062
rect 26424 36780 26476 36786
rect 26424 36722 26476 36728
rect 27712 36780 27764 36786
rect 27712 36722 27764 36728
rect 28908 36780 28960 36786
rect 28908 36722 28960 36728
rect 30012 36780 30064 36786
rect 30012 36722 30064 36728
rect 26608 36712 26660 36718
rect 26608 36654 26660 36660
rect 26332 36168 26384 36174
rect 26332 36110 26384 36116
rect 25228 35624 25280 35630
rect 25228 35566 25280 35572
rect 25504 35624 25556 35630
rect 25504 35566 25556 35572
rect 26240 35624 26292 35630
rect 26240 35566 26292 35572
rect 25136 35556 25188 35562
rect 25136 35498 25188 35504
rect 24768 35148 24820 35154
rect 24768 35090 24820 35096
rect 24676 34740 24728 34746
rect 24676 34682 24728 34688
rect 24492 34604 24544 34610
rect 24492 34546 24544 34552
rect 24216 34060 24268 34066
rect 24216 34002 24268 34008
rect 25228 34060 25280 34066
rect 25228 34002 25280 34008
rect 24124 33992 24176 33998
rect 24124 33934 24176 33940
rect 25136 33992 25188 33998
rect 25136 33934 25188 33940
rect 23572 33856 23624 33862
rect 23572 33798 23624 33804
rect 23204 33516 23256 33522
rect 23204 33458 23256 33464
rect 23216 32910 23244 33458
rect 23204 32904 23256 32910
rect 23204 32846 23256 32852
rect 23216 32434 23244 32846
rect 23204 32428 23256 32434
rect 23204 32370 23256 32376
rect 23480 31816 23532 31822
rect 23480 31758 23532 31764
rect 23492 31414 23520 31758
rect 23584 31414 23612 33798
rect 24136 33658 24164 33934
rect 24400 33856 24452 33862
rect 24400 33798 24452 33804
rect 24860 33856 24912 33862
rect 24860 33798 24912 33804
rect 24124 33652 24176 33658
rect 24124 33594 24176 33600
rect 23756 33312 23808 33318
rect 23756 33254 23808 33260
rect 23480 31408 23532 31414
rect 23480 31350 23532 31356
rect 23572 31408 23624 31414
rect 23572 31350 23624 31356
rect 23572 31272 23624 31278
rect 23768 31260 23796 33254
rect 24412 32978 24440 33798
rect 24492 33652 24544 33658
rect 24492 33594 24544 33600
rect 24504 33454 24532 33594
rect 24872 33522 24900 33798
rect 24860 33516 24912 33522
rect 24860 33458 24912 33464
rect 24492 33448 24544 33454
rect 24492 33390 24544 33396
rect 24400 32972 24452 32978
rect 24400 32914 24452 32920
rect 24400 32224 24452 32230
rect 24400 32166 24452 32172
rect 24412 31822 24440 32166
rect 24400 31816 24452 31822
rect 24400 31758 24452 31764
rect 24032 31680 24084 31686
rect 24032 31622 24084 31628
rect 24044 31278 24072 31622
rect 24216 31408 24268 31414
rect 24216 31350 24268 31356
rect 23624 31232 23796 31260
rect 24032 31272 24084 31278
rect 23572 31214 23624 31220
rect 24032 31214 24084 31220
rect 23020 30728 23072 30734
rect 23020 30670 23072 30676
rect 22836 29232 22888 29238
rect 22836 29174 22888 29180
rect 22848 28082 22876 29174
rect 23032 29034 23060 30670
rect 23204 30184 23256 30190
rect 23204 30126 23256 30132
rect 23020 29028 23072 29034
rect 23020 28970 23072 28976
rect 22836 28076 22888 28082
rect 22836 28018 22888 28024
rect 23216 27470 23244 30126
rect 23296 30116 23348 30122
rect 23296 30058 23348 30064
rect 23308 28626 23336 30058
rect 23388 29708 23440 29714
rect 23388 29650 23440 29656
rect 23296 28620 23348 28626
rect 23296 28562 23348 28568
rect 23020 27464 23072 27470
rect 23020 27406 23072 27412
rect 23204 27464 23256 27470
rect 23204 27406 23256 27412
rect 22928 27396 22980 27402
rect 22928 27338 22980 27344
rect 22836 27328 22888 27334
rect 22836 27270 22888 27276
rect 22848 26926 22876 27270
rect 22940 27130 22968 27338
rect 22928 27124 22980 27130
rect 22928 27066 22980 27072
rect 22836 26920 22888 26926
rect 22836 26862 22888 26868
rect 22848 26450 22876 26862
rect 22836 26444 22888 26450
rect 22836 26386 22888 26392
rect 22744 24336 22796 24342
rect 22744 24278 22796 24284
rect 22848 24070 22876 26386
rect 22928 24744 22980 24750
rect 22928 24686 22980 24692
rect 22836 24064 22888 24070
rect 22836 24006 22888 24012
rect 22940 23866 22968 24686
rect 23032 24342 23060 27406
rect 23020 24336 23072 24342
rect 23020 24278 23072 24284
rect 23308 24274 23336 28562
rect 23296 24268 23348 24274
rect 23296 24210 23348 24216
rect 23204 24064 23256 24070
rect 23204 24006 23256 24012
rect 22928 23860 22980 23866
rect 22928 23802 22980 23808
rect 22940 23186 22968 23802
rect 23020 23656 23072 23662
rect 23020 23598 23072 23604
rect 23032 23322 23060 23598
rect 23216 23322 23244 24006
rect 23020 23316 23072 23322
rect 23020 23258 23072 23264
rect 23204 23316 23256 23322
rect 23204 23258 23256 23264
rect 22928 23180 22980 23186
rect 22928 23122 22980 23128
rect 23032 22574 23060 23258
rect 23308 23050 23336 24210
rect 23400 23730 23428 29650
rect 23480 27328 23532 27334
rect 23480 27270 23532 27276
rect 23492 26450 23520 27270
rect 23480 26444 23532 26450
rect 23480 26386 23532 26392
rect 23584 26314 23612 31214
rect 23664 30796 23716 30802
rect 23664 30738 23716 30744
rect 23676 30054 23704 30738
rect 23940 30184 23992 30190
rect 23940 30126 23992 30132
rect 23664 30048 23716 30054
rect 23664 29990 23716 29996
rect 23676 29578 23704 29990
rect 23664 29572 23716 29578
rect 23664 29514 23716 29520
rect 23676 29102 23704 29514
rect 23664 29096 23716 29102
rect 23664 29038 23716 29044
rect 23572 26308 23624 26314
rect 23572 26250 23624 26256
rect 23480 26240 23532 26246
rect 23480 26182 23532 26188
rect 23492 25498 23520 26182
rect 23676 25838 23704 29038
rect 23848 28620 23900 28626
rect 23848 28562 23900 28568
rect 23756 28484 23808 28490
rect 23756 28426 23808 28432
rect 23768 28014 23796 28426
rect 23756 28008 23808 28014
rect 23756 27950 23808 27956
rect 23860 27606 23888 28562
rect 23952 28098 23980 30126
rect 24044 29714 24072 31214
rect 24228 30802 24256 31350
rect 24216 30796 24268 30802
rect 24216 30738 24268 30744
rect 24032 29708 24084 29714
rect 24032 29650 24084 29656
rect 24216 29708 24268 29714
rect 24216 29650 24268 29656
rect 24228 28762 24256 29650
rect 24412 29102 24440 31758
rect 24400 29096 24452 29102
rect 24400 29038 24452 29044
rect 24504 28778 24532 33390
rect 25148 32910 25176 33934
rect 25240 33114 25268 34002
rect 26252 33930 26280 35566
rect 26344 35494 26372 36110
rect 26620 35494 26648 36654
rect 30012 36576 30064 36582
rect 30012 36518 30064 36524
rect 30024 36242 30052 36518
rect 30012 36236 30064 36242
rect 30012 36178 30064 36184
rect 29644 36168 29696 36174
rect 29644 36110 29696 36116
rect 29736 36168 29788 36174
rect 29736 36110 29788 36116
rect 27344 36032 27396 36038
rect 27344 35974 27396 35980
rect 27356 35630 27384 35974
rect 29656 35834 29684 36110
rect 29644 35828 29696 35834
rect 29644 35770 29696 35776
rect 27712 35760 27764 35766
rect 27712 35702 27764 35708
rect 26792 35624 26844 35630
rect 26792 35566 26844 35572
rect 27344 35624 27396 35630
rect 27620 35624 27672 35630
rect 27344 35566 27396 35572
rect 27540 35572 27620 35578
rect 27540 35566 27672 35572
rect 26332 35488 26384 35494
rect 26332 35430 26384 35436
rect 26608 35488 26660 35494
rect 26608 35430 26660 35436
rect 26344 34950 26372 35430
rect 26620 35086 26648 35430
rect 26804 35154 26832 35566
rect 27068 35556 27120 35562
rect 27068 35498 27120 35504
rect 27540 35550 27660 35566
rect 27080 35154 27108 35498
rect 27540 35154 27568 35550
rect 26792 35148 26844 35154
rect 26792 35090 26844 35096
rect 27068 35148 27120 35154
rect 27068 35090 27120 35096
rect 27252 35148 27304 35154
rect 27252 35090 27304 35096
rect 27528 35148 27580 35154
rect 27528 35090 27580 35096
rect 26608 35080 26660 35086
rect 26608 35022 26660 35028
rect 26332 34944 26384 34950
rect 26332 34886 26384 34892
rect 26344 34542 26372 34886
rect 26332 34536 26384 34542
rect 26332 34478 26384 34484
rect 27080 34134 27108 35090
rect 27264 34610 27292 35090
rect 27724 35018 27752 35702
rect 29748 35630 29776 36110
rect 29736 35624 29788 35630
rect 29736 35566 29788 35572
rect 29748 35154 29776 35566
rect 30668 35222 30696 38218
rect 30944 35850 30972 40200
rect 32968 38214 32996 40200
rect 35176 38298 35204 40200
rect 36082 38720 36138 38729
rect 36082 38655 36138 38664
rect 35176 38270 35296 38298
rect 32956 38208 33008 38214
rect 32956 38150 33008 38156
rect 34940 38108 35236 38128
rect 34996 38106 35020 38108
rect 35076 38106 35100 38108
rect 35156 38106 35180 38108
rect 35018 38054 35020 38106
rect 35082 38054 35094 38106
rect 35156 38054 35158 38106
rect 34996 38052 35020 38054
rect 35076 38052 35100 38054
rect 35156 38052 35180 38054
rect 34940 38032 35236 38052
rect 34612 37868 34664 37874
rect 34612 37810 34664 37816
rect 31484 37800 31536 37806
rect 31484 37742 31536 37748
rect 33600 37800 33652 37806
rect 33600 37742 33652 37748
rect 31024 37732 31076 37738
rect 31024 37674 31076 37680
rect 30852 35822 30972 35850
rect 30852 35766 30880 35822
rect 30840 35760 30892 35766
rect 30840 35702 30892 35708
rect 30748 35488 30800 35494
rect 30748 35430 30800 35436
rect 30656 35216 30708 35222
rect 30656 35158 30708 35164
rect 30760 35154 30788 35430
rect 29736 35148 29788 35154
rect 29736 35090 29788 35096
rect 30748 35148 30800 35154
rect 30748 35090 30800 35096
rect 27712 35012 27764 35018
rect 27712 34954 27764 34960
rect 27252 34604 27304 34610
rect 27252 34546 27304 34552
rect 27264 34202 27292 34546
rect 27252 34196 27304 34202
rect 27252 34138 27304 34144
rect 27068 34128 27120 34134
rect 27068 34070 27120 34076
rect 27264 34066 27292 34138
rect 27724 34066 27752 34954
rect 29552 34944 29604 34950
rect 29552 34886 29604 34892
rect 29564 34610 29592 34886
rect 29552 34604 29604 34610
rect 29552 34546 29604 34552
rect 28172 34536 28224 34542
rect 28172 34478 28224 34484
rect 29368 34536 29420 34542
rect 29420 34484 29500 34490
rect 29368 34478 29500 34484
rect 27252 34060 27304 34066
rect 27252 34002 27304 34008
rect 27712 34060 27764 34066
rect 27712 34002 27764 34008
rect 26240 33924 26292 33930
rect 26240 33866 26292 33872
rect 28184 33862 28212 34478
rect 29380 34462 29500 34478
rect 28356 34400 28408 34406
rect 28356 34342 28408 34348
rect 28368 34134 28396 34342
rect 28356 34128 28408 34134
rect 28356 34070 28408 34076
rect 29472 33998 29500 34462
rect 30656 34400 30708 34406
rect 30656 34342 30708 34348
rect 29460 33992 29512 33998
rect 29460 33934 29512 33940
rect 28172 33856 28224 33862
rect 28172 33798 28224 33804
rect 29472 33522 29500 33934
rect 29552 33652 29604 33658
rect 29552 33594 29604 33600
rect 27160 33516 27212 33522
rect 27160 33458 27212 33464
rect 29460 33516 29512 33522
rect 29460 33458 29512 33464
rect 25228 33108 25280 33114
rect 25228 33050 25280 33056
rect 27172 32910 27200 33458
rect 27620 33448 27672 33454
rect 27620 33390 27672 33396
rect 25136 32904 25188 32910
rect 25136 32846 25188 32852
rect 27160 32904 27212 32910
rect 27160 32846 27212 32852
rect 27436 32904 27488 32910
rect 27436 32846 27488 32852
rect 25596 32768 25648 32774
rect 25596 32710 25648 32716
rect 25608 32434 25636 32710
rect 27448 32570 27476 32846
rect 27632 32774 27660 33390
rect 27896 33312 27948 33318
rect 27896 33254 27948 33260
rect 27620 32768 27672 32774
rect 27620 32710 27672 32716
rect 27436 32564 27488 32570
rect 27436 32506 27488 32512
rect 25596 32428 25648 32434
rect 25596 32370 25648 32376
rect 25780 32360 25832 32366
rect 25780 32302 25832 32308
rect 26056 32360 26108 32366
rect 26056 32302 26108 32308
rect 25792 32026 25820 32302
rect 25780 32020 25832 32026
rect 25780 31962 25832 31968
rect 26068 31822 26096 32302
rect 27160 32224 27212 32230
rect 27160 32166 27212 32172
rect 27172 31890 27200 32166
rect 27252 32020 27304 32026
rect 27252 31962 27304 31968
rect 27160 31884 27212 31890
rect 27160 31826 27212 31832
rect 24676 31816 24728 31822
rect 24676 31758 24728 31764
rect 26056 31816 26108 31822
rect 26056 31758 26108 31764
rect 24584 30796 24636 30802
rect 24584 30738 24636 30744
rect 24596 29782 24624 30738
rect 24584 29776 24636 29782
rect 24584 29718 24636 29724
rect 24584 29164 24636 29170
rect 24584 29106 24636 29112
rect 24216 28756 24268 28762
rect 24216 28698 24268 28704
rect 24320 28750 24532 28778
rect 23952 28070 24072 28098
rect 24228 28082 24256 28698
rect 24044 27946 24072 28070
rect 24216 28076 24268 28082
rect 24216 28018 24268 28024
rect 24032 27940 24084 27946
rect 24032 27882 24084 27888
rect 24044 27606 24072 27882
rect 23848 27600 23900 27606
rect 23848 27542 23900 27548
rect 24032 27600 24084 27606
rect 24032 27542 24084 27548
rect 23848 27328 23900 27334
rect 23848 27270 23900 27276
rect 23860 26858 23888 27270
rect 24124 27056 24176 27062
rect 24124 26998 24176 27004
rect 23848 26852 23900 26858
rect 23848 26794 23900 26800
rect 23860 26246 23888 26794
rect 24136 26382 24164 26998
rect 24216 26444 24268 26450
rect 24216 26386 24268 26392
rect 24124 26376 24176 26382
rect 24124 26318 24176 26324
rect 23848 26240 23900 26246
rect 23848 26182 23900 26188
rect 23664 25832 23716 25838
rect 23664 25774 23716 25780
rect 23480 25492 23532 25498
rect 23480 25434 23532 25440
rect 23756 25152 23808 25158
rect 23756 25094 23808 25100
rect 23664 24812 23716 24818
rect 23664 24754 23716 24760
rect 23572 23860 23624 23866
rect 23572 23802 23624 23808
rect 23388 23724 23440 23730
rect 23388 23666 23440 23672
rect 23296 23044 23348 23050
rect 23296 22986 23348 22992
rect 22836 22568 22888 22574
rect 22836 22510 22888 22516
rect 23020 22568 23072 22574
rect 23020 22510 23072 22516
rect 22848 22098 22876 22510
rect 23584 22506 23612 23802
rect 23676 23186 23704 24754
rect 23768 24274 23796 25094
rect 24228 24818 24256 26386
rect 24216 24812 24268 24818
rect 24216 24754 24268 24760
rect 23848 24744 23900 24750
rect 23848 24686 23900 24692
rect 23756 24268 23808 24274
rect 23756 24210 23808 24216
rect 23860 24154 23888 24686
rect 24320 24614 24348 28750
rect 24400 28620 24452 28626
rect 24400 28562 24452 28568
rect 24412 27878 24440 28562
rect 24596 28150 24624 29106
rect 24688 28558 24716 31758
rect 27172 31278 27200 31826
rect 27264 31822 27292 31962
rect 27344 31952 27396 31958
rect 27344 31894 27396 31900
rect 27252 31816 27304 31822
rect 27252 31758 27304 31764
rect 27356 31482 27384 31894
rect 27620 31816 27672 31822
rect 27620 31758 27672 31764
rect 27344 31476 27396 31482
rect 27344 31418 27396 31424
rect 26240 31272 26292 31278
rect 26240 31214 26292 31220
rect 26424 31272 26476 31278
rect 26424 31214 26476 31220
rect 27160 31272 27212 31278
rect 27160 31214 27212 31220
rect 25320 30796 25372 30802
rect 25320 30738 25372 30744
rect 25228 30184 25280 30190
rect 25228 30126 25280 30132
rect 25240 29238 25268 30126
rect 25332 29850 25360 30738
rect 25596 30592 25648 30598
rect 25596 30534 25648 30540
rect 25320 29844 25372 29850
rect 25320 29786 25372 29792
rect 25412 29844 25464 29850
rect 25412 29786 25464 29792
rect 25320 29708 25372 29714
rect 25424 29696 25452 29786
rect 25372 29668 25452 29696
rect 25320 29650 25372 29656
rect 25228 29232 25280 29238
rect 25228 29174 25280 29180
rect 24768 29096 24820 29102
rect 24768 29038 24820 29044
rect 24780 28762 24808 29038
rect 24768 28756 24820 28762
rect 24768 28698 24820 28704
rect 25424 28626 25452 29668
rect 25608 29102 25636 30534
rect 26252 30394 26280 31214
rect 26240 30388 26292 30394
rect 26240 30330 26292 30336
rect 26056 30252 26108 30258
rect 26056 30194 26108 30200
rect 25596 29096 25648 29102
rect 25596 29038 25648 29044
rect 24768 28620 24820 28626
rect 24768 28562 24820 28568
rect 25412 28620 25464 28626
rect 25412 28562 25464 28568
rect 24676 28552 24728 28558
rect 24676 28494 24728 28500
rect 24780 28218 24808 28562
rect 24768 28212 24820 28218
rect 24768 28154 24820 28160
rect 24584 28144 24636 28150
rect 24584 28086 24636 28092
rect 24584 28008 24636 28014
rect 24584 27950 24636 27956
rect 24400 27872 24452 27878
rect 24400 27814 24452 27820
rect 24412 27538 24440 27814
rect 24596 27606 24624 27950
rect 24676 27940 24728 27946
rect 24676 27882 24728 27888
rect 24688 27674 24716 27882
rect 24676 27668 24728 27674
rect 24676 27610 24728 27616
rect 24584 27600 24636 27606
rect 24584 27542 24636 27548
rect 24400 27532 24452 27538
rect 24400 27474 24452 27480
rect 24492 27532 24544 27538
rect 24492 27474 24544 27480
rect 24504 27130 24532 27474
rect 24492 27124 24544 27130
rect 24492 27066 24544 27072
rect 24596 26586 24624 27542
rect 24584 26580 24636 26586
rect 24584 26522 24636 26528
rect 24400 26376 24452 26382
rect 24400 26318 24452 26324
rect 24412 24954 24440 26318
rect 24688 25906 24716 27610
rect 25424 26874 25452 28562
rect 26068 28082 26096 30194
rect 26436 29102 26464 31214
rect 26884 30728 26936 30734
rect 26884 30670 26936 30676
rect 26976 30728 27028 30734
rect 26976 30670 27028 30676
rect 26896 29646 26924 30670
rect 26988 30394 27016 30670
rect 27632 30666 27660 31758
rect 27712 31408 27764 31414
rect 27712 31350 27764 31356
rect 27724 30802 27752 31350
rect 27908 31210 27936 33254
rect 29564 32978 29592 33594
rect 30668 33522 30696 34342
rect 30656 33516 30708 33522
rect 30656 33458 30708 33464
rect 29552 32972 29604 32978
rect 29552 32914 29604 32920
rect 30380 32972 30432 32978
rect 30380 32914 30432 32920
rect 29276 32904 29328 32910
rect 29276 32846 29328 32852
rect 28080 32496 28132 32502
rect 28080 32438 28132 32444
rect 27896 31204 27948 31210
rect 27896 31146 27948 31152
rect 27712 30796 27764 30802
rect 27712 30738 27764 30744
rect 27620 30660 27672 30666
rect 27620 30602 27672 30608
rect 26976 30388 27028 30394
rect 26976 30330 27028 30336
rect 27344 30184 27396 30190
rect 27344 30126 27396 30132
rect 27356 29782 27384 30126
rect 27344 29776 27396 29782
rect 27344 29718 27396 29724
rect 28092 29714 28120 32438
rect 29288 32434 29316 32846
rect 29276 32428 29328 32434
rect 29276 32370 29328 32376
rect 28632 32360 28684 32366
rect 28632 32302 28684 32308
rect 28816 32360 28868 32366
rect 28816 32302 28868 32308
rect 28644 32042 28672 32302
rect 28644 32014 28764 32042
rect 28448 31680 28500 31686
rect 28448 31622 28500 31628
rect 28460 31142 28488 31622
rect 28540 31204 28592 31210
rect 28540 31146 28592 31152
rect 28448 31136 28500 31142
rect 28448 31078 28500 31084
rect 28552 31090 28580 31146
rect 28552 31062 28672 31090
rect 28172 30796 28224 30802
rect 28172 30738 28224 30744
rect 28080 29708 28132 29714
rect 28080 29650 28132 29656
rect 26884 29640 26936 29646
rect 26884 29582 26936 29588
rect 27252 29572 27304 29578
rect 27252 29514 27304 29520
rect 27264 29102 27292 29514
rect 28080 29164 28132 29170
rect 28080 29106 28132 29112
rect 26424 29096 26476 29102
rect 26424 29038 26476 29044
rect 27252 29096 27304 29102
rect 27252 29038 27304 29044
rect 27264 28762 27292 29038
rect 27712 28960 27764 28966
rect 27712 28902 27764 28908
rect 27252 28756 27304 28762
rect 27252 28698 27304 28704
rect 27264 28626 27292 28698
rect 27252 28620 27304 28626
rect 27252 28562 27304 28568
rect 26608 28416 26660 28422
rect 26608 28358 26660 28364
rect 26056 28076 26108 28082
rect 26056 28018 26108 28024
rect 26068 27962 26096 28018
rect 26240 28008 26292 28014
rect 26068 27934 26188 27962
rect 26240 27950 26292 27956
rect 25596 26920 25648 26926
rect 25424 26846 25544 26874
rect 25596 26862 25648 26868
rect 25412 26784 25464 26790
rect 25412 26726 25464 26732
rect 24952 26444 25004 26450
rect 24952 26386 25004 26392
rect 24860 26240 24912 26246
rect 24860 26182 24912 26188
rect 24676 25900 24728 25906
rect 24676 25842 24728 25848
rect 24584 25832 24636 25838
rect 24584 25774 24636 25780
rect 24400 24948 24452 24954
rect 24400 24890 24452 24896
rect 24308 24608 24360 24614
rect 24308 24550 24360 24556
rect 24032 24268 24084 24274
rect 24032 24210 24084 24216
rect 23768 24126 23888 24154
rect 23664 23180 23716 23186
rect 23664 23122 23716 23128
rect 23768 23032 23796 24126
rect 23848 23656 23900 23662
rect 23848 23598 23900 23604
rect 23676 23004 23796 23032
rect 23572 22500 23624 22506
rect 23572 22442 23624 22448
rect 23676 22438 23704 23004
rect 23860 22574 23888 23598
rect 23940 23180 23992 23186
rect 23940 23122 23992 23128
rect 23952 22642 23980 23122
rect 24044 22642 24072 24210
rect 23940 22636 23992 22642
rect 23940 22578 23992 22584
rect 24032 22636 24084 22642
rect 24032 22578 24084 22584
rect 24216 22636 24268 22642
rect 24216 22578 24268 22584
rect 23756 22568 23808 22574
rect 23756 22510 23808 22516
rect 23848 22568 23900 22574
rect 23848 22510 23900 22516
rect 23664 22432 23716 22438
rect 23664 22374 23716 22380
rect 22744 22092 22796 22098
rect 22744 22034 22796 22040
rect 22836 22092 22888 22098
rect 22836 22034 22888 22040
rect 23388 22092 23440 22098
rect 23388 22034 23440 22040
rect 22652 21956 22704 21962
rect 22652 21898 22704 21904
rect 22560 20936 22612 20942
rect 22560 20878 22612 20884
rect 22572 20466 22600 20878
rect 22560 20460 22612 20466
rect 22560 20402 22612 20408
rect 22560 19712 22612 19718
rect 22560 19654 22612 19660
rect 22468 18828 22520 18834
rect 22572 18816 22600 19654
rect 22520 18788 22600 18816
rect 22468 18770 22520 18776
rect 22572 18222 22600 18788
rect 22560 18216 22612 18222
rect 22560 18158 22612 18164
rect 22572 17116 22600 18158
rect 22664 17270 22692 21898
rect 22756 20806 22784 22034
rect 22928 21888 22980 21894
rect 22928 21830 22980 21836
rect 22940 21434 22968 21830
rect 23400 21690 23428 22034
rect 23388 21684 23440 21690
rect 23388 21626 23440 21632
rect 23400 21486 23428 21626
rect 23572 21616 23624 21622
rect 23572 21558 23624 21564
rect 23480 21548 23532 21554
rect 23480 21490 23532 21496
rect 23388 21480 23440 21486
rect 22940 21406 23060 21434
rect 23388 21422 23440 21428
rect 22928 21344 22980 21350
rect 22928 21286 22980 21292
rect 22940 21146 22968 21286
rect 22928 21140 22980 21146
rect 22928 21082 22980 21088
rect 22836 21004 22888 21010
rect 22836 20946 22888 20952
rect 22848 20806 22876 20946
rect 22744 20800 22796 20806
rect 22744 20742 22796 20748
rect 22836 20800 22888 20806
rect 22836 20742 22888 20748
rect 22756 18222 22784 20742
rect 22848 20398 22876 20742
rect 22836 20392 22888 20398
rect 22836 20334 22888 20340
rect 22928 20392 22980 20398
rect 22928 20334 22980 20340
rect 22940 19718 22968 20334
rect 23032 19961 23060 21406
rect 23204 21412 23256 21418
rect 23204 21354 23256 21360
rect 23216 21146 23244 21354
rect 23112 21140 23164 21146
rect 23112 21082 23164 21088
rect 23204 21140 23256 21146
rect 23204 21082 23256 21088
rect 23018 19952 23074 19961
rect 23018 19887 23074 19896
rect 22928 19712 22980 19718
rect 22928 19654 22980 19660
rect 22928 19168 22980 19174
rect 22928 19110 22980 19116
rect 22836 18828 22888 18834
rect 22836 18770 22888 18776
rect 22848 18426 22876 18770
rect 22836 18420 22888 18426
rect 22836 18362 22888 18368
rect 22744 18216 22796 18222
rect 22744 18158 22796 18164
rect 22756 17814 22784 18158
rect 22744 17808 22796 17814
rect 22744 17750 22796 17756
rect 22940 17746 22968 19110
rect 22928 17740 22980 17746
rect 22928 17682 22980 17688
rect 22652 17264 22704 17270
rect 22652 17206 22704 17212
rect 22744 17196 22796 17202
rect 22744 17138 22796 17144
rect 22572 17088 22692 17116
rect 22560 16516 22612 16522
rect 22560 16458 22612 16464
rect 22572 15570 22600 16458
rect 22664 16046 22692 17088
rect 22756 16658 22784 17138
rect 22744 16652 22796 16658
rect 22744 16594 22796 16600
rect 22940 16046 22968 17682
rect 22652 16040 22704 16046
rect 22652 15982 22704 15988
rect 22928 16040 22980 16046
rect 22928 15982 22980 15988
rect 22664 15570 22692 15982
rect 22560 15564 22612 15570
rect 22560 15506 22612 15512
rect 22652 15564 22704 15570
rect 22652 15506 22704 15512
rect 22940 15366 22968 15982
rect 23032 15910 23060 19887
rect 23020 15904 23072 15910
rect 23020 15846 23072 15852
rect 22928 15360 22980 15366
rect 22928 15302 22980 15308
rect 22744 15088 22796 15094
rect 22744 15030 22796 15036
rect 23020 15088 23072 15094
rect 23020 15030 23072 15036
rect 22560 14884 22612 14890
rect 22560 14826 22612 14832
rect 22572 13938 22600 14826
rect 22756 14414 22784 15030
rect 23032 14482 23060 15030
rect 23124 14958 23152 21082
rect 23492 20398 23520 21490
rect 23584 21078 23612 21558
rect 23572 21072 23624 21078
rect 23572 21014 23624 21020
rect 23480 20392 23532 20398
rect 23480 20334 23532 20340
rect 23204 19236 23256 19242
rect 23204 19178 23256 19184
rect 23216 18970 23244 19178
rect 23204 18964 23256 18970
rect 23204 18906 23256 18912
rect 23204 18828 23256 18834
rect 23204 18770 23256 18776
rect 23216 18698 23244 18770
rect 23204 18692 23256 18698
rect 23204 18634 23256 18640
rect 23204 18148 23256 18154
rect 23204 18090 23256 18096
rect 23112 14952 23164 14958
rect 23112 14894 23164 14900
rect 23124 14482 23152 14894
rect 23020 14476 23072 14482
rect 23020 14418 23072 14424
rect 23112 14476 23164 14482
rect 23112 14418 23164 14424
rect 22744 14408 22796 14414
rect 22744 14350 22796 14356
rect 22560 13932 22612 13938
rect 22560 13874 22612 13880
rect 22468 13796 22520 13802
rect 22468 13738 22520 13744
rect 22480 12374 22508 13738
rect 22560 13388 22612 13394
rect 22560 13330 22612 13336
rect 22572 12442 22600 13330
rect 22652 12640 22704 12646
rect 22652 12582 22704 12588
rect 22560 12436 22612 12442
rect 22560 12378 22612 12384
rect 22468 12368 22520 12374
rect 22468 12310 22520 12316
rect 22664 11762 22692 12582
rect 22652 11756 22704 11762
rect 22652 11698 22704 11704
rect 22468 11280 22520 11286
rect 22468 11222 22520 11228
rect 22480 8430 22508 11222
rect 22836 11212 22888 11218
rect 22836 11154 22888 11160
rect 22848 10674 22876 11154
rect 23124 11082 23152 14418
rect 23112 11076 23164 11082
rect 23112 11018 23164 11024
rect 22836 10668 22888 10674
rect 22836 10610 22888 10616
rect 22652 10600 22704 10606
rect 22652 10542 22704 10548
rect 22664 8430 22692 10542
rect 22848 10266 22876 10610
rect 23216 10606 23244 18090
rect 23480 17332 23532 17338
rect 23480 17274 23532 17280
rect 23492 16046 23520 17274
rect 23572 17128 23624 17134
rect 23572 17070 23624 17076
rect 23584 16522 23612 17070
rect 23572 16516 23624 16522
rect 23572 16458 23624 16464
rect 23480 16040 23532 16046
rect 23480 15982 23532 15988
rect 23296 15564 23348 15570
rect 23296 15506 23348 15512
rect 23308 14278 23336 15506
rect 23388 15360 23440 15366
rect 23388 15302 23440 15308
rect 23400 14550 23428 15302
rect 23676 14822 23704 22374
rect 23768 22234 23796 22510
rect 23756 22228 23808 22234
rect 23756 22170 23808 22176
rect 23940 21480 23992 21486
rect 23940 21422 23992 21428
rect 23848 20256 23900 20262
rect 23848 20198 23900 20204
rect 23860 19904 23888 20198
rect 23768 19876 23888 19904
rect 23768 17610 23796 19876
rect 23848 19780 23900 19786
rect 23848 19722 23900 19728
rect 23860 19310 23888 19722
rect 23848 19304 23900 19310
rect 23848 19246 23900 19252
rect 23860 18902 23888 19246
rect 23848 18896 23900 18902
rect 23848 18838 23900 18844
rect 23848 18692 23900 18698
rect 23848 18634 23900 18640
rect 23860 18290 23888 18634
rect 23952 18358 23980 21422
rect 24124 21072 24176 21078
rect 24124 21014 24176 21020
rect 24032 19440 24084 19446
rect 24032 19382 24084 19388
rect 23940 18352 23992 18358
rect 23940 18294 23992 18300
rect 23848 18284 23900 18290
rect 23848 18226 23900 18232
rect 23860 17746 23888 18226
rect 24044 17882 24072 19382
rect 24032 17876 24084 17882
rect 24032 17818 24084 17824
rect 24136 17762 24164 21014
rect 24228 20942 24256 22578
rect 24400 21004 24452 21010
rect 24400 20946 24452 20952
rect 24216 20936 24268 20942
rect 24216 20878 24268 20884
rect 24228 17814 24256 20878
rect 24412 20398 24440 20946
rect 24400 20392 24452 20398
rect 24400 20334 24452 20340
rect 24308 20256 24360 20262
rect 24308 20198 24360 20204
rect 24320 18766 24348 20198
rect 24400 18828 24452 18834
rect 24400 18770 24452 18776
rect 24308 18760 24360 18766
rect 24308 18702 24360 18708
rect 23848 17740 23900 17746
rect 23848 17682 23900 17688
rect 23952 17734 24164 17762
rect 24216 17808 24268 17814
rect 24216 17750 24268 17756
rect 23756 17604 23808 17610
rect 23756 17546 23808 17552
rect 23768 16658 23796 17546
rect 23756 16652 23808 16658
rect 23756 16594 23808 16600
rect 23952 16538 23980 17734
rect 24320 17542 24348 18702
rect 24124 17536 24176 17542
rect 24124 17478 24176 17484
rect 24308 17536 24360 17542
rect 24308 17478 24360 17484
rect 24032 17264 24084 17270
rect 24032 17206 24084 17212
rect 24044 16726 24072 17206
rect 24032 16720 24084 16726
rect 24032 16662 24084 16668
rect 23768 16510 23980 16538
rect 23664 14816 23716 14822
rect 23664 14758 23716 14764
rect 23676 14618 23704 14758
rect 23664 14612 23716 14618
rect 23664 14554 23716 14560
rect 23388 14544 23440 14550
rect 23388 14486 23440 14492
rect 23296 14272 23348 14278
rect 23296 14214 23348 14220
rect 23572 14272 23624 14278
rect 23572 14214 23624 14220
rect 23294 12744 23350 12753
rect 23294 12679 23296 12688
rect 23348 12679 23350 12688
rect 23296 12650 23348 12656
rect 23388 12640 23440 12646
rect 23388 12582 23440 12588
rect 23400 12306 23428 12582
rect 23388 12300 23440 12306
rect 23388 12242 23440 12248
rect 23480 12164 23532 12170
rect 23480 12106 23532 12112
rect 23388 12096 23440 12102
rect 23388 12038 23440 12044
rect 23400 11830 23428 12038
rect 23492 11898 23520 12106
rect 23480 11892 23532 11898
rect 23480 11834 23532 11840
rect 23388 11824 23440 11830
rect 23388 11766 23440 11772
rect 23296 11688 23348 11694
rect 23296 11630 23348 11636
rect 23308 11218 23336 11630
rect 23388 11552 23440 11558
rect 23388 11494 23440 11500
rect 23296 11212 23348 11218
rect 23296 11154 23348 11160
rect 23204 10600 23256 10606
rect 23204 10542 23256 10548
rect 23308 10538 23336 11154
rect 23296 10532 23348 10538
rect 23296 10474 23348 10480
rect 22836 10260 22888 10266
rect 22836 10202 22888 10208
rect 23400 10130 23428 11494
rect 23388 10124 23440 10130
rect 23388 10066 23440 10072
rect 22744 10056 22796 10062
rect 22744 9998 22796 10004
rect 22756 9722 22784 9998
rect 22744 9716 22796 9722
rect 22744 9658 22796 9664
rect 23296 9648 23348 9654
rect 23296 9590 23348 9596
rect 22836 9512 22888 9518
rect 22836 9454 22888 9460
rect 23112 9512 23164 9518
rect 23112 9454 23164 9460
rect 22848 9081 22876 9454
rect 22834 9072 22890 9081
rect 22834 9007 22890 9016
rect 22468 8424 22520 8430
rect 22468 8366 22520 8372
rect 22652 8424 22704 8430
rect 22652 8366 22704 8372
rect 22480 7750 22508 8366
rect 22468 7744 22520 7750
rect 22468 7686 22520 7692
rect 22296 7534 22416 7562
rect 21916 6656 21968 6662
rect 22192 6656 22244 6662
rect 21916 6598 21968 6604
rect 22112 6616 22192 6644
rect 22112 6322 22140 6616
rect 22192 6598 22244 6604
rect 22100 6316 22152 6322
rect 22100 6258 22152 6264
rect 21732 5772 21784 5778
rect 21732 5714 21784 5720
rect 21640 5704 21692 5710
rect 21640 5646 21692 5652
rect 21824 5704 21876 5710
rect 21824 5646 21876 5652
rect 21652 5574 21680 5646
rect 21640 5568 21692 5574
rect 21640 5510 21692 5516
rect 21732 5228 21784 5234
rect 21732 5170 21784 5176
rect 21548 4616 21600 4622
rect 21548 4558 21600 4564
rect 20720 4548 20772 4554
rect 20720 4490 20772 4496
rect 20444 4140 20496 4146
rect 20444 4082 20496 4088
rect 21744 4078 21772 5170
rect 21836 4690 21864 5646
rect 22100 5160 22152 5166
rect 22100 5102 22152 5108
rect 21824 4684 21876 4690
rect 21824 4626 21876 4632
rect 22112 4214 22140 5102
rect 22192 5092 22244 5098
rect 22192 5034 22244 5040
rect 22100 4208 22152 4214
rect 22100 4150 22152 4156
rect 22204 4078 22232 5034
rect 21732 4072 21784 4078
rect 21732 4014 21784 4020
rect 22192 4072 22244 4078
rect 22192 4014 22244 4020
rect 20996 4004 21048 4010
rect 20996 3946 21048 3952
rect 21008 3738 21036 3946
rect 20996 3732 21048 3738
rect 20996 3674 21048 3680
rect 21364 3596 21416 3602
rect 21364 3538 21416 3544
rect 21376 2582 21404 3538
rect 21744 3534 21772 4014
rect 21732 3528 21784 3534
rect 21732 3470 21784 3476
rect 22100 3528 22152 3534
rect 22100 3470 22152 3476
rect 21548 3392 21600 3398
rect 21548 3334 21600 3340
rect 21364 2576 21416 2582
rect 21364 2518 21416 2524
rect 20076 2100 20128 2106
rect 20076 2042 20128 2048
rect 19892 1964 19944 1970
rect 19892 1906 19944 1912
rect 21560 800 21588 3334
rect 21744 2972 21772 3470
rect 21824 2984 21876 2990
rect 21744 2944 21824 2972
rect 21824 2926 21876 2932
rect 22112 2514 22140 3470
rect 22296 3466 22324 7534
rect 22376 7472 22428 7478
rect 22376 7414 22428 7420
rect 22480 7426 22508 7686
rect 22388 5778 22416 7414
rect 22480 7398 22600 7426
rect 22468 7336 22520 7342
rect 22468 7278 22520 7284
rect 22480 6322 22508 7278
rect 22572 6798 22600 7398
rect 22652 7200 22704 7206
rect 22652 7142 22704 7148
rect 22664 7002 22692 7142
rect 22652 6996 22704 7002
rect 22652 6938 22704 6944
rect 22560 6792 22612 6798
rect 22560 6734 22612 6740
rect 22468 6316 22520 6322
rect 22468 6258 22520 6264
rect 22572 6202 22600 6734
rect 22480 6186 22600 6202
rect 22468 6180 22600 6186
rect 22520 6174 22600 6180
rect 22468 6122 22520 6128
rect 22376 5772 22428 5778
rect 22376 5714 22428 5720
rect 22664 3602 22692 6938
rect 23124 6866 23152 9454
rect 23308 8566 23336 9590
rect 23400 9178 23428 10066
rect 23584 9761 23612 14214
rect 23664 13864 23716 13870
rect 23664 13806 23716 13812
rect 23676 12782 23704 13806
rect 23768 13530 23796 16510
rect 24136 16130 24164 17478
rect 24412 17134 24440 18770
rect 24492 17196 24544 17202
rect 24492 17138 24544 17144
rect 24400 17128 24452 17134
rect 24400 17070 24452 17076
rect 24308 16992 24360 16998
rect 24308 16934 24360 16940
rect 24216 16448 24268 16454
rect 24216 16390 24268 16396
rect 24044 16102 24164 16130
rect 23848 16040 23900 16046
rect 23848 15982 23900 15988
rect 23756 13524 23808 13530
rect 23756 13466 23808 13472
rect 23754 13288 23810 13297
rect 23754 13223 23810 13232
rect 23664 12776 23716 12782
rect 23768 12753 23796 13223
rect 23664 12718 23716 12724
rect 23754 12744 23810 12753
rect 23754 12679 23810 12688
rect 23768 11898 23796 12679
rect 23756 11892 23808 11898
rect 23756 11834 23808 11840
rect 23756 10192 23808 10198
rect 23756 10134 23808 10140
rect 23570 9752 23626 9761
rect 23570 9687 23626 9696
rect 23478 9616 23534 9625
rect 23478 9551 23534 9560
rect 23388 9172 23440 9178
rect 23388 9114 23440 9120
rect 23492 9042 23520 9551
rect 23664 9512 23716 9518
rect 23662 9480 23664 9489
rect 23716 9480 23718 9489
rect 23662 9415 23718 9424
rect 23768 9110 23796 10134
rect 23756 9104 23808 9110
rect 23756 9046 23808 9052
rect 23860 9042 23888 15982
rect 24044 15502 24072 16102
rect 24124 16040 24176 16046
rect 24124 15982 24176 15988
rect 24136 15570 24164 15982
rect 24124 15564 24176 15570
rect 24124 15506 24176 15512
rect 24032 15496 24084 15502
rect 24032 15438 24084 15444
rect 23940 14816 23992 14822
rect 24044 14804 24072 15438
rect 24124 14884 24176 14890
rect 24124 14826 24176 14832
rect 23992 14776 24072 14804
rect 23940 14758 23992 14764
rect 23940 13320 23992 13326
rect 23940 13262 23992 13268
rect 23952 12850 23980 13262
rect 23940 12844 23992 12850
rect 23940 12786 23992 12792
rect 24032 12640 24084 12646
rect 24032 12582 24084 12588
rect 23940 11892 23992 11898
rect 23940 11834 23992 11840
rect 23480 9036 23532 9042
rect 23480 8978 23532 8984
rect 23848 9036 23900 9042
rect 23848 8978 23900 8984
rect 23388 8968 23440 8974
rect 23388 8910 23440 8916
rect 23296 8560 23348 8566
rect 23296 8502 23348 8508
rect 23308 7954 23336 8502
rect 23296 7948 23348 7954
rect 23296 7890 23348 7896
rect 23400 7818 23428 8910
rect 23860 8634 23888 8978
rect 23848 8628 23900 8634
rect 23848 8570 23900 8576
rect 23388 7812 23440 7818
rect 23388 7754 23440 7760
rect 23848 7472 23900 7478
rect 23848 7414 23900 7420
rect 23860 7342 23888 7414
rect 23848 7336 23900 7342
rect 23848 7278 23900 7284
rect 23952 7206 23980 11834
rect 24044 9382 24072 12582
rect 24032 9376 24084 9382
rect 24032 9318 24084 9324
rect 24032 8968 24084 8974
rect 24032 8910 24084 8916
rect 24044 7954 24072 8910
rect 24032 7948 24084 7954
rect 24032 7890 24084 7896
rect 24044 7342 24072 7890
rect 24032 7336 24084 7342
rect 24032 7278 24084 7284
rect 23940 7200 23992 7206
rect 23940 7142 23992 7148
rect 23112 6860 23164 6866
rect 23112 6802 23164 6808
rect 24044 6254 24072 7278
rect 23940 6248 23992 6254
rect 23940 6190 23992 6196
rect 24032 6248 24084 6254
rect 24032 6190 24084 6196
rect 23952 5166 23980 6190
rect 24136 5710 24164 14826
rect 24228 14618 24256 16390
rect 24216 14612 24268 14618
rect 24216 14554 24268 14560
rect 24216 12776 24268 12782
rect 24216 12718 24268 12724
rect 24228 11898 24256 12718
rect 24216 11892 24268 11898
rect 24216 11834 24268 11840
rect 24216 11688 24268 11694
rect 24216 11630 24268 11636
rect 24228 10266 24256 11630
rect 24216 10260 24268 10266
rect 24216 10202 24268 10208
rect 24320 6458 24348 16934
rect 24412 16658 24440 17070
rect 24400 16652 24452 16658
rect 24400 16594 24452 16600
rect 24504 16590 24532 17138
rect 24492 16584 24544 16590
rect 24492 16526 24544 16532
rect 24504 16046 24532 16526
rect 24400 16040 24452 16046
rect 24400 15982 24452 15988
rect 24492 16040 24544 16046
rect 24492 15982 24544 15988
rect 24412 15910 24440 15982
rect 24400 15904 24452 15910
rect 24400 15846 24452 15852
rect 24412 15638 24440 15846
rect 24400 15632 24452 15638
rect 24400 15574 24452 15580
rect 24400 15496 24452 15502
rect 24504 15484 24532 15982
rect 24452 15456 24532 15484
rect 24400 15438 24452 15444
rect 24492 15360 24544 15366
rect 24492 15302 24544 15308
rect 24504 14958 24532 15302
rect 24492 14952 24544 14958
rect 24492 14894 24544 14900
rect 24492 14408 24544 14414
rect 24492 14350 24544 14356
rect 24504 11694 24532 14350
rect 24492 11688 24544 11694
rect 24492 11630 24544 11636
rect 24596 10826 24624 25774
rect 24872 25362 24900 26182
rect 24860 25356 24912 25362
rect 24860 25298 24912 25304
rect 24860 24268 24912 24274
rect 24860 24210 24912 24216
rect 24872 23662 24900 24210
rect 24860 23656 24912 23662
rect 24860 23598 24912 23604
rect 24676 22568 24728 22574
rect 24676 22510 24728 22516
rect 24688 21350 24716 22510
rect 24872 21978 24900 23598
rect 24780 21950 24900 21978
rect 24780 21434 24808 21950
rect 24860 21888 24912 21894
rect 24860 21830 24912 21836
rect 24872 21554 24900 21830
rect 24860 21548 24912 21554
rect 24860 21490 24912 21496
rect 24780 21406 24900 21434
rect 24676 21344 24728 21350
rect 24676 21286 24728 21292
rect 24688 21010 24716 21286
rect 24676 21004 24728 21010
rect 24676 20946 24728 20952
rect 24676 19780 24728 19786
rect 24676 19722 24728 19728
rect 24688 19310 24716 19722
rect 24676 19304 24728 19310
rect 24676 19246 24728 19252
rect 24688 18222 24716 19246
rect 24872 18902 24900 21406
rect 24964 21078 24992 26386
rect 25228 25900 25280 25906
rect 25228 25842 25280 25848
rect 25136 25764 25188 25770
rect 25136 25706 25188 25712
rect 25148 25362 25176 25706
rect 25136 25356 25188 25362
rect 25136 25298 25188 25304
rect 25240 25242 25268 25842
rect 25320 25832 25372 25838
rect 25320 25774 25372 25780
rect 25148 25214 25268 25242
rect 25148 24750 25176 25214
rect 25332 25158 25360 25774
rect 25320 25152 25372 25158
rect 25320 25094 25372 25100
rect 25424 24818 25452 26726
rect 25516 26042 25544 26846
rect 25504 26036 25556 26042
rect 25504 25978 25556 25984
rect 25504 24948 25556 24954
rect 25504 24890 25556 24896
rect 25412 24812 25464 24818
rect 25412 24754 25464 24760
rect 25136 24744 25188 24750
rect 25136 24686 25188 24692
rect 25148 23526 25176 24686
rect 25320 24268 25372 24274
rect 25320 24210 25372 24216
rect 25332 23730 25360 24210
rect 25320 23724 25372 23730
rect 25320 23666 25372 23672
rect 25136 23520 25188 23526
rect 25136 23462 25188 23468
rect 25044 23112 25096 23118
rect 25044 23054 25096 23060
rect 24952 21072 25004 21078
rect 24952 21014 25004 21020
rect 25056 19281 25084 23054
rect 25148 22574 25176 23462
rect 25136 22568 25188 22574
rect 25136 22510 25188 22516
rect 25412 22568 25464 22574
rect 25412 22510 25464 22516
rect 25148 22166 25176 22510
rect 25136 22160 25188 22166
rect 25136 22102 25188 22108
rect 25228 22092 25280 22098
rect 25228 22034 25280 22040
rect 25240 21690 25268 22034
rect 25228 21684 25280 21690
rect 25228 21626 25280 21632
rect 25424 21622 25452 22510
rect 25516 22166 25544 24890
rect 25608 23798 25636 26862
rect 26160 26246 26188 27934
rect 26252 27402 26280 27950
rect 26620 27538 26648 28358
rect 27264 28082 27292 28562
rect 27724 28558 27752 28902
rect 28092 28626 28120 29106
rect 28080 28620 28132 28626
rect 28080 28562 28132 28568
rect 27620 28552 27672 28558
rect 27620 28494 27672 28500
rect 27712 28552 27764 28558
rect 27712 28494 27764 28500
rect 27252 28076 27304 28082
rect 27252 28018 27304 28024
rect 27632 27946 27660 28494
rect 27620 27940 27672 27946
rect 27620 27882 27672 27888
rect 27632 27538 27660 27882
rect 26608 27532 26660 27538
rect 26608 27474 26660 27480
rect 27620 27532 27672 27538
rect 27620 27474 27672 27480
rect 27724 27470 27752 28494
rect 27804 28144 27856 28150
rect 27804 28086 27856 28092
rect 27712 27464 27764 27470
rect 27712 27406 27764 27412
rect 26240 27396 26292 27402
rect 26240 27338 26292 27344
rect 26608 26580 26660 26586
rect 26608 26522 26660 26528
rect 26516 26444 26568 26450
rect 26516 26386 26568 26392
rect 26148 26240 26200 26246
rect 26148 26182 26200 26188
rect 25780 26036 25832 26042
rect 25780 25978 25832 25984
rect 25688 24404 25740 24410
rect 25688 24346 25740 24352
rect 25596 23792 25648 23798
rect 25596 23734 25648 23740
rect 25700 23662 25728 24346
rect 25792 24274 25820 25978
rect 26160 25906 26188 26182
rect 26148 25900 26200 25906
rect 26148 25842 26200 25848
rect 26528 25430 26556 26386
rect 26516 25424 26568 25430
rect 26516 25366 26568 25372
rect 26528 24954 26556 25366
rect 26620 25362 26648 26522
rect 27724 26314 27752 27406
rect 27816 26926 27844 28086
rect 27988 27464 28040 27470
rect 27988 27406 28040 27412
rect 28000 26994 28028 27406
rect 27988 26988 28040 26994
rect 27988 26930 28040 26936
rect 27804 26920 27856 26926
rect 27804 26862 27856 26868
rect 27988 26376 28040 26382
rect 28040 26324 28120 26330
rect 27988 26318 28120 26324
rect 27712 26308 27764 26314
rect 28000 26302 28120 26318
rect 27712 26250 27764 26256
rect 26700 25832 26752 25838
rect 26700 25774 26752 25780
rect 26712 25498 26740 25774
rect 28092 25770 28120 26302
rect 28080 25764 28132 25770
rect 28080 25706 28132 25712
rect 28092 25498 28120 25706
rect 26700 25492 26752 25498
rect 26700 25434 26752 25440
rect 28080 25492 28132 25498
rect 28080 25434 28132 25440
rect 26608 25356 26660 25362
rect 26608 25298 26660 25304
rect 26516 24948 26568 24954
rect 26516 24890 26568 24896
rect 26792 24676 26844 24682
rect 26792 24618 26844 24624
rect 27620 24676 27672 24682
rect 27620 24618 27672 24624
rect 25780 24268 25832 24274
rect 25780 24210 25832 24216
rect 25964 24132 26016 24138
rect 25964 24074 26016 24080
rect 25976 23662 26004 24074
rect 25688 23656 25740 23662
rect 25688 23598 25740 23604
rect 25964 23656 26016 23662
rect 25964 23598 26016 23604
rect 26516 23588 26568 23594
rect 26516 23530 26568 23536
rect 25688 23180 25740 23186
rect 25688 23122 25740 23128
rect 25700 22574 25728 23122
rect 26240 23112 26292 23118
rect 26240 23054 26292 23060
rect 25688 22568 25740 22574
rect 25688 22510 25740 22516
rect 25504 22160 25556 22166
rect 25504 22102 25556 22108
rect 25596 22092 25648 22098
rect 25596 22034 25648 22040
rect 25412 21616 25464 21622
rect 25412 21558 25464 21564
rect 25136 21140 25188 21146
rect 25136 21082 25188 21088
rect 25148 20262 25176 21082
rect 25608 20602 25636 22034
rect 25964 22024 26016 22030
rect 25964 21966 26016 21972
rect 25976 21554 26004 21966
rect 26252 21962 26280 23054
rect 26528 22778 26556 23530
rect 26804 23186 26832 24618
rect 27344 24404 27396 24410
rect 27344 24346 27396 24352
rect 27356 24274 27384 24346
rect 27632 24274 27660 24618
rect 27344 24268 27396 24274
rect 27344 24210 27396 24216
rect 27620 24268 27672 24274
rect 27620 24210 27672 24216
rect 26976 23656 27028 23662
rect 26976 23598 27028 23604
rect 26988 23254 27016 23598
rect 27632 23526 27660 24210
rect 27620 23520 27672 23526
rect 27620 23462 27672 23468
rect 26976 23248 27028 23254
rect 26976 23190 27028 23196
rect 26792 23180 26844 23186
rect 26792 23122 26844 23128
rect 27632 23118 27660 23462
rect 27896 23248 27948 23254
rect 27896 23190 27948 23196
rect 27804 23180 27856 23186
rect 27804 23122 27856 23128
rect 27620 23112 27672 23118
rect 27620 23054 27672 23060
rect 26516 22772 26568 22778
rect 26516 22714 26568 22720
rect 26528 22098 26556 22714
rect 27632 22098 27660 23054
rect 27712 23044 27764 23050
rect 27712 22986 27764 22992
rect 27724 22234 27752 22986
rect 27712 22228 27764 22234
rect 27712 22170 27764 22176
rect 26516 22092 26568 22098
rect 26516 22034 26568 22040
rect 27620 22092 27672 22098
rect 27620 22034 27672 22040
rect 26240 21956 26292 21962
rect 26240 21898 26292 21904
rect 25964 21548 26016 21554
rect 25964 21490 26016 21496
rect 25596 20596 25648 20602
rect 25596 20538 25648 20544
rect 25964 20392 26016 20398
rect 25964 20334 26016 20340
rect 25504 20324 25556 20330
rect 25504 20266 25556 20272
rect 25136 20256 25188 20262
rect 25136 20198 25188 20204
rect 25516 19922 25544 20266
rect 25976 20058 26004 20334
rect 25964 20052 26016 20058
rect 25964 19994 26016 20000
rect 25136 19916 25188 19922
rect 25136 19858 25188 19864
rect 25412 19916 25464 19922
rect 25412 19858 25464 19864
rect 25504 19916 25556 19922
rect 25504 19858 25556 19864
rect 25148 19310 25176 19858
rect 25424 19310 25452 19858
rect 25516 19310 25544 19858
rect 25976 19718 26004 19994
rect 25964 19712 26016 19718
rect 25964 19654 26016 19660
rect 25136 19304 25188 19310
rect 25042 19272 25098 19281
rect 25136 19246 25188 19252
rect 25412 19304 25464 19310
rect 25412 19246 25464 19252
rect 25504 19304 25556 19310
rect 25504 19246 25556 19252
rect 25042 19207 25098 19216
rect 24860 18896 24912 18902
rect 24860 18838 24912 18844
rect 24860 18760 24912 18766
rect 24860 18702 24912 18708
rect 24676 18216 24728 18222
rect 24676 18158 24728 18164
rect 24688 17746 24716 18158
rect 24676 17740 24728 17746
rect 24676 17682 24728 17688
rect 24872 17082 24900 18702
rect 25148 18222 25176 19246
rect 26056 19236 26108 19242
rect 26056 19178 26108 19184
rect 25228 18828 25280 18834
rect 25228 18770 25280 18776
rect 25136 18216 25188 18222
rect 25136 18158 25188 18164
rect 25148 17746 25176 18158
rect 25136 17740 25188 17746
rect 25136 17682 25188 17688
rect 25240 17542 25268 18770
rect 25504 18692 25556 18698
rect 25504 18634 25556 18640
rect 25516 18222 25544 18634
rect 25320 18216 25372 18222
rect 25320 18158 25372 18164
rect 25504 18216 25556 18222
rect 25504 18158 25556 18164
rect 25332 17746 25360 18158
rect 25516 17746 25544 18158
rect 25780 17876 25832 17882
rect 25780 17818 25832 17824
rect 25320 17740 25372 17746
rect 25320 17682 25372 17688
rect 25504 17740 25556 17746
rect 25504 17682 25556 17688
rect 25228 17536 25280 17542
rect 25228 17478 25280 17484
rect 24780 17054 24900 17082
rect 24780 16998 24808 17054
rect 24768 16992 24820 16998
rect 24768 16934 24820 16940
rect 24952 16992 25004 16998
rect 24952 16934 25004 16940
rect 24964 16726 24992 16934
rect 24952 16720 25004 16726
rect 24952 16662 25004 16668
rect 24860 16652 24912 16658
rect 24860 16594 24912 16600
rect 24676 16584 24728 16590
rect 24674 16552 24676 16561
rect 24728 16552 24730 16561
rect 24674 16487 24730 16496
rect 24676 16448 24728 16454
rect 24676 16390 24728 16396
rect 24688 16046 24716 16390
rect 24676 16040 24728 16046
rect 24676 15982 24728 15988
rect 24676 15428 24728 15434
rect 24676 15370 24728 15376
rect 24504 10798 24624 10826
rect 24400 8628 24452 8634
rect 24400 8570 24452 8576
rect 24412 7342 24440 8570
rect 24400 7336 24452 7342
rect 24400 7278 24452 7284
rect 24308 6452 24360 6458
rect 24308 6394 24360 6400
rect 24216 5772 24268 5778
rect 24216 5714 24268 5720
rect 24124 5704 24176 5710
rect 24124 5646 24176 5652
rect 23940 5160 23992 5166
rect 23940 5102 23992 5108
rect 22836 5092 22888 5098
rect 22836 5034 22888 5040
rect 22848 3602 22876 5034
rect 24228 5030 24256 5714
rect 24308 5160 24360 5166
rect 24308 5102 24360 5108
rect 24216 5024 24268 5030
rect 24216 4966 24268 4972
rect 24320 4826 24348 5102
rect 24308 4820 24360 4826
rect 24308 4762 24360 4768
rect 24504 4010 24532 10798
rect 24584 10668 24636 10674
rect 24584 10610 24636 10616
rect 24596 9722 24624 10610
rect 24688 9926 24716 15370
rect 24872 14074 24900 16594
rect 25044 16584 25096 16590
rect 25044 16526 25096 16532
rect 24952 16040 25004 16046
rect 24952 15982 25004 15988
rect 24964 15570 24992 15982
rect 24952 15564 25004 15570
rect 24952 15506 25004 15512
rect 24964 15094 24992 15506
rect 24952 15088 25004 15094
rect 24952 15030 25004 15036
rect 24952 14476 25004 14482
rect 24952 14418 25004 14424
rect 24860 14068 24912 14074
rect 24860 14010 24912 14016
rect 24768 13728 24820 13734
rect 24768 13670 24820 13676
rect 24780 13462 24808 13670
rect 24964 13462 24992 14418
rect 24768 13456 24820 13462
rect 24768 13398 24820 13404
rect 24952 13456 25004 13462
rect 24952 13398 25004 13404
rect 25056 12730 25084 16526
rect 25136 15972 25188 15978
rect 25136 15914 25188 15920
rect 24964 12702 25084 12730
rect 24964 12374 24992 12702
rect 25044 12640 25096 12646
rect 25044 12582 25096 12588
rect 24952 12368 25004 12374
rect 24952 12310 25004 12316
rect 25056 12306 25084 12582
rect 25044 12300 25096 12306
rect 25044 12242 25096 12248
rect 24952 12096 25004 12102
rect 24952 12038 25004 12044
rect 24964 11694 24992 12038
rect 25148 11694 25176 15914
rect 25240 15706 25268 17478
rect 25688 17264 25740 17270
rect 25688 17206 25740 17212
rect 25700 16998 25728 17206
rect 25688 16992 25740 16998
rect 25688 16934 25740 16940
rect 25318 16688 25374 16697
rect 25792 16658 25820 17818
rect 25318 16623 25320 16632
rect 25372 16623 25374 16632
rect 25780 16652 25832 16658
rect 25320 16594 25372 16600
rect 25780 16594 25832 16600
rect 25502 16008 25558 16017
rect 26068 15978 26096 19178
rect 26252 18834 26280 21898
rect 26516 21480 26568 21486
rect 26516 21422 26568 21428
rect 26332 20256 26384 20262
rect 26332 20198 26384 20204
rect 26344 19310 26372 20198
rect 26528 20058 26556 21422
rect 27632 21010 27660 22034
rect 27724 21554 27752 22170
rect 27816 22098 27844 23122
rect 27908 22574 27936 23190
rect 27896 22568 27948 22574
rect 27896 22510 27948 22516
rect 27908 22234 27936 22510
rect 27988 22432 28040 22438
rect 27988 22374 28040 22380
rect 27896 22228 27948 22234
rect 27896 22170 27948 22176
rect 27804 22092 27856 22098
rect 27804 22034 27856 22040
rect 27712 21548 27764 21554
rect 27712 21490 27764 21496
rect 28000 21486 28028 22374
rect 27988 21480 28040 21486
rect 27988 21422 28040 21428
rect 27620 21004 27672 21010
rect 27620 20946 27672 20952
rect 27712 21004 27764 21010
rect 27712 20946 27764 20952
rect 27620 20868 27672 20874
rect 27620 20810 27672 20816
rect 26700 20596 26752 20602
rect 26700 20538 26752 20544
rect 26516 20052 26568 20058
rect 26516 19994 26568 20000
rect 26608 19916 26660 19922
rect 26608 19858 26660 19864
rect 26332 19304 26384 19310
rect 26332 19246 26384 19252
rect 26240 18828 26292 18834
rect 26240 18770 26292 18776
rect 26148 18760 26200 18766
rect 26148 18702 26200 18708
rect 26160 17134 26188 18702
rect 26148 17128 26200 17134
rect 26146 17096 26148 17105
rect 26240 17128 26292 17134
rect 26200 17096 26202 17105
rect 26240 17070 26292 17076
rect 26146 17031 26202 17040
rect 26252 16833 26280 17070
rect 26238 16824 26294 16833
rect 26238 16759 26294 16768
rect 26344 16674 26372 19246
rect 26516 18216 26568 18222
rect 26516 18158 26568 18164
rect 26424 17672 26476 17678
rect 26424 17614 26476 17620
rect 26252 16646 26372 16674
rect 26148 16040 26200 16046
rect 26148 15982 26200 15988
rect 25502 15943 25558 15952
rect 26056 15972 26108 15978
rect 25228 15700 25280 15706
rect 25228 15642 25280 15648
rect 25412 14816 25464 14822
rect 25412 14758 25464 14764
rect 25320 12640 25372 12646
rect 25320 12582 25372 12588
rect 25332 12442 25360 12582
rect 25320 12436 25372 12442
rect 25320 12378 25372 12384
rect 24952 11688 25004 11694
rect 24952 11630 25004 11636
rect 25136 11688 25188 11694
rect 25136 11630 25188 11636
rect 24768 11620 24820 11626
rect 24768 11562 24820 11568
rect 25320 11620 25372 11626
rect 25320 11562 25372 11568
rect 24780 11218 24808 11562
rect 25332 11218 25360 11562
rect 24768 11212 24820 11218
rect 24768 11154 24820 11160
rect 25320 11212 25372 11218
rect 25320 11154 25372 11160
rect 24676 9920 24728 9926
rect 24676 9862 24728 9868
rect 24584 9716 24636 9722
rect 24584 9658 24636 9664
rect 24596 8498 24624 9658
rect 24780 9382 24808 11154
rect 25136 11076 25188 11082
rect 25136 11018 25188 11024
rect 24952 10600 25004 10606
rect 24952 10542 25004 10548
rect 24860 10124 24912 10130
rect 24860 10066 24912 10072
rect 24768 9376 24820 9382
rect 24768 9318 24820 9324
rect 24872 9194 24900 10066
rect 24964 9654 24992 10542
rect 24952 9648 25004 9654
rect 24952 9590 25004 9596
rect 25044 9444 25096 9450
rect 25044 9386 25096 9392
rect 24780 9178 24900 9194
rect 24768 9172 24900 9178
rect 24820 9166 24900 9172
rect 24768 9114 24820 9120
rect 24860 8968 24912 8974
rect 24860 8910 24912 8916
rect 24872 8838 24900 8910
rect 24952 8900 25004 8906
rect 24952 8842 25004 8848
rect 24860 8832 24912 8838
rect 24860 8774 24912 8780
rect 24584 8492 24636 8498
rect 24584 8434 24636 8440
rect 24768 8016 24820 8022
rect 24768 7958 24820 7964
rect 24676 7948 24728 7954
rect 24676 7890 24728 7896
rect 24688 7002 24716 7890
rect 24780 7546 24808 7958
rect 24768 7540 24820 7546
rect 24768 7482 24820 7488
rect 24872 7478 24900 8774
rect 24964 8498 24992 8842
rect 24952 8492 25004 8498
rect 24952 8434 25004 8440
rect 24860 7472 24912 7478
rect 24860 7414 24912 7420
rect 24676 6996 24728 7002
rect 24676 6938 24728 6944
rect 24688 6866 24716 6938
rect 24676 6860 24728 6866
rect 24676 6802 24728 6808
rect 24688 6254 24716 6802
rect 24952 6792 25004 6798
rect 24952 6734 25004 6740
rect 24676 6248 24728 6254
rect 24676 6190 24728 6196
rect 24964 5817 24992 6734
rect 24950 5808 25006 5817
rect 24950 5743 25006 5752
rect 24858 5672 24914 5681
rect 24858 5607 24860 5616
rect 24912 5607 24914 5616
rect 24860 5578 24912 5584
rect 24860 5160 24912 5166
rect 24860 5102 24912 5108
rect 24872 4690 24900 5102
rect 25056 4826 25084 9386
rect 25148 7970 25176 11018
rect 25332 10198 25360 11154
rect 25320 10192 25372 10198
rect 25320 10134 25372 10140
rect 25332 9518 25360 10134
rect 25320 9512 25372 9518
rect 25320 9454 25372 9460
rect 25226 9072 25282 9081
rect 25226 9007 25228 9016
rect 25280 9007 25282 9016
rect 25228 8978 25280 8984
rect 25148 7942 25268 7970
rect 25424 7954 25452 14758
rect 25516 14482 25544 15943
rect 26056 15914 26108 15920
rect 26160 15502 26188 15982
rect 26148 15496 26200 15502
rect 26148 15438 26200 15444
rect 25688 15360 25740 15366
rect 25688 15302 25740 15308
rect 25596 14952 25648 14958
rect 25596 14894 25648 14900
rect 25504 14476 25556 14482
rect 25504 14418 25556 14424
rect 25608 14346 25636 14894
rect 25596 14340 25648 14346
rect 25596 14282 25648 14288
rect 25596 13864 25648 13870
rect 25596 13806 25648 13812
rect 25504 12912 25556 12918
rect 25504 12854 25556 12860
rect 25240 7342 25268 7942
rect 25412 7948 25464 7954
rect 25412 7890 25464 7896
rect 25320 7744 25372 7750
rect 25320 7686 25372 7692
rect 25332 7546 25360 7686
rect 25320 7540 25372 7546
rect 25320 7482 25372 7488
rect 25228 7336 25280 7342
rect 25228 7278 25280 7284
rect 25136 6860 25188 6866
rect 25136 6802 25188 6808
rect 25148 5778 25176 6802
rect 25516 6769 25544 12854
rect 25608 11626 25636 13806
rect 25596 11620 25648 11626
rect 25596 11562 25648 11568
rect 25608 10674 25636 11562
rect 25700 11098 25728 15302
rect 26056 14816 26108 14822
rect 26056 14758 26108 14764
rect 25964 14408 26016 14414
rect 25964 14350 26016 14356
rect 25870 13424 25926 13433
rect 25870 13359 25926 13368
rect 25884 12918 25912 13359
rect 25872 12912 25924 12918
rect 25872 12854 25924 12860
rect 25872 12776 25924 12782
rect 25976 12764 26004 14350
rect 26068 13938 26096 14758
rect 26146 13968 26202 13977
rect 26056 13932 26108 13938
rect 26146 13903 26148 13912
rect 26056 13874 26108 13880
rect 26200 13903 26202 13912
rect 26148 13874 26200 13880
rect 26252 13394 26280 16646
rect 26436 16182 26464 17614
rect 26528 17338 26556 18158
rect 26620 17610 26648 19858
rect 26712 18970 26740 20538
rect 27632 20466 27660 20810
rect 27620 20460 27672 20466
rect 27540 20398 27568 20429
rect 27620 20402 27672 20408
rect 27528 20392 27580 20398
rect 27724 20346 27752 20946
rect 28184 20534 28212 30738
rect 28644 29510 28672 31062
rect 28736 30122 28764 32014
rect 28828 31210 28856 32302
rect 29564 31822 29592 32914
rect 30196 32360 30248 32366
rect 30196 32302 30248 32308
rect 30012 31884 30064 31890
rect 30012 31826 30064 31832
rect 29460 31816 29512 31822
rect 29460 31758 29512 31764
rect 29552 31816 29604 31822
rect 29552 31758 29604 31764
rect 29472 31278 29500 31758
rect 29000 31272 29052 31278
rect 29000 31214 29052 31220
rect 29460 31272 29512 31278
rect 29460 31214 29512 31220
rect 28816 31204 28868 31210
rect 28816 31146 28868 31152
rect 28908 31136 28960 31142
rect 28908 31078 28960 31084
rect 28724 30116 28776 30122
rect 28724 30058 28776 30064
rect 28632 29504 28684 29510
rect 28632 29446 28684 29452
rect 28644 26994 28672 29446
rect 28736 28626 28764 30058
rect 28920 29102 28948 31078
rect 29012 30598 29040 31214
rect 29000 30592 29052 30598
rect 29000 30534 29052 30540
rect 29276 30592 29328 30598
rect 29276 30534 29328 30540
rect 29288 29782 29316 30534
rect 29472 30258 29500 31214
rect 29460 30252 29512 30258
rect 29460 30194 29512 30200
rect 29276 29776 29328 29782
rect 29276 29718 29328 29724
rect 29368 29708 29420 29714
rect 29368 29650 29420 29656
rect 28908 29096 28960 29102
rect 28908 29038 28960 29044
rect 29276 29028 29328 29034
rect 29276 28970 29328 28976
rect 28724 28620 28776 28626
rect 28724 28562 28776 28568
rect 29288 27130 29316 28970
rect 29380 27946 29408 29650
rect 29564 29102 29592 31758
rect 30024 30734 30052 31826
rect 30012 30728 30064 30734
rect 30012 30670 30064 30676
rect 30024 30190 30052 30670
rect 30012 30184 30064 30190
rect 30012 30126 30064 30132
rect 30024 29714 30052 30126
rect 30012 29708 30064 29714
rect 30012 29650 30064 29656
rect 29552 29096 29604 29102
rect 29552 29038 29604 29044
rect 29644 28416 29696 28422
rect 29644 28358 29696 28364
rect 29656 28014 29684 28358
rect 29644 28008 29696 28014
rect 29644 27950 29696 27956
rect 29368 27940 29420 27946
rect 29368 27882 29420 27888
rect 29380 27606 29408 27882
rect 29368 27600 29420 27606
rect 29368 27542 29420 27548
rect 29276 27124 29328 27130
rect 29276 27066 29328 27072
rect 28632 26988 28684 26994
rect 28632 26930 28684 26936
rect 28540 26920 28592 26926
rect 28540 26862 28592 26868
rect 29552 26920 29604 26926
rect 29656 26908 29684 27950
rect 30024 27130 30052 29650
rect 30012 27124 30064 27130
rect 30012 27066 30064 27072
rect 29604 26880 29684 26908
rect 29552 26862 29604 26868
rect 28264 24744 28316 24750
rect 28264 24686 28316 24692
rect 28276 23186 28304 24686
rect 28552 24410 28580 26862
rect 30104 26784 30156 26790
rect 30104 26726 30156 26732
rect 29276 26376 29328 26382
rect 29276 26318 29328 26324
rect 29184 26240 29236 26246
rect 29184 26182 29236 26188
rect 29196 25838 29224 26182
rect 29184 25832 29236 25838
rect 29184 25774 29236 25780
rect 28632 25696 28684 25702
rect 28632 25638 28684 25644
rect 28644 24750 28672 25638
rect 28908 25356 28960 25362
rect 28908 25298 28960 25304
rect 28632 24744 28684 24750
rect 28632 24686 28684 24692
rect 28540 24404 28592 24410
rect 28540 24346 28592 24352
rect 28356 23588 28408 23594
rect 28356 23530 28408 23536
rect 28368 23202 28396 23530
rect 28552 23254 28580 24346
rect 28540 23248 28592 23254
rect 28368 23186 28488 23202
rect 28540 23190 28592 23196
rect 28264 23180 28316 23186
rect 28264 23122 28316 23128
rect 28368 23180 28500 23186
rect 28368 23174 28448 23180
rect 28368 22642 28396 23174
rect 28448 23122 28500 23128
rect 28356 22636 28408 22642
rect 28356 22578 28408 22584
rect 28644 22574 28672 24686
rect 28920 24342 28948 25298
rect 29000 25152 29052 25158
rect 29000 25094 29052 25100
rect 28908 24336 28960 24342
rect 28908 24278 28960 24284
rect 28920 23186 28948 24278
rect 28908 23180 28960 23186
rect 28908 23122 28960 23128
rect 28724 22772 28776 22778
rect 28724 22714 28776 22720
rect 28632 22568 28684 22574
rect 28632 22510 28684 22516
rect 28644 21622 28672 22510
rect 28736 22030 28764 22714
rect 29012 22506 29040 25094
rect 29196 24818 29224 25774
rect 29288 25430 29316 26318
rect 30116 26314 30144 26726
rect 29644 26308 29696 26314
rect 29644 26250 29696 26256
rect 30104 26308 30156 26314
rect 30104 26250 30156 26256
rect 29656 25906 29684 26250
rect 29736 26240 29788 26246
rect 29736 26182 29788 26188
rect 29644 25900 29696 25906
rect 29644 25842 29696 25848
rect 29748 25786 29776 26182
rect 29656 25758 29776 25786
rect 29656 25702 29684 25758
rect 29644 25696 29696 25702
rect 29644 25638 29696 25644
rect 29276 25424 29328 25430
rect 29276 25366 29328 25372
rect 29184 24812 29236 24818
rect 29184 24754 29236 24760
rect 29196 24274 29224 24754
rect 29184 24268 29236 24274
rect 29104 24228 29184 24256
rect 29104 23118 29132 24228
rect 29184 24210 29236 24216
rect 29368 24200 29420 24206
rect 29368 24142 29420 24148
rect 29274 23624 29330 23633
rect 29274 23559 29330 23568
rect 29092 23112 29144 23118
rect 29092 23054 29144 23060
rect 29288 23050 29316 23559
rect 29380 23322 29408 24142
rect 29656 23594 29684 25638
rect 29920 25356 29972 25362
rect 29920 25298 29972 25304
rect 29932 24886 29960 25298
rect 30012 25288 30064 25294
rect 30012 25230 30064 25236
rect 29920 24880 29972 24886
rect 29920 24822 29972 24828
rect 29932 24206 29960 24822
rect 30024 24342 30052 25230
rect 30012 24336 30064 24342
rect 30012 24278 30064 24284
rect 29920 24200 29972 24206
rect 29920 24142 29972 24148
rect 29644 23588 29696 23594
rect 29644 23530 29696 23536
rect 29368 23316 29420 23322
rect 29368 23258 29420 23264
rect 29276 23044 29328 23050
rect 29276 22986 29328 22992
rect 29552 23044 29604 23050
rect 29552 22986 29604 22992
rect 29460 22976 29512 22982
rect 29460 22918 29512 22924
rect 29472 22574 29500 22918
rect 29460 22568 29512 22574
rect 29460 22510 29512 22516
rect 29000 22500 29052 22506
rect 29000 22442 29052 22448
rect 29012 22148 29040 22442
rect 29564 22438 29592 22986
rect 29552 22432 29604 22438
rect 29552 22374 29604 22380
rect 29092 22160 29144 22166
rect 29012 22120 29092 22148
rect 29144 22120 29224 22148
rect 29092 22102 29144 22108
rect 28724 22024 28776 22030
rect 29092 22024 29144 22030
rect 28724 21966 28776 21972
rect 29090 21992 29092 22001
rect 29144 21992 29146 22001
rect 29090 21927 29146 21936
rect 29092 21888 29144 21894
rect 29092 21830 29144 21836
rect 29104 21690 29132 21830
rect 29000 21684 29052 21690
rect 29000 21626 29052 21632
rect 29092 21684 29144 21690
rect 29092 21626 29144 21632
rect 28632 21616 28684 21622
rect 28632 21558 28684 21564
rect 28632 21480 28684 21486
rect 28632 21422 28684 21428
rect 28644 21146 28672 21422
rect 29012 21162 29040 21626
rect 29196 21486 29224 22120
rect 29656 22098 29684 23530
rect 29920 23180 29972 23186
rect 29920 23122 29972 23128
rect 29828 23112 29880 23118
rect 29828 23054 29880 23060
rect 29840 22778 29868 23054
rect 29828 22772 29880 22778
rect 29828 22714 29880 22720
rect 29828 22500 29880 22506
rect 29828 22442 29880 22448
rect 29644 22092 29696 22098
rect 29644 22034 29696 22040
rect 29840 21536 29868 22442
rect 29932 21604 29960 23122
rect 30024 22982 30052 24278
rect 30012 22976 30064 22982
rect 30012 22918 30064 22924
rect 30012 22432 30064 22438
rect 30012 22374 30064 22380
rect 30024 22098 30052 22374
rect 30012 22092 30064 22098
rect 30012 22034 30064 22040
rect 29932 21576 30052 21604
rect 29840 21508 29960 21536
rect 29184 21480 29236 21486
rect 29184 21422 29236 21428
rect 29828 21412 29880 21418
rect 29828 21354 29880 21360
rect 29276 21344 29328 21350
rect 29276 21286 29328 21292
rect 28632 21140 28684 21146
rect 29012 21134 29224 21162
rect 28632 21082 28684 21088
rect 29092 21072 29144 21078
rect 29092 21014 29144 21020
rect 28356 21004 28408 21010
rect 28356 20946 28408 20952
rect 28172 20528 28224 20534
rect 28172 20470 28224 20476
rect 27580 20340 27752 20346
rect 27528 20334 27752 20340
rect 27540 20318 27752 20334
rect 27436 20052 27488 20058
rect 27436 19994 27488 20000
rect 27448 19961 27476 19994
rect 27434 19952 27490 19961
rect 27434 19887 27436 19896
rect 27488 19887 27490 19896
rect 27436 19858 27488 19864
rect 27068 19712 27120 19718
rect 27068 19654 27120 19660
rect 27080 19514 27108 19654
rect 27068 19508 27120 19514
rect 27068 19450 27120 19456
rect 27080 19310 27108 19450
rect 27068 19304 27120 19310
rect 27068 19246 27120 19252
rect 27160 19304 27212 19310
rect 27160 19246 27212 19252
rect 26700 18964 26752 18970
rect 26700 18906 26752 18912
rect 26608 17604 26660 17610
rect 26608 17546 26660 17552
rect 26516 17332 26568 17338
rect 26516 17274 26568 17280
rect 26608 16584 26660 16590
rect 26608 16526 26660 16532
rect 26516 16244 26568 16250
rect 26516 16186 26568 16192
rect 26424 16176 26476 16182
rect 26424 16118 26476 16124
rect 26332 16040 26384 16046
rect 26332 15982 26384 15988
rect 26240 13388 26292 13394
rect 26240 13330 26292 13336
rect 26056 12980 26108 12986
rect 26056 12922 26108 12928
rect 25924 12736 26004 12764
rect 25872 12718 25924 12724
rect 25700 11070 25820 11098
rect 25688 11008 25740 11014
rect 25688 10950 25740 10956
rect 25596 10668 25648 10674
rect 25596 10610 25648 10616
rect 25700 10130 25728 10950
rect 25688 10124 25740 10130
rect 25688 10066 25740 10072
rect 25792 7342 25820 11070
rect 25884 8838 25912 12718
rect 26068 12442 26096 12922
rect 26056 12436 26108 12442
rect 26056 12378 26108 12384
rect 26056 12300 26108 12306
rect 26056 12242 26108 12248
rect 26068 10538 26096 12242
rect 26344 11898 26372 15982
rect 26424 14952 26476 14958
rect 26424 14894 26476 14900
rect 26436 14550 26464 14894
rect 26424 14544 26476 14550
rect 26424 14486 26476 14492
rect 26528 12782 26556 16186
rect 26620 15706 26648 16526
rect 26608 15700 26660 15706
rect 26608 15642 26660 15648
rect 26608 14952 26660 14958
rect 26608 14894 26660 14900
rect 26620 14618 26648 14894
rect 26608 14612 26660 14618
rect 26608 14554 26660 14560
rect 26712 14482 26740 18906
rect 27172 18290 27200 19246
rect 27344 18624 27396 18630
rect 27344 18566 27396 18572
rect 27436 18624 27488 18630
rect 27436 18566 27488 18572
rect 27160 18284 27212 18290
rect 27160 18226 27212 18232
rect 27356 18222 27384 18566
rect 27344 18216 27396 18222
rect 27344 18158 27396 18164
rect 26792 17740 26844 17746
rect 26792 17682 26844 17688
rect 26976 17740 27028 17746
rect 26976 17682 27028 17688
rect 26804 17202 26832 17682
rect 26792 17196 26844 17202
rect 26792 17138 26844 17144
rect 26804 16658 26832 17138
rect 26792 16652 26844 16658
rect 26792 16594 26844 16600
rect 26884 15564 26936 15570
rect 26884 15506 26936 15512
rect 26896 14958 26924 15506
rect 26884 14952 26936 14958
rect 26884 14894 26936 14900
rect 26700 14476 26752 14482
rect 26700 14418 26752 14424
rect 26608 13320 26660 13326
rect 26608 13262 26660 13268
rect 26516 12776 26568 12782
rect 26516 12718 26568 12724
rect 26516 12300 26568 12306
rect 26516 12242 26568 12248
rect 26332 11892 26384 11898
rect 26332 11834 26384 11840
rect 26056 10532 26108 10538
rect 26056 10474 26108 10480
rect 25872 8832 25924 8838
rect 25872 8774 25924 8780
rect 25872 8288 25924 8294
rect 25872 8230 25924 8236
rect 25884 8090 25912 8230
rect 25872 8084 25924 8090
rect 25872 8026 25924 8032
rect 25780 7336 25832 7342
rect 25780 7278 25832 7284
rect 25792 6934 25820 7278
rect 25780 6928 25832 6934
rect 25780 6870 25832 6876
rect 25884 6798 25912 8026
rect 25872 6792 25924 6798
rect 25502 6760 25558 6769
rect 25872 6734 25924 6740
rect 25502 6695 25558 6704
rect 25884 5914 25912 6734
rect 26068 6662 26096 10474
rect 26148 10464 26200 10470
rect 26148 10406 26200 10412
rect 26056 6656 26108 6662
rect 26056 6598 26108 6604
rect 26068 6458 26096 6598
rect 26056 6452 26108 6458
rect 26056 6394 26108 6400
rect 25872 5908 25924 5914
rect 25872 5850 25924 5856
rect 25136 5772 25188 5778
rect 25136 5714 25188 5720
rect 25044 4820 25096 4826
rect 25044 4762 25096 4768
rect 26160 4690 26188 10406
rect 26240 9648 26292 9654
rect 26240 9590 26292 9596
rect 26252 9178 26280 9590
rect 26528 9489 26556 12242
rect 26620 11218 26648 13262
rect 26712 12782 26740 14418
rect 26882 13832 26938 13841
rect 26882 13767 26938 13776
rect 26700 12776 26752 12782
rect 26700 12718 26752 12724
rect 26700 11552 26752 11558
rect 26700 11494 26752 11500
rect 26712 11286 26740 11494
rect 26700 11280 26752 11286
rect 26700 11222 26752 11228
rect 26608 11212 26660 11218
rect 26608 11154 26660 11160
rect 26514 9480 26570 9489
rect 26332 9444 26384 9450
rect 26514 9415 26570 9424
rect 26332 9386 26384 9392
rect 26240 9172 26292 9178
rect 26240 9114 26292 9120
rect 26240 9036 26292 9042
rect 26240 8978 26292 8984
rect 26252 8634 26280 8978
rect 26240 8628 26292 8634
rect 26240 8570 26292 8576
rect 26344 8430 26372 9386
rect 26528 9382 26556 9415
rect 26516 9376 26568 9382
rect 26516 9318 26568 9324
rect 26896 9178 26924 13767
rect 26884 9172 26936 9178
rect 26884 9114 26936 9120
rect 26332 8424 26384 8430
rect 26332 8366 26384 8372
rect 26332 7336 26384 7342
rect 26332 7278 26384 7284
rect 26344 6866 26372 7278
rect 26332 6860 26384 6866
rect 26332 6802 26384 6808
rect 26344 6662 26372 6802
rect 26332 6656 26384 6662
rect 26332 6598 26384 6604
rect 26344 5778 26372 6598
rect 26988 6322 27016 17682
rect 27068 17604 27120 17610
rect 27068 17546 27120 17552
rect 27080 16658 27108 17546
rect 27448 17066 27476 18566
rect 27540 17338 27568 20318
rect 27620 19848 27672 19854
rect 27620 19790 27672 19796
rect 27632 19174 27660 19790
rect 27712 19712 27764 19718
rect 27712 19654 27764 19660
rect 27620 19168 27672 19174
rect 27620 19110 27672 19116
rect 27724 18952 27752 19654
rect 28080 19168 28132 19174
rect 28080 19110 28132 19116
rect 27896 18964 27948 18970
rect 27724 18924 27896 18952
rect 27724 17610 27752 18924
rect 27896 18906 27948 18912
rect 28092 18834 28120 19110
rect 28080 18828 28132 18834
rect 28080 18770 28132 18776
rect 27988 18080 28040 18086
rect 27988 18022 28040 18028
rect 27712 17604 27764 17610
rect 27712 17546 27764 17552
rect 27528 17332 27580 17338
rect 27528 17274 27580 17280
rect 27540 17134 27568 17274
rect 28000 17134 28028 18022
rect 28092 17134 28120 18770
rect 28368 18306 28396 20946
rect 28448 20392 28500 20398
rect 28448 20334 28500 20340
rect 28540 20392 28592 20398
rect 28540 20334 28592 20340
rect 28460 19378 28488 20334
rect 28552 19922 28580 20334
rect 28540 19916 28592 19922
rect 28540 19858 28592 19864
rect 29000 19916 29052 19922
rect 29000 19858 29052 19864
rect 28540 19508 28592 19514
rect 28540 19450 28592 19456
rect 28448 19372 28500 19378
rect 28448 19314 28500 19320
rect 28552 18834 28580 19450
rect 29012 19310 29040 19858
rect 29104 19854 29132 21014
rect 29092 19848 29144 19854
rect 29092 19790 29144 19796
rect 29000 19304 29052 19310
rect 29000 19246 29052 19252
rect 28540 18828 28592 18834
rect 28540 18770 28592 18776
rect 29092 18760 29144 18766
rect 29092 18702 29144 18708
rect 28184 18278 28396 18306
rect 27528 17128 27580 17134
rect 27528 17070 27580 17076
rect 27988 17128 28040 17134
rect 28080 17128 28132 17134
rect 27988 17070 28040 17076
rect 28078 17096 28080 17105
rect 28132 17096 28134 17105
rect 27436 17060 27488 17066
rect 27436 17002 27488 17008
rect 27712 17060 27764 17066
rect 28078 17031 28134 17040
rect 27712 17002 27764 17008
rect 27448 16658 27476 17002
rect 27528 16992 27580 16998
rect 27580 16940 27660 16946
rect 27528 16934 27660 16940
rect 27540 16918 27660 16934
rect 27632 16658 27660 16918
rect 27068 16652 27120 16658
rect 27068 16594 27120 16600
rect 27436 16652 27488 16658
rect 27436 16594 27488 16600
rect 27620 16652 27672 16658
rect 27620 16594 27672 16600
rect 27080 14346 27108 16594
rect 27160 16516 27212 16522
rect 27160 16458 27212 16464
rect 27172 15570 27200 16458
rect 27342 16144 27398 16153
rect 27342 16079 27344 16088
rect 27396 16079 27398 16088
rect 27344 16050 27396 16056
rect 27252 15972 27304 15978
rect 27252 15914 27304 15920
rect 27160 15564 27212 15570
rect 27160 15506 27212 15512
rect 27068 14340 27120 14346
rect 27068 14282 27120 14288
rect 27160 12300 27212 12306
rect 27160 12242 27212 12248
rect 27172 11898 27200 12242
rect 27160 11892 27212 11898
rect 27160 11834 27212 11840
rect 27264 11014 27292 15914
rect 27436 15428 27488 15434
rect 27436 15370 27488 15376
rect 27448 13394 27476 15370
rect 27528 14952 27580 14958
rect 27528 14894 27580 14900
rect 27540 14074 27568 14894
rect 27620 14408 27672 14414
rect 27620 14350 27672 14356
rect 27528 14068 27580 14074
rect 27528 14010 27580 14016
rect 27528 13728 27580 13734
rect 27528 13670 27580 13676
rect 27436 13388 27488 13394
rect 27436 13330 27488 13336
rect 27540 12646 27568 13670
rect 27632 12850 27660 14350
rect 27620 12844 27672 12850
rect 27620 12786 27672 12792
rect 27528 12640 27580 12646
rect 27528 12582 27580 12588
rect 27540 12306 27568 12582
rect 27528 12300 27580 12306
rect 27528 12242 27580 12248
rect 27620 11688 27672 11694
rect 27620 11630 27672 11636
rect 27344 11212 27396 11218
rect 27344 11154 27396 11160
rect 27252 11008 27304 11014
rect 27252 10950 27304 10956
rect 27068 10600 27120 10606
rect 27068 10542 27120 10548
rect 27160 10600 27212 10606
rect 27160 10542 27212 10548
rect 27080 9654 27108 10542
rect 27172 10266 27200 10542
rect 27160 10260 27212 10266
rect 27160 10202 27212 10208
rect 27172 10062 27200 10202
rect 27264 10198 27292 10950
rect 27356 10470 27384 11154
rect 27526 10704 27582 10713
rect 27526 10639 27582 10648
rect 27540 10606 27568 10639
rect 27528 10600 27580 10606
rect 27448 10560 27528 10588
rect 27344 10464 27396 10470
rect 27344 10406 27396 10412
rect 27252 10192 27304 10198
rect 27252 10134 27304 10140
rect 27160 10056 27212 10062
rect 27160 9998 27212 10004
rect 27448 9722 27476 10560
rect 27528 10542 27580 10548
rect 27632 10452 27660 11630
rect 27724 11014 27752 17002
rect 28184 16658 28212 18278
rect 28632 18216 28684 18222
rect 28632 18158 28684 18164
rect 28644 17746 28672 18158
rect 29104 18154 29132 18702
rect 29092 18148 29144 18154
rect 29092 18090 29144 18096
rect 28724 18080 28776 18086
rect 28724 18022 28776 18028
rect 28632 17740 28684 17746
rect 28632 17682 28684 17688
rect 28356 17332 28408 17338
rect 28356 17274 28408 17280
rect 28368 16658 28396 17274
rect 28448 17128 28500 17134
rect 28448 17070 28500 17076
rect 28172 16652 28224 16658
rect 28172 16594 28224 16600
rect 28356 16652 28408 16658
rect 28356 16594 28408 16600
rect 28184 16538 28212 16594
rect 28092 16510 28212 16538
rect 27804 16040 27856 16046
rect 27804 15982 27856 15988
rect 27816 15434 27844 15982
rect 27896 15564 27948 15570
rect 27896 15506 27948 15512
rect 27804 15428 27856 15434
rect 27804 15370 27856 15376
rect 27908 15094 27936 15506
rect 27988 15496 28040 15502
rect 27988 15438 28040 15444
rect 27896 15088 27948 15094
rect 27896 15030 27948 15036
rect 27894 14512 27950 14521
rect 27816 14456 27894 14464
rect 27816 14436 27896 14456
rect 27712 11008 27764 11014
rect 27712 10950 27764 10956
rect 27712 10464 27764 10470
rect 27632 10424 27712 10452
rect 27632 10266 27660 10424
rect 27712 10406 27764 10412
rect 27620 10260 27672 10266
rect 27620 10202 27672 10208
rect 27528 9988 27580 9994
rect 27528 9930 27580 9936
rect 27436 9716 27488 9722
rect 27436 9658 27488 9664
rect 27068 9648 27120 9654
rect 27068 9590 27120 9596
rect 27080 9518 27108 9590
rect 27068 9512 27120 9518
rect 27540 9500 27568 9930
rect 27620 9512 27672 9518
rect 27068 9454 27120 9460
rect 27448 9472 27620 9500
rect 27080 7954 27108 9454
rect 27448 8974 27476 9472
rect 27620 9454 27672 9460
rect 27436 8968 27488 8974
rect 27436 8910 27488 8916
rect 27448 7954 27476 8910
rect 27712 8424 27764 8430
rect 27712 8366 27764 8372
rect 27724 8090 27752 8366
rect 27528 8084 27580 8090
rect 27712 8084 27764 8090
rect 27580 8044 27660 8072
rect 27528 8026 27580 8032
rect 27632 7970 27660 8044
rect 27712 8026 27764 8032
rect 27816 7970 27844 14436
rect 27948 14447 27950 14456
rect 27896 14418 27948 14424
rect 28000 12918 28028 15438
rect 28092 13190 28120 16510
rect 28172 16448 28224 16454
rect 28172 16390 28224 16396
rect 28184 14958 28212 16390
rect 28354 16144 28410 16153
rect 28354 16079 28356 16088
rect 28408 16079 28410 16088
rect 28356 16050 28408 16056
rect 28172 14952 28224 14958
rect 28172 14894 28224 14900
rect 28460 14414 28488 17070
rect 28736 16436 28764 18022
rect 28816 17740 28868 17746
rect 28816 17682 28868 17688
rect 28828 17202 28856 17682
rect 29104 17678 29132 18090
rect 29092 17672 29144 17678
rect 29092 17614 29144 17620
rect 28816 17196 28868 17202
rect 28816 17138 28868 17144
rect 28828 16658 28856 17138
rect 28906 16824 28962 16833
rect 29000 16788 29052 16794
rect 28962 16768 29000 16776
rect 28906 16759 29000 16768
rect 28920 16748 29000 16759
rect 29000 16730 29052 16736
rect 29104 16658 29132 17614
rect 28816 16652 28868 16658
rect 29092 16652 29144 16658
rect 28868 16612 29040 16640
rect 28816 16594 28868 16600
rect 28908 16448 28960 16454
rect 28736 16408 28908 16436
rect 28724 14884 28776 14890
rect 28724 14826 28776 14832
rect 28448 14408 28500 14414
rect 28448 14350 28500 14356
rect 28448 13864 28500 13870
rect 28448 13806 28500 13812
rect 28460 13530 28488 13806
rect 28448 13524 28500 13530
rect 28448 13466 28500 13472
rect 28080 13184 28132 13190
rect 28080 13126 28132 13132
rect 27988 12912 28040 12918
rect 27988 12854 28040 12860
rect 28460 12782 28488 13466
rect 28448 12776 28500 12782
rect 28448 12718 28500 12724
rect 28632 12708 28684 12714
rect 28632 12650 28684 12656
rect 28540 11688 28592 11694
rect 28540 11630 28592 11636
rect 28552 11082 28580 11630
rect 28540 11076 28592 11082
rect 28540 11018 28592 11024
rect 27896 11008 27948 11014
rect 27896 10950 27948 10956
rect 28080 11008 28132 11014
rect 28080 10950 28132 10956
rect 27908 10062 27936 10950
rect 28092 10810 28120 10950
rect 28080 10804 28132 10810
rect 28080 10746 28132 10752
rect 28080 10668 28132 10674
rect 28080 10610 28132 10616
rect 27988 10600 28040 10606
rect 27988 10542 28040 10548
rect 28000 10146 28028 10542
rect 28092 10538 28120 10610
rect 28644 10606 28672 12650
rect 28736 12442 28764 14826
rect 28828 14618 28856 16408
rect 28908 16390 28960 16396
rect 29012 16250 29040 16612
rect 29092 16594 29144 16600
rect 29000 16244 29052 16250
rect 29000 16186 29052 16192
rect 29196 16046 29224 21134
rect 29288 21010 29316 21286
rect 29840 21010 29868 21354
rect 29276 21004 29328 21010
rect 29276 20946 29328 20952
rect 29828 21004 29880 21010
rect 29828 20946 29880 20952
rect 29288 18426 29316 20946
rect 29736 20256 29788 20262
rect 29736 20198 29788 20204
rect 29644 19712 29696 19718
rect 29644 19654 29696 19660
rect 29460 19372 29512 19378
rect 29460 19314 29512 19320
rect 29368 18692 29420 18698
rect 29368 18634 29420 18640
rect 29276 18420 29328 18426
rect 29276 18362 29328 18368
rect 29288 18222 29316 18362
rect 29276 18216 29328 18222
rect 29276 18158 29328 18164
rect 29380 18068 29408 18634
rect 29472 18358 29500 19314
rect 29656 19174 29684 19654
rect 29644 19168 29696 19174
rect 29644 19110 29696 19116
rect 29552 18760 29604 18766
rect 29552 18702 29604 18708
rect 29460 18352 29512 18358
rect 29460 18294 29512 18300
rect 29564 18222 29592 18702
rect 29552 18216 29604 18222
rect 29552 18158 29604 18164
rect 29288 18040 29408 18068
rect 29288 16114 29316 18040
rect 29552 17128 29604 17134
rect 29656 17116 29684 19110
rect 29748 18834 29776 20198
rect 29828 19712 29880 19718
rect 29828 19654 29880 19660
rect 29736 18828 29788 18834
rect 29736 18770 29788 18776
rect 29604 17088 29684 17116
rect 29552 17070 29604 17076
rect 29368 16652 29420 16658
rect 29368 16594 29420 16600
rect 29276 16108 29328 16114
rect 29276 16050 29328 16056
rect 29184 16040 29236 16046
rect 29184 15982 29236 15988
rect 29276 15700 29328 15706
rect 29276 15642 29328 15648
rect 28816 14612 28868 14618
rect 28816 14554 28868 14560
rect 29288 14482 29316 15642
rect 29380 15638 29408 16594
rect 29368 15632 29420 15638
rect 29368 15574 29420 15580
rect 29564 15026 29592 17070
rect 29748 16590 29776 18770
rect 29736 16584 29788 16590
rect 29736 16526 29788 16532
rect 29644 15700 29696 15706
rect 29644 15642 29696 15648
rect 29552 15020 29604 15026
rect 29552 14962 29604 14968
rect 29276 14476 29328 14482
rect 29276 14418 29328 14424
rect 29288 14278 29316 14418
rect 29276 14272 29328 14278
rect 29276 14214 29328 14220
rect 29656 13870 29684 15642
rect 29748 15638 29776 16526
rect 29736 15632 29788 15638
rect 29736 15574 29788 15580
rect 29748 14958 29776 15574
rect 29840 15570 29868 19654
rect 29932 16833 29960 21508
rect 30024 21418 30052 21576
rect 30116 21486 30144 26250
rect 30208 22234 30236 32302
rect 30288 31884 30340 31890
rect 30288 31826 30340 31832
rect 30300 30802 30328 31826
rect 30392 30870 30420 32914
rect 30840 32360 30892 32366
rect 30840 32302 30892 32308
rect 30472 31748 30524 31754
rect 30472 31690 30524 31696
rect 30484 31278 30512 31690
rect 30852 31414 30880 32302
rect 30840 31408 30892 31414
rect 30840 31350 30892 31356
rect 30472 31272 30524 31278
rect 30472 31214 30524 31220
rect 30380 30864 30432 30870
rect 30380 30806 30432 30812
rect 30288 30796 30340 30802
rect 30288 30738 30340 30744
rect 30564 30796 30616 30802
rect 30564 30738 30616 30744
rect 30300 30190 30328 30738
rect 30288 30184 30340 30190
rect 30288 30126 30340 30132
rect 30300 29714 30328 30126
rect 30576 29782 30604 30738
rect 30564 29776 30616 29782
rect 30564 29718 30616 29724
rect 30288 29708 30340 29714
rect 30288 29650 30340 29656
rect 30300 28762 30328 29650
rect 30380 29640 30432 29646
rect 30380 29582 30432 29588
rect 30288 28756 30340 28762
rect 30288 28698 30340 28704
rect 30392 28626 30420 29582
rect 30748 29300 30800 29306
rect 30748 29242 30800 29248
rect 30380 28620 30432 28626
rect 30380 28562 30432 28568
rect 30392 28014 30420 28562
rect 30760 28014 30788 29242
rect 30380 28008 30432 28014
rect 30380 27950 30432 27956
rect 30748 28008 30800 28014
rect 30748 27950 30800 27956
rect 30932 28008 30984 28014
rect 30932 27950 30984 27956
rect 30392 27470 30420 27950
rect 30760 27538 30788 27950
rect 30944 27606 30972 27950
rect 30932 27600 30984 27606
rect 30932 27542 30984 27548
rect 30748 27532 30800 27538
rect 30748 27474 30800 27480
rect 30380 27464 30432 27470
rect 30380 27406 30432 27412
rect 30564 26444 30616 26450
rect 30564 26386 30616 26392
rect 30380 25764 30432 25770
rect 30380 25706 30432 25712
rect 30392 25294 30420 25706
rect 30380 25288 30432 25294
rect 30380 25230 30432 25236
rect 30576 25226 30604 26386
rect 30564 25220 30616 25226
rect 30564 25162 30616 25168
rect 30656 24744 30708 24750
rect 30656 24686 30708 24692
rect 30564 24676 30616 24682
rect 30564 24618 30616 24624
rect 30472 24608 30524 24614
rect 30472 24550 30524 24556
rect 30484 24274 30512 24550
rect 30472 24268 30524 24274
rect 30472 24210 30524 24216
rect 30484 23662 30512 24210
rect 30576 23730 30604 24618
rect 30668 24274 30696 24686
rect 30656 24268 30708 24274
rect 30656 24210 30708 24216
rect 30668 23798 30696 24210
rect 30656 23792 30708 23798
rect 30656 23734 30708 23740
rect 30564 23724 30616 23730
rect 30564 23666 30616 23672
rect 30472 23656 30524 23662
rect 30472 23598 30524 23604
rect 30576 22778 30604 23666
rect 30668 23186 30696 23734
rect 30656 23180 30708 23186
rect 30656 23122 30708 23128
rect 30564 22772 30616 22778
rect 30564 22714 30616 22720
rect 30196 22228 30248 22234
rect 30196 22170 30248 22176
rect 30288 21548 30340 21554
rect 30288 21490 30340 21496
rect 30104 21480 30156 21486
rect 30104 21422 30156 21428
rect 30012 21412 30064 21418
rect 30012 21354 30064 21360
rect 30024 20058 30052 21354
rect 30300 21010 30328 21490
rect 30564 21480 30616 21486
rect 30564 21422 30616 21428
rect 30288 21004 30340 21010
rect 30288 20946 30340 20952
rect 30288 20392 30340 20398
rect 30288 20334 30340 20340
rect 30012 20052 30064 20058
rect 30012 19994 30064 20000
rect 30012 19304 30064 19310
rect 30300 19292 30328 20334
rect 30064 19264 30328 19292
rect 30012 19246 30064 19252
rect 30024 17678 30052 19246
rect 30196 18828 30248 18834
rect 30196 18770 30248 18776
rect 30208 18290 30236 18770
rect 30196 18284 30248 18290
rect 30196 18226 30248 18232
rect 30208 17814 30236 18226
rect 30288 18080 30340 18086
rect 30288 18022 30340 18028
rect 30196 17808 30248 17814
rect 30196 17750 30248 17756
rect 30012 17672 30064 17678
rect 30012 17614 30064 17620
rect 30196 17672 30248 17678
rect 30196 17614 30248 17620
rect 30012 17128 30064 17134
rect 30012 17070 30064 17076
rect 29918 16824 29974 16833
rect 29918 16759 29974 16768
rect 29932 15706 29960 16759
rect 30024 16522 30052 17070
rect 30208 16538 30236 17614
rect 30300 17134 30328 18022
rect 30288 17128 30340 17134
rect 30288 17070 30340 17076
rect 30380 16992 30432 16998
rect 30380 16934 30432 16940
rect 30392 16658 30420 16934
rect 30380 16652 30432 16658
rect 30380 16594 30432 16600
rect 30472 16584 30524 16590
rect 30012 16516 30064 16522
rect 30208 16510 30420 16538
rect 30472 16526 30524 16532
rect 30012 16458 30064 16464
rect 30024 15706 30052 16458
rect 30196 16244 30248 16250
rect 30196 16186 30248 16192
rect 29920 15700 29972 15706
rect 29920 15642 29972 15648
rect 30012 15700 30064 15706
rect 30012 15642 30064 15648
rect 30208 15570 30236 16186
rect 30288 16040 30340 16046
rect 30288 15982 30340 15988
rect 30392 15994 30420 16510
rect 30484 16114 30512 16526
rect 30472 16108 30524 16114
rect 30472 16050 30524 16056
rect 29828 15564 29880 15570
rect 29828 15506 29880 15512
rect 30196 15564 30248 15570
rect 30196 15506 30248 15512
rect 29840 14958 29868 15506
rect 30300 14958 30328 15982
rect 30392 15966 30512 15994
rect 29736 14952 29788 14958
rect 29736 14894 29788 14900
rect 29828 14952 29880 14958
rect 30288 14952 30340 14958
rect 29828 14894 29880 14900
rect 30208 14900 30288 14906
rect 30208 14894 30340 14900
rect 29840 14634 29868 14894
rect 30208 14878 30328 14894
rect 29840 14606 29960 14634
rect 29932 14482 29960 14606
rect 29828 14476 29880 14482
rect 29828 14418 29880 14424
rect 29920 14476 29972 14482
rect 29920 14418 29972 14424
rect 29736 14408 29788 14414
rect 29736 14350 29788 14356
rect 29748 13870 29776 14350
rect 29840 13938 29868 14418
rect 30208 14414 30236 14878
rect 30288 14816 30340 14822
rect 30288 14758 30340 14764
rect 30196 14408 30248 14414
rect 30196 14350 30248 14356
rect 29828 13932 29880 13938
rect 29828 13874 29880 13880
rect 29644 13864 29696 13870
rect 29644 13806 29696 13812
rect 29736 13864 29788 13870
rect 29736 13806 29788 13812
rect 29656 13394 29684 13806
rect 29092 13388 29144 13394
rect 29092 13330 29144 13336
rect 29644 13388 29696 13394
rect 29644 13330 29696 13336
rect 28724 12436 28776 12442
rect 28724 12378 28776 12384
rect 29104 12102 29132 13330
rect 29748 13326 29776 13806
rect 30300 13326 30328 14758
rect 30380 14068 30432 14074
rect 30380 14010 30432 14016
rect 29736 13320 29788 13326
rect 29736 13262 29788 13268
rect 30196 13320 30248 13326
rect 30196 13262 30248 13268
rect 30288 13320 30340 13326
rect 30288 13262 30340 13268
rect 29748 12442 29776 13262
rect 30208 12986 30236 13262
rect 30196 12980 30248 12986
rect 30196 12922 30248 12928
rect 30300 12850 30328 13262
rect 30288 12844 30340 12850
rect 30288 12786 30340 12792
rect 29920 12776 29972 12782
rect 29920 12718 29972 12724
rect 29736 12436 29788 12442
rect 29736 12378 29788 12384
rect 29092 12096 29144 12102
rect 29092 12038 29144 12044
rect 28908 11756 28960 11762
rect 28908 11698 28960 11704
rect 28632 10600 28684 10606
rect 28632 10542 28684 10548
rect 28080 10532 28132 10538
rect 28080 10474 28132 10480
rect 28448 10532 28500 10538
rect 28448 10474 28500 10480
rect 28000 10118 28120 10146
rect 28460 10130 28488 10474
rect 27896 10056 27948 10062
rect 27896 9998 27948 10004
rect 27988 10056 28040 10062
rect 27988 9998 28040 10004
rect 27068 7948 27120 7954
rect 27068 7890 27120 7896
rect 27436 7948 27488 7954
rect 27632 7942 27844 7970
rect 27436 7890 27488 7896
rect 27816 7342 27844 7942
rect 27804 7336 27856 7342
rect 27804 7278 27856 7284
rect 27620 6792 27672 6798
rect 27620 6734 27672 6740
rect 27528 6656 27580 6662
rect 27528 6598 27580 6604
rect 27540 6458 27568 6598
rect 27528 6452 27580 6458
rect 27528 6394 27580 6400
rect 26424 6316 26476 6322
rect 26424 6258 26476 6264
rect 26976 6316 27028 6322
rect 26976 6258 27028 6264
rect 26332 5772 26384 5778
rect 26332 5714 26384 5720
rect 26436 5370 26464 6258
rect 26884 6248 26936 6254
rect 26884 6190 26936 6196
rect 26896 5846 26924 6190
rect 26884 5840 26936 5846
rect 26884 5782 26936 5788
rect 27632 5778 27660 6734
rect 27908 6322 27936 9998
rect 28000 8974 28028 9998
rect 28092 9994 28120 10118
rect 28448 10124 28500 10130
rect 28448 10066 28500 10072
rect 28080 9988 28132 9994
rect 28080 9930 28132 9936
rect 28644 9926 28672 10542
rect 28172 9920 28224 9926
rect 28172 9862 28224 9868
rect 28632 9920 28684 9926
rect 28632 9862 28684 9868
rect 27988 8968 28040 8974
rect 27988 8910 28040 8916
rect 28000 8498 28028 8910
rect 27988 8492 28040 8498
rect 27988 8434 28040 8440
rect 28184 7818 28212 9862
rect 28264 9444 28316 9450
rect 28264 9386 28316 9392
rect 28276 9024 28304 9386
rect 28356 9036 28408 9042
rect 28276 8996 28356 9024
rect 28356 8978 28408 8984
rect 28356 8492 28408 8498
rect 28356 8434 28408 8440
rect 28368 7954 28396 8434
rect 28356 7948 28408 7954
rect 28356 7890 28408 7896
rect 28172 7812 28224 7818
rect 28224 7772 28304 7800
rect 28172 7754 28224 7760
rect 28172 7472 28224 7478
rect 28172 7414 28224 7420
rect 27988 7200 28040 7206
rect 27988 7142 28040 7148
rect 27896 6316 27948 6322
rect 27896 6258 27948 6264
rect 27620 5772 27672 5778
rect 27620 5714 27672 5720
rect 27896 5772 27948 5778
rect 27896 5714 27948 5720
rect 26424 5364 26476 5370
rect 26424 5306 26476 5312
rect 27528 5160 27580 5166
rect 27528 5102 27580 5108
rect 24860 4684 24912 4690
rect 24860 4626 24912 4632
rect 26148 4684 26200 4690
rect 26148 4626 26200 4632
rect 26884 4548 26936 4554
rect 26884 4490 26936 4496
rect 26424 4140 26476 4146
rect 26700 4140 26752 4146
rect 26476 4100 26700 4128
rect 26424 4082 26476 4088
rect 26700 4082 26752 4088
rect 25872 4072 25924 4078
rect 25872 4014 25924 4020
rect 26056 4072 26108 4078
rect 26056 4014 26108 4020
rect 26332 4072 26384 4078
rect 26332 4014 26384 4020
rect 24492 4004 24544 4010
rect 24492 3946 24544 3952
rect 23756 3936 23808 3942
rect 23756 3878 23808 3884
rect 22652 3596 22704 3602
rect 22652 3538 22704 3544
rect 22836 3596 22888 3602
rect 22836 3538 22888 3544
rect 22284 3460 22336 3466
rect 22284 3402 22336 3408
rect 22100 2508 22152 2514
rect 22100 2450 22152 2456
rect 22560 2440 22612 2446
rect 22664 2428 22692 3538
rect 22612 2400 22692 2428
rect 22560 2382 22612 2388
rect 23388 2304 23440 2310
rect 23388 2246 23440 2252
rect 23400 2106 23428 2246
rect 23388 2100 23440 2106
rect 23388 2042 23440 2048
rect 23768 800 23796 3878
rect 25884 3602 25912 4014
rect 25872 3596 25924 3602
rect 25872 3538 25924 3544
rect 23848 3460 23900 3466
rect 23848 3402 23900 3408
rect 23860 3194 23888 3402
rect 24124 3392 24176 3398
rect 24124 3334 24176 3340
rect 24768 3392 24820 3398
rect 24768 3334 24820 3340
rect 23848 3188 23900 3194
rect 23848 3130 23900 3136
rect 24136 3058 24164 3334
rect 24124 3052 24176 3058
rect 24124 2994 24176 3000
rect 24780 2990 24808 3334
rect 26068 3194 26096 4014
rect 26056 3188 26108 3194
rect 26056 3130 26108 3136
rect 26344 2990 26372 4014
rect 26424 3936 26476 3942
rect 26424 3878 26476 3884
rect 26516 3936 26568 3942
rect 26516 3878 26568 3884
rect 24032 2984 24084 2990
rect 24032 2926 24084 2932
rect 24768 2984 24820 2990
rect 24768 2926 24820 2932
rect 26332 2984 26384 2990
rect 26332 2926 26384 2932
rect 24044 2650 24072 2926
rect 26436 2922 26464 3878
rect 26528 3210 26556 3878
rect 26700 3460 26752 3466
rect 26700 3402 26752 3408
rect 26528 3182 26648 3210
rect 24308 2916 24360 2922
rect 24308 2858 24360 2864
rect 26424 2916 26476 2922
rect 26424 2858 26476 2864
rect 24032 2644 24084 2650
rect 24032 2586 24084 2592
rect 24320 2514 24348 2858
rect 26620 2582 26648 3182
rect 26608 2576 26660 2582
rect 26608 2518 26660 2524
rect 24308 2508 24360 2514
rect 24308 2450 24360 2456
rect 26712 2446 26740 3402
rect 26896 3398 26924 4490
rect 27068 4072 27120 4078
rect 27068 4014 27120 4020
rect 27080 3738 27108 4014
rect 27540 4010 27568 5102
rect 27620 5092 27672 5098
rect 27620 5034 27672 5040
rect 27632 4690 27660 5034
rect 27620 4684 27672 4690
rect 27620 4626 27672 4632
rect 27804 4684 27856 4690
rect 27804 4626 27856 4632
rect 27528 4004 27580 4010
rect 27528 3946 27580 3952
rect 27068 3732 27120 3738
rect 27068 3674 27120 3680
rect 27816 3534 27844 4626
rect 27908 3942 27936 5714
rect 27896 3936 27948 3942
rect 27896 3878 27948 3884
rect 27908 3670 27936 3878
rect 27896 3664 27948 3670
rect 27896 3606 27948 3612
rect 28000 3602 28028 7142
rect 28184 6866 28212 7414
rect 28172 6860 28224 6866
rect 28172 6802 28224 6808
rect 28184 6458 28212 6802
rect 28172 6452 28224 6458
rect 28172 6394 28224 6400
rect 28172 5908 28224 5914
rect 28172 5850 28224 5856
rect 28184 5234 28212 5850
rect 28172 5228 28224 5234
rect 28172 5170 28224 5176
rect 28276 5166 28304 7772
rect 28632 6792 28684 6798
rect 28632 6734 28684 6740
rect 28644 5846 28672 6734
rect 28632 5840 28684 5846
rect 28632 5782 28684 5788
rect 28644 5234 28672 5782
rect 28920 5574 28948 11698
rect 29000 9648 29052 9654
rect 29000 9590 29052 9596
rect 29012 8906 29040 9590
rect 29104 9518 29132 12038
rect 29932 11558 29960 12718
rect 30104 12368 30156 12374
rect 30104 12310 30156 12316
rect 29920 11552 29972 11558
rect 29920 11494 29972 11500
rect 29932 11218 29960 11494
rect 29920 11212 29972 11218
rect 29920 11154 29972 11160
rect 30116 11121 30144 12310
rect 30196 12096 30248 12102
rect 30196 12038 30248 12044
rect 30208 11694 30236 12038
rect 30392 11880 30420 14010
rect 30484 13190 30512 15966
rect 30576 15366 30604 21422
rect 30656 19712 30708 19718
rect 30656 19654 30708 19660
rect 30668 18834 30696 19654
rect 30656 18828 30708 18834
rect 30656 18770 30708 18776
rect 30564 15360 30616 15366
rect 30564 15302 30616 15308
rect 30564 14884 30616 14890
rect 30564 14826 30616 14832
rect 30576 14618 30604 14826
rect 30564 14612 30616 14618
rect 30564 14554 30616 14560
rect 30576 13870 30604 14554
rect 30760 14550 30788 27474
rect 31036 27146 31064 37674
rect 31496 36854 31524 37742
rect 33612 37262 33640 37742
rect 33968 37324 34020 37330
rect 33968 37266 34020 37272
rect 33600 37256 33652 37262
rect 33600 37198 33652 37204
rect 31484 36848 31536 36854
rect 31484 36790 31536 36796
rect 31392 36712 31444 36718
rect 31392 36654 31444 36660
rect 31116 36032 31168 36038
rect 31116 35974 31168 35980
rect 31128 35698 31156 35974
rect 31116 35692 31168 35698
rect 31116 35634 31168 35640
rect 31300 35080 31352 35086
rect 31300 35022 31352 35028
rect 31312 34610 31340 35022
rect 31300 34604 31352 34610
rect 31300 34546 31352 34552
rect 31300 34468 31352 34474
rect 31300 34410 31352 34416
rect 31312 33114 31340 34410
rect 31404 34202 31432 36654
rect 33612 36242 33640 37198
rect 33692 36848 33744 36854
rect 33692 36790 33744 36796
rect 32128 36236 32180 36242
rect 32128 36178 32180 36184
rect 33600 36236 33652 36242
rect 33600 36178 33652 36184
rect 32140 35630 32168 36178
rect 32404 36168 32456 36174
rect 32404 36110 32456 36116
rect 32416 35834 32444 36110
rect 33508 36032 33560 36038
rect 33508 35974 33560 35980
rect 32404 35828 32456 35834
rect 32404 35770 32456 35776
rect 33232 35828 33284 35834
rect 33232 35770 33284 35776
rect 32128 35624 32180 35630
rect 32128 35566 32180 35572
rect 33048 35624 33100 35630
rect 33048 35566 33100 35572
rect 31576 35488 31628 35494
rect 31576 35430 31628 35436
rect 31392 34196 31444 34202
rect 31392 34138 31444 34144
rect 31588 33998 31616 35430
rect 32140 35154 32168 35566
rect 32036 35148 32088 35154
rect 32036 35090 32088 35096
rect 32128 35148 32180 35154
rect 32128 35090 32180 35096
rect 32048 34746 32076 35090
rect 33060 34746 33088 35566
rect 32036 34740 32088 34746
rect 32036 34682 32088 34688
rect 33048 34740 33100 34746
rect 33048 34682 33100 34688
rect 32496 34400 32548 34406
rect 32496 34342 32548 34348
rect 32508 34066 32536 34342
rect 32312 34060 32364 34066
rect 32312 34002 32364 34008
rect 32496 34060 32548 34066
rect 32496 34002 32548 34008
rect 31576 33992 31628 33998
rect 31576 33934 31628 33940
rect 31588 33658 31616 33934
rect 31576 33652 31628 33658
rect 31576 33594 31628 33600
rect 31484 33312 31536 33318
rect 31484 33254 31536 33260
rect 31300 33108 31352 33114
rect 31300 33050 31352 33056
rect 31116 30660 31168 30666
rect 31116 30602 31168 30608
rect 31128 30258 31156 30602
rect 31116 30252 31168 30258
rect 31116 30194 31168 30200
rect 31300 29096 31352 29102
rect 31300 29038 31352 29044
rect 31312 27878 31340 29038
rect 31300 27872 31352 27878
rect 31300 27814 31352 27820
rect 31392 27532 31444 27538
rect 31392 27474 31444 27480
rect 30944 27118 31064 27146
rect 30840 26920 30892 26926
rect 30840 26862 30892 26868
rect 30852 26518 30880 26862
rect 30840 26512 30892 26518
rect 30840 26454 30892 26460
rect 30840 24404 30892 24410
rect 30840 24346 30892 24352
rect 30852 24070 30880 24346
rect 30840 24064 30892 24070
rect 30840 24006 30892 24012
rect 30840 23180 30892 23186
rect 30840 23122 30892 23128
rect 30852 22001 30880 23122
rect 30944 22438 30972 27118
rect 31024 25356 31076 25362
rect 31024 25298 31076 25304
rect 31036 24750 31064 25298
rect 31116 25220 31168 25226
rect 31116 25162 31168 25168
rect 31024 24744 31076 24750
rect 31024 24686 31076 24692
rect 31024 24064 31076 24070
rect 31024 24006 31076 24012
rect 31036 23526 31064 24006
rect 31024 23520 31076 23526
rect 31024 23462 31076 23468
rect 31024 23044 31076 23050
rect 31024 22986 31076 22992
rect 31036 22710 31064 22986
rect 31024 22704 31076 22710
rect 31024 22646 31076 22652
rect 30932 22432 30984 22438
rect 30932 22374 30984 22380
rect 31128 22137 31156 25162
rect 31404 23526 31432 27474
rect 31392 23520 31444 23526
rect 31392 23462 31444 23468
rect 31208 23044 31260 23050
rect 31208 22986 31260 22992
rect 31220 22574 31248 22986
rect 31496 22982 31524 33254
rect 32220 32292 32272 32298
rect 32220 32234 32272 32240
rect 32128 32224 32180 32230
rect 32128 32166 32180 32172
rect 32140 31890 32168 32166
rect 32128 31884 32180 31890
rect 32048 31844 32128 31872
rect 31576 31272 31628 31278
rect 31576 31214 31628 31220
rect 31588 30598 31616 31214
rect 31576 30592 31628 30598
rect 31576 30534 31628 30540
rect 31588 29578 31616 30534
rect 32048 30394 32076 31844
rect 32128 31826 32180 31832
rect 32232 31278 32260 32234
rect 32220 31272 32272 31278
rect 32220 31214 32272 31220
rect 32220 30728 32272 30734
rect 32220 30670 32272 30676
rect 32232 30394 32260 30670
rect 32036 30388 32088 30394
rect 32036 30330 32088 30336
rect 32220 30388 32272 30394
rect 32220 30330 32272 30336
rect 32232 29782 32260 30330
rect 32220 29776 32272 29782
rect 32220 29718 32272 29724
rect 31576 29572 31628 29578
rect 31576 29514 31628 29520
rect 31576 29164 31628 29170
rect 31576 29106 31628 29112
rect 31588 28200 31616 29106
rect 32324 29102 32352 34002
rect 32508 33522 32536 34002
rect 33244 33522 33272 35770
rect 33520 35154 33548 35974
rect 33508 35148 33560 35154
rect 33508 35090 33560 35096
rect 32496 33516 32548 33522
rect 32496 33458 32548 33464
rect 33232 33516 33284 33522
rect 33232 33458 33284 33464
rect 32864 32972 32916 32978
rect 32864 32914 32916 32920
rect 32772 32904 32824 32910
rect 32772 32846 32824 32852
rect 32404 32836 32456 32842
rect 32404 32778 32456 32784
rect 32416 31890 32444 32778
rect 32404 31884 32456 31890
rect 32404 31826 32456 31832
rect 32784 30598 32812 32846
rect 32876 32502 32904 32914
rect 33232 32768 33284 32774
rect 33232 32710 33284 32716
rect 32864 32496 32916 32502
rect 32864 32438 32916 32444
rect 32956 32360 33008 32366
rect 32956 32302 33008 32308
rect 32772 30592 32824 30598
rect 32772 30534 32824 30540
rect 32496 30116 32548 30122
rect 32496 30058 32548 30064
rect 32312 29096 32364 29102
rect 32312 29038 32364 29044
rect 32508 28694 32536 30058
rect 32968 29850 32996 32302
rect 33244 31278 33272 32710
rect 33324 32292 33376 32298
rect 33324 32234 33376 32240
rect 33336 31346 33364 32234
rect 33704 32026 33732 36790
rect 33784 34536 33836 34542
rect 33784 34478 33836 34484
rect 33796 33658 33824 34478
rect 33784 33652 33836 33658
rect 33784 33594 33836 33600
rect 33784 32972 33836 32978
rect 33784 32914 33836 32920
rect 33876 32972 33928 32978
rect 33876 32914 33928 32920
rect 33692 32020 33744 32026
rect 33692 31962 33744 31968
rect 33324 31340 33376 31346
rect 33324 31282 33376 31288
rect 33232 31272 33284 31278
rect 33232 31214 33284 31220
rect 33048 31136 33100 31142
rect 33048 31078 33100 31084
rect 33060 30802 33088 31078
rect 33336 30870 33364 31282
rect 33600 31204 33652 31210
rect 33600 31146 33652 31152
rect 33324 30864 33376 30870
rect 33324 30806 33376 30812
rect 33048 30796 33100 30802
rect 33048 30738 33100 30744
rect 33140 30796 33192 30802
rect 33140 30738 33192 30744
rect 33152 30190 33180 30738
rect 33140 30184 33192 30190
rect 33140 30126 33192 30132
rect 32956 29844 33008 29850
rect 32956 29786 33008 29792
rect 32588 29708 32640 29714
rect 32588 29650 32640 29656
rect 32600 29170 32628 29650
rect 32588 29164 32640 29170
rect 32588 29106 32640 29112
rect 32496 28688 32548 28694
rect 32496 28630 32548 28636
rect 32772 28552 32824 28558
rect 32772 28494 32824 28500
rect 32784 28218 32812 28494
rect 31760 28212 31812 28218
rect 31588 28172 31760 28200
rect 31588 26926 31616 28172
rect 31760 28154 31812 28160
rect 32772 28212 32824 28218
rect 32772 28154 32824 28160
rect 32968 28014 32996 29786
rect 33232 29640 33284 29646
rect 33232 29582 33284 29588
rect 33140 29232 33192 29238
rect 33140 29174 33192 29180
rect 33048 28144 33100 28150
rect 33048 28086 33100 28092
rect 32956 28008 33008 28014
rect 32956 27950 33008 27956
rect 33060 27538 33088 28086
rect 33152 28082 33180 29174
rect 33244 29102 33272 29582
rect 33232 29096 33284 29102
rect 33232 29038 33284 29044
rect 33612 28966 33640 31146
rect 33600 28960 33652 28966
rect 33600 28902 33652 28908
rect 33508 28484 33560 28490
rect 33508 28426 33560 28432
rect 33140 28076 33192 28082
rect 33140 28018 33192 28024
rect 33232 28008 33284 28014
rect 33232 27950 33284 27956
rect 33244 27606 33272 27950
rect 33232 27600 33284 27606
rect 33232 27542 33284 27548
rect 32496 27532 32548 27538
rect 32496 27474 32548 27480
rect 33048 27532 33100 27538
rect 33048 27474 33100 27480
rect 31668 27464 31720 27470
rect 31668 27406 31720 27412
rect 31576 26920 31628 26926
rect 31576 26862 31628 26868
rect 31588 26382 31616 26862
rect 31576 26376 31628 26382
rect 31576 26318 31628 26324
rect 31680 26314 31708 27406
rect 32220 27328 32272 27334
rect 32220 27270 32272 27276
rect 31852 26920 31904 26926
rect 31852 26862 31904 26868
rect 31668 26308 31720 26314
rect 31668 26250 31720 26256
rect 31680 24750 31708 26250
rect 31864 25974 31892 26862
rect 32128 26444 32180 26450
rect 32128 26386 32180 26392
rect 32140 26042 32168 26386
rect 32128 26036 32180 26042
rect 32128 25978 32180 25984
rect 31852 25968 31904 25974
rect 31852 25910 31904 25916
rect 32232 25838 32260 27270
rect 32508 27130 32536 27474
rect 33244 27130 33272 27542
rect 33520 27402 33548 28426
rect 33612 28014 33640 28902
rect 33600 28008 33652 28014
rect 33600 27950 33652 27956
rect 33612 27470 33640 27950
rect 33600 27464 33652 27470
rect 33600 27406 33652 27412
rect 33508 27396 33560 27402
rect 33508 27338 33560 27344
rect 32496 27124 32548 27130
rect 32496 27066 32548 27072
rect 33232 27124 33284 27130
rect 33232 27066 33284 27072
rect 32312 26988 32364 26994
rect 32312 26930 32364 26936
rect 32324 25906 32352 26930
rect 33704 26926 33732 31962
rect 33796 31210 33824 32914
rect 33888 32434 33916 32914
rect 33876 32428 33928 32434
rect 33876 32370 33928 32376
rect 33888 31958 33916 32370
rect 33876 31952 33928 31958
rect 33876 31894 33928 31900
rect 33784 31204 33836 31210
rect 33784 31146 33836 31152
rect 33876 30048 33928 30054
rect 33876 29990 33928 29996
rect 33888 29714 33916 29990
rect 33876 29708 33928 29714
rect 33876 29650 33928 29656
rect 33876 28552 33928 28558
rect 33876 28494 33928 28500
rect 33888 27674 33916 28494
rect 33876 27668 33928 27674
rect 33876 27610 33928 27616
rect 33692 26920 33744 26926
rect 33692 26862 33744 26868
rect 33508 26784 33560 26790
rect 33508 26726 33560 26732
rect 33520 26450 33548 26726
rect 33324 26444 33376 26450
rect 33324 26386 33376 26392
rect 33508 26444 33560 26450
rect 33508 26386 33560 26392
rect 32312 25900 32364 25906
rect 32312 25842 32364 25848
rect 32220 25832 32272 25838
rect 32220 25774 32272 25780
rect 31668 24744 31720 24750
rect 31668 24686 31720 24692
rect 32220 24744 32272 24750
rect 32220 24686 32272 24692
rect 32232 24070 32260 24686
rect 32220 24064 32272 24070
rect 32220 24006 32272 24012
rect 31484 22976 31536 22982
rect 31484 22918 31536 22924
rect 31208 22568 31260 22574
rect 31208 22510 31260 22516
rect 31576 22568 31628 22574
rect 31576 22510 31628 22516
rect 31114 22128 31170 22137
rect 31114 22063 31170 22072
rect 30838 21992 30894 22001
rect 30838 21927 30894 21936
rect 31128 21486 31156 22063
rect 31116 21480 31168 21486
rect 31116 21422 31168 21428
rect 31300 21344 31352 21350
rect 31300 21286 31352 21292
rect 31116 20596 31168 20602
rect 31116 20538 31168 20544
rect 30840 18216 30892 18222
rect 30840 18158 30892 18164
rect 30852 16522 30880 18158
rect 31128 17746 31156 20538
rect 31312 20466 31340 21286
rect 31588 20874 31616 22510
rect 32128 22024 32180 22030
rect 32128 21966 32180 21972
rect 31852 21480 31904 21486
rect 31852 21422 31904 21428
rect 32036 21480 32088 21486
rect 32036 21422 32088 21428
rect 31576 20868 31628 20874
rect 31576 20810 31628 20816
rect 31300 20460 31352 20466
rect 31300 20402 31352 20408
rect 31116 17740 31168 17746
rect 31116 17682 31168 17688
rect 31128 16658 31156 17682
rect 31116 16652 31168 16658
rect 31116 16594 31168 16600
rect 30840 16516 30892 16522
rect 30840 16458 30892 16464
rect 31128 16114 31156 16594
rect 31116 16108 31168 16114
rect 31116 16050 31168 16056
rect 31024 16040 31076 16046
rect 31024 15982 31076 15988
rect 30932 15428 30984 15434
rect 30932 15370 30984 15376
rect 30748 14544 30800 14550
rect 30748 14486 30800 14492
rect 30564 13864 30616 13870
rect 30564 13806 30616 13812
rect 30840 13456 30892 13462
rect 30840 13398 30892 13404
rect 30472 13184 30524 13190
rect 30472 13126 30524 13132
rect 30484 12220 30512 13126
rect 30748 12912 30800 12918
rect 30748 12854 30800 12860
rect 30564 12640 30616 12646
rect 30564 12582 30616 12588
rect 30576 12374 30604 12582
rect 30564 12368 30616 12374
rect 30564 12310 30616 12316
rect 30654 12336 30710 12345
rect 30760 12306 30788 12854
rect 30852 12850 30880 13398
rect 30840 12844 30892 12850
rect 30840 12786 30892 12792
rect 30944 12594 30972 15370
rect 30852 12566 30972 12594
rect 30654 12271 30656 12280
rect 30708 12271 30710 12280
rect 30748 12300 30800 12306
rect 30656 12242 30708 12248
rect 30748 12242 30800 12248
rect 30484 12192 30604 12220
rect 30472 11892 30524 11898
rect 30392 11852 30472 11880
rect 30472 11834 30524 11840
rect 30576 11694 30604 12192
rect 30748 12164 30800 12170
rect 30748 12106 30800 12112
rect 30760 11830 30788 12106
rect 30748 11824 30800 11830
rect 30748 11766 30800 11772
rect 30196 11688 30248 11694
rect 30196 11630 30248 11636
rect 30564 11688 30616 11694
rect 30564 11630 30616 11636
rect 30746 11656 30802 11665
rect 30746 11591 30748 11600
rect 30800 11591 30802 11600
rect 30748 11562 30800 11568
rect 30196 11348 30248 11354
rect 30196 11290 30248 11296
rect 30102 11112 30158 11121
rect 30102 11047 30158 11056
rect 29460 10736 29512 10742
rect 29460 10678 29512 10684
rect 29472 10606 29500 10678
rect 29460 10600 29512 10606
rect 29460 10542 29512 10548
rect 29368 9988 29420 9994
rect 29368 9930 29420 9936
rect 29380 9518 29408 9930
rect 30104 9920 30156 9926
rect 30104 9862 30156 9868
rect 29092 9512 29144 9518
rect 29092 9454 29144 9460
rect 29184 9512 29236 9518
rect 29184 9454 29236 9460
rect 29368 9512 29420 9518
rect 29368 9454 29420 9460
rect 29196 9382 29224 9454
rect 29184 9376 29236 9382
rect 29184 9318 29236 9324
rect 29000 8900 29052 8906
rect 29000 8842 29052 8848
rect 29092 8424 29144 8430
rect 29196 8412 29224 9318
rect 29276 8832 29328 8838
rect 29276 8774 29328 8780
rect 29144 8384 29224 8412
rect 29092 8366 29144 8372
rect 29104 7886 29132 8366
rect 29288 7954 29316 8774
rect 29380 8090 29408 9454
rect 30116 9042 30144 9862
rect 30208 9722 30236 11290
rect 30852 11218 30880 12566
rect 30932 12368 30984 12374
rect 30932 12310 30984 12316
rect 30840 11212 30892 11218
rect 30840 11154 30892 11160
rect 30472 10464 30524 10470
rect 30472 10406 30524 10412
rect 30380 10260 30432 10266
rect 30380 10202 30432 10208
rect 30392 9722 30420 10202
rect 30196 9716 30248 9722
rect 30196 9658 30248 9664
rect 30380 9716 30432 9722
rect 30380 9658 30432 9664
rect 30208 9178 30236 9658
rect 30484 9586 30512 10406
rect 30564 10124 30616 10130
rect 30564 10066 30616 10072
rect 30840 10124 30892 10130
rect 30840 10066 30892 10072
rect 30576 9994 30604 10066
rect 30656 10056 30708 10062
rect 30656 9998 30708 10004
rect 30564 9988 30616 9994
rect 30564 9930 30616 9936
rect 30668 9654 30696 9998
rect 30656 9648 30708 9654
rect 30656 9590 30708 9596
rect 30472 9580 30524 9586
rect 30472 9522 30524 9528
rect 30852 9382 30880 10066
rect 30840 9376 30892 9382
rect 30840 9318 30892 9324
rect 30196 9172 30248 9178
rect 30196 9114 30248 9120
rect 30104 9036 30156 9042
rect 30104 8978 30156 8984
rect 29828 8900 29880 8906
rect 29828 8842 29880 8848
rect 29552 8424 29604 8430
rect 29552 8366 29604 8372
rect 29368 8084 29420 8090
rect 29368 8026 29420 8032
rect 29276 7948 29328 7954
rect 29276 7890 29328 7896
rect 29092 7880 29144 7886
rect 29092 7822 29144 7828
rect 29000 7336 29052 7342
rect 29000 7278 29052 7284
rect 29012 6934 29040 7278
rect 29000 6928 29052 6934
rect 29000 6870 29052 6876
rect 29104 6118 29132 7822
rect 29460 7744 29512 7750
rect 29460 7686 29512 7692
rect 29472 7002 29500 7686
rect 29564 7410 29592 8366
rect 29552 7404 29604 7410
rect 29552 7346 29604 7352
rect 29552 7268 29604 7274
rect 29552 7210 29604 7216
rect 29564 7002 29592 7210
rect 29460 6996 29512 7002
rect 29460 6938 29512 6944
rect 29552 6996 29604 7002
rect 29552 6938 29604 6944
rect 29472 6458 29500 6938
rect 29840 6866 29868 8842
rect 30564 7880 30616 7886
rect 30564 7822 30616 7828
rect 30288 7268 30340 7274
rect 30288 7210 30340 7216
rect 29828 6860 29880 6866
rect 29828 6802 29880 6808
rect 29920 6792 29972 6798
rect 29920 6734 29972 6740
rect 29932 6458 29960 6734
rect 29460 6452 29512 6458
rect 29460 6394 29512 6400
rect 29920 6452 29972 6458
rect 29920 6394 29972 6400
rect 29276 6248 29328 6254
rect 29276 6190 29328 6196
rect 29092 6112 29144 6118
rect 29092 6054 29144 6060
rect 29000 5636 29052 5642
rect 29000 5578 29052 5584
rect 28908 5568 28960 5574
rect 28908 5510 28960 5516
rect 28632 5228 28684 5234
rect 28632 5170 28684 5176
rect 28264 5160 28316 5166
rect 28264 5102 28316 5108
rect 29012 4622 29040 5578
rect 29104 5166 29132 6054
rect 29288 5778 29316 6190
rect 29932 5914 29960 6394
rect 30104 6316 30156 6322
rect 30104 6258 30156 6264
rect 29920 5908 29972 5914
rect 29920 5850 29972 5856
rect 29932 5778 29960 5850
rect 30116 5778 30144 6258
rect 29276 5772 29328 5778
rect 29276 5714 29328 5720
rect 29920 5772 29972 5778
rect 29920 5714 29972 5720
rect 30104 5772 30156 5778
rect 30104 5714 30156 5720
rect 29092 5160 29144 5166
rect 29092 5102 29144 5108
rect 29000 4616 29052 4622
rect 29000 4558 29052 4564
rect 27988 3596 28040 3602
rect 27988 3538 28040 3544
rect 28264 3596 28316 3602
rect 28264 3538 28316 3544
rect 27804 3528 27856 3534
rect 27804 3470 27856 3476
rect 27068 3460 27120 3466
rect 27068 3402 27120 3408
rect 26884 3392 26936 3398
rect 26884 3334 26936 3340
rect 26896 2514 26924 3334
rect 27080 2990 27108 3402
rect 27816 3194 27844 3470
rect 28276 3398 28304 3538
rect 29104 3534 29132 5102
rect 29288 4078 29316 5714
rect 29368 5704 29420 5710
rect 29368 5646 29420 5652
rect 29380 4690 29408 5646
rect 29552 5160 29604 5166
rect 30116 5114 30144 5714
rect 29552 5102 29604 5108
rect 29564 4758 29592 5102
rect 30024 5086 30144 5114
rect 30024 5030 30052 5086
rect 30012 5024 30064 5030
rect 30012 4966 30064 4972
rect 29552 4752 29604 4758
rect 29552 4694 29604 4700
rect 29368 4684 29420 4690
rect 29368 4626 29420 4632
rect 29460 4208 29512 4214
rect 29460 4150 29512 4156
rect 29276 4072 29328 4078
rect 29276 4014 29328 4020
rect 29092 3528 29144 3534
rect 29092 3470 29144 3476
rect 29472 3516 29500 4150
rect 30300 3738 30328 7210
rect 30576 6866 30604 7822
rect 30852 7478 30880 9318
rect 30944 7868 30972 12310
rect 31036 9042 31064 15982
rect 31484 14952 31536 14958
rect 31484 14894 31536 14900
rect 31116 14884 31168 14890
rect 31116 14826 31168 14832
rect 31392 14884 31444 14890
rect 31392 14826 31444 14832
rect 31128 14006 31156 14826
rect 31116 14000 31168 14006
rect 31116 13942 31168 13948
rect 31128 13394 31156 13942
rect 31404 13870 31432 14826
rect 31496 14074 31524 14894
rect 31484 14068 31536 14074
rect 31484 14010 31536 14016
rect 31392 13864 31444 13870
rect 31392 13806 31444 13812
rect 31116 13388 31168 13394
rect 31116 13330 31168 13336
rect 31392 12980 31444 12986
rect 31392 12922 31444 12928
rect 31404 12782 31432 12922
rect 31116 12776 31168 12782
rect 31114 12744 31116 12753
rect 31392 12776 31444 12782
rect 31168 12744 31170 12753
rect 31392 12718 31444 12724
rect 31114 12679 31170 12688
rect 31392 12436 31444 12442
rect 31392 12378 31444 12384
rect 31404 12322 31432 12378
rect 31220 12294 31432 12322
rect 31220 11354 31248 12294
rect 31392 12232 31444 12238
rect 31312 12192 31392 12220
rect 31208 11348 31260 11354
rect 31208 11290 31260 11296
rect 31116 11212 31168 11218
rect 31116 11154 31168 11160
rect 31128 10130 31156 11154
rect 31208 10804 31260 10810
rect 31208 10746 31260 10752
rect 31116 10124 31168 10130
rect 31116 10066 31168 10072
rect 31220 9110 31248 10746
rect 31312 10266 31340 12192
rect 31392 12174 31444 12180
rect 31484 11688 31536 11694
rect 31404 11648 31484 11676
rect 31404 11286 31432 11648
rect 31484 11630 31536 11636
rect 31588 11354 31616 20810
rect 31864 19310 31892 21422
rect 32048 21078 32076 21422
rect 32036 21072 32088 21078
rect 32036 21014 32088 21020
rect 32036 19916 32088 19922
rect 32036 19858 32088 19864
rect 32048 19718 32076 19858
rect 32036 19712 32088 19718
rect 32036 19654 32088 19660
rect 32048 19310 32076 19654
rect 31852 19304 31904 19310
rect 31852 19246 31904 19252
rect 32036 19304 32088 19310
rect 32036 19246 32088 19252
rect 31864 18834 31892 19246
rect 32048 18834 32076 19246
rect 31852 18828 31904 18834
rect 31852 18770 31904 18776
rect 32036 18828 32088 18834
rect 32036 18770 32088 18776
rect 31944 18624 31996 18630
rect 31944 18566 31996 18572
rect 31956 17134 31984 18566
rect 32140 17134 32168 21966
rect 32324 21486 32352 25842
rect 32496 25832 32548 25838
rect 32496 25774 32548 25780
rect 32508 25362 32536 25774
rect 33336 25362 33364 26386
rect 33600 25492 33652 25498
rect 33600 25434 33652 25440
rect 32496 25356 32548 25362
rect 32496 25298 32548 25304
rect 33324 25356 33376 25362
rect 33324 25298 33376 25304
rect 33416 25288 33468 25294
rect 33416 25230 33468 25236
rect 32588 24744 32640 24750
rect 32588 24686 32640 24692
rect 32404 24676 32456 24682
rect 32404 24618 32456 24624
rect 32416 24562 32444 24618
rect 32416 24534 32536 24562
rect 32508 24274 32536 24534
rect 32496 24268 32548 24274
rect 32496 24210 32548 24216
rect 32508 23186 32536 24210
rect 32600 24206 32628 24686
rect 33324 24676 33376 24682
rect 33324 24618 33376 24624
rect 33336 24274 33364 24618
rect 33324 24268 33376 24274
rect 33324 24210 33376 24216
rect 32588 24200 32640 24206
rect 32588 24142 32640 24148
rect 33336 23662 33364 24210
rect 32956 23656 33008 23662
rect 32956 23598 33008 23604
rect 33324 23656 33376 23662
rect 33324 23598 33376 23604
rect 32496 23180 32548 23186
rect 32496 23122 32548 23128
rect 32968 23118 32996 23598
rect 33428 23526 33456 25230
rect 33612 24274 33640 25434
rect 33600 24268 33652 24274
rect 33520 24228 33600 24256
rect 33324 23520 33376 23526
rect 33324 23462 33376 23468
rect 33416 23520 33468 23526
rect 33416 23462 33468 23468
rect 33336 23225 33364 23462
rect 33322 23216 33378 23225
rect 33048 23180 33100 23186
rect 33322 23151 33378 23160
rect 33048 23122 33100 23128
rect 32956 23112 33008 23118
rect 32956 23054 33008 23060
rect 32404 22024 32456 22030
rect 32404 21966 32456 21972
rect 32312 21480 32364 21486
rect 32312 21422 32364 21428
rect 32324 17746 32352 21422
rect 32416 21350 32444 21966
rect 32404 21344 32456 21350
rect 32404 21286 32456 21292
rect 32680 21004 32732 21010
rect 32680 20946 32732 20952
rect 32864 21004 32916 21010
rect 32864 20946 32916 20952
rect 32692 20262 32720 20946
rect 32496 20256 32548 20262
rect 32496 20198 32548 20204
rect 32680 20256 32732 20262
rect 32680 20198 32732 20204
rect 32508 19378 32536 20198
rect 32496 19372 32548 19378
rect 32496 19314 32548 19320
rect 32508 18834 32536 19314
rect 32496 18828 32548 18834
rect 32496 18770 32548 18776
rect 32876 18086 32904 20946
rect 33060 20942 33088 23122
rect 33336 22574 33364 23151
rect 33324 22568 33376 22574
rect 33324 22510 33376 22516
rect 33428 22386 33456 23462
rect 33520 22506 33548 24228
rect 33600 24210 33652 24216
rect 33600 24132 33652 24138
rect 33600 24074 33652 24080
rect 33508 22500 33560 22506
rect 33508 22442 33560 22448
rect 33428 22358 33548 22386
rect 33232 22160 33284 22166
rect 33232 22102 33284 22108
rect 33244 21486 33272 22102
rect 33520 21962 33548 22358
rect 33508 21956 33560 21962
rect 33508 21898 33560 21904
rect 33232 21480 33284 21486
rect 33232 21422 33284 21428
rect 33520 21078 33548 21898
rect 33508 21072 33560 21078
rect 33508 21014 33560 21020
rect 33416 21004 33468 21010
rect 33416 20946 33468 20952
rect 33048 20936 33100 20942
rect 33048 20878 33100 20884
rect 33048 20596 33100 20602
rect 33048 20538 33100 20544
rect 33060 20262 33088 20538
rect 33048 20256 33100 20262
rect 33048 20198 33100 20204
rect 32956 19304 33008 19310
rect 32956 19246 33008 19252
rect 32968 18834 32996 19246
rect 33060 18834 33088 20198
rect 33140 19236 33192 19242
rect 33140 19178 33192 19184
rect 32956 18828 33008 18834
rect 32956 18770 33008 18776
rect 33048 18828 33100 18834
rect 33048 18770 33100 18776
rect 32968 18358 32996 18770
rect 33060 18698 33088 18770
rect 33048 18692 33100 18698
rect 33048 18634 33100 18640
rect 32956 18352 33008 18358
rect 32956 18294 33008 18300
rect 33152 18222 33180 19178
rect 33140 18216 33192 18222
rect 33140 18158 33192 18164
rect 32864 18080 32916 18086
rect 32864 18022 32916 18028
rect 32404 17876 32456 17882
rect 32404 17818 32456 17824
rect 32312 17740 32364 17746
rect 32312 17682 32364 17688
rect 31944 17128 31996 17134
rect 31944 17070 31996 17076
rect 32128 17128 32180 17134
rect 32128 17070 32180 17076
rect 31956 13870 31984 17070
rect 32036 15904 32088 15910
rect 32036 15846 32088 15852
rect 32048 15434 32076 15846
rect 32140 15502 32168 17070
rect 32220 16720 32272 16726
rect 32220 16662 32272 16668
rect 32232 16046 32260 16662
rect 32220 16040 32272 16046
rect 32220 15982 32272 15988
rect 32324 15706 32352 17682
rect 32416 17202 32444 17818
rect 32680 17740 32732 17746
rect 32680 17682 32732 17688
rect 32496 17536 32548 17542
rect 32496 17478 32548 17484
rect 32404 17196 32456 17202
rect 32404 17138 32456 17144
rect 32312 15700 32364 15706
rect 32312 15642 32364 15648
rect 32128 15496 32180 15502
rect 32128 15438 32180 15444
rect 32036 15428 32088 15434
rect 32036 15370 32088 15376
rect 32220 14884 32272 14890
rect 32220 14826 32272 14832
rect 31944 13864 31996 13870
rect 31944 13806 31996 13812
rect 32128 13456 32180 13462
rect 32128 13398 32180 13404
rect 32140 13326 32168 13398
rect 32128 13320 32180 13326
rect 32128 13262 32180 13268
rect 32128 12980 32180 12986
rect 32128 12922 32180 12928
rect 31668 12708 31720 12714
rect 31668 12650 31720 12656
rect 31680 12306 31708 12650
rect 32140 12646 32168 12922
rect 32232 12782 32260 14826
rect 32508 13870 32536 17478
rect 32588 14476 32640 14482
rect 32588 14418 32640 14424
rect 32600 14006 32628 14418
rect 32588 14000 32640 14006
rect 32588 13942 32640 13948
rect 32496 13864 32548 13870
rect 32496 13806 32548 13812
rect 32220 12776 32272 12782
rect 32220 12718 32272 12724
rect 32402 12744 32458 12753
rect 32402 12679 32458 12688
rect 32416 12646 32444 12679
rect 32128 12640 32180 12646
rect 32128 12582 32180 12588
rect 32404 12640 32456 12646
rect 32404 12582 32456 12588
rect 32692 12374 32720 17682
rect 33152 17338 33180 18158
rect 33140 17332 33192 17338
rect 33140 17274 33192 17280
rect 32772 17128 32824 17134
rect 32772 17070 32824 17076
rect 32680 12368 32732 12374
rect 32680 12310 32732 12316
rect 31668 12300 31720 12306
rect 31668 12242 31720 12248
rect 32496 12300 32548 12306
rect 32496 12242 32548 12248
rect 31668 12164 31720 12170
rect 31668 12106 31720 12112
rect 31576 11348 31628 11354
rect 31576 11290 31628 11296
rect 31392 11280 31444 11286
rect 31392 11222 31444 11228
rect 31484 11144 31536 11150
rect 31484 11086 31536 11092
rect 31392 10600 31444 10606
rect 31392 10542 31444 10548
rect 31300 10260 31352 10266
rect 31300 10202 31352 10208
rect 31404 9994 31432 10542
rect 31496 10538 31524 11086
rect 31588 10690 31616 11290
rect 31680 11082 31708 12106
rect 32508 11830 32536 12242
rect 32496 11824 32548 11830
rect 32496 11766 32548 11772
rect 32508 11558 32536 11766
rect 32496 11552 32548 11558
rect 32496 11494 32548 11500
rect 31668 11076 31720 11082
rect 31668 11018 31720 11024
rect 31588 10662 31800 10690
rect 31772 10606 31800 10662
rect 31760 10600 31812 10606
rect 31760 10542 31812 10548
rect 32220 10600 32272 10606
rect 32220 10542 32272 10548
rect 31484 10532 31536 10538
rect 31484 10474 31536 10480
rect 31392 9988 31444 9994
rect 31392 9930 31444 9936
rect 31404 9518 31432 9930
rect 31852 9716 31904 9722
rect 31852 9658 31904 9664
rect 31668 9580 31720 9586
rect 31668 9522 31720 9528
rect 31392 9512 31444 9518
rect 31392 9454 31444 9460
rect 31208 9104 31260 9110
rect 31208 9046 31260 9052
rect 31024 9036 31076 9042
rect 31024 8978 31076 8984
rect 31036 8634 31064 8978
rect 31300 8968 31352 8974
rect 31300 8910 31352 8916
rect 31024 8628 31076 8634
rect 31024 8570 31076 8576
rect 31312 8090 31340 8910
rect 31404 8430 31432 9454
rect 31484 9376 31536 9382
rect 31484 9318 31536 9324
rect 31496 9178 31524 9318
rect 31484 9172 31536 9178
rect 31484 9114 31536 9120
rect 31680 8906 31708 9522
rect 31668 8900 31720 8906
rect 31668 8842 31720 8848
rect 31864 8838 31892 9658
rect 32232 9518 32260 10542
rect 32784 10130 32812 17070
rect 33232 16652 33284 16658
rect 33232 16594 33284 16600
rect 32956 16040 33008 16046
rect 32956 15982 33008 15988
rect 32968 15570 32996 15982
rect 32956 15564 33008 15570
rect 32956 15506 33008 15512
rect 33140 15564 33192 15570
rect 33140 15506 33192 15512
rect 33152 15094 33180 15506
rect 33140 15088 33192 15094
rect 33140 15030 33192 15036
rect 33140 14952 33192 14958
rect 33140 14894 33192 14900
rect 32864 14544 32916 14550
rect 32864 14486 32916 14492
rect 32876 13462 32904 14486
rect 33152 13938 33180 14894
rect 33244 14414 33272 16594
rect 33324 14544 33376 14550
rect 33324 14486 33376 14492
rect 33232 14408 33284 14414
rect 33232 14350 33284 14356
rect 33140 13932 33192 13938
rect 33140 13874 33192 13880
rect 33244 13818 33272 14350
rect 33336 13870 33364 14486
rect 32968 13790 33272 13818
rect 33324 13864 33376 13870
rect 33324 13806 33376 13812
rect 32968 13734 32996 13790
rect 32956 13728 33008 13734
rect 32956 13670 33008 13676
rect 33140 13728 33192 13734
rect 33140 13670 33192 13676
rect 32864 13456 32916 13462
rect 32864 13398 32916 13404
rect 32876 10713 32904 13398
rect 32968 13394 32996 13670
rect 32956 13388 33008 13394
rect 32956 13330 33008 13336
rect 32956 13252 33008 13258
rect 32956 13194 33008 13200
rect 32968 12345 32996 13194
rect 33152 12782 33180 13670
rect 33336 12850 33364 13806
rect 33324 12844 33376 12850
rect 33324 12786 33376 12792
rect 33140 12776 33192 12782
rect 33140 12718 33192 12724
rect 33140 12640 33192 12646
rect 33140 12582 33192 12588
rect 32954 12336 33010 12345
rect 32954 12271 33010 12280
rect 33152 11218 33180 12582
rect 33324 11824 33376 11830
rect 33324 11766 33376 11772
rect 33232 11620 33284 11626
rect 33232 11562 33284 11568
rect 33140 11212 33192 11218
rect 33140 11154 33192 11160
rect 32862 10704 32918 10713
rect 32862 10639 32918 10648
rect 33244 10606 33272 11562
rect 33336 11218 33364 11766
rect 33324 11212 33376 11218
rect 33324 11154 33376 11160
rect 33232 10600 33284 10606
rect 33232 10542 33284 10548
rect 33140 10464 33192 10470
rect 33140 10406 33192 10412
rect 33232 10464 33284 10470
rect 33232 10406 33284 10412
rect 32312 10124 32364 10130
rect 32312 10066 32364 10072
rect 32680 10124 32732 10130
rect 32680 10066 32732 10072
rect 32772 10124 32824 10130
rect 32772 10066 32824 10072
rect 32324 9994 32352 10066
rect 32312 9988 32364 9994
rect 32312 9930 32364 9936
rect 32692 9722 32720 10066
rect 32680 9716 32732 9722
rect 32680 9658 32732 9664
rect 32220 9512 32272 9518
rect 32220 9454 32272 9460
rect 31944 9104 31996 9110
rect 31944 9046 31996 9052
rect 31852 8832 31904 8838
rect 31852 8774 31904 8780
rect 31392 8424 31444 8430
rect 31392 8366 31444 8372
rect 31300 8084 31352 8090
rect 31300 8026 31352 8032
rect 30944 7840 31064 7868
rect 30840 7472 30892 7478
rect 30840 7414 30892 7420
rect 31036 7410 31064 7840
rect 31024 7404 31076 7410
rect 31024 7346 31076 7352
rect 31576 7404 31628 7410
rect 31576 7346 31628 7352
rect 30932 7200 30984 7206
rect 30932 7142 30984 7148
rect 30564 6860 30616 6866
rect 30564 6802 30616 6808
rect 30944 6322 30972 7142
rect 30932 6316 30984 6322
rect 30932 6258 30984 6264
rect 30932 6180 30984 6186
rect 30932 6122 30984 6128
rect 30944 4146 30972 6122
rect 31036 5914 31064 7346
rect 31116 7268 31168 7274
rect 31116 7210 31168 7216
rect 31128 6866 31156 7210
rect 31588 7206 31616 7346
rect 31864 7342 31892 8774
rect 31956 8430 31984 9046
rect 32232 8430 32260 9454
rect 33152 9042 33180 10406
rect 33140 9036 33192 9042
rect 33140 8978 33192 8984
rect 33244 8566 33272 10406
rect 33232 8560 33284 8566
rect 33232 8502 33284 8508
rect 31944 8424 31996 8430
rect 31944 8366 31996 8372
rect 32220 8424 32272 8430
rect 32220 8366 32272 8372
rect 31852 7336 31904 7342
rect 31852 7278 31904 7284
rect 31576 7200 31628 7206
rect 31576 7142 31628 7148
rect 31116 6860 31168 6866
rect 31116 6802 31168 6808
rect 31760 6792 31812 6798
rect 31760 6734 31812 6740
rect 31484 6656 31536 6662
rect 31484 6598 31536 6604
rect 31496 6322 31524 6598
rect 31484 6316 31536 6322
rect 31484 6258 31536 6264
rect 31772 6186 31800 6734
rect 31956 6254 31984 8366
rect 33324 8288 33376 8294
rect 33324 8230 33376 8236
rect 32404 7880 32456 7886
rect 32404 7822 32456 7828
rect 32036 7336 32088 7342
rect 32036 7278 32088 7284
rect 32048 6866 32076 7278
rect 32036 6860 32088 6866
rect 32036 6802 32088 6808
rect 32416 6322 32444 7822
rect 33336 7342 33364 8230
rect 33428 7546 33456 20946
rect 33612 19938 33640 24074
rect 33784 23656 33836 23662
rect 33784 23598 33836 23604
rect 33796 23254 33824 23598
rect 33784 23248 33836 23254
rect 33784 23190 33836 23196
rect 33692 22636 33744 22642
rect 33692 22578 33744 22584
rect 33704 22166 33732 22578
rect 33692 22160 33744 22166
rect 33692 22102 33744 22108
rect 33692 21888 33744 21894
rect 33692 21830 33744 21836
rect 33520 19922 33640 19938
rect 33508 19916 33640 19922
rect 33560 19910 33640 19916
rect 33508 19858 33560 19864
rect 33520 18222 33548 19858
rect 33600 18284 33652 18290
rect 33600 18226 33652 18232
rect 33508 18216 33560 18222
rect 33508 18158 33560 18164
rect 33520 16590 33548 18158
rect 33612 17746 33640 18226
rect 33704 18222 33732 21830
rect 33796 21690 33824 23190
rect 33980 23066 34008 37266
rect 34520 36168 34572 36174
rect 34520 36110 34572 36116
rect 34532 35222 34560 36110
rect 34520 35216 34572 35222
rect 34520 35158 34572 35164
rect 34520 34060 34572 34066
rect 34520 34002 34572 34008
rect 34532 33454 34560 34002
rect 34520 33448 34572 33454
rect 34520 33390 34572 33396
rect 34532 32910 34560 33390
rect 34520 32904 34572 32910
rect 34520 32846 34572 32852
rect 34532 32230 34560 32846
rect 34520 32224 34572 32230
rect 34520 32166 34572 32172
rect 34532 31890 34560 32166
rect 34520 31884 34572 31890
rect 34520 31826 34572 31832
rect 34244 30728 34296 30734
rect 34244 30670 34296 30676
rect 34256 30598 34284 30670
rect 34244 30592 34296 30598
rect 34244 30534 34296 30540
rect 34256 30258 34284 30534
rect 34244 30252 34296 30258
rect 34244 30194 34296 30200
rect 34532 29646 34560 31826
rect 34520 29640 34572 29646
rect 34520 29582 34572 29588
rect 34244 28416 34296 28422
rect 34244 28358 34296 28364
rect 34060 27940 34112 27946
rect 34060 27882 34112 27888
rect 34072 27470 34100 27882
rect 34060 27464 34112 27470
rect 34060 27406 34112 27412
rect 34072 25838 34100 27406
rect 34256 26994 34284 28358
rect 34520 28008 34572 28014
rect 34520 27950 34572 27956
rect 34336 27940 34388 27946
rect 34336 27882 34388 27888
rect 34348 27538 34376 27882
rect 34532 27674 34560 27950
rect 34520 27668 34572 27674
rect 34520 27610 34572 27616
rect 34336 27532 34388 27538
rect 34336 27474 34388 27480
rect 34520 27124 34572 27130
rect 34520 27066 34572 27072
rect 34244 26988 34296 26994
rect 34244 26930 34296 26936
rect 34060 25832 34112 25838
rect 34060 25774 34112 25780
rect 34072 25498 34100 25774
rect 34060 25492 34112 25498
rect 34060 25434 34112 25440
rect 34336 25356 34388 25362
rect 34336 25298 34388 25304
rect 34348 24070 34376 25298
rect 34532 24682 34560 27066
rect 34624 26874 34652 37810
rect 34940 37020 35236 37040
rect 34996 37018 35020 37020
rect 35076 37018 35100 37020
rect 35156 37018 35180 37020
rect 35018 36966 35020 37018
rect 35082 36966 35094 37018
rect 35156 36966 35158 37018
rect 34996 36964 35020 36966
rect 35076 36964 35100 36966
rect 35156 36964 35180 36966
rect 34940 36944 35236 36964
rect 35268 36786 35296 38270
rect 35256 36780 35308 36786
rect 35256 36722 35308 36728
rect 35624 36032 35676 36038
rect 35624 35974 35676 35980
rect 34940 35932 35236 35952
rect 34996 35930 35020 35932
rect 35076 35930 35100 35932
rect 35156 35930 35180 35932
rect 35018 35878 35020 35930
rect 35082 35878 35094 35930
rect 35156 35878 35158 35930
rect 34996 35876 35020 35878
rect 35076 35876 35100 35878
rect 35156 35876 35180 35878
rect 34940 35856 35236 35876
rect 35636 34950 35664 35974
rect 35990 35456 36046 35465
rect 35990 35391 36046 35400
rect 36004 35290 36032 35391
rect 35992 35284 36044 35290
rect 35992 35226 36044 35232
rect 35624 34944 35676 34950
rect 35624 34886 35676 34892
rect 34940 34844 35236 34864
rect 34996 34842 35020 34844
rect 35076 34842 35100 34844
rect 35156 34842 35180 34844
rect 35018 34790 35020 34842
rect 35082 34790 35094 34842
rect 35156 34790 35158 34842
rect 34996 34788 35020 34790
rect 35076 34788 35100 34790
rect 35156 34788 35180 34790
rect 34940 34768 35236 34788
rect 34888 34604 34940 34610
rect 34888 34546 34940 34552
rect 34796 34536 34848 34542
rect 34796 34478 34848 34484
rect 34808 32978 34836 34478
rect 34900 34202 34928 34546
rect 34980 34536 35032 34542
rect 34980 34478 35032 34484
rect 34888 34196 34940 34202
rect 34888 34138 34940 34144
rect 34992 34134 35020 34478
rect 35256 34468 35308 34474
rect 35256 34410 35308 34416
rect 34980 34128 35032 34134
rect 34980 34070 35032 34076
rect 34940 33756 35236 33776
rect 34996 33754 35020 33756
rect 35076 33754 35100 33756
rect 35156 33754 35180 33756
rect 35018 33702 35020 33754
rect 35082 33702 35094 33754
rect 35156 33702 35158 33754
rect 34996 33700 35020 33702
rect 35076 33700 35100 33702
rect 35156 33700 35180 33702
rect 34940 33680 35236 33700
rect 35268 33522 35296 34410
rect 36096 34066 36124 38655
rect 37200 38010 37228 40200
rect 37188 38004 37240 38010
rect 37188 37946 37240 37952
rect 39408 37398 39436 40200
rect 39396 37392 39448 37398
rect 39396 37334 39448 37340
rect 36176 34672 36228 34678
rect 36176 34614 36228 34620
rect 36084 34060 36136 34066
rect 36084 34002 36136 34008
rect 35256 33516 35308 33522
rect 35256 33458 35308 33464
rect 34796 32972 34848 32978
rect 34796 32914 34848 32920
rect 34940 32668 35236 32688
rect 34996 32666 35020 32668
rect 35076 32666 35100 32668
rect 35156 32666 35180 32668
rect 35018 32614 35020 32666
rect 35082 32614 35094 32666
rect 35156 32614 35158 32666
rect 34996 32612 35020 32614
rect 35076 32612 35100 32614
rect 35156 32612 35180 32614
rect 34940 32592 35236 32612
rect 36096 32450 36124 34002
rect 36188 32473 36216 34614
rect 37004 33380 37056 33386
rect 37004 33322 37056 33328
rect 36268 32768 36320 32774
rect 36268 32710 36320 32716
rect 36004 32422 36124 32450
rect 36174 32464 36230 32473
rect 34796 32360 34848 32366
rect 34796 32302 34848 32308
rect 34704 31816 34756 31822
rect 34704 31758 34756 31764
rect 34716 30938 34744 31758
rect 34808 31482 34836 32302
rect 35808 32292 35860 32298
rect 35808 32234 35860 32240
rect 34940 31580 35236 31600
rect 34996 31578 35020 31580
rect 35076 31578 35100 31580
rect 35156 31578 35180 31580
rect 35018 31526 35020 31578
rect 35082 31526 35094 31578
rect 35156 31526 35158 31578
rect 34996 31524 35020 31526
rect 35076 31524 35100 31526
rect 35156 31524 35180 31526
rect 34940 31504 35236 31524
rect 34796 31476 34848 31482
rect 34796 31418 34848 31424
rect 34888 31408 34940 31414
rect 34888 31350 34940 31356
rect 34796 31272 34848 31278
rect 34796 31214 34848 31220
rect 34704 30932 34756 30938
rect 34704 30874 34756 30880
rect 34704 30116 34756 30122
rect 34704 30058 34756 30064
rect 34716 29238 34744 30058
rect 34808 29850 34836 31214
rect 34900 30802 34928 31350
rect 35820 31278 35848 32234
rect 35808 31272 35860 31278
rect 35808 31214 35860 31220
rect 35900 31204 35952 31210
rect 35900 31146 35952 31152
rect 34888 30796 34940 30802
rect 34888 30738 34940 30744
rect 34940 30492 35236 30512
rect 34996 30490 35020 30492
rect 35076 30490 35100 30492
rect 35156 30490 35180 30492
rect 35018 30438 35020 30490
rect 35082 30438 35094 30490
rect 35156 30438 35158 30490
rect 34996 30436 35020 30438
rect 35076 30436 35100 30438
rect 35156 30436 35180 30438
rect 34940 30416 35236 30436
rect 35912 30326 35940 31146
rect 35900 30320 35952 30326
rect 35900 30262 35952 30268
rect 35256 30184 35308 30190
rect 35256 30126 35308 30132
rect 34796 29844 34848 29850
rect 34796 29786 34848 29792
rect 34704 29232 34756 29238
rect 34704 29174 34756 29180
rect 34808 29102 34836 29786
rect 34940 29404 35236 29424
rect 34996 29402 35020 29404
rect 35076 29402 35100 29404
rect 35156 29402 35180 29404
rect 35018 29350 35020 29402
rect 35082 29350 35094 29402
rect 35156 29350 35158 29402
rect 34996 29348 35020 29350
rect 35076 29348 35100 29350
rect 35156 29348 35180 29350
rect 34940 29328 35236 29348
rect 34796 29096 34848 29102
rect 34796 29038 34848 29044
rect 35268 28694 35296 30126
rect 35716 30116 35768 30122
rect 35716 30058 35768 30064
rect 35728 29102 35756 30058
rect 35716 29096 35768 29102
rect 35716 29038 35768 29044
rect 35912 29034 35940 30262
rect 35900 29028 35952 29034
rect 35900 28970 35952 28976
rect 35624 28756 35676 28762
rect 35624 28698 35676 28704
rect 35256 28688 35308 28694
rect 35256 28630 35308 28636
rect 34940 28316 35236 28336
rect 34996 28314 35020 28316
rect 35076 28314 35100 28316
rect 35156 28314 35180 28316
rect 35018 28262 35020 28314
rect 35082 28262 35094 28314
rect 35156 28262 35158 28314
rect 34996 28260 35020 28262
rect 35076 28260 35100 28262
rect 35156 28260 35180 28262
rect 34940 28240 35236 28260
rect 35268 27606 35296 28630
rect 35348 28076 35400 28082
rect 35348 28018 35400 28024
rect 35256 27600 35308 27606
rect 35256 27542 35308 27548
rect 35360 27538 35388 28018
rect 35532 28008 35584 28014
rect 35532 27950 35584 27956
rect 35348 27532 35400 27538
rect 35348 27474 35400 27480
rect 34940 27228 35236 27248
rect 34996 27226 35020 27228
rect 35076 27226 35100 27228
rect 35156 27226 35180 27228
rect 35018 27174 35020 27226
rect 35082 27174 35094 27226
rect 35156 27174 35158 27226
rect 34996 27172 35020 27174
rect 35076 27172 35100 27174
rect 35156 27172 35180 27174
rect 34940 27152 35236 27172
rect 34796 26920 34848 26926
rect 34624 26846 34744 26874
rect 34796 26862 34848 26868
rect 34612 26240 34664 26246
rect 34612 26182 34664 26188
rect 34624 25430 34652 26182
rect 34612 25424 34664 25430
rect 34612 25366 34664 25372
rect 34612 24812 34664 24818
rect 34612 24754 34664 24760
rect 34520 24676 34572 24682
rect 34520 24618 34572 24624
rect 34532 24290 34560 24618
rect 34440 24262 34560 24290
rect 34336 24064 34388 24070
rect 34336 24006 34388 24012
rect 34244 23588 34296 23594
rect 34244 23530 34296 23536
rect 34256 23186 34284 23530
rect 34348 23254 34376 24006
rect 34440 23798 34468 24262
rect 34520 24200 34572 24206
rect 34520 24142 34572 24148
rect 34428 23792 34480 23798
rect 34428 23734 34480 23740
rect 34532 23594 34560 24142
rect 34520 23588 34572 23594
rect 34520 23530 34572 23536
rect 34336 23248 34388 23254
rect 34336 23190 34388 23196
rect 34624 23186 34652 24754
rect 34244 23180 34296 23186
rect 34244 23122 34296 23128
rect 34612 23180 34664 23186
rect 34612 23122 34664 23128
rect 33888 23038 34008 23066
rect 33784 21684 33836 21690
rect 33784 21626 33836 21632
rect 33796 21078 33824 21626
rect 33784 21072 33836 21078
rect 33784 21014 33836 21020
rect 33784 20256 33836 20262
rect 33784 20198 33836 20204
rect 33692 18216 33744 18222
rect 33692 18158 33744 18164
rect 33704 17746 33732 18158
rect 33600 17740 33652 17746
rect 33600 17682 33652 17688
rect 33692 17740 33744 17746
rect 33692 17682 33744 17688
rect 33704 16794 33732 17682
rect 33692 16788 33744 16794
rect 33692 16730 33744 16736
rect 33508 16584 33560 16590
rect 33508 16526 33560 16532
rect 33508 16448 33560 16454
rect 33508 16390 33560 16396
rect 33520 15638 33548 16390
rect 33692 16040 33744 16046
rect 33796 16028 33824 20198
rect 33888 16697 33916 23038
rect 34612 22976 34664 22982
rect 34612 22918 34664 22924
rect 34520 22704 34572 22710
rect 34520 22646 34572 22652
rect 34336 21344 34388 21350
rect 34336 21286 34388 21292
rect 34348 21010 34376 21286
rect 34532 21026 34560 22646
rect 34624 22574 34652 22918
rect 34612 22568 34664 22574
rect 34612 22510 34664 22516
rect 34612 22024 34664 22030
rect 34612 21966 34664 21972
rect 34336 21004 34388 21010
rect 34336 20946 34388 20952
rect 34440 20998 34560 21026
rect 34060 20392 34112 20398
rect 34112 20352 34192 20380
rect 34060 20334 34112 20340
rect 33968 19916 34020 19922
rect 33968 19858 34020 19864
rect 33980 19786 34008 19858
rect 33968 19780 34020 19786
rect 33968 19722 34020 19728
rect 33980 19378 34008 19722
rect 33968 19372 34020 19378
rect 33968 19314 34020 19320
rect 34164 18970 34192 20352
rect 34348 19990 34376 20946
rect 34440 20346 34468 20998
rect 34520 20936 34572 20942
rect 34520 20878 34572 20884
rect 34532 20466 34560 20878
rect 34520 20460 34572 20466
rect 34520 20402 34572 20408
rect 34440 20330 34560 20346
rect 34440 20324 34572 20330
rect 34440 20318 34520 20324
rect 34520 20266 34572 20272
rect 34336 19984 34388 19990
rect 34336 19926 34388 19932
rect 34532 19378 34560 20266
rect 34520 19372 34572 19378
rect 34520 19314 34572 19320
rect 34152 18964 34204 18970
rect 34152 18906 34204 18912
rect 33968 16992 34020 16998
rect 33968 16934 34020 16940
rect 33874 16688 33930 16697
rect 33874 16623 33930 16632
rect 33796 16000 33916 16028
rect 33692 15982 33744 15988
rect 33508 15632 33560 15638
rect 33508 15574 33560 15580
rect 33600 14408 33652 14414
rect 33600 14350 33652 14356
rect 33508 13864 33560 13870
rect 33508 13806 33560 13812
rect 33520 13462 33548 13806
rect 33508 13456 33560 13462
rect 33508 13398 33560 13404
rect 33508 12844 33560 12850
rect 33508 12786 33560 12792
rect 33520 12646 33548 12786
rect 33508 12640 33560 12646
rect 33508 12582 33560 12588
rect 33506 12200 33562 12209
rect 33506 12135 33562 12144
rect 33520 12102 33548 12135
rect 33508 12096 33560 12102
rect 33508 12038 33560 12044
rect 33612 11694 33640 14350
rect 33704 14346 33732 15982
rect 33784 15904 33836 15910
rect 33784 15846 33836 15852
rect 33796 15570 33824 15846
rect 33784 15564 33836 15570
rect 33784 15506 33836 15512
rect 33888 15450 33916 16000
rect 33796 15422 33916 15450
rect 33692 14340 33744 14346
rect 33692 14282 33744 14288
rect 33796 13734 33824 15422
rect 33980 14890 34008 16934
rect 34060 16720 34112 16726
rect 34060 16662 34112 16668
rect 33968 14884 34020 14890
rect 33968 14826 34020 14832
rect 33980 14482 34008 14826
rect 33968 14476 34020 14482
rect 33968 14418 34020 14424
rect 33876 13864 33928 13870
rect 33876 13806 33928 13812
rect 33784 13728 33836 13734
rect 33784 13670 33836 13676
rect 33888 13530 33916 13806
rect 33692 13524 33744 13530
rect 33692 13466 33744 13472
rect 33876 13524 33928 13530
rect 33876 13466 33928 13472
rect 33600 11688 33652 11694
rect 33600 11630 33652 11636
rect 33704 10606 33732 13466
rect 33968 13456 34020 13462
rect 33968 13398 34020 13404
rect 33784 13388 33836 13394
rect 33784 13330 33836 13336
rect 33796 12986 33824 13330
rect 33784 12980 33836 12986
rect 33784 12922 33836 12928
rect 33980 12918 34008 13398
rect 33968 12912 34020 12918
rect 33888 12860 33968 12866
rect 33888 12854 34020 12860
rect 33888 12838 34008 12854
rect 33784 12708 33836 12714
rect 33784 12650 33836 12656
rect 33796 12442 33824 12650
rect 33784 12436 33836 12442
rect 33784 12378 33836 12384
rect 33888 12209 33916 12838
rect 33980 12789 34008 12838
rect 33968 12708 34020 12714
rect 33968 12650 34020 12656
rect 33980 12306 34008 12650
rect 33968 12300 34020 12306
rect 33968 12242 34020 12248
rect 33874 12200 33930 12209
rect 33784 12164 33836 12170
rect 33874 12135 33930 12144
rect 33968 12164 34020 12170
rect 33784 12106 33836 12112
rect 33968 12106 34020 12112
rect 33796 11286 33824 12106
rect 33876 11824 33928 11830
rect 33876 11766 33928 11772
rect 33784 11280 33836 11286
rect 33784 11222 33836 11228
rect 33508 10600 33560 10606
rect 33508 10542 33560 10548
rect 33692 10600 33744 10606
rect 33692 10542 33744 10548
rect 33520 10266 33548 10542
rect 33508 10260 33560 10266
rect 33508 10202 33560 10208
rect 33784 10124 33836 10130
rect 33784 10066 33836 10072
rect 33796 9722 33824 10066
rect 33784 9716 33836 9722
rect 33784 9658 33836 9664
rect 33508 8968 33560 8974
rect 33508 8910 33560 8916
rect 33520 7954 33548 8910
rect 33796 8430 33824 9658
rect 33888 8430 33916 11766
rect 33980 9518 34008 12106
rect 34072 9654 34100 16662
rect 34060 9648 34112 9654
rect 34060 9590 34112 9596
rect 33968 9512 34020 9518
rect 33968 9454 34020 9460
rect 34060 9512 34112 9518
rect 34164 9500 34192 18906
rect 34520 18828 34572 18834
rect 34520 18770 34572 18776
rect 34336 18352 34388 18358
rect 34336 18294 34388 18300
rect 34348 17270 34376 18294
rect 34428 18284 34480 18290
rect 34428 18226 34480 18232
rect 34336 17264 34388 17270
rect 34336 17206 34388 17212
rect 34348 16114 34376 17206
rect 34336 16108 34388 16114
rect 34336 16050 34388 16056
rect 34440 15502 34468 18226
rect 34532 18154 34560 18770
rect 34624 18766 34652 21966
rect 34716 21570 34744 26846
rect 34808 25362 34836 26862
rect 35544 26450 35572 27950
rect 35532 26444 35584 26450
rect 35532 26386 35584 26392
rect 34940 26140 35236 26160
rect 34996 26138 35020 26140
rect 35076 26138 35100 26140
rect 35156 26138 35180 26140
rect 35018 26086 35020 26138
rect 35082 26086 35094 26138
rect 35156 26086 35158 26138
rect 34996 26084 35020 26086
rect 35076 26084 35100 26086
rect 35156 26084 35180 26086
rect 34940 26064 35236 26084
rect 35544 25906 35572 26386
rect 35636 26042 35664 28698
rect 35716 28620 35768 28626
rect 35716 28562 35768 28568
rect 35728 27334 35756 28562
rect 35808 28212 35860 28218
rect 35912 28200 35940 28970
rect 35860 28172 35940 28200
rect 35808 28154 35860 28160
rect 35716 27328 35768 27334
rect 35716 27270 35768 27276
rect 35808 27328 35860 27334
rect 35808 27270 35860 27276
rect 35624 26036 35676 26042
rect 35624 25978 35676 25984
rect 35532 25900 35584 25906
rect 35532 25842 35584 25848
rect 35164 25832 35216 25838
rect 35164 25774 35216 25780
rect 35176 25430 35204 25774
rect 35164 25424 35216 25430
rect 35164 25366 35216 25372
rect 35636 25362 35664 25978
rect 34796 25356 34848 25362
rect 34796 25298 34848 25304
rect 35440 25356 35492 25362
rect 35440 25298 35492 25304
rect 35624 25356 35676 25362
rect 35624 25298 35676 25304
rect 34808 21894 34836 25298
rect 34940 25052 35236 25072
rect 34996 25050 35020 25052
rect 35076 25050 35100 25052
rect 35156 25050 35180 25052
rect 35018 24998 35020 25050
rect 35082 24998 35094 25050
rect 35156 24998 35158 25050
rect 34996 24996 35020 24998
rect 35076 24996 35100 24998
rect 35156 24996 35180 24998
rect 34940 24976 35236 24996
rect 35452 24818 35480 25298
rect 34888 24812 34940 24818
rect 34888 24754 34940 24760
rect 35440 24812 35492 24818
rect 35440 24754 35492 24760
rect 34900 24342 34928 24754
rect 35728 24750 35756 27270
rect 35820 27130 35848 27270
rect 35808 27124 35860 27130
rect 35808 27066 35860 27072
rect 35808 26784 35860 26790
rect 35808 26726 35860 26732
rect 35820 26450 35848 26726
rect 35808 26444 35860 26450
rect 35808 26386 35860 26392
rect 35898 26208 35954 26217
rect 35898 26143 35954 26152
rect 35256 24744 35308 24750
rect 35256 24686 35308 24692
rect 35716 24744 35768 24750
rect 35716 24686 35768 24692
rect 35072 24676 35124 24682
rect 35072 24618 35124 24624
rect 34888 24336 34940 24342
rect 34888 24278 34940 24284
rect 35084 24274 35112 24618
rect 35072 24268 35124 24274
rect 35072 24210 35124 24216
rect 34940 23964 35236 23984
rect 34996 23962 35020 23964
rect 35076 23962 35100 23964
rect 35156 23962 35180 23964
rect 35018 23910 35020 23962
rect 35082 23910 35094 23962
rect 35156 23910 35158 23962
rect 34996 23908 35020 23910
rect 35076 23908 35100 23910
rect 35156 23908 35180 23910
rect 34940 23888 35236 23908
rect 35164 23792 35216 23798
rect 35164 23734 35216 23740
rect 35176 23100 35204 23734
rect 35268 23254 35296 24686
rect 35912 24410 35940 26143
rect 35900 24404 35952 24410
rect 35900 24346 35952 24352
rect 35348 24268 35400 24274
rect 35348 24210 35400 24216
rect 35532 24268 35584 24274
rect 35532 24210 35584 24216
rect 35256 23248 35308 23254
rect 35256 23190 35308 23196
rect 35176 23072 35296 23100
rect 34940 22876 35236 22896
rect 34996 22874 35020 22876
rect 35076 22874 35100 22876
rect 35156 22874 35180 22876
rect 35018 22822 35020 22874
rect 35082 22822 35094 22874
rect 35156 22822 35158 22874
rect 34996 22820 35020 22822
rect 35076 22820 35100 22822
rect 35156 22820 35180 22822
rect 34940 22800 35236 22820
rect 35164 22568 35216 22574
rect 35164 22510 35216 22516
rect 35072 22092 35124 22098
rect 35072 22034 35124 22040
rect 35084 21978 35112 22034
rect 35176 22030 35204 22510
rect 35268 22098 35296 23072
rect 35360 22982 35388 24210
rect 35544 23662 35572 24210
rect 35532 23656 35584 23662
rect 35532 23598 35584 23604
rect 35440 23520 35492 23526
rect 35440 23462 35492 23468
rect 35452 23118 35480 23462
rect 35544 23186 35572 23598
rect 35624 23588 35676 23594
rect 35624 23530 35676 23536
rect 35532 23180 35584 23186
rect 35532 23122 35584 23128
rect 35440 23112 35492 23118
rect 35440 23054 35492 23060
rect 35348 22976 35400 22982
rect 35348 22918 35400 22924
rect 35452 22098 35480 23054
rect 35256 22092 35308 22098
rect 35256 22034 35308 22040
rect 35440 22092 35492 22098
rect 35440 22034 35492 22040
rect 34900 21962 35112 21978
rect 35164 22024 35216 22030
rect 35164 21966 35216 21972
rect 34888 21956 35112 21962
rect 34940 21950 35112 21956
rect 34888 21898 34940 21904
rect 34796 21888 34848 21894
rect 34796 21830 34848 21836
rect 34808 21690 34836 21830
rect 34940 21788 35236 21808
rect 34996 21786 35020 21788
rect 35076 21786 35100 21788
rect 35156 21786 35180 21788
rect 35018 21734 35020 21786
rect 35082 21734 35094 21786
rect 35156 21734 35158 21786
rect 34996 21732 35020 21734
rect 35076 21732 35100 21734
rect 35156 21732 35180 21734
rect 34940 21712 35236 21732
rect 34796 21684 34848 21690
rect 34796 21626 34848 21632
rect 35268 21570 35296 22034
rect 34716 21542 34836 21570
rect 34808 19802 34836 21542
rect 34992 21542 35296 21570
rect 34992 21010 35020 21542
rect 35256 21412 35308 21418
rect 35256 21354 35308 21360
rect 34980 21004 35032 21010
rect 34980 20946 35032 20952
rect 34940 20700 35236 20720
rect 34996 20698 35020 20700
rect 35076 20698 35100 20700
rect 35156 20698 35180 20700
rect 35018 20646 35020 20698
rect 35082 20646 35094 20698
rect 35156 20646 35158 20698
rect 34996 20644 35020 20646
rect 35076 20644 35100 20646
rect 35156 20644 35180 20646
rect 34940 20624 35236 20644
rect 35268 20398 35296 21354
rect 35348 21004 35400 21010
rect 35348 20946 35400 20952
rect 35360 20534 35388 20946
rect 35440 20936 35492 20942
rect 35440 20878 35492 20884
rect 35348 20528 35400 20534
rect 35348 20470 35400 20476
rect 35256 20392 35308 20398
rect 35256 20334 35308 20340
rect 35452 19922 35480 20878
rect 35440 19916 35492 19922
rect 35440 19858 35492 19864
rect 35544 19854 35572 23122
rect 35636 20058 35664 23530
rect 35716 22976 35768 22982
rect 35716 22918 35768 22924
rect 35898 22944 35954 22953
rect 35728 21486 35756 22918
rect 35898 22879 35954 22888
rect 35912 22234 35940 22879
rect 35900 22228 35952 22234
rect 35900 22170 35952 22176
rect 35716 21480 35768 21486
rect 35716 21422 35768 21428
rect 35808 21480 35860 21486
rect 35808 21422 35860 21428
rect 35716 21140 35768 21146
rect 35716 21082 35768 21088
rect 35624 20052 35676 20058
rect 35624 19994 35676 20000
rect 35532 19848 35584 19854
rect 34808 19774 35480 19802
rect 35532 19790 35584 19796
rect 35348 19712 35400 19718
rect 35348 19654 35400 19660
rect 34940 19612 35236 19632
rect 34996 19610 35020 19612
rect 35076 19610 35100 19612
rect 35156 19610 35180 19612
rect 35018 19558 35020 19610
rect 35082 19558 35094 19610
rect 35156 19558 35158 19610
rect 34996 19556 35020 19558
rect 35076 19556 35100 19558
rect 35156 19556 35180 19558
rect 34940 19536 35236 19556
rect 34796 19508 34848 19514
rect 34796 19450 34848 19456
rect 34808 18902 34836 19450
rect 34796 18896 34848 18902
rect 34796 18838 34848 18844
rect 34704 18828 34756 18834
rect 34704 18770 34756 18776
rect 34612 18760 34664 18766
rect 34612 18702 34664 18708
rect 34520 18148 34572 18154
rect 34520 18090 34572 18096
rect 34532 17814 34560 18090
rect 34520 17808 34572 17814
rect 34520 17750 34572 17756
rect 34612 17740 34664 17746
rect 34612 17682 34664 17688
rect 34624 17338 34652 17682
rect 34612 17332 34664 17338
rect 34612 17274 34664 17280
rect 34520 17128 34572 17134
rect 34520 17070 34572 17076
rect 34244 15496 34296 15502
rect 34244 15438 34296 15444
rect 34428 15496 34480 15502
rect 34428 15438 34480 15444
rect 34256 14362 34284 15438
rect 34428 14952 34480 14958
rect 34428 14894 34480 14900
rect 34336 14816 34388 14822
rect 34336 14758 34388 14764
rect 34348 14550 34376 14758
rect 34336 14544 34388 14550
rect 34336 14486 34388 14492
rect 34336 14408 34388 14414
rect 34256 14356 34336 14362
rect 34256 14350 34388 14356
rect 34256 14334 34376 14350
rect 34348 14074 34376 14334
rect 34336 14068 34388 14074
rect 34336 14010 34388 14016
rect 34336 13728 34388 13734
rect 34336 13670 34388 13676
rect 34348 12442 34376 13670
rect 34440 12753 34468 14894
rect 34532 13433 34560 17070
rect 34612 16992 34664 16998
rect 34612 16934 34664 16940
rect 34624 16658 34652 16934
rect 34612 16652 34664 16658
rect 34612 16594 34664 16600
rect 34612 14476 34664 14482
rect 34612 14418 34664 14424
rect 34624 13734 34652 14418
rect 34612 13728 34664 13734
rect 34612 13670 34664 13676
rect 34624 13530 34652 13670
rect 34612 13524 34664 13530
rect 34612 13466 34664 13472
rect 34518 13424 34574 13433
rect 34518 13359 34574 13368
rect 34612 13320 34664 13326
rect 34612 13262 34664 13268
rect 34520 12844 34572 12850
rect 34520 12786 34572 12792
rect 34426 12744 34482 12753
rect 34426 12679 34482 12688
rect 34428 12640 34480 12646
rect 34428 12582 34480 12588
rect 34440 12442 34468 12582
rect 34336 12436 34388 12442
rect 34336 12378 34388 12384
rect 34428 12436 34480 12442
rect 34428 12378 34480 12384
rect 34428 12232 34480 12238
rect 34428 12174 34480 12180
rect 34440 11830 34468 12174
rect 34532 12102 34560 12786
rect 34624 12306 34652 13262
rect 34612 12300 34664 12306
rect 34612 12242 34664 12248
rect 34716 12186 34744 18770
rect 34940 18524 35236 18544
rect 34996 18522 35020 18524
rect 35076 18522 35100 18524
rect 35156 18522 35180 18524
rect 35018 18470 35020 18522
rect 35082 18470 35094 18522
rect 35156 18470 35158 18522
rect 34996 18468 35020 18470
rect 35076 18468 35100 18470
rect 35156 18468 35180 18470
rect 34940 18448 35236 18468
rect 34796 18216 34848 18222
rect 34796 18158 34848 18164
rect 34808 17746 34836 18158
rect 35360 17882 35388 19654
rect 35348 17876 35400 17882
rect 35348 17818 35400 17824
rect 34796 17740 34848 17746
rect 34796 17682 34848 17688
rect 34808 17542 34836 17682
rect 34796 17536 34848 17542
rect 34796 17478 34848 17484
rect 34940 17436 35236 17456
rect 34996 17434 35020 17436
rect 35076 17434 35100 17436
rect 35156 17434 35180 17436
rect 35018 17382 35020 17434
rect 35082 17382 35094 17434
rect 35156 17382 35158 17434
rect 34996 17380 35020 17382
rect 35076 17380 35100 17382
rect 35156 17380 35180 17382
rect 34940 17360 35236 17380
rect 35360 17134 35388 17818
rect 35348 17128 35400 17134
rect 35348 17070 35400 17076
rect 34978 16824 35034 16833
rect 34978 16759 34980 16768
rect 35032 16759 35034 16768
rect 34980 16730 35032 16736
rect 34940 16348 35236 16368
rect 34996 16346 35020 16348
rect 35076 16346 35100 16348
rect 35156 16346 35180 16348
rect 35018 16294 35020 16346
rect 35082 16294 35094 16346
rect 35156 16294 35158 16346
rect 34996 16292 35020 16294
rect 35076 16292 35100 16294
rect 35156 16292 35180 16294
rect 34940 16272 35236 16292
rect 35360 15994 35388 17070
rect 35452 16046 35480 19774
rect 35544 19514 35572 19790
rect 35532 19508 35584 19514
rect 35532 19450 35584 19456
rect 35728 18426 35756 21082
rect 35820 19174 35848 21422
rect 35900 20936 35952 20942
rect 35900 20878 35952 20884
rect 35912 20466 35940 20878
rect 35900 20460 35952 20466
rect 35900 20402 35952 20408
rect 36004 19922 36032 32422
rect 36174 32399 36230 32408
rect 36280 32366 36308 32710
rect 36084 32360 36136 32366
rect 36084 32302 36136 32308
rect 36268 32360 36320 32366
rect 36268 32302 36320 32308
rect 36096 31686 36124 32302
rect 36176 32224 36228 32230
rect 36176 32166 36228 32172
rect 36544 32224 36596 32230
rect 36544 32166 36596 32172
rect 36188 31958 36216 32166
rect 36176 31952 36228 31958
rect 36176 31894 36228 31900
rect 36084 31680 36136 31686
rect 36084 31622 36136 31628
rect 36096 31278 36124 31622
rect 36084 31272 36136 31278
rect 36084 31214 36136 31220
rect 36084 30728 36136 30734
rect 36084 30670 36136 30676
rect 36096 30258 36124 30670
rect 36084 30252 36136 30258
rect 36084 30194 36136 30200
rect 36556 29594 36584 32166
rect 36636 31884 36688 31890
rect 36636 31826 36688 31832
rect 36372 29566 36584 29594
rect 36372 29050 36400 29566
rect 36544 29504 36596 29510
rect 36544 29446 36596 29452
rect 36372 29022 36492 29050
rect 36464 28966 36492 29022
rect 36452 28960 36504 28966
rect 36452 28902 36504 28908
rect 36556 28626 36584 29446
rect 36648 28694 36676 31826
rect 36820 31816 36872 31822
rect 36820 31758 36872 31764
rect 36728 31680 36780 31686
rect 36728 31622 36780 31628
rect 36740 30802 36768 31622
rect 36832 31278 36860 31758
rect 36820 31272 36872 31278
rect 36820 31214 36872 31220
rect 36728 30796 36780 30802
rect 36728 30738 36780 30744
rect 36832 30190 36860 31214
rect 36820 30184 36872 30190
rect 36820 30126 36872 30132
rect 36820 29708 36872 29714
rect 36820 29650 36872 29656
rect 36832 29102 36860 29650
rect 36820 29096 36872 29102
rect 36820 29038 36872 29044
rect 36728 28960 36780 28966
rect 36728 28902 36780 28908
rect 36636 28688 36688 28694
rect 36636 28630 36688 28636
rect 36360 28620 36412 28626
rect 36360 28562 36412 28568
rect 36544 28620 36596 28626
rect 36544 28562 36596 28568
rect 36372 24750 36400 28562
rect 36740 28370 36768 28902
rect 36648 28342 36768 28370
rect 36648 27674 36676 28342
rect 36832 28218 36860 29038
rect 36820 28212 36872 28218
rect 36820 28154 36872 28160
rect 36636 27668 36688 27674
rect 36636 27610 36688 27616
rect 36452 27464 36504 27470
rect 36452 27406 36504 27412
rect 36464 25140 36492 27406
rect 36648 26926 36676 27610
rect 36728 27600 36780 27606
rect 36728 27542 36780 27548
rect 36636 26920 36688 26926
rect 36636 26862 36688 26868
rect 36544 26240 36596 26246
rect 36544 26182 36596 26188
rect 36556 25362 36584 26182
rect 36648 25362 36676 26862
rect 36740 26246 36768 27542
rect 37016 26874 37044 33322
rect 39120 32972 39172 32978
rect 39120 32914 39172 32920
rect 38200 32768 38252 32774
rect 38200 32710 38252 32716
rect 37096 31952 37148 31958
rect 37096 31894 37148 31900
rect 37108 29238 37136 31894
rect 38016 31680 38068 31686
rect 38016 31622 38068 31628
rect 37740 31272 37792 31278
rect 37740 31214 37792 31220
rect 37464 30796 37516 30802
rect 37464 30738 37516 30744
rect 37476 30394 37504 30738
rect 37464 30388 37516 30394
rect 37464 30330 37516 30336
rect 37476 29782 37504 30330
rect 37752 30326 37780 31214
rect 37924 30796 37976 30802
rect 37924 30738 37976 30744
rect 37740 30320 37792 30326
rect 37740 30262 37792 30268
rect 37464 29776 37516 29782
rect 37464 29718 37516 29724
rect 37096 29232 37148 29238
rect 37096 29174 37148 29180
rect 37476 29102 37504 29718
rect 37936 29102 37964 30738
rect 38028 30734 38056 31622
rect 38016 30728 38068 30734
rect 38016 30670 38068 30676
rect 38108 30184 38160 30190
rect 38108 30126 38160 30132
rect 38120 29714 38148 30126
rect 38108 29708 38160 29714
rect 38108 29650 38160 29656
rect 38016 29640 38068 29646
rect 38016 29582 38068 29588
rect 38028 29170 38056 29582
rect 38016 29164 38068 29170
rect 38016 29106 38068 29112
rect 37464 29096 37516 29102
rect 37464 29038 37516 29044
rect 37924 29096 37976 29102
rect 37924 29038 37976 29044
rect 37936 28082 37964 29038
rect 37924 28076 37976 28082
rect 37924 28018 37976 28024
rect 37096 28008 37148 28014
rect 37096 27950 37148 27956
rect 37108 27606 37136 27950
rect 37096 27600 37148 27606
rect 37096 27542 37148 27548
rect 37924 27532 37976 27538
rect 37924 27474 37976 27480
rect 37188 27464 37240 27470
rect 37188 27406 37240 27412
rect 37016 26846 37136 26874
rect 36728 26240 36780 26246
rect 36728 26182 36780 26188
rect 36544 25356 36596 25362
rect 36544 25298 36596 25304
rect 36636 25356 36688 25362
rect 36636 25298 36688 25304
rect 36912 25220 36964 25226
rect 36912 25162 36964 25168
rect 36544 25152 36596 25158
rect 36464 25112 36544 25140
rect 36544 25094 36596 25100
rect 36360 24744 36412 24750
rect 36188 24704 36360 24732
rect 36084 24336 36136 24342
rect 36084 24278 36136 24284
rect 36096 23662 36124 24278
rect 36084 23656 36136 23662
rect 36084 23598 36136 23604
rect 36084 21480 36136 21486
rect 36084 21422 36136 21428
rect 36096 20398 36124 21422
rect 36084 20392 36136 20398
rect 36084 20334 36136 20340
rect 35992 19916 36044 19922
rect 35992 19858 36044 19864
rect 36084 19372 36136 19378
rect 36084 19314 36136 19320
rect 35808 19168 35860 19174
rect 35808 19110 35860 19116
rect 35900 18828 35952 18834
rect 35900 18770 35952 18776
rect 35912 18630 35940 18770
rect 35900 18624 35952 18630
rect 35900 18566 35952 18572
rect 35716 18420 35768 18426
rect 35716 18362 35768 18368
rect 35728 18170 35756 18362
rect 35636 18142 35756 18170
rect 35532 17536 35584 17542
rect 35532 17478 35584 17484
rect 35544 16250 35572 17478
rect 35636 16658 35664 18142
rect 35808 17672 35860 17678
rect 35808 17614 35860 17620
rect 35716 17536 35768 17542
rect 35716 17478 35768 17484
rect 35728 17134 35756 17478
rect 35820 17202 35848 17614
rect 35808 17196 35860 17202
rect 35808 17138 35860 17144
rect 35716 17128 35768 17134
rect 35716 17070 35768 17076
rect 35624 16652 35676 16658
rect 35624 16594 35676 16600
rect 35532 16244 35584 16250
rect 35532 16186 35584 16192
rect 35636 16182 35664 16594
rect 35624 16176 35676 16182
rect 35624 16118 35676 16124
rect 35820 16046 35848 17138
rect 35268 15966 35388 15994
rect 35440 16040 35492 16046
rect 35440 15982 35492 15988
rect 35808 16040 35860 16046
rect 35808 15982 35860 15988
rect 34940 15260 35236 15280
rect 34996 15258 35020 15260
rect 35076 15258 35100 15260
rect 35156 15258 35180 15260
rect 35018 15206 35020 15258
rect 35082 15206 35094 15258
rect 35156 15206 35158 15258
rect 34996 15204 35020 15206
rect 35076 15204 35100 15206
rect 35156 15204 35180 15206
rect 34940 15184 35236 15204
rect 35268 14958 35296 15966
rect 35348 15360 35400 15366
rect 35348 15302 35400 15308
rect 35256 14952 35308 14958
rect 35256 14894 35308 14900
rect 34796 14476 34848 14482
rect 34796 14418 34848 14424
rect 34808 13802 34836 14418
rect 34940 14172 35236 14192
rect 34996 14170 35020 14172
rect 35076 14170 35100 14172
rect 35156 14170 35180 14172
rect 35018 14118 35020 14170
rect 35082 14118 35094 14170
rect 35156 14118 35158 14170
rect 34996 14116 35020 14118
rect 35076 14116 35100 14118
rect 35156 14116 35180 14118
rect 34940 14096 35236 14116
rect 34796 13796 34848 13802
rect 34796 13738 34848 13744
rect 34888 13388 34940 13394
rect 34808 13348 34888 13376
rect 34808 12850 34836 13348
rect 34888 13330 34940 13336
rect 35256 13320 35308 13326
rect 35256 13262 35308 13268
rect 34940 13084 35236 13104
rect 34996 13082 35020 13084
rect 35076 13082 35100 13084
rect 35156 13082 35180 13084
rect 35018 13030 35020 13082
rect 35082 13030 35094 13082
rect 35156 13030 35158 13082
rect 34996 13028 35020 13030
rect 35076 13028 35100 13030
rect 35156 13028 35180 13030
rect 34940 13008 35236 13028
rect 34796 12844 34848 12850
rect 34796 12786 34848 12792
rect 35268 12782 35296 13262
rect 35256 12776 35308 12782
rect 34794 12744 34850 12753
rect 35256 12718 35308 12724
rect 34794 12679 34850 12688
rect 34808 12238 34836 12679
rect 34624 12158 34744 12186
rect 34796 12232 34848 12238
rect 34796 12174 34848 12180
rect 34520 12096 34572 12102
rect 34520 12038 34572 12044
rect 34428 11824 34480 11830
rect 34428 11766 34480 11772
rect 34336 10464 34388 10470
rect 34336 10406 34388 10412
rect 34348 9654 34376 10406
rect 34336 9648 34388 9654
rect 34336 9590 34388 9596
rect 34164 9472 34284 9500
rect 34060 9454 34112 9460
rect 34072 8634 34100 9454
rect 34256 9110 34284 9472
rect 34244 9104 34296 9110
rect 34244 9046 34296 9052
rect 34060 8628 34112 8634
rect 34060 8570 34112 8576
rect 33784 8424 33836 8430
rect 33784 8366 33836 8372
rect 33876 8424 33928 8430
rect 33876 8366 33928 8372
rect 33888 8090 33916 8366
rect 34256 8362 34284 9046
rect 34348 8974 34376 9590
rect 34336 8968 34388 8974
rect 34336 8910 34388 8916
rect 34440 8838 34468 11766
rect 34532 11218 34560 12038
rect 34520 11212 34572 11218
rect 34520 11154 34572 11160
rect 34520 9580 34572 9586
rect 34520 9522 34572 9528
rect 34428 8832 34480 8838
rect 34428 8774 34480 8780
rect 34336 8424 34388 8430
rect 34336 8366 34388 8372
rect 34244 8356 34296 8362
rect 34244 8298 34296 8304
rect 33876 8084 33928 8090
rect 33876 8026 33928 8032
rect 34348 8022 34376 8366
rect 34440 8022 34468 8774
rect 34532 8430 34560 9522
rect 34520 8424 34572 8430
rect 34520 8366 34572 8372
rect 34336 8016 34388 8022
rect 34336 7958 34388 7964
rect 34428 8016 34480 8022
rect 34428 7958 34480 7964
rect 33508 7948 33560 7954
rect 33508 7890 33560 7896
rect 33416 7540 33468 7546
rect 33416 7482 33468 7488
rect 33324 7336 33376 7342
rect 33324 7278 33376 7284
rect 32772 7268 32824 7274
rect 32772 7210 32824 7216
rect 32680 7200 32732 7206
rect 32680 7142 32732 7148
rect 32404 6316 32456 6322
rect 32404 6258 32456 6264
rect 31944 6248 31996 6254
rect 31944 6190 31996 6196
rect 31760 6180 31812 6186
rect 31760 6122 31812 6128
rect 31024 5908 31076 5914
rect 31024 5850 31076 5856
rect 31036 4622 31064 5850
rect 31772 5778 31800 6122
rect 32692 5778 32720 7142
rect 32784 6322 32812 7210
rect 33416 6792 33468 6798
rect 33520 6746 33548 7890
rect 33692 7880 33744 7886
rect 33692 7822 33744 7828
rect 33600 7200 33652 7206
rect 33600 7142 33652 7148
rect 33612 6798 33640 7142
rect 33704 6866 33732 7822
rect 33692 6860 33744 6866
rect 33692 6802 33744 6808
rect 33468 6740 33548 6746
rect 33416 6734 33548 6740
rect 33600 6792 33652 6798
rect 33600 6734 33652 6740
rect 34428 6792 34480 6798
rect 34428 6734 34480 6740
rect 33428 6718 33548 6734
rect 32772 6316 32824 6322
rect 32772 6258 32824 6264
rect 33520 6118 33548 6718
rect 33612 6254 33640 6734
rect 33600 6248 33652 6254
rect 33600 6190 33652 6196
rect 33508 6112 33560 6118
rect 33508 6054 33560 6060
rect 31760 5772 31812 5778
rect 31760 5714 31812 5720
rect 32680 5772 32732 5778
rect 32680 5714 32732 5720
rect 33232 5772 33284 5778
rect 33232 5714 33284 5720
rect 31392 4684 31444 4690
rect 31392 4626 31444 4632
rect 31024 4616 31076 4622
rect 31024 4558 31076 4564
rect 30932 4140 30984 4146
rect 30932 4082 30984 4088
rect 31404 3738 31432 4626
rect 31772 4622 31800 5714
rect 32588 5704 32640 5710
rect 32588 5646 32640 5652
rect 32128 5160 32180 5166
rect 32128 5102 32180 5108
rect 32140 4758 32168 5102
rect 32128 4752 32180 4758
rect 32128 4694 32180 4700
rect 32600 4690 32628 5646
rect 33244 5370 33272 5714
rect 33232 5364 33284 5370
rect 33232 5306 33284 5312
rect 32588 4684 32640 4690
rect 32588 4626 32640 4632
rect 31760 4616 31812 4622
rect 31760 4558 31812 4564
rect 31772 4078 31800 4558
rect 32784 4146 33088 4162
rect 31944 4140 31996 4146
rect 31944 4082 31996 4088
rect 32772 4140 33100 4146
rect 32824 4134 33048 4140
rect 32772 4082 32824 4088
rect 33048 4082 33100 4088
rect 31760 4072 31812 4078
rect 31760 4014 31812 4020
rect 31852 4004 31904 4010
rect 31852 3946 31904 3952
rect 30104 3732 30156 3738
rect 30104 3674 30156 3680
rect 30288 3732 30340 3738
rect 30288 3674 30340 3680
rect 30656 3732 30708 3738
rect 30656 3674 30708 3680
rect 31392 3732 31444 3738
rect 31392 3674 31444 3680
rect 29552 3528 29604 3534
rect 29472 3488 29552 3516
rect 28264 3392 28316 3398
rect 28264 3334 28316 3340
rect 27712 3188 27764 3194
rect 27712 3130 27764 3136
rect 27804 3188 27856 3194
rect 27804 3130 27856 3136
rect 28724 3188 28776 3194
rect 28724 3130 28776 3136
rect 27724 2990 27752 3130
rect 27068 2984 27120 2990
rect 27068 2926 27120 2932
rect 27712 2984 27764 2990
rect 27712 2926 27764 2932
rect 27988 2848 28040 2854
rect 27988 2790 28040 2796
rect 26884 2508 26936 2514
rect 26884 2450 26936 2456
rect 26700 2440 26752 2446
rect 26700 2382 26752 2388
rect 25596 2304 25648 2310
rect 25596 2246 25648 2252
rect 25608 2038 25636 2246
rect 25596 2032 25648 2038
rect 25596 1974 25648 1980
rect 25780 1964 25832 1970
rect 25780 1906 25832 1912
rect 25792 800 25820 1906
rect 28000 800 28028 2790
rect 28736 2378 28764 3130
rect 29104 2990 29132 3470
rect 29092 2984 29144 2990
rect 29092 2926 29144 2932
rect 29472 2582 29500 3488
rect 29552 3470 29604 3476
rect 30116 2922 30144 3674
rect 30564 3528 30616 3534
rect 30564 3470 30616 3476
rect 30576 3398 30604 3470
rect 30668 3398 30696 3674
rect 30564 3392 30616 3398
rect 30564 3334 30616 3340
rect 30656 3392 30708 3398
rect 30656 3334 30708 3340
rect 30104 2916 30156 2922
rect 30104 2858 30156 2864
rect 30288 2848 30340 2854
rect 30288 2790 30340 2796
rect 30300 2650 30328 2790
rect 30288 2644 30340 2650
rect 30288 2586 30340 2592
rect 29460 2576 29512 2582
rect 29460 2518 29512 2524
rect 30576 2514 30604 3334
rect 31404 3194 31432 3674
rect 31864 3602 31892 3946
rect 31956 3670 31984 4082
rect 32128 4072 32180 4078
rect 32128 4014 32180 4020
rect 32864 4072 32916 4078
rect 32864 4014 32916 4020
rect 32036 4004 32088 4010
rect 32036 3946 32088 3952
rect 31944 3664 31996 3670
rect 31944 3606 31996 3612
rect 31852 3596 31904 3602
rect 31852 3538 31904 3544
rect 31392 3188 31444 3194
rect 31392 3130 31444 3136
rect 31404 2514 31432 3130
rect 32048 2990 32076 3946
rect 32140 3670 32168 4014
rect 32876 3738 32904 4014
rect 32864 3732 32916 3738
rect 32864 3674 32916 3680
rect 32128 3664 32180 3670
rect 32128 3606 32180 3612
rect 33416 3596 33468 3602
rect 33416 3538 33468 3544
rect 32680 3528 32732 3534
rect 32732 3476 33180 3482
rect 32680 3470 33180 3476
rect 32692 3454 33180 3470
rect 33152 2990 33180 3454
rect 33428 3398 33456 3538
rect 33520 3534 33548 6054
rect 33612 5778 33640 6190
rect 34440 6118 34468 6734
rect 34624 6458 34652 12158
rect 35360 12102 35388 15302
rect 35716 14952 35768 14958
rect 35716 14894 35768 14900
rect 35440 14272 35492 14278
rect 35440 14214 35492 14220
rect 35532 14272 35584 14278
rect 35532 14214 35584 14220
rect 35452 13938 35480 14214
rect 35544 14074 35572 14214
rect 35532 14068 35584 14074
rect 35532 14010 35584 14016
rect 35440 13932 35492 13938
rect 35440 13874 35492 13880
rect 35624 13864 35676 13870
rect 35624 13806 35676 13812
rect 35440 13388 35492 13394
rect 35440 13330 35492 13336
rect 35452 12782 35480 13330
rect 35636 13190 35664 13806
rect 35728 13297 35756 14894
rect 35714 13288 35770 13297
rect 35714 13223 35770 13232
rect 35624 13184 35676 13190
rect 35624 13126 35676 13132
rect 35440 12776 35492 12782
rect 35440 12718 35492 12724
rect 35348 12096 35400 12102
rect 35348 12038 35400 12044
rect 34940 11996 35236 12016
rect 34996 11994 35020 11996
rect 35076 11994 35100 11996
rect 35156 11994 35180 11996
rect 35018 11942 35020 11994
rect 35082 11942 35094 11994
rect 35156 11942 35158 11994
rect 34996 11940 35020 11942
rect 35076 11940 35100 11942
rect 35156 11940 35180 11942
rect 34940 11920 35236 11940
rect 35360 11694 35388 12038
rect 35348 11688 35400 11694
rect 35348 11630 35400 11636
rect 35532 11688 35584 11694
rect 35532 11630 35584 11636
rect 35808 11688 35860 11694
rect 35808 11630 35860 11636
rect 35544 11354 35572 11630
rect 35532 11348 35584 11354
rect 35532 11290 35584 11296
rect 35820 11286 35848 11630
rect 35912 11354 35940 18566
rect 36096 18290 36124 19314
rect 36084 18284 36136 18290
rect 36084 18226 36136 18232
rect 35992 18216 36044 18222
rect 35992 18158 36044 18164
rect 36004 16794 36032 18158
rect 36096 17134 36124 18226
rect 36084 17128 36136 17134
rect 36084 17070 36136 17076
rect 35992 16788 36044 16794
rect 35992 16730 36044 16736
rect 36084 16584 36136 16590
rect 36084 16526 36136 16532
rect 36096 16114 36124 16526
rect 36084 16108 36136 16114
rect 36084 16050 36136 16056
rect 36188 15858 36216 24704
rect 36360 24686 36412 24692
rect 36360 24608 36412 24614
rect 36360 24550 36412 24556
rect 36372 24070 36400 24550
rect 36360 24064 36412 24070
rect 36360 24006 36412 24012
rect 36268 23656 36320 23662
rect 36266 23624 36268 23633
rect 36320 23624 36322 23633
rect 36266 23559 36322 23568
rect 36268 22772 36320 22778
rect 36268 22714 36320 22720
rect 36280 20398 36308 22714
rect 36372 22642 36400 24006
rect 36452 23180 36504 23186
rect 36452 23122 36504 23128
rect 36360 22636 36412 22642
rect 36360 22578 36412 22584
rect 36372 21486 36400 22578
rect 36464 22438 36492 23122
rect 36452 22432 36504 22438
rect 36452 22374 36504 22380
rect 36452 21888 36504 21894
rect 36452 21830 36504 21836
rect 36360 21480 36412 21486
rect 36360 21422 36412 21428
rect 36464 21146 36492 21830
rect 36452 21140 36504 21146
rect 36452 21082 36504 21088
rect 36268 20392 36320 20398
rect 36268 20334 36320 20340
rect 36280 19310 36308 20334
rect 36268 19304 36320 19310
rect 36268 19246 36320 19252
rect 36452 17808 36504 17814
rect 36452 17750 36504 17756
rect 36360 17740 36412 17746
rect 36360 17682 36412 17688
rect 36268 17536 36320 17542
rect 36268 17478 36320 17484
rect 36280 16658 36308 17478
rect 36372 17202 36400 17682
rect 36360 17196 36412 17202
rect 36360 17138 36412 17144
rect 36464 17082 36492 17750
rect 36556 17728 36584 25094
rect 36728 24608 36780 24614
rect 36728 24550 36780 24556
rect 36740 23662 36768 24550
rect 36728 23656 36780 23662
rect 36728 23598 36780 23604
rect 36820 23112 36872 23118
rect 36820 23054 36872 23060
rect 36832 21962 36860 23054
rect 36820 21956 36872 21962
rect 36820 21898 36872 21904
rect 36924 21842 36952 25162
rect 37004 24812 37056 24818
rect 37004 24754 37056 24760
rect 37016 24274 37044 24754
rect 37004 24268 37056 24274
rect 37004 24210 37056 24216
rect 37016 23730 37044 24210
rect 37004 23724 37056 23730
rect 37004 23666 37056 23672
rect 37004 22160 37056 22166
rect 37004 22102 37056 22108
rect 36832 21814 36952 21842
rect 36636 21548 36688 21554
rect 36636 21490 36688 21496
rect 36648 18426 36676 21490
rect 36726 19952 36782 19961
rect 36726 19887 36782 19896
rect 36636 18420 36688 18426
rect 36636 18362 36688 18368
rect 36556 17700 36676 17728
rect 36544 17604 36596 17610
rect 36544 17546 36596 17552
rect 36372 17054 36492 17082
rect 36268 16652 36320 16658
rect 36268 16594 36320 16600
rect 36372 16454 36400 17054
rect 36452 16992 36504 16998
rect 36452 16934 36504 16940
rect 36360 16448 36412 16454
rect 36360 16390 36412 16396
rect 36372 16130 36400 16390
rect 36004 15830 36216 15858
rect 36280 16102 36400 16130
rect 36004 12764 36032 15830
rect 36280 15638 36308 16102
rect 36360 16040 36412 16046
rect 36360 15982 36412 15988
rect 36268 15632 36320 15638
rect 36268 15574 36320 15580
rect 36176 15564 36228 15570
rect 36176 15506 36228 15512
rect 36188 15026 36216 15506
rect 36176 15020 36228 15026
rect 36176 14962 36228 14968
rect 36176 14476 36228 14482
rect 36176 14418 36228 14424
rect 36084 13864 36136 13870
rect 36084 13806 36136 13812
rect 36096 13258 36124 13806
rect 36188 13530 36216 14418
rect 36176 13524 36228 13530
rect 36176 13466 36228 13472
rect 36176 13320 36228 13326
rect 36176 13262 36228 13268
rect 36084 13252 36136 13258
rect 36084 13194 36136 13200
rect 36188 12889 36216 13262
rect 36174 12880 36230 12889
rect 36280 12866 36308 15574
rect 36372 14958 36400 15982
rect 36464 15570 36492 16934
rect 36556 16658 36584 17546
rect 36544 16652 36596 16658
rect 36544 16594 36596 16600
rect 36648 16522 36676 17700
rect 36636 16516 36688 16522
rect 36636 16458 36688 16464
rect 36544 15972 36596 15978
rect 36544 15914 36596 15920
rect 36556 15570 36584 15914
rect 36452 15564 36504 15570
rect 36452 15506 36504 15512
rect 36544 15564 36596 15570
rect 36544 15506 36596 15512
rect 36360 14952 36412 14958
rect 36360 14894 36412 14900
rect 36464 14940 36492 15506
rect 36648 15026 36676 16458
rect 36636 15020 36688 15026
rect 36636 14962 36688 14968
rect 36544 14952 36596 14958
rect 36464 14912 36544 14940
rect 36372 12986 36400 14894
rect 36360 12980 36412 12986
rect 36360 12922 36412 12928
rect 36280 12838 36400 12866
rect 36174 12815 36230 12824
rect 36004 12736 36308 12764
rect 36084 12300 36136 12306
rect 36084 12242 36136 12248
rect 35992 12232 36044 12238
rect 35992 12174 36044 12180
rect 36004 11694 36032 12174
rect 35992 11688 36044 11694
rect 35992 11630 36044 11636
rect 35900 11348 35952 11354
rect 35900 11290 35952 11296
rect 35808 11280 35860 11286
rect 35808 11222 35860 11228
rect 36004 11218 36032 11630
rect 34796 11212 34848 11218
rect 34796 11154 34848 11160
rect 35992 11212 36044 11218
rect 35992 11154 36044 11160
rect 34808 10470 34836 11154
rect 35438 11112 35494 11121
rect 35438 11047 35494 11056
rect 34940 10908 35236 10928
rect 34996 10906 35020 10908
rect 35076 10906 35100 10908
rect 35156 10906 35180 10908
rect 35018 10854 35020 10906
rect 35082 10854 35094 10906
rect 35156 10854 35158 10906
rect 34996 10852 35020 10854
rect 35076 10852 35100 10854
rect 35156 10852 35180 10854
rect 34940 10832 35236 10852
rect 34796 10464 34848 10470
rect 34796 10406 34848 10412
rect 34940 9820 35236 9840
rect 34996 9818 35020 9820
rect 35076 9818 35100 9820
rect 35156 9818 35180 9820
rect 35018 9766 35020 9818
rect 35082 9766 35094 9818
rect 35156 9766 35158 9818
rect 34996 9764 35020 9766
rect 35076 9764 35100 9766
rect 35156 9764 35180 9766
rect 34940 9744 35236 9764
rect 35072 9512 35124 9518
rect 35072 9454 35124 9460
rect 35084 9110 35112 9454
rect 35256 9376 35308 9382
rect 35256 9318 35308 9324
rect 35072 9104 35124 9110
rect 35072 9046 35124 9052
rect 35268 9042 35296 9318
rect 35256 9036 35308 9042
rect 35256 8978 35308 8984
rect 34940 8732 35236 8752
rect 34996 8730 35020 8732
rect 35076 8730 35100 8732
rect 35156 8730 35180 8732
rect 35018 8678 35020 8730
rect 35082 8678 35094 8730
rect 35156 8678 35158 8730
rect 34996 8676 35020 8678
rect 35076 8676 35100 8678
rect 35156 8676 35180 8678
rect 34940 8656 35236 8676
rect 35348 7948 35400 7954
rect 35348 7890 35400 7896
rect 34796 7880 34848 7886
rect 34796 7822 34848 7828
rect 34704 6656 34756 6662
rect 34704 6598 34756 6604
rect 34612 6452 34664 6458
rect 34612 6394 34664 6400
rect 34428 6112 34480 6118
rect 34428 6054 34480 6060
rect 34716 5778 34744 6598
rect 34808 5846 34836 7822
rect 34940 7644 35236 7664
rect 34996 7642 35020 7644
rect 35076 7642 35100 7644
rect 35156 7642 35180 7644
rect 35018 7590 35020 7642
rect 35082 7590 35094 7642
rect 35156 7590 35158 7642
rect 34996 7588 35020 7590
rect 35076 7588 35100 7590
rect 35156 7588 35180 7590
rect 34940 7568 35236 7588
rect 35072 7336 35124 7342
rect 35072 7278 35124 7284
rect 35084 7002 35112 7278
rect 35072 6996 35124 7002
rect 35072 6938 35124 6944
rect 34940 6556 35236 6576
rect 34996 6554 35020 6556
rect 35076 6554 35100 6556
rect 35156 6554 35180 6556
rect 35018 6502 35020 6554
rect 35082 6502 35094 6554
rect 35156 6502 35158 6554
rect 34996 6500 35020 6502
rect 35076 6500 35100 6502
rect 35156 6500 35180 6502
rect 34940 6480 35236 6500
rect 34888 6384 34940 6390
rect 34888 6326 34940 6332
rect 34796 5840 34848 5846
rect 34796 5782 34848 5788
rect 34900 5778 34928 6326
rect 35360 5914 35388 7890
rect 35452 7410 35480 11047
rect 35900 11008 35952 11014
rect 35900 10950 35952 10956
rect 35624 10668 35676 10674
rect 35624 10610 35676 10616
rect 35636 10130 35664 10610
rect 35912 10441 35940 10950
rect 36096 10538 36124 12242
rect 36176 11552 36228 11558
rect 36176 11494 36228 11500
rect 36188 11286 36216 11494
rect 36176 11280 36228 11286
rect 36176 11222 36228 11228
rect 36084 10532 36136 10538
rect 36084 10474 36136 10480
rect 35898 10432 35954 10441
rect 35898 10367 35954 10376
rect 35624 10124 35676 10130
rect 35624 10066 35676 10072
rect 35808 10124 35860 10130
rect 35808 10066 35860 10072
rect 35820 9994 35848 10066
rect 35808 9988 35860 9994
rect 35808 9930 35860 9936
rect 35716 9716 35768 9722
rect 35716 9658 35768 9664
rect 35728 9518 35756 9658
rect 35820 9586 35848 9930
rect 35808 9580 35860 9586
rect 35808 9522 35860 9528
rect 35716 9512 35768 9518
rect 35716 9454 35768 9460
rect 36084 7880 36136 7886
rect 36084 7822 36136 7828
rect 35440 7404 35492 7410
rect 35440 7346 35492 7352
rect 36096 6322 36124 7822
rect 36280 7750 36308 12736
rect 36372 11014 36400 12838
rect 36464 12238 36492 14912
rect 36544 14894 36596 14900
rect 36544 13796 36596 13802
rect 36544 13738 36596 13744
rect 36556 13462 36584 13738
rect 36544 13456 36596 13462
rect 36544 13398 36596 13404
rect 36648 12850 36676 14962
rect 36636 12844 36688 12850
rect 36636 12786 36688 12792
rect 36740 12730 36768 19887
rect 36832 12866 36860 21814
rect 37016 20380 37044 22102
rect 36924 20352 37044 20380
rect 36924 18902 36952 20352
rect 37004 19712 37056 19718
rect 37004 19654 37056 19660
rect 36912 18896 36964 18902
rect 36912 18838 36964 18844
rect 37016 16697 37044 19654
rect 37002 16688 37058 16697
rect 37002 16623 37058 16632
rect 36912 14408 36964 14414
rect 36912 14350 36964 14356
rect 36924 12986 36952 14350
rect 37002 13696 37058 13705
rect 37002 13631 37058 13640
rect 36912 12980 36964 12986
rect 36912 12922 36964 12928
rect 36832 12838 36952 12866
rect 36648 12702 36768 12730
rect 36452 12232 36504 12238
rect 36452 12174 36504 12180
rect 36452 11212 36504 11218
rect 36452 11154 36504 11160
rect 36360 11008 36412 11014
rect 36360 10950 36412 10956
rect 36372 10674 36400 10950
rect 36360 10668 36412 10674
rect 36360 10610 36412 10616
rect 36360 10532 36412 10538
rect 36360 10474 36412 10480
rect 36372 9178 36400 10474
rect 36464 10062 36492 11154
rect 36452 10056 36504 10062
rect 36452 9998 36504 10004
rect 36360 9172 36412 9178
rect 36360 9114 36412 9120
rect 36268 7744 36320 7750
rect 36268 7686 36320 7692
rect 36084 6316 36136 6322
rect 36084 6258 36136 6264
rect 35348 5908 35400 5914
rect 35348 5850 35400 5856
rect 33600 5772 33652 5778
rect 33600 5714 33652 5720
rect 34520 5772 34572 5778
rect 34520 5714 34572 5720
rect 34704 5772 34756 5778
rect 34704 5714 34756 5720
rect 34888 5772 34940 5778
rect 34888 5714 34940 5720
rect 35624 5772 35676 5778
rect 35624 5714 35676 5720
rect 33692 5704 33744 5710
rect 33692 5646 33744 5652
rect 33600 4616 33652 4622
rect 33600 4558 33652 4564
rect 33508 3528 33560 3534
rect 33508 3470 33560 3476
rect 33416 3392 33468 3398
rect 33416 3334 33468 3340
rect 32036 2984 32088 2990
rect 32036 2926 32088 2932
rect 33140 2984 33192 2990
rect 33140 2926 33192 2932
rect 32036 2848 32088 2854
rect 32036 2790 32088 2796
rect 30012 2508 30064 2514
rect 30012 2450 30064 2456
rect 30564 2508 30616 2514
rect 30564 2450 30616 2456
rect 31392 2508 31444 2514
rect 31392 2450 31444 2456
rect 28724 2372 28776 2378
rect 28724 2314 28776 2320
rect 30024 800 30052 2450
rect 32048 1170 32076 2790
rect 33152 2446 33180 2926
rect 33428 2514 33456 3334
rect 33520 2854 33548 3470
rect 33612 3058 33640 4558
rect 33704 3602 33732 5646
rect 34532 5166 34560 5714
rect 34612 5704 34664 5710
rect 34612 5646 34664 5652
rect 34520 5160 34572 5166
rect 34520 5102 34572 5108
rect 34428 5024 34480 5030
rect 34428 4966 34480 4972
rect 34440 4690 34468 4966
rect 34336 4684 34388 4690
rect 34336 4626 34388 4632
rect 34428 4684 34480 4690
rect 34428 4626 34480 4632
rect 33968 4208 34020 4214
rect 33968 4150 34020 4156
rect 33980 4078 34008 4150
rect 33876 4072 33928 4078
rect 33876 4014 33928 4020
rect 33968 4072 34020 4078
rect 33968 4014 34020 4020
rect 34348 4026 34376 4626
rect 34440 4214 34468 4626
rect 34520 4616 34572 4622
rect 34520 4558 34572 4564
rect 34428 4208 34480 4214
rect 34428 4150 34480 4156
rect 34428 4072 34480 4078
rect 34348 4020 34428 4026
rect 34348 4014 34480 4020
rect 33692 3596 33744 3602
rect 33692 3538 33744 3544
rect 33600 3052 33652 3058
rect 33600 2994 33652 3000
rect 33508 2848 33560 2854
rect 33508 2790 33560 2796
rect 33888 2582 33916 4014
rect 33980 3194 34008 4014
rect 34348 3998 34468 4014
rect 34348 3738 34376 3998
rect 34336 3732 34388 3738
rect 34336 3674 34388 3680
rect 33968 3188 34020 3194
rect 33968 3130 34020 3136
rect 34532 3058 34560 4558
rect 34624 4146 34652 5646
rect 34940 5468 35236 5488
rect 34996 5466 35020 5468
rect 35076 5466 35100 5468
rect 35156 5466 35180 5468
rect 35018 5414 35020 5466
rect 35082 5414 35094 5466
rect 35156 5414 35158 5466
rect 34996 5412 35020 5414
rect 35076 5412 35100 5414
rect 35156 5412 35180 5414
rect 34940 5392 35236 5412
rect 35636 5166 35664 5714
rect 36096 5166 36124 6258
rect 36544 5772 36596 5778
rect 36544 5714 36596 5720
rect 36556 5166 36584 5714
rect 35624 5160 35676 5166
rect 35624 5102 35676 5108
rect 36084 5160 36136 5166
rect 36084 5102 36136 5108
rect 36544 5160 36596 5166
rect 36544 5102 36596 5108
rect 35992 5092 36044 5098
rect 35992 5034 36044 5040
rect 35348 4616 35400 4622
rect 35348 4558 35400 4564
rect 34940 4380 35236 4400
rect 34996 4378 35020 4380
rect 35076 4378 35100 4380
rect 35156 4378 35180 4380
rect 35018 4326 35020 4378
rect 35082 4326 35094 4378
rect 35156 4326 35158 4378
rect 34996 4324 35020 4326
rect 35076 4324 35100 4326
rect 35156 4324 35180 4326
rect 34940 4304 35236 4324
rect 34612 4140 34664 4146
rect 34612 4082 34664 4088
rect 35360 3942 35388 4558
rect 35900 4276 35952 4282
rect 35900 4218 35952 4224
rect 35912 4185 35940 4218
rect 35898 4176 35954 4185
rect 36004 4146 36032 5034
rect 36648 4826 36676 12702
rect 36820 11688 36872 11694
rect 36820 11630 36872 11636
rect 36726 10704 36782 10713
rect 36726 10639 36782 10648
rect 36740 10606 36768 10639
rect 36728 10600 36780 10606
rect 36728 10542 36780 10548
rect 36832 8362 36860 11630
rect 36820 8356 36872 8362
rect 36820 8298 36872 8304
rect 36726 7440 36782 7449
rect 36726 7375 36728 7384
rect 36780 7375 36782 7384
rect 36728 7346 36780 7352
rect 36924 6866 36952 12838
rect 37016 12782 37044 13631
rect 37004 12776 37056 12782
rect 37004 12718 37056 12724
rect 36912 6860 36964 6866
rect 36912 6802 36964 6808
rect 36912 6656 36964 6662
rect 36912 6598 36964 6604
rect 36728 6180 36780 6186
rect 36728 6122 36780 6128
rect 36740 5914 36768 6122
rect 36728 5908 36780 5914
rect 36728 5850 36780 5856
rect 36740 5370 36768 5850
rect 36924 5778 36952 6598
rect 37108 6390 37136 26846
rect 37200 22778 37228 27406
rect 37832 27328 37884 27334
rect 37832 27270 37884 27276
rect 37464 26920 37516 26926
rect 37464 26862 37516 26868
rect 37476 25906 37504 26862
rect 37648 26580 37700 26586
rect 37648 26522 37700 26528
rect 37464 25900 37516 25906
rect 37464 25842 37516 25848
rect 37476 24818 37504 25842
rect 37464 24812 37516 24818
rect 37464 24754 37516 24760
rect 37372 24744 37424 24750
rect 37372 24686 37424 24692
rect 37280 24404 37332 24410
rect 37280 24346 37332 24352
rect 37292 23730 37320 24346
rect 37384 23866 37412 24686
rect 37372 23860 37424 23866
rect 37372 23802 37424 23808
rect 37280 23724 37332 23730
rect 37280 23666 37332 23672
rect 37188 22772 37240 22778
rect 37188 22714 37240 22720
rect 37476 22642 37504 24754
rect 37464 22636 37516 22642
rect 37464 22578 37516 22584
rect 37556 21956 37608 21962
rect 37556 21898 37608 21904
rect 37568 21554 37596 21898
rect 37556 21548 37608 21554
rect 37556 21490 37608 21496
rect 37280 21480 37332 21486
rect 37280 21422 37332 21428
rect 37188 20868 37240 20874
rect 37188 20810 37240 20816
rect 37200 19310 37228 20810
rect 37292 20398 37320 21422
rect 37280 20392 37332 20398
rect 37280 20334 37332 20340
rect 37292 19378 37320 20334
rect 37280 19372 37332 19378
rect 37280 19314 37332 19320
rect 37188 19304 37240 19310
rect 37188 19246 37240 19252
rect 37556 17536 37608 17542
rect 37556 17478 37608 17484
rect 37188 17196 37240 17202
rect 37188 17138 37240 17144
rect 37200 16114 37228 17138
rect 37568 16590 37596 17478
rect 37556 16584 37608 16590
rect 37556 16526 37608 16532
rect 37188 16108 37240 16114
rect 37188 16050 37240 16056
rect 37568 13870 37596 16526
rect 37372 13864 37424 13870
rect 37372 13806 37424 13812
rect 37556 13864 37608 13870
rect 37556 13806 37608 13812
rect 37280 13796 37332 13802
rect 37280 13738 37332 13744
rect 37188 13320 37240 13326
rect 37188 13262 37240 13268
rect 37200 12850 37228 13262
rect 37188 12844 37240 12850
rect 37188 12786 37240 12792
rect 37292 12374 37320 13738
rect 37384 13530 37412 13806
rect 37372 13524 37424 13530
rect 37372 13466 37424 13472
rect 37384 13394 37412 13466
rect 37568 13462 37596 13806
rect 37556 13456 37608 13462
rect 37556 13398 37608 13404
rect 37372 13388 37424 13394
rect 37372 13330 37424 13336
rect 37280 12368 37332 12374
rect 37280 12310 37332 12316
rect 37384 11778 37412 13330
rect 37292 11750 37412 11778
rect 37186 11656 37242 11665
rect 37186 11591 37188 11600
rect 37240 11591 37242 11600
rect 37188 11562 37240 11568
rect 37292 10742 37320 11750
rect 37372 11688 37424 11694
rect 37372 11630 37424 11636
rect 37280 10736 37332 10742
rect 37280 10678 37332 10684
rect 37292 10266 37320 10678
rect 37384 10266 37412 11630
rect 37464 10600 37516 10606
rect 37464 10542 37516 10548
rect 37280 10260 37332 10266
rect 37280 10202 37332 10208
rect 37372 10260 37424 10266
rect 37372 10202 37424 10208
rect 37476 9602 37504 10542
rect 37556 10532 37608 10538
rect 37556 10474 37608 10480
rect 37384 9586 37504 9602
rect 37372 9580 37504 9586
rect 37424 9574 37504 9580
rect 37372 9522 37424 9528
rect 37188 9512 37240 9518
rect 37188 9454 37240 9460
rect 37200 9178 37228 9454
rect 37188 9172 37240 9178
rect 37188 9114 37240 9120
rect 37384 7410 37412 9522
rect 37568 9042 37596 10474
rect 37556 9036 37608 9042
rect 37556 8978 37608 8984
rect 37660 7410 37688 26522
rect 37844 25906 37872 27270
rect 37832 25900 37884 25906
rect 37832 25842 37884 25848
rect 37936 24614 37964 27474
rect 38028 26450 38056 29106
rect 38016 26444 38068 26450
rect 38016 26386 38068 26392
rect 38212 25430 38240 32710
rect 38660 32360 38712 32366
rect 38660 32302 38712 32308
rect 38672 31142 38700 32302
rect 38752 32224 38804 32230
rect 38752 32166 38804 32172
rect 38660 31136 38712 31142
rect 38660 31078 38712 31084
rect 38476 29844 38528 29850
rect 38476 29786 38528 29792
rect 38488 28626 38516 29786
rect 38672 29102 38700 31078
rect 38764 30190 38792 32166
rect 38936 31680 38988 31686
rect 38936 31622 38988 31628
rect 38844 30728 38896 30734
rect 38844 30670 38896 30676
rect 38856 30258 38884 30670
rect 38844 30252 38896 30258
rect 38844 30194 38896 30200
rect 38752 30184 38804 30190
rect 38752 30126 38804 30132
rect 38752 29572 38804 29578
rect 38752 29514 38804 29520
rect 38660 29096 38712 29102
rect 38660 29038 38712 29044
rect 38292 28620 38344 28626
rect 38292 28562 38344 28568
rect 38476 28620 38528 28626
rect 38476 28562 38528 28568
rect 38304 28150 38332 28562
rect 38292 28144 38344 28150
rect 38292 28086 38344 28092
rect 38488 28014 38516 28562
rect 38764 28014 38792 29514
rect 38948 29209 38976 31622
rect 39028 29504 39080 29510
rect 39028 29446 39080 29452
rect 38934 29200 38990 29209
rect 38934 29135 38990 29144
rect 38844 28620 38896 28626
rect 38844 28562 38896 28568
rect 38856 28082 38884 28562
rect 38844 28076 38896 28082
rect 38844 28018 38896 28024
rect 38476 28008 38528 28014
rect 38476 27950 38528 27956
rect 38752 28008 38804 28014
rect 38752 27950 38804 27956
rect 38764 27010 38792 27950
rect 38856 27130 38884 28018
rect 38844 27124 38896 27130
rect 38844 27066 38896 27072
rect 38764 26982 38884 27010
rect 38200 25424 38252 25430
rect 38200 25366 38252 25372
rect 37924 24608 37976 24614
rect 37924 24550 37976 24556
rect 38212 24342 38240 25366
rect 38292 25356 38344 25362
rect 38292 25298 38344 25304
rect 38304 24818 38332 25298
rect 38752 25288 38804 25294
rect 38752 25230 38804 25236
rect 38292 24812 38344 24818
rect 38292 24754 38344 24760
rect 38200 24336 38252 24342
rect 38200 24278 38252 24284
rect 38304 24274 38332 24754
rect 37832 24268 37884 24274
rect 37832 24210 37884 24216
rect 38292 24268 38344 24274
rect 38292 24210 38344 24216
rect 37844 22137 37872 24210
rect 38660 23248 38712 23254
rect 38198 23216 38254 23225
rect 38660 23190 38712 23196
rect 38198 23151 38200 23160
rect 38252 23151 38254 23160
rect 38384 23180 38436 23186
rect 38200 23122 38252 23128
rect 38384 23122 38436 23128
rect 38212 22778 38240 23122
rect 38200 22772 38252 22778
rect 38200 22714 38252 22720
rect 37830 22128 37886 22137
rect 37830 22063 37832 22072
rect 37884 22063 37886 22072
rect 37832 22034 37884 22040
rect 37844 21010 37872 22034
rect 37832 21004 37884 21010
rect 37832 20946 37884 20952
rect 37740 20868 37792 20874
rect 37740 20810 37792 20816
rect 37752 20466 37780 20810
rect 38108 20800 38160 20806
rect 38108 20742 38160 20748
rect 37740 20460 37792 20466
rect 37740 20402 37792 20408
rect 38120 20262 38148 20742
rect 38108 20256 38160 20262
rect 38108 20198 38160 20204
rect 38120 19922 38148 20198
rect 38108 19916 38160 19922
rect 38108 19858 38160 19864
rect 38396 19310 38424 23122
rect 38672 21078 38700 23190
rect 38764 22642 38792 25230
rect 38856 23118 38884 26982
rect 39040 26450 39068 29446
rect 39028 26444 39080 26450
rect 39028 26386 39080 26392
rect 39132 26042 39160 32914
rect 39120 26036 39172 26042
rect 39120 25978 39172 25984
rect 38844 23112 38896 23118
rect 38844 23054 38896 23060
rect 38752 22636 38804 22642
rect 38752 22578 38804 22584
rect 38844 22432 38896 22438
rect 38844 22374 38896 22380
rect 38856 21690 38884 22374
rect 38844 21684 38896 21690
rect 38844 21626 38896 21632
rect 38660 21072 38712 21078
rect 38660 21014 38712 21020
rect 38568 21004 38620 21010
rect 38568 20946 38620 20952
rect 38476 20936 38528 20942
rect 38476 20878 38528 20884
rect 38488 19922 38516 20878
rect 38476 19916 38528 19922
rect 38476 19858 38528 19864
rect 38384 19304 38436 19310
rect 38384 19246 38436 19252
rect 38396 18902 38424 19246
rect 38384 18896 38436 18902
rect 38384 18838 38436 18844
rect 38108 18828 38160 18834
rect 38108 18770 38160 18776
rect 38120 17338 38148 18770
rect 38200 18760 38252 18766
rect 38200 18702 38252 18708
rect 38212 18222 38240 18702
rect 38396 18222 38424 18838
rect 38476 18828 38528 18834
rect 38476 18770 38528 18776
rect 38200 18216 38252 18222
rect 38200 18158 38252 18164
rect 38384 18216 38436 18222
rect 38384 18158 38436 18164
rect 38108 17332 38160 17338
rect 38108 17274 38160 17280
rect 37832 17128 37884 17134
rect 37832 17070 37884 17076
rect 37844 15706 37872 17070
rect 38212 16250 38240 18158
rect 38488 18068 38516 18770
rect 38580 18290 38608 20946
rect 38672 19922 38700 21014
rect 38660 19916 38712 19922
rect 38660 19858 38712 19864
rect 38936 19168 38988 19174
rect 38936 19110 38988 19116
rect 38660 18692 38712 18698
rect 38660 18634 38712 18640
rect 38568 18284 38620 18290
rect 38568 18226 38620 18232
rect 38672 18222 38700 18634
rect 38660 18216 38712 18222
rect 38660 18158 38712 18164
rect 38568 18148 38620 18154
rect 38568 18090 38620 18096
rect 38304 18040 38516 18068
rect 38200 16244 38252 16250
rect 38200 16186 38252 16192
rect 37832 15700 37884 15706
rect 37832 15642 37884 15648
rect 37740 14952 37792 14958
rect 37740 14894 37792 14900
rect 37752 14550 37780 14894
rect 37832 14816 37884 14822
rect 37832 14758 37884 14764
rect 37740 14544 37792 14550
rect 37740 14486 37792 14492
rect 37740 14408 37792 14414
rect 37740 14350 37792 14356
rect 37752 13802 37780 14350
rect 37844 14074 37872 14758
rect 37924 14476 37976 14482
rect 37924 14418 37976 14424
rect 38016 14476 38068 14482
rect 38016 14418 38068 14424
rect 37832 14068 37884 14074
rect 37832 14010 37884 14016
rect 37844 13870 37872 14010
rect 37832 13864 37884 13870
rect 37832 13806 37884 13812
rect 37740 13796 37792 13802
rect 37740 13738 37792 13744
rect 37936 12782 37964 14418
rect 37924 12776 37976 12782
rect 37924 12718 37976 12724
rect 37832 12300 37884 12306
rect 37832 12242 37884 12248
rect 37740 12164 37792 12170
rect 37740 12106 37792 12112
rect 37752 10674 37780 12106
rect 37844 11694 37872 12242
rect 37832 11688 37884 11694
rect 37832 11630 37884 11636
rect 37936 11234 37964 12718
rect 37844 11206 37964 11234
rect 37844 11150 37872 11206
rect 37832 11144 37884 11150
rect 37832 11086 37884 11092
rect 37844 10674 37872 11086
rect 37740 10668 37792 10674
rect 37740 10610 37792 10616
rect 37832 10668 37884 10674
rect 37832 10610 37884 10616
rect 37844 8430 37872 10610
rect 38028 10130 38056 14418
rect 38108 14000 38160 14006
rect 38108 13942 38160 13948
rect 38120 13394 38148 13942
rect 38108 13388 38160 13394
rect 38108 13330 38160 13336
rect 38200 12300 38252 12306
rect 38200 12242 38252 12248
rect 38212 11286 38240 12242
rect 38200 11280 38252 11286
rect 38200 11222 38252 11228
rect 38016 10124 38068 10130
rect 38016 10066 38068 10072
rect 38028 9722 38056 10066
rect 38016 9716 38068 9722
rect 38016 9658 38068 9664
rect 38304 8634 38332 18040
rect 38580 17746 38608 18090
rect 38568 17740 38620 17746
rect 38568 17682 38620 17688
rect 38844 17672 38896 17678
rect 38844 17614 38896 17620
rect 38568 17332 38620 17338
rect 38568 17274 38620 17280
rect 38580 16658 38608 17274
rect 38660 17128 38712 17134
rect 38660 17070 38712 17076
rect 38568 16652 38620 16658
rect 38568 16594 38620 16600
rect 38568 14952 38620 14958
rect 38568 14894 38620 14900
rect 38580 14618 38608 14894
rect 38568 14612 38620 14618
rect 38568 14554 38620 14560
rect 38672 14550 38700 17070
rect 38856 16794 38884 17614
rect 38844 16788 38896 16794
rect 38844 16730 38896 16736
rect 38752 16040 38804 16046
rect 38752 15982 38804 15988
rect 38764 15162 38792 15982
rect 38752 15156 38804 15162
rect 38752 15098 38804 15104
rect 38660 14544 38712 14550
rect 38660 14486 38712 14492
rect 38568 13932 38620 13938
rect 38568 13874 38620 13880
rect 38580 13394 38608 13874
rect 38568 13388 38620 13394
rect 38568 13330 38620 13336
rect 38476 13252 38528 13258
rect 38476 13194 38528 13200
rect 38384 11620 38436 11626
rect 38384 11562 38436 11568
rect 38292 8628 38344 8634
rect 38292 8570 38344 8576
rect 38396 8430 38424 11562
rect 38488 9042 38516 13194
rect 38568 12912 38620 12918
rect 38568 12854 38620 12860
rect 38580 12306 38608 12854
rect 38856 12782 38884 16730
rect 38948 15570 38976 19110
rect 39028 18420 39080 18426
rect 39028 18362 39080 18368
rect 39040 15706 39068 18362
rect 39028 15700 39080 15706
rect 39028 15642 39080 15648
rect 38936 15564 38988 15570
rect 38936 15506 38988 15512
rect 38936 14476 38988 14482
rect 38936 14418 38988 14424
rect 38844 12776 38896 12782
rect 38844 12718 38896 12724
rect 38948 12442 38976 14418
rect 38936 12436 38988 12442
rect 38936 12378 38988 12384
rect 38568 12300 38620 12306
rect 38568 12242 38620 12248
rect 38752 12232 38804 12238
rect 38752 12174 38804 12180
rect 38568 11212 38620 11218
rect 38568 11154 38620 11160
rect 38580 10713 38608 11154
rect 38764 10810 38792 12174
rect 38948 11898 38976 12378
rect 38936 11892 38988 11898
rect 38936 11834 38988 11840
rect 38752 10804 38804 10810
rect 38752 10746 38804 10752
rect 38566 10704 38622 10713
rect 38566 10639 38622 10648
rect 38936 10464 38988 10470
rect 38936 10406 38988 10412
rect 38948 10130 38976 10406
rect 38936 10124 38988 10130
rect 38936 10066 38988 10072
rect 38476 9036 38528 9042
rect 38476 8978 38528 8984
rect 37832 8424 37884 8430
rect 37832 8366 37884 8372
rect 38384 8424 38436 8430
rect 38384 8366 38436 8372
rect 37372 7404 37424 7410
rect 37372 7346 37424 7352
rect 37648 7404 37700 7410
rect 37648 7346 37700 7352
rect 37096 6384 37148 6390
rect 37096 6326 37148 6332
rect 37096 6248 37148 6254
rect 37096 6190 37148 6196
rect 36912 5772 36964 5778
rect 36912 5714 36964 5720
rect 36728 5364 36780 5370
rect 36728 5306 36780 5312
rect 37108 5234 37136 6190
rect 37096 5228 37148 5234
rect 37096 5170 37148 5176
rect 36636 4820 36688 4826
rect 36636 4762 36688 4768
rect 35898 4111 35954 4120
rect 35992 4140 36044 4146
rect 35992 4082 36044 4088
rect 35440 4072 35492 4078
rect 35440 4014 35492 4020
rect 35348 3936 35400 3942
rect 35348 3878 35400 3884
rect 34940 3292 35236 3312
rect 34996 3290 35020 3292
rect 35076 3290 35100 3292
rect 35156 3290 35180 3292
rect 35018 3238 35020 3290
rect 35082 3238 35094 3290
rect 35156 3238 35158 3290
rect 34996 3236 35020 3238
rect 35076 3236 35100 3238
rect 35156 3236 35180 3238
rect 34940 3216 35236 3236
rect 35452 3058 35480 4014
rect 36004 3602 36032 4082
rect 35992 3596 36044 3602
rect 35992 3538 36044 3544
rect 35716 3392 35768 3398
rect 35716 3334 35768 3340
rect 34520 3052 34572 3058
rect 34520 2994 34572 3000
rect 35440 3052 35492 3058
rect 35440 2994 35492 3000
rect 35728 2990 35756 3334
rect 35716 2984 35768 2990
rect 35716 2926 35768 2932
rect 36360 2916 36412 2922
rect 36360 2858 36412 2864
rect 33876 2576 33928 2582
rect 33876 2518 33928 2524
rect 33416 2508 33468 2514
rect 33416 2450 33468 2456
rect 33140 2440 33192 2446
rect 33140 2382 33192 2388
rect 34940 2204 35236 2224
rect 34996 2202 35020 2204
rect 35076 2202 35100 2204
rect 35156 2202 35180 2204
rect 35018 2150 35020 2202
rect 35082 2150 35094 2202
rect 35156 2150 35158 2202
rect 34996 2148 35020 2150
rect 35076 2148 35100 2150
rect 35156 2148 35180 2150
rect 34940 2128 35236 2148
rect 34244 2100 34296 2106
rect 34244 2042 34296 2048
rect 32048 1142 32260 1170
rect 32232 800 32260 1142
rect 34256 800 34284 2042
rect 36372 1034 36400 2858
rect 38476 2304 38528 2310
rect 38476 2246 38528 2252
rect 36452 2032 36504 2038
rect 36452 1974 36504 1980
rect 36464 1193 36492 1974
rect 36450 1184 36506 1193
rect 36450 1119 36506 1128
rect 36372 1006 36492 1034
rect 36464 800 36492 1006
rect 38488 800 38516 2246
rect 570 0 626 800
rect 2594 0 2650 800
rect 4618 0 4674 800
rect 6826 0 6882 800
rect 8850 0 8906 800
rect 11058 0 11114 800
rect 13082 0 13138 800
rect 15290 0 15346 800
rect 17314 0 17370 800
rect 19522 0 19578 800
rect 21546 0 21602 800
rect 23754 0 23810 800
rect 25778 0 25834 800
rect 27986 0 28042 800
rect 30010 0 30066 800
rect 32218 0 32274 800
rect 34242 0 34298 800
rect 36450 0 36506 800
rect 38474 0 38530 800
<< via2 >>
rect 1858 38120 1914 38176
rect 9678 38428 9680 38448
rect 9680 38428 9732 38448
rect 9732 38428 9734 38448
rect 9678 38392 9734 38428
rect 4220 38106 4276 38108
rect 4300 38106 4356 38108
rect 4380 38106 4436 38108
rect 4460 38106 4516 38108
rect 4220 38054 4246 38106
rect 4246 38054 4276 38106
rect 4300 38054 4310 38106
rect 4310 38054 4356 38106
rect 4380 38054 4426 38106
rect 4426 38054 4436 38106
rect 4460 38054 4490 38106
rect 4490 38054 4516 38106
rect 4220 38052 4276 38054
rect 4300 38052 4356 38054
rect 4380 38052 4436 38054
rect 4460 38052 4516 38054
rect 4220 37018 4276 37020
rect 4300 37018 4356 37020
rect 4380 37018 4436 37020
rect 4460 37018 4516 37020
rect 4220 36966 4246 37018
rect 4246 36966 4276 37018
rect 4300 36966 4310 37018
rect 4310 36966 4356 37018
rect 4380 36966 4426 37018
rect 4426 36966 4436 37018
rect 4460 36966 4490 37018
rect 4490 36966 4516 37018
rect 4220 36964 4276 36966
rect 4300 36964 4356 36966
rect 4380 36964 4436 36966
rect 4460 36964 4516 36966
rect 4220 35930 4276 35932
rect 4300 35930 4356 35932
rect 4380 35930 4436 35932
rect 4460 35930 4516 35932
rect 4220 35878 4246 35930
rect 4246 35878 4276 35930
rect 4300 35878 4310 35930
rect 4310 35878 4356 35930
rect 4380 35878 4426 35930
rect 4426 35878 4436 35930
rect 4460 35878 4490 35930
rect 4490 35878 4516 35930
rect 4220 35876 4276 35878
rect 4300 35876 4356 35878
rect 4380 35876 4436 35878
rect 4460 35876 4516 35878
rect 3606 35128 3662 35184
rect 2870 31864 2926 31920
rect 3054 28872 3110 28928
rect 1582 22616 1638 22672
rect 2778 19236 2834 19272
rect 2778 19216 2780 19236
rect 2780 19216 2832 19236
rect 2832 19216 2834 19236
rect 3330 16652 3386 16688
rect 3330 16632 3332 16652
rect 3332 16632 3384 16652
rect 3384 16632 3386 16652
rect 2502 14728 2558 14784
rect 2778 10104 2834 10160
rect 4220 34842 4276 34844
rect 4300 34842 4356 34844
rect 4380 34842 4436 34844
rect 4460 34842 4516 34844
rect 4220 34790 4246 34842
rect 4246 34790 4276 34842
rect 4300 34790 4310 34842
rect 4310 34790 4356 34842
rect 4380 34790 4426 34842
rect 4426 34790 4436 34842
rect 4460 34790 4490 34842
rect 4490 34790 4516 34842
rect 4220 34788 4276 34790
rect 4300 34788 4356 34790
rect 4380 34788 4436 34790
rect 4460 34788 4516 34790
rect 4220 33754 4276 33756
rect 4300 33754 4356 33756
rect 4380 33754 4436 33756
rect 4460 33754 4516 33756
rect 4220 33702 4246 33754
rect 4246 33702 4276 33754
rect 4300 33702 4310 33754
rect 4310 33702 4356 33754
rect 4380 33702 4426 33754
rect 4426 33702 4436 33754
rect 4460 33702 4490 33754
rect 4490 33702 4516 33754
rect 4220 33700 4276 33702
rect 4300 33700 4356 33702
rect 4380 33700 4436 33702
rect 4460 33700 4516 33702
rect 4220 32666 4276 32668
rect 4300 32666 4356 32668
rect 4380 32666 4436 32668
rect 4460 32666 4516 32668
rect 4220 32614 4246 32666
rect 4246 32614 4276 32666
rect 4300 32614 4310 32666
rect 4310 32614 4356 32666
rect 4380 32614 4426 32666
rect 4426 32614 4436 32666
rect 4460 32614 4490 32666
rect 4490 32614 4516 32666
rect 4220 32612 4276 32614
rect 4300 32612 4356 32614
rect 4380 32612 4436 32614
rect 4460 32612 4516 32614
rect 4220 31578 4276 31580
rect 4300 31578 4356 31580
rect 4380 31578 4436 31580
rect 4460 31578 4516 31580
rect 4220 31526 4246 31578
rect 4246 31526 4276 31578
rect 4300 31526 4310 31578
rect 4310 31526 4356 31578
rect 4380 31526 4426 31578
rect 4426 31526 4436 31578
rect 4460 31526 4490 31578
rect 4490 31526 4516 31578
rect 4220 31524 4276 31526
rect 4300 31524 4356 31526
rect 4380 31524 4436 31526
rect 4460 31524 4516 31526
rect 4220 30490 4276 30492
rect 4300 30490 4356 30492
rect 4380 30490 4436 30492
rect 4460 30490 4516 30492
rect 4220 30438 4246 30490
rect 4246 30438 4276 30490
rect 4300 30438 4310 30490
rect 4310 30438 4356 30490
rect 4380 30438 4426 30490
rect 4426 30438 4436 30490
rect 4460 30438 4490 30490
rect 4490 30438 4516 30490
rect 4220 30436 4276 30438
rect 4300 30436 4356 30438
rect 4380 30436 4436 30438
rect 4460 30436 4516 30438
rect 4220 29402 4276 29404
rect 4300 29402 4356 29404
rect 4380 29402 4436 29404
rect 4460 29402 4516 29404
rect 4220 29350 4246 29402
rect 4246 29350 4276 29402
rect 4300 29350 4310 29402
rect 4310 29350 4356 29402
rect 4380 29350 4426 29402
rect 4426 29350 4436 29402
rect 4460 29350 4490 29402
rect 4490 29350 4516 29402
rect 4220 29348 4276 29350
rect 4300 29348 4356 29350
rect 4380 29348 4436 29350
rect 4460 29348 4516 29350
rect 4220 28314 4276 28316
rect 4300 28314 4356 28316
rect 4380 28314 4436 28316
rect 4460 28314 4516 28316
rect 4220 28262 4246 28314
rect 4246 28262 4276 28314
rect 4300 28262 4310 28314
rect 4310 28262 4356 28314
rect 4380 28262 4426 28314
rect 4426 28262 4436 28314
rect 4460 28262 4490 28314
rect 4490 28262 4516 28314
rect 4220 28260 4276 28262
rect 4300 28260 4356 28262
rect 4380 28260 4436 28262
rect 4460 28260 4516 28262
rect 4220 27226 4276 27228
rect 4300 27226 4356 27228
rect 4380 27226 4436 27228
rect 4460 27226 4516 27228
rect 4220 27174 4246 27226
rect 4246 27174 4276 27226
rect 4300 27174 4310 27226
rect 4310 27174 4356 27226
rect 4380 27174 4426 27226
rect 4426 27174 4436 27226
rect 4460 27174 4490 27226
rect 4490 27174 4516 27226
rect 4220 27172 4276 27174
rect 4300 27172 4356 27174
rect 4380 27172 4436 27174
rect 4460 27172 4516 27174
rect 4220 26138 4276 26140
rect 4300 26138 4356 26140
rect 4380 26138 4436 26140
rect 4460 26138 4516 26140
rect 4220 26086 4246 26138
rect 4246 26086 4276 26138
rect 4300 26086 4310 26138
rect 4310 26086 4356 26138
rect 4380 26086 4426 26138
rect 4426 26086 4436 26138
rect 4460 26086 4490 26138
rect 4490 26086 4516 26138
rect 4220 26084 4276 26086
rect 4300 26084 4356 26086
rect 4380 26084 4436 26086
rect 4460 26084 4516 26086
rect 3974 25608 4030 25664
rect 4220 25050 4276 25052
rect 4300 25050 4356 25052
rect 4380 25050 4436 25052
rect 4460 25050 4516 25052
rect 4220 24998 4246 25050
rect 4246 24998 4276 25050
rect 4300 24998 4310 25050
rect 4310 24998 4356 25050
rect 4380 24998 4426 25050
rect 4426 24998 4436 25050
rect 4460 24998 4490 25050
rect 4490 24998 4516 25050
rect 4220 24996 4276 24998
rect 4300 24996 4356 24998
rect 4380 24996 4436 24998
rect 4460 24996 4516 24998
rect 4220 23962 4276 23964
rect 4300 23962 4356 23964
rect 4380 23962 4436 23964
rect 4460 23962 4516 23964
rect 4220 23910 4246 23962
rect 4246 23910 4276 23962
rect 4300 23910 4310 23962
rect 4310 23910 4356 23962
rect 4380 23910 4426 23962
rect 4426 23910 4436 23962
rect 4460 23910 4490 23962
rect 4490 23910 4516 23962
rect 4220 23908 4276 23910
rect 4300 23908 4356 23910
rect 4380 23908 4436 23910
rect 4460 23908 4516 23910
rect 4220 22874 4276 22876
rect 4300 22874 4356 22876
rect 4380 22874 4436 22876
rect 4460 22874 4516 22876
rect 4220 22822 4246 22874
rect 4246 22822 4276 22874
rect 4300 22822 4310 22874
rect 4310 22822 4356 22874
rect 4380 22822 4426 22874
rect 4426 22822 4436 22874
rect 4460 22822 4490 22874
rect 4490 22822 4516 22874
rect 4220 22820 4276 22822
rect 4300 22820 4356 22822
rect 4380 22820 4436 22822
rect 4460 22820 4516 22822
rect 4220 21786 4276 21788
rect 4300 21786 4356 21788
rect 4380 21786 4436 21788
rect 4460 21786 4516 21788
rect 4220 21734 4246 21786
rect 4246 21734 4276 21786
rect 4300 21734 4310 21786
rect 4310 21734 4356 21786
rect 4380 21734 4426 21786
rect 4426 21734 4436 21786
rect 4460 21734 4490 21786
rect 4490 21734 4516 21786
rect 4220 21732 4276 21734
rect 4300 21732 4356 21734
rect 4380 21732 4436 21734
rect 4460 21732 4516 21734
rect 4220 20698 4276 20700
rect 4300 20698 4356 20700
rect 4380 20698 4436 20700
rect 4460 20698 4516 20700
rect 4220 20646 4246 20698
rect 4246 20646 4276 20698
rect 4300 20646 4310 20698
rect 4310 20646 4356 20698
rect 4380 20646 4426 20698
rect 4426 20646 4436 20698
rect 4460 20646 4490 20698
rect 4490 20646 4516 20698
rect 4220 20644 4276 20646
rect 4300 20644 4356 20646
rect 4380 20644 4436 20646
rect 4460 20644 4516 20646
rect 3698 19252 3700 19272
rect 3700 19252 3752 19272
rect 3752 19252 3754 19272
rect 3698 19216 3754 19252
rect 4220 19610 4276 19612
rect 4300 19610 4356 19612
rect 4380 19610 4436 19612
rect 4460 19610 4516 19612
rect 4220 19558 4246 19610
rect 4246 19558 4276 19610
rect 4300 19558 4310 19610
rect 4310 19558 4356 19610
rect 4380 19558 4426 19610
rect 4426 19558 4436 19610
rect 4460 19558 4490 19610
rect 4490 19558 4516 19610
rect 4220 19556 4276 19558
rect 4300 19556 4356 19558
rect 4380 19556 4436 19558
rect 4460 19556 4516 19558
rect 4066 19352 4122 19408
rect 4220 18522 4276 18524
rect 4300 18522 4356 18524
rect 4380 18522 4436 18524
rect 4460 18522 4516 18524
rect 4220 18470 4246 18522
rect 4246 18470 4276 18522
rect 4300 18470 4310 18522
rect 4310 18470 4356 18522
rect 4380 18470 4426 18522
rect 4426 18470 4436 18522
rect 4460 18470 4490 18522
rect 4490 18470 4516 18522
rect 4220 18468 4276 18470
rect 4300 18468 4356 18470
rect 4380 18468 4436 18470
rect 4460 18468 4516 18470
rect 4220 17434 4276 17436
rect 4300 17434 4356 17436
rect 4380 17434 4436 17436
rect 4460 17434 4516 17436
rect 4220 17382 4246 17434
rect 4246 17382 4276 17434
rect 4300 17382 4310 17434
rect 4310 17382 4356 17434
rect 4380 17382 4426 17434
rect 4426 17382 4436 17434
rect 4460 17382 4490 17434
rect 4490 17382 4516 17434
rect 4220 17380 4276 17382
rect 4300 17380 4356 17382
rect 4380 17380 4436 17382
rect 4460 17380 4516 17382
rect 4434 16632 4490 16688
rect 4066 16396 4068 16416
rect 4068 16396 4120 16416
rect 4120 16396 4122 16416
rect 4066 16360 4122 16396
rect 4220 16346 4276 16348
rect 4300 16346 4356 16348
rect 4380 16346 4436 16348
rect 4460 16346 4516 16348
rect 4220 16294 4246 16346
rect 4246 16294 4276 16346
rect 4300 16294 4310 16346
rect 4310 16294 4356 16346
rect 4380 16294 4426 16346
rect 4426 16294 4436 16346
rect 4460 16294 4490 16346
rect 4490 16294 4516 16346
rect 4220 16292 4276 16294
rect 4300 16292 4356 16294
rect 4380 16292 4436 16294
rect 4460 16292 4516 16294
rect 4220 15258 4276 15260
rect 4300 15258 4356 15260
rect 4380 15258 4436 15260
rect 4460 15258 4516 15260
rect 4220 15206 4246 15258
rect 4246 15206 4276 15258
rect 4300 15206 4310 15258
rect 4310 15206 4356 15258
rect 4380 15206 4426 15258
rect 4426 15206 4436 15258
rect 4460 15206 4490 15258
rect 4490 15206 4516 15258
rect 4220 15204 4276 15206
rect 4300 15204 4356 15206
rect 4380 15204 4436 15206
rect 4460 15204 4516 15206
rect 4220 14170 4276 14172
rect 4300 14170 4356 14172
rect 4380 14170 4436 14172
rect 4460 14170 4516 14172
rect 4220 14118 4246 14170
rect 4246 14118 4276 14170
rect 4300 14118 4310 14170
rect 4310 14118 4356 14170
rect 4380 14118 4426 14170
rect 4426 14118 4436 14170
rect 4460 14118 4490 14170
rect 4490 14118 4516 14170
rect 4220 14116 4276 14118
rect 4300 14116 4356 14118
rect 4380 14116 4436 14118
rect 4460 14116 4516 14118
rect 5906 20340 5908 20360
rect 5908 20340 5960 20360
rect 5960 20340 5962 20360
rect 5906 20304 5962 20340
rect 6090 17740 6146 17776
rect 6090 17720 6092 17740
rect 6092 17720 6144 17740
rect 6144 17720 6146 17740
rect 7102 17740 7158 17776
rect 7102 17720 7104 17740
rect 7104 17720 7156 17740
rect 7156 17720 7158 17740
rect 5446 14476 5502 14512
rect 5446 14456 5448 14476
rect 5448 14456 5500 14476
rect 5500 14456 5502 14476
rect 4220 13082 4276 13084
rect 4300 13082 4356 13084
rect 4380 13082 4436 13084
rect 4460 13082 4516 13084
rect 4220 13030 4246 13082
rect 4246 13030 4276 13082
rect 4300 13030 4310 13082
rect 4310 13030 4356 13082
rect 4380 13030 4426 13082
rect 4426 13030 4436 13082
rect 4460 13030 4490 13082
rect 4490 13030 4516 13082
rect 4220 13028 4276 13030
rect 4300 13028 4356 13030
rect 4380 13028 4436 13030
rect 4460 13028 4516 13030
rect 4220 11994 4276 11996
rect 4300 11994 4356 11996
rect 4380 11994 4436 11996
rect 4460 11994 4516 11996
rect 4220 11942 4246 11994
rect 4246 11942 4276 11994
rect 4300 11942 4310 11994
rect 4310 11942 4356 11994
rect 4380 11942 4426 11994
rect 4426 11942 4436 11994
rect 4460 11942 4490 11994
rect 4490 11942 4516 11994
rect 4220 11940 4276 11942
rect 4300 11940 4356 11942
rect 4380 11940 4436 11942
rect 4460 11940 4516 11942
rect 4220 10906 4276 10908
rect 4300 10906 4356 10908
rect 4380 10906 4436 10908
rect 4460 10906 4516 10908
rect 4220 10854 4246 10906
rect 4246 10854 4276 10906
rect 4300 10854 4310 10906
rect 4310 10854 4356 10906
rect 4380 10854 4426 10906
rect 4426 10854 4436 10906
rect 4460 10854 4490 10906
rect 4490 10854 4516 10906
rect 4220 10852 4276 10854
rect 4300 10852 4356 10854
rect 4380 10852 4436 10854
rect 4460 10852 4516 10854
rect 4220 9818 4276 9820
rect 4300 9818 4356 9820
rect 4380 9818 4436 9820
rect 4460 9818 4516 9820
rect 4220 9766 4246 9818
rect 4246 9766 4276 9818
rect 4300 9766 4310 9818
rect 4310 9766 4356 9818
rect 4380 9766 4426 9818
rect 4426 9766 4436 9818
rect 4460 9766 4490 9818
rect 4490 9766 4516 9818
rect 4220 9764 4276 9766
rect 4300 9764 4356 9766
rect 4380 9764 4436 9766
rect 4460 9764 4516 9766
rect 2962 6568 3018 6624
rect 4220 8730 4276 8732
rect 4300 8730 4356 8732
rect 4380 8730 4436 8732
rect 4460 8730 4516 8732
rect 4220 8678 4246 8730
rect 4246 8678 4276 8730
rect 4300 8678 4310 8730
rect 4310 8678 4356 8730
rect 4380 8678 4426 8730
rect 4426 8678 4436 8730
rect 4460 8678 4490 8730
rect 4490 8678 4516 8730
rect 4220 8676 4276 8678
rect 4300 8676 4356 8678
rect 4380 8676 4436 8678
rect 4460 8676 4516 8678
rect 4220 7642 4276 7644
rect 4300 7642 4356 7644
rect 4380 7642 4436 7644
rect 4460 7642 4516 7644
rect 4220 7590 4246 7642
rect 4246 7590 4276 7642
rect 4300 7590 4310 7642
rect 4310 7590 4356 7642
rect 4380 7590 4426 7642
rect 4426 7590 4436 7642
rect 4460 7590 4490 7642
rect 4490 7590 4516 7642
rect 4220 7588 4276 7590
rect 4300 7588 4356 7590
rect 4380 7588 4436 7590
rect 4460 7588 4516 7590
rect 4220 6554 4276 6556
rect 4300 6554 4356 6556
rect 4380 6554 4436 6556
rect 4460 6554 4516 6556
rect 4220 6502 4246 6554
rect 4246 6502 4276 6554
rect 4300 6502 4310 6554
rect 4310 6502 4356 6554
rect 4380 6502 4426 6554
rect 4426 6502 4436 6554
rect 4460 6502 4490 6554
rect 4490 6502 4516 6554
rect 4220 6500 4276 6502
rect 4300 6500 4356 6502
rect 4380 6500 4436 6502
rect 4460 6500 4516 6502
rect 4220 5466 4276 5468
rect 4300 5466 4356 5468
rect 4380 5466 4436 5468
rect 4460 5466 4516 5468
rect 4220 5414 4246 5466
rect 4246 5414 4276 5466
rect 4300 5414 4310 5466
rect 4310 5414 4356 5466
rect 4380 5414 4426 5466
rect 4426 5414 4436 5466
rect 4460 5414 4490 5466
rect 4490 5414 4516 5466
rect 4220 5412 4276 5414
rect 4300 5412 4356 5414
rect 4380 5412 4436 5414
rect 4460 5412 4516 5414
rect 5814 13812 5816 13832
rect 5816 13812 5868 13832
rect 5868 13812 5870 13832
rect 5814 13776 5870 13812
rect 4220 4378 4276 4380
rect 4300 4378 4356 4380
rect 4380 4378 4436 4380
rect 4460 4378 4516 4380
rect 4220 4326 4246 4378
rect 4246 4326 4276 4378
rect 4300 4326 4310 4378
rect 4310 4326 4356 4378
rect 4380 4326 4426 4378
rect 4426 4326 4436 4378
rect 4460 4326 4490 4378
rect 4490 4326 4516 4378
rect 4220 4324 4276 4326
rect 4300 4324 4356 4326
rect 4380 4324 4436 4326
rect 4460 4324 4516 4326
rect 4220 3290 4276 3292
rect 4300 3290 4356 3292
rect 4380 3290 4436 3292
rect 4460 3290 4516 3292
rect 4220 3238 4246 3290
rect 4246 3238 4276 3290
rect 4300 3238 4310 3290
rect 4310 3238 4356 3290
rect 4380 3238 4426 3290
rect 4426 3238 4436 3290
rect 4460 3238 4490 3290
rect 4490 3238 4516 3290
rect 4220 3236 4276 3238
rect 4300 3236 4356 3238
rect 4380 3236 4436 3238
rect 4460 3236 4516 3238
rect 9586 30096 9642 30152
rect 8022 20304 8078 20360
rect 10414 19896 10470 19952
rect 9770 18672 9826 18728
rect 7102 4020 7104 4040
rect 7104 4020 7156 4040
rect 7156 4020 7158 4040
rect 7102 3984 7158 4020
rect 8942 14728 8998 14784
rect 8758 5772 8814 5808
rect 8758 5752 8760 5772
rect 8760 5752 8812 5772
rect 8812 5752 8814 5772
rect 4220 2202 4276 2204
rect 4300 2202 4356 2204
rect 4380 2202 4436 2204
rect 4460 2202 4516 2204
rect 4220 2150 4246 2202
rect 4246 2150 4276 2202
rect 4300 2150 4310 2202
rect 4310 2150 4356 2202
rect 4380 2150 4426 2202
rect 4426 2150 4436 2202
rect 4460 2150 4490 2202
rect 4490 2150 4516 2202
rect 4220 2148 4276 2150
rect 4300 2148 4356 2150
rect 4380 2148 4436 2150
rect 4460 2148 4516 2150
rect 12162 23296 12218 23352
rect 12990 24284 12992 24304
rect 12992 24284 13044 24304
rect 13044 24284 13046 24304
rect 12990 24248 13046 24284
rect 10322 14728 10378 14784
rect 9954 13232 10010 13288
rect 9310 4020 9312 4040
rect 9312 4020 9364 4040
rect 9364 4020 9366 4040
rect 9310 3984 9366 4020
rect 9218 3848 9274 3904
rect 11702 15408 11758 15464
rect 11702 14764 11704 14784
rect 11704 14764 11756 14784
rect 11756 14764 11758 14784
rect 11702 14728 11758 14764
rect 12622 15000 12678 15056
rect 11518 5616 11574 5672
rect 12714 11772 12716 11792
rect 12716 11772 12768 11792
rect 12768 11772 12770 11792
rect 12714 11736 12770 11772
rect 13818 20204 13820 20224
rect 13820 20204 13872 20224
rect 13872 20204 13874 20224
rect 13818 20168 13874 20204
rect 13358 5888 13414 5944
rect 15842 30132 15844 30152
rect 15844 30132 15896 30152
rect 15896 30132 15898 30152
rect 15842 30096 15898 30132
rect 14002 6296 14058 6352
rect 12898 3712 12954 3768
rect 15198 14320 15254 14376
rect 15106 11736 15162 11792
rect 19580 38650 19636 38652
rect 19660 38650 19716 38652
rect 19740 38650 19796 38652
rect 19820 38650 19876 38652
rect 19580 38598 19606 38650
rect 19606 38598 19636 38650
rect 19660 38598 19670 38650
rect 19670 38598 19716 38650
rect 19740 38598 19786 38650
rect 19786 38598 19796 38650
rect 19820 38598 19850 38650
rect 19850 38598 19876 38650
rect 19580 38596 19636 38598
rect 19660 38596 19716 38598
rect 19740 38596 19796 38598
rect 19820 38596 19876 38598
rect 19154 38392 19210 38448
rect 16670 19252 16672 19272
rect 16672 19252 16724 19272
rect 16724 19252 16726 19272
rect 16670 19216 16726 19252
rect 16762 18672 16818 18728
rect 15474 12552 15530 12608
rect 15842 6296 15898 6352
rect 16026 5888 16082 5944
rect 17130 15000 17186 15056
rect 17038 13912 17094 13968
rect 17130 13232 17186 13288
rect 17590 20168 17646 20224
rect 17590 19216 17646 19272
rect 16762 6740 16764 6760
rect 16764 6740 16816 6760
rect 16816 6740 16818 6760
rect 16762 6704 16818 6740
rect 18142 15444 18144 15464
rect 18144 15444 18196 15464
rect 18196 15444 18198 15464
rect 18142 15408 18198 15444
rect 18602 29008 18658 29064
rect 19580 37562 19636 37564
rect 19660 37562 19716 37564
rect 19740 37562 19796 37564
rect 19820 37562 19876 37564
rect 19580 37510 19606 37562
rect 19606 37510 19636 37562
rect 19660 37510 19670 37562
rect 19670 37510 19716 37562
rect 19740 37510 19786 37562
rect 19786 37510 19796 37562
rect 19820 37510 19850 37562
rect 19850 37510 19876 37562
rect 19580 37508 19636 37510
rect 19660 37508 19716 37510
rect 19740 37508 19796 37510
rect 19820 37508 19876 37510
rect 19580 36474 19636 36476
rect 19660 36474 19716 36476
rect 19740 36474 19796 36476
rect 19820 36474 19876 36476
rect 19580 36422 19606 36474
rect 19606 36422 19636 36474
rect 19660 36422 19670 36474
rect 19670 36422 19716 36474
rect 19740 36422 19786 36474
rect 19786 36422 19796 36474
rect 19820 36422 19850 36474
rect 19850 36422 19876 36474
rect 19580 36420 19636 36422
rect 19660 36420 19716 36422
rect 19740 36420 19796 36422
rect 19820 36420 19876 36422
rect 19580 35386 19636 35388
rect 19660 35386 19716 35388
rect 19740 35386 19796 35388
rect 19820 35386 19876 35388
rect 19580 35334 19606 35386
rect 19606 35334 19636 35386
rect 19660 35334 19670 35386
rect 19670 35334 19716 35386
rect 19740 35334 19786 35386
rect 19786 35334 19796 35386
rect 19820 35334 19850 35386
rect 19850 35334 19876 35386
rect 19580 35332 19636 35334
rect 19660 35332 19716 35334
rect 19740 35332 19796 35334
rect 19820 35332 19876 35334
rect 19580 34298 19636 34300
rect 19660 34298 19716 34300
rect 19740 34298 19796 34300
rect 19820 34298 19876 34300
rect 19580 34246 19606 34298
rect 19606 34246 19636 34298
rect 19660 34246 19670 34298
rect 19670 34246 19716 34298
rect 19740 34246 19786 34298
rect 19786 34246 19796 34298
rect 19820 34246 19850 34298
rect 19850 34246 19876 34298
rect 19580 34244 19636 34246
rect 19660 34244 19716 34246
rect 19740 34244 19796 34246
rect 19820 34244 19876 34246
rect 19580 33210 19636 33212
rect 19660 33210 19716 33212
rect 19740 33210 19796 33212
rect 19820 33210 19876 33212
rect 19580 33158 19606 33210
rect 19606 33158 19636 33210
rect 19660 33158 19670 33210
rect 19670 33158 19716 33210
rect 19740 33158 19786 33210
rect 19786 33158 19796 33210
rect 19820 33158 19850 33210
rect 19850 33158 19876 33210
rect 19580 33156 19636 33158
rect 19660 33156 19716 33158
rect 19740 33156 19796 33158
rect 19820 33156 19876 33158
rect 19580 32122 19636 32124
rect 19660 32122 19716 32124
rect 19740 32122 19796 32124
rect 19820 32122 19876 32124
rect 19580 32070 19606 32122
rect 19606 32070 19636 32122
rect 19660 32070 19670 32122
rect 19670 32070 19716 32122
rect 19740 32070 19786 32122
rect 19786 32070 19796 32122
rect 19820 32070 19850 32122
rect 19850 32070 19876 32122
rect 19580 32068 19636 32070
rect 19660 32068 19716 32070
rect 19740 32068 19796 32070
rect 19820 32068 19876 32070
rect 19580 31034 19636 31036
rect 19660 31034 19716 31036
rect 19740 31034 19796 31036
rect 19820 31034 19876 31036
rect 19580 30982 19606 31034
rect 19606 30982 19636 31034
rect 19660 30982 19670 31034
rect 19670 30982 19716 31034
rect 19740 30982 19786 31034
rect 19786 30982 19796 31034
rect 19820 30982 19850 31034
rect 19850 30982 19876 31034
rect 19580 30980 19636 30982
rect 19660 30980 19716 30982
rect 19740 30980 19796 30982
rect 19820 30980 19876 30982
rect 18878 28908 18880 28928
rect 18880 28908 18932 28928
rect 18932 28908 18934 28928
rect 18878 28872 18934 28908
rect 18510 28464 18566 28520
rect 19580 29946 19636 29948
rect 19660 29946 19716 29948
rect 19740 29946 19796 29948
rect 19820 29946 19876 29948
rect 19580 29894 19606 29946
rect 19606 29894 19636 29946
rect 19660 29894 19670 29946
rect 19670 29894 19716 29946
rect 19740 29894 19786 29946
rect 19786 29894 19796 29946
rect 19820 29894 19850 29946
rect 19850 29894 19876 29946
rect 19580 29892 19636 29894
rect 19660 29892 19716 29894
rect 19740 29892 19796 29894
rect 19820 29892 19876 29894
rect 19580 28858 19636 28860
rect 19660 28858 19716 28860
rect 19740 28858 19796 28860
rect 19820 28858 19876 28860
rect 19580 28806 19606 28858
rect 19606 28806 19636 28858
rect 19660 28806 19670 28858
rect 19670 28806 19716 28858
rect 19740 28806 19786 28858
rect 19786 28806 19796 28858
rect 19820 28806 19850 28858
rect 19850 28806 19876 28858
rect 19580 28804 19636 28806
rect 19660 28804 19716 28806
rect 19740 28804 19796 28806
rect 19820 28804 19876 28806
rect 19580 27770 19636 27772
rect 19660 27770 19716 27772
rect 19740 27770 19796 27772
rect 19820 27770 19876 27772
rect 19580 27718 19606 27770
rect 19606 27718 19636 27770
rect 19660 27718 19670 27770
rect 19670 27718 19716 27770
rect 19740 27718 19786 27770
rect 19786 27718 19796 27770
rect 19820 27718 19850 27770
rect 19850 27718 19876 27770
rect 19580 27716 19636 27718
rect 19660 27716 19716 27718
rect 19740 27716 19796 27718
rect 19820 27716 19876 27718
rect 19580 26682 19636 26684
rect 19660 26682 19716 26684
rect 19740 26682 19796 26684
rect 19820 26682 19876 26684
rect 19580 26630 19606 26682
rect 19606 26630 19636 26682
rect 19660 26630 19670 26682
rect 19670 26630 19716 26682
rect 19740 26630 19786 26682
rect 19786 26630 19796 26682
rect 19820 26630 19850 26682
rect 19850 26630 19876 26682
rect 19580 26628 19636 26630
rect 19660 26628 19716 26630
rect 19740 26628 19796 26630
rect 19820 26628 19876 26630
rect 19580 25594 19636 25596
rect 19660 25594 19716 25596
rect 19740 25594 19796 25596
rect 19820 25594 19876 25596
rect 19580 25542 19606 25594
rect 19606 25542 19636 25594
rect 19660 25542 19670 25594
rect 19670 25542 19716 25594
rect 19740 25542 19786 25594
rect 19786 25542 19796 25594
rect 19820 25542 19850 25594
rect 19850 25542 19876 25594
rect 19580 25540 19636 25542
rect 19660 25540 19716 25542
rect 19740 25540 19796 25542
rect 19820 25540 19876 25542
rect 19580 24506 19636 24508
rect 19660 24506 19716 24508
rect 19740 24506 19796 24508
rect 19820 24506 19876 24508
rect 19580 24454 19606 24506
rect 19606 24454 19636 24506
rect 19660 24454 19670 24506
rect 19670 24454 19716 24506
rect 19740 24454 19786 24506
rect 19786 24454 19796 24506
rect 19820 24454 19850 24506
rect 19850 24454 19876 24506
rect 19580 24452 19636 24454
rect 19660 24452 19716 24454
rect 19740 24452 19796 24454
rect 19820 24452 19876 24454
rect 18510 24284 18512 24304
rect 18512 24284 18564 24304
rect 18564 24284 18566 24304
rect 18510 24248 18566 24284
rect 19580 23418 19636 23420
rect 19660 23418 19716 23420
rect 19740 23418 19796 23420
rect 19820 23418 19876 23420
rect 19580 23366 19606 23418
rect 19606 23366 19636 23418
rect 19660 23366 19670 23418
rect 19670 23366 19716 23418
rect 19740 23366 19786 23418
rect 19786 23366 19796 23418
rect 19820 23366 19850 23418
rect 19850 23366 19876 23418
rect 19580 23364 19636 23366
rect 19660 23364 19716 23366
rect 19740 23364 19796 23366
rect 19820 23364 19876 23366
rect 18878 23296 18934 23352
rect 18878 23160 18934 23216
rect 18418 19896 18474 19952
rect 19580 22330 19636 22332
rect 19660 22330 19716 22332
rect 19740 22330 19796 22332
rect 19820 22330 19876 22332
rect 19580 22278 19606 22330
rect 19606 22278 19636 22330
rect 19660 22278 19670 22330
rect 19670 22278 19716 22330
rect 19740 22278 19786 22330
rect 19786 22278 19796 22330
rect 19820 22278 19850 22330
rect 19850 22278 19876 22330
rect 19580 22276 19636 22278
rect 19660 22276 19716 22278
rect 19740 22276 19796 22278
rect 19820 22276 19876 22278
rect 19890 21528 19946 21584
rect 19580 21242 19636 21244
rect 19660 21242 19716 21244
rect 19740 21242 19796 21244
rect 19820 21242 19876 21244
rect 19580 21190 19606 21242
rect 19606 21190 19636 21242
rect 19660 21190 19670 21242
rect 19670 21190 19716 21242
rect 19740 21190 19786 21242
rect 19786 21190 19796 21242
rect 19820 21190 19850 21242
rect 19850 21190 19876 21242
rect 19580 21188 19636 21190
rect 19660 21188 19716 21190
rect 19740 21188 19796 21190
rect 19820 21188 19876 21190
rect 19580 20154 19636 20156
rect 19660 20154 19716 20156
rect 19740 20154 19796 20156
rect 19820 20154 19876 20156
rect 19580 20102 19606 20154
rect 19606 20102 19636 20154
rect 19660 20102 19670 20154
rect 19670 20102 19716 20154
rect 19740 20102 19786 20154
rect 19786 20102 19796 20154
rect 19820 20102 19850 20154
rect 19850 20102 19876 20154
rect 19580 20100 19636 20102
rect 19660 20100 19716 20102
rect 19740 20100 19796 20102
rect 19820 20100 19876 20102
rect 19580 19066 19636 19068
rect 19660 19066 19716 19068
rect 19740 19066 19796 19068
rect 19820 19066 19876 19068
rect 19580 19014 19606 19066
rect 19606 19014 19636 19066
rect 19660 19014 19670 19066
rect 19670 19014 19716 19066
rect 19740 19014 19786 19066
rect 19786 19014 19796 19066
rect 19820 19014 19850 19066
rect 19850 19014 19876 19066
rect 19580 19012 19636 19014
rect 19660 19012 19716 19014
rect 19740 19012 19796 19014
rect 19820 19012 19876 19014
rect 18602 14320 18658 14376
rect 18418 12552 18474 12608
rect 19580 17978 19636 17980
rect 19660 17978 19716 17980
rect 19740 17978 19796 17980
rect 19820 17978 19876 17980
rect 19580 17926 19606 17978
rect 19606 17926 19636 17978
rect 19660 17926 19670 17978
rect 19670 17926 19716 17978
rect 19740 17926 19786 17978
rect 19786 17926 19796 17978
rect 19820 17926 19850 17978
rect 19850 17926 19876 17978
rect 19580 17924 19636 17926
rect 19660 17924 19716 17926
rect 19740 17924 19796 17926
rect 19820 17924 19876 17926
rect 19580 16890 19636 16892
rect 19660 16890 19716 16892
rect 19740 16890 19796 16892
rect 19820 16890 19876 16892
rect 19580 16838 19606 16890
rect 19606 16838 19636 16890
rect 19660 16838 19670 16890
rect 19670 16838 19716 16890
rect 19740 16838 19786 16890
rect 19786 16838 19796 16890
rect 19820 16838 19850 16890
rect 19850 16838 19876 16890
rect 19580 16836 19636 16838
rect 19660 16836 19716 16838
rect 19740 16836 19796 16838
rect 19820 16836 19876 16838
rect 20074 21528 20130 21584
rect 19982 15952 20038 16008
rect 19580 15802 19636 15804
rect 19660 15802 19716 15804
rect 19740 15802 19796 15804
rect 19820 15802 19876 15804
rect 19580 15750 19606 15802
rect 19606 15750 19636 15802
rect 19660 15750 19670 15802
rect 19670 15750 19716 15802
rect 19740 15750 19786 15802
rect 19786 15750 19796 15802
rect 19820 15750 19850 15802
rect 19850 15750 19876 15802
rect 19580 15748 19636 15750
rect 19660 15748 19716 15750
rect 19740 15748 19796 15750
rect 19820 15748 19876 15750
rect 18786 13776 18842 13832
rect 17774 4140 17830 4176
rect 17774 4120 17776 4140
rect 17776 4120 17828 4140
rect 17828 4120 17830 4140
rect 19154 14728 19210 14784
rect 19580 14714 19636 14716
rect 19660 14714 19716 14716
rect 19740 14714 19796 14716
rect 19820 14714 19876 14716
rect 19580 14662 19606 14714
rect 19606 14662 19636 14714
rect 19660 14662 19670 14714
rect 19670 14662 19716 14714
rect 19740 14662 19786 14714
rect 19786 14662 19796 14714
rect 19820 14662 19850 14714
rect 19850 14662 19876 14714
rect 19580 14660 19636 14662
rect 19660 14660 19716 14662
rect 19740 14660 19796 14662
rect 19820 14660 19876 14662
rect 19338 14456 19394 14512
rect 19706 14476 19762 14512
rect 19706 14456 19708 14476
rect 19708 14456 19760 14476
rect 19760 14456 19762 14476
rect 19580 13626 19636 13628
rect 19660 13626 19716 13628
rect 19740 13626 19796 13628
rect 19820 13626 19876 13628
rect 19580 13574 19606 13626
rect 19606 13574 19636 13626
rect 19660 13574 19670 13626
rect 19670 13574 19716 13626
rect 19740 13574 19786 13626
rect 19786 13574 19796 13626
rect 19820 13574 19850 13626
rect 19850 13574 19876 13626
rect 19580 13572 19636 13574
rect 19660 13572 19716 13574
rect 19740 13572 19796 13574
rect 19820 13572 19876 13574
rect 19580 12538 19636 12540
rect 19660 12538 19716 12540
rect 19740 12538 19796 12540
rect 19820 12538 19876 12540
rect 19580 12486 19606 12538
rect 19606 12486 19636 12538
rect 19660 12486 19670 12538
rect 19670 12486 19716 12538
rect 19740 12486 19786 12538
rect 19786 12486 19796 12538
rect 19820 12486 19850 12538
rect 19850 12486 19876 12538
rect 19580 12484 19636 12486
rect 19660 12484 19716 12486
rect 19740 12484 19796 12486
rect 19820 12484 19876 12486
rect 19580 11450 19636 11452
rect 19660 11450 19716 11452
rect 19740 11450 19796 11452
rect 19820 11450 19876 11452
rect 19580 11398 19606 11450
rect 19606 11398 19636 11450
rect 19660 11398 19670 11450
rect 19670 11398 19716 11450
rect 19740 11398 19786 11450
rect 19786 11398 19796 11450
rect 19820 11398 19850 11450
rect 19850 11398 19876 11450
rect 19580 11396 19636 11398
rect 19660 11396 19716 11398
rect 19740 11396 19796 11398
rect 19820 11396 19876 11398
rect 19580 10362 19636 10364
rect 19660 10362 19716 10364
rect 19740 10362 19796 10364
rect 19820 10362 19876 10364
rect 19580 10310 19606 10362
rect 19606 10310 19636 10362
rect 19660 10310 19670 10362
rect 19670 10310 19716 10362
rect 19740 10310 19786 10362
rect 19786 10310 19796 10362
rect 19820 10310 19850 10362
rect 19850 10310 19876 10362
rect 19580 10308 19636 10310
rect 19660 10308 19716 10310
rect 19740 10308 19796 10310
rect 19820 10308 19876 10310
rect 19580 9274 19636 9276
rect 19660 9274 19716 9276
rect 19740 9274 19796 9276
rect 19820 9274 19876 9276
rect 19580 9222 19606 9274
rect 19606 9222 19636 9274
rect 19660 9222 19670 9274
rect 19670 9222 19716 9274
rect 19740 9222 19786 9274
rect 19786 9222 19796 9274
rect 19820 9222 19850 9274
rect 19850 9222 19876 9274
rect 19580 9220 19636 9222
rect 19660 9220 19716 9222
rect 19740 9220 19796 9222
rect 19820 9220 19876 9222
rect 19580 8186 19636 8188
rect 19660 8186 19716 8188
rect 19740 8186 19796 8188
rect 19820 8186 19876 8188
rect 19580 8134 19606 8186
rect 19606 8134 19636 8186
rect 19660 8134 19670 8186
rect 19670 8134 19716 8186
rect 19740 8134 19786 8186
rect 19786 8134 19796 8186
rect 19820 8134 19850 8186
rect 19850 8134 19876 8186
rect 19580 8132 19636 8134
rect 19660 8132 19716 8134
rect 19740 8132 19796 8134
rect 19820 8132 19876 8134
rect 19580 7098 19636 7100
rect 19660 7098 19716 7100
rect 19740 7098 19796 7100
rect 19820 7098 19876 7100
rect 19580 7046 19606 7098
rect 19606 7046 19636 7098
rect 19660 7046 19670 7098
rect 19670 7046 19716 7098
rect 19740 7046 19786 7098
rect 19786 7046 19796 7098
rect 19820 7046 19850 7098
rect 19850 7046 19876 7098
rect 19580 7044 19636 7046
rect 19660 7044 19716 7046
rect 19740 7044 19796 7046
rect 19820 7044 19876 7046
rect 19580 6010 19636 6012
rect 19660 6010 19716 6012
rect 19740 6010 19796 6012
rect 19820 6010 19876 6012
rect 19580 5958 19606 6010
rect 19606 5958 19636 6010
rect 19660 5958 19670 6010
rect 19670 5958 19716 6010
rect 19740 5958 19786 6010
rect 19786 5958 19796 6010
rect 19820 5958 19850 6010
rect 19850 5958 19876 6010
rect 19580 5956 19636 5958
rect 19660 5956 19716 5958
rect 19740 5956 19796 5958
rect 19820 5956 19876 5958
rect 19580 4922 19636 4924
rect 19660 4922 19716 4924
rect 19740 4922 19796 4924
rect 19820 4922 19876 4924
rect 19580 4870 19606 4922
rect 19606 4870 19636 4922
rect 19660 4870 19670 4922
rect 19670 4870 19716 4922
rect 19740 4870 19786 4922
rect 19786 4870 19796 4922
rect 19820 4870 19850 4922
rect 19850 4870 19876 4922
rect 19580 4868 19636 4870
rect 19660 4868 19716 4870
rect 19740 4868 19796 4870
rect 19820 4868 19876 4870
rect 19246 4140 19302 4176
rect 19246 4120 19248 4140
rect 19248 4120 19300 4140
rect 19300 4120 19302 4140
rect 19062 3712 19118 3768
rect 19580 3834 19636 3836
rect 19660 3834 19716 3836
rect 19740 3834 19796 3836
rect 19820 3834 19876 3836
rect 19580 3782 19606 3834
rect 19606 3782 19636 3834
rect 19660 3782 19670 3834
rect 19670 3782 19716 3834
rect 19740 3782 19786 3834
rect 19786 3782 19796 3834
rect 19820 3782 19850 3834
rect 19850 3782 19876 3834
rect 19580 3780 19636 3782
rect 19660 3780 19716 3782
rect 19740 3780 19796 3782
rect 19820 3780 19876 3782
rect 19580 2746 19636 2748
rect 19660 2746 19716 2748
rect 19740 2746 19796 2748
rect 19820 2746 19876 2748
rect 19580 2694 19606 2746
rect 19606 2694 19636 2746
rect 19660 2694 19670 2746
rect 19670 2694 19716 2746
rect 19740 2694 19786 2746
rect 19786 2694 19796 2746
rect 19820 2694 19850 2746
rect 19850 2694 19876 2746
rect 19580 2692 19636 2694
rect 19660 2692 19716 2694
rect 19740 2692 19796 2694
rect 19820 2692 19876 2694
rect 20166 13812 20168 13832
rect 20168 13812 20220 13832
rect 20220 13812 20222 13832
rect 20166 13776 20222 13812
rect 20994 13232 21050 13288
rect 21454 16516 21510 16552
rect 21454 16496 21456 16516
rect 21456 16496 21508 16516
rect 21508 16496 21510 16516
rect 22190 13912 22246 13968
rect 21914 10648 21970 10704
rect 36082 38664 36138 38720
rect 34940 38106 34996 38108
rect 35020 38106 35076 38108
rect 35100 38106 35156 38108
rect 35180 38106 35236 38108
rect 34940 38054 34966 38106
rect 34966 38054 34996 38106
rect 35020 38054 35030 38106
rect 35030 38054 35076 38106
rect 35100 38054 35146 38106
rect 35146 38054 35156 38106
rect 35180 38054 35210 38106
rect 35210 38054 35236 38106
rect 34940 38052 34996 38054
rect 35020 38052 35076 38054
rect 35100 38052 35156 38054
rect 35180 38052 35236 38054
rect 23018 19896 23074 19952
rect 23294 12708 23350 12744
rect 23294 12688 23296 12708
rect 23296 12688 23348 12708
rect 23348 12688 23350 12708
rect 22834 9016 22890 9072
rect 23754 13232 23810 13288
rect 23754 12688 23810 12744
rect 23570 9696 23626 9752
rect 23478 9560 23534 9616
rect 23662 9460 23664 9480
rect 23664 9460 23716 9480
rect 23716 9460 23718 9480
rect 23662 9424 23718 9460
rect 25042 19216 25098 19272
rect 24674 16532 24676 16552
rect 24676 16532 24728 16552
rect 24728 16532 24730 16552
rect 24674 16496 24730 16532
rect 25318 16652 25374 16688
rect 25318 16632 25320 16652
rect 25320 16632 25372 16652
rect 25372 16632 25374 16652
rect 25502 15952 25558 16008
rect 26146 17076 26148 17096
rect 26148 17076 26200 17096
rect 26200 17076 26202 17096
rect 26146 17040 26202 17076
rect 26238 16768 26294 16824
rect 24950 5752 25006 5808
rect 24858 5636 24914 5672
rect 24858 5616 24860 5636
rect 24860 5616 24912 5636
rect 24912 5616 24914 5636
rect 25226 9036 25282 9072
rect 25226 9016 25228 9036
rect 25228 9016 25280 9036
rect 25280 9016 25282 9036
rect 25870 13368 25926 13424
rect 26146 13932 26202 13968
rect 26146 13912 26148 13932
rect 26148 13912 26200 13932
rect 26200 13912 26202 13932
rect 29274 23568 29330 23624
rect 29090 21972 29092 21992
rect 29092 21972 29144 21992
rect 29144 21972 29146 21992
rect 29090 21936 29146 21972
rect 27434 19916 27490 19952
rect 27434 19896 27436 19916
rect 27436 19896 27488 19916
rect 27488 19896 27490 19916
rect 25502 6704 25558 6760
rect 26882 13776 26938 13832
rect 26514 9424 26570 9480
rect 28078 17076 28080 17096
rect 28080 17076 28132 17096
rect 28132 17076 28134 17096
rect 28078 17040 28134 17076
rect 27342 16108 27398 16144
rect 27342 16088 27344 16108
rect 27344 16088 27396 16108
rect 27396 16088 27398 16108
rect 27526 10648 27582 10704
rect 27894 14476 27950 14512
rect 27894 14456 27896 14476
rect 27896 14456 27948 14476
rect 27948 14456 27950 14476
rect 28354 16108 28410 16144
rect 28354 16088 28356 16108
rect 28356 16088 28408 16108
rect 28408 16088 28410 16108
rect 28906 16768 28962 16824
rect 29918 16768 29974 16824
rect 31114 22072 31170 22128
rect 30838 21936 30894 21992
rect 30654 12300 30710 12336
rect 30654 12280 30656 12300
rect 30656 12280 30708 12300
rect 30708 12280 30710 12300
rect 30746 11620 30802 11656
rect 30746 11600 30748 11620
rect 30748 11600 30800 11620
rect 30800 11600 30802 11620
rect 30102 11056 30158 11112
rect 31114 12724 31116 12744
rect 31116 12724 31168 12744
rect 31168 12724 31170 12744
rect 31114 12688 31170 12724
rect 33322 23160 33378 23216
rect 32402 12688 32458 12744
rect 32954 12280 33010 12336
rect 32862 10648 32918 10704
rect 34940 37018 34996 37020
rect 35020 37018 35076 37020
rect 35100 37018 35156 37020
rect 35180 37018 35236 37020
rect 34940 36966 34966 37018
rect 34966 36966 34996 37018
rect 35020 36966 35030 37018
rect 35030 36966 35076 37018
rect 35100 36966 35146 37018
rect 35146 36966 35156 37018
rect 35180 36966 35210 37018
rect 35210 36966 35236 37018
rect 34940 36964 34996 36966
rect 35020 36964 35076 36966
rect 35100 36964 35156 36966
rect 35180 36964 35236 36966
rect 34940 35930 34996 35932
rect 35020 35930 35076 35932
rect 35100 35930 35156 35932
rect 35180 35930 35236 35932
rect 34940 35878 34966 35930
rect 34966 35878 34996 35930
rect 35020 35878 35030 35930
rect 35030 35878 35076 35930
rect 35100 35878 35146 35930
rect 35146 35878 35156 35930
rect 35180 35878 35210 35930
rect 35210 35878 35236 35930
rect 34940 35876 34996 35878
rect 35020 35876 35076 35878
rect 35100 35876 35156 35878
rect 35180 35876 35236 35878
rect 35990 35400 36046 35456
rect 34940 34842 34996 34844
rect 35020 34842 35076 34844
rect 35100 34842 35156 34844
rect 35180 34842 35236 34844
rect 34940 34790 34966 34842
rect 34966 34790 34996 34842
rect 35020 34790 35030 34842
rect 35030 34790 35076 34842
rect 35100 34790 35146 34842
rect 35146 34790 35156 34842
rect 35180 34790 35210 34842
rect 35210 34790 35236 34842
rect 34940 34788 34996 34790
rect 35020 34788 35076 34790
rect 35100 34788 35156 34790
rect 35180 34788 35236 34790
rect 34940 33754 34996 33756
rect 35020 33754 35076 33756
rect 35100 33754 35156 33756
rect 35180 33754 35236 33756
rect 34940 33702 34966 33754
rect 34966 33702 34996 33754
rect 35020 33702 35030 33754
rect 35030 33702 35076 33754
rect 35100 33702 35146 33754
rect 35146 33702 35156 33754
rect 35180 33702 35210 33754
rect 35210 33702 35236 33754
rect 34940 33700 34996 33702
rect 35020 33700 35076 33702
rect 35100 33700 35156 33702
rect 35180 33700 35236 33702
rect 34940 32666 34996 32668
rect 35020 32666 35076 32668
rect 35100 32666 35156 32668
rect 35180 32666 35236 32668
rect 34940 32614 34966 32666
rect 34966 32614 34996 32666
rect 35020 32614 35030 32666
rect 35030 32614 35076 32666
rect 35100 32614 35146 32666
rect 35146 32614 35156 32666
rect 35180 32614 35210 32666
rect 35210 32614 35236 32666
rect 34940 32612 34996 32614
rect 35020 32612 35076 32614
rect 35100 32612 35156 32614
rect 35180 32612 35236 32614
rect 34940 31578 34996 31580
rect 35020 31578 35076 31580
rect 35100 31578 35156 31580
rect 35180 31578 35236 31580
rect 34940 31526 34966 31578
rect 34966 31526 34996 31578
rect 35020 31526 35030 31578
rect 35030 31526 35076 31578
rect 35100 31526 35146 31578
rect 35146 31526 35156 31578
rect 35180 31526 35210 31578
rect 35210 31526 35236 31578
rect 34940 31524 34996 31526
rect 35020 31524 35076 31526
rect 35100 31524 35156 31526
rect 35180 31524 35236 31526
rect 34940 30490 34996 30492
rect 35020 30490 35076 30492
rect 35100 30490 35156 30492
rect 35180 30490 35236 30492
rect 34940 30438 34966 30490
rect 34966 30438 34996 30490
rect 35020 30438 35030 30490
rect 35030 30438 35076 30490
rect 35100 30438 35146 30490
rect 35146 30438 35156 30490
rect 35180 30438 35210 30490
rect 35210 30438 35236 30490
rect 34940 30436 34996 30438
rect 35020 30436 35076 30438
rect 35100 30436 35156 30438
rect 35180 30436 35236 30438
rect 34940 29402 34996 29404
rect 35020 29402 35076 29404
rect 35100 29402 35156 29404
rect 35180 29402 35236 29404
rect 34940 29350 34966 29402
rect 34966 29350 34996 29402
rect 35020 29350 35030 29402
rect 35030 29350 35076 29402
rect 35100 29350 35146 29402
rect 35146 29350 35156 29402
rect 35180 29350 35210 29402
rect 35210 29350 35236 29402
rect 34940 29348 34996 29350
rect 35020 29348 35076 29350
rect 35100 29348 35156 29350
rect 35180 29348 35236 29350
rect 34940 28314 34996 28316
rect 35020 28314 35076 28316
rect 35100 28314 35156 28316
rect 35180 28314 35236 28316
rect 34940 28262 34966 28314
rect 34966 28262 34996 28314
rect 35020 28262 35030 28314
rect 35030 28262 35076 28314
rect 35100 28262 35146 28314
rect 35146 28262 35156 28314
rect 35180 28262 35210 28314
rect 35210 28262 35236 28314
rect 34940 28260 34996 28262
rect 35020 28260 35076 28262
rect 35100 28260 35156 28262
rect 35180 28260 35236 28262
rect 34940 27226 34996 27228
rect 35020 27226 35076 27228
rect 35100 27226 35156 27228
rect 35180 27226 35236 27228
rect 34940 27174 34966 27226
rect 34966 27174 34996 27226
rect 35020 27174 35030 27226
rect 35030 27174 35076 27226
rect 35100 27174 35146 27226
rect 35146 27174 35156 27226
rect 35180 27174 35210 27226
rect 35210 27174 35236 27226
rect 34940 27172 34996 27174
rect 35020 27172 35076 27174
rect 35100 27172 35156 27174
rect 35180 27172 35236 27174
rect 33874 16632 33930 16688
rect 33506 12144 33562 12200
rect 33874 12144 33930 12200
rect 34940 26138 34996 26140
rect 35020 26138 35076 26140
rect 35100 26138 35156 26140
rect 35180 26138 35236 26140
rect 34940 26086 34966 26138
rect 34966 26086 34996 26138
rect 35020 26086 35030 26138
rect 35030 26086 35076 26138
rect 35100 26086 35146 26138
rect 35146 26086 35156 26138
rect 35180 26086 35210 26138
rect 35210 26086 35236 26138
rect 34940 26084 34996 26086
rect 35020 26084 35076 26086
rect 35100 26084 35156 26086
rect 35180 26084 35236 26086
rect 34940 25050 34996 25052
rect 35020 25050 35076 25052
rect 35100 25050 35156 25052
rect 35180 25050 35236 25052
rect 34940 24998 34966 25050
rect 34966 24998 34996 25050
rect 35020 24998 35030 25050
rect 35030 24998 35076 25050
rect 35100 24998 35146 25050
rect 35146 24998 35156 25050
rect 35180 24998 35210 25050
rect 35210 24998 35236 25050
rect 34940 24996 34996 24998
rect 35020 24996 35076 24998
rect 35100 24996 35156 24998
rect 35180 24996 35236 24998
rect 35898 26152 35954 26208
rect 34940 23962 34996 23964
rect 35020 23962 35076 23964
rect 35100 23962 35156 23964
rect 35180 23962 35236 23964
rect 34940 23910 34966 23962
rect 34966 23910 34996 23962
rect 35020 23910 35030 23962
rect 35030 23910 35076 23962
rect 35100 23910 35146 23962
rect 35146 23910 35156 23962
rect 35180 23910 35210 23962
rect 35210 23910 35236 23962
rect 34940 23908 34996 23910
rect 35020 23908 35076 23910
rect 35100 23908 35156 23910
rect 35180 23908 35236 23910
rect 34940 22874 34996 22876
rect 35020 22874 35076 22876
rect 35100 22874 35156 22876
rect 35180 22874 35236 22876
rect 34940 22822 34966 22874
rect 34966 22822 34996 22874
rect 35020 22822 35030 22874
rect 35030 22822 35076 22874
rect 35100 22822 35146 22874
rect 35146 22822 35156 22874
rect 35180 22822 35210 22874
rect 35210 22822 35236 22874
rect 34940 22820 34996 22822
rect 35020 22820 35076 22822
rect 35100 22820 35156 22822
rect 35180 22820 35236 22822
rect 34940 21786 34996 21788
rect 35020 21786 35076 21788
rect 35100 21786 35156 21788
rect 35180 21786 35236 21788
rect 34940 21734 34966 21786
rect 34966 21734 34996 21786
rect 35020 21734 35030 21786
rect 35030 21734 35076 21786
rect 35100 21734 35146 21786
rect 35146 21734 35156 21786
rect 35180 21734 35210 21786
rect 35210 21734 35236 21786
rect 34940 21732 34996 21734
rect 35020 21732 35076 21734
rect 35100 21732 35156 21734
rect 35180 21732 35236 21734
rect 34940 20698 34996 20700
rect 35020 20698 35076 20700
rect 35100 20698 35156 20700
rect 35180 20698 35236 20700
rect 34940 20646 34966 20698
rect 34966 20646 34996 20698
rect 35020 20646 35030 20698
rect 35030 20646 35076 20698
rect 35100 20646 35146 20698
rect 35146 20646 35156 20698
rect 35180 20646 35210 20698
rect 35210 20646 35236 20698
rect 34940 20644 34996 20646
rect 35020 20644 35076 20646
rect 35100 20644 35156 20646
rect 35180 20644 35236 20646
rect 35898 22888 35954 22944
rect 34940 19610 34996 19612
rect 35020 19610 35076 19612
rect 35100 19610 35156 19612
rect 35180 19610 35236 19612
rect 34940 19558 34966 19610
rect 34966 19558 34996 19610
rect 35020 19558 35030 19610
rect 35030 19558 35076 19610
rect 35100 19558 35146 19610
rect 35146 19558 35156 19610
rect 35180 19558 35210 19610
rect 35210 19558 35236 19610
rect 34940 19556 34996 19558
rect 35020 19556 35076 19558
rect 35100 19556 35156 19558
rect 35180 19556 35236 19558
rect 34518 13368 34574 13424
rect 34426 12688 34482 12744
rect 34940 18522 34996 18524
rect 35020 18522 35076 18524
rect 35100 18522 35156 18524
rect 35180 18522 35236 18524
rect 34940 18470 34966 18522
rect 34966 18470 34996 18522
rect 35020 18470 35030 18522
rect 35030 18470 35076 18522
rect 35100 18470 35146 18522
rect 35146 18470 35156 18522
rect 35180 18470 35210 18522
rect 35210 18470 35236 18522
rect 34940 18468 34996 18470
rect 35020 18468 35076 18470
rect 35100 18468 35156 18470
rect 35180 18468 35236 18470
rect 34940 17434 34996 17436
rect 35020 17434 35076 17436
rect 35100 17434 35156 17436
rect 35180 17434 35236 17436
rect 34940 17382 34966 17434
rect 34966 17382 34996 17434
rect 35020 17382 35030 17434
rect 35030 17382 35076 17434
rect 35100 17382 35146 17434
rect 35146 17382 35156 17434
rect 35180 17382 35210 17434
rect 35210 17382 35236 17434
rect 34940 17380 34996 17382
rect 35020 17380 35076 17382
rect 35100 17380 35156 17382
rect 35180 17380 35236 17382
rect 34978 16788 35034 16824
rect 34978 16768 34980 16788
rect 34980 16768 35032 16788
rect 35032 16768 35034 16788
rect 34940 16346 34996 16348
rect 35020 16346 35076 16348
rect 35100 16346 35156 16348
rect 35180 16346 35236 16348
rect 34940 16294 34966 16346
rect 34966 16294 34996 16346
rect 35020 16294 35030 16346
rect 35030 16294 35076 16346
rect 35100 16294 35146 16346
rect 35146 16294 35156 16346
rect 35180 16294 35210 16346
rect 35210 16294 35236 16346
rect 34940 16292 34996 16294
rect 35020 16292 35076 16294
rect 35100 16292 35156 16294
rect 35180 16292 35236 16294
rect 36174 32408 36230 32464
rect 34940 15258 34996 15260
rect 35020 15258 35076 15260
rect 35100 15258 35156 15260
rect 35180 15258 35236 15260
rect 34940 15206 34966 15258
rect 34966 15206 34996 15258
rect 35020 15206 35030 15258
rect 35030 15206 35076 15258
rect 35100 15206 35146 15258
rect 35146 15206 35156 15258
rect 35180 15206 35210 15258
rect 35210 15206 35236 15258
rect 34940 15204 34996 15206
rect 35020 15204 35076 15206
rect 35100 15204 35156 15206
rect 35180 15204 35236 15206
rect 34940 14170 34996 14172
rect 35020 14170 35076 14172
rect 35100 14170 35156 14172
rect 35180 14170 35236 14172
rect 34940 14118 34966 14170
rect 34966 14118 34996 14170
rect 35020 14118 35030 14170
rect 35030 14118 35076 14170
rect 35100 14118 35146 14170
rect 35146 14118 35156 14170
rect 35180 14118 35210 14170
rect 35210 14118 35236 14170
rect 34940 14116 34996 14118
rect 35020 14116 35076 14118
rect 35100 14116 35156 14118
rect 35180 14116 35236 14118
rect 34940 13082 34996 13084
rect 35020 13082 35076 13084
rect 35100 13082 35156 13084
rect 35180 13082 35236 13084
rect 34940 13030 34966 13082
rect 34966 13030 34996 13082
rect 35020 13030 35030 13082
rect 35030 13030 35076 13082
rect 35100 13030 35146 13082
rect 35146 13030 35156 13082
rect 35180 13030 35210 13082
rect 35210 13030 35236 13082
rect 34940 13028 34996 13030
rect 35020 13028 35076 13030
rect 35100 13028 35156 13030
rect 35180 13028 35236 13030
rect 34794 12688 34850 12744
rect 35714 13232 35770 13288
rect 34940 11994 34996 11996
rect 35020 11994 35076 11996
rect 35100 11994 35156 11996
rect 35180 11994 35236 11996
rect 34940 11942 34966 11994
rect 34966 11942 34996 11994
rect 35020 11942 35030 11994
rect 35030 11942 35076 11994
rect 35100 11942 35146 11994
rect 35146 11942 35156 11994
rect 35180 11942 35210 11994
rect 35210 11942 35236 11994
rect 34940 11940 34996 11942
rect 35020 11940 35076 11942
rect 35100 11940 35156 11942
rect 35180 11940 35236 11942
rect 36266 23604 36268 23624
rect 36268 23604 36320 23624
rect 36320 23604 36322 23624
rect 36266 23568 36322 23604
rect 36726 19896 36782 19952
rect 36174 12824 36230 12880
rect 35438 11056 35494 11112
rect 34940 10906 34996 10908
rect 35020 10906 35076 10908
rect 35100 10906 35156 10908
rect 35180 10906 35236 10908
rect 34940 10854 34966 10906
rect 34966 10854 34996 10906
rect 35020 10854 35030 10906
rect 35030 10854 35076 10906
rect 35100 10854 35146 10906
rect 35146 10854 35156 10906
rect 35180 10854 35210 10906
rect 35210 10854 35236 10906
rect 34940 10852 34996 10854
rect 35020 10852 35076 10854
rect 35100 10852 35156 10854
rect 35180 10852 35236 10854
rect 34940 9818 34996 9820
rect 35020 9818 35076 9820
rect 35100 9818 35156 9820
rect 35180 9818 35236 9820
rect 34940 9766 34966 9818
rect 34966 9766 34996 9818
rect 35020 9766 35030 9818
rect 35030 9766 35076 9818
rect 35100 9766 35146 9818
rect 35146 9766 35156 9818
rect 35180 9766 35210 9818
rect 35210 9766 35236 9818
rect 34940 9764 34996 9766
rect 35020 9764 35076 9766
rect 35100 9764 35156 9766
rect 35180 9764 35236 9766
rect 34940 8730 34996 8732
rect 35020 8730 35076 8732
rect 35100 8730 35156 8732
rect 35180 8730 35236 8732
rect 34940 8678 34966 8730
rect 34966 8678 34996 8730
rect 35020 8678 35030 8730
rect 35030 8678 35076 8730
rect 35100 8678 35146 8730
rect 35146 8678 35156 8730
rect 35180 8678 35210 8730
rect 35210 8678 35236 8730
rect 34940 8676 34996 8678
rect 35020 8676 35076 8678
rect 35100 8676 35156 8678
rect 35180 8676 35236 8678
rect 34940 7642 34996 7644
rect 35020 7642 35076 7644
rect 35100 7642 35156 7644
rect 35180 7642 35236 7644
rect 34940 7590 34966 7642
rect 34966 7590 34996 7642
rect 35020 7590 35030 7642
rect 35030 7590 35076 7642
rect 35100 7590 35146 7642
rect 35146 7590 35156 7642
rect 35180 7590 35210 7642
rect 35210 7590 35236 7642
rect 34940 7588 34996 7590
rect 35020 7588 35076 7590
rect 35100 7588 35156 7590
rect 35180 7588 35236 7590
rect 34940 6554 34996 6556
rect 35020 6554 35076 6556
rect 35100 6554 35156 6556
rect 35180 6554 35236 6556
rect 34940 6502 34966 6554
rect 34966 6502 34996 6554
rect 35020 6502 35030 6554
rect 35030 6502 35076 6554
rect 35100 6502 35146 6554
rect 35146 6502 35156 6554
rect 35180 6502 35210 6554
rect 35210 6502 35236 6554
rect 34940 6500 34996 6502
rect 35020 6500 35076 6502
rect 35100 6500 35156 6502
rect 35180 6500 35236 6502
rect 35898 10376 35954 10432
rect 37002 16632 37058 16688
rect 37002 13640 37058 13696
rect 34940 5466 34996 5468
rect 35020 5466 35076 5468
rect 35100 5466 35156 5468
rect 35180 5466 35236 5468
rect 34940 5414 34966 5466
rect 34966 5414 34996 5466
rect 35020 5414 35030 5466
rect 35030 5414 35076 5466
rect 35100 5414 35146 5466
rect 35146 5414 35156 5466
rect 35180 5414 35210 5466
rect 35210 5414 35236 5466
rect 34940 5412 34996 5414
rect 35020 5412 35076 5414
rect 35100 5412 35156 5414
rect 35180 5412 35236 5414
rect 34940 4378 34996 4380
rect 35020 4378 35076 4380
rect 35100 4378 35156 4380
rect 35180 4378 35236 4380
rect 34940 4326 34966 4378
rect 34966 4326 34996 4378
rect 35020 4326 35030 4378
rect 35030 4326 35076 4378
rect 35100 4326 35146 4378
rect 35146 4326 35156 4378
rect 35180 4326 35210 4378
rect 35210 4326 35236 4378
rect 34940 4324 34996 4326
rect 35020 4324 35076 4326
rect 35100 4324 35156 4326
rect 35180 4324 35236 4326
rect 35898 4120 35954 4176
rect 36726 10648 36782 10704
rect 36726 7404 36782 7440
rect 36726 7384 36728 7404
rect 36728 7384 36780 7404
rect 36780 7384 36782 7404
rect 37186 11620 37242 11656
rect 37186 11600 37188 11620
rect 37188 11600 37240 11620
rect 37240 11600 37242 11620
rect 38934 29144 38990 29200
rect 38198 23180 38254 23216
rect 38198 23160 38200 23180
rect 38200 23160 38252 23180
rect 38252 23160 38254 23180
rect 37830 22092 37886 22128
rect 37830 22072 37832 22092
rect 37832 22072 37884 22092
rect 37884 22072 37886 22092
rect 38566 10648 38622 10704
rect 34940 3290 34996 3292
rect 35020 3290 35076 3292
rect 35100 3290 35156 3292
rect 35180 3290 35236 3292
rect 34940 3238 34966 3290
rect 34966 3238 34996 3290
rect 35020 3238 35030 3290
rect 35030 3238 35076 3290
rect 35100 3238 35146 3290
rect 35146 3238 35156 3290
rect 35180 3238 35210 3290
rect 35210 3238 35236 3290
rect 34940 3236 34996 3238
rect 35020 3236 35076 3238
rect 35100 3236 35156 3238
rect 35180 3236 35236 3238
rect 34940 2202 34996 2204
rect 35020 2202 35076 2204
rect 35100 2202 35156 2204
rect 35180 2202 35236 2204
rect 34940 2150 34966 2202
rect 34966 2150 34996 2202
rect 35020 2150 35030 2202
rect 35030 2150 35076 2202
rect 35100 2150 35146 2202
rect 35146 2150 35156 2202
rect 35180 2150 35210 2202
rect 35210 2150 35236 2202
rect 34940 2148 34996 2150
rect 35020 2148 35076 2150
rect 35100 2148 35156 2150
rect 35180 2148 35236 2150
rect 36450 1128 36506 1184
<< metal3 >>
rect 36077 38722 36143 38725
rect 40200 38722 41000 38752
rect 36077 38720 41000 38722
rect 36077 38664 36082 38720
rect 36138 38664 41000 38720
rect 36077 38662 41000 38664
rect 36077 38659 36143 38662
rect 19568 38656 19888 38657
rect 19568 38592 19576 38656
rect 19640 38592 19656 38656
rect 19720 38592 19736 38656
rect 19800 38592 19816 38656
rect 19880 38592 19888 38656
rect 40200 38632 41000 38662
rect 19568 38591 19888 38592
rect 9673 38450 9739 38453
rect 19149 38450 19215 38453
rect 9673 38448 19215 38450
rect 9673 38392 9678 38448
rect 9734 38392 19154 38448
rect 19210 38392 19215 38448
rect 9673 38390 19215 38392
rect 9673 38387 9739 38390
rect 19149 38387 19215 38390
rect 0 38178 800 38208
rect 1853 38178 1919 38181
rect 0 38176 1919 38178
rect 0 38120 1858 38176
rect 1914 38120 1919 38176
rect 0 38118 1919 38120
rect 0 38088 800 38118
rect 1853 38115 1919 38118
rect 4208 38112 4528 38113
rect 4208 38048 4216 38112
rect 4280 38048 4296 38112
rect 4360 38048 4376 38112
rect 4440 38048 4456 38112
rect 4520 38048 4528 38112
rect 4208 38047 4528 38048
rect 34928 38112 35248 38113
rect 34928 38048 34936 38112
rect 35000 38048 35016 38112
rect 35080 38048 35096 38112
rect 35160 38048 35176 38112
rect 35240 38048 35248 38112
rect 34928 38047 35248 38048
rect 19568 37568 19888 37569
rect 19568 37504 19576 37568
rect 19640 37504 19656 37568
rect 19720 37504 19736 37568
rect 19800 37504 19816 37568
rect 19880 37504 19888 37568
rect 19568 37503 19888 37504
rect 4208 37024 4528 37025
rect 4208 36960 4216 37024
rect 4280 36960 4296 37024
rect 4360 36960 4376 37024
rect 4440 36960 4456 37024
rect 4520 36960 4528 37024
rect 4208 36959 4528 36960
rect 34928 37024 35248 37025
rect 34928 36960 34936 37024
rect 35000 36960 35016 37024
rect 35080 36960 35096 37024
rect 35160 36960 35176 37024
rect 35240 36960 35248 37024
rect 34928 36959 35248 36960
rect 19568 36480 19888 36481
rect 19568 36416 19576 36480
rect 19640 36416 19656 36480
rect 19720 36416 19736 36480
rect 19800 36416 19816 36480
rect 19880 36416 19888 36480
rect 19568 36415 19888 36416
rect 4208 35936 4528 35937
rect 4208 35872 4216 35936
rect 4280 35872 4296 35936
rect 4360 35872 4376 35936
rect 4440 35872 4456 35936
rect 4520 35872 4528 35936
rect 4208 35871 4528 35872
rect 34928 35936 35248 35937
rect 34928 35872 34936 35936
rect 35000 35872 35016 35936
rect 35080 35872 35096 35936
rect 35160 35872 35176 35936
rect 35240 35872 35248 35936
rect 34928 35871 35248 35872
rect 35985 35458 36051 35461
rect 40200 35458 41000 35488
rect 35985 35456 41000 35458
rect 35985 35400 35990 35456
rect 36046 35400 41000 35456
rect 35985 35398 41000 35400
rect 35985 35395 36051 35398
rect 19568 35392 19888 35393
rect 19568 35328 19576 35392
rect 19640 35328 19656 35392
rect 19720 35328 19736 35392
rect 19800 35328 19816 35392
rect 19880 35328 19888 35392
rect 40200 35368 41000 35398
rect 19568 35327 19888 35328
rect 0 35186 800 35216
rect 3601 35186 3667 35189
rect 0 35184 3667 35186
rect 0 35128 3606 35184
rect 3662 35128 3667 35184
rect 0 35126 3667 35128
rect 0 35096 800 35126
rect 3601 35123 3667 35126
rect 4208 34848 4528 34849
rect 4208 34784 4216 34848
rect 4280 34784 4296 34848
rect 4360 34784 4376 34848
rect 4440 34784 4456 34848
rect 4520 34784 4528 34848
rect 4208 34783 4528 34784
rect 34928 34848 35248 34849
rect 34928 34784 34936 34848
rect 35000 34784 35016 34848
rect 35080 34784 35096 34848
rect 35160 34784 35176 34848
rect 35240 34784 35248 34848
rect 34928 34783 35248 34784
rect 19568 34304 19888 34305
rect 19568 34240 19576 34304
rect 19640 34240 19656 34304
rect 19720 34240 19736 34304
rect 19800 34240 19816 34304
rect 19880 34240 19888 34304
rect 19568 34239 19888 34240
rect 4208 33760 4528 33761
rect 4208 33696 4216 33760
rect 4280 33696 4296 33760
rect 4360 33696 4376 33760
rect 4440 33696 4456 33760
rect 4520 33696 4528 33760
rect 4208 33695 4528 33696
rect 34928 33760 35248 33761
rect 34928 33696 34936 33760
rect 35000 33696 35016 33760
rect 35080 33696 35096 33760
rect 35160 33696 35176 33760
rect 35240 33696 35248 33760
rect 34928 33695 35248 33696
rect 19568 33216 19888 33217
rect 19568 33152 19576 33216
rect 19640 33152 19656 33216
rect 19720 33152 19736 33216
rect 19800 33152 19816 33216
rect 19880 33152 19888 33216
rect 19568 33151 19888 33152
rect 4208 32672 4528 32673
rect 4208 32608 4216 32672
rect 4280 32608 4296 32672
rect 4360 32608 4376 32672
rect 4440 32608 4456 32672
rect 4520 32608 4528 32672
rect 4208 32607 4528 32608
rect 34928 32672 35248 32673
rect 34928 32608 34936 32672
rect 35000 32608 35016 32672
rect 35080 32608 35096 32672
rect 35160 32608 35176 32672
rect 35240 32608 35248 32672
rect 34928 32607 35248 32608
rect 36169 32466 36235 32469
rect 40200 32466 41000 32496
rect 36169 32464 41000 32466
rect 36169 32408 36174 32464
rect 36230 32408 41000 32464
rect 36169 32406 41000 32408
rect 36169 32403 36235 32406
rect 40200 32376 41000 32406
rect 19568 32128 19888 32129
rect 19568 32064 19576 32128
rect 19640 32064 19656 32128
rect 19720 32064 19736 32128
rect 19800 32064 19816 32128
rect 19880 32064 19888 32128
rect 19568 32063 19888 32064
rect 0 31922 800 31952
rect 2865 31922 2931 31925
rect 0 31920 2931 31922
rect 0 31864 2870 31920
rect 2926 31864 2931 31920
rect 0 31862 2931 31864
rect 0 31832 800 31862
rect 2865 31859 2931 31862
rect 4208 31584 4528 31585
rect 4208 31520 4216 31584
rect 4280 31520 4296 31584
rect 4360 31520 4376 31584
rect 4440 31520 4456 31584
rect 4520 31520 4528 31584
rect 4208 31519 4528 31520
rect 34928 31584 35248 31585
rect 34928 31520 34936 31584
rect 35000 31520 35016 31584
rect 35080 31520 35096 31584
rect 35160 31520 35176 31584
rect 35240 31520 35248 31584
rect 34928 31519 35248 31520
rect 19568 31040 19888 31041
rect 19568 30976 19576 31040
rect 19640 30976 19656 31040
rect 19720 30976 19736 31040
rect 19800 30976 19816 31040
rect 19880 30976 19888 31040
rect 19568 30975 19888 30976
rect 4208 30496 4528 30497
rect 4208 30432 4216 30496
rect 4280 30432 4296 30496
rect 4360 30432 4376 30496
rect 4440 30432 4456 30496
rect 4520 30432 4528 30496
rect 4208 30431 4528 30432
rect 34928 30496 35248 30497
rect 34928 30432 34936 30496
rect 35000 30432 35016 30496
rect 35080 30432 35096 30496
rect 35160 30432 35176 30496
rect 35240 30432 35248 30496
rect 34928 30431 35248 30432
rect 9581 30154 9647 30157
rect 15837 30154 15903 30157
rect 9581 30152 15903 30154
rect 9581 30096 9586 30152
rect 9642 30096 15842 30152
rect 15898 30096 15903 30152
rect 9581 30094 15903 30096
rect 9581 30091 9647 30094
rect 15837 30091 15903 30094
rect 19568 29952 19888 29953
rect 19568 29888 19576 29952
rect 19640 29888 19656 29952
rect 19720 29888 19736 29952
rect 19800 29888 19816 29952
rect 19880 29888 19888 29952
rect 19568 29887 19888 29888
rect 4208 29408 4528 29409
rect 4208 29344 4216 29408
rect 4280 29344 4296 29408
rect 4360 29344 4376 29408
rect 4440 29344 4456 29408
rect 4520 29344 4528 29408
rect 4208 29343 4528 29344
rect 34928 29408 35248 29409
rect 34928 29344 34936 29408
rect 35000 29344 35016 29408
rect 35080 29344 35096 29408
rect 35160 29344 35176 29408
rect 35240 29344 35248 29408
rect 34928 29343 35248 29344
rect 38929 29202 38995 29205
rect 40200 29202 41000 29232
rect 38929 29200 41000 29202
rect 38929 29144 38934 29200
rect 38990 29144 41000 29200
rect 38929 29142 41000 29144
rect 38929 29139 38995 29142
rect 40200 29112 41000 29142
rect 18597 29066 18663 29069
rect 18597 29064 18706 29066
rect 18597 29008 18602 29064
rect 18658 29008 18706 29064
rect 18597 29003 18706 29008
rect 0 28930 800 28960
rect 3049 28930 3115 28933
rect 0 28928 3115 28930
rect 0 28872 3054 28928
rect 3110 28872 3115 28928
rect 0 28870 3115 28872
rect 0 28840 800 28870
rect 3049 28867 3115 28870
rect 18505 28522 18571 28525
rect 18646 28522 18706 29003
rect 18873 28932 18939 28933
rect 18822 28868 18828 28932
rect 18892 28930 18939 28932
rect 18892 28928 18984 28930
rect 18934 28872 18984 28928
rect 18892 28870 18984 28872
rect 18892 28868 18939 28870
rect 18873 28867 18939 28868
rect 19568 28864 19888 28865
rect 19568 28800 19576 28864
rect 19640 28800 19656 28864
rect 19720 28800 19736 28864
rect 19800 28800 19816 28864
rect 19880 28800 19888 28864
rect 19568 28799 19888 28800
rect 18505 28520 18706 28522
rect 18505 28464 18510 28520
rect 18566 28464 18706 28520
rect 18505 28462 18706 28464
rect 18505 28459 18571 28462
rect 4208 28320 4528 28321
rect 4208 28256 4216 28320
rect 4280 28256 4296 28320
rect 4360 28256 4376 28320
rect 4440 28256 4456 28320
rect 4520 28256 4528 28320
rect 4208 28255 4528 28256
rect 34928 28320 35248 28321
rect 34928 28256 34936 28320
rect 35000 28256 35016 28320
rect 35080 28256 35096 28320
rect 35160 28256 35176 28320
rect 35240 28256 35248 28320
rect 34928 28255 35248 28256
rect 19568 27776 19888 27777
rect 19568 27712 19576 27776
rect 19640 27712 19656 27776
rect 19720 27712 19736 27776
rect 19800 27712 19816 27776
rect 19880 27712 19888 27776
rect 19568 27711 19888 27712
rect 4208 27232 4528 27233
rect 4208 27168 4216 27232
rect 4280 27168 4296 27232
rect 4360 27168 4376 27232
rect 4440 27168 4456 27232
rect 4520 27168 4528 27232
rect 4208 27167 4528 27168
rect 34928 27232 35248 27233
rect 34928 27168 34936 27232
rect 35000 27168 35016 27232
rect 35080 27168 35096 27232
rect 35160 27168 35176 27232
rect 35240 27168 35248 27232
rect 34928 27167 35248 27168
rect 19568 26688 19888 26689
rect 19568 26624 19576 26688
rect 19640 26624 19656 26688
rect 19720 26624 19736 26688
rect 19800 26624 19816 26688
rect 19880 26624 19888 26688
rect 19568 26623 19888 26624
rect 35893 26210 35959 26213
rect 40200 26210 41000 26240
rect 35893 26208 41000 26210
rect 35893 26152 35898 26208
rect 35954 26152 41000 26208
rect 35893 26150 41000 26152
rect 35893 26147 35959 26150
rect 4208 26144 4528 26145
rect 4208 26080 4216 26144
rect 4280 26080 4296 26144
rect 4360 26080 4376 26144
rect 4440 26080 4456 26144
rect 4520 26080 4528 26144
rect 4208 26079 4528 26080
rect 34928 26144 35248 26145
rect 34928 26080 34936 26144
rect 35000 26080 35016 26144
rect 35080 26080 35096 26144
rect 35160 26080 35176 26144
rect 35240 26080 35248 26144
rect 40200 26120 41000 26150
rect 34928 26079 35248 26080
rect 0 25666 800 25696
rect 3969 25666 4035 25669
rect 0 25664 4035 25666
rect 0 25608 3974 25664
rect 4030 25608 4035 25664
rect 0 25606 4035 25608
rect 0 25576 800 25606
rect 3969 25603 4035 25606
rect 19568 25600 19888 25601
rect 19568 25536 19576 25600
rect 19640 25536 19656 25600
rect 19720 25536 19736 25600
rect 19800 25536 19816 25600
rect 19880 25536 19888 25600
rect 19568 25535 19888 25536
rect 4208 25056 4528 25057
rect 4208 24992 4216 25056
rect 4280 24992 4296 25056
rect 4360 24992 4376 25056
rect 4440 24992 4456 25056
rect 4520 24992 4528 25056
rect 4208 24991 4528 24992
rect 34928 25056 35248 25057
rect 34928 24992 34936 25056
rect 35000 24992 35016 25056
rect 35080 24992 35096 25056
rect 35160 24992 35176 25056
rect 35240 24992 35248 25056
rect 34928 24991 35248 24992
rect 19568 24512 19888 24513
rect 19568 24448 19576 24512
rect 19640 24448 19656 24512
rect 19720 24448 19736 24512
rect 19800 24448 19816 24512
rect 19880 24448 19888 24512
rect 19568 24447 19888 24448
rect 12985 24306 13051 24309
rect 18505 24306 18571 24309
rect 12985 24304 18571 24306
rect 12985 24248 12990 24304
rect 13046 24248 18510 24304
rect 18566 24248 18571 24304
rect 12985 24246 18571 24248
rect 12985 24243 13051 24246
rect 18505 24243 18571 24246
rect 4208 23968 4528 23969
rect 4208 23904 4216 23968
rect 4280 23904 4296 23968
rect 4360 23904 4376 23968
rect 4440 23904 4456 23968
rect 4520 23904 4528 23968
rect 4208 23903 4528 23904
rect 34928 23968 35248 23969
rect 34928 23904 34936 23968
rect 35000 23904 35016 23968
rect 35080 23904 35096 23968
rect 35160 23904 35176 23968
rect 35240 23904 35248 23968
rect 34928 23903 35248 23904
rect 29269 23626 29335 23629
rect 36261 23626 36327 23629
rect 29269 23624 36327 23626
rect 29269 23568 29274 23624
rect 29330 23568 36266 23624
rect 36322 23568 36327 23624
rect 29269 23566 36327 23568
rect 29269 23563 29335 23566
rect 36261 23563 36327 23566
rect 19568 23424 19888 23425
rect 19568 23360 19576 23424
rect 19640 23360 19656 23424
rect 19720 23360 19736 23424
rect 19800 23360 19816 23424
rect 19880 23360 19888 23424
rect 19568 23359 19888 23360
rect 12157 23354 12223 23357
rect 18873 23354 18939 23357
rect 12157 23352 18939 23354
rect 12157 23296 12162 23352
rect 12218 23296 18878 23352
rect 18934 23296 18939 23352
rect 12157 23294 18939 23296
rect 12157 23291 12223 23294
rect 18873 23291 18939 23294
rect 18873 23220 18939 23221
rect 18822 23156 18828 23220
rect 18892 23218 18939 23220
rect 33317 23218 33383 23221
rect 38193 23218 38259 23221
rect 18892 23216 18984 23218
rect 18934 23160 18984 23216
rect 18892 23158 18984 23160
rect 33317 23216 38259 23218
rect 33317 23160 33322 23216
rect 33378 23160 38198 23216
rect 38254 23160 38259 23216
rect 33317 23158 38259 23160
rect 18892 23156 18939 23158
rect 18873 23155 18939 23156
rect 33317 23155 33383 23158
rect 38193 23155 38259 23158
rect 35893 22946 35959 22949
rect 40200 22946 41000 22976
rect 35893 22944 41000 22946
rect 35893 22888 35898 22944
rect 35954 22888 41000 22944
rect 35893 22886 41000 22888
rect 35893 22883 35959 22886
rect 4208 22880 4528 22881
rect 4208 22816 4216 22880
rect 4280 22816 4296 22880
rect 4360 22816 4376 22880
rect 4440 22816 4456 22880
rect 4520 22816 4528 22880
rect 4208 22815 4528 22816
rect 34928 22880 35248 22881
rect 34928 22816 34936 22880
rect 35000 22816 35016 22880
rect 35080 22816 35096 22880
rect 35160 22816 35176 22880
rect 35240 22816 35248 22880
rect 40200 22856 41000 22886
rect 34928 22815 35248 22816
rect 0 22674 800 22704
rect 1577 22674 1643 22677
rect 0 22672 1643 22674
rect 0 22616 1582 22672
rect 1638 22616 1643 22672
rect 0 22614 1643 22616
rect 0 22584 800 22614
rect 1577 22611 1643 22614
rect 19568 22336 19888 22337
rect 19568 22272 19576 22336
rect 19640 22272 19656 22336
rect 19720 22272 19736 22336
rect 19800 22272 19816 22336
rect 19880 22272 19888 22336
rect 19568 22271 19888 22272
rect 31109 22130 31175 22133
rect 37825 22130 37891 22133
rect 31109 22128 37891 22130
rect 31109 22072 31114 22128
rect 31170 22072 37830 22128
rect 37886 22072 37891 22128
rect 31109 22070 37891 22072
rect 31109 22067 31175 22070
rect 37825 22067 37891 22070
rect 29085 21994 29151 21997
rect 30833 21994 30899 21997
rect 29085 21992 30899 21994
rect 29085 21936 29090 21992
rect 29146 21936 30838 21992
rect 30894 21936 30899 21992
rect 29085 21934 30899 21936
rect 29085 21931 29151 21934
rect 30833 21931 30899 21934
rect 4208 21792 4528 21793
rect 4208 21728 4216 21792
rect 4280 21728 4296 21792
rect 4360 21728 4376 21792
rect 4440 21728 4456 21792
rect 4520 21728 4528 21792
rect 4208 21727 4528 21728
rect 34928 21792 35248 21793
rect 34928 21728 34936 21792
rect 35000 21728 35016 21792
rect 35080 21728 35096 21792
rect 35160 21728 35176 21792
rect 35240 21728 35248 21792
rect 34928 21727 35248 21728
rect 19885 21586 19951 21589
rect 20069 21586 20135 21589
rect 19885 21584 20135 21586
rect 19885 21528 19890 21584
rect 19946 21528 20074 21584
rect 20130 21528 20135 21584
rect 19885 21526 20135 21528
rect 19885 21523 19951 21526
rect 20069 21523 20135 21526
rect 19568 21248 19888 21249
rect 19568 21184 19576 21248
rect 19640 21184 19656 21248
rect 19720 21184 19736 21248
rect 19800 21184 19816 21248
rect 19880 21184 19888 21248
rect 19568 21183 19888 21184
rect 4208 20704 4528 20705
rect 4208 20640 4216 20704
rect 4280 20640 4296 20704
rect 4360 20640 4376 20704
rect 4440 20640 4456 20704
rect 4520 20640 4528 20704
rect 4208 20639 4528 20640
rect 34928 20704 35248 20705
rect 34928 20640 34936 20704
rect 35000 20640 35016 20704
rect 35080 20640 35096 20704
rect 35160 20640 35176 20704
rect 35240 20640 35248 20704
rect 34928 20639 35248 20640
rect 5901 20362 5967 20365
rect 8017 20362 8083 20365
rect 5901 20360 8083 20362
rect 5901 20304 5906 20360
rect 5962 20304 8022 20360
rect 8078 20304 8083 20360
rect 5901 20302 8083 20304
rect 5901 20299 5967 20302
rect 8017 20299 8083 20302
rect 13813 20226 13879 20229
rect 17585 20226 17651 20229
rect 13813 20224 17651 20226
rect 13813 20168 13818 20224
rect 13874 20168 17590 20224
rect 17646 20168 17651 20224
rect 13813 20166 17651 20168
rect 13813 20163 13879 20166
rect 17585 20163 17651 20166
rect 19568 20160 19888 20161
rect 19568 20096 19576 20160
rect 19640 20096 19656 20160
rect 19720 20096 19736 20160
rect 19800 20096 19816 20160
rect 19880 20096 19888 20160
rect 19568 20095 19888 20096
rect 10409 19954 10475 19957
rect 18413 19954 18479 19957
rect 10409 19952 18479 19954
rect 10409 19896 10414 19952
rect 10470 19896 18418 19952
rect 18474 19896 18479 19952
rect 10409 19894 18479 19896
rect 10409 19891 10475 19894
rect 18413 19891 18479 19894
rect 23013 19954 23079 19957
rect 27429 19954 27495 19957
rect 23013 19952 27495 19954
rect 23013 19896 23018 19952
rect 23074 19896 27434 19952
rect 27490 19896 27495 19952
rect 23013 19894 27495 19896
rect 23013 19891 23079 19894
rect 27429 19891 27495 19894
rect 36721 19954 36787 19957
rect 40200 19954 41000 19984
rect 36721 19952 41000 19954
rect 36721 19896 36726 19952
rect 36782 19896 41000 19952
rect 36721 19894 41000 19896
rect 36721 19891 36787 19894
rect 40200 19864 41000 19894
rect 4208 19616 4528 19617
rect 4208 19552 4216 19616
rect 4280 19552 4296 19616
rect 4360 19552 4376 19616
rect 4440 19552 4456 19616
rect 4520 19552 4528 19616
rect 4208 19551 4528 19552
rect 34928 19616 35248 19617
rect 34928 19552 34936 19616
rect 35000 19552 35016 19616
rect 35080 19552 35096 19616
rect 35160 19552 35176 19616
rect 35240 19552 35248 19616
rect 34928 19551 35248 19552
rect 0 19410 800 19440
rect 4061 19410 4127 19413
rect 0 19408 4127 19410
rect 0 19352 4066 19408
rect 4122 19352 4127 19408
rect 0 19350 4127 19352
rect 0 19320 800 19350
rect 4061 19347 4127 19350
rect 2773 19274 2839 19277
rect 3693 19274 3759 19277
rect 2773 19272 3759 19274
rect 2773 19216 2778 19272
rect 2834 19216 3698 19272
rect 3754 19216 3759 19272
rect 2773 19214 3759 19216
rect 2773 19211 2839 19214
rect 3693 19211 3759 19214
rect 16665 19274 16731 19277
rect 17585 19274 17651 19277
rect 25037 19274 25103 19277
rect 16665 19272 25103 19274
rect 16665 19216 16670 19272
rect 16726 19216 17590 19272
rect 17646 19216 25042 19272
rect 25098 19216 25103 19272
rect 16665 19214 25103 19216
rect 16665 19211 16731 19214
rect 17585 19211 17651 19214
rect 25037 19211 25103 19214
rect 19568 19072 19888 19073
rect 19568 19008 19576 19072
rect 19640 19008 19656 19072
rect 19720 19008 19736 19072
rect 19800 19008 19816 19072
rect 19880 19008 19888 19072
rect 19568 19007 19888 19008
rect 9765 18730 9831 18733
rect 16757 18730 16823 18733
rect 9765 18728 16823 18730
rect 9765 18672 9770 18728
rect 9826 18672 16762 18728
rect 16818 18672 16823 18728
rect 9765 18670 16823 18672
rect 9765 18667 9831 18670
rect 16757 18667 16823 18670
rect 4208 18528 4528 18529
rect 4208 18464 4216 18528
rect 4280 18464 4296 18528
rect 4360 18464 4376 18528
rect 4440 18464 4456 18528
rect 4520 18464 4528 18528
rect 4208 18463 4528 18464
rect 34928 18528 35248 18529
rect 34928 18464 34936 18528
rect 35000 18464 35016 18528
rect 35080 18464 35096 18528
rect 35160 18464 35176 18528
rect 35240 18464 35248 18528
rect 34928 18463 35248 18464
rect 19568 17984 19888 17985
rect 19568 17920 19576 17984
rect 19640 17920 19656 17984
rect 19720 17920 19736 17984
rect 19800 17920 19816 17984
rect 19880 17920 19888 17984
rect 19568 17919 19888 17920
rect 6085 17778 6151 17781
rect 7097 17778 7163 17781
rect 6085 17776 7163 17778
rect 6085 17720 6090 17776
rect 6146 17720 7102 17776
rect 7158 17720 7163 17776
rect 6085 17718 7163 17720
rect 6085 17715 6151 17718
rect 7097 17715 7163 17718
rect 4208 17440 4528 17441
rect 4208 17376 4216 17440
rect 4280 17376 4296 17440
rect 4360 17376 4376 17440
rect 4440 17376 4456 17440
rect 4520 17376 4528 17440
rect 4208 17375 4528 17376
rect 34928 17440 35248 17441
rect 34928 17376 34936 17440
rect 35000 17376 35016 17440
rect 35080 17376 35096 17440
rect 35160 17376 35176 17440
rect 35240 17376 35248 17440
rect 34928 17375 35248 17376
rect 26141 17098 26207 17101
rect 28073 17098 28139 17101
rect 26141 17096 28139 17098
rect 26141 17040 26146 17096
rect 26202 17040 28078 17096
rect 28134 17040 28139 17096
rect 26141 17038 28139 17040
rect 26141 17035 26207 17038
rect 28073 17035 28139 17038
rect 19568 16896 19888 16897
rect 19568 16832 19576 16896
rect 19640 16832 19656 16896
rect 19720 16832 19736 16896
rect 19800 16832 19816 16896
rect 19880 16832 19888 16896
rect 19568 16831 19888 16832
rect 26233 16826 26299 16829
rect 28901 16826 28967 16829
rect 26233 16824 28967 16826
rect 26233 16768 26238 16824
rect 26294 16768 28906 16824
rect 28962 16768 28967 16824
rect 26233 16766 28967 16768
rect 26233 16763 26299 16766
rect 28901 16763 28967 16766
rect 29913 16826 29979 16829
rect 34973 16826 35039 16829
rect 29913 16824 35039 16826
rect 29913 16768 29918 16824
rect 29974 16768 34978 16824
rect 35034 16768 35039 16824
rect 29913 16766 35039 16768
rect 29913 16763 29979 16766
rect 34973 16763 35039 16766
rect 3325 16690 3391 16693
rect 4429 16690 4495 16693
rect 3325 16688 4495 16690
rect 3325 16632 3330 16688
rect 3386 16632 4434 16688
rect 4490 16632 4495 16688
rect 3325 16630 4495 16632
rect 3325 16627 3391 16630
rect 4429 16627 4495 16630
rect 25313 16690 25379 16693
rect 33869 16690 33935 16693
rect 25313 16688 33935 16690
rect 25313 16632 25318 16688
rect 25374 16632 33874 16688
rect 33930 16632 33935 16688
rect 25313 16630 33935 16632
rect 25313 16627 25379 16630
rect 33869 16627 33935 16630
rect 36997 16690 37063 16693
rect 40200 16690 41000 16720
rect 36997 16688 41000 16690
rect 36997 16632 37002 16688
rect 37058 16632 41000 16688
rect 36997 16630 41000 16632
rect 36997 16627 37063 16630
rect 40200 16600 41000 16630
rect 21449 16554 21515 16557
rect 24669 16554 24735 16557
rect 21449 16552 24735 16554
rect 21449 16496 21454 16552
rect 21510 16496 24674 16552
rect 24730 16496 24735 16552
rect 21449 16494 24735 16496
rect 21449 16491 21515 16494
rect 24669 16491 24735 16494
rect 0 16418 800 16448
rect 4061 16418 4127 16421
rect 0 16416 4127 16418
rect 0 16360 4066 16416
rect 4122 16360 4127 16416
rect 0 16358 4127 16360
rect 0 16328 800 16358
rect 4061 16355 4127 16358
rect 4208 16352 4528 16353
rect 4208 16288 4216 16352
rect 4280 16288 4296 16352
rect 4360 16288 4376 16352
rect 4440 16288 4456 16352
rect 4520 16288 4528 16352
rect 4208 16287 4528 16288
rect 34928 16352 35248 16353
rect 34928 16288 34936 16352
rect 35000 16288 35016 16352
rect 35080 16288 35096 16352
rect 35160 16288 35176 16352
rect 35240 16288 35248 16352
rect 34928 16287 35248 16288
rect 27337 16146 27403 16149
rect 28349 16146 28415 16149
rect 27337 16144 28415 16146
rect 27337 16088 27342 16144
rect 27398 16088 28354 16144
rect 28410 16088 28415 16144
rect 27337 16086 28415 16088
rect 27337 16083 27403 16086
rect 28349 16083 28415 16086
rect 19977 16010 20043 16013
rect 25497 16010 25563 16013
rect 19977 16008 25563 16010
rect 19977 15952 19982 16008
rect 20038 15952 25502 16008
rect 25558 15952 25563 16008
rect 19977 15950 25563 15952
rect 19977 15947 20043 15950
rect 25497 15947 25563 15950
rect 19568 15808 19888 15809
rect 19568 15744 19576 15808
rect 19640 15744 19656 15808
rect 19720 15744 19736 15808
rect 19800 15744 19816 15808
rect 19880 15744 19888 15808
rect 19568 15743 19888 15744
rect 11697 15466 11763 15469
rect 18137 15466 18203 15469
rect 11697 15464 18203 15466
rect 11697 15408 11702 15464
rect 11758 15408 18142 15464
rect 18198 15408 18203 15464
rect 11697 15406 18203 15408
rect 11697 15403 11763 15406
rect 18137 15403 18203 15406
rect 4208 15264 4528 15265
rect 4208 15200 4216 15264
rect 4280 15200 4296 15264
rect 4360 15200 4376 15264
rect 4440 15200 4456 15264
rect 4520 15200 4528 15264
rect 4208 15199 4528 15200
rect 34928 15264 35248 15265
rect 34928 15200 34936 15264
rect 35000 15200 35016 15264
rect 35080 15200 35096 15264
rect 35160 15200 35176 15264
rect 35240 15200 35248 15264
rect 34928 15199 35248 15200
rect 12617 15058 12683 15061
rect 17125 15058 17191 15061
rect 12617 15056 17191 15058
rect 12617 15000 12622 15056
rect 12678 15000 17130 15056
rect 17186 15000 17191 15056
rect 12617 14998 17191 15000
rect 12617 14995 12683 14998
rect 17125 14995 17191 14998
rect 2497 14786 2563 14789
rect 8937 14786 9003 14789
rect 2497 14784 9003 14786
rect 2497 14728 2502 14784
rect 2558 14728 8942 14784
rect 8998 14728 9003 14784
rect 2497 14726 9003 14728
rect 2497 14723 2563 14726
rect 8937 14723 9003 14726
rect 10317 14786 10383 14789
rect 11697 14786 11763 14789
rect 19149 14786 19215 14789
rect 10317 14784 19215 14786
rect 10317 14728 10322 14784
rect 10378 14728 11702 14784
rect 11758 14728 19154 14784
rect 19210 14728 19215 14784
rect 10317 14726 19215 14728
rect 10317 14723 10383 14726
rect 11697 14723 11763 14726
rect 19149 14723 19215 14726
rect 19568 14720 19888 14721
rect 19568 14656 19576 14720
rect 19640 14656 19656 14720
rect 19720 14656 19736 14720
rect 19800 14656 19816 14720
rect 19880 14656 19888 14720
rect 19568 14655 19888 14656
rect 5441 14514 5507 14517
rect 19333 14514 19399 14517
rect 5441 14512 19399 14514
rect 5441 14456 5446 14512
rect 5502 14456 19338 14512
rect 19394 14456 19399 14512
rect 5441 14454 19399 14456
rect 5441 14451 5507 14454
rect 19333 14451 19399 14454
rect 19701 14514 19767 14517
rect 27889 14514 27955 14517
rect 19701 14512 27955 14514
rect 19701 14456 19706 14512
rect 19762 14456 27894 14512
rect 27950 14456 27955 14512
rect 19701 14454 27955 14456
rect 19701 14451 19767 14454
rect 27889 14451 27955 14454
rect 15193 14378 15259 14381
rect 18597 14378 18663 14381
rect 15193 14376 18663 14378
rect 15193 14320 15198 14376
rect 15254 14320 18602 14376
rect 18658 14320 18663 14376
rect 15193 14318 18663 14320
rect 15193 14315 15259 14318
rect 18597 14315 18663 14318
rect 4208 14176 4528 14177
rect 4208 14112 4216 14176
rect 4280 14112 4296 14176
rect 4360 14112 4376 14176
rect 4440 14112 4456 14176
rect 4520 14112 4528 14176
rect 4208 14111 4528 14112
rect 34928 14176 35248 14177
rect 34928 14112 34936 14176
rect 35000 14112 35016 14176
rect 35080 14112 35096 14176
rect 35160 14112 35176 14176
rect 35240 14112 35248 14176
rect 34928 14111 35248 14112
rect 17033 13970 17099 13973
rect 22185 13970 22251 13973
rect 26141 13970 26207 13973
rect 17033 13968 26207 13970
rect 17033 13912 17038 13968
rect 17094 13912 22190 13968
rect 22246 13912 26146 13968
rect 26202 13912 26207 13968
rect 17033 13910 26207 13912
rect 17033 13907 17099 13910
rect 22185 13907 22251 13910
rect 26141 13907 26207 13910
rect 5809 13834 5875 13837
rect 18781 13834 18847 13837
rect 5809 13832 18847 13834
rect 5809 13776 5814 13832
rect 5870 13776 18786 13832
rect 18842 13776 18847 13832
rect 5809 13774 18847 13776
rect 5809 13771 5875 13774
rect 18781 13771 18847 13774
rect 20161 13834 20227 13837
rect 26877 13834 26943 13837
rect 20161 13832 26943 13834
rect 20161 13776 20166 13832
rect 20222 13776 26882 13832
rect 26938 13776 26943 13832
rect 20161 13774 26943 13776
rect 20161 13771 20227 13774
rect 26877 13771 26943 13774
rect 36997 13698 37063 13701
rect 40200 13698 41000 13728
rect 36997 13696 41000 13698
rect 36997 13640 37002 13696
rect 37058 13640 41000 13696
rect 36997 13638 41000 13640
rect 36997 13635 37063 13638
rect 19568 13632 19888 13633
rect 19568 13568 19576 13632
rect 19640 13568 19656 13632
rect 19720 13568 19736 13632
rect 19800 13568 19816 13632
rect 19880 13568 19888 13632
rect 40200 13608 41000 13638
rect 19568 13567 19888 13568
rect 25865 13426 25931 13429
rect 34513 13426 34579 13429
rect 4064 13366 17418 13426
rect 0 13154 800 13184
rect 4064 13154 4124 13366
rect 9949 13290 10015 13293
rect 17125 13290 17191 13293
rect 9949 13288 17191 13290
rect 9949 13232 9954 13288
rect 10010 13232 17130 13288
rect 17186 13232 17191 13288
rect 9949 13230 17191 13232
rect 17358 13290 17418 13366
rect 25865 13424 34579 13426
rect 25865 13368 25870 13424
rect 25926 13368 34518 13424
rect 34574 13368 34579 13424
rect 25865 13366 34579 13368
rect 25865 13363 25931 13366
rect 34513 13363 34579 13366
rect 20989 13290 21055 13293
rect 17358 13288 21055 13290
rect 17358 13232 20994 13288
rect 21050 13232 21055 13288
rect 17358 13230 21055 13232
rect 9949 13227 10015 13230
rect 17125 13227 17191 13230
rect 20989 13227 21055 13230
rect 23749 13290 23815 13293
rect 35709 13290 35775 13293
rect 23749 13288 35775 13290
rect 23749 13232 23754 13288
rect 23810 13232 35714 13288
rect 35770 13232 35775 13288
rect 23749 13230 35775 13232
rect 23749 13227 23815 13230
rect 35709 13227 35775 13230
rect 0 13094 4124 13154
rect 0 13064 800 13094
rect 4208 13088 4528 13089
rect 4208 13024 4216 13088
rect 4280 13024 4296 13088
rect 4360 13024 4376 13088
rect 4440 13024 4456 13088
rect 4520 13024 4528 13088
rect 4208 13023 4528 13024
rect 34928 13088 35248 13089
rect 34928 13024 34936 13088
rect 35000 13024 35016 13088
rect 35080 13024 35096 13088
rect 35160 13024 35176 13088
rect 35240 13024 35248 13088
rect 34928 13023 35248 13024
rect 36169 12882 36235 12885
rect 34286 12880 36235 12882
rect 34286 12824 36174 12880
rect 36230 12824 36235 12880
rect 34286 12822 36235 12824
rect 23289 12746 23355 12749
rect 23749 12746 23815 12749
rect 23289 12744 23815 12746
rect 23289 12688 23294 12744
rect 23350 12688 23754 12744
rect 23810 12688 23815 12744
rect 23289 12686 23815 12688
rect 23289 12683 23355 12686
rect 23749 12683 23815 12686
rect 31109 12746 31175 12749
rect 32397 12746 32463 12749
rect 34286 12746 34346 12822
rect 36169 12819 36235 12822
rect 31109 12744 34346 12746
rect 31109 12688 31114 12744
rect 31170 12688 32402 12744
rect 32458 12688 34346 12744
rect 31109 12686 34346 12688
rect 34421 12746 34487 12749
rect 34789 12746 34855 12749
rect 34421 12744 34855 12746
rect 34421 12688 34426 12744
rect 34482 12688 34794 12744
rect 34850 12688 34855 12744
rect 34421 12686 34855 12688
rect 31109 12683 31175 12686
rect 32397 12683 32463 12686
rect 34421 12683 34487 12686
rect 34789 12683 34855 12686
rect 15469 12610 15535 12613
rect 18413 12610 18479 12613
rect 15469 12608 18479 12610
rect 15469 12552 15474 12608
rect 15530 12552 18418 12608
rect 18474 12552 18479 12608
rect 15469 12550 18479 12552
rect 15469 12547 15535 12550
rect 18413 12547 18479 12550
rect 19568 12544 19888 12545
rect 19568 12480 19576 12544
rect 19640 12480 19656 12544
rect 19720 12480 19736 12544
rect 19800 12480 19816 12544
rect 19880 12480 19888 12544
rect 19568 12479 19888 12480
rect 30649 12338 30715 12341
rect 32949 12338 33015 12341
rect 30649 12336 33015 12338
rect 30649 12280 30654 12336
rect 30710 12280 32954 12336
rect 33010 12280 33015 12336
rect 30649 12278 33015 12280
rect 30649 12275 30715 12278
rect 32949 12275 33015 12278
rect 33501 12202 33567 12205
rect 33869 12202 33935 12205
rect 33501 12200 33935 12202
rect 33501 12144 33506 12200
rect 33562 12144 33874 12200
rect 33930 12144 33935 12200
rect 33501 12142 33935 12144
rect 33501 12139 33567 12142
rect 33869 12139 33935 12142
rect 4208 12000 4528 12001
rect 4208 11936 4216 12000
rect 4280 11936 4296 12000
rect 4360 11936 4376 12000
rect 4440 11936 4456 12000
rect 4520 11936 4528 12000
rect 4208 11935 4528 11936
rect 34928 12000 35248 12001
rect 34928 11936 34936 12000
rect 35000 11936 35016 12000
rect 35080 11936 35096 12000
rect 35160 11936 35176 12000
rect 35240 11936 35248 12000
rect 34928 11935 35248 11936
rect 12709 11794 12775 11797
rect 15101 11794 15167 11797
rect 12709 11792 15167 11794
rect 12709 11736 12714 11792
rect 12770 11736 15106 11792
rect 15162 11736 15167 11792
rect 12709 11734 15167 11736
rect 12709 11731 12775 11734
rect 15101 11731 15167 11734
rect 30741 11658 30807 11661
rect 37181 11658 37247 11661
rect 30741 11656 37247 11658
rect 30741 11600 30746 11656
rect 30802 11600 37186 11656
rect 37242 11600 37247 11656
rect 30741 11598 37247 11600
rect 30741 11595 30807 11598
rect 37181 11595 37247 11598
rect 19568 11456 19888 11457
rect 19568 11392 19576 11456
rect 19640 11392 19656 11456
rect 19720 11392 19736 11456
rect 19800 11392 19816 11456
rect 19880 11392 19888 11456
rect 19568 11391 19888 11392
rect 30097 11114 30163 11117
rect 35433 11114 35499 11117
rect 30097 11112 35499 11114
rect 30097 11056 30102 11112
rect 30158 11056 35438 11112
rect 35494 11056 35499 11112
rect 30097 11054 35499 11056
rect 30097 11051 30163 11054
rect 35433 11051 35499 11054
rect 4208 10912 4528 10913
rect 4208 10848 4216 10912
rect 4280 10848 4296 10912
rect 4360 10848 4376 10912
rect 4440 10848 4456 10912
rect 4520 10848 4528 10912
rect 4208 10847 4528 10848
rect 34928 10912 35248 10913
rect 34928 10848 34936 10912
rect 35000 10848 35016 10912
rect 35080 10848 35096 10912
rect 35160 10848 35176 10912
rect 35240 10848 35248 10912
rect 34928 10847 35248 10848
rect 21909 10706 21975 10709
rect 27521 10706 27587 10709
rect 21909 10704 27587 10706
rect 21909 10648 21914 10704
rect 21970 10648 27526 10704
rect 27582 10648 27587 10704
rect 21909 10646 27587 10648
rect 21909 10643 21975 10646
rect 27521 10643 27587 10646
rect 32857 10706 32923 10709
rect 36721 10706 36787 10709
rect 38561 10706 38627 10709
rect 32857 10704 38627 10706
rect 32857 10648 32862 10704
rect 32918 10648 36726 10704
rect 36782 10648 38566 10704
rect 38622 10648 38627 10704
rect 32857 10646 38627 10648
rect 32857 10643 32923 10646
rect 36721 10643 36787 10646
rect 38561 10643 38627 10646
rect 35893 10434 35959 10437
rect 40200 10434 41000 10464
rect 35893 10432 41000 10434
rect 35893 10376 35898 10432
rect 35954 10376 41000 10432
rect 35893 10374 41000 10376
rect 35893 10371 35959 10374
rect 19568 10368 19888 10369
rect 19568 10304 19576 10368
rect 19640 10304 19656 10368
rect 19720 10304 19736 10368
rect 19800 10304 19816 10368
rect 19880 10304 19888 10368
rect 40200 10344 41000 10374
rect 19568 10303 19888 10304
rect 0 10162 800 10192
rect 2773 10162 2839 10165
rect 0 10160 2839 10162
rect 0 10104 2778 10160
rect 2834 10104 2839 10160
rect 0 10102 2839 10104
rect 0 10072 800 10102
rect 2773 10099 2839 10102
rect 4208 9824 4528 9825
rect 4208 9760 4216 9824
rect 4280 9760 4296 9824
rect 4360 9760 4376 9824
rect 4440 9760 4456 9824
rect 4520 9760 4528 9824
rect 4208 9759 4528 9760
rect 34928 9824 35248 9825
rect 34928 9760 34936 9824
rect 35000 9760 35016 9824
rect 35080 9760 35096 9824
rect 35160 9760 35176 9824
rect 35240 9760 35248 9824
rect 34928 9759 35248 9760
rect 23565 9754 23631 9757
rect 23565 9752 23674 9754
rect 23565 9696 23570 9752
rect 23626 9696 23674 9752
rect 23565 9691 23674 9696
rect 23473 9618 23539 9621
rect 23614 9618 23674 9691
rect 23473 9616 23674 9618
rect 23473 9560 23478 9616
rect 23534 9560 23674 9616
rect 23473 9558 23674 9560
rect 23473 9555 23539 9558
rect 23657 9482 23723 9485
rect 26509 9482 26575 9485
rect 23657 9480 26575 9482
rect 23657 9424 23662 9480
rect 23718 9424 26514 9480
rect 26570 9424 26575 9480
rect 23657 9422 26575 9424
rect 23657 9419 23723 9422
rect 26509 9419 26575 9422
rect 19568 9280 19888 9281
rect 19568 9216 19576 9280
rect 19640 9216 19656 9280
rect 19720 9216 19736 9280
rect 19800 9216 19816 9280
rect 19880 9216 19888 9280
rect 19568 9215 19888 9216
rect 22829 9074 22895 9077
rect 25221 9074 25287 9077
rect 22829 9072 25287 9074
rect 22829 9016 22834 9072
rect 22890 9016 25226 9072
rect 25282 9016 25287 9072
rect 22829 9014 25287 9016
rect 22829 9011 22895 9014
rect 25221 9011 25287 9014
rect 4208 8736 4528 8737
rect 4208 8672 4216 8736
rect 4280 8672 4296 8736
rect 4360 8672 4376 8736
rect 4440 8672 4456 8736
rect 4520 8672 4528 8736
rect 4208 8671 4528 8672
rect 34928 8736 35248 8737
rect 34928 8672 34936 8736
rect 35000 8672 35016 8736
rect 35080 8672 35096 8736
rect 35160 8672 35176 8736
rect 35240 8672 35248 8736
rect 34928 8671 35248 8672
rect 19568 8192 19888 8193
rect 19568 8128 19576 8192
rect 19640 8128 19656 8192
rect 19720 8128 19736 8192
rect 19800 8128 19816 8192
rect 19880 8128 19888 8192
rect 19568 8127 19888 8128
rect 4208 7648 4528 7649
rect 4208 7584 4216 7648
rect 4280 7584 4296 7648
rect 4360 7584 4376 7648
rect 4440 7584 4456 7648
rect 4520 7584 4528 7648
rect 4208 7583 4528 7584
rect 34928 7648 35248 7649
rect 34928 7584 34936 7648
rect 35000 7584 35016 7648
rect 35080 7584 35096 7648
rect 35160 7584 35176 7648
rect 35240 7584 35248 7648
rect 34928 7583 35248 7584
rect 36721 7442 36787 7445
rect 40200 7442 41000 7472
rect 36721 7440 41000 7442
rect 36721 7384 36726 7440
rect 36782 7384 41000 7440
rect 36721 7382 41000 7384
rect 36721 7379 36787 7382
rect 40200 7352 41000 7382
rect 19568 7104 19888 7105
rect 19568 7040 19576 7104
rect 19640 7040 19656 7104
rect 19720 7040 19736 7104
rect 19800 7040 19816 7104
rect 19880 7040 19888 7104
rect 19568 7039 19888 7040
rect 0 6898 800 6928
rect 0 6838 1410 6898
rect 0 6808 800 6838
rect 1350 6626 1410 6838
rect 16757 6762 16823 6765
rect 25497 6762 25563 6765
rect 16757 6760 25563 6762
rect 16757 6704 16762 6760
rect 16818 6704 25502 6760
rect 25558 6704 25563 6760
rect 16757 6702 25563 6704
rect 16757 6699 16823 6702
rect 25497 6699 25563 6702
rect 2957 6626 3023 6629
rect 1350 6624 3023 6626
rect 1350 6568 2962 6624
rect 3018 6568 3023 6624
rect 1350 6566 3023 6568
rect 2957 6563 3023 6566
rect 4208 6560 4528 6561
rect 4208 6496 4216 6560
rect 4280 6496 4296 6560
rect 4360 6496 4376 6560
rect 4440 6496 4456 6560
rect 4520 6496 4528 6560
rect 4208 6495 4528 6496
rect 34928 6560 35248 6561
rect 34928 6496 34936 6560
rect 35000 6496 35016 6560
rect 35080 6496 35096 6560
rect 35160 6496 35176 6560
rect 35240 6496 35248 6560
rect 34928 6495 35248 6496
rect 13997 6354 14063 6357
rect 15837 6354 15903 6357
rect 13997 6352 15903 6354
rect 13997 6296 14002 6352
rect 14058 6296 15842 6352
rect 15898 6296 15903 6352
rect 13997 6294 15903 6296
rect 13997 6291 14063 6294
rect 15837 6291 15903 6294
rect 19568 6016 19888 6017
rect 19568 5952 19576 6016
rect 19640 5952 19656 6016
rect 19720 5952 19736 6016
rect 19800 5952 19816 6016
rect 19880 5952 19888 6016
rect 19568 5951 19888 5952
rect 13353 5946 13419 5949
rect 16021 5946 16087 5949
rect 13353 5944 16087 5946
rect 13353 5888 13358 5944
rect 13414 5888 16026 5944
rect 16082 5888 16087 5944
rect 13353 5886 16087 5888
rect 13353 5883 13419 5886
rect 16021 5883 16087 5886
rect 8753 5810 8819 5813
rect 24945 5810 25011 5813
rect 8753 5808 25011 5810
rect 8753 5752 8758 5808
rect 8814 5752 24950 5808
rect 25006 5752 25011 5808
rect 8753 5750 25011 5752
rect 8753 5747 8819 5750
rect 24945 5747 25011 5750
rect 11513 5674 11579 5677
rect 24853 5674 24919 5677
rect 11513 5672 24919 5674
rect 11513 5616 11518 5672
rect 11574 5616 24858 5672
rect 24914 5616 24919 5672
rect 11513 5614 24919 5616
rect 11513 5611 11579 5614
rect 24853 5611 24919 5614
rect 4208 5472 4528 5473
rect 4208 5408 4216 5472
rect 4280 5408 4296 5472
rect 4360 5408 4376 5472
rect 4440 5408 4456 5472
rect 4520 5408 4528 5472
rect 4208 5407 4528 5408
rect 34928 5472 35248 5473
rect 34928 5408 34936 5472
rect 35000 5408 35016 5472
rect 35080 5408 35096 5472
rect 35160 5408 35176 5472
rect 35240 5408 35248 5472
rect 34928 5407 35248 5408
rect 19568 4928 19888 4929
rect 19568 4864 19576 4928
rect 19640 4864 19656 4928
rect 19720 4864 19736 4928
rect 19800 4864 19816 4928
rect 19880 4864 19888 4928
rect 19568 4863 19888 4864
rect 4208 4384 4528 4385
rect 4208 4320 4216 4384
rect 4280 4320 4296 4384
rect 4360 4320 4376 4384
rect 4440 4320 4456 4384
rect 4520 4320 4528 4384
rect 4208 4319 4528 4320
rect 34928 4384 35248 4385
rect 34928 4320 34936 4384
rect 35000 4320 35016 4384
rect 35080 4320 35096 4384
rect 35160 4320 35176 4384
rect 35240 4320 35248 4384
rect 34928 4319 35248 4320
rect 17769 4178 17835 4181
rect 19241 4178 19307 4181
rect 17769 4176 19307 4178
rect 17769 4120 17774 4176
rect 17830 4120 19246 4176
rect 19302 4120 19307 4176
rect 17769 4118 19307 4120
rect 17769 4115 17835 4118
rect 19241 4115 19307 4118
rect 35893 4178 35959 4181
rect 40200 4178 41000 4208
rect 35893 4176 41000 4178
rect 35893 4120 35898 4176
rect 35954 4120 41000 4176
rect 35893 4118 41000 4120
rect 35893 4115 35959 4118
rect 40200 4088 41000 4118
rect 7097 4042 7163 4045
rect 9305 4042 9371 4045
rect 7097 4040 9371 4042
rect 7097 3984 7102 4040
rect 7158 3984 9310 4040
rect 9366 3984 9371 4040
rect 7097 3982 9371 3984
rect 7097 3979 7163 3982
rect 9305 3979 9371 3982
rect 0 3906 800 3936
rect 9213 3906 9279 3909
rect 0 3904 9279 3906
rect 0 3848 9218 3904
rect 9274 3848 9279 3904
rect 0 3846 9279 3848
rect 0 3816 800 3846
rect 9213 3843 9279 3846
rect 19568 3840 19888 3841
rect 19568 3776 19576 3840
rect 19640 3776 19656 3840
rect 19720 3776 19736 3840
rect 19800 3776 19816 3840
rect 19880 3776 19888 3840
rect 19568 3775 19888 3776
rect 12893 3770 12959 3773
rect 19057 3770 19123 3773
rect 12893 3768 19123 3770
rect 12893 3712 12898 3768
rect 12954 3712 19062 3768
rect 19118 3712 19123 3768
rect 12893 3710 19123 3712
rect 12893 3707 12959 3710
rect 19057 3707 19123 3710
rect 4208 3296 4528 3297
rect 4208 3232 4216 3296
rect 4280 3232 4296 3296
rect 4360 3232 4376 3296
rect 4440 3232 4456 3296
rect 4520 3232 4528 3296
rect 4208 3231 4528 3232
rect 34928 3296 35248 3297
rect 34928 3232 34936 3296
rect 35000 3232 35016 3296
rect 35080 3232 35096 3296
rect 35160 3232 35176 3296
rect 35240 3232 35248 3296
rect 34928 3231 35248 3232
rect 19568 2752 19888 2753
rect 19568 2688 19576 2752
rect 19640 2688 19656 2752
rect 19720 2688 19736 2752
rect 19800 2688 19816 2752
rect 19880 2688 19888 2752
rect 19568 2687 19888 2688
rect 4208 2208 4528 2209
rect 4208 2144 4216 2208
rect 4280 2144 4296 2208
rect 4360 2144 4376 2208
rect 4440 2144 4456 2208
rect 4520 2144 4528 2208
rect 4208 2143 4528 2144
rect 34928 2208 35248 2209
rect 34928 2144 34936 2208
rect 35000 2144 35016 2208
rect 35080 2144 35096 2208
rect 35160 2144 35176 2208
rect 35240 2144 35248 2208
rect 34928 2143 35248 2144
rect 36445 1186 36511 1189
rect 40200 1186 41000 1216
rect 36445 1184 41000 1186
rect 36445 1128 36450 1184
rect 36506 1128 41000 1184
rect 36445 1126 41000 1128
rect 36445 1123 36511 1126
rect 40200 1096 41000 1126
<< via3 >>
rect 19576 38652 19640 38656
rect 19576 38596 19580 38652
rect 19580 38596 19636 38652
rect 19636 38596 19640 38652
rect 19576 38592 19640 38596
rect 19656 38652 19720 38656
rect 19656 38596 19660 38652
rect 19660 38596 19716 38652
rect 19716 38596 19720 38652
rect 19656 38592 19720 38596
rect 19736 38652 19800 38656
rect 19736 38596 19740 38652
rect 19740 38596 19796 38652
rect 19796 38596 19800 38652
rect 19736 38592 19800 38596
rect 19816 38652 19880 38656
rect 19816 38596 19820 38652
rect 19820 38596 19876 38652
rect 19876 38596 19880 38652
rect 19816 38592 19880 38596
rect 4216 38108 4280 38112
rect 4216 38052 4220 38108
rect 4220 38052 4276 38108
rect 4276 38052 4280 38108
rect 4216 38048 4280 38052
rect 4296 38108 4360 38112
rect 4296 38052 4300 38108
rect 4300 38052 4356 38108
rect 4356 38052 4360 38108
rect 4296 38048 4360 38052
rect 4376 38108 4440 38112
rect 4376 38052 4380 38108
rect 4380 38052 4436 38108
rect 4436 38052 4440 38108
rect 4376 38048 4440 38052
rect 4456 38108 4520 38112
rect 4456 38052 4460 38108
rect 4460 38052 4516 38108
rect 4516 38052 4520 38108
rect 4456 38048 4520 38052
rect 34936 38108 35000 38112
rect 34936 38052 34940 38108
rect 34940 38052 34996 38108
rect 34996 38052 35000 38108
rect 34936 38048 35000 38052
rect 35016 38108 35080 38112
rect 35016 38052 35020 38108
rect 35020 38052 35076 38108
rect 35076 38052 35080 38108
rect 35016 38048 35080 38052
rect 35096 38108 35160 38112
rect 35096 38052 35100 38108
rect 35100 38052 35156 38108
rect 35156 38052 35160 38108
rect 35096 38048 35160 38052
rect 35176 38108 35240 38112
rect 35176 38052 35180 38108
rect 35180 38052 35236 38108
rect 35236 38052 35240 38108
rect 35176 38048 35240 38052
rect 19576 37564 19640 37568
rect 19576 37508 19580 37564
rect 19580 37508 19636 37564
rect 19636 37508 19640 37564
rect 19576 37504 19640 37508
rect 19656 37564 19720 37568
rect 19656 37508 19660 37564
rect 19660 37508 19716 37564
rect 19716 37508 19720 37564
rect 19656 37504 19720 37508
rect 19736 37564 19800 37568
rect 19736 37508 19740 37564
rect 19740 37508 19796 37564
rect 19796 37508 19800 37564
rect 19736 37504 19800 37508
rect 19816 37564 19880 37568
rect 19816 37508 19820 37564
rect 19820 37508 19876 37564
rect 19876 37508 19880 37564
rect 19816 37504 19880 37508
rect 4216 37020 4280 37024
rect 4216 36964 4220 37020
rect 4220 36964 4276 37020
rect 4276 36964 4280 37020
rect 4216 36960 4280 36964
rect 4296 37020 4360 37024
rect 4296 36964 4300 37020
rect 4300 36964 4356 37020
rect 4356 36964 4360 37020
rect 4296 36960 4360 36964
rect 4376 37020 4440 37024
rect 4376 36964 4380 37020
rect 4380 36964 4436 37020
rect 4436 36964 4440 37020
rect 4376 36960 4440 36964
rect 4456 37020 4520 37024
rect 4456 36964 4460 37020
rect 4460 36964 4516 37020
rect 4516 36964 4520 37020
rect 4456 36960 4520 36964
rect 34936 37020 35000 37024
rect 34936 36964 34940 37020
rect 34940 36964 34996 37020
rect 34996 36964 35000 37020
rect 34936 36960 35000 36964
rect 35016 37020 35080 37024
rect 35016 36964 35020 37020
rect 35020 36964 35076 37020
rect 35076 36964 35080 37020
rect 35016 36960 35080 36964
rect 35096 37020 35160 37024
rect 35096 36964 35100 37020
rect 35100 36964 35156 37020
rect 35156 36964 35160 37020
rect 35096 36960 35160 36964
rect 35176 37020 35240 37024
rect 35176 36964 35180 37020
rect 35180 36964 35236 37020
rect 35236 36964 35240 37020
rect 35176 36960 35240 36964
rect 19576 36476 19640 36480
rect 19576 36420 19580 36476
rect 19580 36420 19636 36476
rect 19636 36420 19640 36476
rect 19576 36416 19640 36420
rect 19656 36476 19720 36480
rect 19656 36420 19660 36476
rect 19660 36420 19716 36476
rect 19716 36420 19720 36476
rect 19656 36416 19720 36420
rect 19736 36476 19800 36480
rect 19736 36420 19740 36476
rect 19740 36420 19796 36476
rect 19796 36420 19800 36476
rect 19736 36416 19800 36420
rect 19816 36476 19880 36480
rect 19816 36420 19820 36476
rect 19820 36420 19876 36476
rect 19876 36420 19880 36476
rect 19816 36416 19880 36420
rect 4216 35932 4280 35936
rect 4216 35876 4220 35932
rect 4220 35876 4276 35932
rect 4276 35876 4280 35932
rect 4216 35872 4280 35876
rect 4296 35932 4360 35936
rect 4296 35876 4300 35932
rect 4300 35876 4356 35932
rect 4356 35876 4360 35932
rect 4296 35872 4360 35876
rect 4376 35932 4440 35936
rect 4376 35876 4380 35932
rect 4380 35876 4436 35932
rect 4436 35876 4440 35932
rect 4376 35872 4440 35876
rect 4456 35932 4520 35936
rect 4456 35876 4460 35932
rect 4460 35876 4516 35932
rect 4516 35876 4520 35932
rect 4456 35872 4520 35876
rect 34936 35932 35000 35936
rect 34936 35876 34940 35932
rect 34940 35876 34996 35932
rect 34996 35876 35000 35932
rect 34936 35872 35000 35876
rect 35016 35932 35080 35936
rect 35016 35876 35020 35932
rect 35020 35876 35076 35932
rect 35076 35876 35080 35932
rect 35016 35872 35080 35876
rect 35096 35932 35160 35936
rect 35096 35876 35100 35932
rect 35100 35876 35156 35932
rect 35156 35876 35160 35932
rect 35096 35872 35160 35876
rect 35176 35932 35240 35936
rect 35176 35876 35180 35932
rect 35180 35876 35236 35932
rect 35236 35876 35240 35932
rect 35176 35872 35240 35876
rect 19576 35388 19640 35392
rect 19576 35332 19580 35388
rect 19580 35332 19636 35388
rect 19636 35332 19640 35388
rect 19576 35328 19640 35332
rect 19656 35388 19720 35392
rect 19656 35332 19660 35388
rect 19660 35332 19716 35388
rect 19716 35332 19720 35388
rect 19656 35328 19720 35332
rect 19736 35388 19800 35392
rect 19736 35332 19740 35388
rect 19740 35332 19796 35388
rect 19796 35332 19800 35388
rect 19736 35328 19800 35332
rect 19816 35388 19880 35392
rect 19816 35332 19820 35388
rect 19820 35332 19876 35388
rect 19876 35332 19880 35388
rect 19816 35328 19880 35332
rect 4216 34844 4280 34848
rect 4216 34788 4220 34844
rect 4220 34788 4276 34844
rect 4276 34788 4280 34844
rect 4216 34784 4280 34788
rect 4296 34844 4360 34848
rect 4296 34788 4300 34844
rect 4300 34788 4356 34844
rect 4356 34788 4360 34844
rect 4296 34784 4360 34788
rect 4376 34844 4440 34848
rect 4376 34788 4380 34844
rect 4380 34788 4436 34844
rect 4436 34788 4440 34844
rect 4376 34784 4440 34788
rect 4456 34844 4520 34848
rect 4456 34788 4460 34844
rect 4460 34788 4516 34844
rect 4516 34788 4520 34844
rect 4456 34784 4520 34788
rect 34936 34844 35000 34848
rect 34936 34788 34940 34844
rect 34940 34788 34996 34844
rect 34996 34788 35000 34844
rect 34936 34784 35000 34788
rect 35016 34844 35080 34848
rect 35016 34788 35020 34844
rect 35020 34788 35076 34844
rect 35076 34788 35080 34844
rect 35016 34784 35080 34788
rect 35096 34844 35160 34848
rect 35096 34788 35100 34844
rect 35100 34788 35156 34844
rect 35156 34788 35160 34844
rect 35096 34784 35160 34788
rect 35176 34844 35240 34848
rect 35176 34788 35180 34844
rect 35180 34788 35236 34844
rect 35236 34788 35240 34844
rect 35176 34784 35240 34788
rect 19576 34300 19640 34304
rect 19576 34244 19580 34300
rect 19580 34244 19636 34300
rect 19636 34244 19640 34300
rect 19576 34240 19640 34244
rect 19656 34300 19720 34304
rect 19656 34244 19660 34300
rect 19660 34244 19716 34300
rect 19716 34244 19720 34300
rect 19656 34240 19720 34244
rect 19736 34300 19800 34304
rect 19736 34244 19740 34300
rect 19740 34244 19796 34300
rect 19796 34244 19800 34300
rect 19736 34240 19800 34244
rect 19816 34300 19880 34304
rect 19816 34244 19820 34300
rect 19820 34244 19876 34300
rect 19876 34244 19880 34300
rect 19816 34240 19880 34244
rect 4216 33756 4280 33760
rect 4216 33700 4220 33756
rect 4220 33700 4276 33756
rect 4276 33700 4280 33756
rect 4216 33696 4280 33700
rect 4296 33756 4360 33760
rect 4296 33700 4300 33756
rect 4300 33700 4356 33756
rect 4356 33700 4360 33756
rect 4296 33696 4360 33700
rect 4376 33756 4440 33760
rect 4376 33700 4380 33756
rect 4380 33700 4436 33756
rect 4436 33700 4440 33756
rect 4376 33696 4440 33700
rect 4456 33756 4520 33760
rect 4456 33700 4460 33756
rect 4460 33700 4516 33756
rect 4516 33700 4520 33756
rect 4456 33696 4520 33700
rect 34936 33756 35000 33760
rect 34936 33700 34940 33756
rect 34940 33700 34996 33756
rect 34996 33700 35000 33756
rect 34936 33696 35000 33700
rect 35016 33756 35080 33760
rect 35016 33700 35020 33756
rect 35020 33700 35076 33756
rect 35076 33700 35080 33756
rect 35016 33696 35080 33700
rect 35096 33756 35160 33760
rect 35096 33700 35100 33756
rect 35100 33700 35156 33756
rect 35156 33700 35160 33756
rect 35096 33696 35160 33700
rect 35176 33756 35240 33760
rect 35176 33700 35180 33756
rect 35180 33700 35236 33756
rect 35236 33700 35240 33756
rect 35176 33696 35240 33700
rect 19576 33212 19640 33216
rect 19576 33156 19580 33212
rect 19580 33156 19636 33212
rect 19636 33156 19640 33212
rect 19576 33152 19640 33156
rect 19656 33212 19720 33216
rect 19656 33156 19660 33212
rect 19660 33156 19716 33212
rect 19716 33156 19720 33212
rect 19656 33152 19720 33156
rect 19736 33212 19800 33216
rect 19736 33156 19740 33212
rect 19740 33156 19796 33212
rect 19796 33156 19800 33212
rect 19736 33152 19800 33156
rect 19816 33212 19880 33216
rect 19816 33156 19820 33212
rect 19820 33156 19876 33212
rect 19876 33156 19880 33212
rect 19816 33152 19880 33156
rect 4216 32668 4280 32672
rect 4216 32612 4220 32668
rect 4220 32612 4276 32668
rect 4276 32612 4280 32668
rect 4216 32608 4280 32612
rect 4296 32668 4360 32672
rect 4296 32612 4300 32668
rect 4300 32612 4356 32668
rect 4356 32612 4360 32668
rect 4296 32608 4360 32612
rect 4376 32668 4440 32672
rect 4376 32612 4380 32668
rect 4380 32612 4436 32668
rect 4436 32612 4440 32668
rect 4376 32608 4440 32612
rect 4456 32668 4520 32672
rect 4456 32612 4460 32668
rect 4460 32612 4516 32668
rect 4516 32612 4520 32668
rect 4456 32608 4520 32612
rect 34936 32668 35000 32672
rect 34936 32612 34940 32668
rect 34940 32612 34996 32668
rect 34996 32612 35000 32668
rect 34936 32608 35000 32612
rect 35016 32668 35080 32672
rect 35016 32612 35020 32668
rect 35020 32612 35076 32668
rect 35076 32612 35080 32668
rect 35016 32608 35080 32612
rect 35096 32668 35160 32672
rect 35096 32612 35100 32668
rect 35100 32612 35156 32668
rect 35156 32612 35160 32668
rect 35096 32608 35160 32612
rect 35176 32668 35240 32672
rect 35176 32612 35180 32668
rect 35180 32612 35236 32668
rect 35236 32612 35240 32668
rect 35176 32608 35240 32612
rect 19576 32124 19640 32128
rect 19576 32068 19580 32124
rect 19580 32068 19636 32124
rect 19636 32068 19640 32124
rect 19576 32064 19640 32068
rect 19656 32124 19720 32128
rect 19656 32068 19660 32124
rect 19660 32068 19716 32124
rect 19716 32068 19720 32124
rect 19656 32064 19720 32068
rect 19736 32124 19800 32128
rect 19736 32068 19740 32124
rect 19740 32068 19796 32124
rect 19796 32068 19800 32124
rect 19736 32064 19800 32068
rect 19816 32124 19880 32128
rect 19816 32068 19820 32124
rect 19820 32068 19876 32124
rect 19876 32068 19880 32124
rect 19816 32064 19880 32068
rect 4216 31580 4280 31584
rect 4216 31524 4220 31580
rect 4220 31524 4276 31580
rect 4276 31524 4280 31580
rect 4216 31520 4280 31524
rect 4296 31580 4360 31584
rect 4296 31524 4300 31580
rect 4300 31524 4356 31580
rect 4356 31524 4360 31580
rect 4296 31520 4360 31524
rect 4376 31580 4440 31584
rect 4376 31524 4380 31580
rect 4380 31524 4436 31580
rect 4436 31524 4440 31580
rect 4376 31520 4440 31524
rect 4456 31580 4520 31584
rect 4456 31524 4460 31580
rect 4460 31524 4516 31580
rect 4516 31524 4520 31580
rect 4456 31520 4520 31524
rect 34936 31580 35000 31584
rect 34936 31524 34940 31580
rect 34940 31524 34996 31580
rect 34996 31524 35000 31580
rect 34936 31520 35000 31524
rect 35016 31580 35080 31584
rect 35016 31524 35020 31580
rect 35020 31524 35076 31580
rect 35076 31524 35080 31580
rect 35016 31520 35080 31524
rect 35096 31580 35160 31584
rect 35096 31524 35100 31580
rect 35100 31524 35156 31580
rect 35156 31524 35160 31580
rect 35096 31520 35160 31524
rect 35176 31580 35240 31584
rect 35176 31524 35180 31580
rect 35180 31524 35236 31580
rect 35236 31524 35240 31580
rect 35176 31520 35240 31524
rect 19576 31036 19640 31040
rect 19576 30980 19580 31036
rect 19580 30980 19636 31036
rect 19636 30980 19640 31036
rect 19576 30976 19640 30980
rect 19656 31036 19720 31040
rect 19656 30980 19660 31036
rect 19660 30980 19716 31036
rect 19716 30980 19720 31036
rect 19656 30976 19720 30980
rect 19736 31036 19800 31040
rect 19736 30980 19740 31036
rect 19740 30980 19796 31036
rect 19796 30980 19800 31036
rect 19736 30976 19800 30980
rect 19816 31036 19880 31040
rect 19816 30980 19820 31036
rect 19820 30980 19876 31036
rect 19876 30980 19880 31036
rect 19816 30976 19880 30980
rect 4216 30492 4280 30496
rect 4216 30436 4220 30492
rect 4220 30436 4276 30492
rect 4276 30436 4280 30492
rect 4216 30432 4280 30436
rect 4296 30492 4360 30496
rect 4296 30436 4300 30492
rect 4300 30436 4356 30492
rect 4356 30436 4360 30492
rect 4296 30432 4360 30436
rect 4376 30492 4440 30496
rect 4376 30436 4380 30492
rect 4380 30436 4436 30492
rect 4436 30436 4440 30492
rect 4376 30432 4440 30436
rect 4456 30492 4520 30496
rect 4456 30436 4460 30492
rect 4460 30436 4516 30492
rect 4516 30436 4520 30492
rect 4456 30432 4520 30436
rect 34936 30492 35000 30496
rect 34936 30436 34940 30492
rect 34940 30436 34996 30492
rect 34996 30436 35000 30492
rect 34936 30432 35000 30436
rect 35016 30492 35080 30496
rect 35016 30436 35020 30492
rect 35020 30436 35076 30492
rect 35076 30436 35080 30492
rect 35016 30432 35080 30436
rect 35096 30492 35160 30496
rect 35096 30436 35100 30492
rect 35100 30436 35156 30492
rect 35156 30436 35160 30492
rect 35096 30432 35160 30436
rect 35176 30492 35240 30496
rect 35176 30436 35180 30492
rect 35180 30436 35236 30492
rect 35236 30436 35240 30492
rect 35176 30432 35240 30436
rect 19576 29948 19640 29952
rect 19576 29892 19580 29948
rect 19580 29892 19636 29948
rect 19636 29892 19640 29948
rect 19576 29888 19640 29892
rect 19656 29948 19720 29952
rect 19656 29892 19660 29948
rect 19660 29892 19716 29948
rect 19716 29892 19720 29948
rect 19656 29888 19720 29892
rect 19736 29948 19800 29952
rect 19736 29892 19740 29948
rect 19740 29892 19796 29948
rect 19796 29892 19800 29948
rect 19736 29888 19800 29892
rect 19816 29948 19880 29952
rect 19816 29892 19820 29948
rect 19820 29892 19876 29948
rect 19876 29892 19880 29948
rect 19816 29888 19880 29892
rect 4216 29404 4280 29408
rect 4216 29348 4220 29404
rect 4220 29348 4276 29404
rect 4276 29348 4280 29404
rect 4216 29344 4280 29348
rect 4296 29404 4360 29408
rect 4296 29348 4300 29404
rect 4300 29348 4356 29404
rect 4356 29348 4360 29404
rect 4296 29344 4360 29348
rect 4376 29404 4440 29408
rect 4376 29348 4380 29404
rect 4380 29348 4436 29404
rect 4436 29348 4440 29404
rect 4376 29344 4440 29348
rect 4456 29404 4520 29408
rect 4456 29348 4460 29404
rect 4460 29348 4516 29404
rect 4516 29348 4520 29404
rect 4456 29344 4520 29348
rect 34936 29404 35000 29408
rect 34936 29348 34940 29404
rect 34940 29348 34996 29404
rect 34996 29348 35000 29404
rect 34936 29344 35000 29348
rect 35016 29404 35080 29408
rect 35016 29348 35020 29404
rect 35020 29348 35076 29404
rect 35076 29348 35080 29404
rect 35016 29344 35080 29348
rect 35096 29404 35160 29408
rect 35096 29348 35100 29404
rect 35100 29348 35156 29404
rect 35156 29348 35160 29404
rect 35096 29344 35160 29348
rect 35176 29404 35240 29408
rect 35176 29348 35180 29404
rect 35180 29348 35236 29404
rect 35236 29348 35240 29404
rect 35176 29344 35240 29348
rect 18828 28928 18892 28932
rect 18828 28872 18878 28928
rect 18878 28872 18892 28928
rect 18828 28868 18892 28872
rect 19576 28860 19640 28864
rect 19576 28804 19580 28860
rect 19580 28804 19636 28860
rect 19636 28804 19640 28860
rect 19576 28800 19640 28804
rect 19656 28860 19720 28864
rect 19656 28804 19660 28860
rect 19660 28804 19716 28860
rect 19716 28804 19720 28860
rect 19656 28800 19720 28804
rect 19736 28860 19800 28864
rect 19736 28804 19740 28860
rect 19740 28804 19796 28860
rect 19796 28804 19800 28860
rect 19736 28800 19800 28804
rect 19816 28860 19880 28864
rect 19816 28804 19820 28860
rect 19820 28804 19876 28860
rect 19876 28804 19880 28860
rect 19816 28800 19880 28804
rect 4216 28316 4280 28320
rect 4216 28260 4220 28316
rect 4220 28260 4276 28316
rect 4276 28260 4280 28316
rect 4216 28256 4280 28260
rect 4296 28316 4360 28320
rect 4296 28260 4300 28316
rect 4300 28260 4356 28316
rect 4356 28260 4360 28316
rect 4296 28256 4360 28260
rect 4376 28316 4440 28320
rect 4376 28260 4380 28316
rect 4380 28260 4436 28316
rect 4436 28260 4440 28316
rect 4376 28256 4440 28260
rect 4456 28316 4520 28320
rect 4456 28260 4460 28316
rect 4460 28260 4516 28316
rect 4516 28260 4520 28316
rect 4456 28256 4520 28260
rect 34936 28316 35000 28320
rect 34936 28260 34940 28316
rect 34940 28260 34996 28316
rect 34996 28260 35000 28316
rect 34936 28256 35000 28260
rect 35016 28316 35080 28320
rect 35016 28260 35020 28316
rect 35020 28260 35076 28316
rect 35076 28260 35080 28316
rect 35016 28256 35080 28260
rect 35096 28316 35160 28320
rect 35096 28260 35100 28316
rect 35100 28260 35156 28316
rect 35156 28260 35160 28316
rect 35096 28256 35160 28260
rect 35176 28316 35240 28320
rect 35176 28260 35180 28316
rect 35180 28260 35236 28316
rect 35236 28260 35240 28316
rect 35176 28256 35240 28260
rect 19576 27772 19640 27776
rect 19576 27716 19580 27772
rect 19580 27716 19636 27772
rect 19636 27716 19640 27772
rect 19576 27712 19640 27716
rect 19656 27772 19720 27776
rect 19656 27716 19660 27772
rect 19660 27716 19716 27772
rect 19716 27716 19720 27772
rect 19656 27712 19720 27716
rect 19736 27772 19800 27776
rect 19736 27716 19740 27772
rect 19740 27716 19796 27772
rect 19796 27716 19800 27772
rect 19736 27712 19800 27716
rect 19816 27772 19880 27776
rect 19816 27716 19820 27772
rect 19820 27716 19876 27772
rect 19876 27716 19880 27772
rect 19816 27712 19880 27716
rect 4216 27228 4280 27232
rect 4216 27172 4220 27228
rect 4220 27172 4276 27228
rect 4276 27172 4280 27228
rect 4216 27168 4280 27172
rect 4296 27228 4360 27232
rect 4296 27172 4300 27228
rect 4300 27172 4356 27228
rect 4356 27172 4360 27228
rect 4296 27168 4360 27172
rect 4376 27228 4440 27232
rect 4376 27172 4380 27228
rect 4380 27172 4436 27228
rect 4436 27172 4440 27228
rect 4376 27168 4440 27172
rect 4456 27228 4520 27232
rect 4456 27172 4460 27228
rect 4460 27172 4516 27228
rect 4516 27172 4520 27228
rect 4456 27168 4520 27172
rect 34936 27228 35000 27232
rect 34936 27172 34940 27228
rect 34940 27172 34996 27228
rect 34996 27172 35000 27228
rect 34936 27168 35000 27172
rect 35016 27228 35080 27232
rect 35016 27172 35020 27228
rect 35020 27172 35076 27228
rect 35076 27172 35080 27228
rect 35016 27168 35080 27172
rect 35096 27228 35160 27232
rect 35096 27172 35100 27228
rect 35100 27172 35156 27228
rect 35156 27172 35160 27228
rect 35096 27168 35160 27172
rect 35176 27228 35240 27232
rect 35176 27172 35180 27228
rect 35180 27172 35236 27228
rect 35236 27172 35240 27228
rect 35176 27168 35240 27172
rect 19576 26684 19640 26688
rect 19576 26628 19580 26684
rect 19580 26628 19636 26684
rect 19636 26628 19640 26684
rect 19576 26624 19640 26628
rect 19656 26684 19720 26688
rect 19656 26628 19660 26684
rect 19660 26628 19716 26684
rect 19716 26628 19720 26684
rect 19656 26624 19720 26628
rect 19736 26684 19800 26688
rect 19736 26628 19740 26684
rect 19740 26628 19796 26684
rect 19796 26628 19800 26684
rect 19736 26624 19800 26628
rect 19816 26684 19880 26688
rect 19816 26628 19820 26684
rect 19820 26628 19876 26684
rect 19876 26628 19880 26684
rect 19816 26624 19880 26628
rect 4216 26140 4280 26144
rect 4216 26084 4220 26140
rect 4220 26084 4276 26140
rect 4276 26084 4280 26140
rect 4216 26080 4280 26084
rect 4296 26140 4360 26144
rect 4296 26084 4300 26140
rect 4300 26084 4356 26140
rect 4356 26084 4360 26140
rect 4296 26080 4360 26084
rect 4376 26140 4440 26144
rect 4376 26084 4380 26140
rect 4380 26084 4436 26140
rect 4436 26084 4440 26140
rect 4376 26080 4440 26084
rect 4456 26140 4520 26144
rect 4456 26084 4460 26140
rect 4460 26084 4516 26140
rect 4516 26084 4520 26140
rect 4456 26080 4520 26084
rect 34936 26140 35000 26144
rect 34936 26084 34940 26140
rect 34940 26084 34996 26140
rect 34996 26084 35000 26140
rect 34936 26080 35000 26084
rect 35016 26140 35080 26144
rect 35016 26084 35020 26140
rect 35020 26084 35076 26140
rect 35076 26084 35080 26140
rect 35016 26080 35080 26084
rect 35096 26140 35160 26144
rect 35096 26084 35100 26140
rect 35100 26084 35156 26140
rect 35156 26084 35160 26140
rect 35096 26080 35160 26084
rect 35176 26140 35240 26144
rect 35176 26084 35180 26140
rect 35180 26084 35236 26140
rect 35236 26084 35240 26140
rect 35176 26080 35240 26084
rect 19576 25596 19640 25600
rect 19576 25540 19580 25596
rect 19580 25540 19636 25596
rect 19636 25540 19640 25596
rect 19576 25536 19640 25540
rect 19656 25596 19720 25600
rect 19656 25540 19660 25596
rect 19660 25540 19716 25596
rect 19716 25540 19720 25596
rect 19656 25536 19720 25540
rect 19736 25596 19800 25600
rect 19736 25540 19740 25596
rect 19740 25540 19796 25596
rect 19796 25540 19800 25596
rect 19736 25536 19800 25540
rect 19816 25596 19880 25600
rect 19816 25540 19820 25596
rect 19820 25540 19876 25596
rect 19876 25540 19880 25596
rect 19816 25536 19880 25540
rect 4216 25052 4280 25056
rect 4216 24996 4220 25052
rect 4220 24996 4276 25052
rect 4276 24996 4280 25052
rect 4216 24992 4280 24996
rect 4296 25052 4360 25056
rect 4296 24996 4300 25052
rect 4300 24996 4356 25052
rect 4356 24996 4360 25052
rect 4296 24992 4360 24996
rect 4376 25052 4440 25056
rect 4376 24996 4380 25052
rect 4380 24996 4436 25052
rect 4436 24996 4440 25052
rect 4376 24992 4440 24996
rect 4456 25052 4520 25056
rect 4456 24996 4460 25052
rect 4460 24996 4516 25052
rect 4516 24996 4520 25052
rect 4456 24992 4520 24996
rect 34936 25052 35000 25056
rect 34936 24996 34940 25052
rect 34940 24996 34996 25052
rect 34996 24996 35000 25052
rect 34936 24992 35000 24996
rect 35016 25052 35080 25056
rect 35016 24996 35020 25052
rect 35020 24996 35076 25052
rect 35076 24996 35080 25052
rect 35016 24992 35080 24996
rect 35096 25052 35160 25056
rect 35096 24996 35100 25052
rect 35100 24996 35156 25052
rect 35156 24996 35160 25052
rect 35096 24992 35160 24996
rect 35176 25052 35240 25056
rect 35176 24996 35180 25052
rect 35180 24996 35236 25052
rect 35236 24996 35240 25052
rect 35176 24992 35240 24996
rect 19576 24508 19640 24512
rect 19576 24452 19580 24508
rect 19580 24452 19636 24508
rect 19636 24452 19640 24508
rect 19576 24448 19640 24452
rect 19656 24508 19720 24512
rect 19656 24452 19660 24508
rect 19660 24452 19716 24508
rect 19716 24452 19720 24508
rect 19656 24448 19720 24452
rect 19736 24508 19800 24512
rect 19736 24452 19740 24508
rect 19740 24452 19796 24508
rect 19796 24452 19800 24508
rect 19736 24448 19800 24452
rect 19816 24508 19880 24512
rect 19816 24452 19820 24508
rect 19820 24452 19876 24508
rect 19876 24452 19880 24508
rect 19816 24448 19880 24452
rect 4216 23964 4280 23968
rect 4216 23908 4220 23964
rect 4220 23908 4276 23964
rect 4276 23908 4280 23964
rect 4216 23904 4280 23908
rect 4296 23964 4360 23968
rect 4296 23908 4300 23964
rect 4300 23908 4356 23964
rect 4356 23908 4360 23964
rect 4296 23904 4360 23908
rect 4376 23964 4440 23968
rect 4376 23908 4380 23964
rect 4380 23908 4436 23964
rect 4436 23908 4440 23964
rect 4376 23904 4440 23908
rect 4456 23964 4520 23968
rect 4456 23908 4460 23964
rect 4460 23908 4516 23964
rect 4516 23908 4520 23964
rect 4456 23904 4520 23908
rect 34936 23964 35000 23968
rect 34936 23908 34940 23964
rect 34940 23908 34996 23964
rect 34996 23908 35000 23964
rect 34936 23904 35000 23908
rect 35016 23964 35080 23968
rect 35016 23908 35020 23964
rect 35020 23908 35076 23964
rect 35076 23908 35080 23964
rect 35016 23904 35080 23908
rect 35096 23964 35160 23968
rect 35096 23908 35100 23964
rect 35100 23908 35156 23964
rect 35156 23908 35160 23964
rect 35096 23904 35160 23908
rect 35176 23964 35240 23968
rect 35176 23908 35180 23964
rect 35180 23908 35236 23964
rect 35236 23908 35240 23964
rect 35176 23904 35240 23908
rect 19576 23420 19640 23424
rect 19576 23364 19580 23420
rect 19580 23364 19636 23420
rect 19636 23364 19640 23420
rect 19576 23360 19640 23364
rect 19656 23420 19720 23424
rect 19656 23364 19660 23420
rect 19660 23364 19716 23420
rect 19716 23364 19720 23420
rect 19656 23360 19720 23364
rect 19736 23420 19800 23424
rect 19736 23364 19740 23420
rect 19740 23364 19796 23420
rect 19796 23364 19800 23420
rect 19736 23360 19800 23364
rect 19816 23420 19880 23424
rect 19816 23364 19820 23420
rect 19820 23364 19876 23420
rect 19876 23364 19880 23420
rect 19816 23360 19880 23364
rect 18828 23216 18892 23220
rect 18828 23160 18878 23216
rect 18878 23160 18892 23216
rect 18828 23156 18892 23160
rect 4216 22876 4280 22880
rect 4216 22820 4220 22876
rect 4220 22820 4276 22876
rect 4276 22820 4280 22876
rect 4216 22816 4280 22820
rect 4296 22876 4360 22880
rect 4296 22820 4300 22876
rect 4300 22820 4356 22876
rect 4356 22820 4360 22876
rect 4296 22816 4360 22820
rect 4376 22876 4440 22880
rect 4376 22820 4380 22876
rect 4380 22820 4436 22876
rect 4436 22820 4440 22876
rect 4376 22816 4440 22820
rect 4456 22876 4520 22880
rect 4456 22820 4460 22876
rect 4460 22820 4516 22876
rect 4516 22820 4520 22876
rect 4456 22816 4520 22820
rect 34936 22876 35000 22880
rect 34936 22820 34940 22876
rect 34940 22820 34996 22876
rect 34996 22820 35000 22876
rect 34936 22816 35000 22820
rect 35016 22876 35080 22880
rect 35016 22820 35020 22876
rect 35020 22820 35076 22876
rect 35076 22820 35080 22876
rect 35016 22816 35080 22820
rect 35096 22876 35160 22880
rect 35096 22820 35100 22876
rect 35100 22820 35156 22876
rect 35156 22820 35160 22876
rect 35096 22816 35160 22820
rect 35176 22876 35240 22880
rect 35176 22820 35180 22876
rect 35180 22820 35236 22876
rect 35236 22820 35240 22876
rect 35176 22816 35240 22820
rect 19576 22332 19640 22336
rect 19576 22276 19580 22332
rect 19580 22276 19636 22332
rect 19636 22276 19640 22332
rect 19576 22272 19640 22276
rect 19656 22332 19720 22336
rect 19656 22276 19660 22332
rect 19660 22276 19716 22332
rect 19716 22276 19720 22332
rect 19656 22272 19720 22276
rect 19736 22332 19800 22336
rect 19736 22276 19740 22332
rect 19740 22276 19796 22332
rect 19796 22276 19800 22332
rect 19736 22272 19800 22276
rect 19816 22332 19880 22336
rect 19816 22276 19820 22332
rect 19820 22276 19876 22332
rect 19876 22276 19880 22332
rect 19816 22272 19880 22276
rect 4216 21788 4280 21792
rect 4216 21732 4220 21788
rect 4220 21732 4276 21788
rect 4276 21732 4280 21788
rect 4216 21728 4280 21732
rect 4296 21788 4360 21792
rect 4296 21732 4300 21788
rect 4300 21732 4356 21788
rect 4356 21732 4360 21788
rect 4296 21728 4360 21732
rect 4376 21788 4440 21792
rect 4376 21732 4380 21788
rect 4380 21732 4436 21788
rect 4436 21732 4440 21788
rect 4376 21728 4440 21732
rect 4456 21788 4520 21792
rect 4456 21732 4460 21788
rect 4460 21732 4516 21788
rect 4516 21732 4520 21788
rect 4456 21728 4520 21732
rect 34936 21788 35000 21792
rect 34936 21732 34940 21788
rect 34940 21732 34996 21788
rect 34996 21732 35000 21788
rect 34936 21728 35000 21732
rect 35016 21788 35080 21792
rect 35016 21732 35020 21788
rect 35020 21732 35076 21788
rect 35076 21732 35080 21788
rect 35016 21728 35080 21732
rect 35096 21788 35160 21792
rect 35096 21732 35100 21788
rect 35100 21732 35156 21788
rect 35156 21732 35160 21788
rect 35096 21728 35160 21732
rect 35176 21788 35240 21792
rect 35176 21732 35180 21788
rect 35180 21732 35236 21788
rect 35236 21732 35240 21788
rect 35176 21728 35240 21732
rect 19576 21244 19640 21248
rect 19576 21188 19580 21244
rect 19580 21188 19636 21244
rect 19636 21188 19640 21244
rect 19576 21184 19640 21188
rect 19656 21244 19720 21248
rect 19656 21188 19660 21244
rect 19660 21188 19716 21244
rect 19716 21188 19720 21244
rect 19656 21184 19720 21188
rect 19736 21244 19800 21248
rect 19736 21188 19740 21244
rect 19740 21188 19796 21244
rect 19796 21188 19800 21244
rect 19736 21184 19800 21188
rect 19816 21244 19880 21248
rect 19816 21188 19820 21244
rect 19820 21188 19876 21244
rect 19876 21188 19880 21244
rect 19816 21184 19880 21188
rect 4216 20700 4280 20704
rect 4216 20644 4220 20700
rect 4220 20644 4276 20700
rect 4276 20644 4280 20700
rect 4216 20640 4280 20644
rect 4296 20700 4360 20704
rect 4296 20644 4300 20700
rect 4300 20644 4356 20700
rect 4356 20644 4360 20700
rect 4296 20640 4360 20644
rect 4376 20700 4440 20704
rect 4376 20644 4380 20700
rect 4380 20644 4436 20700
rect 4436 20644 4440 20700
rect 4376 20640 4440 20644
rect 4456 20700 4520 20704
rect 4456 20644 4460 20700
rect 4460 20644 4516 20700
rect 4516 20644 4520 20700
rect 4456 20640 4520 20644
rect 34936 20700 35000 20704
rect 34936 20644 34940 20700
rect 34940 20644 34996 20700
rect 34996 20644 35000 20700
rect 34936 20640 35000 20644
rect 35016 20700 35080 20704
rect 35016 20644 35020 20700
rect 35020 20644 35076 20700
rect 35076 20644 35080 20700
rect 35016 20640 35080 20644
rect 35096 20700 35160 20704
rect 35096 20644 35100 20700
rect 35100 20644 35156 20700
rect 35156 20644 35160 20700
rect 35096 20640 35160 20644
rect 35176 20700 35240 20704
rect 35176 20644 35180 20700
rect 35180 20644 35236 20700
rect 35236 20644 35240 20700
rect 35176 20640 35240 20644
rect 19576 20156 19640 20160
rect 19576 20100 19580 20156
rect 19580 20100 19636 20156
rect 19636 20100 19640 20156
rect 19576 20096 19640 20100
rect 19656 20156 19720 20160
rect 19656 20100 19660 20156
rect 19660 20100 19716 20156
rect 19716 20100 19720 20156
rect 19656 20096 19720 20100
rect 19736 20156 19800 20160
rect 19736 20100 19740 20156
rect 19740 20100 19796 20156
rect 19796 20100 19800 20156
rect 19736 20096 19800 20100
rect 19816 20156 19880 20160
rect 19816 20100 19820 20156
rect 19820 20100 19876 20156
rect 19876 20100 19880 20156
rect 19816 20096 19880 20100
rect 4216 19612 4280 19616
rect 4216 19556 4220 19612
rect 4220 19556 4276 19612
rect 4276 19556 4280 19612
rect 4216 19552 4280 19556
rect 4296 19612 4360 19616
rect 4296 19556 4300 19612
rect 4300 19556 4356 19612
rect 4356 19556 4360 19612
rect 4296 19552 4360 19556
rect 4376 19612 4440 19616
rect 4376 19556 4380 19612
rect 4380 19556 4436 19612
rect 4436 19556 4440 19612
rect 4376 19552 4440 19556
rect 4456 19612 4520 19616
rect 4456 19556 4460 19612
rect 4460 19556 4516 19612
rect 4516 19556 4520 19612
rect 4456 19552 4520 19556
rect 34936 19612 35000 19616
rect 34936 19556 34940 19612
rect 34940 19556 34996 19612
rect 34996 19556 35000 19612
rect 34936 19552 35000 19556
rect 35016 19612 35080 19616
rect 35016 19556 35020 19612
rect 35020 19556 35076 19612
rect 35076 19556 35080 19612
rect 35016 19552 35080 19556
rect 35096 19612 35160 19616
rect 35096 19556 35100 19612
rect 35100 19556 35156 19612
rect 35156 19556 35160 19612
rect 35096 19552 35160 19556
rect 35176 19612 35240 19616
rect 35176 19556 35180 19612
rect 35180 19556 35236 19612
rect 35236 19556 35240 19612
rect 35176 19552 35240 19556
rect 19576 19068 19640 19072
rect 19576 19012 19580 19068
rect 19580 19012 19636 19068
rect 19636 19012 19640 19068
rect 19576 19008 19640 19012
rect 19656 19068 19720 19072
rect 19656 19012 19660 19068
rect 19660 19012 19716 19068
rect 19716 19012 19720 19068
rect 19656 19008 19720 19012
rect 19736 19068 19800 19072
rect 19736 19012 19740 19068
rect 19740 19012 19796 19068
rect 19796 19012 19800 19068
rect 19736 19008 19800 19012
rect 19816 19068 19880 19072
rect 19816 19012 19820 19068
rect 19820 19012 19876 19068
rect 19876 19012 19880 19068
rect 19816 19008 19880 19012
rect 4216 18524 4280 18528
rect 4216 18468 4220 18524
rect 4220 18468 4276 18524
rect 4276 18468 4280 18524
rect 4216 18464 4280 18468
rect 4296 18524 4360 18528
rect 4296 18468 4300 18524
rect 4300 18468 4356 18524
rect 4356 18468 4360 18524
rect 4296 18464 4360 18468
rect 4376 18524 4440 18528
rect 4376 18468 4380 18524
rect 4380 18468 4436 18524
rect 4436 18468 4440 18524
rect 4376 18464 4440 18468
rect 4456 18524 4520 18528
rect 4456 18468 4460 18524
rect 4460 18468 4516 18524
rect 4516 18468 4520 18524
rect 4456 18464 4520 18468
rect 34936 18524 35000 18528
rect 34936 18468 34940 18524
rect 34940 18468 34996 18524
rect 34996 18468 35000 18524
rect 34936 18464 35000 18468
rect 35016 18524 35080 18528
rect 35016 18468 35020 18524
rect 35020 18468 35076 18524
rect 35076 18468 35080 18524
rect 35016 18464 35080 18468
rect 35096 18524 35160 18528
rect 35096 18468 35100 18524
rect 35100 18468 35156 18524
rect 35156 18468 35160 18524
rect 35096 18464 35160 18468
rect 35176 18524 35240 18528
rect 35176 18468 35180 18524
rect 35180 18468 35236 18524
rect 35236 18468 35240 18524
rect 35176 18464 35240 18468
rect 19576 17980 19640 17984
rect 19576 17924 19580 17980
rect 19580 17924 19636 17980
rect 19636 17924 19640 17980
rect 19576 17920 19640 17924
rect 19656 17980 19720 17984
rect 19656 17924 19660 17980
rect 19660 17924 19716 17980
rect 19716 17924 19720 17980
rect 19656 17920 19720 17924
rect 19736 17980 19800 17984
rect 19736 17924 19740 17980
rect 19740 17924 19796 17980
rect 19796 17924 19800 17980
rect 19736 17920 19800 17924
rect 19816 17980 19880 17984
rect 19816 17924 19820 17980
rect 19820 17924 19876 17980
rect 19876 17924 19880 17980
rect 19816 17920 19880 17924
rect 4216 17436 4280 17440
rect 4216 17380 4220 17436
rect 4220 17380 4276 17436
rect 4276 17380 4280 17436
rect 4216 17376 4280 17380
rect 4296 17436 4360 17440
rect 4296 17380 4300 17436
rect 4300 17380 4356 17436
rect 4356 17380 4360 17436
rect 4296 17376 4360 17380
rect 4376 17436 4440 17440
rect 4376 17380 4380 17436
rect 4380 17380 4436 17436
rect 4436 17380 4440 17436
rect 4376 17376 4440 17380
rect 4456 17436 4520 17440
rect 4456 17380 4460 17436
rect 4460 17380 4516 17436
rect 4516 17380 4520 17436
rect 4456 17376 4520 17380
rect 34936 17436 35000 17440
rect 34936 17380 34940 17436
rect 34940 17380 34996 17436
rect 34996 17380 35000 17436
rect 34936 17376 35000 17380
rect 35016 17436 35080 17440
rect 35016 17380 35020 17436
rect 35020 17380 35076 17436
rect 35076 17380 35080 17436
rect 35016 17376 35080 17380
rect 35096 17436 35160 17440
rect 35096 17380 35100 17436
rect 35100 17380 35156 17436
rect 35156 17380 35160 17436
rect 35096 17376 35160 17380
rect 35176 17436 35240 17440
rect 35176 17380 35180 17436
rect 35180 17380 35236 17436
rect 35236 17380 35240 17436
rect 35176 17376 35240 17380
rect 19576 16892 19640 16896
rect 19576 16836 19580 16892
rect 19580 16836 19636 16892
rect 19636 16836 19640 16892
rect 19576 16832 19640 16836
rect 19656 16892 19720 16896
rect 19656 16836 19660 16892
rect 19660 16836 19716 16892
rect 19716 16836 19720 16892
rect 19656 16832 19720 16836
rect 19736 16892 19800 16896
rect 19736 16836 19740 16892
rect 19740 16836 19796 16892
rect 19796 16836 19800 16892
rect 19736 16832 19800 16836
rect 19816 16892 19880 16896
rect 19816 16836 19820 16892
rect 19820 16836 19876 16892
rect 19876 16836 19880 16892
rect 19816 16832 19880 16836
rect 4216 16348 4280 16352
rect 4216 16292 4220 16348
rect 4220 16292 4276 16348
rect 4276 16292 4280 16348
rect 4216 16288 4280 16292
rect 4296 16348 4360 16352
rect 4296 16292 4300 16348
rect 4300 16292 4356 16348
rect 4356 16292 4360 16348
rect 4296 16288 4360 16292
rect 4376 16348 4440 16352
rect 4376 16292 4380 16348
rect 4380 16292 4436 16348
rect 4436 16292 4440 16348
rect 4376 16288 4440 16292
rect 4456 16348 4520 16352
rect 4456 16292 4460 16348
rect 4460 16292 4516 16348
rect 4516 16292 4520 16348
rect 4456 16288 4520 16292
rect 34936 16348 35000 16352
rect 34936 16292 34940 16348
rect 34940 16292 34996 16348
rect 34996 16292 35000 16348
rect 34936 16288 35000 16292
rect 35016 16348 35080 16352
rect 35016 16292 35020 16348
rect 35020 16292 35076 16348
rect 35076 16292 35080 16348
rect 35016 16288 35080 16292
rect 35096 16348 35160 16352
rect 35096 16292 35100 16348
rect 35100 16292 35156 16348
rect 35156 16292 35160 16348
rect 35096 16288 35160 16292
rect 35176 16348 35240 16352
rect 35176 16292 35180 16348
rect 35180 16292 35236 16348
rect 35236 16292 35240 16348
rect 35176 16288 35240 16292
rect 19576 15804 19640 15808
rect 19576 15748 19580 15804
rect 19580 15748 19636 15804
rect 19636 15748 19640 15804
rect 19576 15744 19640 15748
rect 19656 15804 19720 15808
rect 19656 15748 19660 15804
rect 19660 15748 19716 15804
rect 19716 15748 19720 15804
rect 19656 15744 19720 15748
rect 19736 15804 19800 15808
rect 19736 15748 19740 15804
rect 19740 15748 19796 15804
rect 19796 15748 19800 15804
rect 19736 15744 19800 15748
rect 19816 15804 19880 15808
rect 19816 15748 19820 15804
rect 19820 15748 19876 15804
rect 19876 15748 19880 15804
rect 19816 15744 19880 15748
rect 4216 15260 4280 15264
rect 4216 15204 4220 15260
rect 4220 15204 4276 15260
rect 4276 15204 4280 15260
rect 4216 15200 4280 15204
rect 4296 15260 4360 15264
rect 4296 15204 4300 15260
rect 4300 15204 4356 15260
rect 4356 15204 4360 15260
rect 4296 15200 4360 15204
rect 4376 15260 4440 15264
rect 4376 15204 4380 15260
rect 4380 15204 4436 15260
rect 4436 15204 4440 15260
rect 4376 15200 4440 15204
rect 4456 15260 4520 15264
rect 4456 15204 4460 15260
rect 4460 15204 4516 15260
rect 4516 15204 4520 15260
rect 4456 15200 4520 15204
rect 34936 15260 35000 15264
rect 34936 15204 34940 15260
rect 34940 15204 34996 15260
rect 34996 15204 35000 15260
rect 34936 15200 35000 15204
rect 35016 15260 35080 15264
rect 35016 15204 35020 15260
rect 35020 15204 35076 15260
rect 35076 15204 35080 15260
rect 35016 15200 35080 15204
rect 35096 15260 35160 15264
rect 35096 15204 35100 15260
rect 35100 15204 35156 15260
rect 35156 15204 35160 15260
rect 35096 15200 35160 15204
rect 35176 15260 35240 15264
rect 35176 15204 35180 15260
rect 35180 15204 35236 15260
rect 35236 15204 35240 15260
rect 35176 15200 35240 15204
rect 19576 14716 19640 14720
rect 19576 14660 19580 14716
rect 19580 14660 19636 14716
rect 19636 14660 19640 14716
rect 19576 14656 19640 14660
rect 19656 14716 19720 14720
rect 19656 14660 19660 14716
rect 19660 14660 19716 14716
rect 19716 14660 19720 14716
rect 19656 14656 19720 14660
rect 19736 14716 19800 14720
rect 19736 14660 19740 14716
rect 19740 14660 19796 14716
rect 19796 14660 19800 14716
rect 19736 14656 19800 14660
rect 19816 14716 19880 14720
rect 19816 14660 19820 14716
rect 19820 14660 19876 14716
rect 19876 14660 19880 14716
rect 19816 14656 19880 14660
rect 4216 14172 4280 14176
rect 4216 14116 4220 14172
rect 4220 14116 4276 14172
rect 4276 14116 4280 14172
rect 4216 14112 4280 14116
rect 4296 14172 4360 14176
rect 4296 14116 4300 14172
rect 4300 14116 4356 14172
rect 4356 14116 4360 14172
rect 4296 14112 4360 14116
rect 4376 14172 4440 14176
rect 4376 14116 4380 14172
rect 4380 14116 4436 14172
rect 4436 14116 4440 14172
rect 4376 14112 4440 14116
rect 4456 14172 4520 14176
rect 4456 14116 4460 14172
rect 4460 14116 4516 14172
rect 4516 14116 4520 14172
rect 4456 14112 4520 14116
rect 34936 14172 35000 14176
rect 34936 14116 34940 14172
rect 34940 14116 34996 14172
rect 34996 14116 35000 14172
rect 34936 14112 35000 14116
rect 35016 14172 35080 14176
rect 35016 14116 35020 14172
rect 35020 14116 35076 14172
rect 35076 14116 35080 14172
rect 35016 14112 35080 14116
rect 35096 14172 35160 14176
rect 35096 14116 35100 14172
rect 35100 14116 35156 14172
rect 35156 14116 35160 14172
rect 35096 14112 35160 14116
rect 35176 14172 35240 14176
rect 35176 14116 35180 14172
rect 35180 14116 35236 14172
rect 35236 14116 35240 14172
rect 35176 14112 35240 14116
rect 19576 13628 19640 13632
rect 19576 13572 19580 13628
rect 19580 13572 19636 13628
rect 19636 13572 19640 13628
rect 19576 13568 19640 13572
rect 19656 13628 19720 13632
rect 19656 13572 19660 13628
rect 19660 13572 19716 13628
rect 19716 13572 19720 13628
rect 19656 13568 19720 13572
rect 19736 13628 19800 13632
rect 19736 13572 19740 13628
rect 19740 13572 19796 13628
rect 19796 13572 19800 13628
rect 19736 13568 19800 13572
rect 19816 13628 19880 13632
rect 19816 13572 19820 13628
rect 19820 13572 19876 13628
rect 19876 13572 19880 13628
rect 19816 13568 19880 13572
rect 4216 13084 4280 13088
rect 4216 13028 4220 13084
rect 4220 13028 4276 13084
rect 4276 13028 4280 13084
rect 4216 13024 4280 13028
rect 4296 13084 4360 13088
rect 4296 13028 4300 13084
rect 4300 13028 4356 13084
rect 4356 13028 4360 13084
rect 4296 13024 4360 13028
rect 4376 13084 4440 13088
rect 4376 13028 4380 13084
rect 4380 13028 4436 13084
rect 4436 13028 4440 13084
rect 4376 13024 4440 13028
rect 4456 13084 4520 13088
rect 4456 13028 4460 13084
rect 4460 13028 4516 13084
rect 4516 13028 4520 13084
rect 4456 13024 4520 13028
rect 34936 13084 35000 13088
rect 34936 13028 34940 13084
rect 34940 13028 34996 13084
rect 34996 13028 35000 13084
rect 34936 13024 35000 13028
rect 35016 13084 35080 13088
rect 35016 13028 35020 13084
rect 35020 13028 35076 13084
rect 35076 13028 35080 13084
rect 35016 13024 35080 13028
rect 35096 13084 35160 13088
rect 35096 13028 35100 13084
rect 35100 13028 35156 13084
rect 35156 13028 35160 13084
rect 35096 13024 35160 13028
rect 35176 13084 35240 13088
rect 35176 13028 35180 13084
rect 35180 13028 35236 13084
rect 35236 13028 35240 13084
rect 35176 13024 35240 13028
rect 19576 12540 19640 12544
rect 19576 12484 19580 12540
rect 19580 12484 19636 12540
rect 19636 12484 19640 12540
rect 19576 12480 19640 12484
rect 19656 12540 19720 12544
rect 19656 12484 19660 12540
rect 19660 12484 19716 12540
rect 19716 12484 19720 12540
rect 19656 12480 19720 12484
rect 19736 12540 19800 12544
rect 19736 12484 19740 12540
rect 19740 12484 19796 12540
rect 19796 12484 19800 12540
rect 19736 12480 19800 12484
rect 19816 12540 19880 12544
rect 19816 12484 19820 12540
rect 19820 12484 19876 12540
rect 19876 12484 19880 12540
rect 19816 12480 19880 12484
rect 4216 11996 4280 12000
rect 4216 11940 4220 11996
rect 4220 11940 4276 11996
rect 4276 11940 4280 11996
rect 4216 11936 4280 11940
rect 4296 11996 4360 12000
rect 4296 11940 4300 11996
rect 4300 11940 4356 11996
rect 4356 11940 4360 11996
rect 4296 11936 4360 11940
rect 4376 11996 4440 12000
rect 4376 11940 4380 11996
rect 4380 11940 4436 11996
rect 4436 11940 4440 11996
rect 4376 11936 4440 11940
rect 4456 11996 4520 12000
rect 4456 11940 4460 11996
rect 4460 11940 4516 11996
rect 4516 11940 4520 11996
rect 4456 11936 4520 11940
rect 34936 11996 35000 12000
rect 34936 11940 34940 11996
rect 34940 11940 34996 11996
rect 34996 11940 35000 11996
rect 34936 11936 35000 11940
rect 35016 11996 35080 12000
rect 35016 11940 35020 11996
rect 35020 11940 35076 11996
rect 35076 11940 35080 11996
rect 35016 11936 35080 11940
rect 35096 11996 35160 12000
rect 35096 11940 35100 11996
rect 35100 11940 35156 11996
rect 35156 11940 35160 11996
rect 35096 11936 35160 11940
rect 35176 11996 35240 12000
rect 35176 11940 35180 11996
rect 35180 11940 35236 11996
rect 35236 11940 35240 11996
rect 35176 11936 35240 11940
rect 19576 11452 19640 11456
rect 19576 11396 19580 11452
rect 19580 11396 19636 11452
rect 19636 11396 19640 11452
rect 19576 11392 19640 11396
rect 19656 11452 19720 11456
rect 19656 11396 19660 11452
rect 19660 11396 19716 11452
rect 19716 11396 19720 11452
rect 19656 11392 19720 11396
rect 19736 11452 19800 11456
rect 19736 11396 19740 11452
rect 19740 11396 19796 11452
rect 19796 11396 19800 11452
rect 19736 11392 19800 11396
rect 19816 11452 19880 11456
rect 19816 11396 19820 11452
rect 19820 11396 19876 11452
rect 19876 11396 19880 11452
rect 19816 11392 19880 11396
rect 4216 10908 4280 10912
rect 4216 10852 4220 10908
rect 4220 10852 4276 10908
rect 4276 10852 4280 10908
rect 4216 10848 4280 10852
rect 4296 10908 4360 10912
rect 4296 10852 4300 10908
rect 4300 10852 4356 10908
rect 4356 10852 4360 10908
rect 4296 10848 4360 10852
rect 4376 10908 4440 10912
rect 4376 10852 4380 10908
rect 4380 10852 4436 10908
rect 4436 10852 4440 10908
rect 4376 10848 4440 10852
rect 4456 10908 4520 10912
rect 4456 10852 4460 10908
rect 4460 10852 4516 10908
rect 4516 10852 4520 10908
rect 4456 10848 4520 10852
rect 34936 10908 35000 10912
rect 34936 10852 34940 10908
rect 34940 10852 34996 10908
rect 34996 10852 35000 10908
rect 34936 10848 35000 10852
rect 35016 10908 35080 10912
rect 35016 10852 35020 10908
rect 35020 10852 35076 10908
rect 35076 10852 35080 10908
rect 35016 10848 35080 10852
rect 35096 10908 35160 10912
rect 35096 10852 35100 10908
rect 35100 10852 35156 10908
rect 35156 10852 35160 10908
rect 35096 10848 35160 10852
rect 35176 10908 35240 10912
rect 35176 10852 35180 10908
rect 35180 10852 35236 10908
rect 35236 10852 35240 10908
rect 35176 10848 35240 10852
rect 19576 10364 19640 10368
rect 19576 10308 19580 10364
rect 19580 10308 19636 10364
rect 19636 10308 19640 10364
rect 19576 10304 19640 10308
rect 19656 10364 19720 10368
rect 19656 10308 19660 10364
rect 19660 10308 19716 10364
rect 19716 10308 19720 10364
rect 19656 10304 19720 10308
rect 19736 10364 19800 10368
rect 19736 10308 19740 10364
rect 19740 10308 19796 10364
rect 19796 10308 19800 10364
rect 19736 10304 19800 10308
rect 19816 10364 19880 10368
rect 19816 10308 19820 10364
rect 19820 10308 19876 10364
rect 19876 10308 19880 10364
rect 19816 10304 19880 10308
rect 4216 9820 4280 9824
rect 4216 9764 4220 9820
rect 4220 9764 4276 9820
rect 4276 9764 4280 9820
rect 4216 9760 4280 9764
rect 4296 9820 4360 9824
rect 4296 9764 4300 9820
rect 4300 9764 4356 9820
rect 4356 9764 4360 9820
rect 4296 9760 4360 9764
rect 4376 9820 4440 9824
rect 4376 9764 4380 9820
rect 4380 9764 4436 9820
rect 4436 9764 4440 9820
rect 4376 9760 4440 9764
rect 4456 9820 4520 9824
rect 4456 9764 4460 9820
rect 4460 9764 4516 9820
rect 4516 9764 4520 9820
rect 4456 9760 4520 9764
rect 34936 9820 35000 9824
rect 34936 9764 34940 9820
rect 34940 9764 34996 9820
rect 34996 9764 35000 9820
rect 34936 9760 35000 9764
rect 35016 9820 35080 9824
rect 35016 9764 35020 9820
rect 35020 9764 35076 9820
rect 35076 9764 35080 9820
rect 35016 9760 35080 9764
rect 35096 9820 35160 9824
rect 35096 9764 35100 9820
rect 35100 9764 35156 9820
rect 35156 9764 35160 9820
rect 35096 9760 35160 9764
rect 35176 9820 35240 9824
rect 35176 9764 35180 9820
rect 35180 9764 35236 9820
rect 35236 9764 35240 9820
rect 35176 9760 35240 9764
rect 19576 9276 19640 9280
rect 19576 9220 19580 9276
rect 19580 9220 19636 9276
rect 19636 9220 19640 9276
rect 19576 9216 19640 9220
rect 19656 9276 19720 9280
rect 19656 9220 19660 9276
rect 19660 9220 19716 9276
rect 19716 9220 19720 9276
rect 19656 9216 19720 9220
rect 19736 9276 19800 9280
rect 19736 9220 19740 9276
rect 19740 9220 19796 9276
rect 19796 9220 19800 9276
rect 19736 9216 19800 9220
rect 19816 9276 19880 9280
rect 19816 9220 19820 9276
rect 19820 9220 19876 9276
rect 19876 9220 19880 9276
rect 19816 9216 19880 9220
rect 4216 8732 4280 8736
rect 4216 8676 4220 8732
rect 4220 8676 4276 8732
rect 4276 8676 4280 8732
rect 4216 8672 4280 8676
rect 4296 8732 4360 8736
rect 4296 8676 4300 8732
rect 4300 8676 4356 8732
rect 4356 8676 4360 8732
rect 4296 8672 4360 8676
rect 4376 8732 4440 8736
rect 4376 8676 4380 8732
rect 4380 8676 4436 8732
rect 4436 8676 4440 8732
rect 4376 8672 4440 8676
rect 4456 8732 4520 8736
rect 4456 8676 4460 8732
rect 4460 8676 4516 8732
rect 4516 8676 4520 8732
rect 4456 8672 4520 8676
rect 34936 8732 35000 8736
rect 34936 8676 34940 8732
rect 34940 8676 34996 8732
rect 34996 8676 35000 8732
rect 34936 8672 35000 8676
rect 35016 8732 35080 8736
rect 35016 8676 35020 8732
rect 35020 8676 35076 8732
rect 35076 8676 35080 8732
rect 35016 8672 35080 8676
rect 35096 8732 35160 8736
rect 35096 8676 35100 8732
rect 35100 8676 35156 8732
rect 35156 8676 35160 8732
rect 35096 8672 35160 8676
rect 35176 8732 35240 8736
rect 35176 8676 35180 8732
rect 35180 8676 35236 8732
rect 35236 8676 35240 8732
rect 35176 8672 35240 8676
rect 19576 8188 19640 8192
rect 19576 8132 19580 8188
rect 19580 8132 19636 8188
rect 19636 8132 19640 8188
rect 19576 8128 19640 8132
rect 19656 8188 19720 8192
rect 19656 8132 19660 8188
rect 19660 8132 19716 8188
rect 19716 8132 19720 8188
rect 19656 8128 19720 8132
rect 19736 8188 19800 8192
rect 19736 8132 19740 8188
rect 19740 8132 19796 8188
rect 19796 8132 19800 8188
rect 19736 8128 19800 8132
rect 19816 8188 19880 8192
rect 19816 8132 19820 8188
rect 19820 8132 19876 8188
rect 19876 8132 19880 8188
rect 19816 8128 19880 8132
rect 4216 7644 4280 7648
rect 4216 7588 4220 7644
rect 4220 7588 4276 7644
rect 4276 7588 4280 7644
rect 4216 7584 4280 7588
rect 4296 7644 4360 7648
rect 4296 7588 4300 7644
rect 4300 7588 4356 7644
rect 4356 7588 4360 7644
rect 4296 7584 4360 7588
rect 4376 7644 4440 7648
rect 4376 7588 4380 7644
rect 4380 7588 4436 7644
rect 4436 7588 4440 7644
rect 4376 7584 4440 7588
rect 4456 7644 4520 7648
rect 4456 7588 4460 7644
rect 4460 7588 4516 7644
rect 4516 7588 4520 7644
rect 4456 7584 4520 7588
rect 34936 7644 35000 7648
rect 34936 7588 34940 7644
rect 34940 7588 34996 7644
rect 34996 7588 35000 7644
rect 34936 7584 35000 7588
rect 35016 7644 35080 7648
rect 35016 7588 35020 7644
rect 35020 7588 35076 7644
rect 35076 7588 35080 7644
rect 35016 7584 35080 7588
rect 35096 7644 35160 7648
rect 35096 7588 35100 7644
rect 35100 7588 35156 7644
rect 35156 7588 35160 7644
rect 35096 7584 35160 7588
rect 35176 7644 35240 7648
rect 35176 7588 35180 7644
rect 35180 7588 35236 7644
rect 35236 7588 35240 7644
rect 35176 7584 35240 7588
rect 19576 7100 19640 7104
rect 19576 7044 19580 7100
rect 19580 7044 19636 7100
rect 19636 7044 19640 7100
rect 19576 7040 19640 7044
rect 19656 7100 19720 7104
rect 19656 7044 19660 7100
rect 19660 7044 19716 7100
rect 19716 7044 19720 7100
rect 19656 7040 19720 7044
rect 19736 7100 19800 7104
rect 19736 7044 19740 7100
rect 19740 7044 19796 7100
rect 19796 7044 19800 7100
rect 19736 7040 19800 7044
rect 19816 7100 19880 7104
rect 19816 7044 19820 7100
rect 19820 7044 19876 7100
rect 19876 7044 19880 7100
rect 19816 7040 19880 7044
rect 4216 6556 4280 6560
rect 4216 6500 4220 6556
rect 4220 6500 4276 6556
rect 4276 6500 4280 6556
rect 4216 6496 4280 6500
rect 4296 6556 4360 6560
rect 4296 6500 4300 6556
rect 4300 6500 4356 6556
rect 4356 6500 4360 6556
rect 4296 6496 4360 6500
rect 4376 6556 4440 6560
rect 4376 6500 4380 6556
rect 4380 6500 4436 6556
rect 4436 6500 4440 6556
rect 4376 6496 4440 6500
rect 4456 6556 4520 6560
rect 4456 6500 4460 6556
rect 4460 6500 4516 6556
rect 4516 6500 4520 6556
rect 4456 6496 4520 6500
rect 34936 6556 35000 6560
rect 34936 6500 34940 6556
rect 34940 6500 34996 6556
rect 34996 6500 35000 6556
rect 34936 6496 35000 6500
rect 35016 6556 35080 6560
rect 35016 6500 35020 6556
rect 35020 6500 35076 6556
rect 35076 6500 35080 6556
rect 35016 6496 35080 6500
rect 35096 6556 35160 6560
rect 35096 6500 35100 6556
rect 35100 6500 35156 6556
rect 35156 6500 35160 6556
rect 35096 6496 35160 6500
rect 35176 6556 35240 6560
rect 35176 6500 35180 6556
rect 35180 6500 35236 6556
rect 35236 6500 35240 6556
rect 35176 6496 35240 6500
rect 19576 6012 19640 6016
rect 19576 5956 19580 6012
rect 19580 5956 19636 6012
rect 19636 5956 19640 6012
rect 19576 5952 19640 5956
rect 19656 6012 19720 6016
rect 19656 5956 19660 6012
rect 19660 5956 19716 6012
rect 19716 5956 19720 6012
rect 19656 5952 19720 5956
rect 19736 6012 19800 6016
rect 19736 5956 19740 6012
rect 19740 5956 19796 6012
rect 19796 5956 19800 6012
rect 19736 5952 19800 5956
rect 19816 6012 19880 6016
rect 19816 5956 19820 6012
rect 19820 5956 19876 6012
rect 19876 5956 19880 6012
rect 19816 5952 19880 5956
rect 4216 5468 4280 5472
rect 4216 5412 4220 5468
rect 4220 5412 4276 5468
rect 4276 5412 4280 5468
rect 4216 5408 4280 5412
rect 4296 5468 4360 5472
rect 4296 5412 4300 5468
rect 4300 5412 4356 5468
rect 4356 5412 4360 5468
rect 4296 5408 4360 5412
rect 4376 5468 4440 5472
rect 4376 5412 4380 5468
rect 4380 5412 4436 5468
rect 4436 5412 4440 5468
rect 4376 5408 4440 5412
rect 4456 5468 4520 5472
rect 4456 5412 4460 5468
rect 4460 5412 4516 5468
rect 4516 5412 4520 5468
rect 4456 5408 4520 5412
rect 34936 5468 35000 5472
rect 34936 5412 34940 5468
rect 34940 5412 34996 5468
rect 34996 5412 35000 5468
rect 34936 5408 35000 5412
rect 35016 5468 35080 5472
rect 35016 5412 35020 5468
rect 35020 5412 35076 5468
rect 35076 5412 35080 5468
rect 35016 5408 35080 5412
rect 35096 5468 35160 5472
rect 35096 5412 35100 5468
rect 35100 5412 35156 5468
rect 35156 5412 35160 5468
rect 35096 5408 35160 5412
rect 35176 5468 35240 5472
rect 35176 5412 35180 5468
rect 35180 5412 35236 5468
rect 35236 5412 35240 5468
rect 35176 5408 35240 5412
rect 19576 4924 19640 4928
rect 19576 4868 19580 4924
rect 19580 4868 19636 4924
rect 19636 4868 19640 4924
rect 19576 4864 19640 4868
rect 19656 4924 19720 4928
rect 19656 4868 19660 4924
rect 19660 4868 19716 4924
rect 19716 4868 19720 4924
rect 19656 4864 19720 4868
rect 19736 4924 19800 4928
rect 19736 4868 19740 4924
rect 19740 4868 19796 4924
rect 19796 4868 19800 4924
rect 19736 4864 19800 4868
rect 19816 4924 19880 4928
rect 19816 4868 19820 4924
rect 19820 4868 19876 4924
rect 19876 4868 19880 4924
rect 19816 4864 19880 4868
rect 4216 4380 4280 4384
rect 4216 4324 4220 4380
rect 4220 4324 4276 4380
rect 4276 4324 4280 4380
rect 4216 4320 4280 4324
rect 4296 4380 4360 4384
rect 4296 4324 4300 4380
rect 4300 4324 4356 4380
rect 4356 4324 4360 4380
rect 4296 4320 4360 4324
rect 4376 4380 4440 4384
rect 4376 4324 4380 4380
rect 4380 4324 4436 4380
rect 4436 4324 4440 4380
rect 4376 4320 4440 4324
rect 4456 4380 4520 4384
rect 4456 4324 4460 4380
rect 4460 4324 4516 4380
rect 4516 4324 4520 4380
rect 4456 4320 4520 4324
rect 34936 4380 35000 4384
rect 34936 4324 34940 4380
rect 34940 4324 34996 4380
rect 34996 4324 35000 4380
rect 34936 4320 35000 4324
rect 35016 4380 35080 4384
rect 35016 4324 35020 4380
rect 35020 4324 35076 4380
rect 35076 4324 35080 4380
rect 35016 4320 35080 4324
rect 35096 4380 35160 4384
rect 35096 4324 35100 4380
rect 35100 4324 35156 4380
rect 35156 4324 35160 4380
rect 35096 4320 35160 4324
rect 35176 4380 35240 4384
rect 35176 4324 35180 4380
rect 35180 4324 35236 4380
rect 35236 4324 35240 4380
rect 35176 4320 35240 4324
rect 19576 3836 19640 3840
rect 19576 3780 19580 3836
rect 19580 3780 19636 3836
rect 19636 3780 19640 3836
rect 19576 3776 19640 3780
rect 19656 3836 19720 3840
rect 19656 3780 19660 3836
rect 19660 3780 19716 3836
rect 19716 3780 19720 3836
rect 19656 3776 19720 3780
rect 19736 3836 19800 3840
rect 19736 3780 19740 3836
rect 19740 3780 19796 3836
rect 19796 3780 19800 3836
rect 19736 3776 19800 3780
rect 19816 3836 19880 3840
rect 19816 3780 19820 3836
rect 19820 3780 19876 3836
rect 19876 3780 19880 3836
rect 19816 3776 19880 3780
rect 4216 3292 4280 3296
rect 4216 3236 4220 3292
rect 4220 3236 4276 3292
rect 4276 3236 4280 3292
rect 4216 3232 4280 3236
rect 4296 3292 4360 3296
rect 4296 3236 4300 3292
rect 4300 3236 4356 3292
rect 4356 3236 4360 3292
rect 4296 3232 4360 3236
rect 4376 3292 4440 3296
rect 4376 3236 4380 3292
rect 4380 3236 4436 3292
rect 4436 3236 4440 3292
rect 4376 3232 4440 3236
rect 4456 3292 4520 3296
rect 4456 3236 4460 3292
rect 4460 3236 4516 3292
rect 4516 3236 4520 3292
rect 4456 3232 4520 3236
rect 34936 3292 35000 3296
rect 34936 3236 34940 3292
rect 34940 3236 34996 3292
rect 34996 3236 35000 3292
rect 34936 3232 35000 3236
rect 35016 3292 35080 3296
rect 35016 3236 35020 3292
rect 35020 3236 35076 3292
rect 35076 3236 35080 3292
rect 35016 3232 35080 3236
rect 35096 3292 35160 3296
rect 35096 3236 35100 3292
rect 35100 3236 35156 3292
rect 35156 3236 35160 3292
rect 35096 3232 35160 3236
rect 35176 3292 35240 3296
rect 35176 3236 35180 3292
rect 35180 3236 35236 3292
rect 35236 3236 35240 3292
rect 35176 3232 35240 3236
rect 19576 2748 19640 2752
rect 19576 2692 19580 2748
rect 19580 2692 19636 2748
rect 19636 2692 19640 2748
rect 19576 2688 19640 2692
rect 19656 2748 19720 2752
rect 19656 2692 19660 2748
rect 19660 2692 19716 2748
rect 19716 2692 19720 2748
rect 19656 2688 19720 2692
rect 19736 2748 19800 2752
rect 19736 2692 19740 2748
rect 19740 2692 19796 2748
rect 19796 2692 19800 2748
rect 19736 2688 19800 2692
rect 19816 2748 19880 2752
rect 19816 2692 19820 2748
rect 19820 2692 19876 2748
rect 19876 2692 19880 2748
rect 19816 2688 19880 2692
rect 4216 2204 4280 2208
rect 4216 2148 4220 2204
rect 4220 2148 4276 2204
rect 4276 2148 4280 2204
rect 4216 2144 4280 2148
rect 4296 2204 4360 2208
rect 4296 2148 4300 2204
rect 4300 2148 4356 2204
rect 4356 2148 4360 2204
rect 4296 2144 4360 2148
rect 4376 2204 4440 2208
rect 4376 2148 4380 2204
rect 4380 2148 4436 2204
rect 4436 2148 4440 2204
rect 4376 2144 4440 2148
rect 4456 2204 4520 2208
rect 4456 2148 4460 2204
rect 4460 2148 4516 2204
rect 4516 2148 4520 2204
rect 4456 2144 4520 2148
rect 34936 2204 35000 2208
rect 34936 2148 34940 2204
rect 34940 2148 34996 2204
rect 34996 2148 35000 2204
rect 34936 2144 35000 2148
rect 35016 2204 35080 2208
rect 35016 2148 35020 2204
rect 35020 2148 35076 2204
rect 35076 2148 35080 2204
rect 35016 2144 35080 2148
rect 35096 2204 35160 2208
rect 35096 2148 35100 2204
rect 35100 2148 35156 2204
rect 35156 2148 35160 2204
rect 35096 2144 35160 2148
rect 35176 2204 35240 2208
rect 35176 2148 35180 2204
rect 35180 2148 35236 2204
rect 35236 2148 35240 2204
rect 35176 2144 35240 2148
<< metal4 >>
rect 4208 38112 4528 38672
rect 19568 38656 19888 38672
rect 4208 38048 4216 38112
rect 4280 38048 4296 38112
rect 4360 38048 4376 38112
rect 4440 38048 4456 38112
rect 4520 38048 4528 38112
rect 4208 37024 4528 38048
rect 4208 36960 4216 37024
rect 4280 36960 4296 37024
rect 4360 36960 4376 37024
rect 4440 36960 4456 37024
rect 4520 36960 4528 37024
rect 4208 35936 4528 36960
rect 4208 35872 4216 35936
rect 4280 35872 4296 35936
rect 4360 35872 4376 35936
rect 4440 35872 4456 35936
rect 4520 35872 4528 35936
rect 4208 34848 4528 35872
rect 4208 34784 4216 34848
rect 4280 34784 4296 34848
rect 4360 34784 4376 34848
rect 4440 34784 4456 34848
rect 4520 34784 4528 34848
rect 4208 33760 4528 34784
rect 4208 33696 4216 33760
rect 4280 33696 4296 33760
rect 4360 33696 4376 33760
rect 4440 33696 4456 33760
rect 4520 33696 4528 33760
rect 4208 32672 4528 33696
rect 4208 32608 4216 32672
rect 4280 32608 4296 32672
rect 4360 32608 4376 32672
rect 4440 32608 4456 32672
rect 4520 32608 4528 32672
rect 4208 31584 4528 32608
rect 4208 31520 4216 31584
rect 4280 31520 4296 31584
rect 4360 31520 4376 31584
rect 4440 31520 4456 31584
rect 4520 31520 4528 31584
rect 4208 30496 4528 31520
rect 4208 30432 4216 30496
rect 4280 30432 4296 30496
rect 4360 30432 4376 30496
rect 4440 30432 4456 30496
rect 4520 30432 4528 30496
rect 4208 29408 4528 30432
rect 4208 29344 4216 29408
rect 4280 29344 4296 29408
rect 4360 29344 4376 29408
rect 4440 29344 4456 29408
rect 4520 29344 4528 29408
rect 4208 28320 4528 29344
rect 4208 28256 4216 28320
rect 4280 28256 4296 28320
rect 4360 28256 4376 28320
rect 4440 28256 4456 28320
rect 4520 28256 4528 28320
rect 4208 27232 4528 28256
rect 4208 27168 4216 27232
rect 4280 27168 4296 27232
rect 4360 27168 4376 27232
rect 4440 27168 4456 27232
rect 4520 27168 4528 27232
rect 4208 26144 4528 27168
rect 4208 26080 4216 26144
rect 4280 26080 4296 26144
rect 4360 26080 4376 26144
rect 4440 26080 4456 26144
rect 4520 26080 4528 26144
rect 4208 25056 4528 26080
rect 4208 24992 4216 25056
rect 4280 24992 4296 25056
rect 4360 24992 4376 25056
rect 4440 24992 4456 25056
rect 4520 24992 4528 25056
rect 4208 23968 4528 24992
rect 4208 23904 4216 23968
rect 4280 23904 4296 23968
rect 4360 23904 4376 23968
rect 4440 23904 4456 23968
rect 4520 23904 4528 23968
rect 4208 22880 4528 23904
rect 4208 22816 4216 22880
rect 4280 22816 4296 22880
rect 4360 22816 4376 22880
rect 4440 22816 4456 22880
rect 4520 22816 4528 22880
rect 4208 21792 4528 22816
rect 4208 21728 4216 21792
rect 4280 21728 4296 21792
rect 4360 21728 4376 21792
rect 4440 21728 4456 21792
rect 4520 21728 4528 21792
rect 4208 20704 4528 21728
rect 4208 20640 4216 20704
rect 4280 20640 4296 20704
rect 4360 20640 4376 20704
rect 4440 20640 4456 20704
rect 4520 20640 4528 20704
rect 4208 19616 4528 20640
rect 4208 19552 4216 19616
rect 4280 19552 4296 19616
rect 4360 19552 4376 19616
rect 4440 19552 4456 19616
rect 4520 19552 4528 19616
rect 4208 18528 4528 19552
rect 4208 18464 4216 18528
rect 4280 18464 4296 18528
rect 4360 18464 4376 18528
rect 4440 18464 4456 18528
rect 4520 18464 4528 18528
rect 4208 17440 4528 18464
rect 4208 17376 4216 17440
rect 4280 17376 4296 17440
rect 4360 17376 4376 17440
rect 4440 17376 4456 17440
rect 4520 17376 4528 17440
rect 4208 16352 4528 17376
rect 4208 16288 4216 16352
rect 4280 16288 4296 16352
rect 4360 16288 4376 16352
rect 4440 16288 4456 16352
rect 4520 16288 4528 16352
rect 4208 15264 4528 16288
rect 4208 15200 4216 15264
rect 4280 15200 4296 15264
rect 4360 15200 4376 15264
rect 4440 15200 4456 15264
rect 4520 15200 4528 15264
rect 4208 14176 4528 15200
rect 4208 14112 4216 14176
rect 4280 14112 4296 14176
rect 4360 14112 4376 14176
rect 4440 14112 4456 14176
rect 4520 14112 4528 14176
rect 4208 13088 4528 14112
rect 4208 13024 4216 13088
rect 4280 13024 4296 13088
rect 4360 13024 4376 13088
rect 4440 13024 4456 13088
rect 4520 13024 4528 13088
rect 4208 12000 4528 13024
rect 4208 11936 4216 12000
rect 4280 11936 4296 12000
rect 4360 11936 4376 12000
rect 4440 11936 4456 12000
rect 4520 11936 4528 12000
rect 4208 10912 4528 11936
rect 4208 10848 4216 10912
rect 4280 10848 4296 10912
rect 4360 10848 4376 10912
rect 4440 10848 4456 10912
rect 4520 10848 4528 10912
rect 4208 9824 4528 10848
rect 4208 9760 4216 9824
rect 4280 9760 4296 9824
rect 4360 9760 4376 9824
rect 4440 9760 4456 9824
rect 4520 9760 4528 9824
rect 4208 8736 4528 9760
rect 4208 8672 4216 8736
rect 4280 8672 4296 8736
rect 4360 8672 4376 8736
rect 4440 8672 4456 8736
rect 4520 8672 4528 8736
rect 4208 7648 4528 8672
rect 4208 7584 4216 7648
rect 4280 7584 4296 7648
rect 4360 7584 4376 7648
rect 4440 7584 4456 7648
rect 4520 7584 4528 7648
rect 4208 6560 4528 7584
rect 4208 6496 4216 6560
rect 4280 6496 4296 6560
rect 4360 6496 4376 6560
rect 4440 6496 4456 6560
rect 4520 6496 4528 6560
rect 4208 5472 4528 6496
rect 4208 5408 4216 5472
rect 4280 5408 4296 5472
rect 4360 5408 4376 5472
rect 4440 5408 4456 5472
rect 4520 5408 4528 5472
rect 4208 4384 4528 5408
rect 4208 4320 4216 4384
rect 4280 4320 4296 4384
rect 4360 4320 4376 4384
rect 4440 4320 4456 4384
rect 4520 4320 4528 4384
rect 4208 3296 4528 4320
rect 4208 3232 4216 3296
rect 4280 3232 4296 3296
rect 4360 3232 4376 3296
rect 4440 3232 4456 3296
rect 4520 3232 4528 3296
rect 4208 2208 4528 3232
rect 4208 2144 4216 2208
rect 4280 2144 4296 2208
rect 4360 2144 4376 2208
rect 4440 2144 4456 2208
rect 4520 2144 4528 2208
rect 4868 2176 5188 38624
rect 5528 2176 5848 38624
rect 6188 2176 6508 38624
rect 19568 38592 19576 38656
rect 19640 38592 19656 38656
rect 19720 38592 19736 38656
rect 19800 38592 19816 38656
rect 19880 38592 19888 38656
rect 19568 37568 19888 38592
rect 19568 37504 19576 37568
rect 19640 37504 19656 37568
rect 19720 37504 19736 37568
rect 19800 37504 19816 37568
rect 19880 37504 19888 37568
rect 19568 36480 19888 37504
rect 19568 36416 19576 36480
rect 19640 36416 19656 36480
rect 19720 36416 19736 36480
rect 19800 36416 19816 36480
rect 19880 36416 19888 36480
rect 19568 35392 19888 36416
rect 19568 35328 19576 35392
rect 19640 35328 19656 35392
rect 19720 35328 19736 35392
rect 19800 35328 19816 35392
rect 19880 35328 19888 35392
rect 19568 34304 19888 35328
rect 19568 34240 19576 34304
rect 19640 34240 19656 34304
rect 19720 34240 19736 34304
rect 19800 34240 19816 34304
rect 19880 34240 19888 34304
rect 19568 33216 19888 34240
rect 19568 33152 19576 33216
rect 19640 33152 19656 33216
rect 19720 33152 19736 33216
rect 19800 33152 19816 33216
rect 19880 33152 19888 33216
rect 19568 32128 19888 33152
rect 19568 32064 19576 32128
rect 19640 32064 19656 32128
rect 19720 32064 19736 32128
rect 19800 32064 19816 32128
rect 19880 32064 19888 32128
rect 19568 31040 19888 32064
rect 19568 30976 19576 31040
rect 19640 30976 19656 31040
rect 19720 30976 19736 31040
rect 19800 30976 19816 31040
rect 19880 30976 19888 31040
rect 19568 29952 19888 30976
rect 19568 29888 19576 29952
rect 19640 29888 19656 29952
rect 19720 29888 19736 29952
rect 19800 29888 19816 29952
rect 19880 29888 19888 29952
rect 18827 28932 18893 28933
rect 18827 28868 18828 28932
rect 18892 28868 18893 28932
rect 18827 28867 18893 28868
rect 18830 23221 18890 28867
rect 19568 28864 19888 29888
rect 19568 28800 19576 28864
rect 19640 28800 19656 28864
rect 19720 28800 19736 28864
rect 19800 28800 19816 28864
rect 19880 28800 19888 28864
rect 19568 27776 19888 28800
rect 19568 27712 19576 27776
rect 19640 27712 19656 27776
rect 19720 27712 19736 27776
rect 19800 27712 19816 27776
rect 19880 27712 19888 27776
rect 19568 26688 19888 27712
rect 19568 26624 19576 26688
rect 19640 26624 19656 26688
rect 19720 26624 19736 26688
rect 19800 26624 19816 26688
rect 19880 26624 19888 26688
rect 19568 25600 19888 26624
rect 19568 25536 19576 25600
rect 19640 25536 19656 25600
rect 19720 25536 19736 25600
rect 19800 25536 19816 25600
rect 19880 25536 19888 25600
rect 19568 24512 19888 25536
rect 19568 24448 19576 24512
rect 19640 24448 19656 24512
rect 19720 24448 19736 24512
rect 19800 24448 19816 24512
rect 19880 24448 19888 24512
rect 19568 23424 19888 24448
rect 19568 23360 19576 23424
rect 19640 23360 19656 23424
rect 19720 23360 19736 23424
rect 19800 23360 19816 23424
rect 19880 23360 19888 23424
rect 18827 23220 18893 23221
rect 18827 23156 18828 23220
rect 18892 23156 18893 23220
rect 18827 23155 18893 23156
rect 19568 22336 19888 23360
rect 19568 22272 19576 22336
rect 19640 22272 19656 22336
rect 19720 22272 19736 22336
rect 19800 22272 19816 22336
rect 19880 22272 19888 22336
rect 19568 21248 19888 22272
rect 19568 21184 19576 21248
rect 19640 21184 19656 21248
rect 19720 21184 19736 21248
rect 19800 21184 19816 21248
rect 19880 21184 19888 21248
rect 19568 20160 19888 21184
rect 19568 20096 19576 20160
rect 19640 20096 19656 20160
rect 19720 20096 19736 20160
rect 19800 20096 19816 20160
rect 19880 20096 19888 20160
rect 19568 19072 19888 20096
rect 19568 19008 19576 19072
rect 19640 19008 19656 19072
rect 19720 19008 19736 19072
rect 19800 19008 19816 19072
rect 19880 19008 19888 19072
rect 19568 17984 19888 19008
rect 19568 17920 19576 17984
rect 19640 17920 19656 17984
rect 19720 17920 19736 17984
rect 19800 17920 19816 17984
rect 19880 17920 19888 17984
rect 19568 16896 19888 17920
rect 19568 16832 19576 16896
rect 19640 16832 19656 16896
rect 19720 16832 19736 16896
rect 19800 16832 19816 16896
rect 19880 16832 19888 16896
rect 19568 15808 19888 16832
rect 19568 15744 19576 15808
rect 19640 15744 19656 15808
rect 19720 15744 19736 15808
rect 19800 15744 19816 15808
rect 19880 15744 19888 15808
rect 19568 14720 19888 15744
rect 19568 14656 19576 14720
rect 19640 14656 19656 14720
rect 19720 14656 19736 14720
rect 19800 14656 19816 14720
rect 19880 14656 19888 14720
rect 19568 13632 19888 14656
rect 19568 13568 19576 13632
rect 19640 13568 19656 13632
rect 19720 13568 19736 13632
rect 19800 13568 19816 13632
rect 19880 13568 19888 13632
rect 19568 12544 19888 13568
rect 19568 12480 19576 12544
rect 19640 12480 19656 12544
rect 19720 12480 19736 12544
rect 19800 12480 19816 12544
rect 19880 12480 19888 12544
rect 19568 11456 19888 12480
rect 19568 11392 19576 11456
rect 19640 11392 19656 11456
rect 19720 11392 19736 11456
rect 19800 11392 19816 11456
rect 19880 11392 19888 11456
rect 19568 10368 19888 11392
rect 19568 10304 19576 10368
rect 19640 10304 19656 10368
rect 19720 10304 19736 10368
rect 19800 10304 19816 10368
rect 19880 10304 19888 10368
rect 19568 9280 19888 10304
rect 19568 9216 19576 9280
rect 19640 9216 19656 9280
rect 19720 9216 19736 9280
rect 19800 9216 19816 9280
rect 19880 9216 19888 9280
rect 19568 8192 19888 9216
rect 19568 8128 19576 8192
rect 19640 8128 19656 8192
rect 19720 8128 19736 8192
rect 19800 8128 19816 8192
rect 19880 8128 19888 8192
rect 19568 7104 19888 8128
rect 19568 7040 19576 7104
rect 19640 7040 19656 7104
rect 19720 7040 19736 7104
rect 19800 7040 19816 7104
rect 19880 7040 19888 7104
rect 19568 6016 19888 7040
rect 19568 5952 19576 6016
rect 19640 5952 19656 6016
rect 19720 5952 19736 6016
rect 19800 5952 19816 6016
rect 19880 5952 19888 6016
rect 19568 4928 19888 5952
rect 19568 4864 19576 4928
rect 19640 4864 19656 4928
rect 19720 4864 19736 4928
rect 19800 4864 19816 4928
rect 19880 4864 19888 4928
rect 19568 3840 19888 4864
rect 19568 3776 19576 3840
rect 19640 3776 19656 3840
rect 19720 3776 19736 3840
rect 19800 3776 19816 3840
rect 19880 3776 19888 3840
rect 19568 2752 19888 3776
rect 19568 2688 19576 2752
rect 19640 2688 19656 2752
rect 19720 2688 19736 2752
rect 19800 2688 19816 2752
rect 19880 2688 19888 2752
rect 4208 2128 4528 2144
rect 19568 2128 19888 2688
rect 20228 2176 20548 38624
rect 20888 2176 21208 38624
rect 21548 2176 21868 38624
rect 34928 38112 35248 38672
rect 34928 38048 34936 38112
rect 35000 38048 35016 38112
rect 35080 38048 35096 38112
rect 35160 38048 35176 38112
rect 35240 38048 35248 38112
rect 34928 37024 35248 38048
rect 34928 36960 34936 37024
rect 35000 36960 35016 37024
rect 35080 36960 35096 37024
rect 35160 36960 35176 37024
rect 35240 36960 35248 37024
rect 34928 35936 35248 36960
rect 34928 35872 34936 35936
rect 35000 35872 35016 35936
rect 35080 35872 35096 35936
rect 35160 35872 35176 35936
rect 35240 35872 35248 35936
rect 34928 34848 35248 35872
rect 34928 34784 34936 34848
rect 35000 34784 35016 34848
rect 35080 34784 35096 34848
rect 35160 34784 35176 34848
rect 35240 34784 35248 34848
rect 34928 33760 35248 34784
rect 34928 33696 34936 33760
rect 35000 33696 35016 33760
rect 35080 33696 35096 33760
rect 35160 33696 35176 33760
rect 35240 33696 35248 33760
rect 34928 32672 35248 33696
rect 34928 32608 34936 32672
rect 35000 32608 35016 32672
rect 35080 32608 35096 32672
rect 35160 32608 35176 32672
rect 35240 32608 35248 32672
rect 34928 31584 35248 32608
rect 34928 31520 34936 31584
rect 35000 31520 35016 31584
rect 35080 31520 35096 31584
rect 35160 31520 35176 31584
rect 35240 31520 35248 31584
rect 34928 30496 35248 31520
rect 34928 30432 34936 30496
rect 35000 30432 35016 30496
rect 35080 30432 35096 30496
rect 35160 30432 35176 30496
rect 35240 30432 35248 30496
rect 34928 29408 35248 30432
rect 34928 29344 34936 29408
rect 35000 29344 35016 29408
rect 35080 29344 35096 29408
rect 35160 29344 35176 29408
rect 35240 29344 35248 29408
rect 34928 28320 35248 29344
rect 34928 28256 34936 28320
rect 35000 28256 35016 28320
rect 35080 28256 35096 28320
rect 35160 28256 35176 28320
rect 35240 28256 35248 28320
rect 34928 27232 35248 28256
rect 34928 27168 34936 27232
rect 35000 27168 35016 27232
rect 35080 27168 35096 27232
rect 35160 27168 35176 27232
rect 35240 27168 35248 27232
rect 34928 26144 35248 27168
rect 34928 26080 34936 26144
rect 35000 26080 35016 26144
rect 35080 26080 35096 26144
rect 35160 26080 35176 26144
rect 35240 26080 35248 26144
rect 34928 25056 35248 26080
rect 34928 24992 34936 25056
rect 35000 24992 35016 25056
rect 35080 24992 35096 25056
rect 35160 24992 35176 25056
rect 35240 24992 35248 25056
rect 34928 23968 35248 24992
rect 34928 23904 34936 23968
rect 35000 23904 35016 23968
rect 35080 23904 35096 23968
rect 35160 23904 35176 23968
rect 35240 23904 35248 23968
rect 34928 22880 35248 23904
rect 34928 22816 34936 22880
rect 35000 22816 35016 22880
rect 35080 22816 35096 22880
rect 35160 22816 35176 22880
rect 35240 22816 35248 22880
rect 34928 21792 35248 22816
rect 34928 21728 34936 21792
rect 35000 21728 35016 21792
rect 35080 21728 35096 21792
rect 35160 21728 35176 21792
rect 35240 21728 35248 21792
rect 34928 20704 35248 21728
rect 34928 20640 34936 20704
rect 35000 20640 35016 20704
rect 35080 20640 35096 20704
rect 35160 20640 35176 20704
rect 35240 20640 35248 20704
rect 34928 19616 35248 20640
rect 34928 19552 34936 19616
rect 35000 19552 35016 19616
rect 35080 19552 35096 19616
rect 35160 19552 35176 19616
rect 35240 19552 35248 19616
rect 34928 18528 35248 19552
rect 34928 18464 34936 18528
rect 35000 18464 35016 18528
rect 35080 18464 35096 18528
rect 35160 18464 35176 18528
rect 35240 18464 35248 18528
rect 34928 17440 35248 18464
rect 34928 17376 34936 17440
rect 35000 17376 35016 17440
rect 35080 17376 35096 17440
rect 35160 17376 35176 17440
rect 35240 17376 35248 17440
rect 34928 16352 35248 17376
rect 34928 16288 34936 16352
rect 35000 16288 35016 16352
rect 35080 16288 35096 16352
rect 35160 16288 35176 16352
rect 35240 16288 35248 16352
rect 34928 15264 35248 16288
rect 34928 15200 34936 15264
rect 35000 15200 35016 15264
rect 35080 15200 35096 15264
rect 35160 15200 35176 15264
rect 35240 15200 35248 15264
rect 34928 14176 35248 15200
rect 34928 14112 34936 14176
rect 35000 14112 35016 14176
rect 35080 14112 35096 14176
rect 35160 14112 35176 14176
rect 35240 14112 35248 14176
rect 34928 13088 35248 14112
rect 34928 13024 34936 13088
rect 35000 13024 35016 13088
rect 35080 13024 35096 13088
rect 35160 13024 35176 13088
rect 35240 13024 35248 13088
rect 34928 12000 35248 13024
rect 34928 11936 34936 12000
rect 35000 11936 35016 12000
rect 35080 11936 35096 12000
rect 35160 11936 35176 12000
rect 35240 11936 35248 12000
rect 34928 10912 35248 11936
rect 34928 10848 34936 10912
rect 35000 10848 35016 10912
rect 35080 10848 35096 10912
rect 35160 10848 35176 10912
rect 35240 10848 35248 10912
rect 34928 9824 35248 10848
rect 34928 9760 34936 9824
rect 35000 9760 35016 9824
rect 35080 9760 35096 9824
rect 35160 9760 35176 9824
rect 35240 9760 35248 9824
rect 34928 8736 35248 9760
rect 34928 8672 34936 8736
rect 35000 8672 35016 8736
rect 35080 8672 35096 8736
rect 35160 8672 35176 8736
rect 35240 8672 35248 8736
rect 34928 7648 35248 8672
rect 34928 7584 34936 7648
rect 35000 7584 35016 7648
rect 35080 7584 35096 7648
rect 35160 7584 35176 7648
rect 35240 7584 35248 7648
rect 34928 6560 35248 7584
rect 34928 6496 34936 6560
rect 35000 6496 35016 6560
rect 35080 6496 35096 6560
rect 35160 6496 35176 6560
rect 35240 6496 35248 6560
rect 34928 5472 35248 6496
rect 34928 5408 34936 5472
rect 35000 5408 35016 5472
rect 35080 5408 35096 5472
rect 35160 5408 35176 5472
rect 35240 5408 35248 5472
rect 34928 4384 35248 5408
rect 34928 4320 34936 4384
rect 35000 4320 35016 4384
rect 35080 4320 35096 4384
rect 35160 4320 35176 4384
rect 35240 4320 35248 4384
rect 34928 3296 35248 4320
rect 34928 3232 34936 3296
rect 35000 3232 35016 3296
rect 35080 3232 35096 3296
rect 35160 3232 35176 3296
rect 35240 3232 35248 3296
rect 34928 2208 35248 3232
rect 34928 2144 34936 2208
rect 35000 2144 35016 2208
rect 35080 2144 35096 2208
rect 35160 2144 35176 2208
rect 35240 2144 35248 2208
rect 35588 2176 35908 38624
rect 36248 2176 36568 38624
rect 36908 2176 37228 38624
rect 34928 2128 35248 2144
use sky130_fd_sc_hd__fill_1  FILLER_1_7 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 1748 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 1380 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_15 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 2484 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_3
timestamp 1608254825
transform 1 0 1380 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1608254825
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _2500_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 1840 0 1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_1_39 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 4692 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_1_27
timestamp 1608254825
transform 1 0 3588 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27
timestamp 1608254825
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2509_
timestamp 1608254825
transform 1 0 4048 0 -1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_1_57
timestamp 1608254825
transform 1 0 6348 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_47
timestamp 1608254825
transform 1 0 5428 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51
timestamp 1608254825
transform 1 0 5796 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_4  _2343_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 5520 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_1_62
timestamp 1608254825
transform 1 0 6808 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_59
timestamp 1608254825
transform 1 0 6532 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1608254825
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1608254825
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2533_
timestamp 1608254825
transform 1 0 6900 0 -1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _2530_
timestamp 1608254825
transform 1 0 7176 0 1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_1_85
timestamp 1608254825
transform 1 0 8924 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_89
timestamp 1608254825
transform 1 0 9292 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_82
timestamp 1608254825
transform 1 0 8648 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2528_
timestamp 1608254825
transform 1 0 9292 0 1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_2  _2342_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 9016 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_108
timestamp 1608254825
transform 1 0 11040 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_100
timestamp 1608254825
transform 1 0 10304 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_94 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 9752 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1608254825
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2526_
timestamp 1608254825
transform 1 0 10396 0 -1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_1_120 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 12144 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_125
timestamp 1608254825
transform 1 0 12604 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_120
timestamp 1608254825
transform 1 0 12144 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1608254825
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1608254825
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _1931_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 12420 0 1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_1_134
timestamp 1608254825
transform 1 0 13432 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_130
timestamp 1608254825
transform 1 0 13064 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_131
timestamp 1608254825
transform 1 0 13156 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2537_
timestamp 1608254825
transform 1 0 13248 0 -1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _2527_
timestamp 1608254825
transform 1 0 13524 0 1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_1_154
timestamp 1608254825
transform 1 0 15272 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_156
timestamp 1608254825
transform 1 0 15456 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_151
timestamp 1608254825
transform 1 0 14996 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1608254825
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2525_
timestamp 1608254825
transform 1 0 15548 0 -1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__and2_4  _1922_
timestamp 1608254825
transform 1 0 15640 0 1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_1_182
timestamp 1608254825
transform 1 0 17848 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_176
timestamp 1608254825
transform 1 0 17296 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_165
timestamp 1608254825
transform 1 0 16284 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_176
timestamp 1608254825
transform 1 0 17296 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__and2_4  _1932_
timestamp 1608254825
transform 1 0 16652 0 1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_1_194
timestamp 1608254825
transform 1 0 18952 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_184
timestamp 1608254825
transform 1 0 18032 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_190
timestamp 1608254825
transform 1 0 18584 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_184
timestamp 1608254825
transform 1 0 18032 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1608254825
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1608254825
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _1936_
timestamp 1608254825
transform 1 0 18124 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1622_
timestamp 1608254825
transform 1 0 18308 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _2522_
timestamp 1608254825
transform 1 0 18952 0 -1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _2520_
timestamp 1608254825
transform 1 0 19504 0 1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_1_219
timestamp 1608254825
transform 1 0 21252 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_224
timestamp 1608254825
transform 1 0 21712 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_218
timestamp 1608254825
transform 1 0 21160 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_213
timestamp 1608254825
transform 1 0 20700 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1608254825
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2514_
timestamp 1608254825
transform 1 0 21804 0 -1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__and2_4  _1934_
timestamp 1608254825
transform 1 0 21620 0 1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_1_242
timestamp 1608254825
transform 1 0 23368 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_230
timestamp 1608254825
transform 1 0 22264 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_244
timestamp 1608254825
transform 1 0 23552 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1608254825
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1608254825
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2512_
timestamp 1608254825
transform 1 0 24012 0 -1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__and2_4  _1953_
timestamp 1608254825
transform 1 0 23644 0 1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_1_258
timestamp 1608254825
transform 1 0 24840 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_252
timestamp 1608254825
transform 1 0 24288 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_268
timestamp 1608254825
transform 1 0 25760 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _2523_
timestamp 1608254825
transform 1 0 24932 0 1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_1_278
timestamp 1608254825
transform 1 0 26680 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_276
timestamp 1608254825
transform 1 0 26496 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1608254825
transform 1 0 26772 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2578_
timestamp 1608254825
transform 1 0 27048 0 1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _2531_
timestamp 1608254825
transform 1 0 26864 0 -1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_1_306
timestamp 1608254825
transform 1 0 29256 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_301
timestamp 1608254825
transform 1 0 28796 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_306
timestamp 1608254825
transform 1 0 29256 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_299
timestamp 1608254825
transform 1 0 28612 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1608254825
transform 1 0 29164 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1608254825
transform 1 0 29624 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2576_
timestamp 1608254825
transform 1 0 29992 0 1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__conb_1  _2357_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 28980 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_4  _1814_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 29716 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_333
timestamp 1608254825
transform 1 0 31740 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_335
timestamp 1608254825
transform 1 0 31924 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_323
timestamp 1608254825
transform 1 0 30820 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1608254825
transform 1 0 32476 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2575_
timestamp 1608254825
transform 1 0 32108 0 1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__o21a_4  _1818_
timestamp 1608254825
transform 1 0 32568 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_364
timestamp 1608254825
transform 1 0 34592 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_356
timestamp 1608254825
transform 1 0 33856 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_0_354
timestamp 1608254825
transform 1 0 33672 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_379
timestamp 1608254825
transform 1 0 35972 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_385
timestamp 1608254825
transform 1 0 36524 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_373
timestamp 1608254825
transform 1 0 35420 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_366
timestamp 1608254825
transform 1 0 34776 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1608254825
transform 1 0 34776 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1608254825
transform 1 0 35328 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_4  _1820_
timestamp 1608254825
transform 1 0 34868 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_403
timestamp 1608254825
transform 1 0 38180 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_391
timestamp 1608254825
transform 1 0 37076 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_407
timestamp 1608254825
transform 1 0 38548 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_397
timestamp 1608254825
transform 1 0 37628 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1608254825
transform 1 0 38180 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _2358_
timestamp 1608254825
transform 1 0 38272 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_415
timestamp 1608254825
transform 1 0 39284 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_415
timestamp 1608254825
transform 1 0 39284 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1608254825
transform -1 0 39836 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1608254825
transform -1 0 39836 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_15
timestamp 1608254825
transform 1 0 2484 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1608254825
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1608254825
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_32
timestamp 1608254825
transform 1 0 4048 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_27
timestamp 1608254825
transform 1 0 3588 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1608254825
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _1919_
timestamp 1608254825
transform 1 0 5152 0 -1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_2_61
timestamp 1608254825
transform 1 0 6716 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_51
timestamp 1608254825
transform 1 0 5796 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_4  _2344_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 7084 0 -1 3808
box -38 -48 1234 592
use sky130_fd_sc_hd__buf_2  _1950_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 6348 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_86
timestamp 1608254825
transform 1 0 9016 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_78
timestamp 1608254825
transform 1 0 8280 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1912_
timestamp 1608254825
transform 1 0 8648 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_113
timestamp 1608254825
transform 1 0 11500 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_109
timestamp 1608254825
transform 1 0 11132 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_102
timestamp 1608254825
transform 1 0 10488 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1608254825
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2529_
timestamp 1608254825
transform 1 0 11592 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_2  _1927_
timestamp 1608254825
transform 1 0 10856 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_4  _1924_
timestamp 1608254825
transform 1 0 9660 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_2_133
timestamp 1608254825
transform 1 0 13340 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_4  _1914_
timestamp 1608254825
transform 1 0 13708 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_2_154
timestamp 1608254825
transform 1 0 15272 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_152
timestamp 1608254825
transform 1 0 15088 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_146
timestamp 1608254825
transform 1 0 14536 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1608254825
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_180
timestamp 1608254825
transform 1 0 17664 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_160
timestamp 1608254825
transform 1 0 15824 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2426_
timestamp 1608254825
transform 1 0 15916 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_2_203
timestamp 1608254825
transform 1 0 19780 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _2524_
timestamp 1608254825
transform 1 0 18032 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_2_226
timestamp 1608254825
transform 1 0 21896 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_215
timestamp 1608254825
transform 1 0 20884 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_2_211
timestamp 1608254825
transform 1 0 20516 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1608254825
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _1951_
timestamp 1608254825
transform 1 0 21252 0 -1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_2_232
timestamp 1608254825
transform 1 0 22448 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2510_
timestamp 1608254825
transform 1 0 22540 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_2_271
timestamp 1608254825
transform 1 0 26036 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_258
timestamp 1608254825
transform 1 0 24840 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_252
timestamp 1608254825
transform 1 0 24288 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_4  _1812_
timestamp 1608254825
transform 1 0 24932 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_284
timestamp 1608254825
transform 1 0 27232 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_276
timestamp 1608254825
transform 1 0 26496 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1608254825
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_4  _1811_
timestamp 1608254825
transform 1 0 27416 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_298
timestamp 1608254825
transform 1 0 28520 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2577_
timestamp 1608254825
transform 1 0 28888 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  FILLER_2_333
timestamp 1608254825
transform 1 0 31740 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_321
timestamp 1608254825
transform 1 0 30636 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1608254825
transform 1 0 32016 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_4  _1816_
timestamp 1608254825
transform 1 0 32108 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_349
timestamp 1608254825
transform 1 0 33212 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2574_
timestamp 1608254825
transform 1 0 33580 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_2_380
timestamp 1608254825
transform 1 0 36064 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_372
timestamp 1608254825
transform 1 0 35328 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1810_
timestamp 1608254825
transform 1 0 35696 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_410
timestamp 1608254825
transform 1 0 38824 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_2_398
timestamp 1608254825
transform 1 0 37720 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_396
timestamp 1608254825
transform 1 0 37536 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_392
timestamp 1608254825
transform 1 0 37168 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1608254825
transform 1 0 37628 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1608254825
transform -1 0 39836 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_15
timestamp 1608254825
transform 1 0 2484 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1608254825
transform 1 0 1380 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1608254825
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_27
timestamp 1608254825
transform 1 0 3588 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2539_
timestamp 1608254825
transform 1 0 3680 0 1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_3_57
timestamp 1608254825
transform 1 0 6348 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_47
timestamp 1608254825
transform 1 0 5428 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1608254825
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _1940_
timestamp 1608254825
transform 1 0 6808 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _1935_
timestamp 1608254825
transform 1 0 5980 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_79
timestamp 1608254825
transform 1 0 8372 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_71
timestamp 1608254825
transform 1 0 7636 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2412_
timestamp 1608254825
transform 1 0 8740 0 1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  _1921_
timestamp 1608254825
transform 1 0 8004 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_102
timestamp 1608254825
transform 1 0 10488 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_4  _1926_
timestamp 1608254825
transform 1 0 11040 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_3_123
timestamp 1608254825
transform 1 0 12420 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_121
timestamp 1608254825
transform 1 0 12236 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_117
timestamp 1608254825
transform 1 0 11868 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1608254825
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _1930_
timestamp 1608254825
transform 1 0 12972 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_3_144
timestamp 1608254825
transform 1 0 14352 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_138
timestamp 1608254825
transform 1 0 13800 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  _2425_
timestamp 1608254825
transform 1 0 14444 0 1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_3_179
timestamp 1608254825
transform 1 0 17572 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_164
timestamp 1608254825
transform 1 0 16192 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_4  _1942_
timestamp 1608254825
transform 1 0 16744 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_3_199
timestamp 1608254825
transform 1 0 19412 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_3_184
timestamp 1608254825
transform 1 0 18032 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1608254825
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2518_
timestamp 1608254825
transform 1 0 19964 0 1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__nor2_4  _1939_
timestamp 1608254825
transform 1 0 18584 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_3_224
timestamp 1608254825
transform 1 0 21712 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__and2_4  _1952_
timestamp 1608254825
transform 1 0 22080 0 1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_3_245
timestamp 1608254825
transform 1 0 23644 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_243
timestamp 1608254825
transform 1 0 23460 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_235
timestamp 1608254825
transform 1 0 22724 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1608254825
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_272
timestamp 1608254825
transform 1 0 26128 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_3_257
timestamp 1608254825
transform 1 0 24748 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_4  _1815_
timestamp 1608254825
transform 1 0 25024 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_295
timestamp 1608254825
transform 1 0 28244 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _2579_
timestamp 1608254825
transform 1 0 26496 0 1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_3_310
timestamp 1608254825
transform 1 0 29624 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_303
timestamp 1608254825
transform 1 0 28980 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1608254825
transform 1 0 29164 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1813_
timestamp 1608254825
transform 1 0 29256 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_4  _1801_
timestamp 1608254825
transform 1 0 30360 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_330
timestamp 1608254825
transform 1 0 31464 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_4  _1817_
timestamp 1608254825
transform 1 0 31832 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_362
timestamp 1608254825
transform 1 0 34408 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_346
timestamp 1608254825
transform 1 0 32936 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_4  _1819_
timestamp 1608254825
transform 1 0 33304 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_379
timestamp 1608254825
transform 1 0 35972 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1608254825
transform 1 0 34776 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_4  _1822_
timestamp 1608254825
transform 1 0 34868 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_403
timestamp 1608254825
transform 1 0 38180 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_391
timestamp 1608254825
transform 1 0 37076 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_415
timestamp 1608254825
transform 1 0 39284 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1608254825
transform -1 0 39836 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1608254825
transform 1 0 2484 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1608254825
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1608254825
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_40
timestamp 1608254825
transform 1 0 4784 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_4_32
timestamp 1608254825
transform 1 0 4048 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_27
timestamp 1608254825
transform 1 0 3588 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1608254825
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1915_
timestamp 1608254825
transform 1 0 5060 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_47
timestamp 1608254825
transform 1 0 5428 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2519_
timestamp 1608254825
transform 1 0 5796 0 -1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_4_88
timestamp 1608254825
transform 1 0 9200 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_70
timestamp 1608254825
transform 1 0 7544 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_0_0_addressalyzerBlock.SPI_CLK $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 8096 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_4  _1928_
timestamp 1608254825
transform 1 0 8372 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_4_93
timestamp 1608254825
transform 1 0 9660 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1608254825
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2413_
timestamp 1608254825
transform 1 0 10212 0 -1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_4_118
timestamp 1608254825
transform 1 0 11960 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2411_
timestamp 1608254825
transform 1 0 12328 0 -1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  FILLER_4_154
timestamp 1608254825
transform 1 0 15272 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_152
timestamp 1608254825
transform 1 0 15088 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_148
timestamp 1608254825
transform 1 0 14720 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_141
timestamp 1608254825
transform 1 0 14076 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1608254825
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__o32ai_4  _2269_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 15548 0 -1 4896
box -38 -48 2062 592
use sky130_fd_sc_hd__inv_2  _1929_
timestamp 1608254825
transform 1 0 14444 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_179
timestamp 1608254825
transform 1 0 17572 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_202
timestamp 1608254825
transform 1 0 19688 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2424_
timestamp 1608254825
transform 1 0 17940 0 -1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_4_228
timestamp 1608254825
transform 1 0 22080 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_213
timestamp 1608254825
transform 1 0 20700 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_209
timestamp 1608254825
transform 1 0 20332 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1608254825
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_4  _2129_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 20884 0 -1 4896
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _1847_
timestamp 1608254825
transform 1 0 20056 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_236
timestamp 1608254825
transform 1 0 22816 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2586_
timestamp 1608254825
transform 1 0 22908 0 -1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_4_274
timestamp 1608254825
transform 1 0 26312 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_266
timestamp 1608254825
transform 1 0 25576 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_262
timestamp 1608254825
transform 1 0 25208 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_256
timestamp 1608254825
transform 1 0 24656 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _2223_
timestamp 1608254825
transform 1 0 25300 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_4_294
timestamp 1608254825
transform 1 0 28152 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_4_276
timestamp 1608254825
transform 1 0 26496 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1608254825
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_4  _1794_
timestamp 1608254825
transform 1 0 27048 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_317
timestamp 1608254825
transform 1 0 30268 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_302
timestamp 1608254825
transform 1 0 28888 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_4  _1798_
timestamp 1608254825
transform 1 0 29164 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_335
timestamp 1608254825
transform 1 0 31924 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_329
timestamp 1608254825
transform 1 0 31372 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1608254825
transform 1 0 32016 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_4  _1803_
timestamp 1608254825
transform 1 0 32108 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_365
timestamp 1608254825
transform 1 0 34684 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_349
timestamp 1608254825
transform 1 0 33212 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_4  _1821_
timestamp 1608254825
transform 1 0 33580 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_388
timestamp 1608254825
transform 1 0 36800 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _2513_
timestamp 1608254825
transform 1 0 35052 0 -1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_4_410
timestamp 1608254825
transform 1 0 38824 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_4_398
timestamp 1608254825
transform 1 0 37720 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_396
timestamp 1608254825
transform 1 0 37536 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1608254825
transform 1 0 37628 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1608254825
transform -1 0 39836 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_15
timestamp 1608254825
transform 1 0 2484 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1608254825
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1608254825
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_37
timestamp 1608254825
transform 1 0 4508 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_33
timestamp 1608254825
transform 1 0 4140 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_23
timestamp 1608254825
transform 1 0 3220 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2433_
timestamp 1608254825
transform 1 0 4600 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__nor2_4  _1909_
timestamp 1608254825
transform 1 0 3312 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_5_62
timestamp 1608254825
transform 1 0 6808 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_57
timestamp 1608254825
transform 1 0 6348 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1608254825
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2414_
timestamp 1608254825
transform 1 0 6992 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_5_83
timestamp 1608254825
transform 1 0 8740 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__o32ai_4  _2287_
timestamp 1608254825
transform 1 0 9108 0 1 4896
box -38 -48 2062 592
use sky130_fd_sc_hd__decap_4  FILLER_5_109
timestamp 1608254825
transform 1 0 11132 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1925_
timestamp 1608254825
transform 1 0 11500 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_123
timestamp 1608254825
transform 1 0 12420 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_5_116
timestamp 1608254825
transform 1 0 11776 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1608254825
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__o32ai_4  _2288_
timestamp 1608254825
transform 1 0 12604 0 1 4896
box -38 -48 2062 592
use sky130_fd_sc_hd__fill_1  FILLER_5_153
timestamp 1608254825
transform 1 0 15180 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_147
timestamp 1608254825
transform 1 0 14628 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__o32ai_4  _2265_
timestamp 1608254825
transform 1 0 15272 0 1 4896
box -38 -48 2062 592
use sky130_fd_sc_hd__decap_4  FILLER_5_176
timestamp 1608254825
transform 1 0 17296 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_5_0_m1_clk_local
timestamp 1608254825
transform 1 0 17664 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_200
timestamp 1608254825
transform 1 0 19504 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_187
timestamp 1608254825
transform 1 0 18308 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1608254825
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2521_
timestamp 1608254825
transform 1 0 19872 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__nor2_4  _1938_
timestamp 1608254825
transform 1 0 18676 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1937_
timestamp 1608254825
transform 1 0 18032 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_223
timestamp 1608254825
transform 1 0 21620 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__and2_4  _1955_
timestamp 1608254825
transform 1 0 21988 0 1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_5_245
timestamp 1608254825
transform 1 0 23644 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_242
timestamp 1608254825
transform 1 0 23368 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_234
timestamp 1608254825
transform 1 0 22632 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1608254825
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1459_
timestamp 1608254825
transform 1 0 24012 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_257
timestamp 1608254825
transform 1 0 24748 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_253
timestamp 1608254825
transform 1 0 24380 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2583_
timestamp 1608254825
transform 1 0 24840 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  FILLER_5_285
timestamp 1608254825
transform 1 0 27324 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_277
timestamp 1608254825
transform 1 0 26588 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_4  _1793_
timestamp 1608254825
transform 1 0 27600 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_304
timestamp 1608254825
transform 1 0 29072 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_300
timestamp 1608254825
transform 1 0 28704 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1608254825
transform 1 0 29164 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2584_
timestamp 1608254825
transform 1 0 29256 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_5_325
timestamp 1608254825
transform 1 0 31004 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  _2582_
timestamp 1608254825
transform 1 0 31556 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_5_365
timestamp 1608254825
transform 1 0 34684 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_361
timestamp 1608254825
transform 1 0 34316 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_356
timestamp 1608254825
transform 1 0 33856 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_350
timestamp 1608254825
transform 1 0 33304 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _1809_
timestamp 1608254825
transform 1 0 33948 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_388
timestamp 1608254825
transform 1 0 36800 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_381
timestamp 1608254825
transform 1 0 36156 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_367
timestamp 1608254825
transform 1 0 34868 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1608254825
transform 1 0 34776 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_4  _1827_
timestamp 1608254825
transform 1 0 35052 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1808_
timestamp 1608254825
transform 1 0 36524 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_400
timestamp 1608254825
transform 1 0 37904 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_412
timestamp 1608254825
transform 1 0 39008 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1608254825
transform -1 0 39836 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1608254825
transform 1 0 2484 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1608254825
transform 1 0 1380 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1608254825
transform 1 0 2484 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1608254825
transform 1 0 1380 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1608254825
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1608254825
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_27
timestamp 1608254825
transform 1 0 3588 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_27
timestamp 1608254825
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1608254825
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2429_
timestamp 1608254825
transform 1 0 4048 0 -1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__o32ai_4  _2256_
timestamp 1608254825
transform 1 0 3680 0 1 5984
box -38 -48 2062 592
use sky130_fd_sc_hd__decap_4  FILLER_7_57
timestamp 1608254825
transform 1 0 6348 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_50
timestamp 1608254825
transform 1 0 5704 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_51
timestamp 1608254825
transform 1 0 5796 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__and2_4  _1954_
timestamp 1608254825
transform 1 0 6164 0 -1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1709_
timestamp 1608254825
transform 1 0 6072 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_62
timestamp 1608254825
transform 1 0 6808 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_62
timestamp 1608254825
transform 1 0 6808 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1608254825
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__o32ai_4  _2285_
timestamp 1608254825
transform 1 0 7176 0 -1 5984
box -38 -48 2062 592
use sky130_fd_sc_hd__o32ai_4  _2282_
timestamp 1608254825
transform 1 0 7084 0 1 5984
box -38 -48 2062 592
use sky130_fd_sc_hd__decap_6  FILLER_7_87
timestamp 1608254825
transform 1 0 9108 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_88
timestamp 1608254825
transform 1 0 9200 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_105
timestamp 1608254825
transform 1 0 10764 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_97
timestamp 1608254825
transform 1 0 10028 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_96
timestamp 1608254825
transform 1 0 9936 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1608254825
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__o32ai_4  _2286_
timestamp 1608254825
transform 1 0 10304 0 -1 5984
box -38 -48 2062 592
use sky130_fd_sc_hd__buf_2  _2278_
timestamp 1608254825
transform 1 0 9660 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _2276_
timestamp 1608254825
transform 1 0 10396 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__and2_4  _1933_
timestamp 1608254825
transform 1 0 11132 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1923_
timestamp 1608254825
transform 1 0 9660 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_123
timestamp 1608254825
transform 1 0 12420 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_116
timestamp 1608254825
transform 1 0 11776 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_122
timestamp 1608254825
transform 1 0 12328 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1608254825
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__o32ai_4  _2261_
timestamp 1608254825
transform 1 0 12604 0 1 5984
box -38 -48 2062 592
use sky130_fd_sc_hd__a21oi_4  _2220_
timestamp 1608254825
transform 1 0 12696 0 -1 5984
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_7_147
timestamp 1608254825
transform 1 0 14628 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_146
timestamp 1608254825
transform 1 0 14536 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_139
timestamp 1608254825
transform 1 0 13892 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_addressalyzerBlock.SPI_CLK
timestamp 1608254825
transform 1 0 14260 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_4_0_m1_clk_local
timestamp 1608254825
transform 1 0 14904 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1608254825
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__o32ai_4  _2267_
timestamp 1608254825
transform 1 0 15272 0 -1 5984
box -38 -48 2062 592
use sky130_fd_sc_hd__nor2_4  _1710_
timestamp 1608254825
transform 1 0 14996 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_7_179
timestamp 1608254825
transform 1 0 17572 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_160
timestamp 1608254825
transform 1 0 15824 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_176
timestamp 1608254825
transform 1 0 17296 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2409_
timestamp 1608254825
transform 1 0 17664 0 -1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__o21ai_4  _2296_
timestamp 1608254825
transform 1 0 16376 0 1 5984
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_2  FILLER_7_198
timestamp 1608254825
transform 1 0 19320 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_191
timestamp 1608254825
transform 1 0 18676 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_184
timestamp 1608254825
transform 1 0 18032 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_199
timestamp 1608254825
transform 1 0 19412 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_2_0_addressalyzerBlock.SPI_CLK
timestamp 1608254825
transform 1 0 19044 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_m1_clk_local
timestamp 1608254825
transform 1 0 18400 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_188
timestamp 1608254825
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2445_
timestamp 1608254825
transform 1 0 19504 0 1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_7_219
timestamp 1608254825
transform 1 0 21252 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_218
timestamp 1608254825
transform 1 0 21160 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_6_211
timestamp 1608254825
transform 1 0 20516 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_6_0_m1_clk_local
timestamp 1608254825
transform 1 0 21528 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1608254825
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2446_
timestamp 1608254825
transform 1 0 21804 0 -1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_2  _2239_
timestamp 1608254825
transform 1 0 20884 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_4  _2125_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 21804 0 1 5984
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_1  FILLER_7_243
timestamp 1608254825
transform 1 0 23460 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_239
timestamp 1608254825
transform 1 0 23092 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_251
timestamp 1608254825
transform 1 0 24196 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_244
timestamp 1608254825
transform 1 0 23552 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_189
timestamp 1608254825
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _2266_
timestamp 1608254825
transform 1 0 23920 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_4  _2127_
timestamp 1608254825
transform 1 0 23644 0 1 5984
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_7_273
timestamp 1608254825
transform 1 0 26220 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_267
timestamp 1608254825
transform 1 0 25668 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_259
timestamp 1608254825
transform 1 0 24932 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_271
timestamp 1608254825
transform 1 0 26036 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_4  _2255_
timestamp 1608254825
transform 1 0 24748 0 -1 5984
box -38 -48 1326 592
use sky130_fd_sc_hd__buf_2  _1497_
timestamp 1608254825
transform 1 0 25852 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_296
timestamp 1608254825
transform 1 0 28336 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_294
timestamp 1608254825
transform 1 0 28152 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_276
timestamp 1608254825
transform 1 0 26496 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1608254825
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2587_
timestamp 1608254825
transform 1 0 26588 0 1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__o21a_4  _1792_
timestamp 1608254825
transform 1 0 27048 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_304
timestamp 1608254825
transform 1 0 29072 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_306
timestamp 1608254825
transform 1 0 29256 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_302
timestamp 1608254825
transform 1 0 28888 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_190
timestamp 1608254825
transform 1 0 29164 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1838_
timestamp 1608254825
transform 1 0 29256 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1790_
timestamp 1608254825
transform 1 0 28520 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_318
timestamp 1608254825
transform 1 0 30360 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_310
timestamp 1608254825
transform 1 0 29624 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_6_319
timestamp 1608254825
transform 1 0 30452 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_4  _1800_
timestamp 1608254825
transform 1 0 30452 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__o21a_4  _1797_
timestamp 1608254825
transform 1 0 29348 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_337
timestamp 1608254825
transform 1 0 32108 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_331
timestamp 1608254825
transform 1 0 31556 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_332
timestamp 1608254825
transform 1 0 31648 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_327
timestamp 1608254825
transform 1 0 31188 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1608254825
transform 1 0 32016 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_4  _1807_
timestamp 1608254825
transform 1 0 32200 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__o21a_4  _1802_
timestamp 1608254825
transform 1 0 32108 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _1787_
timestamp 1608254825
transform 1 0 31280 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_365
timestamp 1608254825
transform 1 0 34684 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_357
timestamp 1608254825
transform 1 0 33948 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_7_350
timestamp 1608254825
transform 1 0 33304 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_353
timestamp 1608254825
transform 1 0 33580 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_349
timestamp 1608254825
transform 1 0 33212 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_4  _1823_
timestamp 1608254825
transform 1 0 33672 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1786_
timestamp 1608254825
transform 1 0 33672 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_386
timestamp 1608254825
transform 1 0 36616 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_382
timestamp 1608254825
transform 1 0 36248 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_366
timestamp 1608254825
transform 1 0 34776 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_191
timestamp 1608254825
transform 1 0 34776 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2572_
timestamp 1608254825
transform 1 0 34868 0 1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__o21a_4  _1825_
timestamp 1608254825
transform 1 0 35144 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_402
timestamp 1608254825
transform 1 0 38088 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_410
timestamp 1608254825
transform 1 0 38824 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_6_398
timestamp 1608254825
transform 1 0 37720 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_394
timestamp 1608254825
transform 1 0 37352 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1608254825
transform 1 0 37628 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_4  _1828_
timestamp 1608254825
transform 1 0 36984 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_414
timestamp 1608254825
transform 1 0 39192 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1608254825
transform -1 0 39836 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1608254825
transform -1 0 39836 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_19
timestamp 1608254825
transform 1 0 2852 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_11
timestamp 1608254825
transform 1 0 2116 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_3
timestamp 1608254825
transform 1 0 1380 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1608254825
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__and2_4  _1917_
timestamp 1608254825
transform 1 0 2208 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_8_37
timestamp 1608254825
transform 1 0 4508 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_32
timestamp 1608254825
transform 1 0 4048 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_192
timestamp 1608254825
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__o32ai_4  _2250_
timestamp 1608254825
transform 1 0 4876 0 -1 7072
box -38 -48 2062 592
use sky130_fd_sc_hd__inv_2  _1908_
timestamp 1608254825
transform 1 0 4232 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_63
timestamp 1608254825
transform 1 0 6900 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2417_
timestamp 1608254825
transform 1 0 7268 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_8_86
timestamp 1608254825
transform 1 0 9016 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_112
timestamp 1608254825
transform 1 0 11408 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_93
timestamp 1608254825
transform 1 0 9660 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_193
timestamp 1608254825
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_4  _1849_
timestamp 1608254825
transform 1 0 10212 0 -1 7072
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_8_135
timestamp 1608254825
transform 1 0 13524 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2427_
timestamp 1608254825
transform 1 0 11776 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_8_158
timestamp 1608254825
transform 1 0 15640 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_154
timestamp 1608254825
transform 1 0 15272 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_149
timestamp 1608254825
transform 1 0 14812 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_142
timestamp 1608254825
transform 1 0 14168 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_194
timestamp 1608254825
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_4  _2294_
timestamp 1608254825
transform 1 0 15732 0 -1 7072
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _2277_
timestamp 1608254825
transform 1 0 14536 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1913_
timestamp 1608254825
transform 1 0 13892 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_172
timestamp 1608254825
transform 1 0 16928 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_4  _2295_
timestamp 1608254825
transform 1 0 17296 0 -1 7072
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_6  FILLER_8_190
timestamp 1608254825
transform 1 0 18584 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_4  _2241_
timestamp 1608254825
transform 1 0 19136 0 -1 7072
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_8_210
timestamp 1608254825
transform 1 0 20424 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_195
timestamp 1608254825
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__nand3_4  _2128_
timestamp 1608254825
transform 1 0 20884 0 -1 7072
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_8_250
timestamp 1608254825
transform 1 0 24104 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_229
timestamp 1608254825
transform 1 0 22172 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_7_0_m1_clk_local
timestamp 1608254825
transform 1 0 22540 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_4  _2260_
timestamp 1608254825
transform 1 0 22816 0 -1 7072
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_1  FILLER_8_274
timestamp 1608254825
transform 1 0 26312 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_268
timestamp 1608254825
transform 1 0 25760 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_4  _2253_
timestamp 1608254825
transform 1 0 24472 0 -1 7072
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_1  FILLER_8_286
timestamp 1608254825
transform 1 0 27416 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_280
timestamp 1608254825
transform 1 0 26864 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_196
timestamp 1608254825
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1824_
timestamp 1608254825
transform 1 0 26496 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_4  _1791_
timestamp 1608254825
transform 1 0 27508 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_319
timestamp 1608254825
transform 1 0 30452 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_315
timestamp 1608254825
transform 1 0 30084 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_299
timestamp 1608254825
transform 1 0 28612 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_4  _1795_
timestamp 1608254825
transform 1 0 28980 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_341
timestamp 1608254825
transform 1 0 32476 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_8_332
timestamp 1608254825
transform 1 0 31648 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_197
timestamp 1608254825
transform 1 0 32016 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_4  _1805_
timestamp 1608254825
transform 1 0 30544 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _1788_
timestamp 1608254825
transform 1 0 32108 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_349
timestamp 1608254825
transform 1 0 33212 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _2573_
timestamp 1608254825
transform 1 0 33396 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_8_370
timestamp 1608254825
transform 1 0 35144 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2461_
timestamp 1608254825
transform 1 0 35512 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_8_410
timestamp 1608254825
transform 1 0 38824 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_8_398
timestamp 1608254825
transform 1 0 37720 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_393
timestamp 1608254825
transform 1 0 37260 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_198
timestamp 1608254825
transform 1 0 37628 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1608254825
transform -1 0 39836 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_19
timestamp 1608254825
transform 1 0 2852 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_9
timestamp 1608254825
transform 1 0 1932 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_3
timestamp 1608254825
transform 1 0 1380 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1608254825
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_4  _1905_
timestamp 1608254825
transform 1 0 2024 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_9_42
timestamp 1608254825
transform 1 0 4968 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2432_
timestamp 1608254825
transform 1 0 3220 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_9_66
timestamp 1608254825
transform 1 0 7176 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_9_58
timestamp 1608254825
transform 1 0 6440 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_50
timestamp 1608254825
transform 1 0 5704 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_199
timestamp 1608254825
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _2249_
timestamp 1608254825
transform 1 0 5336 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _2244_
timestamp 1608254825
transform 1 0 6808 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_83
timestamp 1608254825
transform 1 0 8740 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_75
timestamp 1608254825
transform 1 0 8004 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__o32ai_4  _2281_
timestamp 1608254825
transform 1 0 9108 0 1 7072
box -38 -48 2062 592
use sky130_fd_sc_hd__buf_2  _2280_
timestamp 1608254825
transform 1 0 8372 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1705_
timestamp 1608254825
transform 1 0 7728 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_109
timestamp 1608254825
transform 1 0 11132 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1619_
timestamp 1608254825
transform 1 0 11500 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_130
timestamp 1608254825
transform 1 0 13064 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_9_123
timestamp 1608254825
transform 1 0 12420 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_116
timestamp 1608254825
transform 1 0 11776 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_addressalyzerBlock.SPI_CLK
timestamp 1608254825
transform 1 0 12788 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_200
timestamp 1608254825
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_152
timestamp 1608254825
transform 1 0 15088 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_138
timestamp 1608254825
transform 1 0 13800 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_addressalyzerBlock.SPI_CLK
timestamp 1608254825
transform 1 0 15456 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _2410_
timestamp 1608254825
transform 1 0 15732 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__a21oi_4  _1626_
timestamp 1608254825
transform 1 0 13892 0 1 7072
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_1  FILLER_9_182
timestamp 1608254825
transform 1 0 17848 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_178
timestamp 1608254825
transform 1 0 17480 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_190
timestamp 1608254825
transform 1 0 18584 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_184
timestamp 1608254825
transform 1 0 18032 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_201
timestamp 1608254825
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2434_
timestamp 1608254825
transform 1 0 18952 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  _2240_
timestamp 1608254825
transform 1 0 18216 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_220
timestamp 1608254825
transform 1 0 21344 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_213
timestamp 1608254825
transform 1 0 20700 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_m1_clk_local
timestamp 1608254825
transform 1 0 21068 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_4  _2126_
timestamp 1608254825
transform 1 0 21528 0 1 7072
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_1  FILLER_9_243
timestamp 1608254825
transform 1 0 23460 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_235
timestamp 1608254825
transform 1 0 22724 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_202
timestamp 1608254825
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__nand3_4  _2122_
timestamp 1608254825
transform 1 0 23644 0 1 7072
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_9_259
timestamp 1608254825
transform 1 0 24932 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_4  _2257_
timestamp 1608254825
transform 1 0 25300 0 1 7072
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_9_291
timestamp 1608254825
transform 1 0 27876 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_285
timestamp 1608254825
transform 1 0 27324 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_277
timestamp 1608254825
transform 1 0 26588 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _2124_
timestamp 1608254825
transform 1 0 28244 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1799_
timestamp 1608254825
transform 1 0 27508 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_318
timestamp 1608254825
transform 1 0 30360 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_9_299
timestamp 1608254825
transform 1 0 28612 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_203
timestamp 1608254825
transform 1 0 29164 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_4  _1796_
timestamp 1608254825
transform 1 0 29256 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_337
timestamp 1608254825
transform 1 0 32108 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_324
timestamp 1608254825
transform 1 0 30912 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_4  _1806_
timestamp 1608254825
transform 1 0 32476 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__o21a_4  _1804_
timestamp 1608254825
transform 1 0 31004 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_365
timestamp 1608254825
transform 1 0 34684 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_353
timestamp 1608254825
transform 1 0 33580 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_388
timestamp 1608254825
transform 1 0 36800 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_9_367
timestamp 1608254825
transform 1 0 34868 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_204
timestamp 1608254825
transform 1 0 34776 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2502_
timestamp 1608254825
transform 1 0 35052 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _2591_
timestamp 1608254825
transform 1 0 37352 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_9_417
timestamp 1608254825
transform 1 0 39468 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_413
timestamp 1608254825
transform 1 0 39100 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1608254825
transform -1 0 39836 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_10_22
timestamp 1608254825
transform 1 0 3128 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1608254825
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _2535_
timestamp 1608254825
transform 1 0 1380 0 -1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_10_30
timestamp 1608254825
transform 1 0 3864 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_205
timestamp 1608254825
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__o32ai_4  _2251_
timestamp 1608254825
transform 1 0 4048 0 -1 8160
box -38 -48 2062 592
use sky130_fd_sc_hd__decap_4  FILLER_10_54
timestamp 1608254825
transform 1 0 6072 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2416_
timestamp 1608254825
transform 1 0 6440 0 -1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_10_84
timestamp 1608254825
transform 1 0 8832 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_10_77
timestamp 1608254825
transform 1 0 8188 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1844_
timestamp 1608254825
transform 1 0 8556 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_112
timestamp 1608254825
transform 1 0 11408 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_206
timestamp 1608254825
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2418_
timestamp 1608254825
transform 1 0 9660 0 -1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_10_129
timestamp 1608254825
transform 1 0 12972 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_4  _1848_
timestamp 1608254825
transform 1 0 11776 0 -1 8160
box -38 -48 1234 592
use sky130_fd_sc_hd__o21ai_4  _1627_
timestamp 1608254825
transform 1 0 13340 0 -1 8160
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_1  FILLER_10_152
timestamp 1608254825
transform 1 0 15088 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_146
timestamp 1608254825
transform 1 0 14536 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_207
timestamp 1608254825
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _1706_
timestamp 1608254825
transform 1 0 15272 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_10_163
timestamp 1608254825
transform 1 0 16100 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_3_0_addressalyzerBlock.SPI_CLK
timestamp 1608254825
transform 1 0 16652 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_4  _2293_
timestamp 1608254825
transform 1 0 16928 0 -1 8160
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_2  FILLER_10_193
timestamp 1608254825
transform 1 0 18860 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_186
timestamp 1608254825
transform 1 0 18216 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_m1_clk_local
timestamp 1608254825
transform 1 0 18584 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_4  _2242_
timestamp 1608254825
transform 1 0 19044 0 -1 8160
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_2  FILLER_10_215
timestamp 1608254825
transform 1 0 20884 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_208
timestamp 1608254825
transform 1 0 20240 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_208
timestamp 1608254825
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2444_
timestamp 1608254825
transform 1 0 21068 0 -1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_10_240
timestamp 1608254825
transform 1 0 23184 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_236
timestamp 1608254825
transform 1 0 22816 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_4  _2130_
timestamp 1608254825
transform 1 0 23276 0 -1 8160
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_10_271
timestamp 1608254825
transform 1 0 26036 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_263
timestamp 1608254825
transform 1 0 25300 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_255
timestamp 1608254825
transform 1 0 24564 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1789_
timestamp 1608254825
transform 1 0 25668 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1554_
timestamp 1608254825
transform 1 0 24932 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_292
timestamp 1608254825
transform 1 0 27968 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_209
timestamp 1608254825
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _2315_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 26496 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  _1713_
timestamp 1608254825
transform 1 0 28336 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_309
timestamp 1608254825
transform 1 0 29532 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_305
timestamp 1608254825
transform 1 0 29164 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_299
timestamp 1608254825
transform 1 0 28612 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  _2581_
timestamp 1608254825
transform 1 0 29900 0 -1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_2  _1765_
timestamp 1608254825
transform 1 0 29256 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_332
timestamp 1608254825
transform 1 0 31648 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_210
timestamp 1608254825
transform 1 0 32016 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2580_
timestamp 1608254825
transform 1 0 32108 0 -1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_10_356
timestamp 1608254825
transform 1 0 33856 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_4  _1826_
timestamp 1608254825
transform 1 0 34224 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_379
timestamp 1608254825
transform 1 0 35972 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_372
timestamp 1608254825
transform 1 0 35328 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1512_
timestamp 1608254825
transform 1 0 35696 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_10_410
timestamp 1608254825
transform 1 0 38824 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_10_398
timestamp 1608254825
transform 1 0 37720 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_391
timestamp 1608254825
transform 1 0 37076 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_211
timestamp 1608254825
transform 1 0 37628 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1608254825
transform -1 0 39836 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_22
timestamp 1608254825
transform 1 0 3128 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1608254825
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _2541_
timestamp 1608254825
transform 1 0 1380 0 1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_11_34
timestamp 1608254825
transform 1 0 4232 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_30
timestamp 1608254825
transform 1 0 3864 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2431_
timestamp 1608254825
transform 1 0 4600 0 1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_2  _1902_
timestamp 1608254825
transform 1 0 3956 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_62
timestamp 1608254825
transform 1 0 6808 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_57
timestamp 1608254825
transform 1 0 6348 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_212
timestamp 1608254825
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__o32ai_4  _2283_
timestamp 1608254825
transform 1 0 7084 0 1 8160
box -38 -48 2062 592
use sky130_fd_sc_hd__decap_8  FILLER_11_87
timestamp 1608254825
transform 1 0 9108 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_113
timestamp 1608254825
transform 1 0 11500 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_106
timestamp 1608254825
transform 1 0 10856 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_95
timestamp 1608254825
transform 1 0 9844 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_1_0_addressalyzerBlock.SPI_CLK
timestamp 1608254825
transform 1 0 11224 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_4  _1620_
timestamp 1608254825
transform 1 0 10028 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_11_123
timestamp 1608254825
transform 1 0 12420 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_11_118
timestamp 1608254825
transform 1 0 11960 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_213
timestamp 1608254825
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__a211o_4  _1621_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 12972 0 1 8160
box -38 -48 1326 592
use sky130_fd_sc_hd__inv_2  _1617_
timestamp 1608254825
transform 1 0 11684 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_155
timestamp 1608254825
transform 1 0 15364 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_143
timestamp 1608254825
transform 1 0 14260 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__a211o_4  _1707_
timestamp 1608254825
transform 1 0 15456 0 1 8160
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_11_179
timestamp 1608254825
transform 1 0 17572 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_170
timestamp 1608254825
transform 1 0 16744 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _2268_
timestamp 1608254825
transform 1 0 17296 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_199
timestamp 1608254825
transform 1 0 19412 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_193
timestamp 1608254825
transform 1 0 18860 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_214
timestamp 1608254825
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _1714_
timestamp 1608254825
transform 1 0 19504 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  _1712_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 18032 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_11_222
timestamp 1608254825
transform 1 0 21528 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_209
timestamp 1608254825
transform 1 0 20332 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_4  _2131_
timestamp 1608254825
transform 1 0 21896 0 1 8160
box -38 -48 1326 592
use sky130_fd_sc_hd__nor2_4  _1851_
timestamp 1608254825
transform 1 0 20700 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_11_245
timestamp 1608254825
transform 1 0 23644 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_240
timestamp 1608254825
transform 1 0 23184 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_215
timestamp 1608254825
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1873_
timestamp 1608254825
transform 1 0 23920 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_252
timestamp 1608254825
transform 1 0 24288 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2402_
timestamp 1608254825
transform 1 0 24656 0 1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_11_275
timestamp 1608254825
transform 1 0 26404 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2401_
timestamp 1608254825
transform 1 0 26772 0 1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_11_304
timestamp 1608254825
transform 1 0 29072 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_298
timestamp 1608254825
transform 1 0 28520 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_216
timestamp 1608254825
transform 1 0 29164 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2585_
timestamp 1608254825
transform 1 0 29256 0 1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_11_342
timestamp 1608254825
transform 1 0 32568 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_325
timestamp 1608254825
transform 1 0 31004 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_4  _1498_
timestamp 1608254825
transform 1 0 31372 0 1 8160
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_8  FILLER_11_358
timestamp 1608254825
transform 1 0 34040 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_4  _1516_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 32936 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_377
timestamp 1608254825
transform 1 0 35788 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_371
timestamp 1608254825
transform 1 0 35236 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_217
timestamp 1608254825
transform 1 0 34776 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__xor2_4  _1768_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 35880 0 1 8160
box -38 -48 2062 592
use sky130_fd_sc_hd__buf_2  _1520_
timestamp 1608254825
transform 1 0 34868 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_408
timestamp 1608254825
transform 1 0 38640 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_404
timestamp 1608254825
transform 1 0 38272 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_400
timestamp 1608254825
transform 1 0 37904 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1770_
timestamp 1608254825
transform 1 0 38364 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_416
timestamp 1608254825
transform 1 0 39376 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1608254825
transform -1 0 39836 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_12_22
timestamp 1608254825
transform 1 0 3128 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1608254825
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _2542_
timestamp 1608254825
transform 1 0 1380 0 -1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_12_32
timestamp 1608254825
transform 1 0 4048 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_1_0_m1_clk_local
timestamp 1608254825
transform 1 0 3680 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_218
timestamp 1608254825
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__o32ai_4  _2252_
timestamp 1608254825
transform 1 0 4416 0 -1 9248
box -38 -48 2062 592
use sky130_fd_sc_hd__decap_8  FILLER_12_58
timestamp 1608254825
transform 1 0 6440 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__o32ai_4  _2284_
timestamp 1608254825
transform 1 0 7176 0 -1 9248
box -38 -48 2062 592
use sky130_fd_sc_hd__decap_4  FILLER_12_88
timestamp 1608254825
transform 1 0 9200 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_111
timestamp 1608254825
transform 1 0 11316 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_93
timestamp 1608254825
transform 1 0 9660 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_219
timestamp 1608254825
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__a21o_4  _1850_
timestamp 1608254825
transform 1 0 10212 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_129
timestamp 1608254825
transform 1 0 12972 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_4  _2218_
timestamp 1608254825
transform 1 0 13340 0 -1 9248
box -38 -48 1234 592
use sky130_fd_sc_hd__a211o_4  _1846_
timestamp 1608254825
transform 1 0 11684 0 -1 9248
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_1  FILLER_12_152
timestamp 1608254825
transform 1 0 15088 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_146
timestamp 1608254825
transform 1 0 14536 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_220
timestamp 1608254825
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__a211o_4  _1711_
timestamp 1608254825
transform 1 0 15272 0 -1 9248
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_12_168
timestamp 1608254825
transform 1 0 16560 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2408_
timestamp 1608254825
transform 1 0 16928 0 -1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1608254825
transform 1 0 19044 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_191
timestamp 1608254825
transform 1 0 18676 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_4  _1715_
timestamp 1608254825
transform 1 0 19136 0 -1 9248
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_12_215
timestamp 1608254825
transform 1 0 20884 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_210
timestamp 1608254825
transform 1 0 20424 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_221
timestamp 1608254825
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_4  _2132_
timestamp 1608254825
transform 1 0 21252 0 -1 9248
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_12_251
timestamp 1608254825
transform 1 0 24196 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_236
timestamp 1608254825
transform 1 0 22816 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_232
timestamp 1608254825
transform 1 0 22448 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_4  _2133_
timestamp 1608254825
transform 1 0 22908 0 -1 9248
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_12_271
timestamp 1608254825
transform 1 0 26036 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_4  _2314_
timestamp 1608254825
transform 1 0 24564 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_12_288
timestamp 1608254825
transform 1 0 27600 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_279
timestamp 1608254825
transform 1 0 26772 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_222
timestamp 1608254825
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2400_
timestamp 1608254825
transform 1 0 27968 0 -1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_2  _2142_
timestamp 1608254825
transform 1 0 27324 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1636_
timestamp 1608254825
transform 1 0 26496 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_318
timestamp 1608254825
transform 1 0 30360 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_311
timestamp 1608254825
transform 1 0 29716 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1750_
timestamp 1608254825
transform 1 0 30084 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_341
timestamp 1608254825
transform 1 0 32476 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_334
timestamp 1608254825
transform 1 0 31832 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_326
timestamp 1608254825
transform 1 0 31096 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_223
timestamp 1608254825
transform 1 0 32016 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1514_
timestamp 1608254825
transform 1 0 32108 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1477_
timestamp 1608254825
transform 1 0 30728 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_364
timestamp 1608254825
transform 1 0 34592 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2606_
timestamp 1608254825
transform 1 0 32844 0 -1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_12_387
timestamp 1608254825
transform 1 0 36708 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _2608_
timestamp 1608254825
transform 1 0 34960 0 -1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_12_411
timestamp 1608254825
transform 1 0 38916 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_12_395
timestamp 1608254825
transform 1 0 37444 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_224
timestamp 1608254825
transform 1 0 37628 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_4  _1480_
timestamp 1608254825
transform 1 0 37720 0 -1 9248
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_1  FILLER_12_417
timestamp 1608254825
transform 1 0 39468 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1608254825
transform -1 0 39836 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_22
timestamp 1608254825
transform 1 0 3128 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_21
timestamp 1608254825
transform 1 0 3036 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_11
timestamp 1608254825
transform 1 0 2116 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_3
timestamp 1608254825
transform 1 0 1380 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1608254825
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1608254825
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _2536_
timestamp 1608254825
transform 1 0 1380 0 -1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__nor2_4  _1903_
timestamp 1608254825
transform 1 0 2208 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_14_30
timestamp 1608254825
transform 1 0 3864 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_231
timestamp 1608254825
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2430_
timestamp 1608254825
transform 1 0 4048 0 -1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__o32ai_4  _2254_
timestamp 1608254825
transform 1 0 3404 0 1 9248
box -38 -48 2062 592
use sky130_fd_sc_hd__decap_4  FILLER_14_51
timestamp 1608254825
transform 1 0 5796 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_54
timestamp 1608254825
transform 1 0 6072 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_47
timestamp 1608254825
transform 1 0 5428 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _2247_
timestamp 1608254825
transform 1 0 6164 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1904_
timestamp 1608254825
transform 1 0 5796 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_14_67
timestamp 1608254825
transform 1 0 7268 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_59
timestamp 1608254825
transform 1 0 6532 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_62
timestamp 1608254825
transform 1 0 6808 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_60
timestamp 1608254825
transform 1 0 6624 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_225
timestamp 1608254825
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2415_
timestamp 1608254825
transform 1 0 6992 0 1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_14_88
timestamp 1608254825
transform 1 0 9200 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1608254825
transform 1 0 8740 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_79
timestamp 1608254825
transform 1 0 8372 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_90
timestamp 1608254825
transform 1 0 9384 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_83
timestamp 1608254825
transform 1 0 8740 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_4  _2199_
timestamp 1608254825
transform 1 0 7544 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1743_
timestamp 1608254825
transform 1 0 9108 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1624_
timestamp 1608254825
transform 1 0 8832 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_109
timestamp 1608254825
transform 1 0 11132 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_93
timestamp 1608254825
transform 1 0 9660 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_109
timestamp 1608254825
transform 1 0 11132 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_232
timestamp 1608254825
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_4  _1748_
timestamp 1608254825
transform 1 0 9936 0 -1 10336
box -38 -48 1234 592
use sky130_fd_sc_hd__a21oi_4  _1747_
timestamp 1608254825
transform 1 0 9936 0 1 9248
box -38 -48 1234 592
use sky130_fd_sc_hd__buf_2  _1625_
timestamp 1608254825
transform 1 0 11500 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_117
timestamp 1608254825
transform 1 0 11868 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_123
timestamp 1608254825
transform 1 0 12420 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_121
timestamp 1608254825
transform 1 0 12236 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_117
timestamp 1608254825
transform 1 0 11868 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_226
timestamp 1608254825
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _1744_
timestamp 1608254825
transform 1 0 12052 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _1704_
timestamp 1608254825
transform 1 0 12604 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_128
timestamp 1608254825
transform 1 0 12880 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_129
timestamp 1608254825
transform 1 0 12972 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_4  _1853_
timestamp 1608254825
transform 1 0 13248 0 -1 10336
box -38 -48 1234 592
use sky130_fd_sc_hd__a21oi_4  _1639_
timestamp 1608254825
transform 1 0 13340 0 1 9248
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_8  FILLER_14_145
timestamp 1608254825
transform 1 0 14444 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_146
timestamp 1608254825
transform 1 0 14536 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_233
timestamp 1608254825
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__a211o_4  _1745_
timestamp 1608254825
transform 1 0 15272 0 -1 10336
box -38 -48 1326 592
use sky130_fd_sc_hd__a21o_4  _1629_
timestamp 1608254825
transform 1 0 14904 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_172
timestamp 1608254825
transform 1 0 16928 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_168
timestamp 1608254825
transform 1 0 16560 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_179
timestamp 1608254825
transform 1 0 17572 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_162
timestamp 1608254825
transform 1 0 16008 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_4  _2299_
timestamp 1608254825
transform 1 0 16376 0 1 9248
box -38 -48 1234 592
use sky130_fd_sc_hd__nand3_4  _2298_
timestamp 1608254825
transform 1 0 17020 0 -1 10336
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_14_200
timestamp 1608254825
transform 1 0 19504 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_187
timestamp 1608254825
transform 1 0 18308 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_199
timestamp 1608254825
transform 1 0 19412 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_184
timestamp 1608254825
transform 1 0 18032 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_227
timestamp 1608254825
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_4  _1717_
timestamp 1608254825
transform 1 0 18216 0 1 9248
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_4  _1716_
timestamp 1608254825
transform 1 0 18676 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _1633_
timestamp 1608254825
transform 1 0 19872 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1631_
timestamp 1608254825
transform 1 0 19780 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_208
timestamp 1608254825
transform 1 0 20240 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_226
timestamp 1608254825
transform 1 0 21896 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_211
timestamp 1608254825
transform 1 0 20516 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_207
timestamp 1608254825
transform 1 0 20148 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_234
timestamp 1608254825
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__a211o_4  _1852_
timestamp 1608254825
transform 1 0 20884 0 -1 10336
box -38 -48 1326 592
use sky130_fd_sc_hd__a211o_4  _1638_
timestamp 1608254825
transform 1 0 20608 0 1 9248
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_6  FILLER_14_229
timestamp 1608254825
transform 1 0 22172 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_245
timestamp 1608254825
transform 1 0 23644 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_243
timestamp 1608254825
transform 1 0 23460 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_239
timestamp 1608254825
transform 1 0 23092 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_228
timestamp 1608254825
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2443_
timestamp 1608254825
transform 1 0 22724 0 -1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__a2bb2o_4  _2321_
timestamp 1608254825
transform 1 0 24012 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__nor2_4  _1637_
timestamp 1608254825
transform 1 0 22264 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_14_271
timestamp 1608254825
transform 1 0 26036 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_254
timestamp 1608254825
transform 1 0 24472 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_273
timestamp 1608254825
transform 1 0 26220 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_265
timestamp 1608254825
transform 1 0 25484 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _2313_
timestamp 1608254825
transform 1 0 25852 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_4  _2135_
timestamp 1608254825
transform 1 0 24840 0 -1 10336
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_6  FILLER_14_280
timestamp 1608254825
transform 1 0 26864 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1608254825
transform 1 0 26772 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_235
timestamp 1608254825
transform 1 0 26404 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _2311_
timestamp 1608254825
transform 1 0 26496 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_290
timestamp 1608254825
transform 1 0 27784 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_286
timestamp 1608254825
transform 1 0 27416 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_296
timestamp 1608254825
transform 1 0 28336 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1773_
timestamp 1608254825
transform 1 0 27508 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _2399_
timestamp 1608254825
transform 1 0 28152 0 -1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__a2bb2o_4  _2316_
timestamp 1608254825
transform 1 0 26864 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_14_313
timestamp 1608254825
transform 1 0 29900 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_8_0_addressalyzerBlock.SPI_CLK
timestamp 1608254825
transform 1 0 28888 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_229
timestamp 1608254825
transform 1 0 29164 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2398_
timestamp 1608254825
transform 1 0 29256 0 1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__a21oi_4  _1521_
timestamp 1608254825
transform 1 0 30452 0 -1 10336
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_14_332
timestamp 1608254825
transform 1 0 31648 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_342
timestamp 1608254825
transform 1 0 32568 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_325
timestamp 1608254825
transform 1 0 31004 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_236
timestamp 1608254825
transform 1 0 32016 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_4  _1515_
timestamp 1608254825
transform 1 0 32108 0 -1 10336
box -38 -48 1234 592
use sky130_fd_sc_hd__a21oi_4  _1478_
timestamp 1608254825
transform 1 0 31372 0 1 9248
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_8  FILLER_14_358
timestamp 1608254825
transform 1 0 34040 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_14_350
timestamp 1608254825
transform 1 0 33304 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_362
timestamp 1608254825
transform 1 0 34408 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_348
timestamp 1608254825
transform 1 0 33120 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_4  _1502_
timestamp 1608254825
transform 1 0 33212 0 1 9248
box -38 -48 1234 592
use sky130_fd_sc_hd__buf_2  _1462_
timestamp 1608254825
transform 1 0 33672 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_388
timestamp 1608254825
transform 1 0 36800 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_384
timestamp 1608254825
transform 1 0 36432 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_366
timestamp 1608254825
transform 1 0 34776 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_387
timestamp 1608254825
transform 1 0 36708 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_379
timestamp 1608254825
transform 1 0 35972 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_230
timestamp 1608254825
transform 1 0 34776 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__a22oi_4  _1775_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 34868 0 -1 10336
box -38 -48 1602 592
use sky130_fd_sc_hd__a21o_4  _1501_
timestamp 1608254825
transform 1 0 34868 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_407
timestamp 1608254825
transform 1 0 38548 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_393
timestamp 1608254825
transform 1 0 37260 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_408
timestamp 1608254825
transform 1 0 38640 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_237
timestamp 1608254825
transform 1 0 37628 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2610_
timestamp 1608254825
transform 1 0 36892 0 1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__nor2_4  _1766_
timestamp 1608254825
transform 1 0 37720 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1499_
timestamp 1608254825
transform 1 0 38916 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1456_
timestamp 1608254825
transform 1 0 36892 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_414
timestamp 1608254825
transform 1 0 39192 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_416
timestamp 1608254825
transform 1 0 39376 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1608254825
transform -1 0 39836 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1608254825
transform -1 0 39836 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_19
timestamp 1608254825
transform 1 0 2852 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_11
timestamp 1608254825
transform 1 0 2116 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_3
timestamp 1608254825
transform 1 0 1380 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1608254825
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__and2_4  _1916_
timestamp 1608254825
transform 1 0 2208 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_15_37
timestamp 1608254825
transform 1 0 4508 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_26
timestamp 1608254825
transform 1 0 3496 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_0_0_m1_clk_local
timestamp 1608254825
transform 1 0 3220 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1906_
timestamp 1608254825
transform 1 0 4232 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_66
timestamp 1608254825
transform 1 0 7176 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_49
timestamp 1608254825
transform 1 0 5612 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_238
timestamp 1608254825
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _2258_
timestamp 1608254825
transform 1 0 6808 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_88
timestamp 1608254825
transform 1 0 9200 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_80
timestamp 1608254825
transform 1 0 8464 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_70
timestamp 1608254825
transform 1 0 7544 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_4  _2154_
timestamp 1608254825
transform 1 0 7636 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _2150_
timestamp 1608254825
transform 1 0 8832 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_101
timestamp 1608254825
transform 1 0 10396 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_4  _2174_
timestamp 1608254825
transform 1 0 11132 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_4  _1845_
timestamp 1608254825
transform 1 0 9568 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_15_136
timestamp 1608254825
transform 1 0 13616 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_118
timestamp 1608254825
transform 1 0 11960 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_239
timestamp 1608254825
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_4  _2219_
timestamp 1608254825
transform 1 0 12420 0 1 10336
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_15_152
timestamp 1608254825
transform 1 0 15088 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_4  _1749_
timestamp 1608254825
transform 1 0 13984 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _1630_
timestamp 1608254825
transform 1 0 15456 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_179
timestamp 1608254825
transform 1 0 17572 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_164
timestamp 1608254825
transform 1 0 16192 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_160
timestamp 1608254825
transform 1 0 15824 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_4  _2300_
timestamp 1608254825
transform 1 0 16284 0 1 10336
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_1  FILLER_15_192
timestamp 1608254825
transform 1 0 18768 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_188
timestamp 1608254825
transform 1 0 18400 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_240
timestamp 1608254825
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__a211o_4  _2225_
timestamp 1608254825
transform 1 0 18860 0 1 10336
box -38 -48 1326 592
use sky130_fd_sc_hd__buf_2  _1703_
timestamp 1608254825
transform 1 0 18032 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_215
timestamp 1608254825
transform 1 0 20884 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_207
timestamp 1608254825
transform 1 0 20148 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_4  _1752_
timestamp 1608254825
transform 1 0 20976 0 1 10336
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_8  FILLER_15_248
timestamp 1608254825
transform 1 0 23920 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_15_238
timestamp 1608254825
transform 1 0 23000 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_230
timestamp 1608254825
transform 1 0 22264 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_241
timestamp 1608254825
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _2123_
timestamp 1608254825
transform 1 0 22632 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2119_
timestamp 1608254825
transform 1 0 23644 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _2395_
timestamp 1608254825
transform 1 0 24656 0 1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_15_296
timestamp 1608254825
transform 1 0 28336 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_279
timestamp 1608254825
transform 1 0 26772 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_275
timestamp 1608254825
transform 1 0 26404 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_4  _2317_
timestamp 1608254825
transform 1 0 26864 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_15_304
timestamp 1608254825
transform 1 0 29072 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_242
timestamp 1608254825
transform 1 0 29164 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _2318_
timestamp 1608254825
transform 1 0 29256 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_15_339
timestamp 1608254825
transform 1 0 32292 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_322
timestamp 1608254825
transform 1 0 30728 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_4  _1463_
timestamp 1608254825
transform 1 0 31096 0 1 10336
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_3  FILLER_15_363
timestamp 1608254825
transform 1 0 34500 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_356
timestamp 1608254825
transform 1 0 33856 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_10_0_addressalyzerBlock.SPI_CLK
timestamp 1608254825
transform 1 0 34224 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_4  _1517_
timestamp 1608254825
transform 1 0 32660 0 1 10336
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_15_374
timestamp 1608254825
transform 1 0 35512 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_15_367
timestamp 1608254825
transform 1 0 34868 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_243
timestamp 1608254825
transform 1 0 34776 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1481_
timestamp 1608254825
transform 1 0 35144 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_4  _1479_
timestamp 1608254825
transform 1 0 35880 0 1 10336
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_15_391
timestamp 1608254825
transform 1 0 37076 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2611_
timestamp 1608254825
transform 1 0 37444 0 1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_15_414
timestamp 1608254825
transform 1 0 39192 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1608254825
transform -1 0 39836 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_16_15
timestamp 1608254825
transform 1 0 2484 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_3
timestamp 1608254825
transform 1 0 1380 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1608254825
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_4  _1907_
timestamp 1608254825
transform 1 0 2760 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_16_39
timestamp 1608254825
transform 1 0 4692 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_32
timestamp 1608254825
transform 1 0 4048 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_27
timestamp 1608254825
transform 1 0 3588 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_m1_clk_local
timestamp 1608254825
transform 1 0 4416 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_244
timestamp 1608254825
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__o32ai_4  _2259_
timestamp 1608254825
transform 1 0 5244 0 -1 11424
box -38 -48 2062 592
use sky130_fd_sc_hd__decap_4  FILLER_16_67
timestamp 1608254825
transform 1 0 7268 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_80
timestamp 1608254825
transform 1 0 8464 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_4  _2177_
timestamp 1608254825
transform 1 0 7636 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_16_109
timestamp 1608254825
transform 1 0 11132 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_102
timestamp 1608254825
transform 1 0 10488 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_245
timestamp 1608254825
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_4  _2221_
timestamp 1608254825
transform 1 0 11500 0 -1 11424
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_4  _2151_
timestamp 1608254825
transform 1 0 9660 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1623_
timestamp 1608254825
transform 1 0 10856 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_126
timestamp 1608254825
transform 1 0 12696 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_4  _1753_
timestamp 1608254825
transform 1 0 13064 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_158
timestamp 1608254825
transform 1 0 15640 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_149
timestamp 1608254825
transform 1 0 14812 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_142
timestamp 1608254825
transform 1 0 14168 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_246
timestamp 1608254825
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1941_
timestamp 1608254825
transform 1 0 14536 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1616_
timestamp 1608254825
transform 1 0 15272 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2407_
timestamp 1608254825
transform 1 0 16192 0 -1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_16_197
timestamp 1608254825
transform 1 0 19228 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_187
timestamp 1608254825
transform 1 0 18308 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_183
timestamp 1608254825
transform 1 0 17940 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_4  _2203_
timestamp 1608254825
transform 1 0 18400 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_4  _2158_
timestamp 1608254825
transform 1 0 19596 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_16_219
timestamp 1608254825
transform 1 0 21252 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_215
timestamp 1608254825
transform 1 0 20884 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_210
timestamp 1608254825
transform 1 0 20424 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_247
timestamp 1608254825
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _1751_
timestamp 1608254825
transform 1 0 21344 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_16_247
timestamp 1608254825
transform 1 0 23828 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_16_229
timestamp 1608254825
transform 1 0 22172 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_4  _2134_
timestamp 1608254825
transform 1 0 22540 0 -1 11424
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_16_271
timestamp 1608254825
transform 1 0 26036 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_4  _2320_
timestamp 1608254825
transform 1 0 24564 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_16_296
timestamp 1608254825
transform 1 0 28336 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_276
timestamp 1608254825
transform 1 0 26496 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_248
timestamp 1608254825
transform 1 0 26404 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2396_
timestamp 1608254825
transform 1 0 26588 0 -1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__xor2_4  _1767_
timestamp 1608254825
transform 1 0 28704 0 -1 11424
box -38 -48 2062 592
use sky130_fd_sc_hd__fill_2  FILLER_16_337
timestamp 1608254825
transform 1 0 32108 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_332
timestamp 1608254825
transform 1 0 31648 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_322
timestamp 1608254825
transform 1 0 30728 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_249
timestamp 1608254825
transform 1 0 32016 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__a22oi_4  _1776_
timestamp 1608254825
transform 1 0 32292 0 -1 11424
box -38 -48 1602 592
use sky130_fd_sc_hd__buf_2  _1461_
timestamp 1608254825
transform 1 0 31280 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_356
timestamp 1608254825
transform 1 0 33856 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__a22oi_4  _1774_
timestamp 1608254825
transform 1 0 34224 0 -1 11424
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_16_377
timestamp 1608254825
transform 1 0 35788 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__and4_4  _1777_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 36156 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_16_411
timestamp 1608254825
transform 1 0 38916 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_396
timestamp 1608254825
transform 1 0 37536 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_390
timestamp 1608254825
transform 1 0 36984 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_250
timestamp 1608254825
transform 1 0 37628 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_4  _1464_
timestamp 1608254825
transform 1 0 37720 0 -1 11424
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_1  FILLER_16_417
timestamp 1608254825
transform 1 0 39468 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1608254825
transform -1 0 39836 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_17_15
timestamp 1608254825
transform 1 0 2484 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1608254825
transform 1 0 1380 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1608254825
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _2540_
timestamp 1608254825
transform 1 0 3036 0 1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_17_40
timestamp 1608254825
transform 1 0 4784 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_68
timestamp 1608254825
transform 1 0 7360 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_17_62
timestamp 1608254825
transform 1 0 6808 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_57
timestamp 1608254825
transform 1 0 6348 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_52
timestamp 1608254825
transform 1 0 5888 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_251
timestamp 1608254825
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1944_
timestamp 1608254825
transform 1 0 7084 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1910_
timestamp 1608254825
transform 1 0 6072 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_86
timestamp 1608254825
transform 1 0 9016 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_4  _2156_
timestamp 1608254825
transform 1 0 7728 0 1 11424
box -38 -48 1326 592
use sky130_fd_sc_hd__nand3_4  _2153_
timestamp 1608254825
transform 1 0 9384 0 1 11424
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_17_104
timestamp 1608254825
transform 1 0 10672 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_4  _2196_
timestamp 1608254825
transform 1 0 11040 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_17_135
timestamp 1608254825
transform 1 0 13524 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_121
timestamp 1608254825
transform 1 0 12236 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_117
timestamp 1608254825
transform 1 0 11868 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_252
timestamp 1608254825
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__a21o_4  _2222_
timestamp 1608254825
transform 1 0 12420 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_159
timestamp 1608254825
transform 1 0 15732 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_142
timestamp 1608254825
transform 1 0 14168 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2243_
timestamp 1608254825
transform 1 0 13892 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_4  _2226_
timestamp 1608254825
transform 1 0 14536 0 1 11424
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_6  FILLER_17_177
timestamp 1608254825
transform 1 0 17388 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_163
timestamp 1608254825
transform 1 0 16100 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_4  _2301_
timestamp 1608254825
transform 1 0 16192 0 1 11424
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_17_198
timestamp 1608254825
transform 1 0 19320 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_188
timestamp 1608254825
transform 1 0 18400 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_184
timestamp 1608254825
transform 1 0 18032 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_253
timestamp 1608254825
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _2181_
timestamp 1608254825
transform 1 0 18492 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_4  _2159_
timestamp 1608254825
transform 1 0 19688 0 1 11424
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_8  FILLER_17_223
timestamp 1608254825
transform 1 0 21620 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_17_216
timestamp 1608254825
transform 1 0 20976 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1632_
timestamp 1608254825
transform 1 0 21344 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_248
timestamp 1608254825
transform 1 0 23920 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_243
timestamp 1608254825
transform 1 0 23460 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_237
timestamp 1608254825
transform 1 0 22908 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_17_231
timestamp 1608254825
transform 1 0 22356 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_254
timestamp 1608254825
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _2120_
timestamp 1608254825
transform 1 0 22540 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1490_
timestamp 1608254825
transform 1 0 23644 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_268
timestamp 1608254825
transform 1 0 25760 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2397_
timestamp 1608254825
transform 1 0 26128 0 1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__a2bb2o_4  _2319_
timestamp 1608254825
transform 1 0 24288 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_17_291
timestamp 1608254825
transform 1 0 27876 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_313
timestamp 1608254825
transform 1 0 29900 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_306
timestamp 1608254825
transform 1 0 29256 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_301
timestamp 1608254825
transform 1 0 28796 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_297
timestamp 1608254825
transform 1 0 28428 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_255
timestamp 1608254825
transform 1 0 29164 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1764_
timestamp 1608254825
transform 1 0 28520 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1511_
timestamp 1608254825
transform 1 0 29624 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1503_
timestamp 1608254825
transform 1 0 30268 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_320
timestamp 1608254825
transform 1 0 30544 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2605_
timestamp 1608254825
transform 1 0 30912 0 1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_17_360
timestamp 1608254825
transform 1 0 34224 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_347
timestamp 1608254825
transform 1 0 33028 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_343
timestamp 1608254825
transform 1 0 32660 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_4  _1513_
timestamp 1608254825
transform 1 0 33120 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_387
timestamp 1608254825
transform 1 0 36708 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_381
timestamp 1608254825
transform 1 0 36156 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_256
timestamp 1608254825
transform 1 0 34776 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_4  _1772_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 34868 0 1 11424
box -38 -48 1326 592
use sky130_fd_sc_hd__a2111o_4  _1769_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 36800 0 1 11424
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_17_405
timestamp 1608254825
transform 1 0 38364 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1485_
timestamp 1608254825
transform 1 0 38732 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_417
timestamp 1608254825
transform 1 0 39468 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_413
timestamp 1608254825
transform 1 0 39100 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1608254825
transform -1 0 39836 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_14
timestamp 1608254825
transform 1 0 2392 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_9
timestamp 1608254825
transform 1 0 1932 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_3
timestamp 1608254825
transform 1 0 1380 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1608254825
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_4  _1911_
timestamp 1608254825
transform 1 0 2760 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _1901_
timestamp 1608254825
transform 1 0 2024 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_32
timestamp 1608254825
transform 1 0 4048 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_27
timestamp 1608254825
transform 1 0 3588 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_257
timestamp 1608254825
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2428_
timestamp 1608254825
transform 1 0 5152 0 -1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_18_67
timestamp 1608254825
transform 1 0 7268 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_63
timestamp 1608254825
transform 1 0 6900 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_4  _2179_
timestamp 1608254825
transform 1 0 7360 0 -1 12512
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_2  FILLER_18_90
timestamp 1608254825
transform 1 0 9384 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_82
timestamp 1608254825
transform 1 0 8648 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_18_105
timestamp 1608254825
transform 1 0 10764 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_258
timestamp 1608254825
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__a21o_4  _2180_
timestamp 1608254825
transform 1 0 11316 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__a21o_4  _2157_
timestamp 1608254825
transform 1 0 9660 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_129
timestamp 1608254825
transform 1 0 12972 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_123
timestamp 1608254825
transform 1 0 12420 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  _2422_
timestamp 1608254825
transform 1 0 13064 0 -1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_18_149
timestamp 1608254825
transform 1 0 14812 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_259
timestamp 1608254825
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__o32ai_4  _2272_
timestamp 1608254825
transform 1 0 15272 0 -1 12512
box -38 -48 2062 592
use sky130_fd_sc_hd__decap_4  FILLER_18_176
timestamp 1608254825
transform 1 0 17296 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _2262_
timestamp 1608254825
transform 1 0 17664 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_192
timestamp 1608254825
transform 1 0 18768 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_184
timestamp 1608254825
transform 1 0 18032 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_4  _2182_
timestamp 1608254825
transform 1 0 19136 0 -1 12512
box -38 -48 1326 592
use sky130_fd_sc_hd__buf_2  _1635_
timestamp 1608254825
transform 1 0 18400 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_215
timestamp 1608254825
transform 1 0 20884 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_210
timestamp 1608254825
transform 1 0 20424 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_260
timestamp 1608254825
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__o32ai_4  _2140_
timestamp 1608254825
transform 1 0 21252 0 -1 12512
box -38 -48 2062 592
use sky130_fd_sc_hd__decap_8  FILLER_18_248
timestamp 1608254825
transform 1 0 23920 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_18_241
timestamp 1608254825
transform 1 0 23276 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1960_
timestamp 1608254825
transform 1 0 23644 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_18_274
timestamp 1608254825
transform 1 0 26312 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_270
timestamp 1608254825
transform 1 0 25944 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_263
timestamp 1608254825
transform 1 0 25300 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2136_
timestamp 1608254825
transform 1 0 25668 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__and2_4  _1968_
timestamp 1608254825
transform 1 0 24656 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_18_294
timestamp 1608254825
transform 1 0 28152 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_286
timestamp 1608254825
transform 1 0 27416 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_279
timestamp 1608254825
transform 1 0 26772 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_261
timestamp 1608254825
transform 1 0 26404 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _2144_
timestamp 1608254825
transform 1 0 26496 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1771_
timestamp 1608254825
transform 1 0 27140 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1471_
timestamp 1608254825
transform 1 0 27784 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_317
timestamp 1608254825
transform 1 0 30268 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_310
timestamp 1608254825
transform 1 0 29624 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_302
timestamp 1608254825
transform 1 0 28888 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_addressalyzerBlock.SPI_CLK
timestamp 1608254825
transform 1 0 29992 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_4  _1523_
timestamp 1608254825
transform 1 0 30452 0 -1 12512
box -38 -48 1234 592
use sky130_fd_sc_hd__buf_2  _1472_
timestamp 1608254825
transform 1 0 29256 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1430_
timestamp 1608254825
transform 1 0 28520 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_342
timestamp 1608254825
transform 1 0 32568 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_337
timestamp 1608254825
transform 1 0 32108 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_332
timestamp 1608254825
transform 1 0 31648 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_262
timestamp 1608254825
transform 1 0 32016 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1484_
timestamp 1608254825
transform 1 0 32200 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_354
timestamp 1608254825
transform 1 0 33672 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_350
timestamp 1608254825
transform 1 0 33304 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_4  _1496_
timestamp 1608254825
transform 1 0 33764 0 -1 12512
box -38 -48 1234 592
use sky130_fd_sc_hd__buf_2  _1437_
timestamp 1608254825
transform 1 0 32936 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_387
timestamp 1608254825
transform 1 0 36708 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_376
timestamp 1608254825
transform 1 0 35696 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_368
timestamp 1608254825
transform 1 0 34960 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__and4_4  _1436_
timestamp 1608254825
transform 1 0 35880 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_18_398
timestamp 1608254825
transform 1 0 37720 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_395
timestamp 1608254825
transform 1 0 37444 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_263
timestamp 1608254825
transform 1 0 37628 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_4  _1465_
timestamp 1608254825
transform 1 0 37904 0 -1 12512
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_1  FILLER_18_417
timestamp 1608254825
transform 1 0 39468 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_413
timestamp 1608254825
transform 1 0 39100 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1608254825
transform -1 0 39836 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_13
timestamp 1608254825
transform 1 0 2300 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_3
timestamp 1608254825
transform 1 0 1380 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_22
timestamp 1608254825
transform 1 0 3128 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1608254825
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1608254825
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _2517_
timestamp 1608254825
transform 1 0 1380 0 1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__and2_4  _1970_
timestamp 1608254825
transform 1 0 1656 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _1957_
timestamp 1608254825
transform 1 0 2668 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_20_38
timestamp 1608254825
transform 1 0 4600 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_32
timestamp 1608254825
transform 1 0 4048 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_30
timestamp 1608254825
transform 1 0 3864 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_24
timestamp 1608254825
transform 1 0 3312 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_45
timestamp 1608254825
transform 1 0 5244 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_270
timestamp 1608254825
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2538_
timestamp 1608254825
transform 1 0 3496 0 1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _2423_
timestamp 1608254825
transform 1 0 4968 0 -1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  _1956_
timestamp 1608254825
transform 1 0 4232 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_61
timestamp 1608254825
transform 1 0 6716 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_65
timestamp 1608254825
transform 1 0 7084 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_60
timestamp 1608254825
transform 1 0 6624 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_56
timestamp 1608254825
transform 1 0 6256 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_264
timestamp 1608254825
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _1945_
timestamp 1608254825
transform 1 0 7084 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__and2_4  _1918_
timestamp 1608254825
transform 1 0 5612 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1746_
timestamp 1608254825
transform 1 0 6808 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_20_91
timestamp 1608254825
transform 1 0 9476 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_87
timestamp 1608254825
transform 1 0 9108 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_74
timestamp 1608254825
transform 1 0 7912 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_83
timestamp 1608254825
transform 1 0 8740 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_4  _2201_
timestamp 1608254825
transform 1 0 7452 0 1 12512
box -38 -48 1326 592
use sky130_fd_sc_hd__nand2_4  _2200_
timestamp 1608254825
transform 1 0 8280 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  _2155_
timestamp 1608254825
transform 1 0 9108 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_20_102
timestamp 1608254825
transform 1 0 10488 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_19_96
timestamp 1608254825
transform 1 0 9936 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_271
timestamp 1608254825
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__nand3_4  _2198_
timestamp 1608254825
transform 1 0 10672 0 1 12512
box -38 -48 1326 592
use sky130_fd_sc_hd__nand3_4  _2176_
timestamp 1608254825
transform 1 0 11224 0 -1 13600
box -38 -48 1326 592
use sky130_fd_sc_hd__nand2_4  _2152_
timestamp 1608254825
transform 1 0 9660 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_20_137
timestamp 1608254825
transform 1 0 13708 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_124
timestamp 1608254825
transform 1 0 12512 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_135
timestamp 1608254825
transform 1 0 13524 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_118
timestamp 1608254825
transform 1 0 11960 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_265
timestamp 1608254825
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__a21o_4  _2202_
timestamp 1608254825
transform 1 0 12420 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_4  _2197_
timestamp 1608254825
transform 1 0 12880 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_20_158
timestamp 1608254825
transform 1 0 15640 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_145
timestamp 1608254825
transform 1 0 14444 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_272
timestamp 1608254825
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__o32ai_4  _2271_
timestamp 1608254825
transform 1 0 14260 0 1 12512
box -38 -48 2062 592
use sky130_fd_sc_hd__buf_2  _1634_
timestamp 1608254825
transform 1 0 15272 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1628_
timestamp 1608254825
transform 1 0 14076 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_181
timestamp 1608254825
transform 1 0 17756 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_165
timestamp 1608254825
transform 1 0 16284 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_181
timestamp 1608254825
transform 1 0 17756 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_173
timestamp 1608254825
transform 1 0 17020 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_165
timestamp 1608254825
transform 1 0 16284 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_addressalyzerBlock.SPI_CLK
timestamp 1608254825
transform 1 0 16008 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_4  _2160_
timestamp 1608254825
transform 1 0 16560 0 -1 13600
box -38 -48 1234 592
use sky130_fd_sc_hd__buf_2  _1708_
timestamp 1608254825
transform 1 0 16652 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_205
timestamp 1608254825
transform 1 0 19964 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_198
timestamp 1608254825
transform 1 0 19320 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_200
timestamp 1608254825
transform 1 0 19504 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_184
timestamp 1608254825
transform 1 0 18032 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_266
timestamp 1608254825
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _2224_
timestamp 1608254825
transform 1 0 19872 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_4  _2205_
timestamp 1608254825
transform 1 0 18124 0 -1 13600
box -38 -48 1234 592
use sky130_fd_sc_hd__a211o_4  _2204_
timestamp 1608254825
transform 1 0 18216 0 1 12512
box -38 -48 1326 592
use sky130_fd_sc_hd__inv_2  _1533_
timestamp 1608254825
transform 1 0 19688 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_223
timestamp 1608254825
transform 1 0 21620 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_219
timestamp 1608254825
transform 1 0 21252 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_215
timestamp 1608254825
transform 1 0 20884 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_213
timestamp 1608254825
transform 1 0 20700 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_213
timestamp 1608254825
transform 1 0 20700 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_273
timestamp 1608254825
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2442_
timestamp 1608254825
transform 1 0 21252 0 1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_2  _1962_
timestamp 1608254825
transform 1 0 21344 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_4  _1961_
timestamp 1608254825
transform 1 0 21988 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_20_251
timestamp 1608254825
transform 1 0 24196 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_243
timestamp 1608254825
transform 1 0 23460 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_236
timestamp 1608254825
transform 1 0 22816 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_238
timestamp 1608254825
transform 1 0 23000 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_267
timestamp 1608254825
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2506_
timestamp 1608254825
transform 1 0 23644 0 1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_2  _1964_
timestamp 1608254825
transform 1 0 23184 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_20_274
timestamp 1608254825
transform 1 0 26312 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_268
timestamp 1608254825
transform 1 0 25760 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_261
timestamp 1608254825
transform 1 0 25116 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_271
timestamp 1608254825
transform 1 0 26036 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_264
timestamp 1608254825
transform 1 0 25392 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1966_
timestamp 1608254825
transform 1 0 25484 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_4  _1607_
timestamp 1608254825
transform 1 0 24288 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1420_
timestamp 1608254825
transform 1 0 25760 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_279
timestamp 1608254825
transform 1 0 26772 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_278
timestamp 1608254825
transform 1 0 26680 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_274
timestamp 1608254825
transform 1 0 26404 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2603_
timestamp 1608254825
transform 1 0 27140 0 -1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_2  _2138_
timestamp 1608254825
transform 1 0 26404 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1691_
timestamp 1608254825
transform 1 0 26496 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_4  _1540_
timestamp 1608254825
transform 1 0 27232 0 1 12512
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_1  FILLER_20_309
timestamp 1608254825
transform 1 0 29532 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_302
timestamp 1608254825
transform 1 0 28888 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_315
timestamp 1608254825
transform 1 0 30084 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_19_297
timestamp 1608254825
transform 1 0 28428 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_9_0_addressalyzerBlock.SPI_CLK
timestamp 1608254825
transform 1 0 29256 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_268
timestamp 1608254825
transform 1 0 29164 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__a41oi_4  _1518_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 29624 0 -1 13600
box -38 -48 2062 592
use sky130_fd_sc_hd__and4_4  _1483_
timestamp 1608254825
transform 1 0 29256 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_20_332
timestamp 1608254825
transform 1 0 31648 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_342
timestamp 1608254825
transform 1 0 32568 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_334
timestamp 1608254825
transform 1 0 31832 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_275
timestamp 1608254825
transform 1 0 32016 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_4  _1522_
timestamp 1608254825
transform 1 0 32108 0 -1 13600
box -38 -48 1234 592
use sky130_fd_sc_hd__o21ai_4  _1519_
timestamp 1608254825
transform 1 0 30636 0 1 12512
box -38 -48 1234 592
use sky130_fd_sc_hd__buf_2  _1433_
timestamp 1608254825
transform 1 0 32200 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_357
timestamp 1608254825
transform 1 0 33948 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_350
timestamp 1608254825
transform 1 0 33304 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_358
timestamp 1608254825
transform 1 0 34040 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_addressalyzerBlock.SPI_CLK
timestamp 1608254825
transform 1 0 33672 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_addressalyzerBlock.SPI_CLK
timestamp 1608254825
transform 1 0 32936 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__a41oi_4  _1495_
timestamp 1608254825
transform 1 0 34040 0 -1 13600
box -38 -48 2062 592
use sky130_fd_sc_hd__and4_4  _1494_
timestamp 1608254825
transform 1 0 33212 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_20_380
timestamp 1608254825
transform 1 0 36064 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_385
timestamp 1608254825
transform 1 0 36524 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_367
timestamp 1608254825
transform 1 0 34868 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_269
timestamp 1608254825
transform 1 0 34776 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__nand4_4  _1487_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 34960 0 1 12512
box -38 -48 1602 592
use sky130_fd_sc_hd__and4_4  _1457_
timestamp 1608254825
transform 1 0 36432 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_20_411
timestamp 1608254825
transform 1 0 38916 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_393
timestamp 1608254825
transform 1 0 37260 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_396
timestamp 1608254825
transform 1 0 37536 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_276
timestamp 1608254825
transform 1 0 37628 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _2114_
timestamp 1608254825
transform 1 0 36892 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_4  _1476_
timestamp 1608254825
transform 1 0 37720 0 -1 13600
box -38 -48 1234 592
use sky130_fd_sc_hd__o21ai_4  _1458_
timestamp 1608254825
transform 1 0 37904 0 1 12512
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_1  FILLER_20_417
timestamp 1608254825
transform 1 0 39468 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_417
timestamp 1608254825
transform 1 0 39468 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_413
timestamp 1608254825
transform 1 0 39100 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1608254825
transform -1 0 39836 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1608254825
transform -1 0 39836 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_3
timestamp 1608254825
transform 1 0 1380 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1608254825
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _2504_
timestamp 1608254825
transform 1 0 1564 0 1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_21_41
timestamp 1608254825
transform 1 0 4876 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_28
timestamp 1608254825
transform 1 0 3680 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_24
timestamp 1608254825
transform 1 0 3312 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_m1_clk_local
timestamp 1608254825
transform 1 0 3772 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_4  _2090_
timestamp 1608254825
transform 1 0 4048 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__and2_4  _1920_
timestamp 1608254825
transform 1 0 5244 0 1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_21_62
timestamp 1608254825
transform 1 0 6808 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_60
timestamp 1608254825
transform 1 0 6624 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_52
timestamp 1608254825
transform 1 0 5888 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_277
timestamp 1608254825
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_4  _2178_
timestamp 1608254825
transform 1 0 6992 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_21_73
timestamp 1608254825
transform 1 0 7820 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__o32ai_4  _2273_
timestamp 1608254825
transform 1 0 8188 0 1 13600
box -38 -48 2062 592
use sky130_fd_sc_hd__fill_2  FILLER_21_107
timestamp 1608254825
transform 1 0 10948 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_99
timestamp 1608254825
transform 1 0 10212 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_4  _2175_
timestamp 1608254825
transform 1 0 11132 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_21_123
timestamp 1608254825
transform 1 0 12420 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_118
timestamp 1608254825
transform 1 0 11960 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_278
timestamp 1608254825
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2404_
timestamp 1608254825
transform 1 0 12512 0 1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_21_143
timestamp 1608254825
transform 1 0 14260 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_4  _2306_
timestamp 1608254825
transform 1 0 14628 0 1 13600
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_1  FILLER_21_182
timestamp 1608254825
transform 1 0 17848 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_178
timestamp 1608254825
transform 1 0 17480 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_161
timestamp 1608254825
transform 1 0 15916 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_4  _2183_
timestamp 1608254825
transform 1 0 16284 0 1 13600
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_2  FILLER_21_184
timestamp 1608254825
transform 1 0 18032 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_279
timestamp 1608254825
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__o32ai_4  _2143_
timestamp 1608254825
transform 1 0 18216 0 1 13600
box -38 -48 2062 592
use sky130_fd_sc_hd__decap_4  FILLER_21_208
timestamp 1608254825
transform 1 0 20240 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__o32ai_4  _2141_
timestamp 1608254825
transform 1 0 20608 0 1 13600
box -38 -48 2062 592
use sky130_fd_sc_hd__fill_2  FILLER_21_242
timestamp 1608254825
transform 1 0 23368 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_234
timestamp 1608254825
transform 1 0 22632 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_280
timestamp 1608254825
transform 1 0 23552 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2505_
timestamp 1608254825
transform 1 0 23644 0 1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_21_264
timestamp 1608254825
transform 1 0 25392 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2604_
timestamp 1608254825
transform 1 0 25760 0 1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_21_295
timestamp 1608254825
transform 1 0 28244 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_287
timestamp 1608254825
transform 1 0 27508 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_306
timestamp 1608254825
transform 1 0 29256 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_301
timestamp 1608254825
transform 1 0 28796 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_281
timestamp 1608254825
transform 1 0 29164 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__a41oi_4  _1524_
timestamp 1608254825
transform 1 0 29440 0 1 13600
box -38 -48 2062 592
use sky130_fd_sc_hd__buf_2  _1431_
timestamp 1608254825
transform 1 0 28428 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_337
timestamp 1608254825
transform 1 0 32108 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_330
timestamp 1608254825
transform 1 0 31464 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__nand4_4  _1505_
timestamp 1608254825
transform 1 0 32476 0 1 13600
box -38 -48 1602 592
use sky130_fd_sc_hd__inv_2  _1447_
timestamp 1608254825
transform 1 0 31832 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_21_365
timestamp 1608254825
transform 1 0 34684 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_358
timestamp 1608254825
transform 1 0 34040 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_11_0_addressalyzerBlock.SPI_CLK
timestamp 1608254825
transform 1 0 34408 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_382
timestamp 1608254825
transform 1 0 36248 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_367
timestamp 1608254825
transform 1 0 34868 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_282
timestamp 1608254825
transform 1 0 34776 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__a41oi_4  _1475_
timestamp 1608254825
transform 1 0 36616 0 1 13600
box -38 -48 2062 592
use sky130_fd_sc_hd__and4_4  _1473_
timestamp 1608254825
transform 1 0 35420 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_21_408
timestamp 1608254825
transform 1 0 38640 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_416
timestamp 1608254825
transform 1 0 39376 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1608254825
transform -1 0 39836 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_22_22
timestamp 1608254825
transform 1 0 3128 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_18
timestamp 1608254825
transform 1 0 2760 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_3
timestamp 1608254825
transform 1 0 1380 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1608254825
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_4  _1965_
timestamp 1608254825
transform 1 0 1932 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_22_41
timestamp 1608254825
transform 1 0 4876 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_22_27
timestamp 1608254825
transform 1 0 3588 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_283
timestamp 1608254825
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _1967_
timestamp 1608254825
transform 1 0 4048 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _1255_
timestamp 1608254825
transform 1 0 3220 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_22_49
timestamp 1608254825
transform 1 0 5612 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _2421_
timestamp 1608254825
transform 1 0 5888 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_22_91
timestamp 1608254825
transform 1 0 9476 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_85
timestamp 1608254825
transform 1 0 8924 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_75
timestamp 1608254825
transform 1 0 8004 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_71
timestamp 1608254825
transform 1 0 7636 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_4  _1947_
timestamp 1608254825
transform 1 0 8096 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_22_93
timestamp 1608254825
transform 1 0 9660 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_284
timestamp 1608254825
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2419_
timestamp 1608254825
transform 1 0 10212 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_22_126
timestamp 1608254825
transform 1 0 12696 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_118
timestamp 1608254825
transform 1 0 11960 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_4  _2307_
timestamp 1608254825
transform 1 0 12880 0 -1 14688
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_22_149
timestamp 1608254825
transform 1 0 14812 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_141
timestamp 1608254825
transform 1 0 14076 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_285
timestamp 1608254825
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2406_
timestamp 1608254825
transform 1 0 15272 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  _2264_
timestamp 1608254825
transform 1 0 14444 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_173
timestamp 1608254825
transform 1 0 17020 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _2440_
timestamp 1608254825
transform 1 0 17756 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_22_200
timestamp 1608254825
transform 1 0 19504 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1601_
timestamp 1608254825
transform 1 0 19872 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_208
timestamp 1608254825
transform 1 0 20240 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_286
timestamp 1608254825
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2441_
timestamp 1608254825
transform 1 0 20884 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_22_242
timestamp 1608254825
transform 1 0 23368 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_234
timestamp 1608254825
transform 1 0 22632 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__and4_4  _2312_
timestamp 1608254825
transform 1 0 23736 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _2121_
timestamp 1608254825
transform 1 0 23000 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_271
timestamp 1608254825
transform 1 0 26036 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_255
timestamp 1608254825
transform 1 0 24564 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_4  _1535_
timestamp 1608254825
transform 1 0 24932 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_289
timestamp 1608254825
transform 1 0 27692 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_287
timestamp 1608254825
transform 1 0 26404 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1555_
timestamp 1608254825
transform 1 0 28060 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_4  _1532_
timestamp 1608254825
transform 1 0 26496 0 -1 14688
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_22_315
timestamp 1608254825
transform 1 0 30084 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_301
timestamp 1608254825
transform 1 0 28796 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_297
timestamp 1608254825
transform 1 0 28428 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_4  _1525_
timestamp 1608254825
transform 1 0 28888 0 -1 14688
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_4  _1429_
timestamp 1608254825
transform 1 0 30452 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_22_328
timestamp 1608254825
transform 1 0 31280 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_288
timestamp 1608254825
transform 1 0 32016 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__a21o_4  _1509_
timestamp 1608254825
transform 1 0 32108 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_349
timestamp 1608254825
transform 1 0 33212 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__a41o_4  _1508_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 33580 0 -1 14688
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_22_370
timestamp 1608254825
transform 1 0 35144 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2450_
timestamp 1608254825
transform 1 0 35512 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_22_407
timestamp 1608254825
transform 1 0 38548 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_393
timestamp 1608254825
transform 1 0 37260 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_289
timestamp 1608254825
transform 1 0 37628 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1504_
timestamp 1608254825
transform 1 0 38916 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__and4_4  _1438_
timestamp 1608254825
transform 1 0 37720 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_22_414
timestamp 1608254825
transform 1 0 39192 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1608254825
transform -1 0 39836 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_23_22
timestamp 1608254825
transform 1 0 3128 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1608254825
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _2515_
timestamp 1608254825
transform 1 0 1380 0 1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_23_30
timestamp 1608254825
transform 1 0 3864 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _2469_
timestamp 1608254825
transform 1 0 4048 0 1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_23_62
timestamp 1608254825
transform 1 0 6808 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_59
timestamp 1608254825
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_51
timestamp 1608254825
transform 1 0 5796 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_290
timestamp 1608254825
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _1949_
timestamp 1608254825
transform 1 0 6992 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_23_73
timestamp 1608254825
transform 1 0 7820 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__o32ai_4  _2274_
timestamp 1608254825
transform 1 0 8372 0 1 14688
box -38 -48 2062 592
use sky130_fd_sc_hd__decap_4  FILLER_23_109
timestamp 1608254825
transform 1 0 11132 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_101
timestamp 1608254825
transform 1 0 10396 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1943_
timestamp 1608254825
transform 1 0 11500 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1618_
timestamp 1608254825
transform 1 0 10764 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_127
timestamp 1608254825
transform 1 0 12788 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_121
timestamp 1608254825
transform 1 0 12236 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_117
timestamp 1608254825
transform 1 0 11868 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_m1_clk_local
timestamp 1608254825
transform 1 0 13340 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_291
timestamp 1608254825
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__nand3_4  _2308_
timestamp 1608254825
transform 1 0 13616 0 1 14688
box -38 -48 1326 592
use sky130_fd_sc_hd__buf_2  _2270_
timestamp 1608254825
transform 1 0 12420 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_158
timestamp 1608254825
transform 1 0 15640 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_150
timestamp 1608254825
transform 1 0 14904 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_182
timestamp 1608254825
transform 1 0 17848 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_174
timestamp 1608254825
transform 1 0 17112 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__nand3_4  _2302_
timestamp 1608254825
transform 1 0 15824 0 1 14688
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_23_188
timestamp 1608254825
transform 1 0 18400 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_292
timestamp 1608254825
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _2297_
timestamp 1608254825
transform 1 0 18032 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__o32ai_4  _2145_
timestamp 1608254825
transform 1 0 18768 0 1 14688
box -38 -48 2062 592
use sky130_fd_sc_hd__decap_4  FILLER_23_221
timestamp 1608254825
transform 1 0 21436 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_214
timestamp 1608254825
transform 1 0 20792 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_4  _1963_
timestamp 1608254825
transform 1 0 21804 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1603_
timestamp 1608254825
transform 1 0 21160 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_242
timestamp 1608254825
transform 1 0 23368 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_234
timestamp 1608254825
transform 1 0 22632 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_293
timestamp 1608254825
transform 1 0 23552 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__and4_4  _2238_
timestamp 1608254825
transform 1 0 23644 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_23_262
timestamp 1608254825
transform 1 0 25208 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_254
timestamp 1608254825
transform 1 0 24472 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1695_
timestamp 1608254825
transform 1 0 24840 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_4  _1536_
timestamp 1608254825
transform 1 0 25576 0 1 14688
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_1  FILLER_23_287
timestamp 1608254825
transform 1 0 27508 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_279
timestamp 1608254825
transform 1 0 26772 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_4  _1539_
timestamp 1608254825
transform 1 0 27600 0 1 14688
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_2  FILLER_23_306
timestamp 1608254825
transform 1 0 29256 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_301
timestamp 1608254825
transform 1 0 28796 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_294
timestamp 1608254825
transform 1 0 29164 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__nor3_4  _1482_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 29440 0 1 14688
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_1  FILLER_23_338
timestamp 1608254825
transform 1 0 32200 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_334
timestamp 1608254825
transform 1 0 31832 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_321
timestamp 1608254825
transform 1 0 30636 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_4  _1506_
timestamp 1608254825
transform 1 0 32292 0 1 14688
box -38 -48 1234 592
use sky130_fd_sc_hd__and4_4  _1432_
timestamp 1608254825
transform 1 0 31004 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_23_362
timestamp 1608254825
transform 1 0 34408 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_352
timestamp 1608254825
transform 1 0 33488 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _1486_
timestamp 1608254825
transform 1 0 34040 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_367
timestamp 1608254825
transform 1 0 34868 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_295
timestamp 1608254825
transform 1 0 34776 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__o32ai_4  _1491_
timestamp 1608254825
transform 1 0 35236 0 1 14688
box -38 -48 2062 592
use sky130_fd_sc_hd__decap_4  FILLER_23_402
timestamp 1608254825
transform 1 0 38088 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_397
timestamp 1608254825
transform 1 0 37628 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_393
timestamp 1608254825
transform 1 0 37260 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__and2_4  _2113_
timestamp 1608254825
transform 1 0 38456 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _1470_
timestamp 1608254825
transform 1 0 37720 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_417
timestamp 1608254825
transform 1 0 39468 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_413
timestamp 1608254825
transform 1 0 39100 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1608254825
transform -1 0 39836 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_24_21
timestamp 1608254825
transform 1 0 3036 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_24_11
timestamp 1608254825
transform 1 0 2116 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_24_3
timestamp 1608254825
transform 1 0 1380 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1608254825
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__and2_4  _1959_
timestamp 1608254825
transform 1 0 2392 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1608254825
transform 1 0 3588 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_m1_clk_local
timestamp 1608254825
transform 1 0 3680 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_296
timestamp 1608254825
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2503_
timestamp 1608254825
transform 1 0 4048 0 -1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_24_57
timestamp 1608254825
transform 1 0 6348 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_51
timestamp 1608254825
transform 1 0 5796 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  _2420_
timestamp 1608254825
transform 1 0 6440 0 -1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_24_91
timestamp 1608254825
transform 1 0 9476 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_85
timestamp 1608254825
transform 1 0 8924 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_77
timestamp 1608254825
transform 1 0 8188 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1254_
timestamp 1608254825
transform 1 0 8556 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_96
timestamp 1608254825
transform 1 0 9936 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_297
timestamp 1608254825
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__o32ai_4  _2275_
timestamp 1608254825
transform 1 0 10304 0 -1 15776
box -38 -48 2062 592
use sky130_fd_sc_hd__inv_2  _1946_
timestamp 1608254825
transform 1 0 9660 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_122
timestamp 1608254825
transform 1 0 12328 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2403_
timestamp 1608254825
transform 1 0 12696 0 -1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_24_154
timestamp 1608254825
transform 1 0 15272 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_145
timestamp 1608254825
transform 1 0 14444 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_298
timestamp 1608254825
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_4  _2303_
timestamp 1608254825
transform 1 0 15456 0 -1 15776
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_24_169
timestamp 1608254825
transform 1 0 16652 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_4  _2304_
timestamp 1608254825
transform 1 0 17020 0 -1 15776
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_24_187
timestamp 1608254825
transform 1 0 18308 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2439_
timestamp 1608254825
transform 1 0 18676 0 -1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_24_219
timestamp 1608254825
transform 1 0 21252 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_215
timestamp 1608254825
transform 1 0 20884 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_210
timestamp 1608254825
transform 1 0 20424 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_299
timestamp 1608254825
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__a41o_4  _2139_
timestamp 1608254825
transform 1 0 21620 0 -1 15776
box -38 -48 1602 592
use sky130_fd_sc_hd__inv_2  _1562_
timestamp 1608254825
transform 1 0 20976 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_240
timestamp 1608254825
transform 1 0 23184 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__a41o_4  _2248_
timestamp 1608254825
transform 1 0 23552 0 -1 15776
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_6  FILLER_24_269
timestamp 1608254825
transform 1 0 25852 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_261
timestamp 1608254825
transform 1 0 25116 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1696_
timestamp 1608254825
transform 1 0 25484 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_296
timestamp 1608254825
transform 1 0 28336 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_279
timestamp 1608254825
transform 1 0 26772 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_300
timestamp 1608254825
transform 1 0 26404 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_4  _1543_
timestamp 1608254825
transform 1 0 27140 0 -1 15776
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _1466_
timestamp 1608254825
transform 1 0 26496 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_24_302
timestamp 1608254825
transform 1 0 28888 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__nor4_4  _1469_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 28980 0 -1 15776
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_2  FILLER_24_337
timestamp 1608254825
transform 1 0 32108 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_328
timestamp 1608254825
transform 1 0 31280 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_24_320
timestamp 1608254825
transform 1 0 30544 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_301
timestamp 1608254825
transform 1 0 32016 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1537_
timestamp 1608254825
transform 1 0 30912 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_4  _1507_
timestamp 1608254825
transform 1 0 32292 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_24_348
timestamp 1608254825
transform 1 0 33120 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2607_
timestamp 1608254825
transform 1 0 33488 0 -1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_24_371
timestamp 1608254825
transform 1 0 35236 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__a22oi_4  _1492_
timestamp 1608254825
transform 1 0 35604 0 -1 15776
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_24_407
timestamp 1608254825
transform 1 0 38548 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_396
timestamp 1608254825
transform 1 0 37536 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_392
timestamp 1608254825
transform 1 0 37168 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_302
timestamp 1608254825
transform 1 0 37628 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1529_
timestamp 1608254825
transform 1 0 38916 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_4  _1493_
timestamp 1608254825
transform 1 0 37720 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_24_414
timestamp 1608254825
transform 1 0 39192 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1608254825
transform -1 0 39836 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_22
timestamp 1608254825
transform 1 0 3128 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1608254825
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _2507_
timestamp 1608254825
transform 1 0 1380 0 1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_25_34
timestamp 1608254825
transform 1 0 4232 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_26
timestamp 1608254825
transform 1 0 3496 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2644_
timestamp 1608254825
transform 1 0 4600 0 1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__and2_4  _1971_
timestamp 1608254825
transform 1 0 3588 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_25_57
timestamp 1608254825
transform 1 0 6348 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_303
timestamp 1608254825
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _2088_
timestamp 1608254825
transform 1 0 6808 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_25_77
timestamp 1608254825
transform 1 0 8188 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_69
timestamp 1608254825
transform 1 0 7452 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _2516_
timestamp 1608254825
transform 1 0 8372 0 1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_25_109
timestamp 1608254825
transform 1 0 11132 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_98
timestamp 1608254825
transform 1 0 10120 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__and2_4  _1958_
timestamp 1608254825
transform 1 0 10488 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1948_
timestamp 1608254825
transform 1 0 11500 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_25_123
timestamp 1608254825
transform 1 0 12420 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_25_116
timestamp 1608254825
transform 1 0 11776 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_304
timestamp 1608254825
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_4  _2309_
timestamp 1608254825
transform 1 0 12696 0 1 15776
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_1  FILLER_25_145
timestamp 1608254825
transform 1 0 14444 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_139
timestamp 1608254825
transform 1 0 13892 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  _2447_
timestamp 1608254825
transform 1 0 14536 0 1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_25_181
timestamp 1608254825
transform 1 0 17756 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_173
timestamp 1608254825
transform 1 0 17020 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_25_165
timestamp 1608254825
transform 1 0 16284 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _2291_
timestamp 1608254825
transform 1 0 16652 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_203
timestamp 1608254825
transform 1 0 19780 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_305
timestamp 1608254825
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2405_
timestamp 1608254825
transform 1 0 18032 0 1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_25_217
timestamp 1608254825
transform 1 0 21068 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_207
timestamp 1608254825
transform 1 0 20148 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__a41o_4  _2263_
timestamp 1608254825
transform 1 0 21436 0 1 15776
box -38 -48 1602 592
use sky130_fd_sc_hd__nor2_4  _2137_
timestamp 1608254825
transform 1 0 20240 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_25_238
timestamp 1608254825
transform 1 0 23000 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_306
timestamp 1608254825
transform 1 0 23552 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__a41o_4  _2310_
timestamp 1608254825
transform 1 0 23644 0 1 15776
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_25_262
timestamp 1608254825
transform 1 0 25208 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_4  _1578_
timestamp 1608254825
transform 1 0 25576 0 1 15776
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_8  FILLER_25_296
timestamp 1608254825
transform 1 0 28336 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_25_279
timestamp 1608254825
transform 1 0 26772 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_4  _1588_
timestamp 1608254825
transform 1 0 27140 0 1 15776
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_25_315
timestamp 1608254825
transform 1 0 30084 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_310
timestamp 1608254825
transform 1 0 29624 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_306
timestamp 1608254825
transform 1 0 29256 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_304
timestamp 1608254825
transform 1 0 29072 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_307
timestamp 1608254825
transform 1 0 29164 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_4  _1547_
timestamp 1608254825
transform 1 0 30452 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _1468_
timestamp 1608254825
transform 1 0 29716 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_339
timestamp 1608254825
transform 1 0 32292 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_331
timestamp 1608254825
transform 1 0 31556 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1460_
timestamp 1608254825
transform 1 0 31924 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_358
timestamp 1608254825
transform 1 0 34040 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_4  _1510_
timestamp 1608254825
transform 1 0 32844 0 1 15776
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_25_384
timestamp 1608254825
transform 1 0 36432 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_371
timestamp 1608254825
transform 1 0 35236 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_367
timestamp 1608254825
transform 1 0 34868 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_308
timestamp 1608254825
transform 1 0 34776 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__a21o_4  _1489_
timestamp 1608254825
transform 1 0 35328 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1435_
timestamp 1608254825
transform 1 0 36800 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_391
timestamp 1608254825
transform 1 0 37076 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2451_
timestamp 1608254825
transform 1 0 37444 0 1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_25_414
timestamp 1608254825
transform 1 0 39192 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1608254825
transform -1 0 39836 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_26_11
timestamp 1608254825
transform 1 0 2116 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_26_3
timestamp 1608254825
transform 1 0 1380 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1608254825
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1608254825
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_16
timestamp 1608254825
transform 1 0 2576 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_20
timestamp 1608254825
transform 1 0 2944 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_2_0_m1_clk_local
timestamp 1608254825
transform 1 0 2392 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1290_
timestamp 1608254825
transform 1 0 2668 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_4  _1289_
timestamp 1608254825
transform 1 0 2944 0 1 16864
box -38 -48 1326 592
use sky130_fd_sc_hd__nor3_4  _1286_
timestamp 1608254825
transform 1 0 1380 0 1 16864
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_6  FILLER_27_34
timestamp 1608254825
transform 1 0 4232 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_27
timestamp 1608254825
transform 1 0 3588 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_309
timestamp 1608254825
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2639_
timestamp 1608254825
transform 1 0 4048 0 -1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_2  _1264_
timestamp 1608254825
transform 1 0 3312 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__nand4_4  _1262_
timestamp 1608254825
transform 1 0 4784 0 1 16864
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_8  FILLER_27_65
timestamp 1608254825
transform 1 0 7084 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_27_57
timestamp 1608254825
transform 1 0 6348 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_51
timestamp 1608254825
transform 1 0 5796 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_316
timestamp 1608254825
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__nand3_4  _1263_
timestamp 1608254825
transform 1 0 6164 0 -1 16864
box -38 -48 1326 592
use sky130_fd_sc_hd__inv_2  _1251_
timestamp 1608254825
transform 1 0 6808 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_90
timestamp 1608254825
transform 1 0 9384 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_82
timestamp 1608254825
transform 1 0 8648 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_69
timestamp 1608254825
transform 1 0 7452 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2643_
timestamp 1608254825
transform 1 0 7820 0 1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__and3_4  _1271_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 7820 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_27_103
timestamp 1608254825
transform 1 0 10580 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_27_92
timestamp 1608254825
transform 1 0 9568 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_97
timestamp 1608254825
transform 1 0 10028 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_93
timestamp 1608254825
transform 1 0 9660 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_310
timestamp 1608254825
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2566_
timestamp 1608254825
transform 1 0 10120 0 -1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__and2_4  _1882_
timestamp 1608254825
transform 1 0 11316 0 1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _1875_
timestamp 1608254825
transform 1 0 9936 0 1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_27_137
timestamp 1608254825
transform 1 0 13708 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_123
timestamp 1608254825
transform 1 0 12420 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_118
timestamp 1608254825
transform 1 0 11960 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_125
timestamp 1608254825
transform 1 0 12604 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_117
timestamp 1608254825
transform 1 0 11868 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_317
timestamp 1608254825
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2448_
timestamp 1608254825
transform 1 0 12788 0 -1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__o21ai_4  _1615_
timestamp 1608254825
transform 1 0 12512 0 1 16864
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_27_146
timestamp 1608254825
transform 1 0 14536 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_141
timestamp 1608254825
transform 1 0 14076 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_154
timestamp 1608254825
transform 1 0 15272 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_152
timestamp 1608254825
transform 1 0 15088 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_146
timestamp 1608254825
transform 1 0 14536 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_311
timestamp 1608254825
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _2292_
timestamp 1608254825
transform 1 0 14168 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__and2_4  _1883_
timestamp 1608254825
transform 1 0 15456 0 -1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_4  _1718_
timestamp 1608254825
transform 1 0 14904 0 1 16864
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_1  FILLER_27_182
timestamp 1608254825
transform 1 0 17848 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_176
timestamp 1608254825
transform 1 0 17296 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_163
timestamp 1608254825
transform 1 0 16100 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_163
timestamp 1608254825
transform 1 0 16100 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_4  _2305_
timestamp 1608254825
transform 1 0 16836 0 -1 16864
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_4  _1701_
timestamp 1608254825
transform 1 0 16468 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_27_192
timestamp 1608254825
transform 1 0 18768 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_188
timestamp 1608254825
transform 1 0 18400 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_192
timestamp 1608254825
transform 1 0 18768 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_184
timestamp 1608254825
transform 1 0 18032 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_318
timestamp 1608254825
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2449_
timestamp 1608254825
transform 1 0 18860 0 1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  _1874_
timestamp 1608254825
transform 1 0 18032 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_4  _1602_
timestamp 1608254825
transform 1 0 19136 0 -1 16864
box -38 -48 1326 592
use sky130_fd_sc_hd__buf_2  _1534_
timestamp 1608254825
transform 1 0 18400 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_218
timestamp 1608254825
transform 1 0 21160 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_212
timestamp 1608254825
transform 1 0 20608 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_26_215
timestamp 1608254825
transform 1 0 20884 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_210
timestamp 1608254825
transform 1 0 20424 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_312
timestamp 1608254825
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__nor4_4  _2289_
timestamp 1608254825
transform 1 0 21252 0 1 16864
box -38 -48 1602 592
use sky130_fd_sc_hd__nor3_4  _2245_
timestamp 1608254825
transform 1 0 21160 0 -1 16864
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_8  FILLER_27_236
timestamp 1608254825
transform 1 0 22816 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_231
timestamp 1608254825
transform 1 0 22356 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1580_
timestamp 1608254825
transform 1 0 22724 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_245
timestamp 1608254825
transform 1 0 23644 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_243
timestamp 1608254825
transform 1 0 23460 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_239
timestamp 1608254825
transform 1 0 23092 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_319
timestamp 1608254825
transform 1 0 23552 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_4  _1600_
timestamp 1608254825
transform 1 0 23552 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_27_249
timestamp 1608254825
transform 1 0 24012 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1581_
timestamp 1608254825
transform 1 0 24104 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_261
timestamp 1608254825
transform 1 0 25116 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_254
timestamp 1608254825
transform 1 0 24472 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_271
timestamp 1608254825
transform 1 0 26036 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_264
timestamp 1608254825
transform 1 0 25392 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_253
timestamp 1608254825
transform 1 0 24380 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__and2_4  _1969_
timestamp 1608254825
transform 1 0 24748 0 -1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_4  _1599_
timestamp 1608254825
transform 1 0 25484 0 1 16864
box -38 -48 1326 592
use sky130_fd_sc_hd__inv_2  _1549_
timestamp 1608254825
transform 1 0 24840 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1527_
timestamp 1608254825
transform 1 0 25760 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_27_279
timestamp 1608254825
transform 1 0 26772 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_289
timestamp 1608254825
transform 1 0 27692 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_276
timestamp 1608254825
transform 1 0 26496 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_313
timestamp 1608254825
transform 1 0 26404 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__a211o_4  _1553_
timestamp 1608254825
transform 1 0 27324 0 1 16864
box -38 -48 1326 592
use sky130_fd_sc_hd__a21o_4  _1542_
timestamp 1608254825
transform 1 0 26588 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__o41a_4  _1538_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 28060 0 -1 16864
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_6  FILLER_27_299
timestamp 1608254825
transform 1 0 28612 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_310
timestamp 1608254825
transform 1 0 29624 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_320
timestamp 1608254825
transform 1 0 29164 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_4  _1550_
timestamp 1608254825
transform 1 0 29992 0 -1 16864
box -38 -48 1234 592
use sky130_fd_sc_hd__nor4_4  _1548_
timestamp 1608254825
transform 1 0 29256 0 1 16864
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_27_333
timestamp 1608254825
transform 1 0 31740 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_323
timestamp 1608254825
transform 1 0 30820 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_335
timestamp 1608254825
transform 1 0 31924 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_327
timestamp 1608254825
transform 1 0 31188 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_314
timestamp 1608254825
transform 1 0 32016 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2494_
timestamp 1608254825
transform 1 0 32108 0 1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__o21a_4  _1598_
timestamp 1608254825
transform 1 0 32108 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _1450_
timestamp 1608254825
transform 1 0 31372 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_364
timestamp 1608254825
transform 1 0 34592 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_356
timestamp 1608254825
transform 1 0 33856 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_365
timestamp 1608254825
transform 1 0 34684 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_357
timestamp 1608254825
transform 1 0 33948 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_349
timestamp 1608254825
transform 1 0 33212 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1448_
timestamp 1608254825
transform 1 0 33580 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_384
timestamp 1608254825
transform 1 0 36432 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_380
timestamp 1608254825
transform 1 0 36064 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_387
timestamp 1608254825
transform 1 0 36708 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_370
timestamp 1608254825
transform 1 0 35144 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_321
timestamp 1608254825
transform 1 0 34776 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2609_
timestamp 1608254825
transform 1 0 36524 0 1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  _1474_
timestamp 1608254825
transform 1 0 34776 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_4  _1455_
timestamp 1608254825
transform 1 0 35512 0 -1 16864
box -38 -48 1234 592
use sky130_fd_sc_hd__o21ai_4  _1441_
timestamp 1608254825
transform 1 0 34868 0 1 16864
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_27_404
timestamp 1608254825
transform 1 0 38272 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_411
timestamp 1608254825
transform 1 0 38916 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_26_395
timestamp 1608254825
transform 1 0 37444 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_315
timestamp 1608254825
transform 1 0 37628 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_4  _1452_
timestamp 1608254825
transform 1 0 37720 0 -1 16864
box -38 -48 1234 592
use sky130_fd_sc_hd__buf_2  _1439_
timestamp 1608254825
transform 1 0 38640 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_412
timestamp 1608254825
transform 1 0 39008 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_417
timestamp 1608254825
transform 1 0 39468 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1608254825
transform -1 0 39836 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1608254825
transform -1 0 39836 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_28_3
timestamp 1608254825
transform 1 0 1380 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1608254825
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _2640_
timestamp 1608254825
transform 1 0 1472 0 -1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_28_35
timestamp 1608254825
transform 1 0 4324 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_23
timestamp 1608254825
transform 1 0 3220 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_322
timestamp 1608254825
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1287_
timestamp 1608254825
transform 1 0 4048 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__nand4_4  _1266_
timestamp 1608254825
transform 1 0 4692 0 -1 17952
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_28_56
timestamp 1608254825
transform 1 0 6256 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__nand4_4  _1250_
timestamp 1608254825
transform 1 0 6624 0 -1 17952
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_8  FILLER_28_84
timestamp 1608254825
transform 1 0 8832 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_28_77
timestamp 1608254825
transform 1 0 8188 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1249_
timestamp 1608254825
transform 1 0 8556 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_107
timestamp 1608254825
transform 1 0 10948 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_96
timestamp 1608254825
transform 1 0 9936 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_323
timestamp 1608254825
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2558_
timestamp 1608254825
transform 1 0 11316 0 -1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__and2_4  _1884_
timestamp 1608254825
transform 1 0 10304 0 -1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1267_
timestamp 1608254825
transform 1 0 9660 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_130
timestamp 1608254825
transform 1 0 13064 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_4  _1642_
timestamp 1608254825
transform 1 0 13432 0 -1 17952
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_6  FILLER_28_147
timestamp 1608254825
transform 1 0 14628 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_324
timestamp 1608254825
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2557_
timestamp 1608254825
transform 1 0 15272 0 -1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_28_173
timestamp 1608254825
transform 1 0 17020 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__and2_4  _1871_
timestamp 1608254825
transform 1 0 17572 0 -1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_28_197
timestamp 1608254825
transform 1 0 19228 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_186
timestamp 1608254825
transform 1 0 18216 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__and2_4  _1881_
timestamp 1608254825
transform 1 0 19596 0 -1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _1879_
timestamp 1608254825
transform 1 0 18584 0 -1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_28_219
timestamp 1608254825
transform 1 0 21252 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_215
timestamp 1608254825
transform 1 0 20884 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_208
timestamp 1608254825
transform 1 0 20240 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_325
timestamp 1608254825
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__a41o_4  _2279_
timestamp 1608254825
transform 1 0 21344 0 -1 17952
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_2  FILLER_28_245
timestamp 1608254825
transform 1 0 23644 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_237
timestamp 1608254825
transform 1 0 22908 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__a41oi_4  _2115_
timestamp 1608254825
transform 1 0 23828 0 -1 17952
box -38 -48 2062 592
use sky130_fd_sc_hd__decap_6  FILLER_28_269
timestamp 1608254825
transform 1 0 25852 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_326
timestamp 1608254825
transform 1 0 26404 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__a32oi_4  _1563_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 26496 0 -1 17952
box -38 -48 2062 592
use sky130_fd_sc_hd__decap_8  FILLER_28_315
timestamp 1608254825
transform 1 0 30084 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_28_298
timestamp 1608254825
transform 1 0 28520 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_4  _1544_
timestamp 1608254825
transform 1 0 28888 0 -1 17952
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_28_332
timestamp 1608254825
transform 1 0 31648 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_327
timestamp 1608254825
transform 1 0 32016 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _1983_
timestamp 1608254825
transform 1 0 32108 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_4  _1526_
timestamp 1608254825
transform 1 0 30820 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_28_360
timestamp 1608254825
transform 1 0 34224 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_356
timestamp 1608254825
transform 1 0 33856 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_346
timestamp 1608254825
transform 1 0 32936 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__nand4_4  _1440_
timestamp 1608254825
transform 1 0 34316 0 -1 17952
box -38 -48 1602 592
use sky130_fd_sc_hd__buf_2  _1422_
timestamp 1608254825
transform 1 0 33488 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_378
timestamp 1608254825
transform 1 0 35880 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_4  _1449_
timestamp 1608254825
transform 1 0 36248 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_28_411
timestamp 1608254825
transform 1 0 38916 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_28_391
timestamp 1608254825
transform 1 0 37076 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_328
timestamp 1608254825
transform 1 0 37628 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_4  _1453_
timestamp 1608254825
transform 1 0 37720 0 -1 17952
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_1  FILLER_28_417
timestamp 1608254825
transform 1 0 39468 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1608254825
transform -1 0 39836 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_29_15
timestamp 1608254825
transform 1 0 2484 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_3
timestamp 1608254825
transform 1 0 1380 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1608254825
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__nor4_4  _1261_
timestamp 1608254825
transform 1 0 2760 0 1 17952
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_29_35
timestamp 1608254825
transform 1 0 4324 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_4  _1288_
timestamp 1608254825
transform 1 0 4692 0 1 17952
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_2  FILLER_29_59
timestamp 1608254825
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_52
timestamp 1608254825
transform 1 0 5888 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_3_0_m1_clk_local
timestamp 1608254825
transform 1 0 6256 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_329
timestamp 1608254825
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_4  _1252_
timestamp 1608254825
transform 1 0 6808 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_29_88
timestamp 1608254825
transform 1 0 9200 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_84
timestamp 1608254825
transform 1 0 8832 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_71
timestamp 1608254825
transform 1 0 7636 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2564_
timestamp 1608254825
transform 1 0 9292 0 1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__nand2_4  _1268_
timestamp 1608254825
transform 1 0 8004 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_29_108
timestamp 1608254825
transform 1 0 11040 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_5_0_addressalyzerBlock.SPI_CLK
timestamp 1608254825
transform 1 0 11408 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_128
timestamp 1608254825
transform 1 0 12880 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_123
timestamp 1608254825
transform 1 0 12420 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_118
timestamp 1608254825
transform 1 0 11960 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_330
timestamp 1608254825
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _2117_
timestamp 1608254825
transform 1 0 11684 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2089_
timestamp 1608254825
transform 1 0 12604 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__or2_4  _1641_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 13248 0 1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_29_146
timestamp 1608254825
transform 1 0 14536 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_139
timestamp 1608254825
transform 1 0 13892 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2565_
timestamp 1608254825
transform 1 0 14904 0 1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_2  _1702_
timestamp 1608254825
transform 1 0 14260 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_179
timestamp 1608254825
transform 1 0 17572 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_169
timestamp 1608254825
transform 1 0 16652 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _1880_
timestamp 1608254825
transform 1 0 17204 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_331
timestamp 1608254825
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2560_
timestamp 1608254825
transform 1 0 18032 0 1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  _1594_
timestamp 1608254825
transform 1 0 19780 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_226
timestamp 1608254825
transform 1 0 21896 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2597_
timestamp 1608254825
transform 1 0 20148 0 1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_29_245
timestamp 1608254825
transform 1 0 23644 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_243
timestamp 1608254825
transform 1 0 23460 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_239
timestamp 1608254825
transform 1 0 23092 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_332
timestamp 1608254825
transform 1 0 23552 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__a41oi_4  _1587_
timestamp 1608254825
transform 1 0 23828 0 1 17952
box -38 -48 2062 592
use sky130_fd_sc_hd__nand2_4  _1561_
timestamp 1608254825
transform 1 0 22264 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_29_269
timestamp 1608254825
transform 1 0 25852 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_284
timestamp 1608254825
transform 1 0 27232 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__and3_4  _1557_
timestamp 1608254825
transform 1 0 26404 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_4  _1552_
timestamp 1608254825
transform 1 0 27600 0 1 17952
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_8  FILLER_29_319
timestamp 1608254825
transform 1 0 30452 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_29_301
timestamp 1608254825
transform 1 0 28796 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_333
timestamp 1608254825
transform 1 0 29164 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_4  _1551_
timestamp 1608254825
transform 1 0 29256 0 1 17952
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_29_339
timestamp 1608254825
transform 1 0 32292 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_332
timestamp 1608254825
transform 1 0 31648 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_327
timestamp 1608254825
transform 1 0 31188 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1451_
timestamp 1608254825
transform 1 0 31280 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1423_
timestamp 1608254825
transform 1 0 32016 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_362
timestamp 1608254825
transform 1 0 34408 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_355
timestamp 1608254825
transform 1 0 33764 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_4  _1442_
timestamp 1608254825
transform 1 0 32660 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1421_
timestamp 1608254825
transform 1 0 34132 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_29_375
timestamp 1608254825
transform 1 0 35604 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_371
timestamp 1608254825
transform 1 0 35236 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_334
timestamp 1608254825
transform 1 0 34776 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2612_
timestamp 1608254825
transform 1 0 35696 0 1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  _1488_
timestamp 1608254825
transform 1 0 34868 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_399
timestamp 1608254825
transform 1 0 37812 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_395
timestamp 1608254825
transform 1 0 37444 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_4  _1779_
timestamp 1608254825
transform 1 0 37904 0 1 17952
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_29_414
timestamp 1608254825
transform 1 0 39192 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1608254825
transform -1 0 39836 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_30_9
timestamp 1608254825
transform 1 0 1932 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_3
timestamp 1608254825
transform 1 0 1380 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1608254825
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__o41a_4  _1285_
timestamp 1608254825
transform 1 0 2024 0 -1 19040
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_30_42
timestamp 1608254825
transform 1 0 4968 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_32
timestamp 1608254825
transform 1 0 4048 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_27
timestamp 1608254825
transform 1 0 3588 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_335
timestamp 1608254825
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1225_
timestamp 1608254825
transform 1 0 4600 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_63
timestamp 1608254825
transform 1 0 6900 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__nand4_4  _1272_
timestamp 1608254825
transform 1 0 5336 0 -1 19040
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_1  FILLER_30_91
timestamp 1608254825
transform 1 0 9476 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_85
timestamp 1608254825
transform 1 0 8924 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_78
timestamp 1608254825
transform 1 0 8280 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_4  _1248_
timestamp 1608254825
transform 1 0 7452 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1224_
timestamp 1608254825
transform 1 0 8648 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_30_104
timestamp 1608254825
transform 1 0 10672 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_100
timestamp 1608254825
transform 1 0 10304 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_336
timestamp 1608254825
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2556_
timestamp 1608254825
transform 1 0 10764 0 -1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__and2_4  _1876_
timestamp 1608254825
transform 1 0 9660 0 -1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_30_124
timestamp 1608254825
transform 1 0 12512 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_4  _1843_
timestamp 1608254825
transform 1 0 12880 0 -1 19040
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_30_149
timestamp 1608254825
transform 1 0 14812 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_141
timestamp 1608254825
transform 1 0 14076 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_337
timestamp 1608254825
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _2148_
timestamp 1608254825
transform 1 0 14444 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__or2_4  _1719_
timestamp 1608254825
transform 1 0 15272 0 -1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_30_169
timestamp 1608254825
transform 1 0 16652 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_161
timestamp 1608254825
transform 1 0 15916 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _2559_
timestamp 1608254825
transform 1 0 16744 0 -1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  FILLER_30_189
timestamp 1608254825
transform 1 0 18492 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_4  _2195_
timestamp 1608254825
transform 1 0 18768 0 -1 19040
box -38 -48 1234 592
use sky130_fd_sc_hd__and2_4  _1889_
timestamp 1608254825
transform 1 0 19964 0 -1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_30_212
timestamp 1608254825
transform 1 0 20608 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_338
timestamp 1608254825
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__and4_4  _2118_
timestamp 1608254825
transform 1 0 21252 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_4  _1595_
timestamp 1608254825
transform 1 0 22080 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _1427_
timestamp 1608254825
transform 1 0 20884 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_4  _1586_
timestamp 1608254825
transform 1 0 23184 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_269
timestamp 1608254825
transform 1 0 25852 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_252
timestamp 1608254825
transform 1 0 24288 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_4  _1582_
timestamp 1608254825
transform 1 0 24656 0 -1 19040
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_30_293
timestamp 1608254825
transform 1 0 28060 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_280
timestamp 1608254825
transform 1 0 26864 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_339
timestamp 1608254825
transform 1 0 26404 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_4  _1556_
timestamp 1608254825
transform 1 0 27232 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _1531_
timestamp 1608254825
transform 1 0 26496 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_301
timestamp 1608254825
transform 1 0 28796 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__a41o_4  _1546_
timestamp 1608254825
transform 1 0 29532 0 -1 19040
box -38 -48 1602 592
use sky130_fd_sc_hd__buf_2  _1541_
timestamp 1608254825
transform 1 0 28428 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_334
timestamp 1608254825
transform 1 0 31832 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_326
timestamp 1608254825
transform 1 0 31096 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_340
timestamp 1608254825
transform 1 0 32016 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__nand3_4  _1446_
timestamp 1608254825
transform 1 0 32108 0 -1 19040
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_30_351
timestamp 1608254825
transform 1 0 33396 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__nand4_4  _2326_
timestamp 1608254825
transform 1 0 33764 0 -1 19040
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_30_372
timestamp 1608254825
transform 1 0 35328 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__nand4_4  _1783_
timestamp 1608254825
transform 1 0 35696 0 -1 19040
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_6  FILLER_30_411
timestamp 1608254825
transform 1 0 38916 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_398
timestamp 1608254825
transform 1 0 37720 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_393
timestamp 1608254825
transform 1 0 37260 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_341
timestamp 1608254825
transform 1 0 37628 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__a21o_4  _1778_
timestamp 1608254825
transform 1 0 37812 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_417
timestamp 1608254825
transform 1 0 39468 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1608254825
transform -1 0 39836 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_15
timestamp 1608254825
transform 1 0 2484 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_7
timestamp 1608254825
transform 1 0 1748 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_3
timestamp 1608254825
transform 1 0 1380 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1608254825
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1297_
timestamp 1608254825
transform 1 0 1472 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1257_
timestamp 1608254825
transform 1 0 2116 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__nor4_4  _1247_
timestamp 1608254825
transform 1 0 2852 0 1 19040
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_1  FILLER_31_44
timestamp 1608254825
transform 1 0 5152 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_36
timestamp 1608254825
transform 1 0 4416 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_4  _1265_
timestamp 1608254825
transform 1 0 5244 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_31_62
timestamp 1608254825
transform 1 0 6808 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_60
timestamp 1608254825
transform 1 0 6624 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_54
timestamp 1608254825
transform 1 0 6072 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_342
timestamp 1608254825
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__nand4_4  _1277_
timestamp 1608254825
transform 1 0 6992 0 1 19040
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_8  FILLER_31_81
timestamp 1608254825
transform 1 0 8556 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _2563_
timestamp 1608254825
transform 1 0 9292 0 1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_31_108
timestamp 1608254825
transform 1 0 11040 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1280_
timestamp 1608254825
transform 1 0 11408 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_123
timestamp 1608254825
transform 1 0 12420 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_115
timestamp 1608254825
transform 1 0 11684 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_4_0_addressalyzerBlock.SPI_CLK
timestamp 1608254825
transform 1 0 12052 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_343
timestamp 1608254825
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_4  _1855_
timestamp 1608254825
transform 1 0 12604 0 1 19040
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_31_138
timestamp 1608254825
transform 1 0 13800 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2551_
timestamp 1608254825
transform 1 0 14168 0 1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_31_179
timestamp 1608254825
transform 1 0 17572 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_172
timestamp 1608254825
transform 1 0 16928 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_161
timestamp 1608254825
transform 1 0 15916 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__and2_4  _1872_
timestamp 1608254825
transform 1 0 16284 0 1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1591_
timestamp 1608254825
transform 1 0 17296 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_31_188
timestamp 1608254825
transform 1 0 18400 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_344
timestamp 1608254825
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2552_
timestamp 1608254825
transform 1 0 18676 0 1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  _1886_
timestamp 1608254825
transform 1 0 18032 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_210
timestamp 1608254825
transform 1 0 20424 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_addressalyzerBlock.SPI_CLK $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 20792 0 1 19040
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_3  FILLER_31_245
timestamp 1608254825
transform 1 0 23644 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_31_241
timestamp 1608254825
transform 1 0 23276 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_345
timestamp 1608254825
transform 1 0 23552 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__a41oi_4  _2116_
timestamp 1608254825
transform 1 0 23920 0 1 19040
box -38 -48 2062 592
use sky130_fd_sc_hd__and2_4  _1890_
timestamp 1608254825
transform 1 0 22632 0 1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_31_270
timestamp 1608254825
transform 1 0 25944 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1694_
timestamp 1608254825
transform 1 0 26312 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_278
timestamp 1608254825
transform 1 0 26680 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2601_
timestamp 1608254825
transform 1 0 27048 0 1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_31_301
timestamp 1608254825
transform 1 0 28796 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_346
timestamp 1608254825
transform 1 0 29164 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2602_
timestamp 1608254825
transform 1 0 29256 0 1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_31_325
timestamp 1608254825
transform 1 0 31004 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_4  _1530_
timestamp 1608254825
transform 1 0 31372 0 1 19040
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_31_362
timestamp 1608254825
transform 1 0 34408 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_351
timestamp 1608254825
transform 1 0 33396 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_343
timestamp 1608254825
transform 1 0 32660 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_4  _1528_
timestamp 1608254825
transform 1 0 33580 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_31_388
timestamp 1608254825
transform 1 0 36800 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_384
timestamp 1608254825
transform 1 0 36432 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_371
timestamp 1608254825
transform 1 0 35236 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_347
timestamp 1608254825
transform 1 0 34776 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _1679_
timestamp 1608254825
transform 1 0 35604 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _1184_
timestamp 1608254825
transform 1 0 34868 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_408
timestamp 1608254825
transform 1 0 38640 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _2595_
timestamp 1608254825
transform 1 0 36892 0 1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_31_416
timestamp 1608254825
transform 1 0 39376 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1608254825
transform -1 0 39836 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_32_22
timestamp 1608254825
transform 1 0 3128 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1608254825
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _2638_
timestamp 1608254825
transform 1 0 1380 0 -1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_32_35
timestamp 1608254825
transform 1 0 4324 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_30
timestamp 1608254825
transform 1 0 3864 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_348
timestamp 1608254825
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__o41ai_4  _1281_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 4692 0 -1 20128
box -38 -48 2062 592
use sky130_fd_sc_hd__inv_2  _1256_
timestamp 1608254825
transform 1 0 4048 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_32_61
timestamp 1608254825
transform 1 0 6716 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_32_88
timestamp 1608254825
transform 1 0 9200 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2642_
timestamp 1608254825
transform 1 0 7452 0 -1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_32_102
timestamp 1608254825
transform 1 0 10488 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_96
timestamp 1608254825
transform 1 0 9936 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_349
timestamp 1608254825
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2555_
timestamp 1608254825
transform 1 0 10580 0 -1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_2  _1273_
timestamp 1608254825
transform 1 0 9660 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_122
timestamp 1608254825
transform 1 0 12328 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_4  _1756_
timestamp 1608254825
transform 1 0 12696 0 -1 20128
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_32_149
timestamp 1608254825
transform 1 0 14812 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_139
timestamp 1608254825
transform 1 0 13892 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_350
timestamp 1608254825
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _1854_
timestamp 1608254825
transform 1 0 15272 0 -1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _1640_
timestamp 1608254825
transform 1 0 14444 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_161
timestamp 1608254825
transform 1 0 15916 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__a2bb2oi_4  _2206_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 16468 0 -1 20128
box -38 -48 1970 592
use sky130_fd_sc_hd__fill_1  FILLER_32_192
timestamp 1608254825
transform 1 0 18768 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_188
timestamp 1608254825
transform 1 0 18400 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__nand4_4  _1613_
timestamp 1608254825
transform 1 0 18860 0 -1 20128
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_32_210
timestamp 1608254825
transform 1 0 20424 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_351
timestamp 1608254825
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2598_
timestamp 1608254825
transform 1 0 20884 0 -1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_32_242
timestamp 1608254825
transform 1 0 23368 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_234
timestamp 1608254825
transform 1 0 22632 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__a41oi_4  _1596_
timestamp 1608254825
transform 1 0 23920 0 -1 20128
box -38 -48 2062 592
use sky130_fd_sc_hd__buf_2  _1560_
timestamp 1608254825
transform 1 0 23000 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_274
timestamp 1608254825
transform 1 0 26312 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_270
timestamp 1608254825
transform 1 0 25944 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_291
timestamp 1608254825
transform 1 0 27876 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_283
timestamp 1608254825
transform 1 0 27140 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_352
timestamp 1608254825
transform 1 0 26404 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _1564_
timestamp 1608254825
transform 1 0 26496 0 -1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _1500_
timestamp 1608254825
transform 1 0 27508 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_314
timestamp 1608254825
transform 1 0 29992 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_32_307
timestamp 1608254825
transform 1 0 29348 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_297
timestamp 1608254825
transform 1 0 28428 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _1608_
timestamp 1608254825
transform 1 0 28520 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1424_
timestamp 1608254825
transform 1 0 29716 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_32_337
timestamp 1608254825
transform 1 0 32108 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_335
timestamp 1608254825
transform 1 0 31924 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_327
timestamp 1608254825
transform 1 0 31188 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_322
timestamp 1608254825
transform 1 0 30728 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_353
timestamp 1608254825
transform 1 0 32016 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1545_
timestamp 1608254825
transform 1 0 30820 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_360
timestamp 1608254825
transform 1 0 34224 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__a41o_4  _1576_
timestamp 1608254825
transform 1 0 34592 0 -1 20128
box -38 -48 1602 592
use sky130_fd_sc_hd__nand4_4  _1445_
timestamp 1608254825
transform 1 0 32660 0 -1 20128
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_8  FILLER_32_381
timestamp 1608254825
transform 1 0 36156 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_32_411
timestamp 1608254825
transform 1 0 38916 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_398
timestamp 1608254825
transform 1 0 37720 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_393
timestamp 1608254825
transform 1 0 37260 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_354
timestamp 1608254825
transform 1 0 37628 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _2360_
timestamp 1608254825
transform 1 0 36892 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_4  _1780_
timestamp 1608254825
transform 1 0 38088 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_32_417
timestamp 1608254825
transform 1 0 39468 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1608254825
transform -1 0 39836 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_34_22
timestamp 1608254825
transform 1 0 3128 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_33_11
timestamp 1608254825
transform 1 0 2116 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_7
timestamp 1608254825
transform 1 0 1748 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_3
timestamp 1608254825
transform 1 0 1380 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1608254825
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1608254825
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _2637_
timestamp 1608254825
transform 1 0 1380 0 -1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_2  _1293_
timestamp 1608254825
transform 1 0 1840 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_4  _1227_
timestamp 1608254825
transform 1 0 2484 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_34_30
timestamp 1608254825
transform 1 0 3864 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_41
timestamp 1608254825
transform 1 0 4876 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_24
timestamp 1608254825
transform 1 0 3312 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_361
timestamp 1608254825
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_4  _1294_
timestamp 1608254825
transform 1 0 3680 0 1 20128
box -38 -48 1234 592
use sky130_fd_sc_hd__nand3_4  _1292_
timestamp 1608254825
transform 1 0 4048 0 -1 21216
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_34_67
timestamp 1608254825
transform 1 0 7268 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_46
timestamp 1608254825
transform 1 0 5336 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_57
timestamp 1608254825
transform 1 0 6348 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_47
timestamp 1608254825
transform 1 0 5428 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_355
timestamp 1608254825
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2641_
timestamp 1608254825
transform 1 0 6808 0 1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__and3_4  _1282_
timestamp 1608254825
transform 1 0 5520 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__nand4_4  _1260_
timestamp 1608254825
transform 1 0 5704 0 -1 21216
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_1  FILLER_34_91
timestamp 1608254825
transform 1 0 9476 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_87
timestamp 1608254825
transform 1 0 9108 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_80
timestamp 1608254825
transform 1 0 8464 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_81
timestamp 1608254825
transform 1 0 8556 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1279_
timestamp 1608254825
transform 1 0 8832 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_4  _1278_
timestamp 1608254825
transform 1 0 7636 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_4  _1276_
timestamp 1608254825
transform 1 0 8924 0 1 20128
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_34_112
timestamp 1608254825
transform 1 0 11408 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_98
timestamp 1608254825
transform 1 0 10120 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_362
timestamp 1608254825
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2631_
timestamp 1608254825
transform 1 0 9660 0 -1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__o21a_4  _1754_
timestamp 1608254825
transform 1 0 10856 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_120
timestamp 1608254825
transform 1 0 12144 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_136
timestamp 1608254825
transform 1 0 13616 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_33_118
timestamp 1608254825
transform 1 0 11960 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_356
timestamp 1608254825
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2oi_4  _2227_
timestamp 1608254825
transform 1 0 12512 0 -1 21216
box -38 -48 1970 592
use sky130_fd_sc_hd__o21ai_4  _1755_
timestamp 1608254825
transform 1 0 12420 0 1 20128
box -38 -48 1234 592
use sky130_fd_sc_hd__buf_2  _1328_
timestamp 1608254825
transform 1 0 11776 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_154
timestamp 1608254825
transform 1 0 15272 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_34_145
timestamp 1608254825
transform 1 0 14444 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_33_158
timestamp 1608254825
transform 1 0 15640 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_144
timestamp 1608254825
transform 1 0 14352 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_363
timestamp 1608254825
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_4  _2217_
timestamp 1608254825
transform 1 0 14444 0 1 20128
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_8  FILLER_34_181
timestamp 1608254825
transform 1 0 17756 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_162
timestamp 1608254825
transform 1 0 16008 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_6_0_addressalyzerBlock.SPI_CLK
timestamp 1608254825
transform 1 0 16100 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_4  _2207_
timestamp 1608254825
transform 1 0 16376 0 1 20128
box -38 -48 1234 592
use sky130_fd_sc_hd__a2bb2oi_4  _2184_
timestamp 1608254825
transform 1 0 15824 0 -1 21216
box -38 -48 1970 592
use sky130_fd_sc_hd__buf_2  _1614_
timestamp 1608254825
transform 1 0 17572 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_193
timestamp 1608254825
transform 1 0 18860 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_184
timestamp 1608254825
transform 1 0 18032 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_m1_clk_local
timestamp 1608254825
transform 1 0 18400 0 1 20128
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_357
timestamp 1608254825
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1650_
timestamp 1608254825
transform 1 0 18492 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__and4_4  _1643_
timestamp 1608254825
transform 1 0 19228 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_34_215
timestamp 1608254825
transform 1 0 20884 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_34_206
timestamp 1608254825
transform 1 0 20056 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_33_208
timestamp 1608254825
transform 1 0 20240 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_364
timestamp 1608254825
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _1592_
timestamp 1608254825
transform 1 0 20792 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_34_221
timestamp 1608254825
transform 1 0 21436 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_223
timestamp 1608254825
transform 1 0 21620 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_4  _1590_
timestamp 1608254825
transform 1 0 21804 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _1426_
timestamp 1608254825
transform 1 0 21068 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_4  _1669_
timestamp 1608254825
transform 1 0 21988 0 1 20128
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_34_247
timestamp 1608254825
transform 1 0 23828 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_234
timestamp 1608254825
transform 1 0 22632 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_249
timestamp 1608254825
transform 1 0 24012 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_240
timestamp 1608254825
transform 1 0 23184 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_358
timestamp 1608254825
transform 1 0 23552 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__and4_4  _1667_
timestamp 1608254825
transform 1 0 24196 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_4  _1606_
timestamp 1608254825
transform 1 0 23000 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _1597_
timestamp 1608254825
transform 1 0 23644 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_274
timestamp 1608254825
transform 1 0 26312 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_34_268
timestamp 1608254825
transform 1 0 25760 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_260
timestamp 1608254825
transform 1 0 25024 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_266
timestamp 1608254825
transform 1 0 25576 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2594_
timestamp 1608254825
transform 1 0 25944 0 1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__o21ai_4  _1593_
timestamp 1608254825
transform 1 0 24380 0 1 20128
box -38 -48 1234 592
use sky130_fd_sc_hd__buf_2  _1583_
timestamp 1608254825
transform 1 0 25392 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_285
timestamp 1608254825
transform 1 0 27324 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_34_279
timestamp 1608254825
transform 1 0 26772 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_33_289
timestamp 1608254825
transform 1 0 27692 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_addressalyzerBlock.SPI_CLK
timestamp 1608254825
transform 1 0 28244 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_365
timestamp 1608254825
transform 1 0 26404 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1692_
timestamp 1608254825
transform 1 0 27416 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  _1589_
timestamp 1608254825
transform 1 0 26496 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_302
timestamp 1608254825
transform 1 0 28888 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_306
timestamp 1608254825
transform 1 0 29256 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_301
timestamp 1608254825
transform 1 0 28796 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_359
timestamp 1608254825
transform 1 0 29164 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1467_
timestamp 1608254825
transform 1 0 28520 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_319
timestamp 1608254825
transform 1 0 30452 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_314
timestamp 1608254825
transform 1 0 29992 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_310
timestamp 1608254825
transform 1 0 29624 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1443_
timestamp 1608254825
transform 1 0 29716 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _2389_
timestamp 1608254825
transform 1 0 30360 0 1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__a21oi_4  _1699_
timestamp 1608254825
transform 1 0 29256 0 -1 21216
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_34_332
timestamp 1608254825
transform 1 0 31648 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_337
timestamp 1608254825
transform 1 0 32108 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_366
timestamp 1608254825
transform 1 0 32016 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__nand4_4  _2335_
timestamp 1608254825
transform 1 0 32108 0 -1 21216
box -38 -48 1602 592
use sky130_fd_sc_hd__nand2_4  _2333_
timestamp 1608254825
transform 1 0 30820 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _1577_
timestamp 1608254825
transform 1 0 32476 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_354
timestamp 1608254825
transform 1 0 33672 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_362
timestamp 1608254825
transform 1 0 34408 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_349
timestamp 1608254825
transform 1 0 33212 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_345
timestamp 1608254825
transform 1 0 32844 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_4  _1685_
timestamp 1608254825
transform 1 0 33304 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__nand3_4  _1684_
timestamp 1608254825
transform 1 0 34040 0 -1 21216
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_8  FILLER_34_372
timestamp 1608254825
transform 1 0 35328 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_367
timestamp 1608254825
transform 1 0 34868 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_360
timestamp 1608254825
transform 1 0 34776 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_4  _1686_
timestamp 1608254825
transform 1 0 36064 0 -1 21216
box -38 -48 1234 592
use sky130_fd_sc_hd__o41ai_4  _1682_
timestamp 1608254825
transform 1 0 35052 0 1 20128
box -38 -48 2062 592
use sky130_fd_sc_hd__fill_1  FILLER_34_398
timestamp 1608254825
transform 1 0 37720 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_393
timestamp 1608254825
transform 1 0 37260 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_391
timestamp 1608254825
transform 1 0 37076 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_367
timestamp 1608254825
transform 1 0 37628 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2589_
timestamp 1608254825
transform 1 0 37444 0 1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__a21oi_4  _1782_
timestamp 1608254825
transform 1 0 37812 0 -1 21216
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_6  FILLER_34_412
timestamp 1608254825
transform 1 0 39008 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_414
timestamp 1608254825
transform 1 0 39192 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1608254825
transform -1 0 39836 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1608254825
transform -1 0 39836 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_9
timestamp 1608254825
transform 1 0 1932 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_35_3
timestamp 1608254825
transform 1 0 1380 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1608254825
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__nand4_4  _1295_
timestamp 1608254825
transform 1 0 2300 0 1 21216
box -38 -48 1602 592
use sky130_fd_sc_hd__inv_2  _1259_
timestamp 1608254825
transform 1 0 1656 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_35_38
timestamp 1608254825
transform 1 0 4600 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_30
timestamp 1608254825
transform 1 0 3864 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__nand3_4  _1301_
timestamp 1608254825
transform 1 0 4692 0 1 21216
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_3  FILLER_35_62
timestamp 1608254825
transform 1 0 6808 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_35_53
timestamp 1608254825
transform 1 0 5980 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_368
timestamp 1608254825
transform 1 0 6716 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1339_
timestamp 1608254825
transform 1 0 7084 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_83
timestamp 1608254825
transform 1 0 8740 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_77
timestamp 1608254825
transform 1 0 8188 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_69
timestamp 1608254825
transform 1 0 7452 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__a41oi_4  _1340_
timestamp 1608254825
transform 1 0 8832 0 1 21216
box -38 -48 2062 592
use sky130_fd_sc_hd__buf_2  _1303_
timestamp 1608254825
transform 1 0 7820 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_106
timestamp 1608254825
transform 1 0 10856 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__and2_4  _1885_
timestamp 1608254825
transform 1 0 11224 0 1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_35_132
timestamp 1608254825
transform 1 0 13248 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_121
timestamp 1608254825
transform 1 0 12236 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_117
timestamp 1608254825
transform 1 0 11868 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_addressalyzerBlock.SPI_CLK
timestamp 1608254825
transform 1 0 13616 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_369
timestamp 1608254825
transform 1 0 12328 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__and3_4  _1652_
timestamp 1608254825
transform 1 0 12420 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_35_155
timestamp 1608254825
transform 1 0 15364 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_35_139
timestamp 1608254825
transform 1 0 13892 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_4  _2185_
timestamp 1608254825
transform 1 0 15732 0 1 21216
box -38 -48 1234 592
use sky130_fd_sc_hd__a21oi_4  _1720_
timestamp 1608254825
transform 1 0 14168 0 1 21216
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_35_179
timestamp 1608254825
transform 1 0 17572 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_172
timestamp 1608254825
transform 1 0 16928 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2246_
timestamp 1608254825
transform 1 0 17296 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_202
timestamp 1608254825
transform 1 0 19688 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_192
timestamp 1608254825
transform 1 0 18768 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_188
timestamp 1608254825
transform 1 0 18400 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_370
timestamp 1608254825
transform 1 0 17940 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1644_
timestamp 1608254825
transform 1 0 18032 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__and4_4  _1609_
timestamp 1608254825
transform 1 0 18860 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_35_215
timestamp 1608254825
transform 1 0 20884 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_4  _1664_
timestamp 1608254825
transform 1 0 21252 0 1 21216
box -38 -48 1326 592
use sky130_fd_sc_hd__nand2_4  _1647_
timestamp 1608254825
transform 1 0 20056 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_35_240
timestamp 1608254825
transform 1 0 23184 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_233
timestamp 1608254825
transform 1 0 22540 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_371
timestamp 1608254825
transform 1 0 23552 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2599_
timestamp 1608254825
transform 1 0 23644 0 1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_2  _1558_
timestamp 1608254825
transform 1 0 22908 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_264
timestamp 1608254825
transform 1 0 25392 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_4  _1573_
timestamp 1608254825
transform 1 0 25760 0 1 21216
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_1  FILLER_35_287
timestamp 1608254825
transform 1 0 27508 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_281
timestamp 1608254825
transform 1 0 26956 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_4  _1693_
timestamp 1608254825
transform 1 0 27600 0 1 21216
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_35_301
timestamp 1608254825
transform 1 0 28796 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_372
timestamp 1608254825
transform 1 0 29164 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__nand4_4  _1698_
timestamp 1608254825
transform 1 0 29256 0 1 21216
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_35_340
timestamp 1608254825
transform 1 0 32384 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_323
timestamp 1608254825
transform 1 0 30820 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_4  _2334_
timestamp 1608254825
transform 1 0 31188 0 1 21216
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_1  FILLER_35_365
timestamp 1608254825
transform 1 0 34684 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_361
timestamp 1608254825
transform 1 0 34316 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_353
timestamp 1608254825
transform 1 0 33580 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_4  _2331_
timestamp 1608254825
transform 1 0 32752 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _1221_
timestamp 1608254825
transform 1 0 33948 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_386
timestamp 1608254825
transform 1 0 36616 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_379
timestamp 1608254825
transform 1 0 35972 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_373
timestamp 1608254825
transform 1 0 34776 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_4  _1681_
timestamp 1608254825
transform 1 0 34868 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1444_
timestamp 1608254825
transform 1 0 36340 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_35_392
timestamp 1608254825
transform 1 0 37168 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2588_
timestamp 1608254825
transform 1 0 37260 0 1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_35_412
timestamp 1608254825
transform 1 0 39008 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1608254825
transform -1 0 39836 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_14
timestamp 1608254825
transform 1 0 2392 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_7
timestamp 1608254825
transform 1 0 1748 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_3
timestamp 1608254825
transform 1 0 1380 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1608254825
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1302_
timestamp 1608254825
transform 1 0 1472 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1291_
timestamp 1608254825
transform 1 0 2116 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_4  _1226_
timestamp 1608254825
transform 1 0 2760 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_36_41
timestamp 1608254825
transform 1 0 4876 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_27
timestamp 1608254825
transform 1 0 3588 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_374
timestamp 1608254825
transform 1 0 3956 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_4  _1300_
timestamp 1608254825
transform 1 0 5244 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  _1296_
timestamp 1608254825
transform 1 0 4048 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_36_54
timestamp 1608254825
transform 1 0 6072 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__nand4_4  _1246_
timestamp 1608254825
transform 1 0 6440 0 -1 22304
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_36_88
timestamp 1608254825
transform 1 0 9200 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_75
timestamp 1608254825
transform 1 0 8004 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__and4_4  _1338_
timestamp 1608254825
transform 1 0 8372 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_36_105
timestamp 1608254825
transform 1 0 10764 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_375
timestamp 1608254825
transform 1 0 9568 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_4  _1341_
timestamp 1608254825
transform 1 0 9660 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__and4_4  _1330_
timestamp 1608254825
transform 1 0 11132 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_36_126
timestamp 1608254825
transform 1 0 12696 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_118
timestamp 1608254825
transform 1 0 11960 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_4  _1653_
timestamp 1608254825
transform 1 0 13064 0 -1 22304
box -38 -48 1234 592
use sky130_fd_sc_hd__buf_2  _1334_
timestamp 1608254825
transform 1 0 12328 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_157
timestamp 1608254825
transform 1 0 15548 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_36_150
timestamp 1608254825
transform 1 0 14904 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_143
timestamp 1608254825
transform 1 0 14260 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_addressalyzerBlock.SPI_CLK
timestamp 1608254825
transform 1 0 14628 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_376
timestamp 1608254825
transform 1 0 15180 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _2290_
timestamp 1608254825
transform 1 0 15272 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_182
timestamp 1608254825
transform 1 0 17848 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2oi_4  _2161_
timestamp 1608254825
transform 1 0 15916 0 -1 22304
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_4  FILLER_36_203
timestamp 1608254825
transform 1 0 19780 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_190
timestamp 1608254825
transform 1 0 18584 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1651_
timestamp 1608254825
transform 1 0 18216 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_4  _1649_
timestamp 1608254825
transform 1 0 18952 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_36_227
timestamp 1608254825
transform 1 0 21988 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_219
timestamp 1608254825
transform 1 0 21252 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_210
timestamp 1608254825
transform 1 0 20424 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_377
timestamp 1608254825
transform 1 0 20792 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1648_
timestamp 1608254825
transform 1 0 20148 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1579_
timestamp 1608254825
transform 1 0 20884 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1220_
timestamp 1608254825
transform 1 0 21620 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_248
timestamp 1608254825
transform 1 0 23920 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__nand4_4  _1428_
timestamp 1608254825
transform 1 0 22356 0 -1 22304
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_36_271
timestamp 1608254825
transform 1 0 26036 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_256
timestamp 1608254825
transform 1 0 24656 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__o21ai_4  _1572_
timestamp 1608254825
transform 1 0 24840 0 -1 22304
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_6  FILLER_36_280
timestamp 1608254825
transform 1 0 26864 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_378
timestamp 1608254825
transform 1 0 26404 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__nor3_4  _1688_
timestamp 1608254825
transform 1 0 27416 0 -1 22304
box -38 -48 1234 592
use sky130_fd_sc_hd__buf_2  _1425_
timestamp 1608254825
transform 1 0 26496 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_306
timestamp 1608254825
transform 1 0 29256 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_299
timestamp 1608254825
transform 1 0 28612 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2393_
timestamp 1608254825
transform 1 0 29624 0 -1 22304
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_2  _1575_
timestamp 1608254825
transform 1 0 28980 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_36_335
timestamp 1608254825
transform 1 0 31924 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_329
timestamp 1608254825
transform 1 0 31372 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_379
timestamp 1608254825
transform 1 0 32016 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2390_
timestamp 1608254825
transform 1 0 32108 0 -1 22304
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_36_362
timestamp 1608254825
transform 1 0 34408 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_356
timestamp 1608254825
transform 1 0 33856 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__o41ai_4  _2327_
timestamp 1608254825
transform 1 0 34500 0 -1 22304
box -38 -48 2062 592
use sky130_fd_sc_hd__decap_4  FILLER_36_385
timestamp 1608254825
transform 1 0 36524 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_411
timestamp 1608254825
transform 1 0 38916 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_36_393
timestamp 1608254825
transform 1 0 37260 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_380
timestamp 1608254825
transform 1 0 37628 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_4  _1785_
timestamp 1608254825
transform 1 0 37720 0 -1 22304
box -38 -48 1234 592
use sky130_fd_sc_hd__buf_2  _1454_
timestamp 1608254825
transform 1 0 36892 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_417
timestamp 1608254825
transform 1 0 39468 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1608254825
transform -1 0 39836 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_17
timestamp 1608254825
transform 1 0 2668 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_9
timestamp 1608254825
transform 1 0 1932 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_37_3
timestamp 1608254825
transform 1 0 1380 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1608254825
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1314_
timestamp 1608254825
transform 1 0 1656 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_4  _1308_
timestamp 1608254825
transform 1 0 3036 0 1 22304
box -38 -48 1326 592
use sky130_fd_sc_hd__buf_2  _1304_
timestamp 1608254825
transform 1 0 2300 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_42
timestamp 1608254825
transform 1 0 4968 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_35
timestamp 1608254825
transform 1 0 4324 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1299_
timestamp 1608254825
transform 1 0 4692 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_57
timestamp 1608254825
transform 1 0 6348 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_49
timestamp 1608254825
transform 1 0 5612 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_381
timestamp 1608254825
transform 1 0 6716 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1311_
timestamp 1608254825
transform 1 0 5980 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__and4_4  _1305_
timestamp 1608254825
transform 1 0 6808 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1245_
timestamp 1608254825
transform 1 0 5336 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_37_71
timestamp 1608254825
transform 1 0 7636 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  _2630_
timestamp 1608254825
transform 1 0 8188 0 1 22304
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  FILLER_37_104
timestamp 1608254825
transform 1 0 10672 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_37_96
timestamp 1608254825
transform 1 0 9936 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__and4_4  _1242_
timestamp 1608254825
transform 1 0 10948 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_37_126
timestamp 1608254825
transform 1 0 12696 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_116
timestamp 1608254825
transform 1 0 11776 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_382
timestamp 1608254825
transform 1 0 12328 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_4  _1857_
timestamp 1608254825
transform 1 0 13064 0 1 22304
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _1337_
timestamp 1608254825
transform 1 0 12420 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_143
timestamp 1608254825
transform 1 0 14260 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_4  _2228_
timestamp 1608254825
transform 1 0 14628 0 1 22304
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_1  FILLER_37_182
timestamp 1608254825
transform 1 0 17848 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_178
timestamp 1608254825
transform 1 0 17480 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_164
timestamp 1608254825
transform 1 0 16192 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_160
timestamp 1608254825
transform 1 0 15824 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_4  _2162_
timestamp 1608254825
transform 1 0 16284 0 1 22304
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_6  FILLER_37_197
timestamp 1608254825
transform 1 0 19228 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_383
timestamp 1608254825
transform 1 0 17940 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_4  _2149_
timestamp 1608254825
transform 1 0 18032 0 1 22304
box -38 -48 1234 592
use sky130_fd_sc_hd__buf_2  _1605_
timestamp 1608254825
transform 1 0 19780 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_215
timestamp 1608254825
transform 1 0 20884 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_207
timestamp 1608254825
transform 1 0 20148 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1584_
timestamp 1608254825
transform 1 0 20516 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_4  _1567_
timestamp 1608254825
transform 1 0 21252 0 1 22304
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_37_240
timestamp 1608254825
transform 1 0 23184 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_233
timestamp 1608254825
transform 1 0 22540 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_384
timestamp 1608254825
transform 1 0 23552 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _1559_
timestamp 1608254825
transform 1 0 23644 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1189_
timestamp 1608254825
transform 1 0 22908 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_37_260
timestamp 1608254825
transform 1 0 25024 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_37_254
timestamp 1608254825
transform 1 0 24472 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  _2600_
timestamp 1608254825
transform 1 0 25116 0 1 22304
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_37_280
timestamp 1608254825
transform 1 0 26864 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__nor3_4  _1690_
timestamp 1608254825
transform 1 0 27600 0 1 22304
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_2  FILLER_37_306
timestamp 1608254825
transform 1 0 29256 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_301
timestamp 1608254825
transform 1 0 28796 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_385
timestamp 1608254825
transform 1 0 29164 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__nor3_4  _2340_
timestamp 1608254825
transform 1 0 29440 0 1 22304
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_2  FILLER_37_339
timestamp 1608254825
transform 1 0 32292 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_331
timestamp 1608254825
transform 1 0 31556 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_37_321
timestamp 1608254825
transform 1 0 30636 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__a22oi_4  _2330_
timestamp 1608254825
transform 1 0 32476 0 1 22304
box -38 -48 1602 592
use sky130_fd_sc_hd__buf_2  _1585_
timestamp 1608254825
transform 1 0 31188 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_358
timestamp 1608254825
transform 1 0 34040 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_37_386
timestamp 1608254825
transform 1 0 36616 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_386
timestamp 1608254825
transform 1 0 34776 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2387_
timestamp 1608254825
transform 1 0 34868 0 1 22304
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_37_394
timestamp 1608254825
transform 1 0 37352 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2463_
timestamp 1608254825
transform 1 0 37444 0 1 22304
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_37_414
timestamp 1608254825
transform 1 0 39192 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1608254825
transform -1 0 39836 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_38_22
timestamp 1608254825
transform 1 0 3128 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1608254825
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _2635_
timestamp 1608254825
transform 1 0 1380 0 -1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_38_32
timestamp 1608254825
transform 1 0 4048 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_30
timestamp 1608254825
transform 1 0 3864 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_387
timestamp 1608254825
transform 1 0 3956 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__a41oi_4  _1312_
timestamp 1608254825
transform 1 0 4600 0 -1 23392
box -38 -48 2062 592
use sky130_fd_sc_hd__decap_4  FILLER_38_60
timestamp 1608254825
transform 1 0 6624 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_4  _1307_
timestamp 1608254825
transform 1 0 6992 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_84
timestamp 1608254825
transform 1 0 8832 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_38_76
timestamp 1608254825
transform 1 0 8096 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1243_
timestamp 1608254825
transform 1 0 8464 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_93
timestamp 1608254825
transform 1 0 9660 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_388
timestamp 1608254825
transform 1 0 9568 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__nand4_4  _1335_
timestamp 1608254825
transform 1 0 10212 0 -1 23392
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_38_132
timestamp 1608254825
transform 1 0 13248 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_116
timestamp 1608254825
transform 1 0 11776 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_4  _2208_
timestamp 1608254825
transform 1 0 12144 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__o21a_4  _2186_
timestamp 1608254825
transform 1 0 13616 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_152
timestamp 1608254825
transform 1 0 15088 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_148
timestamp 1608254825
transform 1 0 14720 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_389
timestamp 1608254825
transform 1 0 15180 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__a21o_4  _2187_
timestamp 1608254825
transform 1 0 15272 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_178
timestamp 1608254825
transform 1 0 17480 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_173
timestamp 1608254825
transform 1 0 17020 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_166
timestamp 1608254825
transform 1 0 16376 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_addressalyzerBlock.SPI_CLK
timestamp 1608254825
transform 1 0 16744 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_4  _2173_
timestamp 1608254825
transform 1 0 17848 0 -1 23392
box -38 -48 1234 592
use sky130_fd_sc_hd__buf_2  _1610_
timestamp 1608254825
transform 1 0 17112 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_195
timestamp 1608254825
transform 1 0 19044 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_4  _2189_
timestamp 1608254825
transform 1 0 19596 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_38_215
timestamp 1608254825
transform 1 0 20884 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_210
timestamp 1608254825
transform 1 0 20424 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_390
timestamp 1608254825
transform 1 0 20792 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__nor3_4  _1665_
timestamp 1608254825
transform 1 0 20976 0 -1 23392
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_38_247
timestamp 1608254825
transform 1 0 23828 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_233
timestamp 1608254825
transform 1 0 22540 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_229
timestamp 1608254825
transform 1 0 22172 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_4  _1671_
timestamp 1608254825
transform 1 0 22632 0 -1 23392
box -38 -48 1234 592
use sky130_fd_sc_hd__buf_2  _1219_
timestamp 1608254825
transform 1 0 24196 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_271
timestamp 1608254825
transform 1 0 26036 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_255
timestamp 1608254825
transform 1 0 24564 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_4  _2325_
timestamp 1608254825
transform 1 0 24932 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_288
timestamp 1608254825
transform 1 0 27600 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_391
timestamp 1608254825
transform 1 0 26404 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__nor3_4  _1728_
timestamp 1608254825
transform 1 0 28336 0 -1 23392
box -38 -48 1234 592
use sky130_fd_sc_hd__o21a_4  _1569_
timestamp 1608254825
transform 1 0 26496 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_319
timestamp 1608254825
transform 1 0 30452 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_309
timestamp 1608254825
transform 1 0 29532 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _2101_
timestamp 1608254825
transform 1 0 30084 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_335
timestamp 1608254825
transform 1 0 31924 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_327
timestamp 1608254825
transform 1 0 31188 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_392
timestamp 1608254825
transform 1 0 32016 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_4  _2336_
timestamp 1608254825
transform 1 0 32108 0 -1 23392
box -38 -48 1234 592
use sky130_fd_sc_hd__buf_2  _1566_
timestamp 1608254825
transform 1 0 30820 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_358
timestamp 1608254825
transform 1 0 34040 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_350
timestamp 1608254825
transform 1 0 33304 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__and3_4  _2338_
timestamp 1608254825
transform 1 0 34132 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_38_383
timestamp 1608254825
transform 1 0 36340 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_379
timestamp 1608254825
transform 1 0 35972 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_368
timestamp 1608254825
transform 1 0 34960 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_4  _1784_
timestamp 1608254825
transform 1 0 36432 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__or2_4  _1680_
timestamp 1608254825
transform 1 0 35328 0 -1 23392
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_38_407
timestamp 1608254825
transform 1 0 38548 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_393
timestamp 1608254825
transform 1 0 37260 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_393
timestamp 1608254825
transform 1 0 37628 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _1736_
timestamp 1608254825
transform 1 0 37720 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1678_
timestamp 1608254825
transform 1 0 38916 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_414
timestamp 1608254825
transform 1 0 39192 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1608254825
transform -1 0 39836 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_40_7
timestamp 1608254825
transform 1 0 1748 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_3
timestamp 1608254825
transform 1 0 1380 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_7
timestamp 1608254825
transform 1 0 1748 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_3
timestamp 1608254825
transform 1 0 1380 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1608254825
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1608254825
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_20
timestamp 1608254825
transform 1 0 2944 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_21
timestamp 1608254825
transform 1 0 3036 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_4  _2086_
timestamp 1608254825
transform 1 0 1840 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__o21ai_4  _1313_
timestamp 1608254825
transform 1 0 1840 0 1 23392
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_1  FILLER_40_45
timestamp 1608254825
transform 1 0 5244 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_41
timestamp 1608254825
transform 1 0 4876 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_27
timestamp 1608254825
transform 1 0 3588 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_44
timestamp 1608254825
transform 1 0 5152 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_400
timestamp 1608254825
transform 1 0 3956 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2636_
timestamp 1608254825
transform 1 0 3404 0 1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_2  _1310_
timestamp 1608254825
transform 1 0 3312 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_4  _1309_
timestamp 1608254825
transform 1 0 4048 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_40_59
timestamp 1608254825
transform 1 0 6532 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_62
timestamp 1608254825
transform 1 0 6808 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_57
timestamp 1608254825
transform 1 0 6348 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_394
timestamp 1608254825
transform 1 0 6716 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_4  _1343_
timestamp 1608254825
transform 1 0 6900 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__o21ai_4  _1326_
timestamp 1608254825
transform 1 0 5336 0 -1 24480
box -38 -48 1234 592
use sky130_fd_sc_hd__nand3_4  _1322_
timestamp 1608254825
transform 1 0 6900 0 -1 24480
box -38 -48 1326 592
use sky130_fd_sc_hd__nand2_4  _1244_
timestamp 1608254825
transform 1 0 5520 0 1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_40_91
timestamp 1608254825
transform 1 0 9476 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_40_85
timestamp 1608254825
transform 1 0 8924 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_40_77
timestamp 1608254825
transform 1 0 8188 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_75
timestamp 1608254825
transform 1 0 8004 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__a41oi_4  _1342_
timestamp 1608254825
transform 1 0 8372 0 1 23392
box -38 -48 2062 592
use sky130_fd_sc_hd__buf_2  _1321_
timestamp 1608254825
transform 1 0 8556 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_113
timestamp 1608254825
transform 1 0 11500 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_40_105
timestamp 1608254825
transform 1 0 10764 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_105
timestamp 1608254825
transform 1 0 10764 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_101
timestamp 1608254825
transform 1 0 10396 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_401
timestamp 1608254825
transform 1 0 9568 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__a21o_4  _1344_
timestamp 1608254825
transform 1 0 9660 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__o21a_4  _1331_
timestamp 1608254825
transform 1 0 10856 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _1329_
timestamp 1608254825
transform 1 0 11132 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_133
timestamp 1608254825
transform 1 0 13340 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_119
timestamp 1608254825
transform 1 0 12052 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_118
timestamp 1608254825
transform 1 0 11960 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_395
timestamp 1608254825
transform 1 0 12328 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2632_
timestamp 1608254825
transform 1 0 12420 0 1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__o21a_4  _2163_
timestamp 1608254825
transform 1 0 13708 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__o21ai_4  _1742_
timestamp 1608254825
transform 1 0 12144 0 -1 24480
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_40_157
timestamp 1608254825
transform 1 0 15548 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_149
timestamp 1608254825
transform 1 0 14812 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_150
timestamp 1608254825
transform 1 0 14904 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_142
timestamp 1608254825
transform 1 0 14168 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_402
timestamp 1608254825
transform 1 0 15180 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_4  _2188_
timestamp 1608254825
transform 1 0 15272 0 1 23392
box -38 -48 1234 592
use sky130_fd_sc_hd__buf_2  _1646_
timestamp 1608254825
transform 1 0 14536 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1645_
timestamp 1608254825
transform 1 0 15272 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_177
timestamp 1608254825
transform 1 0 17388 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_182
timestamp 1608254825
transform 1 0 17848 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_176
timestamp 1608254825
transform 1 0 17296 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_171
timestamp 1608254825
transform 1 0 16836 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_167
timestamp 1608254825
transform 1 0 16468 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_7_0_addressalyzerBlock.SPI_CLK
timestamp 1608254825
transform 1 0 15916 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_4  _2209_
timestamp 1608254825
transform 1 0 17756 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__a21oi_4  _2165_
timestamp 1608254825
transform 1 0 16192 0 -1 24480
box -38 -48 1234 592
use sky130_fd_sc_hd__buf_2  _1655_
timestamp 1608254825
transform 1 0 16928 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_205
timestamp 1608254825
transform 1 0 19964 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_201
timestamp 1608254825
transform 1 0 19596 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_193
timestamp 1608254825
transform 1 0 18860 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_197
timestamp 1608254825
transform 1 0 19228 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_396
timestamp 1608254825
transform 1 0 17940 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_4  _2210_
timestamp 1608254825
transform 1 0 18032 0 1 23392
box -38 -48 1234 592
use sky130_fd_sc_hd__nor3_4  _1654_
timestamp 1608254825
transform 1 0 19596 0 1 23392
box -38 -48 1234 592
use sky130_fd_sc_hd__buf_2  _1405_
timestamp 1608254825
transform 1 0 19228 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_226
timestamp 1608254825
transform 1 0 21896 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_215
timestamp 1608254825
transform 1 0 20884 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_210
timestamp 1608254825
transform 1 0 20424 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_214
timestamp 1608254825
transform 1 0 20792 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_403
timestamp 1608254825
transform 1 0 20792 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_4  _2211_
timestamp 1608254825
transform 1 0 21068 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_4  _2190_
timestamp 1608254825
transform 1 0 21160 0 1 23392
box -38 -48 1234 592
use sky130_fd_sc_hd__buf_2  _1659_
timestamp 1608254825
transform 1 0 20056 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_234
timestamp 1608254825
transform 1 0 22632 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_239
timestamp 1608254825
transform 1 0 23092 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_231
timestamp 1608254825
transform 1 0 22356 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1570_
timestamp 1608254825
transform 1 0 22724 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1568_
timestamp 1608254825
transform 1 0 22264 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_245
timestamp 1608254825
transform 1 0 23644 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_39_243
timestamp 1608254825
transform 1 0 23460 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_397
timestamp 1608254825
transform 1 0 23552 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _1604_
timestamp 1608254825
transform 1 0 23828 0 1 23392
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_4  _1724_
timestamp 1608254825
transform 1 0 23000 0 -1 24480
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_40_271
timestamp 1608254825
transform 1 0 26036 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_252
timestamp 1608254825
transform 1 0 24288 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_274
timestamp 1608254825
transform 1 0 26312 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_260
timestamp 1608254825
transform 1 0 25024 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_254
timestamp 1608254825
transform 1 0 24472 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_4  _1733_
timestamp 1608254825
transform 1 0 25116 0 1 23392
box -38 -48 1234 592
use sky130_fd_sc_hd__a21oi_4  _1732_
timestamp 1608254825
transform 1 0 24840 0 -1 24480
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_40_295
timestamp 1608254825
transform 1 0 28244 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_276
timestamp 1608254825
transform 1 0 26496 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_404
timestamp 1608254825
transform 1 0 26404 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2394_
timestamp 1608254825
transform 1 0 26680 0 1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__nor3_4  _1731_
timestamp 1608254825
transform 1 0 27048 0 -1 24480
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_40_313
timestamp 1608254825
transform 1 0 29900 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_317
timestamp 1608254825
transform 1 0 30268 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_310
timestamp 1608254825
transform 1 0 29624 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_297
timestamp 1608254825
transform 1 0 28428 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_398
timestamp 1608254825
transform 1 0 29164 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__a211o_4  _1730_
timestamp 1608254825
transform 1 0 28612 0 -1 24480
box -38 -48 1326 592
use sky130_fd_sc_hd__inv_2  _1574_
timestamp 1608254825
transform 1 0 29992 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1565_
timestamp 1608254825
transform 1 0 29256 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_4  _1434_
timestamp 1608254825
transform 1 0 30268 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_40_337
timestamp 1608254825
transform 1 0 32108 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_334
timestamp 1608254825
transform 1 0 31832 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_40_326
timestamp 1608254825
transform 1 0 31096 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_39_340
timestamp 1608254825
transform 1 0 32384 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_405
timestamp 1608254825
transform 1 0 32016 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2388_
timestamp 1608254825
transform 1 0 30636 0 1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__o32ai_4  _2329_
timestamp 1608254825
transform 1 0 32384 0 -1 24480
box -38 -48 2062 592
use sky130_fd_sc_hd__decap_4  FILLER_40_362
timestamp 1608254825
transform 1 0 34408 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_362
timestamp 1608254825
transform 1 0 34408 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_4  _2337_
timestamp 1608254825
transform 1 0 33120 0 1 23392
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_40_385
timestamp 1608254825
transform 1 0 36524 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_386
timestamp 1608254825
transform 1 0 36616 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_371
timestamp 1608254825
transform 1 0 35236 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_399
timestamp 1608254825
transform 1 0 34776 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2385_
timestamp 1608254825
transform 1 0 34776 0 -1 24480
box -38 -48 1786 592
use sky130_fd_sc_hd__nand2_4  _2111_
timestamp 1608254825
transform 1 0 35788 0 1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _1217_
timestamp 1608254825
transform 1 0 34868 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_411
timestamp 1608254825
transform 1 0 38916 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_396
timestamp 1608254825
transform 1 0 37536 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_392
timestamp 1608254825
transform 1 0 37168 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_409
timestamp 1608254825
transform 1 0 38732 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_406
timestamp 1608254825
transform 1 0 37628 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2462_
timestamp 1608254825
transform 1 0 36984 0 1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__nor3_4  _2100_
timestamp 1608254825
transform 1 0 37720 0 -1 24480
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _1185_
timestamp 1608254825
transform 1 0 36892 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_40_417
timestamp 1608254825
transform 1 0 39468 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_39_417
timestamp 1608254825
transform 1 0 39468 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1608254825
transform -1 0 39836 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1608254825
transform -1 0 39836 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_41_8
timestamp 1608254825
transform 1 0 1840 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_3
timestamp 1608254825
transform 1 0 1380 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1608254825
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2345_
timestamp 1608254825
transform 1 0 1564 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_4  _2085_
timestamp 1608254825
transform 1 0 2208 0 1 24480
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_1  FILLER_41_31
timestamp 1608254825
transform 1 0 3956 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_41_25
timestamp 1608254825
transform 1 0 3404 0 1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  _2633_
timestamp 1608254825
transform 1 0 4048 0 1 24480
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_41_59
timestamp 1608254825
transform 1 0 6532 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_41_51
timestamp 1608254825
transform 1 0 5796 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_407
timestamp 1608254825
transform 1 0 6716 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__a41oi_4  _1325_
timestamp 1608254825
transform 1 0 6808 0 1 24480
box -38 -48 2062 592
use sky130_fd_sc_hd__decap_4  FILLER_41_84
timestamp 1608254825
transform 1 0 8832 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_4  _1347_
timestamp 1608254825
transform 1 0 9200 0 1 24480
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_41_102
timestamp 1608254825
transform 1 0 10488 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_4  _1336_
timestamp 1608254825
transform 1 0 10856 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_41_134
timestamp 1608254825
transform 1 0 13432 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_126
timestamp 1608254825
transform 1 0 12696 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_121
timestamp 1608254825
transform 1 0 12236 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_41_115
timestamp 1608254825
transform 1 0 11684 0 1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_408
timestamp 1608254825
transform 1 0 12328 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__a21o_4  _1700_
timestamp 1608254825
transform 1 0 13524 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1348_
timestamp 1608254825
transform 1 0 12420 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_41_159
timestamp 1608254825
transform 1 0 15732 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_155
timestamp 1608254825
transform 1 0 15364 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_147
timestamp 1608254825
transform 1 0 14628 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1611_
timestamp 1608254825
transform 1 0 14996 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_179
timestamp 1608254825
transform 1 0 17572 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_172
timestamp 1608254825
transform 1 0 16928 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_4  _2164_
timestamp 1608254825
transform 1 0 15824 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _2146_
timestamp 1608254825
transform 1 0 17296 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_41_201
timestamp 1608254825
transform 1 0 19596 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_41_193
timestamp 1608254825
transform 1 0 18860 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_409
timestamp 1608254825
transform 1 0 17940 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__o41ai_4  _2172_
timestamp 1608254825
transform 1 0 19780 0 1 24480
box -38 -48 2062 592
use sky130_fd_sc_hd__and3_4  _1419_
timestamp 1608254825
transform 1 0 18032 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_41_225
timestamp 1608254825
transform 1 0 21804 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_245
timestamp 1608254825
transform 1 0 23644 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_240
timestamp 1608254825
transform 1 0 23184 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_232
timestamp 1608254825
transform 1 0 22448 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_410
timestamp 1608254825
transform 1 0 23552 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1670_
timestamp 1608254825
transform 1 0 22172 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1571_
timestamp 1608254825
transform 1 0 22816 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1190_
timestamp 1608254825
transform 1 0 24012 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_253
timestamp 1608254825
transform 1 0 24380 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _2592_
timestamp 1608254825
transform 1 0 25116 0 1 24480
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_41_280
timestamp 1608254825
transform 1 0 26864 0 1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_4  _2324_
timestamp 1608254825
transform 1 0 27416 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_319
timestamp 1608254825
transform 1 0 30452 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_304
timestamp 1608254825
transform 1 0 29072 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_41_298
timestamp 1608254825
transform 1 0 28520 0 1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_411
timestamp 1608254825
transform 1 0 29164 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__nor3_4  _1729_
timestamp 1608254825
transform 1 0 29256 0 1 24480
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_41_335
timestamp 1608254825
transform 1 0 31924 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2386_
timestamp 1608254825
transform 1 0 32292 0 1 24480
box -38 -48 1786 592
use sky130_fd_sc_hd__a21o_4  _2328_
timestamp 1608254825
transform 1 0 30820 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_358
timestamp 1608254825
transform 1 0 34040 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_41_381
timestamp 1608254825
transform 1 0 36156 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_412
timestamp 1608254825
transform 1 0 34776 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__a211o_4  _2339_
timestamp 1608254825
transform 1 0 34868 0 1 24480
box -38 -48 1326 592
use sky130_fd_sc_hd__buf_2  _1870_
timestamp 1608254825
transform 1 0 36524 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_389
timestamp 1608254825
transform 1 0 36892 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2453_
timestamp 1608254825
transform 1 0 37260 0 1 24480
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_41_412
timestamp 1608254825
transform 1 0 39008 0 1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1608254825
transform -1 0 39836 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_42_22
timestamp 1608254825
transform 1 0 3128 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1608254825
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _2472_
timestamp 1608254825
transform 1 0 1380 0 -1 25568
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_42_45
timestamp 1608254825
transform 1 0 5244 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_41
timestamp 1608254825
transform 1 0 4876 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_30
timestamp 1608254825
transform 1 0 3864 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_413
timestamp 1608254825
transform 1 0 3956 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _2087_
timestamp 1608254825
transform 1 0 4048 0 -1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_42_67
timestamp 1608254825
transform 1 0 7268 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_63
timestamp 1608254825
transform 1 0 6900 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__nand4_4  _1318_
timestamp 1608254825
transform 1 0 5336 0 -1 25568
box -38 -48 1602 592
use sky130_fd_sc_hd__and4_4  _1316_
timestamp 1608254825
transform 1 0 7360 0 -1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_42_84
timestamp 1608254825
transform 1 0 8832 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_42_77
timestamp 1608254825
transform 1 0 8188 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1241_
timestamp 1608254825
transform 1 0 8556 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_42_114
timestamp 1608254825
transform 1 0 11592 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_93
timestamp 1608254825
transform 1 0 9660 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_414
timestamp 1608254825
transform 1 0 9568 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2629_
timestamp 1608254825
transform 1 0 9844 0 -1 25568
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_42_136
timestamp 1608254825
transform 1 0 13616 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_122
timestamp 1608254825
transform 1 0 12328 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_4  _1758_
timestamp 1608254825
transform 1 0 12420 0 -1 25568
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_42_149
timestamp 1608254825
transform 1 0 14812 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_144
timestamp 1608254825
transform 1 0 14352 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_415
timestamp 1608254825
transform 1 0 15180 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_4  _2229_
timestamp 1608254825
transform 1 0 15272 0 -1 25568
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _1741_
timestamp 1608254825
transform 1 0 14536 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_42_173
timestamp 1608254825
transform 1 0 17020 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_167
timestamp 1608254825
transform 1 0 16468 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  _2613_
timestamp 1608254825
transform 1 0 17112 0 -1 25568
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_42_204
timestamp 1608254825
transform 1 0 19872 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_42_193
timestamp 1608254825
transform 1 0 18860 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__or2_4  _1411_
timestamp 1608254825
transform 1 0 19228 0 -1 25568
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_42_212
timestamp 1608254825
transform 1 0 20608 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_416
timestamp 1608254825
transform 1 0 20792 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__o41ai_4  _2194_
timestamp 1608254825
transform 1 0 20884 0 -1 25568
box -38 -48 2062 592
use sky130_fd_sc_hd__decap_8  FILLER_42_245
timestamp 1608254825
transform 1 0 23644 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_42_237
timestamp 1608254825
transform 1 0 22908 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1660_
timestamp 1608254825
transform 1 0 23276 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_271
timestamp 1608254825
transform 1 0 26036 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_264
timestamp 1608254825
transform 1 0 25392 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_253
timestamp 1608254825
transform 1 0 24380 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__nand2_4  _2235_
timestamp 1608254825
transform 1 0 24564 0 -1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1662_
timestamp 1608254825
transform 1 0 25760 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_42_289
timestamp 1608254825
transform 1 0 27692 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_417
timestamp 1608254825
transform 1 0 26404 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_4  _2237_
timestamp 1608254825
transform 1 0 26496 0 -1 25568
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_42_302
timestamp 1608254825
transform 1 0 28888 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_297
timestamp 1608254825
transform 1 0 28428 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__a211o_4  _2332_
timestamp 1608254825
transform 1 0 29256 0 -1 25568
box -38 -48 1326 592
use sky130_fd_sc_hd__inv_2  _1687_
timestamp 1608254825
transform 1 0 28612 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_42_328
timestamp 1608254825
transform 1 0 31280 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_42_320
timestamp 1608254825
transform 1 0 30544 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_418
timestamp 1608254825
transform 1 0 32016 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1781_
timestamp 1608254825
transform 1 0 30912 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_4  _1218_
timestamp 1608254825
transform 1 0 32108 0 -1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_42_362
timestamp 1608254825
transform 1 0 34408 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_354
timestamp 1608254825
transform 1 0 33672 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_42_346
timestamp 1608254825
transform 1 0 32936 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__or2_4  _2105_
timestamp 1608254825
transform 1 0 34500 0 -1 25568
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _1212_
timestamp 1608254825
transform 1 0 33304 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_370
timestamp 1608254825
transform 1 0 35144 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__nor4_4  _2102_
timestamp 1608254825
transform 1 0 35512 0 -1 25568
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_8  FILLER_42_410
timestamp 1608254825
transform 1 0 38824 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_42_398
timestamp 1608254825
transform 1 0 37720 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_42_391
timestamp 1608254825
transform 1 0 37076 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_419
timestamp 1608254825
transform 1 0 37628 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__and3_4  _2099_
timestamp 1608254825
transform 1 0 37996 0 -1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1608254825
transform -1 0 39836 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_43_15
timestamp 1608254825
transform 1 0 2484 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_3
timestamp 1608254825
transform 1 0 1380 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1608254825
transform 1 0 1104 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _2471_
timestamp 1608254825
transform 1 0 2576 0 1 25568
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_43_43
timestamp 1608254825
transform 1 0 5060 0 1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_35
timestamp 1608254825
transform 1 0 4324 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _2078_
timestamp 1608254825
transform 1 0 4692 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_43_62
timestamp 1608254825
transform 1 0 6808 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_43_60
timestamp 1608254825
transform 1 0 6624 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_43_54
timestamp 1608254825
transform 1 0 6072 0 1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_49
timestamp 1608254825
transform 1 0 5612 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_420
timestamp 1608254825
transform 1 0 6716 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1324_
timestamp 1608254825
transform 1 0 7084 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1315_
timestamp 1608254825
transform 1 0 5704 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_86
timestamp 1608254825
transform 1 0 9016 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_69
timestamp 1608254825
transform 1 0 7452 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1323_
timestamp 1608254825
transform 1 0 9384 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_4  _1258_
timestamp 1608254825
transform 1 0 7820 0 1 25568
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_8  FILLER_43_93
timestamp 1608254825
transform 1 0 9660 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__nor4_4  _1333_
timestamp 1608254825
transform 1 0 10396 0 1 25568
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_1  FILLER_43_136
timestamp 1608254825
transform 1 0 13616 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_132
timestamp 1608254825
transform 1 0 13248 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_118
timestamp 1608254825
transform 1 0 11960 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_421
timestamp 1608254825
transform 1 0 12328 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__and3_4  _1856_
timestamp 1608254825
transform 1 0 12420 0 1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_4  _1722_
timestamp 1608254825
transform 1 0 13708 0 1 25568
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_43_150
timestamp 1608254825
transform 1 0 14904 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_4  _2231_
timestamp 1608254825
transform 1 0 15272 0 1 25568
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_43_179
timestamp 1608254825
transform 1 0 17572 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_171
timestamp 1608254825
transform 1 0 16836 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_167
timestamp 1608254825
transform 1 0 16468 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__or2_4  _1418_
timestamp 1608254825
transform 1 0 16928 0 1 25568
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_43_204
timestamp 1608254825
transform 1 0 19872 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_43_184
timestamp 1608254825
transform 1 0 18032 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_422
timestamp 1608254825
transform 1 0 17940 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__nand4_4  _1232_
timestamp 1608254825
transform 1 0 18308 0 1 25568
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_6  FILLER_43_221
timestamp 1608254825
transform 1 0 21436 0 1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_4  _2233_
timestamp 1608254825
transform 1 0 21988 0 1 25568
box -38 -48 1234 592
use sky130_fd_sc_hd__o21ai_4  _2212_
timestamp 1608254825
transform 1 0 20240 0 1 25568
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_43_240
timestamp 1608254825
transform 1 0 23184 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_423
timestamp 1608254825
transform 1 0 23552 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__a21boi_4  _2232_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 23644 0 1 25568
box -38 -48 1418 592
use sky130_fd_sc_hd__fill_1  FILLER_43_274
timestamp 1608254825
transform 1 0 26312 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_43_268
timestamp 1608254825
transform 1 0 25760 0 1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_260
timestamp 1608254825
transform 1 0 25024 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1663_
timestamp 1608254825
transform 1 0 25392 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_294
timestamp 1608254825
transform 1 0 28152 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2435_
timestamp 1608254825
transform 1 0 26404 0 1 25568
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_43_306
timestamp 1608254825
transform 1 0 29256 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_301
timestamp 1608254825
transform 1 0 28796 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_424
timestamp 1608254825
transform 1 0 29164 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2392_
timestamp 1608254825
transform 1 0 29348 0 1 25568
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_2  _1689_
timestamp 1608254825
transform 1 0 28520 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_43_330
timestamp 1608254825
transform 1 0 31464 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_326
timestamp 1608254825
transform 1 0 31096 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_4  _1223_
timestamp 1608254825
transform 1 0 31556 0 1 25568
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_1  FILLER_43_365
timestamp 1608254825
transform 1 0 34684 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_357
timestamp 1608254825
transform 1 0 33948 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_43_344
timestamp 1608254825
transform 1 0 32752 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_4  _2322_
timestamp 1608254825
transform 1 0 33120 0 1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_43_386
timestamp 1608254825
transform 1 0 36616 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_425
timestamp 1608254825
transform 1 0 34776 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2459_
timestamp 1608254825
transform 1 0 34868 0 1 25568
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_43_394
timestamp 1608254825
transform 1 0 37352 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2452_
timestamp 1608254825
transform 1 0 37444 0 1 25568
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_43_414
timestamp 1608254825
transform 1 0 39192 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1608254825
transform -1 0 39836 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_44_21
timestamp 1608254825
transform 1 0 3036 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_44_3
timestamp 1608254825
transform 1 0 1380 0 -1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1608254825
transform 1 0 1104 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_4  _2083_
timestamp 1608254825
transform 1 0 1932 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_43
timestamp 1608254825
transform 1 0 5060 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_36
timestamp 1608254825
transform 1 0 4416 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_29
timestamp 1608254825
transform 1 0 3772 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_426
timestamp 1608254825
transform 1 0 3956 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1320_
timestamp 1608254825
transform 1 0 4784 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1284_
timestamp 1608254825
transform 1 0 4048 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_66
timestamp 1608254825
transform 1 0 7176 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _2634_
timestamp 1608254825
transform 1 0 5428 0 -1 26656
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_44_84
timestamp 1608254825
transform 1 0 8832 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_74
timestamp 1608254825
transform 1 0 7912 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _1239_
timestamp 1608254825
transform 1 0 8004 0 -1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_44_113
timestamp 1608254825
transform 1 0 11500 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_100
timestamp 1608254825
transform 1 0 10304 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_96
timestamp 1608254825
transform 1 0 9936 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_427
timestamp 1608254825
transform 1 0 9568 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_4  _1352_
timestamp 1608254825
transform 1 0 10396 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1345_
timestamp 1608254825
transform 1 0 9660 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_44_126
timestamp 1608254825
transform 1 0 12696 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_44_120
timestamp 1608254825
transform 1 0 12144 0 -1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_4  _1757_
timestamp 1608254825
transform 1 0 12788 0 -1 26656
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _1332_
timestamp 1608254825
transform 1 0 11868 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_44_152
timestamp 1608254825
transform 1 0 15088 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_148
timestamp 1608254825
transform 1 0 14720 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_140
timestamp 1608254825
transform 1 0 13984 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_428
timestamp 1608254825
transform 1 0 15180 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__a21o_4  _2230_
timestamp 1608254825
transform 1 0 15272 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _1612_
timestamp 1608254825
transform 1 0 14352 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_179
timestamp 1608254825
transform 1 0 17572 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_166
timestamp 1608254825
transform 1 0 16376 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_4  _1414_
timestamp 1608254825
transform 1 0 16744 0 -1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_44_197
timestamp 1608254825
transform 1 0 19228 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__and3_4  _1412_
timestamp 1608254825
transform 1 0 19596 0 -1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__nand3_4  _1409_
timestamp 1608254825
transform 1 0 17940 0 -1 26656
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_6  FILLER_44_219
timestamp 1608254825
transform 1 0 21252 0 -1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_44_210
timestamp 1608254825
transform 1 0 20424 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_429
timestamp 1608254825
transform 1 0 20792 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__o41ai_4  _2216_
timestamp 1608254825
transform 1 0 21804 0 -1 26656
box -38 -48 2062 592
use sky130_fd_sc_hd__buf_2  _1406_
timestamp 1608254825
transform 1 0 20884 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_247
timestamp 1608254825
transform 1 0 23828 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__or4_4  _2234_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 24196 0 -1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_44_274
timestamp 1608254825
transform 1 0 26312 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_44_268
timestamp 1608254825
transform 1 0 25760 0 -1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_44_260
timestamp 1608254825
transform 1 0 25024 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1668_
timestamp 1608254825
transform 1 0 25392 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_289
timestamp 1608254825
transform 1 0 27692 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_285
timestamp 1608254825
transform 1 0 27324 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_430
timestamp 1608254825
transform 1 0 26404 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2391_
timestamp 1608254825
transform 1 0 27784 0 -1 26656
box -38 -48 1786 592
use sky130_fd_sc_hd__nor2_4  _2236_
timestamp 1608254825
transform 1 0 26496 0 -1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_44_309
timestamp 1608254825
transform 1 0 29532 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_4  _2323_
timestamp 1608254825
transform 1 0 29900 0 -1 26656
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_2  FILLER_44_337
timestamp 1608254825
transform 1 0 32108 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_334
timestamp 1608254825
transform 1 0 31832 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_44_326
timestamp 1608254825
transform 1 0 31096 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_431
timestamp 1608254825
transform 1 0 32016 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1186_
timestamp 1608254825
transform 1 0 32292 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_44_343
timestamp 1608254825
transform 1 0 32660 0 -1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  _2458_
timestamp 1608254825
transform 1 0 33212 0 -1 26656
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_44_368
timestamp 1608254825
transform 1 0 34960 0 -1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  _2468_
timestamp 1608254825
transform 1 0 35512 0 -1 26656
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_44_408
timestamp 1608254825
transform 1 0 38640 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_398
timestamp 1608254825
transform 1 0 37720 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_393
timestamp 1608254825
transform 1 0 37260 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_432
timestamp 1608254825
transform 1 0 37628 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _1738_
timestamp 1608254825
transform 1 0 37812 0 -1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_44_416
timestamp 1608254825
transform 1 0 39376 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1608254825
transform -1 0 39836 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_45_11
timestamp 1608254825
transform 1 0 2116 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_3
timestamp 1608254825
transform 1 0 1380 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1608254825
transform 1 0 1104 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_4  _2079_
timestamp 1608254825
transform 1 0 2208 0 1 26656
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_45_44
timestamp 1608254825
transform 1 0 5152 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_37
timestamp 1608254825
transform 1 0 4508 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_26
timestamp 1608254825
transform 1 0 3496 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__or2_4  _2081_
timestamp 1608254825
transform 1 0 3864 0 1 26656
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1327_
timestamp 1608254825
transform 1 0 4876 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_45_57
timestamp 1608254825
transform 1 0 6348 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_433
timestamp 1608254825
transform 1 0 6716 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_4  _1319_
timestamp 1608254825
transform 1 0 5520 0 1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_4  _1317_
timestamp 1608254825
transform 1 0 6808 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_88
timestamp 1608254825
transform 1 0 9200 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_78
timestamp 1608254825
transform 1 0 8280 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_74
timestamp 1608254825
transform 1 0 7912 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_4  _1240_
timestamp 1608254825
transform 1 0 8372 0 1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_45_113
timestamp 1608254825
transform 1 0 11500 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_45_106
timestamp 1608254825
transform 1 0 10856 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_4  _1353_
timestamp 1608254825
transform 1 0 9568 0 1 26656
box -38 -48 1326 592
use sky130_fd_sc_hd__inv_2  _1349_
timestamp 1608254825
transform 1 0 11224 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_45_130
timestamp 1608254825
transform 1 0 13064 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_126
timestamp 1608254825
transform 1 0 12696 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_121
timestamp 1608254825
transform 1 0 12236 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_434
timestamp 1608254825
transform 1 0 12328 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_4  _1658_
timestamp 1608254825
transform 1 0 13156 0 1 26656
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _1369_
timestamp 1608254825
transform 1 0 12420 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_45_159
timestamp 1608254825
transform 1 0 15732 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_151
timestamp 1608254825
transform 1 0 14996 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_144
timestamp 1608254825
transform 1 0 14352 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1656_
timestamp 1608254825
transform 1 0 15364 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1417_
timestamp 1608254825
transform 1 0 14720 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_45_182
timestamp 1608254825
transform 1 0 17848 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_45_176
timestamp 1608254825
transform 1 0 17296 0 1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_4  _1416_
timestamp 1608254825
transform 1 0 16100 0 1 26656
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_6  FILLER_45_184
timestamp 1608254825
transform 1 0 18032 0 1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_435
timestamp 1608254825
transform 1 0 17940 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__a41oi_4  _1407_
timestamp 1608254825
transform 1 0 18584 0 1 26656
box -38 -48 2062 592
use sky130_fd_sc_hd__decap_4  FILLER_45_212
timestamp 1608254825
transform 1 0 20608 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__o41ai_4  _2147_
timestamp 1608254825
transform 1 0 20976 0 1 26656
box -38 -48 2062 592
use sky130_fd_sc_hd__fill_2  FILLER_45_245
timestamp 1608254825
transform 1 0 23644 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_45_238
timestamp 1608254825
transform 1 0 23000 0 1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_436
timestamp 1608254825
transform 1 0 23552 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__or4_4  _1661_
timestamp 1608254825
transform 1 0 23828 0 1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_45_269
timestamp 1608254825
transform 1 0 25852 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_264
timestamp 1608254825
transform 1 0 25392 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_45_256
timestamp 1608254825
transform 1 0 24656 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1734_
timestamp 1608254825
transform 1 0 25576 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_45_294
timestamp 1608254825
transform 1 0 28152 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_281
timestamp 1608254825
transform 1 0 26956 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_4  _1727_
timestamp 1608254825
transform 1 0 27324 0 1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_45_315
timestamp 1608254825
transform 1 0 30084 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_45_301
timestamp 1608254825
transform 1 0 28796 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_437
timestamp 1608254825
transform 1 0 29164 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_4  _2214_
timestamp 1608254825
transform 1 0 29256 0 1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1697_
timestamp 1608254825
transform 1 0 28520 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_45_327
timestamp 1608254825
transform 1 0 31188 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2645_
timestamp 1608254825
transform 1 0 31556 0 1 26656
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  _1188_
timestamp 1608254825
transform 1 0 30820 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_365
timestamp 1608254825
transform 1 0 34684 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_361
timestamp 1608254825
transform 1 0 34316 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_350
timestamp 1608254825
transform 1 0 33304 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__or2_4  _2106_
timestamp 1608254825
transform 1 0 33672 0 1 26656
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_45_385
timestamp 1608254825
transform 1 0 36524 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_375
timestamp 1608254825
transform 1 0 35604 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_371
timestamp 1608254825
transform 1 0 35236 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_438
timestamp 1608254825
transform 1 0 34776 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _2092_
timestamp 1608254825
transform 1 0 35696 0 1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _1222_
timestamp 1608254825
transform 1 0 34868 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_393
timestamp 1608254825
transform 1 0 37260 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _2570_
timestamp 1608254825
transform 1 0 37444 0 1 26656
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_45_414
timestamp 1608254825
transform 1 0 39192 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1608254825
transform -1 0 39836 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_47_12
timestamp 1608254825
transform 1 0 2208 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_3
timestamp 1608254825
transform 1 0 1380 0 1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_46_22
timestamp 1608254825
transform 1 0 3128 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1608254825
transform 1 0 1104 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1608254825
transform 1 0 1104 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _2473_
timestamp 1608254825
transform 1 0 1380 0 -1 27744
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_2  _2080_
timestamp 1608254825
transform 1 0 1932 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__nand4_4  _1991_
timestamp 1608254825
transform 1 0 2576 0 1 27744
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_47_40
timestamp 1608254825
transform 1 0 4784 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_33
timestamp 1608254825
transform 1 0 4140 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_30
timestamp 1608254825
transform 1 0 3864 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_439
timestamp 1608254825
transform 1 0 3956 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2474_
timestamp 1608254825
transform 1 0 4048 0 -1 27744
box -38 -48 1786 592
use sky130_fd_sc_hd__a21oi_4  _2077_
timestamp 1608254825
transform 1 0 5152 0 1 27744
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _1359_
timestamp 1608254825
transform 1 0 4508 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_46_51
timestamp 1608254825
transform 1 0 5796 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_57
timestamp 1608254825
transform 1 0 6348 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_59
timestamp 1608254825
transform 1 0 6532 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1275_
timestamp 1608254825
transform 1 0 6164 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_66
timestamp 1608254825
transform 1 0 7176 0 1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_63
timestamp 1608254825
transform 1 0 6900 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_446
timestamp 1608254825
transform 1 0 6716 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1391_
timestamp 1608254825
transform 1 0 6808 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1253_
timestamp 1608254825
transform 1 0 6992 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_46_67
timestamp 1608254825
transform 1 0 7268 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_91
timestamp 1608254825
transform 1 0 9476 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_88
timestamp 1608254825
transform 1 0 9200 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_75
timestamp 1608254825
transform 1 0 8004 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2627_
timestamp 1608254825
transform 1 0 7728 0 1 27744
box -38 -48 1786 592
use sky130_fd_sc_hd__nand2_4  _1354_
timestamp 1608254825
transform 1 0 8372 0 -1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _1274_
timestamp 1608254825
transform 1 0 7636 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_109
timestamp 1608254825
transform 1 0 11132 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_104
timestamp 1608254825
transform 1 0 10672 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_93
timestamp 1608254825
transform 1 0 9660 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_440
timestamp 1608254825
transform 1 0 9568 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2628_
timestamp 1608254825
transform 1 0 11040 0 -1 27744
box -38 -48 1786 592
use sky130_fd_sc_hd__nand3_4  _1358_
timestamp 1608254825
transform 1 0 9844 0 1 27744
box -38 -48 1326 592
use sky130_fd_sc_hd__inv_2  _1355_
timestamp 1608254825
transform 1 0 11500 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_4  _1228_
timestamp 1608254825
transform 1 0 9844 0 -1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_47_126
timestamp 1608254825
transform 1 0 12696 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_47_116
timestamp 1608254825
transform 1 0 11776 0 1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_46_127
timestamp 1608254825
transform 1 0 12788 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_447
timestamp 1608254825
transform 1 0 12328 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_4  _1721_
timestamp 1608254825
transform 1 0 13432 0 1 27744
box -38 -48 1234 592
use sky130_fd_sc_hd__a21oi_4  _1657_
timestamp 1608254825
transform 1 0 13156 0 -1 27744
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _1356_
timestamp 1608254825
transform 1 0 12420 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_47_158
timestamp 1608254825
transform 1 0 15640 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_147
timestamp 1608254825
transform 1 0 14628 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_154
timestamp 1608254825
transform 1 0 15272 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_46_152
timestamp 1608254825
transform 1 0 15088 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_144
timestamp 1608254825
transform 1 0 14352 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_441
timestamp 1608254825
transform 1 0 15180 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1413_
timestamp 1608254825
transform 1 0 15548 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1378_
timestamp 1608254825
transform 1 0 15364 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_47_179
timestamp 1608254825
transform 1 0 17572 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_162
timestamp 1608254825
transform 1 0 16008 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_160
timestamp 1608254825
transform 1 0 15824 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_m1_clk_local
timestamp 1608254825
transform 1 0 16100 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _2614_
timestamp 1608254825
transform 1 0 16192 0 -1 27744
box -38 -48 1786 592
use sky130_fd_sc_hd__a21oi_4  _1415_
timestamp 1608254825
transform 1 0 16376 0 1 27744
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_47_194
timestamp 1608254825
transform 1 0 18952 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_184
timestamp 1608254825
transform 1 0 18032 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_46_191
timestamp 1608254825
transform 1 0 18676 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_183
timestamp 1608254825
transform 1 0 17940 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_448
timestamp 1608254825
transform 1 0 17940 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_4  _2166_
timestamp 1608254825
transform 1 0 18124 0 1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_4  _1401_
timestamp 1608254825
transform 1 0 18768 0 -1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_46_201
timestamp 1608254825
transform 1 0 19596 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1396_
timestamp 1608254825
transform 1 0 19964 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _2615_
timestamp 1608254825
transform 1 0 19320 0 1 27744
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_47_225
timestamp 1608254825
transform 1 0 21804 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_47_217
timestamp 1608254825
transform 1 0 21068 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_46_219
timestamp 1608254825
transform 1 0 21252 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_208
timestamp 1608254825
transform 1 0 20240 0 -1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_442
timestamp 1608254825
transform 1 0 20792 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_4  _1760_
timestamp 1608254825
transform 1 0 21988 0 1 27744
box -38 -48 1234 592
use sky130_fd_sc_hd__a21o_4  _1725_
timestamp 1608254825
transform 1 0 21620 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _1666_
timestamp 1608254825
transform 1 0 20884 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_240
timestamp 1608254825
transform 1 0 23184 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_248
timestamp 1608254825
transform 1 0 23920 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_235
timestamp 1608254825
transform 1 0 22724 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_449
timestamp 1608254825
transform 1 0 23552 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__or4_4  _1860_
timestamp 1608254825
transform 1 0 23092 0 -1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__nor4_4  _1673_
timestamp 1608254825
transform 1 0 23644 0 1 27744
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_1  FILLER_47_268
timestamp 1608254825
transform 1 0 25760 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_47_262
timestamp 1608254825
transform 1 0 25208 0 1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_46_267
timestamp 1608254825
transform 1 0 25668 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_252
timestamp 1608254825
transform 1 0 24288 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2596_
timestamp 1608254825
transform 1 0 25852 0 1 27744
box -38 -48 1786 592
use sky130_fd_sc_hd__nand3_4  _1674_
timestamp 1608254825
transform 1 0 24380 0 -1 27744
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_47_288
timestamp 1608254825
transform 1 0 27600 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_285
timestamp 1608254825
transform 1 0 27324 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_443
timestamp 1608254825
transform 1 0 26404 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2593_
timestamp 1608254825
transform 1 0 27692 0 -1 27744
box -38 -48 1786 592
use sky130_fd_sc_hd__nand2_4  _1726_
timestamp 1608254825
transform 1 0 27968 0 1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  _1677_
timestamp 1608254825
transform 1 0 26496 0 -1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_47_306
timestamp 1608254825
transform 1 0 29256 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_301
timestamp 1608254825
transform 1 0 28796 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_308
timestamp 1608254825
transform 1 0 29440 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_450
timestamp 1608254825
transform 1 0 29164 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_4  _2355_
timestamp 1608254825
transform 1 0 29808 0 -1 27744
box -38 -48 1234 592
use sky130_fd_sc_hd__o21ai_4  _1214_
timestamp 1608254825
transform 1 0 29624 0 1 27744
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_47_340
timestamp 1608254825
transform 1 0 32384 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_323
timestamp 1608254825
transform 1 0 30820 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_332
timestamp 1608254825
transform 1 0 31648 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_325
timestamp 1608254825
transform 1 0 31004 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_444
timestamp 1608254825
transform 1 0 32016 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_4  _2356_
timestamp 1608254825
transform 1 0 31188 0 1 27744
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _1839_
timestamp 1608254825
transform 1 0 31372 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_4  _1216_
timestamp 1608254825
transform 1 0 32108 0 -1 27744
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_47_362
timestamp 1608254825
transform 1 0 34408 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_347
timestamp 1608254825
transform 1 0 33028 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_351
timestamp 1608254825
transform 1 0 33396 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_14_0_addressalyzerBlock.SPI_CLK
timestamp 1608254825
transform 1 0 32752 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_4  _1215_
timestamp 1608254825
transform 1 0 33764 0 -1 27744
box -38 -48 1234 592
use sky130_fd_sc_hd__o21ai_4  _1211_
timestamp 1608254825
transform 1 0 33212 0 1 27744
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_6  FILLER_47_371
timestamp 1608254825
transform 1 0 35236 0 1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_367
timestamp 1608254825
transform 1 0 34868 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_379
timestamp 1608254825
transform 1 0 35972 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_368
timestamp 1608254825
transform 1 0 34960 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_451
timestamp 1608254825
transform 1 0 34776 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2460_
timestamp 1608254825
transform 1 0 35788 0 1 27744
box -38 -48 1786 592
use sky130_fd_sc_hd__and4_4  _2104_
timestamp 1608254825
transform 1 0 36340 0 -1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__or2_4  _1210_
timestamp 1608254825
transform 1 0 35328 0 -1 27744
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1180_
timestamp 1608254825
transform 1 0 34960 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_47_396
timestamp 1608254825
transform 1 0 37536 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_407
timestamp 1608254825
transform 1 0 38548 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_396
timestamp 1608254825
transform 1 0 37536 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_392
timestamp 1608254825
transform 1 0 37168 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_445
timestamp 1608254825
transform 1 0 37628 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_4  _2112_
timestamp 1608254825
transform 1 0 37720 0 -1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_4  _1835_
timestamp 1608254825
transform 1 0 37904 0 1 27744
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _1683_
timestamp 1608254825
transform 1 0 38916 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_47_417
timestamp 1608254825
transform 1 0 39468 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_413
timestamp 1608254825
transform 1 0 39100 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_414
timestamp 1608254825
transform 1 0 39192 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1608254825
transform -1 0 39836 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1608254825
transform -1 0 39836 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_48_18
timestamp 1608254825
transform 1 0 2760 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_3
timestamp 1608254825
transform 1 0 1380 0 -1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1608254825
transform 1 0 1104 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__and3_4  _2084_
timestamp 1608254825
transform 1 0 1932 0 -1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _2058_
timestamp 1608254825
transform 1 0 3128 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_41
timestamp 1608254825
transform 1 0 4876 0 -1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_30
timestamp 1608254825
transform 1 0 3864 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_26
timestamp 1608254825
transform 1 0 3496 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_452
timestamp 1608254825
transform 1 0 3956 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__and3_4  _2082_
timestamp 1608254825
transform 1 0 4048 0 -1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_48_66
timestamp 1608254825
transform 1 0 7176 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2475_
timestamp 1608254825
transform 1 0 5428 0 -1 28832
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_48_88
timestamp 1608254825
transform 1 0 9200 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_74
timestamp 1608254825
transform 1 0 7912 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_48_70
timestamp 1608254825
transform 1 0 7544 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_m1_clk_local
timestamp 1608254825
transform 1 0 7636 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_4  _1357_
timestamp 1608254825
transform 1 0 8004 0 -1 28832
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_2  FILLER_48_114
timestamp 1608254825
transform 1 0 11592 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_107
timestamp 1608254825
transform 1 0 10948 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_93
timestamp 1608254825
transform 1 0 9660 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_9_0_m1_clk_local
timestamp 1608254825
transform 1 0 11316 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_453
timestamp 1608254825
transform 1 0 9568 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__nor3_4  _1351_
timestamp 1608254825
transform 1 0 9752 0 -1 28832
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_48_129
timestamp 1608254825
transform 1 0 12972 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_4  _1859_
timestamp 1608254825
transform 1 0 11776 0 -1 28832
box -38 -48 1234 592
use sky130_fd_sc_hd__a21oi_4  _1858_
timestamp 1608254825
transform 1 0 13340 0 -1 28832
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_1  FILLER_48_152
timestamp 1608254825
transform 1 0 15088 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_48_146
timestamp 1608254825
transform 1 0 14536 0 -1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_454
timestamp 1608254825
transform 1 0 15180 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2624_
timestamp 1608254825
transform 1 0 15272 0 -1 28832
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_48_182
timestamp 1608254825
transform 1 0 17848 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_173
timestamp 1608254825
transform 1 0 17020 0 -1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1410_
timestamp 1608254825
transform 1 0 17572 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_48_205
timestamp 1608254825
transform 1 0 19964 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _2616_
timestamp 1608254825
transform 1 0 18216 0 -1 28832
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_48_219
timestamp 1608254825
transform 1 0 21252 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_215
timestamp 1608254825
transform 1 0 20884 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_213
timestamp 1608254825
transform 1 0 20700 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_455
timestamp 1608254825
transform 1 0 20792 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_4  _1723_
timestamp 1608254825
transform 1 0 21344 0 -1 28832
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_48_245
timestamp 1608254825
transform 1 0 23644 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_233
timestamp 1608254825
transform 1 0 22540 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__nand3_4  _1861_
timestamp 1608254825
transform 1 0 24012 0 -1 28832
box -38 -48 1326 592
use sky130_fd_sc_hd__buf_2  _1672_
timestamp 1608254825
transform 1 0 23276 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_271
timestamp 1608254825
transform 1 0 26036 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_263
timestamp 1608254825
transform 1 0 25300 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1675_
timestamp 1608254825
transform 1 0 25668 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_289
timestamp 1608254825
transform 1 0 27692 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_285
timestamp 1608254825
transform 1 0 27324 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_456
timestamp 1608254825
transform 1 0 26404 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2436_
timestamp 1608254825
transform 1 0 27784 0 -1 28832
box -38 -48 1786 592
use sky130_fd_sc_hd__nand2_4  _1676_
timestamp 1608254825
transform 1 0 26496 0 -1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_48_309
timestamp 1608254825
transform 1 0 29532 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_4  _1208_
timestamp 1608254825
transform 1 0 29900 0 -1 28832
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_48_342
timestamp 1608254825
transform 1 0 32568 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_337
timestamp 1608254825
transform 1 0 32108 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_334
timestamp 1608254825
transform 1 0 31832 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_48_326
timestamp 1608254825
transform 1 0 31096 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_457
timestamp 1608254825
transform 1 0 32016 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _2103_
timestamp 1608254825
transform 1 0 32292 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_48_349
timestamp 1608254825
transform 1 0 33212 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2646_
timestamp 1608254825
transform 1 0 33580 0 -1 28832
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_2  _1837_
timestamp 1608254825
transform 1 0 32936 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_48_372
timestamp 1608254825
transform 1 0 35328 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_4  _1840_
timestamp 1608254825
transform 1 0 35696 0 -1 28832
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_6  FILLER_48_411
timestamp 1608254825
transform 1 0 38916 0 -1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_398
timestamp 1608254825
transform 1 0 37720 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_48_396
timestamp 1608254825
transform 1 0 37536 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_48_390
timestamp 1608254825
transform 1 0 36984 0 -1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_458
timestamp 1608254825
transform 1 0 37628 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__a21o_4  _1836_
timestamp 1608254825
transform 1 0 37812 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_417
timestamp 1608254825
transform 1 0 39468 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1608254825
transform -1 0 39836 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_49_10
timestamp 1608254825
transform 1 0 2024 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_3
timestamp 1608254825
transform 1 0 1380 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1608254825
transform 1 0 1104 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2070_
timestamp 1608254825
transform 1 0 1748 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_4  _2053_
timestamp 1608254825
transform 1 0 2392 0 1 28832
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_6  FILLER_49_44
timestamp 1608254825
transform 1 0 5152 0 1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_49_27
timestamp 1608254825
transform 1 0 3588 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_4  _2069_
timestamp 1608254825
transform 1 0 3956 0 1 28832
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_49_66
timestamp 1608254825
transform 1 0 7176 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_57
timestamp 1608254825
transform 1 0 6348 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_8_0_m1_clk_local
timestamp 1608254825
transform 1 0 5704 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_459
timestamp 1608254825
transform 1 0 6716 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1374_
timestamp 1608254825
transform 1 0 5980 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1306_
timestamp 1608254825
transform 1 0 6808 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_90
timestamp 1608254825
transform 1 0 9384 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_74
timestamp 1608254825
transform 1 0 7912 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_4  _1362_
timestamp 1608254825
transform 1 0 8280 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _1283_
timestamp 1608254825
transform 1 0 7544 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_107
timestamp 1608254825
transform 1 0 10948 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _2027_
timestamp 1608254825
transform 1 0 11316 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_4  _1371_
timestamp 1608254825
transform 1 0 9752 0 1 28832
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_1  FILLER_49_121
timestamp 1608254825
transform 1 0 12236 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_49_115
timestamp 1608254825
transform 1 0 11684 0 1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_460
timestamp 1608254825
transform 1 0 12328 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2626_
timestamp 1608254825
transform 1 0 12420 0 1 28832
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_49_149
timestamp 1608254825
transform 1 0 14812 0 1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_49_142
timestamp 1608254825
transform 1 0 14168 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__and4_4  _1373_
timestamp 1608254825
transform 1 0 15364 0 1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1237_
timestamp 1608254825
transform 1 0 14536 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_49_179
timestamp 1608254825
transform 1 0 17572 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_172
timestamp 1608254825
transform 1 0 16928 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_164
timestamp 1608254825
transform 1 0 16192 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1404_
timestamp 1608254825
transform 1 0 17296 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1388_
timestamp 1608254825
transform 1 0 16560 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_203
timestamp 1608254825
transform 1 0 19780 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_49_197
timestamp 1608254825
transform 1 0 19228 0 1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_461
timestamp 1608254825
transform 1 0 17940 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_4  _2167_
timestamp 1608254825
transform 1 0 19872 0 1 28832
box -38 -48 1234 592
use sky130_fd_sc_hd__nor3_4  _1408_
timestamp 1608254825
transform 1 0 18032 0 1 28832
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_49_217
timestamp 1608254825
transform 1 0 21068 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_4  _1759_
timestamp 1608254825
transform 1 0 21436 0 1 28832
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_2  FILLER_49_242
timestamp 1608254825
transform 1 0 23368 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_49_234
timestamp 1608254825
transform 1 0 22632 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_462
timestamp 1608254825
transform 1 0 23552 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__a22oi_4  _2213_
timestamp 1608254825
transform 1 0 23644 0 1 28832
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_49_262
timestamp 1608254825
transform 1 0 25208 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_4  _1763_
timestamp 1608254825
transform 1 0 25576 0 1 28832
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_49_296
timestamp 1608254825
transform 1 0 28336 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_279
timestamp 1608254825
transform 1 0 26772 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_4  _2215_
timestamp 1608254825
transform 1 0 27140 0 1 28832
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_49_313
timestamp 1608254825
transform 1 0 29900 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_49_306
timestamp 1608254825
transform 1 0 29256 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_49_303
timestamp 1608254825
transform 1 0 28980 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_12_0_addressalyzerBlock.SPI_CLK
timestamp 1608254825
transform 1 0 28704 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_463
timestamp 1608254825
transform 1 0 29164 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2652_
timestamp 1608254825
transform 1 0 30268 0 1 28832
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  _1213_
timestamp 1608254825
transform 1 0 29532 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_336
timestamp 1608254825
transform 1 0 32016 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_4  _2354_
timestamp 1608254825
transform 1 0 32384 0 1 28832
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_1  FILLER_49_365
timestamp 1608254825
transform 1 0 34684 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_361
timestamp 1608254825
transform 1 0 34316 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_353
timestamp 1608254825
transform 1 0 33580 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1181_
timestamp 1608254825
transform 1 0 33948 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_388
timestamp 1608254825
transform 1 0 36800 0 1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_49_380
timestamp 1608254825
transform 1 0 36064 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_464
timestamp 1608254825
transform 1 0 34776 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_4  _1207_
timestamp 1608254825
transform 1 0 34868 0 1 28832
box -38 -48 1234 592
use sky130_fd_sc_hd__buf_2  _1178_
timestamp 1608254825
transform 1 0 36432 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_411
timestamp 1608254825
transform 1 0 38916 0 1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__nand4_4  _1735_
timestamp 1608254825
transform 1 0 37352 0 1 28832
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_1  FILLER_49_417
timestamp 1608254825
transform 1 0 39468 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1608254825
transform -1 0 39836 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_50_22
timestamp 1608254825
transform 1 0 3128 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1608254825
transform 1 0 1104 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _2477_
timestamp 1608254825
transform 1 0 1380 0 -1 29920
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_50_45
timestamp 1608254825
transform 1 0 5244 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_30
timestamp 1608254825
transform 1 0 3864 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_465
timestamp 1608254825
transform 1 0 3956 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_4  _2068_
timestamp 1608254825
transform 1 0 4048 0 -1 29920
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_50_62
timestamp 1608254825
transform 1 0 6808 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_4  _2076_
timestamp 1608254825
transform 1 0 5612 0 -1 29920
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_4  _1990_
timestamp 1608254825
transform 1 0 7176 0 -1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_50_91
timestamp 1608254825
transform 1 0 9476 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_83
timestamp 1608254825
transform 1 0 8740 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_50_75
timestamp 1608254825
transform 1 0 8004 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1269_
timestamp 1608254825
transform 1 0 8372 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_50_113
timestamp 1608254825
transform 1 0 11500 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_93
timestamp 1608254825
transform 1 0 9660 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_466
timestamp 1608254825
transform 1 0 9568 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2625_
timestamp 1608254825
transform 1 0 9752 0 -1 29920
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_50_121
timestamp 1608254825
transform 1 0 12236 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__nand4_4  _1367_
timestamp 1608254825
transform 1 0 12328 0 -1 29920
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_6  FILLER_50_147
timestamp 1608254825
transform 1 0 14628 0 -1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_50_139
timestamp 1608254825
transform 1 0 13892 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_467
timestamp 1608254825
transform 1 0 15180 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__nand3_4  _1376_
timestamp 1608254825
transform 1 0 15272 0 -1 29920
box -38 -48 1326 592
use sky130_fd_sc_hd__buf_2  _1372_
timestamp 1608254825
transform 1 0 14260 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_172
timestamp 1608254825
transform 1 0 16928 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_168
timestamp 1608254825
transform 1 0 16560 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_4  _1402_
timestamp 1608254825
transform 1 0 17020 0 -1 29920
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_50_203
timestamp 1608254825
transform 1 0 19780 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_186
timestamp 1608254825
transform 1 0 18216 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_4  _1403_
timestamp 1608254825
transform 1 0 18584 0 -1 29920
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_8  FILLER_50_228
timestamp 1608254825
transform 1 0 22080 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_50_210
timestamp 1608254825
transform 1 0 20424 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_468
timestamp 1608254825
transform 1 0 20792 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_4  _1398_
timestamp 1608254825
transform 1 0 20884 0 -1 29920
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _1230_
timestamp 1608254825
transform 1 0 20148 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_50_236
timestamp 1608254825
transform 1 0 22816 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__a22oi_4  _2191_
timestamp 1608254825
transform 1 0 23000 0 -1 29920
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_1  FILLER_50_274
timestamp 1608254825
transform 1 0 26312 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_50_268
timestamp 1608254825
transform 1 0 25760 0 -1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_50_255
timestamp 1608254825
transform 1 0 24564 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_4  _1739_
timestamp 1608254825
transform 1 0 24932 0 -1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_50_293
timestamp 1608254825
transform 1 0 28060 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_276
timestamp 1608254825
transform 1 0 26496 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_469
timestamp 1608254825
transform 1 0 26404 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_4  _2193_
timestamp 1608254825
transform 1 0 26864 0 -1 29920
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_1  FILLER_50_307
timestamp 1608254825
transform 1 0 29348 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_50_301
timestamp 1608254825
transform 1 0 28796 0 -1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _1761_
timestamp 1608254825
transform 1 0 28428 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_4  _1192_
timestamp 1608254825
transform 1 0 29440 0 -1 29920
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_50_337
timestamp 1608254825
transform 1 0 32108 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_332
timestamp 1608254825
transform 1 0 31648 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_321
timestamp 1608254825
transform 1 0 30636 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_addressalyzerBlock.SPI_CLK
timestamp 1608254825
transform 1 0 31004 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_470
timestamp 1608254825
transform 1 0 32016 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _2353_
timestamp 1608254825
transform 1 0 32476 0 -1 29920
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _1187_
timestamp 1608254825
transform 1 0 31280 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_352
timestamp 1608254825
transform 1 0 33488 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_348
timestamp 1608254825
transform 1 0 33120 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2647_
timestamp 1608254825
transform 1 0 33580 0 -1 29920
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_50_380
timestamp 1608254825
transform 1 0 36064 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_376
timestamp 1608254825
transform 1 0 35696 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_372
timestamp 1608254825
transform 1 0 35328 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1834_
timestamp 1608254825
transform 1 0 35788 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_4  _1833_
timestamp 1608254825
transform 1 0 36432 0 -1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_50_407
timestamp 1608254825
transform 1 0 38548 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_393
timestamp 1608254825
transform 1 0 37260 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_471
timestamp 1608254825
transform 1 0 37628 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_4  _1831_
timestamp 1608254825
transform 1 0 37720 0 -1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1737_
timestamp 1608254825
transform 1 0 38916 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_50_414
timestamp 1608254825
transform 1 0 39192 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1608254825
transform -1 0 39836 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_51_9
timestamp 1608254825
transform 1 0 1932 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_51_3
timestamp 1608254825
transform 1 0 1380 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1608254825
transform 1 0 1104 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__nor4_4  _1992_
timestamp 1608254825
transform 1 0 2300 0 1 29920
box -38 -48 1602 592
use sky130_fd_sc_hd__inv_2  _1988_
timestamp 1608254825
transform 1 0 1656 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_51_43
timestamp 1608254825
transform 1 0 5060 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_30
timestamp 1608254825
transform 1 0 3864 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_4  _2060_
timestamp 1608254825
transform 1 0 4232 0 1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_51_57
timestamp 1608254825
transform 1 0 6348 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_47
timestamp 1608254825
transform 1 0 5428 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_472
timestamp 1608254825
transform 1 0 6716 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_4  _2073_
timestamp 1608254825
transform 1 0 6808 0 1 29920
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_4  _2072_
timestamp 1608254825
transform 1 0 5520 0 1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_51_90
timestamp 1608254825
transform 1 0 9384 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_83
timestamp 1608254825
transform 1 0 8740 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_75
timestamp 1608254825
transform 1 0 8004 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_m1_clk_local
timestamp 1608254825
transform 1 0 9108 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_4  _1370_
timestamp 1608254825
transform 1 0 9476 0 1 29920
box -38 -48 1234 592
use sky130_fd_sc_hd__buf_2  _1270_
timestamp 1608254825
transform 1 0 8372 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_104
timestamp 1608254825
transform 1 0 10672 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_4  _1361_
timestamp 1608254825
transform 1 0 11040 0 1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_51_132
timestamp 1608254825
transform 1 0 13248 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_121
timestamp 1608254825
transform 1 0 12236 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_117
timestamp 1608254825
transform 1 0 11868 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_473
timestamp 1608254825
transform 1 0 12328 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_4  _1368_
timestamp 1608254825
transform 1 0 12420 0 1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__nand4_4  _1238_
timestamp 1608254825
transform 1 0 13616 0 1 29920
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_51_153
timestamp 1608254825
transform 1 0 15180 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_4  _1375_
timestamp 1608254825
transform 1 0 15548 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_179
timestamp 1608254825
transform 1 0 17572 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_175
timestamp 1608254825
transform 1 0 17204 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_51_169
timestamp 1608254825
transform 1 0 16652 0 1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1229_
timestamp 1608254825
transform 1 0 17296 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_51_203
timestamp 1608254825
transform 1 0 19780 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_474
timestamp 1608254825
transform 1 0 17940 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2617_
timestamp 1608254825
transform 1 0 18032 0 1 29920
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_51_220
timestamp 1608254825
transform 1 0 21344 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_4  _1399_
timestamp 1608254825
transform 1 0 21712 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__nor3_4  _1397_
timestamp 1608254825
transform 1 0 20148 0 1 29920
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_8  FILLER_51_236
timestamp 1608254825
transform 1 0 22816 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_475
timestamp 1608254825
transform 1 0 23552 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _2168_
timestamp 1608254825
transform 1 0 23644 0 1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_51_258
timestamp 1608254825
transform 1 0 24840 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_254
timestamp 1608254825
transform 1 0 24472 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2590_
timestamp 1608254825
transform 1 0 24932 0 1 29920
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_51_278
timestamp 1608254825
transform 1 0 26680 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2437_
timestamp 1608254825
transform 1 0 27048 0 1 29920
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_51_319
timestamp 1608254825
transform 1 0 30452 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_301
timestamp 1608254825
transform 1 0 28796 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_476
timestamp 1608254825
transform 1 0 29164 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_4  _1204_
timestamp 1608254825
transform 1 0 29256 0 1 29920
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_6  FILLER_51_342
timestamp 1608254825
transform 1 0 32568 0 1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  _2651_
timestamp 1608254825
transform 1 0 30820 0 1 29920
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_51_362
timestamp 1608254825
transform 1 0 34408 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_348
timestamp 1608254825
transform 1 0 33120 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_4  _1209_
timestamp 1608254825
transform 1 0 33212 0 1 29920
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_51_374
timestamp 1608254825
transform 1 0 35512 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_477
timestamp 1608254825
transform 1 0 34776 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2569_
timestamp 1608254825
transform 1 0 35880 0 1 29920
box -38 -48 1786 592
use sky130_fd_sc_hd__or2_4  _1206_
timestamp 1608254825
transform 1 0 34868 0 1 29920
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_51_397
timestamp 1608254825
transform 1 0 37628 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_4  _1832_
timestamp 1608254825
transform 1 0 37996 0 1 29920
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_51_414
timestamp 1608254825
transform 1 0 39192 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1608254825
transform -1 0 39836 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_53_22
timestamp 1608254825
transform 1 0 3128 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_10
timestamp 1608254825
transform 1 0 2024 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_3
timestamp 1608254825
transform 1 0 1380 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1608254825
transform 1 0 1104 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1608254825
transform 1 0 1104 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _2478_
timestamp 1608254825
transform 1 0 1380 0 1 31008
box -38 -48 1786 592
use sky130_fd_sc_hd__nor3_4  _2067_
timestamp 1608254825
transform 1 0 2392 0 -1 31008
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _1989_
timestamp 1608254825
transform 1 0 1748 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_53_39
timestamp 1608254825
transform 1 0 4692 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_42
timestamp 1608254825
transform 1 0 4968 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_52_36
timestamp 1608254825
transform 1 0 4416 0 -1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_52_27
timestamp 1608254825
transform 1 0 3588 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_478
timestamp 1608254825
transform 1 0 3956 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2476_
timestamp 1608254825
transform 1 0 5060 0 -1 31008
box -38 -48 1786 592
use sky130_fd_sc_hd__a21oi_4  _2066_
timestamp 1608254825
transform 1 0 3496 0 1 31008
box -38 -48 1234 592
use sky130_fd_sc_hd__buf_2  _2059_
timestamp 1608254825
transform 1 0 4048 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_57
timestamp 1608254825
transform 1 0 6348 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_50
timestamp 1608254825
transform 1 0 5704 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2071_
timestamp 1608254825
transform 1 0 5428 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2039_
timestamp 1608254825
transform 1 0 6072 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_53_66
timestamp 1608254825
transform 1 0 7176 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_62
timestamp 1608254825
transform 1 0 6808 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_62
timestamp 1608254825
transform 1 0 6808 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_485
timestamp 1608254825
transform 1 0 6716 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2486_
timestamp 1608254825
transform 1 0 7268 0 1 31008
box -38 -48 1786 592
use sky130_fd_sc_hd__a21o_4  _2074_
timestamp 1608254825
transform 1 0 7176 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_86
timestamp 1608254825
transform 1 0 9016 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_52_86
timestamp 1608254825
transform 1 0 9016 0 -1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_52_78
timestamp 1608254825
transform 1 0 8280 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_4  _1995_
timestamp 1608254825
transform 1 0 9384 0 1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _1298_
timestamp 1608254825
transform 1 0 8648 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_105
timestamp 1608254825
transform 1 0 10764 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_53_99
timestamp 1608254825
transform 1 0 10212 0 1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_52_113
timestamp 1608254825
transform 1 0 11500 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_52_105
timestamp 1608254825
transform 1 0 10764 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_52_97
timestamp 1608254825
transform 1 0 10028 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_479
timestamp 1608254825
transform 1 0 9568 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_4  _1382_
timestamp 1608254825
transform 1 0 10856 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _1350_
timestamp 1608254825
transform 1 0 10396 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1346_
timestamp 1608254825
transform 1 0 9660 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_118
timestamp 1608254825
transform 1 0 11960 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_134
timestamp 1608254825
transform 1 0 13432 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_486
timestamp 1608254825
transform 1 0 12328 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2623_
timestamp 1608254825
transform 1 0 11684 0 -1 31008
box -38 -48 1786 592
use sky130_fd_sc_hd__a41oi_4  _1381_
timestamp 1608254825
transform 1 0 12420 0 1 31008
box -38 -48 2062 592
use sky130_fd_sc_hd__decap_4  FILLER_53_158
timestamp 1608254825
transform 1 0 15640 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_145
timestamp 1608254825
transform 1 0 14444 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_52_158
timestamp 1608254825
transform 1 0 15640 0 -1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_52_147
timestamp 1608254825
transform 1 0 14628 0 -1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_480
timestamp 1608254825
transform 1 0 15180 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_4  _1377_
timestamp 1608254825
transform 1 0 14812 0 1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _1364_
timestamp 1608254825
transform 1 0 15272 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_4  _1236_
timestamp 1608254825
transform 1 0 13800 0 -1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_53_179
timestamp 1608254825
transform 1 0 17572 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_171
timestamp 1608254825
transform 1 0 16836 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_52_181
timestamp 1608254825
transform 1 0 17756 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_52_173
timestamp 1608254825
transform 1 0 17020 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1380_
timestamp 1608254825
transform 1 0 17204 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1366_
timestamp 1608254825
transform 1 0 17388 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__and4_4  _1365_
timestamp 1608254825
transform 1 0 16008 0 1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  _1234_
timestamp 1608254825
transform 1 0 16192 0 -1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_53_189
timestamp 1608254825
transform 1 0 18492 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_184
timestamp 1608254825
transform 1 0 18032 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_487
timestamp 1608254825
transform 1 0 17940 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1379_
timestamp 1608254825
transform 1 0 18124 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_4  _1363_
timestamp 1608254825
transform 1 0 18860 0 1 31008
box -38 -48 1234 592
use sky130_fd_sc_hd__nor4_4  _1233_
timestamp 1608254825
transform 1 0 18492 0 -1 31008
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_53_226
timestamp 1608254825
transform 1 0 21896 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_219
timestamp 1608254825
transform 1 0 21252 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_206
timestamp 1608254825
transform 1 0 20056 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_215
timestamp 1608254825
transform 1 0 20884 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_52_206
timestamp 1608254825
transform 1 0 20056 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_481
timestamp 1608254825
transform 1 0 20792 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2618_
timestamp 1608254825
transform 1 0 21252 0 -1 31008
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_2  _1400_
timestamp 1608254825
transform 1 0 21620 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_4  _1231_
timestamp 1608254825
transform 1 0 20424 0 1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_53_245
timestamp 1608254825
transform 1 0 23644 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_240
timestamp 1608254825
transform 1 0 23184 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_230
timestamp 1608254825
transform 1 0 22264 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_238
timestamp 1608254825
transform 1 0 23000 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_488
timestamp 1608254825
transform 1 0 23552 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__or3_4  _2352_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 22356 0 1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__or3_4  _2351_
timestamp 1608254825
transform 1 0 23828 0 1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__a22oi_4  _2169_
timestamp 1608254825
transform 1 0 23368 0 -1 31008
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_3  FILLER_53_268
timestamp 1608254825
transform 1 0 25760 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_53_256
timestamp 1608254825
transform 1 0 24656 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_274
timestamp 1608254825
transform 1 0 26312 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_266
timestamp 1608254825
transform 1 0 25576 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_52_259
timestamp 1608254825
transform 1 0 24932 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_4  _1762_
timestamp 1608254825
transform 1 0 26036 0 1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1740_
timestamp 1608254825
transform 1 0 25300 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_53_293
timestamp 1608254825
transform 1 0 28060 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_280
timestamp 1608254825
transform 1 0 26864 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_52_292
timestamp 1608254825
transform 1 0 27968 0 -1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_52_276
timestamp 1608254825
transform 1 0 26496 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_482
timestamp 1608254825
transform 1 0 26404 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_4  _2171_
timestamp 1608254825
transform 1 0 26772 0 -1 31008
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_4  _1862_
timestamp 1608254825
transform 1 0 27232 0 1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_53_304
timestamp 1608254825
transform 1 0 29072 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_300
timestamp 1608254825
transform 1 0 28704 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_298
timestamp 1608254825
transform 1 0 28520 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_addressalyzerBlock.SPI_CLK
timestamp 1608254825
transform 1 0 28428 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_addressalyzerBlock.SPI_CLK
timestamp 1608254825
transform 1 0 28612 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_489
timestamp 1608254825
transform 1 0 29164 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_4  _2170_
timestamp 1608254825
transform 1 0 29256 0 1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_53_315
timestamp 1608254825
transform 1 0 30084 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_315
timestamp 1608254825
transform 1 0 30084 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_4  _1200_
timestamp 1608254825
transform 1 0 28888 0 -1 31008
box -38 -48 1234 592
use sky130_fd_sc_hd__a21oi_4  _1197_
timestamp 1608254825
transform 1 0 30452 0 1 31008
box -38 -48 1234 592
use sky130_fd_sc_hd__a21oi_4  _1193_
timestamp 1608254825
transform 1 0 30452 0 -1 31008
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_6  FILLER_53_332
timestamp 1608254825
transform 1 0 31648 0 1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_52_332
timestamp 1608254825
transform 1 0 31648 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_483
timestamp 1608254825
transform 1 0 32016 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_4  _1195_
timestamp 1608254825
transform 1 0 32200 0 1 31008
box -38 -48 1234 592
use sky130_fd_sc_hd__o21ai_4  _1183_
timestamp 1608254825
transform 1 0 32108 0 -1 31008
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_53_362
timestamp 1608254825
transform 1 0 34408 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_351
timestamp 1608254825
transform 1 0 33396 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_358
timestamp 1608254825
transform 1 0 34040 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_350
timestamp 1608254825
transform 1 0 33304 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_4  _1205_
timestamp 1608254825
transform 1 0 34132 0 -1 31008
box -38 -48 1234 592
use sky130_fd_sc_hd__or2_4  _1182_
timestamp 1608254825
transform 1 0 33764 0 1 31008
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_53_380
timestamp 1608254825
transform 1 0 36064 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_52_372
timestamp 1608254825
transform 1 0 35328 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_490
timestamp 1608254825
transform 1 0 34776 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_4  _1842_
timestamp 1608254825
transform 1 0 36064 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__o21ai_4  _1203_
timestamp 1608254825
transform 1 0 34868 0 1 31008
box -38 -48 1234 592
use sky130_fd_sc_hd__or2_4  _1198_
timestamp 1608254825
transform 1 0 36432 0 1 31008
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_53_391
timestamp 1608254825
transform 1 0 37076 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_396
timestamp 1608254825
transform 1 0 37536 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_392
timestamp 1608254825
transform 1 0 37168 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_484
timestamp 1608254825
transform 1 0 37628 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2571_
timestamp 1608254825
transform 1 0 37444 0 1 31008
box -38 -48 1786 592
use sky130_fd_sc_hd__nand3_4  _1830_
timestamp 1608254825
transform 1 0 37720 0 -1 31008
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_53_414
timestamp 1608254825
transform 1 0 39192 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_52_412
timestamp 1608254825
transform 1 0 39008 0 -1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1608254825
transform -1 0 39836 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1608254825
transform -1 0 39836 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_54_11
timestamp 1608254825
transform 1 0 2116 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_3
timestamp 1608254825
transform 1 0 1380 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1608254825
transform 1 0 1104 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_4  _2063_
timestamp 1608254825
transform 1 0 2208 0 -1 32096
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_12  FILLER_54_36
timestamp 1608254825
transform 1 0 4416 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_25
timestamp 1608254825
transform 1 0 3404 0 -1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_491
timestamp 1608254825
transform 1 0 3956 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _2054_
timestamp 1608254825
transform 1 0 4048 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_66
timestamp 1608254825
transform 1 0 7176 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_54_51
timestamp 1608254825
transform 1 0 5796 0 -1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _2075_
timestamp 1608254825
transform 1 0 5520 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_4  _2038_
timestamp 1608254825
transform 1 0 6348 0 -1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_54_91
timestamp 1608254825
transform 1 0 9476 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_87
timestamp 1608254825
transform 1 0 9108 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__nand4_4  _2037_
timestamp 1608254825
transform 1 0 7544 0 -1 32096
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_54_114
timestamp 1608254825
transform 1 0 11592 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_54_93
timestamp 1608254825
transform 1 0 9660 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_492
timestamp 1608254825
transform 1 0 9568 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2487_
timestamp 1608254825
transform 1 0 9844 0 -1 32096
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_54_121
timestamp 1608254825
transform 1 0 12236 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_4  _1392_
timestamp 1608254825
transform 1 0 12972 0 -1 32096
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _1360_
timestamp 1608254825
transform 1 0 11960 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_54_149
timestamp 1608254825
transform 1 0 14812 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_142
timestamp 1608254825
transform 1 0 14168 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_493
timestamp 1608254825
transform 1 0 15180 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_4  _1389_
timestamp 1608254825
transform 1 0 15272 0 -1 32096
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _1235_
timestamp 1608254825
transform 1 0 14536 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_54_167
timestamp 1608254825
transform 1 0 16468 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_4  _1384_
timestamp 1608254825
transform 1 0 16836 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_196
timestamp 1608254825
transform 1 0 19136 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_183
timestamp 1608254825
transform 1 0 17940 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_4  _1394_
timestamp 1608254825
transform 1 0 19504 0 -1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__and4_4  _1383_
timestamp 1608254825
transform 1 0 18308 0 -1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_54_224
timestamp 1608254825
transform 1 0 21712 0 -1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_213
timestamp 1608254825
transform 1 0 20700 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_209
timestamp 1608254825
transform 1 0 20332 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 21528 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_494
timestamp 1608254825
transform 1 0 20792 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _1893_
timestamp 1608254825
transform 1 0 20884 0 -1 32096
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_54_250
timestamp 1608254825
transform 1 0 24104 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_230
timestamp 1608254825
transform 1 0 22264 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2545_
timestamp 1608254825
transform 1 0 22356 0 -1 32096
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_54_274
timestamp 1608254825
transform 1 0 26312 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_270
timestamp 1608254825
transform 1 0 25944 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_54_258
timestamp 1608254825
transform 1 0 24840 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_4  _1863_
timestamp 1608254825
transform 1 0 25116 0 -1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_54_283
timestamp 1608254825
transform 1 0 27140 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_276
timestamp 1608254825
transform 1 0 26496 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_13_0_addressalyzerBlock.SPI_CLK
timestamp 1608254825
transform 1 0 26864 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_495
timestamp 1608254825
transform 1 0 26404 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2438_
timestamp 1608254825
transform 1 0 27232 0 -1 32096
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_54_303
timestamp 1608254825
transform 1 0 28980 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_4  _1196_
timestamp 1608254825
transform 1 0 29348 0 -1 32096
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_8  FILLER_54_328
timestamp 1608254825
transform 1 0 31280 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_54_320
timestamp 1608254825
transform 1 0 30544 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_496
timestamp 1608254825
transform 1 0 32016 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2649_
timestamp 1608254825
transform 1 0 32108 0 -1 32096
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  _1191_
timestamp 1608254825
transform 1 0 30912 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_362
timestamp 1608254825
transform 1 0 34408 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_54_356
timestamp 1608254825
transform 1 0 33856 0 -1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  _2648_
timestamp 1608254825
transform 1 0 34500 0 -1 32096
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_54_382
timestamp 1608254825
transform 1 0 36248 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1841_
timestamp 1608254825
transform 1 0 36616 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_54_408
timestamp 1608254825
transform 1 0 38640 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_54_402
timestamp 1608254825
transform 1 0 38088 0 -1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_54_389
timestamp 1608254825
transform 1 0 36892 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_497
timestamp 1608254825
transform 1 0 37628 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _2362_
timestamp 1608254825
transform 1 0 38732 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1179_
timestamp 1608254825
transform 1 0 37720 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_417
timestamp 1608254825
transform 1 0 39468 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_413
timestamp 1608254825
transform 1 0 39100 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1608254825
transform -1 0 39836 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_55_18
timestamp 1608254825
transform 1 0 2760 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_55_3
timestamp 1608254825
transform 1 0 1380 0 1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1608254825
transform 1 0 1104 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__and4_4  _2062_
timestamp 1608254825
transform 1 0 1932 0 1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__a41oi_4  _2061_
timestamp 1608254825
transform 1 0 3128 0 1 32096
box -38 -48 2062 592
use sky130_fd_sc_hd__decap_4  FILLER_55_44
timestamp 1608254825
transform 1 0 5152 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_68
timestamp 1608254825
transform 1 0 7360 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_55_62
timestamp 1608254825
transform 1 0 6808 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_55_57
timestamp 1608254825
transform 1 0 6348 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_498
timestamp 1608254825
transform 1 0 6716 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__and3_4  _2044_
timestamp 1608254825
transform 1 0 5520 0 1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1996_
timestamp 1608254825
transform 1 0 7084 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_55_84
timestamp 1608254825
transform 1 0 8832 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_4  _2036_
timestamp 1608254825
transform 1 0 7728 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_114
timestamp 1608254825
transform 1 0 11592 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__a41oi_4  _2033_
timestamp 1608254825
transform 1 0 9568 0 1 32096
box -38 -48 2062 592
use sky130_fd_sc_hd__decap_8  FILLER_55_123
timestamp 1608254825
transform 1 0 12420 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_499
timestamp 1608254825
transform 1 0 12328 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2620_
timestamp 1608254825
transform 1 0 13156 0 1 32096
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_55_150
timestamp 1608254825
transform 1 0 14904 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__nand4_4  _1385_
timestamp 1608254825
transform 1 0 15640 0 1 32096
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_1  FILLER_55_179
timestamp 1608254825
transform 1 0 17572 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_175
timestamp 1608254825
transform 1 0 17204 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_12_0_m1_clk_local
timestamp 1608254825
transform 1 0 17664 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_55_197
timestamp 1608254825
transform 1 0 19228 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_500
timestamp 1608254825
transform 1 0 17940 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__nor3_4  _1395_
timestamp 1608254825
transform 1 0 18032 0 1 32096
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_1  FILLER_55_209
timestamp 1608254825
transform 1 0 20332 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2549_
timestamp 1608254825
transform 1 0 20424 0 1 32096
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_55_240
timestamp 1608254825
transform 1 0 23184 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_229
timestamp 1608254825
transform 1 0 22172 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_501
timestamp 1608254825
transform 1 0 23552 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2544_
timestamp 1608254825
transform 1 0 23644 0 1 32096
box -38 -48 1786 592
use sky130_fd_sc_hd__and2_4  _1897_
timestamp 1608254825
transform 1 0 22540 0 1 32096
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_55_264
timestamp 1608254825
transform 1 0 25392 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2568_
timestamp 1608254825
transform 1 0 25760 0 1 32096
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_55_291
timestamp 1608254825
transform 1 0 27876 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_287
timestamp 1608254825
transform 1 0 27508 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_4  _2192_
timestamp 1608254825
transform 1 0 27968 0 1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_55_319
timestamp 1608254825
transform 1 0 30452 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_55_313
timestamp 1608254825
transform 1 0 29900 0 1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_55_301
timestamp 1608254825
transform 1 0 28796 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_502
timestamp 1608254825
transform 1 0 29164 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _2095_
timestamp 1608254825
transform 1 0 29256 0 1 32096
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_55_339
timestamp 1608254825
transform 1 0 32292 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2650_
timestamp 1608254825
transform 1 0 30544 0 1 32096
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_55_362
timestamp 1608254825
transform 1 0 34408 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_55_347
timestamp 1608254825
transform 1 0 33028 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_55_343
timestamp 1608254825
transform 1 0 32660 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_15_0_addressalyzerBlock.SPI_CLK
timestamp 1608254825
transform 1 0 32752 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_4  _1199_
timestamp 1608254825
transform 1 0 33212 0 1 32096
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_12  FILLER_55_385
timestamp 1608254825
transform 1 0 36524 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_378
timestamp 1608254825
transform 1 0 35880 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_367
timestamp 1608254825
transform 1 0 34868 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_503
timestamp 1608254825
transform 1 0 34776 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _2091_
timestamp 1608254825
transform 1 0 36248 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__or2_4  _1202_
timestamp 1608254825
transform 1 0 35236 0 1 32096
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_55_411
timestamp 1608254825
transform 1 0 38916 0 1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_55_405
timestamp 1608254825
transform 1 0 38364 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_55_397
timestamp 1608254825
transform 1 0 37628 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1829_
timestamp 1608254825
transform 1 0 38640 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_55_417
timestamp 1608254825
transform 1 0 39468 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1608254825
transform -1 0 39836 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_56_22
timestamp 1608254825
transform 1 0 3128 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1608254825
transform 1 0 1104 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _2480_
timestamp 1608254825
transform 1 0 1380 0 -1 33184
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_56_30
timestamp 1608254825
transform 1 0 3864 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_504
timestamp 1608254825
transform 1 0 3956 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__a41oi_4  _2064_
timestamp 1608254825
transform 1 0 4048 0 -1 33184
box -38 -48 2062 592
use sky130_fd_sc_hd__decap_4  FILLER_56_54
timestamp 1608254825
transform 1 0 6072 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2485_
timestamp 1608254825
transform 1 0 6440 0 -1 33184
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_56_85
timestamp 1608254825
transform 1 0 8924 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_77
timestamp 1608254825
transform 1 0 8188 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_m1_clk_local
timestamp 1608254825
transform 1 0 9292 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _2031_
timestamp 1608254825
transform 1 0 8556 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_105
timestamp 1608254825
transform 1 0 10764 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_505
timestamp 1608254825
transform 1 0 9568 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_4  _2034_
timestamp 1608254825
transform 1 0 9660 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__and4_4  _2032_
timestamp 1608254825
transform 1 0 11132 0 -1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_56_130
timestamp 1608254825
transform 1 0 13064 0 -1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_56_118
timestamp 1608254825
transform 1 0 11960 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__nor3_4  _1390_
timestamp 1608254825
transform 1 0 13616 0 -1 33184
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_1  FILLER_56_154
timestamp 1608254825
transform 1 0 15272 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_149
timestamp 1608254825
transform 1 0 14812 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_506
timestamp 1608254825
transform 1 0 15180 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_4  _1386_
timestamp 1608254825
transform 1 0 15364 0 -1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_56_164
timestamp 1608254825
transform 1 0 16192 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2622_
timestamp 1608254825
transform 1 0 16560 0 -1 33184
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_56_187
timestamp 1608254825
transform 1 0 18308 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2619_
timestamp 1608254825
transform 1 0 18676 0 -1 33184
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_56_210
timestamp 1608254825
transform 1 0 20424 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_507
timestamp 1608254825
transform 1 0 20792 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2548_
timestamp 1608254825
transform 1 0 20884 0 -1 33184
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_56_234
timestamp 1608254825
transform 1 0 22632 0 -1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  _2547_
timestamp 1608254825
transform 1 0 23184 0 -1 33184
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_56_274
timestamp 1608254825
transform 1 0 26312 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_270
timestamp 1608254825
transform 1 0 25944 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_259
timestamp 1608254825
transform 1 0 24932 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__and2_4  _1899_
timestamp 1608254825
transform 1 0 25300 0 -1 33184
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_56_282
timestamp 1608254825
transform 1 0 27048 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_56_276
timestamp 1608254825
transform 1 0 26496 0 -1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_508
timestamp 1608254825
transform 1 0 26404 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2465_
timestamp 1608254825
transform 1 0 27140 0 -1 33184
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_56_313
timestamp 1608254825
transform 1 0 29900 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_302
timestamp 1608254825
transform 1 0 28888 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__and2_4  _2094_
timestamp 1608254825
transform 1 0 29256 0 -1 33184
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _1898_
timestamp 1608254825
transform 1 0 30268 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_56_333
timestamp 1608254825
transform 1 0 31740 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_56_321
timestamp 1608254825
transform 1 0 30636 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_509
timestamp 1608254825
transform 1 0 32016 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_4  _1201_
timestamp 1608254825
transform 1 0 32108 0 -1 33184
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_56_361
timestamp 1608254825
transform 1 0 34316 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_350
timestamp 1608254825
transform 1 0 33304 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2467_
timestamp 1608254825
transform 1 0 34684 0 -1 33184
box -38 -48 1786 592
use sky130_fd_sc_hd__or2_4  _1194_
timestamp 1608254825
transform 1 0 33672 0 -1 33184
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_56_384
timestamp 1608254825
transform 1 0 36432 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_398
timestamp 1608254825
transform 1 0 37720 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_396
timestamp 1608254825
transform 1 0 37536 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_510
timestamp 1608254825
transform 1 0 37628 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _2098_
timestamp 1608254825
transform 1 0 38824 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_56_417
timestamp 1608254825
transform 1 0 39468 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_413
timestamp 1608254825
transform 1 0 39100 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1608254825
transform -1 0 39836 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_57_15
timestamp 1608254825
transform 1 0 2484 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_57_3
timestamp 1608254825
transform 1 0 1380 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1608254825
transform 1 0 1104 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__nand4_4  _1993_
timestamp 1608254825
transform 1 0 2760 0 1 33184
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_57_43
timestamp 1608254825
transform 1 0 5060 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_35
timestamp 1608254825
transform 1 0 4324 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _2055_
timestamp 1608254825
transform 1 0 4692 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_57
timestamp 1608254825
transform 1 0 6348 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_47
timestamp 1608254825
transform 1 0 5428 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_511
timestamp 1608254825
transform 1 0 6716 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__nand4_4  _2043_
timestamp 1608254825
transform 1 0 6808 0 1 33184
box -38 -48 1602 592
use sky130_fd_sc_hd__and4_4  _2035_
timestamp 1608254825
transform 1 0 5520 0 1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_57_79
timestamp 1608254825
transform 1 0 8372 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__and3_4  _2028_
timestamp 1608254825
transform 1 0 8740 0 1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_57_113
timestamp 1608254825
transform 1 0 11500 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_57_92
timestamp 1608254825
transform 1 0 9568 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__a41o_4  _2026_
timestamp 1608254825
transform 1 0 9936 0 1 33184
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_1  FILLER_57_129
timestamp 1608254825
transform 1 0 12972 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_57_123
timestamp 1608254825
transform 1 0 12420 0 1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_121
timestamp 1608254825
transform 1 0 12236 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_512
timestamp 1608254825
transform 1 0 12328 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_4  _1393_
timestamp 1608254825
transform 1 0 13064 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_57_148
timestamp 1608254825
transform 1 0 14720 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_57_142
timestamp 1608254825
transform 1 0 14168 0 1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  _2621_
timestamp 1608254825
transform 1 0 14812 0 1 33184
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_57_182
timestamp 1608254825
transform 1 0 17848 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_57_176
timestamp 1608254825
transform 1 0 17296 0 1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_172
timestamp 1608254825
transform 1 0 16928 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_168
timestamp 1608254825
transform 1 0 16560 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1387_
timestamp 1608254825
transform 1 0 17020 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_57_200
timestamp 1608254825
transform 1 0 19504 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_57_196
timestamp 1608254825
transform 1 0 19136 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_184
timestamp 1608254825
transform 1 0 18032 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_m1_clk_local
timestamp 1608254825
transform 1 0 19228 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_513
timestamp 1608254825
transform 1 0 17940 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _1891_
timestamp 1608254825
transform 1 0 19688 0 1 33184
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_57_220
timestamp 1608254825
transform 1 0 21344 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_209
timestamp 1608254825
transform 1 0 20332 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__and2_4  _1896_
timestamp 1608254825
transform 1 0 21712 0 1 33184
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _1894_
timestamp 1608254825
transform 1 0 20700 0 1 33184
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_57_249
timestamp 1608254825
transform 1 0 24012 0 1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_243
timestamp 1608254825
transform 1 0 23460 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_231
timestamp 1608254825
transform 1 0 22356 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_514
timestamp 1608254825
transform 1 0 23552 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1892_
timestamp 1608254825
transform 1 0 23644 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_274
timestamp 1608254825
transform 1 0 26312 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2543_
timestamp 1608254825
transform 1 0 24564 0 1 33184
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _2466_
timestamp 1608254825
transform 1 0 26680 0 1 33184
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_57_297
timestamp 1608254825
transform 1 0 28428 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_515
timestamp 1608254825
transform 1 0 29164 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2384_
timestamp 1608254825
transform 1 0 29256 0 1 33184
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_57_333
timestamp 1608254825
transform 1 0 31740 0 1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_57_325
timestamp 1608254825
transform 1 0 31004 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2457_
timestamp 1608254825
transform 1 0 32292 0 1 33184
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  _2096_
timestamp 1608254825
transform 1 0 31372 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_57_358
timestamp 1608254825
transform 1 0 34040 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_57_386
timestamp 1608254825
transform 1 0 36616 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_516
timestamp 1608254825
transform 1 0 34776 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2455_
timestamp 1608254825
transform 1 0 34868 0 1 33184
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_57_410
timestamp 1608254825
transform 1 0 38824 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_57_398
timestamp 1608254825
transform 1 0 37720 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1608254825
transform -1 0 39836 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_58_9
timestamp 1608254825
transform 1 0 1932 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_58_3
timestamp 1608254825
transform 1 0 1380 0 -1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1608254825
transform 1 0 1104 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__a41o_4  _2056_
timestamp 1608254825
transform 1 0 2024 0 -1 34272
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_58_44
timestamp 1608254825
transform 1 0 5152 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_27
timestamp 1608254825
transform 1 0 3588 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_517
timestamp 1608254825
transform 1 0 3956 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_4  _2065_
timestamp 1608254825
transform 1 0 4048 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_48
timestamp 1608254825
transform 1 0 5520 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_10_0_m1_clk_local
timestamp 1608254825
transform 1 0 5612 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__a41o_4  _2042_
timestamp 1608254825
transform 1 0 5888 0 -1 34272
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_58_88
timestamp 1608254825
transform 1 0 9200 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_58_69
timestamp 1608254825
transform 1 0 7452 0 -1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_4  _2046_
timestamp 1608254825
transform 1 0 8004 0 -1 34272
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_58_103
timestamp 1608254825
transform 1 0 10580 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_93
timestamp 1608254825
transform 1 0 9660 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_518
timestamp 1608254825
transform 1 0 9568 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2488_
timestamp 1608254825
transform 1 0 10948 0 -1 34272
box -38 -48 1786 592
use sky130_fd_sc_hd__and4_4  _2017_
timestamp 1608254825
transform 1 0 9752 0 -1 34272
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_58_126
timestamp 1608254825
transform 1 0 12696 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_4  _2019_
timestamp 1608254825
transform 1 0 13064 0 -1 34272
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_12  FILLER_58_154
timestamp 1608254825
transform 1 0 15272 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_58_151
timestamp 1608254825
transform 1 0 14996 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_58_143
timestamp 1608254825
transform 1 0 14260 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_519
timestamp 1608254825
transform 1 0 15180 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_58_166
timestamp 1608254825
transform 1 0 16376 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _2554_
timestamp 1608254825
transform 1 0 16560 0 -1 34272
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_58_187
timestamp 1608254825
transform 1 0 18308 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2553_
timestamp 1608254825
transform 1 0 18676 0 -1 34272
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_58_223
timestamp 1608254825
transform 1 0 21620 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_215
timestamp 1608254825
transform 1 0 20884 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_58_210
timestamp 1608254825
transform 1 0 20424 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_m1_clk_local
timestamp 1608254825
transform 1 0 21712 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_520
timestamp 1608254825
transform 1 0 20792 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2546_
timestamp 1608254825
transform 1 0 21988 0 -1 34272
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_58_246
timestamp 1608254825
transform 1 0 23736 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__and2_4  _1895_
timestamp 1608254825
transform 1 0 24104 0 -1 34272
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_58_274
timestamp 1608254825
transform 1 0 26312 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_58_268
timestamp 1608254825
transform 1 0 25760 0 -1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_58_257
timestamp 1608254825
transform 1 0 24748 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__and2_4  _1900_
timestamp 1608254825
transform 1 0 25116 0 -1 34272
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_58_285
timestamp 1608254825
transform 1 0 27324 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_521
timestamp 1608254825
transform 1 0 26404 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__and3_4  _1980_
timestamp 1608254825
transform 1 0 27692 0 -1 34272
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  _1866_
timestamp 1608254825
transform 1 0 26496 0 -1 34272
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_58_309
timestamp 1608254825
transform 1 0 29532 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_298
timestamp 1608254825
transform 1 0 28520 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2464_
timestamp 1608254825
transform 1 0 29900 0 -1 34272
box -38 -48 1786 592
use sky130_fd_sc_hd__or2_4  _1979_
timestamp 1608254825
transform 1 0 28888 0 -1 34272
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_58_332
timestamp 1608254825
transform 1 0 31648 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_522
timestamp 1608254825
transform 1 0 32016 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _2097_
timestamp 1608254825
transform 1 0 32108 0 -1 34272
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_58_344
timestamp 1608254825
transform 1 0 32752 0 -1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  _2454_
timestamp 1608254825
transform 1 0 33304 0 -1 34272
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_58_380
timestamp 1608254825
transform 1 0 36064 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_369
timestamp 1608254825
transform 1 0 35052 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__and2_4  _2110_
timestamp 1608254825
transform 1 0 35420 0 -1 34272
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_58_410
timestamp 1608254825
transform 1 0 38824 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_58_398
timestamp 1608254825
transform 1 0 37720 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_396
timestamp 1608254825
transform 1 0 37536 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_392
timestamp 1608254825
transform 1 0 37168 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_523
timestamp 1608254825
transform 1 0 37628 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1608254825
transform -1 0 39836 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_60_22
timestamp 1608254825
transform 1 0 3128 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_59_15
timestamp 1608254825
transform 1 0 2484 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_59_3
timestamp 1608254825
transform 1 0 1380 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1608254825
transform 1 0 1104 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1608254825
transform 1 0 1104 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _2481_
timestamp 1608254825
transform 1 0 1380 0 -1 35360
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _2479_
timestamp 1608254825
transform 1 0 2852 0 1 34272
box -38 -48 1786 592
use sky130_fd_sc_hd__and3_4  _2057_
timestamp 1608254825
transform 1 0 1656 0 1 34272
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_60_35
timestamp 1608254825
transform 1 0 4324 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_30
timestamp 1608254825
transform 1 0 3864 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_38
timestamp 1608254825
transform 1 0 4600 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_530
timestamp 1608254825
transform 1 0 3956 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2482_
timestamp 1608254825
transform 1 0 4692 0 -1 35360
box -38 -48 1786 592
use sky130_fd_sc_hd__o21ai_4  _2051_
timestamp 1608254825
transform 1 0 4968 0 1 34272
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _2041_
timestamp 1608254825
transform 1 0 4048 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_60_58
timestamp 1608254825
transform 1 0 6440 0 -1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_62
timestamp 1608254825
transform 1 0 6808 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_59_55
timestamp 1608254825
transform 1 0 6164 0 1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_524
timestamp 1608254825
transform 1 0 6716 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _2029_
timestamp 1608254825
transform 1 0 6900 0 1 34272
box -38 -48 866 592
use sky130_fd_sc_hd__nor4_4  _1994_
timestamp 1608254825
transform 1 0 6992 0 -1 35360
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_60_88
timestamp 1608254825
transform 1 0 9200 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_81
timestamp 1608254825
transform 1 0 8556 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_90
timestamp 1608254825
transform 1 0 9384 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_76
timestamp 1608254825
transform 1 0 8096 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_72
timestamp 1608254825
transform 1 0 7728 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_4  _2045_
timestamp 1608254825
transform 1 0 8188 0 1 34272
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _1985_
timestamp 1608254825
transform 1 0 8924 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_60_110
timestamp 1608254825
transform 1 0 11224 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_93
timestamp 1608254825
transform 1 0 9660 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_59_114
timestamp 1608254825
transform 1 0 11592 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_11_0_m1_clk_local
timestamp 1608254825
transform 1 0 9752 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_531
timestamp 1608254825
transform 1 0 9568 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_4  _2024_
timestamp 1608254825
transform 1 0 10028 0 -1 35360
box -38 -48 1234 592
use sky130_fd_sc_hd__buf_2  _2012_
timestamp 1608254825
transform 1 0 11592 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__nand4_4  _1997_
timestamp 1608254825
transform 1 0 10028 0 1 34272
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_1  FILLER_60_126
timestamp 1608254825
transform 1 0 12696 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_60_118
timestamp 1608254825
transform 1 0 11960 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_525
timestamp 1608254825
transform 1 0 12328 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2489_
timestamp 1608254825
transform 1 0 12788 0 -1 35360
box -38 -48 1786 592
use sky130_fd_sc_hd__a41oi_4  _2018_
timestamp 1608254825
transform 1 0 12420 0 1 34272
box -38 -48 2062 592
use sky130_fd_sc_hd__fill_1  FILLER_60_152
timestamp 1608254825
transform 1 0 15088 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_60_146
timestamp 1608254825
transform 1 0 14536 0 -1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_59_145
timestamp 1608254825
transform 1 0 14444 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_532
timestamp 1608254825
transform 1 0 15180 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2562_
timestamp 1608254825
transform 1 0 15272 0 -1 35360
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _2491_
timestamp 1608254825
transform 1 0 14812 0 1 34272
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_60_173
timestamp 1608254825
transform 1 0 17020 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_59_179
timestamp 1608254825
transform 1 0 17572 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_168
timestamp 1608254825
transform 1 0 16560 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2561_
timestamp 1608254825
transform 1 0 17756 0 -1 35360
box -38 -48 1786 592
use sky130_fd_sc_hd__and2_4  _1887_
timestamp 1608254825
transform 1 0 16928 0 1 34272
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_60_200
timestamp 1608254825
transform 1 0 19504 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_200
timestamp 1608254825
transform 1 0 19504 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_192
timestamp 1608254825
transform 1 0 18768 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_184
timestamp 1608254825
transform 1 0 18032 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_526
timestamp 1608254825
transform 1 0 17940 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2550_
timestamp 1608254825
transform 1 0 19872 0 1 34272
box -38 -48 1786 592
use sky130_fd_sc_hd__and2_4  _1888_
timestamp 1608254825
transform 1 0 18860 0 1 34272
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_60_221
timestamp 1608254825
transform 1 0 21436 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_60_215
timestamp 1608254825
transform 1 0 20884 0 -1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_60_212
timestamp 1608254825
transform 1 0 20608 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_223
timestamp 1608254825
transform 1 0 21620 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_533
timestamp 1608254825
transform 1 0 20792 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_4  _2347_
timestamp 1608254825
transform 1 0 21528 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_4  _2346_
timestamp 1608254825
transform 1 0 21988 0 1 34272
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_60_238
timestamp 1608254825
transform 1 0 23000 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_234
timestamp 1608254825
transform 1 0 22632 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_236
timestamp 1608254825
transform 1 0 22816 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__or3_4  _1981_
timestamp 1608254825
transform 1 0 23092 0 -1 35360
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_60_248
timestamp 1608254825
transform 1 0 23920 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_59_245
timestamp 1608254825
transform 1 0 23644 0 1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_240
timestamp 1608254825
transform 1 0 23184 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_m1_clk_local
timestamp 1608254825
transform 1 0 23276 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_527
timestamp 1608254825
transform 1 0 23552 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2495_
timestamp 1608254825
transform 1 0 24196 0 1 34272
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_60_268
timestamp 1608254825
transform 1 0 25760 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_261
timestamp 1608254825
transform 1 0 25116 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_59_270
timestamp 1608254825
transform 1 0 25944 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_15_0_m1_clk_local
timestamp 1608254825
transform 1 0 26128 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1982_
timestamp 1608254825
transform 1 0 25484 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_4  _1976_
timestamp 1608254825
transform 1 0 24288 0 -1 35360
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_60_290
timestamp 1608254825
transform 1 0 27784 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_59_278
timestamp 1608254825
transform 1 0 26680 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_534
timestamp 1608254825
transform 1 0 26404 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2496_
timestamp 1608254825
transform 1 0 26772 0 1 34272
box -38 -48 1786 592
use sky130_fd_sc_hd__nand3_4  _1972_
timestamp 1608254825
transform 1 0 26496 0 -1 35360
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_60_318
timestamp 1608254825
transform 1 0 30360 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_298
timestamp 1608254825
transform 1 0 28520 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_59_304
timestamp 1608254825
transform 1 0 29072 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_59_298
timestamp 1608254825
transform 1 0 28520 0 1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_528
timestamp 1608254825
transform 1 0 29164 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2383_
timestamp 1608254825
transform 1 0 29256 0 1 34272
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _2381_
timestamp 1608254825
transform 1 0 28612 0 -1 35360
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_60_337
timestamp 1608254825
transform 1 0 32108 0 -1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_335
timestamp 1608254825
transform 1 0 31924 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_60_329
timestamp 1608254825
transform 1 0 31372 0 -1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_59_325
timestamp 1608254825
transform 1 0 31004 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_535
timestamp 1608254825
transform 1 0 32016 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2456_
timestamp 1608254825
transform 1 0 31372 0 1 34272
box -38 -48 1786 592
use sky130_fd_sc_hd__and2_4  _2108_
timestamp 1608254825
transform 1 0 30728 0 -1 35360
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_60_363
timestamp 1608254825
transform 1 0 34500 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_343
timestamp 1608254825
transform 1 0 32660 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_59_365
timestamp 1608254825
transform 1 0 34684 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_361
timestamp 1608254825
transform 1 0 34316 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_59_348
timestamp 1608254825
transform 1 0 33120 0 1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  _2379_
timestamp 1608254825
transform 1 0 32752 0 -1 35360
box -38 -48 1786 592
use sky130_fd_sc_hd__and2_4  _2093_
timestamp 1608254825
transform 1 0 33672 0 1 34272
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_60_387
timestamp 1608254825
transform 1 0 36708 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_60_375
timestamp 1608254825
transform 1 0 35604 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_386
timestamp 1608254825
transform 1 0 36616 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_374
timestamp 1608254825
transform 1 0 35512 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_529
timestamp 1608254825
transform 1 0 34776 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _2109_
timestamp 1608254825
transform 1 0 34868 0 1 34272
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_60_410
timestamp 1608254825
transform 1 0 38824 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_60_398
timestamp 1608254825
transform 1 0 37720 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_60_395
timestamp 1608254825
transform 1 0 37444 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_59_410
timestamp 1608254825
transform 1 0 38824 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_59_398
timestamp 1608254825
transform 1 0 37720 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_536
timestamp 1608254825
transform 1 0 37628 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1608254825
transform -1 0 39836 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1608254825
transform -1 0 39836 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_61_11
timestamp 1608254825
transform 1 0 2116 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_3
timestamp 1608254825
transform 1 0 1380 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1608254825
transform 1 0 1104 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _2359_
timestamp 1608254825
transform 1 0 1748 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_41
timestamp 1608254825
transform 1 0 4876 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_33
timestamp 1608254825
transform 1 0 4140 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_61_23
timestamp 1608254825
transform 1 0 3220 0 1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_4  _2048_
timestamp 1608254825
transform 1 0 4968 0 1 35360
box -38 -48 1234 592
use sky130_fd_sc_hd__buf_2  _2040_
timestamp 1608254825
transform 1 0 3772 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_61_66
timestamp 1608254825
transform 1 0 7176 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_61_55
timestamp 1608254825
transform 1 0 6164 0 1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_537
timestamp 1608254825
transform 1 0 6716 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _2014_
timestamp 1608254825
transform 1 0 6808 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_74
timestamp 1608254825
transform 1 0 7912 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2484_
timestamp 1608254825
transform 1 0 8004 0 1 35360
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_61_113
timestamp 1608254825
transform 1 0 11500 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_61_94
timestamp 1608254825
transform 1 0 9752 0 1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_4  _2004_
timestamp 1608254825
transform 1 0 10304 0 1 35360
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_6  FILLER_61_136
timestamp 1608254825
transform 1 0 13616 0 1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_121
timestamp 1608254825
transform 1 0 12236 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_538
timestamp 1608254825
transform 1 0 12328 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_4  _2025_
timestamp 1608254825
transform 1 0 12420 0 1 35360
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_61_150
timestamp 1608254825
transform 1 0 14904 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_142
timestamp 1608254825
transform 1 0 14168 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2382_
timestamp 1608254825
transform 1 0 15272 0 1 35360
box -38 -48 1786 592
use sky130_fd_sc_hd__and2_4  _1877_
timestamp 1608254825
transform 1 0 14260 0 1 35360
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_61_181
timestamp 1608254825
transform 1 0 17756 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_61_173
timestamp 1608254825
transform 1 0 17020 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_61_198
timestamp 1608254825
transform 1 0 19320 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_191
timestamp 1608254825
transform 1 0 18676 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_13_0_m1_clk_local
timestamp 1608254825
transform 1 0 19044 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_539
timestamp 1608254825
transform 1 0 17940 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _1878_
timestamp 1608254825
transform 1 0 18032 0 1 35360
box -38 -48 682 592
use sky130_fd_sc_hd__nor3_4  _1865_
timestamp 1608254825
transform 1 0 19688 0 1 35360
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_61_215
timestamp 1608254825
transform 1 0 20884 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2567_
timestamp 1608254825
transform 1 0 21252 0 1 35360
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_61_238
timestamp 1608254825
transform 1 0 23000 0 1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_540
timestamp 1608254825
transform 1 0 23552 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__nor3_4  _1975_
timestamp 1608254825
transform 1 0 23644 0 1 35360
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_1  FILLER_61_262
timestamp 1608254825
transform 1 0 25208 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_258
timestamp 1608254825
transform 1 0 24840 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_4  _1867_
timestamp 1608254825
transform 1 0 25300 0 1 35360
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_12  FILLER_61_292
timestamp 1608254825
transform 1 0 27968 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_276
timestamp 1608254825
transform 1 0 26496 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_4  _1977_
timestamp 1608254825
transform 1 0 26864 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_315
timestamp 1608254825
transform 1 0 30084 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_304
timestamp 1608254825
transform 1 0 29072 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_541
timestamp 1608254825
transform 1 0 29164 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__and3_4  _1978_
timestamp 1608254825
transform 1 0 29256 0 1 35360
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_61_342
timestamp 1608254825
transform 1 0 32568 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2377_
timestamp 1608254825
transform 1 0 30820 0 1 35360
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_61_365
timestamp 1608254825
transform 1 0 34684 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_353
timestamp 1608254825
transform 1 0 33580 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__and2_4  _2107_
timestamp 1608254825
transform 1 0 32936 0 1 35360
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_61_379
timestamp 1608254825
transform 1 0 35972 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_367
timestamp 1608254825
transform 1 0 34868 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_542
timestamp 1608254825
transform 1 0 34776 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_403
timestamp 1608254825
transform 1 0 38180 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_391
timestamp 1608254825
transform 1 0 37076 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_61_415
timestamp 1608254825
transform 1 0 39284 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1608254825
transform -1 0 39836 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_62_15
timestamp 1608254825
transform 1 0 2484 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_3
timestamp 1608254825
transform 1 0 1380 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1608254825
transform 1 0 1104 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_62_32
timestamp 1608254825
transform 1 0 4048 0 -1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_62_27
timestamp 1608254825
transform 1 0 3588 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_543
timestamp 1608254825
transform 1 0 3956 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_4  _2052_
timestamp 1608254825
transform 1 0 4600 0 -1 36448
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_8  FILLER_62_51
timestamp 1608254825
transform 1 0 5796 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__nor3_4  _2015_
timestamp 1608254825
transform 1 0 6532 0 -1 36448
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_62_88
timestamp 1608254825
transform 1 0 9200 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 1608254825
transform 1 0 8740 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_79
timestamp 1608254825
transform 1 0 8372 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_72
timestamp 1608254825
transform 1 0 7728 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _2016_
timestamp 1608254825
transform 1 0 8832 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1986_
timestamp 1608254825
transform 1 0 8096 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_62_107
timestamp 1608254825
transform 1 0 10948 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_93
timestamp 1608254825
transform 1 0 9660 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_544
timestamp 1608254825
transform 1 0 9568 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_4  _2021_
timestamp 1608254825
transform 1 0 9752 0 -1 36448
box -38 -48 1234 592
use sky130_fd_sc_hd__nor4_4  _2013_
timestamp 1608254825
transform 1 0 11316 0 -1 36448
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_6  FILLER_62_128
timestamp 1608254825
transform 1 0 12880 0 -1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_4  _1998_
timestamp 1608254825
transform 1 0 13432 0 -1 36448
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_62_157
timestamp 1608254825
transform 1 0 15548 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_62_151
timestamp 1608254825
transform 1 0 14996 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_62_143
timestamp 1608254825
transform 1 0 14260 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_545
timestamp 1608254825
transform 1 0 15180 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1984_
timestamp 1608254825
transform 1 0 15272 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_62_165
timestamp 1608254825
transform 1 0 16284 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2363_
timestamp 1608254825
transform 1 0 16376 0 -1 36448
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_62_185
timestamp 1608254825
transform 1 0 18124 0 -1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  _2365_
timestamp 1608254825
transform 1 0 18676 0 -1 36448
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_62_218
timestamp 1608254825
transform 1 0 21160 0 -1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_62_210
timestamp 1608254825
transform 1 0 20424 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_546
timestamp 1608254825
transform 1 0 20792 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__xnor2_4  _1868_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 21712 0 -1 36448
box -38 -48 2062 592
use sky130_fd_sc_hd__inv_2  _1864_
timestamp 1608254825
transform 1 0 20884 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_62_246
timestamp 1608254825
transform 1 0 23736 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2498_
timestamp 1608254825
transform 1 0 24104 0 -1 36448
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_62_269
timestamp 1608254825
transform 1 0 25852 0 -1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_284
timestamp 1608254825
transform 1 0 27232 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_276
timestamp 1608254825
transform 1 0 26496 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_547
timestamp 1608254825
transform 1 0 26404 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2497_
timestamp 1608254825
transform 1 0 27324 0 -1 36448
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_62_310
timestamp 1608254825
transform 1 0 29624 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_62_304
timestamp 1608254825
transform 1 0 29072 0 -1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  _2376_
timestamp 1608254825
transform 1 0 29716 0 -1 36448
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_62_330
timestamp 1608254825
transform 1 0 31464 0 -1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_548
timestamp 1608254825
transform 1 0 32016 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2378_
timestamp 1608254825
transform 1 0 32108 0 -1 36448
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_62_356
timestamp 1608254825
transform 1 0 33856 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2380_
timestamp 1608254825
transform 1 0 34224 0 -1 36448
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_62_379
timestamp 1608254825
transform 1 0 35972 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_410
timestamp 1608254825
transform 1 0 38824 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_62_398
timestamp 1608254825
transform 1 0 37720 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_391
timestamp 1608254825
transform 1 0 37076 0 -1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_549
timestamp 1608254825
transform 1 0 37628 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1608254825
transform -1 0 39836 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_63_15
timestamp 1608254825
transform 1 0 2484 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_3
timestamp 1608254825
transform 1 0 1380 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1608254825
transform 1 0 1104 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_63_39
timestamp 1608254825
transform 1 0 4692 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_63_27
timestamp 1608254825
transform 1 0 3588 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__nand3_4  _2049_
timestamp 1608254825
transform 1 0 5060 0 1 36448
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_63_62
timestamp 1608254825
transform 1 0 6808 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_57
timestamp 1608254825
transform 1 0 6348 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_550
timestamp 1608254825
transform 1 0 6716 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _2030_
timestamp 1608254825
transform 1 0 7176 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_90
timestamp 1608254825
transform 1 0 9384 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_77
timestamp 1608254825
transform 1 0 8188 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_70
timestamp 1608254825
transform 1 0 7544 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_4  _2001_
timestamp 1608254825
transform 1 0 8556 0 1 36448
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1987_
timestamp 1608254825
transform 1 0 7912 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_63_114
timestamp 1608254825
transform 1 0 11592 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_63_108
timestamp 1608254825
transform 1 0 11040 0 1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_4  _2022_
timestamp 1608254825
transform 1 0 9752 0 1 36448
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_63_130
timestamp 1608254825
transform 1 0 13064 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_63_123
timestamp 1608254825
transform 1 0 12420 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_63_118
timestamp 1608254825
transform 1 0 11960 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_551
timestamp 1608254825
transform 1 0 12328 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__a41o_4  _2009_
timestamp 1608254825
transform 1 0 13432 0 1 36448
box -38 -48 1602 592
use sky130_fd_sc_hd__inv_2  _2003_
timestamp 1608254825
transform 1 0 11684 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _2002_
timestamp 1608254825
transform 1 0 12696 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_151
timestamp 1608254825
transform 1 0 14996 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__and3_4  _2010_
timestamp 1608254825
transform 1 0 15364 0 1 36448
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_63_182
timestamp 1608254825
transform 1 0 17848 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_63_176
timestamp 1608254825
transform 1 0 17296 0 1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_63_164
timestamp 1608254825
transform 1 0 16192 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_203
timestamp 1608254825
transform 1 0 19780 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_552
timestamp 1608254825
transform 1 0 17940 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2364_
timestamp 1608254825
transform 1 0 18032 0 1 36448
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_63_226
timestamp 1608254825
transform 1 0 21896 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2366_
timestamp 1608254825
transform 1 0 20148 0 1 36448
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_63_245
timestamp 1608254825
transform 1 0 23644 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_243
timestamp 1608254825
transform 1 0 23460 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_239
timestamp 1608254825
transform 1 0 23092 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_553
timestamp 1608254825
transform 1 0 23552 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _1869_
timestamp 1608254825
transform 1 0 22264 0 1 36448
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_63_274
timestamp 1608254825
transform 1 0 26312 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_63_258
timestamp 1608254825
transform 1 0 24840 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_63_253
timestamp 1608254825
transform 1 0 24380 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_14_0_m1_clk_local
timestamp 1608254825
transform 1 0 24564 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_4  _1974_
timestamp 1608254825
transform 1 0 25116 0 1 36448
box -38 -48 1234 592
use sky130_fd_sc_hd__dfxtp_4  _2373_
timestamp 1608254825
transform 1 0 27048 0 1 36448
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_63_301
timestamp 1608254825
transform 1 0 28796 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_554
timestamp 1608254825
transform 1 0 29164 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2375_
timestamp 1608254825
transform 1 0 29256 0 1 36448
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_63_332
timestamp 1608254825
transform 1 0 31648 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_325
timestamp 1608254825
transform 1 0 31004 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2348_
timestamp 1608254825
transform 1 0 31372 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_63_364
timestamp 1608254825
transform 1 0 34592 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_63_356
timestamp 1608254825
transform 1 0 33856 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_63_344
timestamp 1608254825
transform 1 0 32752 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_379
timestamp 1608254825
transform 1 0 35972 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_367
timestamp 1608254825
transform 1 0 34868 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_555
timestamp 1608254825
transform 1 0 34776 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_403
timestamp 1608254825
transform 1 0 38180 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_391
timestamp 1608254825
transform 1 0 37076 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_63_415
timestamp 1608254825
transform 1 0 39284 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1608254825
transform -1 0 39836 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_11
timestamp 1608254825
transform 1 0 2116 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_64_3
timestamp 1608254825
transform 1 0 1380 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_1
timestamp 1608254825
transform 1 0 1564 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1608254825
transform 1 0 1104 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _2361_
timestamp 1608254825
transform 1 0 1748 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_45
timestamp 1608254825
transform 1 0 5244 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_40
timestamp 1608254825
transform 1 0 4784 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_32
timestamp 1608254825
transform 1 0 4048 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_64_23
timestamp 1608254825
transform 1 0 3220 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_556
timestamp 1608254825
transform 1 0 3956 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _2050_
timestamp 1608254825
transform 1 0 4968 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_64_68
timestamp 1608254825
transform 1 0 7360 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  _2483_
timestamp 1608254825
transform 1 0 5612 0 -1 37536
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_64_88
timestamp 1608254825
transform 1 0 9200 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_4  _2006_
timestamp 1608254825
transform 1 0 7912 0 -1 37536
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_1  FILLER_64_104
timestamp 1608254825
transform 1 0 10672 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_96
timestamp 1608254825
transform 1 0 9936 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_557
timestamp 1608254825
transform 1 0 9568 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2490_
timestamp 1608254825
transform 1 0 10764 0 -1 37536
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_2  _2000_
timestamp 1608254825
transform 1 0 9660 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_64_124
timestamp 1608254825
transform 1 0 12512 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__nand4_4  _1999_
timestamp 1608254825
transform 1 0 13064 0 -1 37536
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_64_157
timestamp 1608254825
transform 1 0 15548 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_147
timestamp 1608254825
transform 1 0 14628 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_558
timestamp 1608254825
transform 1 0 15180 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _2008_
timestamp 1608254825
transform 1 0 15272 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_64_172
timestamp 1608254825
transform 1 0 16928 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_64_164
timestamp 1608254825
transform 1 0 16192 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _2534_
timestamp 1608254825
transform 1 0 17204 0 -1 37536
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_2  _2341_
timestamp 1608254825
transform 1 0 15916 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_194
timestamp 1608254825
transform 1 0 18952 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_206
timestamp 1608254825
transform 1 0 20056 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_559
timestamp 1608254825
transform 1 0 20792 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2367_
timestamp 1608254825
transform 1 0 20884 0 -1 37536
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_64_234
timestamp 1608254825
transform 1 0 22632 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2369_
timestamp 1608254825
transform 1 0 23000 0 -1 37536
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_64_271
timestamp 1608254825
transform 1 0 26036 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_261
timestamp 1608254825
transform 1 0 25116 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_257
timestamp 1608254825
transform 1 0 24748 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_4  _1973_
timestamp 1608254825
transform 1 0 25208 0 -1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_64_295
timestamp 1608254825
transform 1 0 28244 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_560
timestamp 1608254825
transform 1 0 26404 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2372_
timestamp 1608254825
transform 1 0 26496 0 -1 37536
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_64_318
timestamp 1608254825
transform 1 0 30360 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _2374_
timestamp 1608254825
transform 1 0 28612 0 -1 37536
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_64_337
timestamp 1608254825
transform 1 0 32108 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_330
timestamp 1608254825
transform 1 0 31464 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_561
timestamp 1608254825
transform 1 0 32016 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_349
timestamp 1608254825
transform 1 0 33212 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_2
timestamp 1608254825
transform 1 0 33396 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _2501_
timestamp 1608254825
transform 1 0 33580 0 -1 37536
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_64_384
timestamp 1608254825
transform 1 0 36432 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_372
timestamp 1608254825
transform 1 0 35328 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_410
timestamp 1608254825
transform 1 0 38824 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_64_398
timestamp 1608254825
transform 1 0 37720 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_396
timestamp 1608254825
transform 1 0 37536 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_562
timestamp 1608254825
transform 1 0 37628 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1608254825
transform -1 0 39836 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_65_15
timestamp 1608254825
transform 1 0 2484 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_3
timestamp 1608254825
transform 1 0 1380 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1608254825
transform 1 0 1104 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_65_35
timestamp 1608254825
transform 1 0 4324 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_65_27
timestamp 1608254825
transform 1 0 3588 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _2499_
timestamp 1608254825
transform 1 0 4600 0 1 37536
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_65_65
timestamp 1608254825
transform 1 0 7084 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_65_57
timestamp 1608254825
transform 1 0 6348 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_563
timestamp 1608254825
transform 1 0 6716 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _2047_
timestamp 1608254825
transform 1 0 6808 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _2493_
timestamp 1608254825
transform 1 0 7820 0 1 37536
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_65_113
timestamp 1608254825
transform 1 0 11500 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_65_92
timestamp 1608254825
transform 1 0 9568 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__nand4_4  _2005_
timestamp 1608254825
transform 1 0 9936 0 1 37536
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_1  FILLER_65_121
timestamp 1608254825
transform 1 0 12236 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_564
timestamp 1608254825
transform 1 0 12328 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2470_
timestamp 1608254825
transform 1 0 12420 0 1 37536
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_65_142
timestamp 1608254825
transform 1 0 14168 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2492_
timestamp 1608254825
transform 1 0 14536 0 1 37536
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_65_177
timestamp 1608254825
transform 1 0 17388 0 1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_65_165
timestamp 1608254825
transform 1 0 16284 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_65_192
timestamp 1608254825
transform 1 0 18768 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_65_184
timestamp 1608254825
transform 1 0 18032 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_3
timestamp 1608254825
transform 1 0 19044 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_565
timestamp 1608254825
transform 1 0 17940 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2532_
timestamp 1608254825
transform 1 0 19228 0 1 37536
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_65_220
timestamp 1608254825
transform 1 0 21344 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_216
timestamp 1608254825
transform 1 0 20976 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2368_
timestamp 1608254825
transform 1 0 21436 0 1 37536
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  FILLER_65_245
timestamp 1608254825
transform 1 0 23644 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_65_240
timestamp 1608254825
transform 1 0 23184 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_566
timestamp 1608254825
transform 1 0 23552 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2370_
timestamp 1608254825
transform 1 0 23920 0 1 37536
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_65_267
timestamp 1608254825
transform 1 0 25668 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2371_
timestamp 1608254825
transform 1 0 26036 0 1 37536
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_65_290
timestamp 1608254825
transform 1 0 27784 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_65_310
timestamp 1608254825
transform 1 0 29624 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_306
timestamp 1608254825
transform 1 0 29256 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_65_302
timestamp 1608254825
transform 1 0 28888 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_567
timestamp 1608254825
transform 1 0 29164 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_4  _2350_
timestamp 1608254825
transform 1 0 29716 0 1 37536
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_12  FILLER_65_336
timestamp 1608254825
transform 1 0 32016 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_324
timestamp 1608254825
transform 1 0 30912 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_360
timestamp 1608254825
transform 1 0 34224 0 1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_65_348
timestamp 1608254825
transform 1 0 33120 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_386
timestamp 1608254825
transform 1 0 36616 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_568
timestamp 1608254825
transform 1 0 34776 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2508_
timestamp 1608254825
transform 1 0 34868 0 1 37536
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_65_410
timestamp 1608254825
transform 1 0 38824 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_65_398
timestamp 1608254825
transform 1 0 37720 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1608254825
transform -1 0 39836 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_66_15
timestamp 1608254825
transform 1 0 2484 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_3
timestamp 1608254825
transform 1 0 1380 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1608254825
transform 1 0 1104 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_66_44
timestamp 1608254825
transform 1 0 5152 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_32
timestamp 1608254825
transform 1 0 4048 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_66_27
timestamp 1608254825
transform 1 0 3588 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_569
timestamp 1608254825
transform 1 0 3956 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_66_56
timestamp 1608254825
transform 1 0 6256 0 -1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_570
timestamp 1608254825
transform 1 0 6808 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2511_
timestamp 1608254825
transform 1 0 6900 0 -1 38624
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_66_89
timestamp 1608254825
transform 1 0 9292 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_82
timestamp 1608254825
transform 1 0 8648 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2007_
timestamp 1608254825
transform 1 0 9016 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_66_114
timestamp 1608254825
transform 1 0 11592 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_66_107
timestamp 1608254825
transform 1 0 10948 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_66_102
timestamp 1608254825
transform 1 0 10488 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_66_94
timestamp 1608254825
transform 1 0 9752 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_571
timestamp 1608254825
transform 1 0 9660 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _2023_
timestamp 1608254825
transform 1 0 11316 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2020_
timestamp 1608254825
transform 1 0 10672 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_66_128
timestamp 1608254825
transform 1 0 12880 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_66_122
timestamp 1608254825
transform 1 0 12328 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_572
timestamp 1608254825
transform 1 0 12512 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _2011_
timestamp 1608254825
transform 1 0 12604 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_66_156
timestamp 1608254825
transform 1 0 15456 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_66_152
timestamp 1608254825
transform 1 0 15088 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_66_140
timestamp 1608254825
transform 1 0 13984 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_573
timestamp 1608254825
transform 1 0 15364 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_66_180
timestamp 1608254825
transform 1 0 17664 0 -1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_66_168
timestamp 1608254825
transform 1 0 16560 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_199
timestamp 1608254825
transform 1 0 19412 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_187
timestamp 1608254825
transform 1 0 18308 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_574
timestamp 1608254825
transform 1 0 18216 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_218
timestamp 1608254825
transform 1 0 21160 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_211
timestamp 1608254825
transform 1 0 20516 0 -1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_575
timestamp 1608254825
transform 1 0 21068 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_249
timestamp 1608254825
transform 1 0 24012 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_242
timestamp 1608254825
transform 1 0 23368 0 -1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_66_230
timestamp 1608254825
transform 1 0 22264 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_576
timestamp 1608254825
transform 1 0 23920 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_66_273
timestamp 1608254825
transform 1 0 26220 0 -1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_66_261
timestamp 1608254825
transform 1 0 25116 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_292
timestamp 1608254825
transform 1 0 27968 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_280
timestamp 1608254825
transform 1 0 26864 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_577
timestamp 1608254825
transform 1 0 26772 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_66_304
timestamp 1608254825
transform 1 0 29072 0 -1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_578
timestamp 1608254825
transform 1 0 29624 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _2349_
timestamp 1608254825
transform 1 0 29716 0 -1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_66_342
timestamp 1608254825
transform 1 0 32568 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_340
timestamp 1608254825
transform 1 0 32384 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_66_332
timestamp 1608254825
transform 1 0 31648 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_66_320
timestamp 1608254825
transform 1 0 30544 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_579
timestamp 1608254825
transform 1 0 32476 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_354
timestamp 1608254825
transform 1 0 33672 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_385
timestamp 1608254825
transform 1 0 36524 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_373
timestamp 1608254825
transform 1 0 35420 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_366
timestamp 1608254825
transform 1 0 34776 0 -1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_580
timestamp 1608254825
transform 1 0 35328 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_404
timestamp 1608254825
transform 1 0 38272 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_397
timestamp 1608254825
transform 1 0 37628 0 -1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_581
timestamp 1608254825
transform 1 0 38180 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_66_416
timestamp 1608254825
transform 1 0 39376 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1608254825
transform -1 0 39836 0 -1 38624
box -38 -48 314 592
<< labels >>
rlabel metal2 s 3330 40200 3386 41000 6 CLK_LED
port 0 nsew signal tristate
rlabel metal2 s 22466 40200 22522 41000 6 DATA_AVAILABLE[0]
port 1 nsew signal input
rlabel metal2 s 18234 40200 18290 41000 6 DATA_AVAILABLE[1]
port 2 nsew signal input
rlabel metal3 s 0 13064 800 13184 6 DATA_AVAILABLE[2]
port 3 nsew signal input
rlabel metal2 s 35162 40200 35218 41000 6 DATA_AVAILABLE[3]
port 4 nsew signal input
rlabel metal2 s 19522 0 19578 800 6 DATA_FROM_HASH[0]
port 5 nsew signal input
rlabel metal2 s 23754 0 23810 800 6 DATA_FROM_HASH[1]
port 6 nsew signal input
rlabel metal2 s 30930 40200 30986 41000 6 DATA_FROM_HASH[2]
port 7 nsew signal input
rlabel metal2 s 5538 40200 5594 41000 6 DATA_FROM_HASH[3]
port 8 nsew signal input
rlabel metal3 s 0 19320 800 19440 6 DATA_FROM_HASH[4]
port 9 nsew signal input
rlabel metal3 s 40200 10344 41000 10464 6 DATA_FROM_HASH[5]
port 10 nsew signal input
rlabel metal2 s 16026 40200 16082 41000 6 DATA_FROM_HASH[6]
port 11 nsew signal input
rlabel metal2 s 25778 0 25834 800 6 DATA_FROM_HASH[7]
port 12 nsew signal input
rlabel metal3 s 0 28840 800 28960 6 DATA_TO_HASH[0]
port 13 nsew signal tristate
rlabel metal2 s 37186 40200 37242 41000 6 DATA_TO_HASH[1]
port 14 nsew signal tristate
rlabel metal2 s 4618 0 4674 800 6 DATA_TO_HASH[2]
port 15 nsew signal tristate
rlabel metal2 s 36450 0 36506 800 6 DATA_TO_HASH[3]
port 16 nsew signal tristate
rlabel metal2 s 7562 40200 7618 41000 6 DATA_TO_HASH[4]
port 17 nsew signal tristate
rlabel metal3 s 40200 1096 41000 1216 6 DATA_TO_HASH[5]
port 18 nsew signal tristate
rlabel metal3 s 40200 19864 41000 19984 6 DATA_TO_HASH[6]
port 19 nsew signal tristate
rlabel metal2 s 34242 0 34298 800 6 DATA_TO_HASH[7]
port 20 nsew signal tristate
rlabel metal2 s 24490 40200 24546 41000 6 EXT_RESET_N_fromHost
port 21 nsew signal input
rlabel metal3 s 0 31832 800 31952 6 EXT_RESET_N_toClient
port 22 nsew signal tristate
rlabel metal2 s 32218 0 32274 800 6 HASH_ADDR[0]
port 23 nsew signal tristate
rlabel metal2 s 32954 40200 33010 41000 6 HASH_ADDR[1]
port 24 nsew signal tristate
rlabel metal2 s 11058 0 11114 800 6 HASH_ADDR[2]
port 25 nsew signal tristate
rlabel metal2 s 28722 40200 28778 41000 6 HASH_ADDR[3]
port 26 nsew signal tristate
rlabel metal3 s 0 6808 800 6928 6 HASH_ADDR[4]
port 27 nsew signal tristate
rlabel metal3 s 0 10072 800 10192 6 HASH_ADDR[5]
port 28 nsew signal tristate
rlabel metal2 s 14002 40200 14058 41000 6 HASH_EN
port 29 nsew signal tristate
rlabel metal3 s 0 16328 800 16448 6 HASH_LED
port 30 nsew signal tristate
rlabel metal3 s 40200 13608 41000 13728 6 ID_fromClient
port 31 nsew signal input
rlabel metal3 s 0 35096 800 35216 6 ID_toHost
port 32 nsew signal tristate
rlabel metal3 s 40200 22856 41000 22976 6 IRQ_OUT_fromClient
port 33 nsew signal input
rlabel metal3 s 0 3816 800 3936 6 IRQ_OUT_toHost
port 34 nsew signal tristate
rlabel metal2 s 8850 0 8906 800 6 M1_CLK_IN
port 35 nsew signal input
rlabel metal2 s 6826 0 6882 800 6 M1_CLK_SELECT
port 36 nsew signal input
rlabel metal2 s 27986 0 28042 800 6 MACRO_RD_SELECT[0]
port 37 nsew signal tristate
rlabel metal2 s 21546 0 21602 800 6 MACRO_RD_SELECT[1]
port 38 nsew signal tristate
rlabel metal2 s 17314 0 17370 800 6 MACRO_RD_SELECT[2]
port 39 nsew signal tristate
rlabel metal2 s 13082 0 13138 800 6 MACRO_RD_SELECT[3]
port 40 nsew signal tristate
rlabel metal2 s 9770 40200 9826 41000 6 MACRO_WR_SELECT[0]
port 41 nsew signal tristate
rlabel metal2 s 2594 0 2650 800 6 MACRO_WR_SELECT[1]
port 42 nsew signal tristate
rlabel metal2 s 39394 40200 39450 41000 6 MACRO_WR_SELECT[2]
port 43 nsew signal tristate
rlabel metal3 s 40200 7352 41000 7472 6 MACRO_WR_SELECT[3]
port 44 nsew signal tristate
rlabel metal2 s 1306 40200 1362 41000 6 MISO_fromClient
port 45 nsew signal input
rlabel metal2 s 26698 40200 26754 41000 6 MISO_toHost
port 46 nsew signal tristate
rlabel metal3 s 40200 38632 41000 38752 6 MOSI_fromHost
port 47 nsew signal input
rlabel metal3 s 40200 16600 41000 16720 6 MOSI_toClient
port 48 nsew signal tristate
rlabel metal3 s 40200 4088 41000 4208 6 PLL_INPUT
port 49 nsew signal input
rlabel metal3 s 0 22584 800 22704 6 S1_CLK_IN
port 50 nsew signal input
rlabel metal3 s 40200 35368 41000 35488 6 S1_CLK_SELECT
port 51 nsew signal input
rlabel metal3 s 40200 32376 41000 32496 6 SCLK_fromHost
port 52 nsew signal input
rlabel metal3 s 0 38088 800 38208 6 SCLK_toClient
port 53 nsew signal tristate
rlabel metal2 s 20258 40200 20314 41000 6 SCSN_fromHost
port 54 nsew signal input
rlabel metal3 s 40200 29112 41000 29232 6 SCSN_toClient
port 55 nsew signal tristate
rlabel metal2 s 570 0 626 800 6 THREAD_COUNT[0]
port 56 nsew signal input
rlabel metal3 s 40200 26120 41000 26240 6 THREAD_COUNT[1]
port 57 nsew signal input
rlabel metal2 s 15290 0 15346 800 6 THREAD_COUNT[2]
port 58 nsew signal input
rlabel metal2 s 11794 40200 11850 41000 6 THREAD_COUNT[3]
port 59 nsew signal input
rlabel metal3 s 0 25576 800 25696 6 m1_clk_local
port 60 nsew signal tristate
rlabel metal2 s 30010 0 30066 800 6 one
port 61 nsew signal tristate
rlabel metal2 s 38474 0 38530 800 6 zero
port 62 nsew signal tristate
rlabel metal4 s 34928 2128 35248 38672 6 vccd1
port 63 nsew power bidirectional
rlabel metal4 s 4208 2128 4528 38672 6 vccd1
port 64 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 38672 6 vssd1
port 65 nsew ground bidirectional
rlabel metal4 s 35588 2176 35908 38624 6 vccd2
port 66 nsew power bidirectional
rlabel metal4 s 4868 2176 5188 38624 6 vccd2
port 67 nsew power bidirectional
rlabel metal4 s 20228 2176 20548 38624 6 vssd2
port 68 nsew ground bidirectional
rlabel metal4 s 36248 2176 36568 38624 6 vdda1
port 69 nsew power bidirectional
rlabel metal4 s 5528 2176 5848 38624 6 vdda1
port 70 nsew power bidirectional
rlabel metal4 s 20888 2176 21208 38624 6 vssa1
port 71 nsew ground bidirectional
rlabel metal4 s 36908 2176 37228 38624 6 vdda2
port 72 nsew power bidirectional
rlabel metal4 s 6188 2176 6508 38624 6 vdda2
port 73 nsew power bidirectional
rlabel metal4 s 21548 2176 21868 38624 6 vssa2
port 74 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 41000 41000
<< end >>

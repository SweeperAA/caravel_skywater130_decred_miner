VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_project_wrapper
  CLASS BLOCK ;
  FOREIGN user_project_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 2920.000 BY 3520.000 ;
  PIN analog_io[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 28.980 2924.800 30.180 ;
    END
  END analog_io[0]
  PIN analog_io[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 2374.980 2924.800 2376.180 ;
    END
  END analog_io[10]
  PIN analog_io[11]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 2609.580 2924.800 2610.780 ;
    END
  END analog_io[11]
  PIN analog_io[12]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 2844.180 2924.800 2845.380 ;
    END
  END analog_io[12]
  PIN analog_io[13]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 3078.780 2924.800 3079.980 ;
    END
  END analog_io[13]
  PIN analog_io[14]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 3313.380 2924.800 3314.580 ;
    END
  END analog_io[14]
  PIN analog_io[15]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2879.090 3519.700 2879.650 3524.800 ;
    END
  END analog_io[15]
  PIN analog_io[16]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2554.790 3519.700 2555.350 3524.800 ;
    END
  END analog_io[16]
  PIN analog_io[17]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2230.490 3519.700 2231.050 3524.800 ;
    END
  END analog_io[17]
  PIN analog_io[18]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1905.730 3519.700 1906.290 3524.800 ;
    END
  END analog_io[18]
  PIN analog_io[19]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1581.430 3519.700 1581.990 3524.800 ;
    END
  END analog_io[19]
  PIN analog_io[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 263.580 2924.800 264.780 ;
    END
  END analog_io[1]
  PIN analog_io[20]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1257.130 3519.700 1257.690 3524.800 ;
    END
  END analog_io[20]
  PIN analog_io[21]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 932.370 3519.700 932.930 3524.800 ;
    END
  END analog_io[21]
  PIN analog_io[22]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 608.070 3519.700 608.630 3524.800 ;
    END
  END analog_io[22]
  PIN analog_io[23]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.770 3519.700 284.330 3524.800 ;
    END
  END analog_io[23]
  PIN analog_io[24]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3482.700 0.300 3483.900 ;
    END
  END analog_io[24]
  PIN analog_io[25]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3195.060 0.300 3196.260 ;
    END
  END analog_io[25]
  PIN analog_io[26]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2908.100 0.300 2909.300 ;
    END
  END analog_io[26]
  PIN analog_io[27]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2620.460 0.300 2621.660 ;
    END
  END analog_io[27]
  PIN analog_io[28]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2333.500 0.300 2334.700 ;
    END
  END analog_io[28]
  PIN analog_io[29]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2045.860 0.300 2047.060 ;
    END
  END analog_io[29]
  PIN analog_io[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 498.180 2924.800 499.380 ;
    END
  END analog_io[2]
  PIN analog_io[30]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1758.900 0.300 1760.100 ;
    END
  END analog_io[30]
  PIN analog_io[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 732.780 2924.800 733.980 ;
    END
  END analog_io[3]
  PIN analog_io[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 967.380 2924.800 968.580 ;
    END
  END analog_io[4]
  PIN analog_io[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 1201.980 2924.800 1203.180 ;
    END
  END analog_io[5]
  PIN analog_io[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 1436.580 2924.800 1437.780 ;
    END
  END analog_io[6]
  PIN analog_io[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 1671.180 2924.800 1672.380 ;
    END
  END analog_io[7]
  PIN analog_io[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 1905.780 2924.800 1906.980 ;
    END
  END analog_io[8]
  PIN analog_io[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 2140.380 2924.800 2141.580 ;
    END
  END analog_io[9]
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 87.460 2924.800 88.660 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 2433.460 2924.800 2434.660 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 2668.740 2924.800 2669.940 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 2903.340 2924.800 2904.540 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 3137.940 2924.800 3139.140 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 3372.540 2924.800 3373.740 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2798.130 3519.700 2798.690 3524.800 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2473.830 3519.700 2474.390 3524.800 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2149.070 3519.700 2149.630 3524.800 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1824.770 3519.700 1825.330 3524.800 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1500.470 3519.700 1501.030 3524.800 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 322.060 2924.800 323.260 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1175.710 3519.700 1176.270 3524.800 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 851.410 3519.700 851.970 3524.800 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 527.110 3519.700 527.670 3524.800 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.350 3519.700 202.910 3524.800 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3410.620 0.300 3411.820 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3123.660 0.300 3124.860 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2836.020 0.300 2837.220 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2549.060 0.300 2550.260 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2261.420 0.300 2262.620 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1974.460 0.300 1975.660 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 556.660 2924.800 557.860 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1686.820 0.300 1688.020 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1471.260 0.300 1472.460 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1255.700 0.300 1256.900 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1040.140 0.300 1041.340 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 824.580 0.300 825.780 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 609.700 0.300 610.900 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 394.140 0.300 395.340 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 178.580 0.300 179.780 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 791.260 2924.800 792.460 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 1025.860 2924.800 1027.060 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 1260.460 2924.800 1261.660 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 1495.060 2924.800 1496.260 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 1729.660 2924.800 1730.860 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 1964.260 2924.800 1965.460 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 2198.860 2924.800 2200.060 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 204.420 2924.800 205.620 ;
    END
  END io_oeb[0]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 439.020 2924.800 440.220 ;
    END
  END io_oeb[1]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2117.940 0.300 2119.140 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1830.300 0.300 1831.500 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 673.620 2924.800 674.820 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1543.340 0.300 1544.540 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1327.780 0.300 1328.980 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1112.220 0.300 1113.420 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 896.660 0.300 897.860 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 681.100 0.300 682.300 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 465.540 0.300 466.740 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 249.980 0.300 251.180 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 35.100 0.300 36.300 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 908.900 2924.800 910.100 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 1143.500 2924.800 1144.700 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 1378.100 2924.800 1379.300 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 1612.700 2924.800 1613.900 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 1847.300 2924.800 1848.500 ;
    END
  END io_oeb[7]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 145.940 2924.800 147.140 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 2492.620 2924.800 2493.820 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 2727.220 2924.800 2728.420 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 2961.820 2924.800 2963.020 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 3196.420 2924.800 3197.620 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 3431.020 2924.800 3432.220 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2717.170 3519.700 2717.730 3524.800 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2392.410 3519.700 2392.970 3524.800 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2068.110 3519.700 2068.670 3524.800 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1743.810 3519.700 1744.370 3524.800 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1419.050 3519.700 1419.610 3524.800 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 380.540 2924.800 381.740 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1094.750 3519.700 1095.310 3524.800 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 770.450 3519.700 771.010 3524.800 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 445.690 3519.700 446.250 3524.800 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.390 3519.700 121.950 3524.800 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3339.220 0.300 3340.420 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3051.580 0.300 3052.780 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2764.620 0.300 2765.820 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2476.980 0.300 2478.180 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2189.340 0.300 2190.540 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1902.380 0.300 1903.580 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 615.140 2924.800 616.340 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1614.740 0.300 1615.940 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1399.860 0.300 1401.060 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1184.300 0.300 1185.500 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 968.740 0.300 969.940 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 753.180 0.300 754.380 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 537.620 0.300 538.820 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 322.060 0.300 323.260 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 106.500 0.300 107.700 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 849.740 2924.800 850.940 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 1084.340 2924.800 1085.540 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 1318.940 2924.800 1320.140 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 1553.540 2924.800 1554.740 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 1788.820 2924.800 1790.020 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 2023.420 2924.800 2024.620 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 2258.020 2924.800 2259.220 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 632.910 -4.800 633.470 0.300 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2417.250 -4.800 2417.810 0.300 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2434.730 -4.800 2435.290 0.300 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2452.670 -4.800 2453.230 0.300 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2470.610 -4.800 2471.170 0.300 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2488.550 -4.800 2489.110 0.300 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2506.030 -4.800 2506.590 0.300 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2523.970 -4.800 2524.530 0.300 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2541.910 -4.800 2542.470 0.300 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2559.850 -4.800 2560.410 0.300 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2577.790 -4.800 2578.350 0.300 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 811.390 -4.800 811.950 0.300 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2595.270 -4.800 2595.830 0.300 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2613.210 -4.800 2613.770 0.300 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2631.150 -4.800 2631.710 0.300 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2649.090 -4.800 2649.650 0.300 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2667.030 -4.800 2667.590 0.300 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2684.510 -4.800 2685.070 0.300 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2702.450 -4.800 2703.010 0.300 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2720.390 -4.800 2720.950 0.300 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2738.330 -4.800 2738.890 0.300 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2755.810 -4.800 2756.370 0.300 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 829.330 -4.800 829.890 0.300 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2773.750 -4.800 2774.310 0.300 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2791.690 -4.800 2792.250 0.300 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2809.630 -4.800 2810.190 0.300 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2827.570 -4.800 2828.130 0.300 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2845.050 -4.800 2845.610 0.300 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2862.990 -4.800 2863.550 0.300 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2880.930 -4.800 2881.490 0.300 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2898.870 -4.800 2899.430 0.300 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 846.810 -4.800 847.370 0.300 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 864.750 -4.800 865.310 0.300 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 882.690 -4.800 883.250 0.300 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 900.630 -4.800 901.190 0.300 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 918.570 -4.800 919.130 0.300 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 936.050 -4.800 936.610 0.300 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 953.990 -4.800 954.550 0.300 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 971.930 -4.800 972.490 0.300 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 650.850 -4.800 651.410 0.300 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 989.870 -4.800 990.430 0.300 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1007.350 -4.800 1007.910 0.300 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1025.290 -4.800 1025.850 0.300 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1043.230 -4.800 1043.790 0.300 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1061.170 -4.800 1061.730 0.300 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1079.110 -4.800 1079.670 0.300 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1096.590 -4.800 1097.150 0.300 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1114.530 -4.800 1115.090 0.300 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1132.470 -4.800 1133.030 0.300 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1150.410 -4.800 1150.970 0.300 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 668.790 -4.800 669.350 0.300 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1168.350 -4.800 1168.910 0.300 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1185.830 -4.800 1186.390 0.300 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1203.770 -4.800 1204.330 0.300 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1221.710 -4.800 1222.270 0.300 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1239.650 -4.800 1240.210 0.300 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1257.130 -4.800 1257.690 0.300 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1275.070 -4.800 1275.630 0.300 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1293.010 -4.800 1293.570 0.300 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1310.950 -4.800 1311.510 0.300 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1328.890 -4.800 1329.450 0.300 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 686.270 -4.800 686.830 0.300 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1346.370 -4.800 1346.930 0.300 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1364.310 -4.800 1364.870 0.300 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1382.250 -4.800 1382.810 0.300 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1400.190 -4.800 1400.750 0.300 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1418.130 -4.800 1418.690 0.300 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1435.610 -4.800 1436.170 0.300 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1453.550 -4.800 1454.110 0.300 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1471.490 -4.800 1472.050 0.300 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1489.430 -4.800 1489.990 0.300 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1506.910 -4.800 1507.470 0.300 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 704.210 -4.800 704.770 0.300 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1524.850 -4.800 1525.410 0.300 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1542.790 -4.800 1543.350 0.300 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1560.730 -4.800 1561.290 0.300 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1578.670 -4.800 1579.230 0.300 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1596.150 -4.800 1596.710 0.300 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1614.090 -4.800 1614.650 0.300 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1632.030 -4.800 1632.590 0.300 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1649.970 -4.800 1650.530 0.300 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1667.910 -4.800 1668.470 0.300 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1685.390 -4.800 1685.950 0.300 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 722.150 -4.800 722.710 0.300 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1703.330 -4.800 1703.890 0.300 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1721.270 -4.800 1721.830 0.300 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1739.210 -4.800 1739.770 0.300 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1756.690 -4.800 1757.250 0.300 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1774.630 -4.800 1775.190 0.300 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1792.570 -4.800 1793.130 0.300 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1810.510 -4.800 1811.070 0.300 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1828.450 -4.800 1829.010 0.300 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1845.930 -4.800 1846.490 0.300 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1863.870 -4.800 1864.430 0.300 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 740.090 -4.800 740.650 0.300 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1881.810 -4.800 1882.370 0.300 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1899.750 -4.800 1900.310 0.300 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1917.690 -4.800 1918.250 0.300 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1935.170 -4.800 1935.730 0.300 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1953.110 -4.800 1953.670 0.300 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1971.050 -4.800 1971.610 0.300 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1988.990 -4.800 1989.550 0.300 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2006.470 -4.800 2007.030 0.300 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2024.410 -4.800 2024.970 0.300 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2042.350 -4.800 2042.910 0.300 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 757.570 -4.800 758.130 0.300 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2060.290 -4.800 2060.850 0.300 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2078.230 -4.800 2078.790 0.300 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2095.710 -4.800 2096.270 0.300 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2113.650 -4.800 2114.210 0.300 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2131.590 -4.800 2132.150 0.300 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2149.530 -4.800 2150.090 0.300 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2167.470 -4.800 2168.030 0.300 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2184.950 -4.800 2185.510 0.300 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2202.890 -4.800 2203.450 0.300 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2220.830 -4.800 2221.390 0.300 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 775.510 -4.800 776.070 0.300 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2238.770 -4.800 2239.330 0.300 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2256.250 -4.800 2256.810 0.300 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2274.190 -4.800 2274.750 0.300 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2292.130 -4.800 2292.690 0.300 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2310.070 -4.800 2310.630 0.300 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2328.010 -4.800 2328.570 0.300 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2345.490 -4.800 2346.050 0.300 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2363.430 -4.800 2363.990 0.300 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2381.370 -4.800 2381.930 0.300 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2399.310 -4.800 2399.870 0.300 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 793.450 -4.800 794.010 0.300 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 638.890 -4.800 639.450 0.300 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2422.770 -4.800 2423.330 0.300 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2440.710 -4.800 2441.270 0.300 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2458.650 -4.800 2459.210 0.300 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2476.590 -4.800 2477.150 0.300 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2494.530 -4.800 2495.090 0.300 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2512.010 -4.800 2512.570 0.300 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2529.950 -4.800 2530.510 0.300 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2547.890 -4.800 2548.450 0.300 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2565.830 -4.800 2566.390 0.300 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2583.770 -4.800 2584.330 0.300 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 817.370 -4.800 817.930 0.300 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2601.250 -4.800 2601.810 0.300 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2619.190 -4.800 2619.750 0.300 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2637.130 -4.800 2637.690 0.300 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2655.070 -4.800 2655.630 0.300 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2672.550 -4.800 2673.110 0.300 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2690.490 -4.800 2691.050 0.300 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2708.430 -4.800 2708.990 0.300 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2726.370 -4.800 2726.930 0.300 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2744.310 -4.800 2744.870 0.300 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2761.790 -4.800 2762.350 0.300 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 835.310 -4.800 835.870 0.300 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2779.730 -4.800 2780.290 0.300 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2797.670 -4.800 2798.230 0.300 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2815.610 -4.800 2816.170 0.300 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2833.550 -4.800 2834.110 0.300 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2851.030 -4.800 2851.590 0.300 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2868.970 -4.800 2869.530 0.300 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2886.910 -4.800 2887.470 0.300 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2904.850 -4.800 2905.410 0.300 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 852.790 -4.800 853.350 0.300 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 870.730 -4.800 871.290 0.300 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 888.670 -4.800 889.230 0.300 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 906.610 -4.800 907.170 0.300 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 924.090 -4.800 924.650 0.300 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 942.030 -4.800 942.590 0.300 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 959.970 -4.800 960.530 0.300 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 977.910 -4.800 978.470 0.300 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 656.830 -4.800 657.390 0.300 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 995.850 -4.800 996.410 0.300 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1013.330 -4.800 1013.890 0.300 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1031.270 -4.800 1031.830 0.300 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1049.210 -4.800 1049.770 0.300 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1067.150 -4.800 1067.710 0.300 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1085.090 -4.800 1085.650 0.300 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1102.570 -4.800 1103.130 0.300 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1120.510 -4.800 1121.070 0.300 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1138.450 -4.800 1139.010 0.300 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1156.390 -4.800 1156.950 0.300 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 674.310 -4.800 674.870 0.300 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1173.870 -4.800 1174.430 0.300 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1191.810 -4.800 1192.370 0.300 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1209.750 -4.800 1210.310 0.300 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1227.690 -4.800 1228.250 0.300 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1245.630 -4.800 1246.190 0.300 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1263.110 -4.800 1263.670 0.300 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1281.050 -4.800 1281.610 0.300 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1298.990 -4.800 1299.550 0.300 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1316.930 -4.800 1317.490 0.300 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1334.870 -4.800 1335.430 0.300 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 692.250 -4.800 692.810 0.300 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1352.350 -4.800 1352.910 0.300 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1370.290 -4.800 1370.850 0.300 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1388.230 -4.800 1388.790 0.300 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1406.170 -4.800 1406.730 0.300 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1423.650 -4.800 1424.210 0.300 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1441.590 -4.800 1442.150 0.300 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1459.530 -4.800 1460.090 0.300 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1477.470 -4.800 1478.030 0.300 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1495.410 -4.800 1495.970 0.300 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1512.890 -4.800 1513.450 0.300 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 710.190 -4.800 710.750 0.300 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1530.830 -4.800 1531.390 0.300 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1548.770 -4.800 1549.330 0.300 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1566.710 -4.800 1567.270 0.300 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1584.650 -4.800 1585.210 0.300 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1602.130 -4.800 1602.690 0.300 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1620.070 -4.800 1620.630 0.300 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1638.010 -4.800 1638.570 0.300 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1655.950 -4.800 1656.510 0.300 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1673.430 -4.800 1673.990 0.300 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1691.370 -4.800 1691.930 0.300 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 728.130 -4.800 728.690 0.300 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1709.310 -4.800 1709.870 0.300 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1727.250 -4.800 1727.810 0.300 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1745.190 -4.800 1745.750 0.300 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1762.670 -4.800 1763.230 0.300 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1780.610 -4.800 1781.170 0.300 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1798.550 -4.800 1799.110 0.300 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1816.490 -4.800 1817.050 0.300 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1834.430 -4.800 1834.990 0.300 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1851.910 -4.800 1852.470 0.300 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1869.850 -4.800 1870.410 0.300 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 746.070 -4.800 746.630 0.300 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1887.790 -4.800 1888.350 0.300 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1905.730 -4.800 1906.290 0.300 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1923.210 -4.800 1923.770 0.300 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1941.150 -4.800 1941.710 0.300 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1959.090 -4.800 1959.650 0.300 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1977.030 -4.800 1977.590 0.300 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1994.970 -4.800 1995.530 0.300 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2012.450 -4.800 2013.010 0.300 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2030.390 -4.800 2030.950 0.300 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2048.330 -4.800 2048.890 0.300 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 763.550 -4.800 764.110 0.300 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2066.270 -4.800 2066.830 0.300 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2084.210 -4.800 2084.770 0.300 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2101.690 -4.800 2102.250 0.300 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2119.630 -4.800 2120.190 0.300 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2137.570 -4.800 2138.130 0.300 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2155.510 -4.800 2156.070 0.300 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2172.990 -4.800 2173.550 0.300 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2190.930 -4.800 2191.490 0.300 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2208.870 -4.800 2209.430 0.300 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2226.810 -4.800 2227.370 0.300 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 781.490 -4.800 782.050 0.300 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2244.750 -4.800 2245.310 0.300 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2262.230 -4.800 2262.790 0.300 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2280.170 -4.800 2280.730 0.300 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2298.110 -4.800 2298.670 0.300 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2316.050 -4.800 2316.610 0.300 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2333.990 -4.800 2334.550 0.300 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2351.470 -4.800 2352.030 0.300 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2369.410 -4.800 2369.970 0.300 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2387.350 -4.800 2387.910 0.300 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2405.290 -4.800 2405.850 0.300 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 799.430 -4.800 799.990 0.300 ;
    END
  END la_data_out[9]
  PIN la_oen[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 644.870 -4.800 645.430 0.300 ;
    END
  END la_oen[0]
  PIN la_oen[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2428.750 -4.800 2429.310 0.300 ;
    END
  END la_oen[100]
  PIN la_oen[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2446.690 -4.800 2447.250 0.300 ;
    END
  END la_oen[101]
  PIN la_oen[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2464.630 -4.800 2465.190 0.300 ;
    END
  END la_oen[102]
  PIN la_oen[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2482.570 -4.800 2483.130 0.300 ;
    END
  END la_oen[103]
  PIN la_oen[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2500.510 -4.800 2501.070 0.300 ;
    END
  END la_oen[104]
  PIN la_oen[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2517.990 -4.800 2518.550 0.300 ;
    END
  END la_oen[105]
  PIN la_oen[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2535.930 -4.800 2536.490 0.300 ;
    END
  END la_oen[106]
  PIN la_oen[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2553.870 -4.800 2554.430 0.300 ;
    END
  END la_oen[107]
  PIN la_oen[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2571.810 -4.800 2572.370 0.300 ;
    END
  END la_oen[108]
  PIN la_oen[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2589.290 -4.800 2589.850 0.300 ;
    END
  END la_oen[109]
  PIN la_oen[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 823.350 -4.800 823.910 0.300 ;
    END
  END la_oen[10]
  PIN la_oen[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2607.230 -4.800 2607.790 0.300 ;
    END
  END la_oen[110]
  PIN la_oen[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2625.170 -4.800 2625.730 0.300 ;
    END
  END la_oen[111]
  PIN la_oen[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2643.110 -4.800 2643.670 0.300 ;
    END
  END la_oen[112]
  PIN la_oen[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2661.050 -4.800 2661.610 0.300 ;
    END
  END la_oen[113]
  PIN la_oen[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2678.530 -4.800 2679.090 0.300 ;
    END
  END la_oen[114]
  PIN la_oen[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2696.470 -4.800 2697.030 0.300 ;
    END
  END la_oen[115]
  PIN la_oen[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2714.410 -4.800 2714.970 0.300 ;
    END
  END la_oen[116]
  PIN la_oen[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2732.350 -4.800 2732.910 0.300 ;
    END
  END la_oen[117]
  PIN la_oen[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2750.290 -4.800 2750.850 0.300 ;
    END
  END la_oen[118]
  PIN la_oen[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2767.770 -4.800 2768.330 0.300 ;
    END
  END la_oen[119]
  PIN la_oen[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 840.830 -4.800 841.390 0.300 ;
    END
  END la_oen[11]
  PIN la_oen[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2785.710 -4.800 2786.270 0.300 ;
    END
  END la_oen[120]
  PIN la_oen[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2803.650 -4.800 2804.210 0.300 ;
    END
  END la_oen[121]
  PIN la_oen[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2821.590 -4.800 2822.150 0.300 ;
    END
  END la_oen[122]
  PIN la_oen[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2839.070 -4.800 2839.630 0.300 ;
    END
  END la_oen[123]
  PIN la_oen[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2857.010 -4.800 2857.570 0.300 ;
    END
  END la_oen[124]
  PIN la_oen[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2874.950 -4.800 2875.510 0.300 ;
    END
  END la_oen[125]
  PIN la_oen[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2892.890 -4.800 2893.450 0.300 ;
    END
  END la_oen[126]
  PIN la_oen[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2910.830 -4.800 2911.390 0.300 ;
    END
  END la_oen[127]
  PIN la_oen[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 858.770 -4.800 859.330 0.300 ;
    END
  END la_oen[12]
  PIN la_oen[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 876.710 -4.800 877.270 0.300 ;
    END
  END la_oen[13]
  PIN la_oen[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 894.650 -4.800 895.210 0.300 ;
    END
  END la_oen[14]
  PIN la_oen[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 912.590 -4.800 913.150 0.300 ;
    END
  END la_oen[15]
  PIN la_oen[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 930.070 -4.800 930.630 0.300 ;
    END
  END la_oen[16]
  PIN la_oen[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 948.010 -4.800 948.570 0.300 ;
    END
  END la_oen[17]
  PIN la_oen[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 965.950 -4.800 966.510 0.300 ;
    END
  END la_oen[18]
  PIN la_oen[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 983.890 -4.800 984.450 0.300 ;
    END
  END la_oen[19]
  PIN la_oen[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 662.810 -4.800 663.370 0.300 ;
    END
  END la_oen[1]
  PIN la_oen[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1001.830 -4.800 1002.390 0.300 ;
    END
  END la_oen[20]
  PIN la_oen[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1019.310 -4.800 1019.870 0.300 ;
    END
  END la_oen[21]
  PIN la_oen[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1037.250 -4.800 1037.810 0.300 ;
    END
  END la_oen[22]
  PIN la_oen[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1055.190 -4.800 1055.750 0.300 ;
    END
  END la_oen[23]
  PIN la_oen[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1073.130 -4.800 1073.690 0.300 ;
    END
  END la_oen[24]
  PIN la_oen[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1090.610 -4.800 1091.170 0.300 ;
    END
  END la_oen[25]
  PIN la_oen[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1108.550 -4.800 1109.110 0.300 ;
    END
  END la_oen[26]
  PIN la_oen[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1126.490 -4.800 1127.050 0.300 ;
    END
  END la_oen[27]
  PIN la_oen[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1144.430 -4.800 1144.990 0.300 ;
    END
  END la_oen[28]
  PIN la_oen[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1162.370 -4.800 1162.930 0.300 ;
    END
  END la_oen[29]
  PIN la_oen[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 680.290 -4.800 680.850 0.300 ;
    END
  END la_oen[2]
  PIN la_oen[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1179.850 -4.800 1180.410 0.300 ;
    END
  END la_oen[30]
  PIN la_oen[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1197.790 -4.800 1198.350 0.300 ;
    END
  END la_oen[31]
  PIN la_oen[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1215.730 -4.800 1216.290 0.300 ;
    END
  END la_oen[32]
  PIN la_oen[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1233.670 -4.800 1234.230 0.300 ;
    END
  END la_oen[33]
  PIN la_oen[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1251.610 -4.800 1252.170 0.300 ;
    END
  END la_oen[34]
  PIN la_oen[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1269.090 -4.800 1269.650 0.300 ;
    END
  END la_oen[35]
  PIN la_oen[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1287.030 -4.800 1287.590 0.300 ;
    END
  END la_oen[36]
  PIN la_oen[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1304.970 -4.800 1305.530 0.300 ;
    END
  END la_oen[37]
  PIN la_oen[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1322.910 -4.800 1323.470 0.300 ;
    END
  END la_oen[38]
  PIN la_oen[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1340.390 -4.800 1340.950 0.300 ;
    END
  END la_oen[39]
  PIN la_oen[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 698.230 -4.800 698.790 0.300 ;
    END
  END la_oen[3]
  PIN la_oen[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1358.330 -4.800 1358.890 0.300 ;
    END
  END la_oen[40]
  PIN la_oen[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1376.270 -4.800 1376.830 0.300 ;
    END
  END la_oen[41]
  PIN la_oen[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1394.210 -4.800 1394.770 0.300 ;
    END
  END la_oen[42]
  PIN la_oen[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1412.150 -4.800 1412.710 0.300 ;
    END
  END la_oen[43]
  PIN la_oen[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1429.630 -4.800 1430.190 0.300 ;
    END
  END la_oen[44]
  PIN la_oen[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1447.570 -4.800 1448.130 0.300 ;
    END
  END la_oen[45]
  PIN la_oen[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1465.510 -4.800 1466.070 0.300 ;
    END
  END la_oen[46]
  PIN la_oen[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1483.450 -4.800 1484.010 0.300 ;
    END
  END la_oen[47]
  PIN la_oen[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1501.390 -4.800 1501.950 0.300 ;
    END
  END la_oen[48]
  PIN la_oen[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1518.870 -4.800 1519.430 0.300 ;
    END
  END la_oen[49]
  PIN la_oen[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 716.170 -4.800 716.730 0.300 ;
    END
  END la_oen[4]
  PIN la_oen[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1536.810 -4.800 1537.370 0.300 ;
    END
  END la_oen[50]
  PIN la_oen[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1554.750 -4.800 1555.310 0.300 ;
    END
  END la_oen[51]
  PIN la_oen[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1572.690 -4.800 1573.250 0.300 ;
    END
  END la_oen[52]
  PIN la_oen[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1590.170 -4.800 1590.730 0.300 ;
    END
  END la_oen[53]
  PIN la_oen[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1608.110 -4.800 1608.670 0.300 ;
    END
  END la_oen[54]
  PIN la_oen[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1626.050 -4.800 1626.610 0.300 ;
    END
  END la_oen[55]
  PIN la_oen[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1643.990 -4.800 1644.550 0.300 ;
    END
  END la_oen[56]
  PIN la_oen[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1661.930 -4.800 1662.490 0.300 ;
    END
  END la_oen[57]
  PIN la_oen[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1679.410 -4.800 1679.970 0.300 ;
    END
  END la_oen[58]
  PIN la_oen[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1697.350 -4.800 1697.910 0.300 ;
    END
  END la_oen[59]
  PIN la_oen[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 734.110 -4.800 734.670 0.300 ;
    END
  END la_oen[5]
  PIN la_oen[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1715.290 -4.800 1715.850 0.300 ;
    END
  END la_oen[60]
  PIN la_oen[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1733.230 -4.800 1733.790 0.300 ;
    END
  END la_oen[61]
  PIN la_oen[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1751.170 -4.800 1751.730 0.300 ;
    END
  END la_oen[62]
  PIN la_oen[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1768.650 -4.800 1769.210 0.300 ;
    END
  END la_oen[63]
  PIN la_oen[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1786.590 -4.800 1787.150 0.300 ;
    END
  END la_oen[64]
  PIN la_oen[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1804.530 -4.800 1805.090 0.300 ;
    END
  END la_oen[65]
  PIN la_oen[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1822.470 -4.800 1823.030 0.300 ;
    END
  END la_oen[66]
  PIN la_oen[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1839.950 -4.800 1840.510 0.300 ;
    END
  END la_oen[67]
  PIN la_oen[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1857.890 -4.800 1858.450 0.300 ;
    END
  END la_oen[68]
  PIN la_oen[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1875.830 -4.800 1876.390 0.300 ;
    END
  END la_oen[69]
  PIN la_oen[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 752.050 -4.800 752.610 0.300 ;
    END
  END la_oen[6]
  PIN la_oen[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1893.770 -4.800 1894.330 0.300 ;
    END
  END la_oen[70]
  PIN la_oen[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1911.710 -4.800 1912.270 0.300 ;
    END
  END la_oen[71]
  PIN la_oen[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1929.190 -4.800 1929.750 0.300 ;
    END
  END la_oen[72]
  PIN la_oen[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1947.130 -4.800 1947.690 0.300 ;
    END
  END la_oen[73]
  PIN la_oen[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1965.070 -4.800 1965.630 0.300 ;
    END
  END la_oen[74]
  PIN la_oen[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1983.010 -4.800 1983.570 0.300 ;
    END
  END la_oen[75]
  PIN la_oen[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2000.950 -4.800 2001.510 0.300 ;
    END
  END la_oen[76]
  PIN la_oen[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2018.430 -4.800 2018.990 0.300 ;
    END
  END la_oen[77]
  PIN la_oen[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2036.370 -4.800 2036.930 0.300 ;
    END
  END la_oen[78]
  PIN la_oen[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2054.310 -4.800 2054.870 0.300 ;
    END
  END la_oen[79]
  PIN la_oen[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 769.530 -4.800 770.090 0.300 ;
    END
  END la_oen[7]
  PIN la_oen[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2072.250 -4.800 2072.810 0.300 ;
    END
  END la_oen[80]
  PIN la_oen[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2089.730 -4.800 2090.290 0.300 ;
    END
  END la_oen[81]
  PIN la_oen[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2107.670 -4.800 2108.230 0.300 ;
    END
  END la_oen[82]
  PIN la_oen[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2125.610 -4.800 2126.170 0.300 ;
    END
  END la_oen[83]
  PIN la_oen[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2143.550 -4.800 2144.110 0.300 ;
    END
  END la_oen[84]
  PIN la_oen[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2161.490 -4.800 2162.050 0.300 ;
    END
  END la_oen[85]
  PIN la_oen[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2178.970 -4.800 2179.530 0.300 ;
    END
  END la_oen[86]
  PIN la_oen[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2196.910 -4.800 2197.470 0.300 ;
    END
  END la_oen[87]
  PIN la_oen[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2214.850 -4.800 2215.410 0.300 ;
    END
  END la_oen[88]
  PIN la_oen[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2232.790 -4.800 2233.350 0.300 ;
    END
  END la_oen[89]
  PIN la_oen[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 787.470 -4.800 788.030 0.300 ;
    END
  END la_oen[8]
  PIN la_oen[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2250.730 -4.800 2251.290 0.300 ;
    END
  END la_oen[90]
  PIN la_oen[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2268.210 -4.800 2268.770 0.300 ;
    END
  END la_oen[91]
  PIN la_oen[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2286.150 -4.800 2286.710 0.300 ;
    END
  END la_oen[92]
  PIN la_oen[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2304.090 -4.800 2304.650 0.300 ;
    END
  END la_oen[93]
  PIN la_oen[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2322.030 -4.800 2322.590 0.300 ;
    END
  END la_oen[94]
  PIN la_oen[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2339.510 -4.800 2340.070 0.300 ;
    END
  END la_oen[95]
  PIN la_oen[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2357.450 -4.800 2358.010 0.300 ;
    END
  END la_oen[96]
  PIN la_oen[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2375.390 -4.800 2375.950 0.300 ;
    END
  END la_oen[97]
  PIN la_oen[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2393.330 -4.800 2393.890 0.300 ;
    END
  END la_oen[98]
  PIN la_oen[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2411.270 -4.800 2411.830 0.300 ;
    END
  END la_oen[99]
  PIN la_oen[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 805.410 -4.800 805.970 0.300 ;
    END
  END la_oen[9]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1662.390 3519.700 1662.950 3524.800 ;
        RECT 1987.150 3519.700 1987.710 3524.800 ;
        RECT 2311.450 3519.700 2312.010 3524.800 ;
        RECT 2635.750 3519.700 2636.310 3524.800 ;
      LAYER met3 ;
        RECT 2919.700 3489.500 2924.800 3490.700 ;
        RECT 2919.700 3254.900 2924.800 3256.100 ;
        RECT 2919.700 3020.300 2924.800 3021.500 ;
        RECT 2919.700 2785.700 2924.800 2786.900 ;
        RECT 2919.700 2551.100 2924.800 2552.300 ;
        RECT 2919.700 2316.500 2924.800 2317.700 ;
        RECT 2919.700 2081.900 2924.800 2083.100 ;
    END
  END io_oeb[10]
  PIN user_clock2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2916.810 -4.800 2917.370 0.300 ;
    END
  END user_clock2
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.710 -4.800 3.270 0.300 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.230 -4.800 8.790 0.300 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.210 -4.800 14.770 0.300 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.130 -4.800 38.690 0.300 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 240.530 -4.800 241.090 0.300 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 258.010 -4.800 258.570 0.300 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 275.950 -4.800 276.510 0.300 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.890 -4.800 294.450 0.300 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.830 -4.800 312.390 0.300 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 329.770 -4.800 330.330 0.300 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.250 -4.800 347.810 0.300 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 365.190 -4.800 365.750 0.300 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 383.130 -4.800 383.690 0.300 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 401.070 -4.800 401.630 0.300 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.050 -4.800 62.610 0.300 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 419.010 -4.800 419.570 0.300 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 436.490 -4.800 437.050 0.300 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 454.430 -4.800 454.990 0.300 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 472.370 -4.800 472.930 0.300 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 490.310 -4.800 490.870 0.300 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 507.790 -4.800 508.350 0.300 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 525.730 -4.800 526.290 0.300 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 543.670 -4.800 544.230 0.300 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 561.610 -4.800 562.170 0.300 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 579.550 -4.800 580.110 0.300 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.970 -4.800 86.530 0.300 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 597.030 -4.800 597.590 0.300 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 614.970 -4.800 615.530 0.300 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.430 -4.800 109.990 0.300 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.350 -4.800 133.910 0.300 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.290 -4.800 151.850 0.300 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 169.230 -4.800 169.790 0.300 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.710 -4.800 187.270 0.300 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 204.650 -4.800 205.210 0.300 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.590 -4.800 223.150 0.300 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.190 -4.800 20.750 0.300 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.110 -4.800 44.670 0.300 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 246.510 -4.800 247.070 0.300 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 263.990 -4.800 264.550 0.300 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 281.930 -4.800 282.490 0.300 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.870 -4.800 300.430 0.300 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.810 -4.800 318.370 0.300 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 335.750 -4.800 336.310 0.300 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 353.230 -4.800 353.790 0.300 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 371.170 -4.800 371.730 0.300 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 389.110 -4.800 389.670 0.300 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 407.050 -4.800 407.610 0.300 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.030 -4.800 68.590 0.300 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 424.530 -4.800 425.090 0.300 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 442.470 -4.800 443.030 0.300 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 460.410 -4.800 460.970 0.300 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 478.350 -4.800 478.910 0.300 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 496.290 -4.800 496.850 0.300 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 513.770 -4.800 514.330 0.300 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 531.710 -4.800 532.270 0.300 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 549.650 -4.800 550.210 0.300 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 567.590 -4.800 568.150 0.300 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 585.530 -4.800 586.090 0.300 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.490 -4.800 92.050 0.300 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 603.010 -4.800 603.570 0.300 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 620.950 -4.800 621.510 0.300 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.410 -4.800 115.970 0.300 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.330 -4.800 139.890 0.300 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.270 -4.800 157.830 0.300 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.750 -4.800 175.310 0.300 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.690 -4.800 193.250 0.300 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 210.630 -4.800 211.190 0.300 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.570 -4.800 229.130 0.300 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.090 -4.800 50.650 0.300 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 252.490 -4.800 253.050 0.300 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 269.970 -4.800 270.530 0.300 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 287.910 -4.800 288.470 0.300 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.850 -4.800 306.410 0.300 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.790 -4.800 324.350 0.300 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.270 -4.800 341.830 0.300 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 359.210 -4.800 359.770 0.300 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 377.150 -4.800 377.710 0.300 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 395.090 -4.800 395.650 0.300 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 413.030 -4.800 413.590 0.300 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.010 -4.800 74.570 0.300 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 430.510 -4.800 431.070 0.300 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 448.450 -4.800 449.010 0.300 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.390 -4.800 466.950 0.300 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 484.330 -4.800 484.890 0.300 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 502.270 -4.800 502.830 0.300 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 519.750 -4.800 520.310 0.300 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 537.690 -4.800 538.250 0.300 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 555.630 -4.800 556.190 0.300 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 573.570 -4.800 574.130 0.300 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 591.050 -4.800 591.610 0.300 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.470 -4.800 98.030 0.300 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 608.990 -4.800 609.550 0.300 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 626.930 -4.800 627.490 0.300 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.390 -4.800 121.950 0.300 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.310 -4.800 145.870 0.300 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.250 -4.800 163.810 0.300 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.730 -4.800 181.290 0.300 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.670 -4.800 199.230 0.300 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.610 -4.800 217.170 0.300 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 234.550 -4.800 235.110 0.300 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.070 -4.800 56.630 0.300 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.990 -4.800 80.550 0.300 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.450 -4.800 104.010 0.300 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.370 -4.800 127.930 0.300 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.170 -4.800 26.730 0.300 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.150 -4.800 32.710 0.300 ;
    END
  END wbs_we_i
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.430 3519.700 40.990 3524.800 ;
        RECT 364.730 3519.700 365.290 3524.800 ;
        RECT 689.030 3519.700 689.590 3524.800 ;
        RECT 1013.790 3519.700 1014.350 3524.800 ;
        RECT 1338.090 3519.700 1338.650 3524.800 ;
      LAYER met3 ;
        RECT -4.800 3267.140 0.300 3268.340 ;
        RECT -4.800 2979.500 0.300 2980.700 ;
        RECT -4.800 2692.540 0.300 2693.740 ;
        RECT -4.800 2404.900 0.300 2406.100 ;
    END
  END io_oeb[19]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -9.980 -4.620 -6.980 3524.300 ;
        RECT 4.020 3519.700 7.020 3529.000 ;
        RECT 184.020 3519.700 187.020 3529.000 ;
        RECT 364.020 3519.700 367.020 3529.000 ;
        RECT 544.020 3519.700 547.020 3529.000 ;
        RECT 724.020 3519.700 727.020 3529.000 ;
        RECT 904.020 3519.700 907.020 3529.000 ;
        RECT 1084.020 3519.700 1087.020 3529.000 ;
        RECT 1264.020 3519.700 1267.020 3529.000 ;
        RECT 1444.020 3519.700 1447.020 3529.000 ;
        RECT 1624.020 3519.700 1627.020 3529.000 ;
        RECT 1804.020 3519.700 1807.020 3529.000 ;
        RECT 1984.020 3519.700 1987.020 3529.000 ;
        RECT 2164.020 3519.700 2167.020 3529.000 ;
        RECT 2344.020 3519.700 2347.020 3529.000 ;
        RECT 2524.020 3519.700 2527.020 3529.000 ;
        RECT 2704.020 3519.700 2707.020 3529.000 ;
        RECT 2884.020 3519.700 2887.020 3529.000 ;
        RECT 4.020 -9.320 7.020 0.300 ;
        RECT 184.020 -9.320 187.020 0.300 ;
        RECT 364.020 -9.320 367.020 0.300 ;
        RECT 544.020 -9.320 547.020 0.300 ;
        RECT 724.020 -9.320 727.020 0.300 ;
        RECT 904.020 -9.320 907.020 0.300 ;
        RECT 1084.020 -9.320 1087.020 0.300 ;
        RECT 1264.020 -9.320 1267.020 0.300 ;
        RECT 1444.020 -9.320 1447.020 0.300 ;
        RECT 1624.020 -9.320 1627.020 0.300 ;
        RECT 1804.020 -9.320 1807.020 0.300 ;
        RECT 1984.020 -9.320 1987.020 0.300 ;
        RECT 2164.020 -9.320 2167.020 0.300 ;
        RECT 2344.020 -9.320 2347.020 0.300 ;
        RECT 2524.020 -9.320 2527.020 0.300 ;
        RECT 2704.020 -9.320 2707.020 0.300 ;
        RECT 2884.020 -9.320 2887.020 0.300 ;
        RECT 2926.600 -4.620 2929.600 3524.300 ;
      LAYER via4 ;
        RECT -9.070 3523.010 -7.890 3524.190 ;
        RECT -9.070 3521.410 -7.890 3522.590 ;
        RECT 4.930 3523.010 6.110 3524.190 ;
        RECT 4.930 3521.410 6.110 3522.590 ;
        RECT 184.930 3523.010 186.110 3524.190 ;
        RECT 184.930 3521.410 186.110 3522.590 ;
        RECT 364.930 3523.010 366.110 3524.190 ;
        RECT 364.930 3521.410 366.110 3522.590 ;
        RECT 544.930 3523.010 546.110 3524.190 ;
        RECT 544.930 3521.410 546.110 3522.590 ;
        RECT 724.930 3523.010 726.110 3524.190 ;
        RECT 724.930 3521.410 726.110 3522.590 ;
        RECT 904.930 3523.010 906.110 3524.190 ;
        RECT 904.930 3521.410 906.110 3522.590 ;
        RECT 1084.930 3523.010 1086.110 3524.190 ;
        RECT 1084.930 3521.410 1086.110 3522.590 ;
        RECT 1264.930 3523.010 1266.110 3524.190 ;
        RECT 1264.930 3521.410 1266.110 3522.590 ;
        RECT 1444.930 3523.010 1446.110 3524.190 ;
        RECT 1444.930 3521.410 1446.110 3522.590 ;
        RECT 1624.930 3523.010 1626.110 3524.190 ;
        RECT 1624.930 3521.410 1626.110 3522.590 ;
        RECT 1804.930 3523.010 1806.110 3524.190 ;
        RECT 1804.930 3521.410 1806.110 3522.590 ;
        RECT 1984.930 3523.010 1986.110 3524.190 ;
        RECT 1984.930 3521.410 1986.110 3522.590 ;
        RECT 2164.930 3523.010 2166.110 3524.190 ;
        RECT 2164.930 3521.410 2166.110 3522.590 ;
        RECT 2344.930 3523.010 2346.110 3524.190 ;
        RECT 2344.930 3521.410 2346.110 3522.590 ;
        RECT 2524.930 3523.010 2526.110 3524.190 ;
        RECT 2524.930 3521.410 2526.110 3522.590 ;
        RECT 2704.930 3523.010 2706.110 3524.190 ;
        RECT 2704.930 3521.410 2706.110 3522.590 ;
        RECT 2884.930 3523.010 2886.110 3524.190 ;
        RECT 2884.930 3521.410 2886.110 3522.590 ;
        RECT 2927.510 3523.010 2928.690 3524.190 ;
        RECT 2927.510 3521.410 2928.690 3522.590 ;
        RECT -9.070 3431.090 -7.890 3432.270 ;
        RECT -9.070 3429.490 -7.890 3430.670 ;
        RECT -9.070 3251.090 -7.890 3252.270 ;
        RECT -9.070 3249.490 -7.890 3250.670 ;
        RECT -9.070 3071.090 -7.890 3072.270 ;
        RECT -9.070 3069.490 -7.890 3070.670 ;
        RECT -9.070 2891.090 -7.890 2892.270 ;
        RECT -9.070 2889.490 -7.890 2890.670 ;
        RECT -9.070 2711.090 -7.890 2712.270 ;
        RECT -9.070 2709.490 -7.890 2710.670 ;
        RECT -9.070 2531.090 -7.890 2532.270 ;
        RECT -9.070 2529.490 -7.890 2530.670 ;
        RECT -9.070 2351.090 -7.890 2352.270 ;
        RECT -9.070 2349.490 -7.890 2350.670 ;
        RECT -9.070 2171.090 -7.890 2172.270 ;
        RECT -9.070 2169.490 -7.890 2170.670 ;
        RECT -9.070 1991.090 -7.890 1992.270 ;
        RECT -9.070 1989.490 -7.890 1990.670 ;
        RECT -9.070 1811.090 -7.890 1812.270 ;
        RECT -9.070 1809.490 -7.890 1810.670 ;
        RECT -9.070 1631.090 -7.890 1632.270 ;
        RECT -9.070 1629.490 -7.890 1630.670 ;
        RECT -9.070 1451.090 -7.890 1452.270 ;
        RECT -9.070 1449.490 -7.890 1450.670 ;
        RECT -9.070 1271.090 -7.890 1272.270 ;
        RECT -9.070 1269.490 -7.890 1270.670 ;
        RECT -9.070 1091.090 -7.890 1092.270 ;
        RECT -9.070 1089.490 -7.890 1090.670 ;
        RECT -9.070 911.090 -7.890 912.270 ;
        RECT -9.070 909.490 -7.890 910.670 ;
        RECT -9.070 731.090 -7.890 732.270 ;
        RECT -9.070 729.490 -7.890 730.670 ;
        RECT -9.070 551.090 -7.890 552.270 ;
        RECT -9.070 549.490 -7.890 550.670 ;
        RECT -9.070 371.090 -7.890 372.270 ;
        RECT -9.070 369.490 -7.890 370.670 ;
        RECT -9.070 191.090 -7.890 192.270 ;
        RECT -9.070 189.490 -7.890 190.670 ;
        RECT -9.070 11.090 -7.890 12.270 ;
        RECT -9.070 9.490 -7.890 10.670 ;
        RECT 2927.510 3431.090 2928.690 3432.270 ;
        RECT 2927.510 3429.490 2928.690 3430.670 ;
        RECT 2927.510 3251.090 2928.690 3252.270 ;
        RECT 2927.510 3249.490 2928.690 3250.670 ;
        RECT 2927.510 3071.090 2928.690 3072.270 ;
        RECT 2927.510 3069.490 2928.690 3070.670 ;
        RECT 2927.510 2891.090 2928.690 2892.270 ;
        RECT 2927.510 2889.490 2928.690 2890.670 ;
        RECT 2927.510 2711.090 2928.690 2712.270 ;
        RECT 2927.510 2709.490 2928.690 2710.670 ;
        RECT 2927.510 2531.090 2928.690 2532.270 ;
        RECT 2927.510 2529.490 2928.690 2530.670 ;
        RECT 2927.510 2351.090 2928.690 2352.270 ;
        RECT 2927.510 2349.490 2928.690 2350.670 ;
        RECT 2927.510 2171.090 2928.690 2172.270 ;
        RECT 2927.510 2169.490 2928.690 2170.670 ;
        RECT 2927.510 1991.090 2928.690 1992.270 ;
        RECT 2927.510 1989.490 2928.690 1990.670 ;
        RECT 2927.510 1811.090 2928.690 1812.270 ;
        RECT 2927.510 1809.490 2928.690 1810.670 ;
        RECT 2927.510 1631.090 2928.690 1632.270 ;
        RECT 2927.510 1629.490 2928.690 1630.670 ;
        RECT 2927.510 1451.090 2928.690 1452.270 ;
        RECT 2927.510 1449.490 2928.690 1450.670 ;
        RECT 2927.510 1271.090 2928.690 1272.270 ;
        RECT 2927.510 1269.490 2928.690 1270.670 ;
        RECT 2927.510 1091.090 2928.690 1092.270 ;
        RECT 2927.510 1089.490 2928.690 1090.670 ;
        RECT 2927.510 911.090 2928.690 912.270 ;
        RECT 2927.510 909.490 2928.690 910.670 ;
        RECT 2927.510 731.090 2928.690 732.270 ;
        RECT 2927.510 729.490 2928.690 730.670 ;
        RECT 2927.510 551.090 2928.690 552.270 ;
        RECT 2927.510 549.490 2928.690 550.670 ;
        RECT 2927.510 371.090 2928.690 372.270 ;
        RECT 2927.510 369.490 2928.690 370.670 ;
        RECT 2927.510 191.090 2928.690 192.270 ;
        RECT 2927.510 189.490 2928.690 190.670 ;
        RECT 2927.510 11.090 2928.690 12.270 ;
        RECT 2927.510 9.490 2928.690 10.670 ;
        RECT -9.070 -2.910 -7.890 -1.730 ;
        RECT -9.070 -4.510 -7.890 -3.330 ;
        RECT 4.930 -2.910 6.110 -1.730 ;
        RECT 4.930 -4.510 6.110 -3.330 ;
        RECT 184.930 -2.910 186.110 -1.730 ;
        RECT 184.930 -4.510 186.110 -3.330 ;
        RECT 364.930 -2.910 366.110 -1.730 ;
        RECT 364.930 -4.510 366.110 -3.330 ;
        RECT 544.930 -2.910 546.110 -1.730 ;
        RECT 544.930 -4.510 546.110 -3.330 ;
        RECT 724.930 -2.910 726.110 -1.730 ;
        RECT 724.930 -4.510 726.110 -3.330 ;
        RECT 904.930 -2.910 906.110 -1.730 ;
        RECT 904.930 -4.510 906.110 -3.330 ;
        RECT 1084.930 -2.910 1086.110 -1.730 ;
        RECT 1084.930 -4.510 1086.110 -3.330 ;
        RECT 1264.930 -2.910 1266.110 -1.730 ;
        RECT 1264.930 -4.510 1266.110 -3.330 ;
        RECT 1444.930 -2.910 1446.110 -1.730 ;
        RECT 1444.930 -4.510 1446.110 -3.330 ;
        RECT 1624.930 -2.910 1626.110 -1.730 ;
        RECT 1624.930 -4.510 1626.110 -3.330 ;
        RECT 1804.930 -2.910 1806.110 -1.730 ;
        RECT 1804.930 -4.510 1806.110 -3.330 ;
        RECT 1984.930 -2.910 1986.110 -1.730 ;
        RECT 1984.930 -4.510 1986.110 -3.330 ;
        RECT 2164.930 -2.910 2166.110 -1.730 ;
        RECT 2164.930 -4.510 2166.110 -3.330 ;
        RECT 2344.930 -2.910 2346.110 -1.730 ;
        RECT 2344.930 -4.510 2346.110 -3.330 ;
        RECT 2524.930 -2.910 2526.110 -1.730 ;
        RECT 2524.930 -4.510 2526.110 -3.330 ;
        RECT 2704.930 -2.910 2706.110 -1.730 ;
        RECT 2704.930 -4.510 2706.110 -3.330 ;
        RECT 2884.930 -2.910 2886.110 -1.730 ;
        RECT 2884.930 -4.510 2886.110 -3.330 ;
        RECT 2927.510 -2.910 2928.690 -1.730 ;
        RECT 2927.510 -4.510 2928.690 -3.330 ;
      LAYER met5 ;
        RECT -9.980 3524.300 -6.980 3524.310 ;
        RECT 4.020 3524.300 7.020 3524.310 ;
        RECT 184.020 3524.300 187.020 3524.310 ;
        RECT 364.020 3524.300 367.020 3524.310 ;
        RECT 544.020 3524.300 547.020 3524.310 ;
        RECT 724.020 3524.300 727.020 3524.310 ;
        RECT 904.020 3524.300 907.020 3524.310 ;
        RECT 1084.020 3524.300 1087.020 3524.310 ;
        RECT 1264.020 3524.300 1267.020 3524.310 ;
        RECT 1444.020 3524.300 1447.020 3524.310 ;
        RECT 1624.020 3524.300 1627.020 3524.310 ;
        RECT 1804.020 3524.300 1807.020 3524.310 ;
        RECT 1984.020 3524.300 1987.020 3524.310 ;
        RECT 2164.020 3524.300 2167.020 3524.310 ;
        RECT 2344.020 3524.300 2347.020 3524.310 ;
        RECT 2524.020 3524.300 2527.020 3524.310 ;
        RECT 2704.020 3524.300 2707.020 3524.310 ;
        RECT 2884.020 3524.300 2887.020 3524.310 ;
        RECT 2926.600 3524.300 2929.600 3524.310 ;
        RECT -9.980 3521.300 2929.600 3524.300 ;
        RECT -9.980 3521.290 -6.980 3521.300 ;
        RECT 4.020 3521.290 7.020 3521.300 ;
        RECT 184.020 3521.290 187.020 3521.300 ;
        RECT 364.020 3521.290 367.020 3521.300 ;
        RECT 544.020 3521.290 547.020 3521.300 ;
        RECT 724.020 3521.290 727.020 3521.300 ;
        RECT 904.020 3521.290 907.020 3521.300 ;
        RECT 1084.020 3521.290 1087.020 3521.300 ;
        RECT 1264.020 3521.290 1267.020 3521.300 ;
        RECT 1444.020 3521.290 1447.020 3521.300 ;
        RECT 1624.020 3521.290 1627.020 3521.300 ;
        RECT 1804.020 3521.290 1807.020 3521.300 ;
        RECT 1984.020 3521.290 1987.020 3521.300 ;
        RECT 2164.020 3521.290 2167.020 3521.300 ;
        RECT 2344.020 3521.290 2347.020 3521.300 ;
        RECT 2524.020 3521.290 2527.020 3521.300 ;
        RECT 2704.020 3521.290 2707.020 3521.300 ;
        RECT 2884.020 3521.290 2887.020 3521.300 ;
        RECT 2926.600 3521.290 2929.600 3521.300 ;
        RECT -9.980 3432.380 -6.980 3432.390 ;
        RECT 2926.600 3432.380 2929.600 3432.390 ;
        RECT -14.680 3429.380 0.300 3432.380 ;
        RECT 2919.700 3429.380 2934.300 3432.380 ;
        RECT -9.980 3429.370 -6.980 3429.380 ;
        RECT 2926.600 3429.370 2929.600 3429.380 ;
        RECT -9.980 3252.380 -6.980 3252.390 ;
        RECT 2926.600 3252.380 2929.600 3252.390 ;
        RECT -14.680 3249.380 0.300 3252.380 ;
        RECT 2919.700 3249.380 2934.300 3252.380 ;
        RECT -9.980 3249.370 -6.980 3249.380 ;
        RECT 2926.600 3249.370 2929.600 3249.380 ;
        RECT -9.980 3072.380 -6.980 3072.390 ;
        RECT 2926.600 3072.380 2929.600 3072.390 ;
        RECT -14.680 3069.380 0.300 3072.380 ;
        RECT 2919.700 3069.380 2934.300 3072.380 ;
        RECT -9.980 3069.370 -6.980 3069.380 ;
        RECT 2926.600 3069.370 2929.600 3069.380 ;
        RECT -9.980 2892.380 -6.980 2892.390 ;
        RECT 2926.600 2892.380 2929.600 2892.390 ;
        RECT -14.680 2889.380 0.300 2892.380 ;
        RECT 2919.700 2889.380 2934.300 2892.380 ;
        RECT -9.980 2889.370 -6.980 2889.380 ;
        RECT 2926.600 2889.370 2929.600 2889.380 ;
        RECT -9.980 2712.380 -6.980 2712.390 ;
        RECT 2926.600 2712.380 2929.600 2712.390 ;
        RECT -14.680 2709.380 0.300 2712.380 ;
        RECT 2919.700 2709.380 2934.300 2712.380 ;
        RECT -9.980 2709.370 -6.980 2709.380 ;
        RECT 2926.600 2709.370 2929.600 2709.380 ;
        RECT -9.980 2532.380 -6.980 2532.390 ;
        RECT 2926.600 2532.380 2929.600 2532.390 ;
        RECT -14.680 2529.380 0.300 2532.380 ;
        RECT 2919.700 2529.380 2934.300 2532.380 ;
        RECT -9.980 2529.370 -6.980 2529.380 ;
        RECT 2926.600 2529.370 2929.600 2529.380 ;
        RECT -9.980 2352.380 -6.980 2352.390 ;
        RECT 2926.600 2352.380 2929.600 2352.390 ;
        RECT -14.680 2349.380 0.300 2352.380 ;
        RECT 2919.700 2349.380 2934.300 2352.380 ;
        RECT -9.980 2349.370 -6.980 2349.380 ;
        RECT 2926.600 2349.370 2929.600 2349.380 ;
        RECT -9.980 2172.380 -6.980 2172.390 ;
        RECT 2926.600 2172.380 2929.600 2172.390 ;
        RECT -14.680 2169.380 0.300 2172.380 ;
        RECT 2919.700 2169.380 2934.300 2172.380 ;
        RECT -9.980 2169.370 -6.980 2169.380 ;
        RECT 2926.600 2169.370 2929.600 2169.380 ;
        RECT -9.980 1992.380 -6.980 1992.390 ;
        RECT 2926.600 1992.380 2929.600 1992.390 ;
        RECT -14.680 1989.380 0.300 1992.380 ;
        RECT 2919.700 1989.380 2934.300 1992.380 ;
        RECT -9.980 1989.370 -6.980 1989.380 ;
        RECT 2926.600 1989.370 2929.600 1989.380 ;
        RECT -9.980 1812.380 -6.980 1812.390 ;
        RECT 2926.600 1812.380 2929.600 1812.390 ;
        RECT -14.680 1809.380 0.300 1812.380 ;
        RECT 2919.700 1809.380 2934.300 1812.380 ;
        RECT -9.980 1809.370 -6.980 1809.380 ;
        RECT 2926.600 1809.370 2929.600 1809.380 ;
        RECT -9.980 1632.380 -6.980 1632.390 ;
        RECT 2926.600 1632.380 2929.600 1632.390 ;
        RECT -14.680 1629.380 0.300 1632.380 ;
        RECT 2919.700 1629.380 2934.300 1632.380 ;
        RECT -9.980 1629.370 -6.980 1629.380 ;
        RECT 2926.600 1629.370 2929.600 1629.380 ;
        RECT -9.980 1452.380 -6.980 1452.390 ;
        RECT 2926.600 1452.380 2929.600 1452.390 ;
        RECT -14.680 1449.380 0.300 1452.380 ;
        RECT 2919.700 1449.380 2934.300 1452.380 ;
        RECT -9.980 1449.370 -6.980 1449.380 ;
        RECT 2926.600 1449.370 2929.600 1449.380 ;
        RECT -9.980 1272.380 -6.980 1272.390 ;
        RECT 2926.600 1272.380 2929.600 1272.390 ;
        RECT -14.680 1269.380 0.300 1272.380 ;
        RECT 2919.700 1269.380 2934.300 1272.380 ;
        RECT -9.980 1269.370 -6.980 1269.380 ;
        RECT 2926.600 1269.370 2929.600 1269.380 ;
        RECT -9.980 1092.380 -6.980 1092.390 ;
        RECT 2926.600 1092.380 2929.600 1092.390 ;
        RECT -14.680 1089.380 0.300 1092.380 ;
        RECT 2919.700 1089.380 2934.300 1092.380 ;
        RECT -9.980 1089.370 -6.980 1089.380 ;
        RECT 2926.600 1089.370 2929.600 1089.380 ;
        RECT -9.980 912.380 -6.980 912.390 ;
        RECT 2926.600 912.380 2929.600 912.390 ;
        RECT -14.680 909.380 0.300 912.380 ;
        RECT 2919.700 909.380 2934.300 912.380 ;
        RECT -9.980 909.370 -6.980 909.380 ;
        RECT 2926.600 909.370 2929.600 909.380 ;
        RECT -9.980 732.380 -6.980 732.390 ;
        RECT 2926.600 732.380 2929.600 732.390 ;
        RECT -14.680 729.380 0.300 732.380 ;
        RECT 2919.700 729.380 2934.300 732.380 ;
        RECT -9.980 729.370 -6.980 729.380 ;
        RECT 2926.600 729.370 2929.600 729.380 ;
        RECT -9.980 552.380 -6.980 552.390 ;
        RECT 2926.600 552.380 2929.600 552.390 ;
        RECT -14.680 549.380 0.300 552.380 ;
        RECT 2919.700 549.380 2934.300 552.380 ;
        RECT -9.980 549.370 -6.980 549.380 ;
        RECT 2926.600 549.370 2929.600 549.380 ;
        RECT -9.980 372.380 -6.980 372.390 ;
        RECT 2926.600 372.380 2929.600 372.390 ;
        RECT -14.680 369.380 0.300 372.380 ;
        RECT 2919.700 369.380 2934.300 372.380 ;
        RECT -9.980 369.370 -6.980 369.380 ;
        RECT 2926.600 369.370 2929.600 369.380 ;
        RECT -9.980 192.380 -6.980 192.390 ;
        RECT 2926.600 192.380 2929.600 192.390 ;
        RECT -14.680 189.380 0.300 192.380 ;
        RECT 2919.700 189.380 2934.300 192.380 ;
        RECT -9.980 189.370 -6.980 189.380 ;
        RECT 2926.600 189.370 2929.600 189.380 ;
        RECT -9.980 12.380 -6.980 12.390 ;
        RECT 2926.600 12.380 2929.600 12.390 ;
        RECT -14.680 9.380 0.300 12.380 ;
        RECT 2919.700 9.380 2934.300 12.380 ;
        RECT -9.980 9.370 -6.980 9.380 ;
        RECT 2926.600 9.370 2929.600 9.380 ;
        RECT -9.980 -1.620 -6.980 -1.610 ;
        RECT 4.020 -1.620 7.020 -1.610 ;
        RECT 184.020 -1.620 187.020 -1.610 ;
        RECT 364.020 -1.620 367.020 -1.610 ;
        RECT 544.020 -1.620 547.020 -1.610 ;
        RECT 724.020 -1.620 727.020 -1.610 ;
        RECT 904.020 -1.620 907.020 -1.610 ;
        RECT 1084.020 -1.620 1087.020 -1.610 ;
        RECT 1264.020 -1.620 1267.020 -1.610 ;
        RECT 1444.020 -1.620 1447.020 -1.610 ;
        RECT 1624.020 -1.620 1627.020 -1.610 ;
        RECT 1804.020 -1.620 1807.020 -1.610 ;
        RECT 1984.020 -1.620 1987.020 -1.610 ;
        RECT 2164.020 -1.620 2167.020 -1.610 ;
        RECT 2344.020 -1.620 2347.020 -1.610 ;
        RECT 2524.020 -1.620 2527.020 -1.610 ;
        RECT 2704.020 -1.620 2707.020 -1.610 ;
        RECT 2884.020 -1.620 2887.020 -1.610 ;
        RECT 2926.600 -1.620 2929.600 -1.610 ;
        RECT -9.980 -4.620 2929.600 -1.620 ;
        RECT -9.980 -4.630 -6.980 -4.620 ;
        RECT 4.020 -4.630 7.020 -4.620 ;
        RECT 184.020 -4.630 187.020 -4.620 ;
        RECT 364.020 -4.630 367.020 -4.620 ;
        RECT 544.020 -4.630 547.020 -4.620 ;
        RECT 724.020 -4.630 727.020 -4.620 ;
        RECT 904.020 -4.630 907.020 -4.620 ;
        RECT 1084.020 -4.630 1087.020 -4.620 ;
        RECT 1264.020 -4.630 1267.020 -4.620 ;
        RECT 1444.020 -4.630 1447.020 -4.620 ;
        RECT 1624.020 -4.630 1627.020 -4.620 ;
        RECT 1804.020 -4.630 1807.020 -4.620 ;
        RECT 1984.020 -4.630 1987.020 -4.620 ;
        RECT 2164.020 -4.630 2167.020 -4.620 ;
        RECT 2344.020 -4.630 2347.020 -4.620 ;
        RECT 2524.020 -4.630 2527.020 -4.620 ;
        RECT 2704.020 -4.630 2707.020 -4.620 ;
        RECT 2884.020 -4.630 2887.020 -4.620 ;
        RECT 2926.600 -4.630 2929.600 -4.620 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -14.680 -9.320 -11.680 3529.000 ;
        RECT 94.020 3519.700 97.020 3529.000 ;
        RECT 274.020 3519.700 277.020 3529.000 ;
        RECT 454.020 3519.700 457.020 3529.000 ;
        RECT 634.020 3519.700 637.020 3529.000 ;
        RECT 814.020 3519.700 817.020 3529.000 ;
        RECT 994.020 3519.700 997.020 3529.000 ;
        RECT 1174.020 3519.700 1177.020 3529.000 ;
        RECT 1354.020 3519.700 1357.020 3529.000 ;
        RECT 1534.020 3519.700 1537.020 3529.000 ;
        RECT 1714.020 3519.700 1717.020 3529.000 ;
        RECT 1894.020 3519.700 1897.020 3529.000 ;
        RECT 2074.020 3519.700 2077.020 3529.000 ;
        RECT 2254.020 3519.700 2257.020 3529.000 ;
        RECT 2434.020 3519.700 2437.020 3529.000 ;
        RECT 2614.020 3519.700 2617.020 3529.000 ;
        RECT 2794.020 3519.700 2797.020 3529.000 ;
        RECT 94.020 -9.320 97.020 0.300 ;
        RECT 274.020 -9.320 277.020 0.300 ;
        RECT 454.020 -9.320 457.020 0.300 ;
        RECT 634.020 -9.320 637.020 0.300 ;
        RECT 814.020 -9.320 817.020 0.300 ;
        RECT 994.020 -9.320 997.020 0.300 ;
        RECT 1174.020 -9.320 1177.020 0.300 ;
        RECT 1354.020 -9.320 1357.020 0.300 ;
        RECT 1534.020 -9.320 1537.020 0.300 ;
        RECT 1714.020 -9.320 1717.020 0.300 ;
        RECT 1894.020 -9.320 1897.020 0.300 ;
        RECT 2074.020 -9.320 2077.020 0.300 ;
        RECT 2254.020 -9.320 2257.020 0.300 ;
        RECT 2434.020 -9.320 2437.020 0.300 ;
        RECT 2614.020 -9.320 2617.020 0.300 ;
        RECT 2794.020 -9.320 2797.020 0.300 ;
        RECT 2931.300 -9.320 2934.300 3529.000 ;
      LAYER via4 ;
        RECT -13.770 3527.710 -12.590 3528.890 ;
        RECT -13.770 3526.110 -12.590 3527.290 ;
        RECT 94.930 3527.710 96.110 3528.890 ;
        RECT 94.930 3526.110 96.110 3527.290 ;
        RECT 274.930 3527.710 276.110 3528.890 ;
        RECT 274.930 3526.110 276.110 3527.290 ;
        RECT 454.930 3527.710 456.110 3528.890 ;
        RECT 454.930 3526.110 456.110 3527.290 ;
        RECT 634.930 3527.710 636.110 3528.890 ;
        RECT 634.930 3526.110 636.110 3527.290 ;
        RECT 814.930 3527.710 816.110 3528.890 ;
        RECT 814.930 3526.110 816.110 3527.290 ;
        RECT 994.930 3527.710 996.110 3528.890 ;
        RECT 994.930 3526.110 996.110 3527.290 ;
        RECT 1174.930 3527.710 1176.110 3528.890 ;
        RECT 1174.930 3526.110 1176.110 3527.290 ;
        RECT 1354.930 3527.710 1356.110 3528.890 ;
        RECT 1354.930 3526.110 1356.110 3527.290 ;
        RECT 1534.930 3527.710 1536.110 3528.890 ;
        RECT 1534.930 3526.110 1536.110 3527.290 ;
        RECT 1714.930 3527.710 1716.110 3528.890 ;
        RECT 1714.930 3526.110 1716.110 3527.290 ;
        RECT 1894.930 3527.710 1896.110 3528.890 ;
        RECT 1894.930 3526.110 1896.110 3527.290 ;
        RECT 2074.930 3527.710 2076.110 3528.890 ;
        RECT 2074.930 3526.110 2076.110 3527.290 ;
        RECT 2254.930 3527.710 2256.110 3528.890 ;
        RECT 2254.930 3526.110 2256.110 3527.290 ;
        RECT 2434.930 3527.710 2436.110 3528.890 ;
        RECT 2434.930 3526.110 2436.110 3527.290 ;
        RECT 2614.930 3527.710 2616.110 3528.890 ;
        RECT 2614.930 3526.110 2616.110 3527.290 ;
        RECT 2794.930 3527.710 2796.110 3528.890 ;
        RECT 2794.930 3526.110 2796.110 3527.290 ;
        RECT 2932.210 3527.710 2933.390 3528.890 ;
        RECT 2932.210 3526.110 2933.390 3527.290 ;
        RECT -13.770 3341.090 -12.590 3342.270 ;
        RECT -13.770 3339.490 -12.590 3340.670 ;
        RECT -13.770 3161.090 -12.590 3162.270 ;
        RECT -13.770 3159.490 -12.590 3160.670 ;
        RECT -13.770 2981.090 -12.590 2982.270 ;
        RECT -13.770 2979.490 -12.590 2980.670 ;
        RECT -13.770 2801.090 -12.590 2802.270 ;
        RECT -13.770 2799.490 -12.590 2800.670 ;
        RECT -13.770 2621.090 -12.590 2622.270 ;
        RECT -13.770 2619.490 -12.590 2620.670 ;
        RECT -13.770 2441.090 -12.590 2442.270 ;
        RECT -13.770 2439.490 -12.590 2440.670 ;
        RECT -13.770 2261.090 -12.590 2262.270 ;
        RECT -13.770 2259.490 -12.590 2260.670 ;
        RECT -13.770 2081.090 -12.590 2082.270 ;
        RECT -13.770 2079.490 -12.590 2080.670 ;
        RECT -13.770 1901.090 -12.590 1902.270 ;
        RECT -13.770 1899.490 -12.590 1900.670 ;
        RECT -13.770 1721.090 -12.590 1722.270 ;
        RECT -13.770 1719.490 -12.590 1720.670 ;
        RECT -13.770 1541.090 -12.590 1542.270 ;
        RECT -13.770 1539.490 -12.590 1540.670 ;
        RECT -13.770 1361.090 -12.590 1362.270 ;
        RECT -13.770 1359.490 -12.590 1360.670 ;
        RECT -13.770 1181.090 -12.590 1182.270 ;
        RECT -13.770 1179.490 -12.590 1180.670 ;
        RECT -13.770 1001.090 -12.590 1002.270 ;
        RECT -13.770 999.490 -12.590 1000.670 ;
        RECT -13.770 821.090 -12.590 822.270 ;
        RECT -13.770 819.490 -12.590 820.670 ;
        RECT -13.770 641.090 -12.590 642.270 ;
        RECT -13.770 639.490 -12.590 640.670 ;
        RECT -13.770 461.090 -12.590 462.270 ;
        RECT -13.770 459.490 -12.590 460.670 ;
        RECT -13.770 281.090 -12.590 282.270 ;
        RECT -13.770 279.490 -12.590 280.670 ;
        RECT -13.770 101.090 -12.590 102.270 ;
        RECT -13.770 99.490 -12.590 100.670 ;
        RECT 2932.210 3341.090 2933.390 3342.270 ;
        RECT 2932.210 3339.490 2933.390 3340.670 ;
        RECT 2932.210 3161.090 2933.390 3162.270 ;
        RECT 2932.210 3159.490 2933.390 3160.670 ;
        RECT 2932.210 2981.090 2933.390 2982.270 ;
        RECT 2932.210 2979.490 2933.390 2980.670 ;
        RECT 2932.210 2801.090 2933.390 2802.270 ;
        RECT 2932.210 2799.490 2933.390 2800.670 ;
        RECT 2932.210 2621.090 2933.390 2622.270 ;
        RECT 2932.210 2619.490 2933.390 2620.670 ;
        RECT 2932.210 2441.090 2933.390 2442.270 ;
        RECT 2932.210 2439.490 2933.390 2440.670 ;
        RECT 2932.210 2261.090 2933.390 2262.270 ;
        RECT 2932.210 2259.490 2933.390 2260.670 ;
        RECT 2932.210 2081.090 2933.390 2082.270 ;
        RECT 2932.210 2079.490 2933.390 2080.670 ;
        RECT 2932.210 1901.090 2933.390 1902.270 ;
        RECT 2932.210 1899.490 2933.390 1900.670 ;
        RECT 2932.210 1721.090 2933.390 1722.270 ;
        RECT 2932.210 1719.490 2933.390 1720.670 ;
        RECT 2932.210 1541.090 2933.390 1542.270 ;
        RECT 2932.210 1539.490 2933.390 1540.670 ;
        RECT 2932.210 1361.090 2933.390 1362.270 ;
        RECT 2932.210 1359.490 2933.390 1360.670 ;
        RECT 2932.210 1181.090 2933.390 1182.270 ;
        RECT 2932.210 1179.490 2933.390 1180.670 ;
        RECT 2932.210 1001.090 2933.390 1002.270 ;
        RECT 2932.210 999.490 2933.390 1000.670 ;
        RECT 2932.210 821.090 2933.390 822.270 ;
        RECT 2932.210 819.490 2933.390 820.670 ;
        RECT 2932.210 641.090 2933.390 642.270 ;
        RECT 2932.210 639.490 2933.390 640.670 ;
        RECT 2932.210 461.090 2933.390 462.270 ;
        RECT 2932.210 459.490 2933.390 460.670 ;
        RECT 2932.210 281.090 2933.390 282.270 ;
        RECT 2932.210 279.490 2933.390 280.670 ;
        RECT 2932.210 101.090 2933.390 102.270 ;
        RECT 2932.210 99.490 2933.390 100.670 ;
        RECT -13.770 -7.610 -12.590 -6.430 ;
        RECT -13.770 -9.210 -12.590 -8.030 ;
        RECT 94.930 -7.610 96.110 -6.430 ;
        RECT 94.930 -9.210 96.110 -8.030 ;
        RECT 274.930 -7.610 276.110 -6.430 ;
        RECT 274.930 -9.210 276.110 -8.030 ;
        RECT 454.930 -7.610 456.110 -6.430 ;
        RECT 454.930 -9.210 456.110 -8.030 ;
        RECT 634.930 -7.610 636.110 -6.430 ;
        RECT 634.930 -9.210 636.110 -8.030 ;
        RECT 814.930 -7.610 816.110 -6.430 ;
        RECT 814.930 -9.210 816.110 -8.030 ;
        RECT 994.930 -7.610 996.110 -6.430 ;
        RECT 994.930 -9.210 996.110 -8.030 ;
        RECT 1174.930 -7.610 1176.110 -6.430 ;
        RECT 1174.930 -9.210 1176.110 -8.030 ;
        RECT 1354.930 -7.610 1356.110 -6.430 ;
        RECT 1354.930 -9.210 1356.110 -8.030 ;
        RECT 1534.930 -7.610 1536.110 -6.430 ;
        RECT 1534.930 -9.210 1536.110 -8.030 ;
        RECT 1714.930 -7.610 1716.110 -6.430 ;
        RECT 1714.930 -9.210 1716.110 -8.030 ;
        RECT 1894.930 -7.610 1896.110 -6.430 ;
        RECT 1894.930 -9.210 1896.110 -8.030 ;
        RECT 2074.930 -7.610 2076.110 -6.430 ;
        RECT 2074.930 -9.210 2076.110 -8.030 ;
        RECT 2254.930 -7.610 2256.110 -6.430 ;
        RECT 2254.930 -9.210 2256.110 -8.030 ;
        RECT 2434.930 -7.610 2436.110 -6.430 ;
        RECT 2434.930 -9.210 2436.110 -8.030 ;
        RECT 2614.930 -7.610 2616.110 -6.430 ;
        RECT 2614.930 -9.210 2616.110 -8.030 ;
        RECT 2794.930 -7.610 2796.110 -6.430 ;
        RECT 2794.930 -9.210 2796.110 -8.030 ;
        RECT 2932.210 -7.610 2933.390 -6.430 ;
        RECT 2932.210 -9.210 2933.390 -8.030 ;
      LAYER met5 ;
        RECT -14.680 3529.000 -11.680 3529.010 ;
        RECT 94.020 3529.000 97.020 3529.010 ;
        RECT 274.020 3529.000 277.020 3529.010 ;
        RECT 454.020 3529.000 457.020 3529.010 ;
        RECT 634.020 3529.000 637.020 3529.010 ;
        RECT 814.020 3529.000 817.020 3529.010 ;
        RECT 994.020 3529.000 997.020 3529.010 ;
        RECT 1174.020 3529.000 1177.020 3529.010 ;
        RECT 1354.020 3529.000 1357.020 3529.010 ;
        RECT 1534.020 3529.000 1537.020 3529.010 ;
        RECT 1714.020 3529.000 1717.020 3529.010 ;
        RECT 1894.020 3529.000 1897.020 3529.010 ;
        RECT 2074.020 3529.000 2077.020 3529.010 ;
        RECT 2254.020 3529.000 2257.020 3529.010 ;
        RECT 2434.020 3529.000 2437.020 3529.010 ;
        RECT 2614.020 3529.000 2617.020 3529.010 ;
        RECT 2794.020 3529.000 2797.020 3529.010 ;
        RECT 2931.300 3529.000 2934.300 3529.010 ;
        RECT -14.680 3526.000 2934.300 3529.000 ;
        RECT -14.680 3525.990 -11.680 3526.000 ;
        RECT 94.020 3525.990 97.020 3526.000 ;
        RECT 274.020 3525.990 277.020 3526.000 ;
        RECT 454.020 3525.990 457.020 3526.000 ;
        RECT 634.020 3525.990 637.020 3526.000 ;
        RECT 814.020 3525.990 817.020 3526.000 ;
        RECT 994.020 3525.990 997.020 3526.000 ;
        RECT 1174.020 3525.990 1177.020 3526.000 ;
        RECT 1354.020 3525.990 1357.020 3526.000 ;
        RECT 1534.020 3525.990 1537.020 3526.000 ;
        RECT 1714.020 3525.990 1717.020 3526.000 ;
        RECT 1894.020 3525.990 1897.020 3526.000 ;
        RECT 2074.020 3525.990 2077.020 3526.000 ;
        RECT 2254.020 3525.990 2257.020 3526.000 ;
        RECT 2434.020 3525.990 2437.020 3526.000 ;
        RECT 2614.020 3525.990 2617.020 3526.000 ;
        RECT 2794.020 3525.990 2797.020 3526.000 ;
        RECT 2931.300 3525.990 2934.300 3526.000 ;
        RECT -14.680 3342.380 -11.680 3342.390 ;
        RECT 2931.300 3342.380 2934.300 3342.390 ;
        RECT -14.680 3339.380 0.300 3342.380 ;
        RECT 2919.700 3339.380 2934.300 3342.380 ;
        RECT -14.680 3339.370 -11.680 3339.380 ;
        RECT 2931.300 3339.370 2934.300 3339.380 ;
        RECT -14.680 3162.380 -11.680 3162.390 ;
        RECT 2931.300 3162.380 2934.300 3162.390 ;
        RECT -14.680 3159.380 0.300 3162.380 ;
        RECT 2919.700 3159.380 2934.300 3162.380 ;
        RECT -14.680 3159.370 -11.680 3159.380 ;
        RECT 2931.300 3159.370 2934.300 3159.380 ;
        RECT -14.680 2982.380 -11.680 2982.390 ;
        RECT 2931.300 2982.380 2934.300 2982.390 ;
        RECT -14.680 2979.380 0.300 2982.380 ;
        RECT 2919.700 2979.380 2934.300 2982.380 ;
        RECT -14.680 2979.370 -11.680 2979.380 ;
        RECT 2931.300 2979.370 2934.300 2979.380 ;
        RECT -14.680 2802.380 -11.680 2802.390 ;
        RECT 2931.300 2802.380 2934.300 2802.390 ;
        RECT -14.680 2799.380 0.300 2802.380 ;
        RECT 2919.700 2799.380 2934.300 2802.380 ;
        RECT -14.680 2799.370 -11.680 2799.380 ;
        RECT 2931.300 2799.370 2934.300 2799.380 ;
        RECT -14.680 2622.380 -11.680 2622.390 ;
        RECT 2931.300 2622.380 2934.300 2622.390 ;
        RECT -14.680 2619.380 0.300 2622.380 ;
        RECT 2919.700 2619.380 2934.300 2622.380 ;
        RECT -14.680 2619.370 -11.680 2619.380 ;
        RECT 2931.300 2619.370 2934.300 2619.380 ;
        RECT -14.680 2442.380 -11.680 2442.390 ;
        RECT 2931.300 2442.380 2934.300 2442.390 ;
        RECT -14.680 2439.380 0.300 2442.380 ;
        RECT 2919.700 2439.380 2934.300 2442.380 ;
        RECT -14.680 2439.370 -11.680 2439.380 ;
        RECT 2931.300 2439.370 2934.300 2439.380 ;
        RECT -14.680 2262.380 -11.680 2262.390 ;
        RECT 2931.300 2262.380 2934.300 2262.390 ;
        RECT -14.680 2259.380 0.300 2262.380 ;
        RECT 2919.700 2259.380 2934.300 2262.380 ;
        RECT -14.680 2259.370 -11.680 2259.380 ;
        RECT 2931.300 2259.370 2934.300 2259.380 ;
        RECT -14.680 2082.380 -11.680 2082.390 ;
        RECT 2931.300 2082.380 2934.300 2082.390 ;
        RECT -14.680 2079.380 0.300 2082.380 ;
        RECT 2919.700 2079.380 2934.300 2082.380 ;
        RECT -14.680 2079.370 -11.680 2079.380 ;
        RECT 2931.300 2079.370 2934.300 2079.380 ;
        RECT -14.680 1902.380 -11.680 1902.390 ;
        RECT 2931.300 1902.380 2934.300 1902.390 ;
        RECT -14.680 1899.380 0.300 1902.380 ;
        RECT 2919.700 1899.380 2934.300 1902.380 ;
        RECT -14.680 1899.370 -11.680 1899.380 ;
        RECT 2931.300 1899.370 2934.300 1899.380 ;
        RECT -14.680 1722.380 -11.680 1722.390 ;
        RECT 2931.300 1722.380 2934.300 1722.390 ;
        RECT -14.680 1719.380 0.300 1722.380 ;
        RECT 2919.700 1719.380 2934.300 1722.380 ;
        RECT -14.680 1719.370 -11.680 1719.380 ;
        RECT 2931.300 1719.370 2934.300 1719.380 ;
        RECT -14.680 1542.380 -11.680 1542.390 ;
        RECT 2931.300 1542.380 2934.300 1542.390 ;
        RECT -14.680 1539.380 0.300 1542.380 ;
        RECT 2919.700 1539.380 2934.300 1542.380 ;
        RECT -14.680 1539.370 -11.680 1539.380 ;
        RECT 2931.300 1539.370 2934.300 1539.380 ;
        RECT -14.680 1362.380 -11.680 1362.390 ;
        RECT 2931.300 1362.380 2934.300 1362.390 ;
        RECT -14.680 1359.380 0.300 1362.380 ;
        RECT 2919.700 1359.380 2934.300 1362.380 ;
        RECT -14.680 1359.370 -11.680 1359.380 ;
        RECT 2931.300 1359.370 2934.300 1359.380 ;
        RECT -14.680 1182.380 -11.680 1182.390 ;
        RECT 2931.300 1182.380 2934.300 1182.390 ;
        RECT -14.680 1179.380 0.300 1182.380 ;
        RECT 2919.700 1179.380 2934.300 1182.380 ;
        RECT -14.680 1179.370 -11.680 1179.380 ;
        RECT 2931.300 1179.370 2934.300 1179.380 ;
        RECT -14.680 1002.380 -11.680 1002.390 ;
        RECT 2931.300 1002.380 2934.300 1002.390 ;
        RECT -14.680 999.380 0.300 1002.380 ;
        RECT 2919.700 999.380 2934.300 1002.380 ;
        RECT -14.680 999.370 -11.680 999.380 ;
        RECT 2931.300 999.370 2934.300 999.380 ;
        RECT -14.680 822.380 -11.680 822.390 ;
        RECT 2931.300 822.380 2934.300 822.390 ;
        RECT -14.680 819.380 0.300 822.380 ;
        RECT 2919.700 819.380 2934.300 822.380 ;
        RECT -14.680 819.370 -11.680 819.380 ;
        RECT 2931.300 819.370 2934.300 819.380 ;
        RECT -14.680 642.380 -11.680 642.390 ;
        RECT 2931.300 642.380 2934.300 642.390 ;
        RECT -14.680 639.380 0.300 642.380 ;
        RECT 2919.700 639.380 2934.300 642.380 ;
        RECT -14.680 639.370 -11.680 639.380 ;
        RECT 2931.300 639.370 2934.300 639.380 ;
        RECT -14.680 462.380 -11.680 462.390 ;
        RECT 2931.300 462.380 2934.300 462.390 ;
        RECT -14.680 459.380 0.300 462.380 ;
        RECT 2919.700 459.380 2934.300 462.380 ;
        RECT -14.680 459.370 -11.680 459.380 ;
        RECT 2931.300 459.370 2934.300 459.380 ;
        RECT -14.680 282.380 -11.680 282.390 ;
        RECT 2931.300 282.380 2934.300 282.390 ;
        RECT -14.680 279.380 0.300 282.380 ;
        RECT 2919.700 279.380 2934.300 282.380 ;
        RECT -14.680 279.370 -11.680 279.380 ;
        RECT 2931.300 279.370 2934.300 279.380 ;
        RECT -14.680 102.380 -11.680 102.390 ;
        RECT 2931.300 102.380 2934.300 102.390 ;
        RECT -14.680 99.380 0.300 102.380 ;
        RECT 2919.700 99.380 2934.300 102.380 ;
        RECT -14.680 99.370 -11.680 99.380 ;
        RECT 2931.300 99.370 2934.300 99.380 ;
        RECT -14.680 -6.320 -11.680 -6.310 ;
        RECT 94.020 -6.320 97.020 -6.310 ;
        RECT 274.020 -6.320 277.020 -6.310 ;
        RECT 454.020 -6.320 457.020 -6.310 ;
        RECT 634.020 -6.320 637.020 -6.310 ;
        RECT 814.020 -6.320 817.020 -6.310 ;
        RECT 994.020 -6.320 997.020 -6.310 ;
        RECT 1174.020 -6.320 1177.020 -6.310 ;
        RECT 1354.020 -6.320 1357.020 -6.310 ;
        RECT 1534.020 -6.320 1537.020 -6.310 ;
        RECT 1714.020 -6.320 1717.020 -6.310 ;
        RECT 1894.020 -6.320 1897.020 -6.310 ;
        RECT 2074.020 -6.320 2077.020 -6.310 ;
        RECT 2254.020 -6.320 2257.020 -6.310 ;
        RECT 2434.020 -6.320 2437.020 -6.310 ;
        RECT 2614.020 -6.320 2617.020 -6.310 ;
        RECT 2794.020 -6.320 2797.020 -6.310 ;
        RECT 2931.300 -6.320 2934.300 -6.310 ;
        RECT -14.680 -9.320 2934.300 -6.320 ;
        RECT -14.680 -9.330 -11.680 -9.320 ;
        RECT 94.020 -9.330 97.020 -9.320 ;
        RECT 274.020 -9.330 277.020 -9.320 ;
        RECT 454.020 -9.330 457.020 -9.320 ;
        RECT 634.020 -9.330 637.020 -9.320 ;
        RECT 814.020 -9.330 817.020 -9.320 ;
        RECT 994.020 -9.330 997.020 -9.320 ;
        RECT 1174.020 -9.330 1177.020 -9.320 ;
        RECT 1354.020 -9.330 1357.020 -9.320 ;
        RECT 1534.020 -9.330 1537.020 -9.320 ;
        RECT 1714.020 -9.330 1717.020 -9.320 ;
        RECT 1894.020 -9.330 1897.020 -9.320 ;
        RECT 2074.020 -9.330 2077.020 -9.320 ;
        RECT 2254.020 -9.330 2257.020 -9.320 ;
        RECT 2434.020 -9.330 2437.020 -9.320 ;
        RECT 2614.020 -9.330 2617.020 -9.320 ;
        RECT 2794.020 -9.330 2797.020 -9.320 ;
        RECT 2931.300 -9.330 2934.300 -9.320 ;
    END
  END vssd1
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -19.380 -14.020 -16.380 3533.700 ;
        RECT 2936.000 -14.020 2939.000 3533.700 ;
      LAYER via4 ;
        RECT -18.470 3532.410 -17.290 3533.590 ;
        RECT -18.470 3530.810 -17.290 3531.990 ;
        RECT -18.470 -12.310 -17.290 -11.130 ;
        RECT -18.470 -13.910 -17.290 -12.730 ;
        RECT 2936.910 3532.410 2938.090 3533.590 ;
        RECT 2936.910 3530.810 2938.090 3531.990 ;
        RECT 2936.910 -12.310 2938.090 -11.130 ;
        RECT 2936.910 -13.910 2938.090 -12.730 ;
      LAYER met5 ;
        RECT -19.380 3533.700 -16.380 3533.710 ;
        RECT 2936.000 3533.700 2939.000 3533.710 ;
        RECT -19.380 3530.700 2939.000 3533.700 ;
        RECT -19.380 3530.690 -16.380 3530.700 ;
        RECT 2936.000 3530.690 2939.000 3530.700 ;
        RECT -19.380 -11.020 -16.380 -11.010 ;
        RECT 2936.000 -11.020 2939.000 -11.010 ;
        RECT -19.380 -14.020 2939.000 -11.020 ;
        RECT -19.380 -14.030 -16.380 -14.020 ;
        RECT 2936.000 -14.030 2939.000 -14.020 ;
    END
  END vccd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -24.080 -18.720 -21.080 3538.400 ;
        RECT 2940.700 -18.720 2943.700 3538.400 ;
      LAYER via4 ;
        RECT -23.170 3537.110 -21.990 3538.290 ;
        RECT -23.170 3535.510 -21.990 3536.690 ;
        RECT -23.170 -17.010 -21.990 -15.830 ;
        RECT -23.170 -18.610 -21.990 -17.430 ;
        RECT 2941.610 3537.110 2942.790 3538.290 ;
        RECT 2941.610 3535.510 2942.790 3536.690 ;
        RECT 2941.610 -17.010 2942.790 -15.830 ;
        RECT 2941.610 -18.610 2942.790 -17.430 ;
      LAYER met5 ;
        RECT -24.080 3538.400 -21.080 3538.410 ;
        RECT 2940.700 3538.400 2943.700 3538.410 ;
        RECT -24.080 3535.400 2943.700 3538.400 ;
        RECT -24.080 3535.390 -21.080 3535.400 ;
        RECT 2940.700 3535.390 2943.700 3535.400 ;
        RECT -24.080 -15.720 -21.080 -15.710 ;
        RECT 2940.700 -15.720 2943.700 -15.710 ;
        RECT -24.080 -18.720 2943.700 -15.720 ;
        RECT -24.080 -18.730 -21.080 -18.720 ;
        RECT 2940.700 -18.730 2943.700 -18.720 ;
    END
  END vssd2
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -28.780 -23.420 -25.780 3543.100 ;
        RECT 2945.400 -23.420 2948.400 3543.100 ;
      LAYER via4 ;
        RECT -27.870 3541.810 -26.690 3542.990 ;
        RECT -27.870 3540.210 -26.690 3541.390 ;
        RECT -27.870 -21.710 -26.690 -20.530 ;
        RECT -27.870 -23.310 -26.690 -22.130 ;
        RECT 2946.310 3541.810 2947.490 3542.990 ;
        RECT 2946.310 3540.210 2947.490 3541.390 ;
        RECT 2946.310 -21.710 2947.490 -20.530 ;
        RECT 2946.310 -23.310 2947.490 -22.130 ;
      LAYER met5 ;
        RECT -28.780 3543.100 -25.780 3543.110 ;
        RECT 2945.400 3543.100 2948.400 3543.110 ;
        RECT -28.780 3540.100 2948.400 3543.100 ;
        RECT -28.780 3540.090 -25.780 3540.100 ;
        RECT 2945.400 3540.090 2948.400 3540.100 ;
        RECT -28.780 -20.420 -25.780 -20.410 ;
        RECT 2945.400 -20.420 2948.400 -20.410 ;
        RECT -28.780 -23.420 2948.400 -20.420 ;
        RECT -28.780 -23.430 -25.780 -23.420 ;
        RECT 2945.400 -23.430 2948.400 -23.420 ;
    END
  END vdda1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -33.480 -28.120 -30.480 3547.800 ;
        RECT 2950.100 -28.120 2953.100 3547.800 ;
      LAYER via4 ;
        RECT -32.570 3546.510 -31.390 3547.690 ;
        RECT -32.570 3544.910 -31.390 3546.090 ;
        RECT -32.570 -26.410 -31.390 -25.230 ;
        RECT -32.570 -28.010 -31.390 -26.830 ;
        RECT 2951.010 3546.510 2952.190 3547.690 ;
        RECT 2951.010 3544.910 2952.190 3546.090 ;
        RECT 2951.010 -26.410 2952.190 -25.230 ;
        RECT 2951.010 -28.010 2952.190 -26.830 ;
      LAYER met5 ;
        RECT -33.480 3547.800 -30.480 3547.810 ;
        RECT 2950.100 3547.800 2953.100 3547.810 ;
        RECT -33.480 3544.800 2953.100 3547.800 ;
        RECT -33.480 3544.790 -30.480 3544.800 ;
        RECT 2950.100 3544.790 2953.100 3544.800 ;
        RECT -33.480 -25.120 -30.480 -25.110 ;
        RECT 2950.100 -25.120 2953.100 -25.110 ;
        RECT -33.480 -28.120 2953.100 -25.120 ;
        RECT -33.480 -28.130 -30.480 -28.120 ;
        RECT 2950.100 -28.130 2953.100 -28.120 ;
    END
  END vssa1
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -38.180 -32.820 -35.180 3552.500 ;
        RECT 2954.800 -32.820 2957.800 3552.500 ;
      LAYER via4 ;
        RECT -37.270 3551.210 -36.090 3552.390 ;
        RECT -37.270 3549.610 -36.090 3550.790 ;
        RECT -37.270 -31.110 -36.090 -29.930 ;
        RECT -37.270 -32.710 -36.090 -31.530 ;
        RECT 2955.710 3551.210 2956.890 3552.390 ;
        RECT 2955.710 3549.610 2956.890 3550.790 ;
        RECT 2955.710 -31.110 2956.890 -29.930 ;
        RECT 2955.710 -32.710 2956.890 -31.530 ;
      LAYER met5 ;
        RECT -38.180 3552.500 -35.180 3552.510 ;
        RECT 2954.800 3552.500 2957.800 3552.510 ;
        RECT -38.180 3549.500 2957.800 3552.500 ;
        RECT -38.180 3549.490 -35.180 3549.500 ;
        RECT 2954.800 3549.490 2957.800 3549.500 ;
        RECT -38.180 -29.820 -35.180 -29.810 ;
        RECT 2954.800 -29.820 2957.800 -29.810 ;
        RECT -38.180 -32.820 2957.800 -29.820 ;
        RECT -38.180 -32.830 -35.180 -32.820 ;
        RECT 2954.800 -32.830 2957.800 -32.820 ;
    END
  END vdda2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -42.880 -37.520 -39.880 3557.200 ;
        RECT 2959.500 -37.520 2962.500 3557.200 ;
      LAYER via4 ;
        RECT -41.970 3555.910 -40.790 3557.090 ;
        RECT -41.970 3554.310 -40.790 3555.490 ;
        RECT -41.970 -35.810 -40.790 -34.630 ;
        RECT -41.970 -37.410 -40.790 -36.230 ;
        RECT 2960.410 3555.910 2961.590 3557.090 ;
        RECT 2960.410 3554.310 2961.590 3555.490 ;
        RECT 2960.410 -35.810 2961.590 -34.630 ;
        RECT 2960.410 -37.410 2961.590 -36.230 ;
      LAYER met5 ;
        RECT -42.880 3557.200 -39.880 3557.210 ;
        RECT 2959.500 3557.200 2962.500 3557.210 ;
        RECT -42.880 3554.200 2962.500 3557.200 ;
        RECT -42.880 3554.190 -39.880 3554.200 ;
        RECT 2959.500 3554.190 2962.500 3554.200 ;
        RECT -42.880 -34.520 -39.880 -34.510 ;
        RECT 2959.500 -34.520 2962.500 -34.510 ;
        RECT -42.880 -37.520 2962.500 -34.520 ;
        RECT -42.880 -37.530 -39.880 -37.520 ;
        RECT 2959.500 -37.530 2962.500 -37.520 ;
    END
  END vssa2
  OBS
      LAYER li1 ;
        RECT 139.120 380.555 2788.400 2908.785 ;
      LAYER met1 ;
        RECT 14.790 18.060 2917.250 3503.320 ;
      LAYER met2 ;
        RECT 2.710 0.300 2917.370 3519.700 ;
      LAYER met3 ;
        RECT 0.300 28.980 2919.700 3490.700 ;
      LAYER met4 ;
        RECT 4.020 0.300 2887.020 3519.700 ;
      LAYER met5 ;
        RECT 0.300 9.370 2919.700 3432.390 ;
  END
END user_project_wrapper
END LIBRARY


* NGSPICE file created from decred_controller.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_4 abstract view
.subckt sky130_fd_sc_hd__nand4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_4 abstract view
.subckt sky130_fd_sc_hd__and4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_4 abstract view
.subckt sky130_fd_sc_hd__o32ai_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_4 abstract view
.subckt sky130_fd_sc_hd__a211o_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_4 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41oi_4 abstract view
.subckt sky130_fd_sc_hd__a41oi_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_4 abstract view
.subckt sky130_fd_sc_hd__nor4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_4 abstract view
.subckt sky130_fd_sc_hd__a41o_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41ai_4 abstract view
.subckt sky130_fd_sc_hd__o41ai_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2oi_4 abstract view
.subckt sky130_fd_sc_hd__a2bb2oi_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_4 abstract view
.subckt sky130_fd_sc_hd__o41a_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_4 abstract view
.subckt sky130_fd_sc_hd__a32oi_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_4 abstract view
.subckt sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_4 abstract view
.subckt sky130_fd_sc_hd__a21boi_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_4 abstract view
.subckt sky130_fd_sc_hd__a2111o_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

.subckt decred_controller CLK_LED DATA_AVAILABLE[0] DATA_AVAILABLE[1] DATA_AVAILABLE[2]
+ DATA_AVAILABLE[3] DATA_FROM_HASH[0] DATA_FROM_HASH[1] DATA_FROM_HASH[2] DATA_FROM_HASH[3]
+ DATA_FROM_HASH[4] DATA_FROM_HASH[5] DATA_FROM_HASH[6] DATA_FROM_HASH[7] DATA_TO_HASH[0]
+ DATA_TO_HASH[1] DATA_TO_HASH[2] DATA_TO_HASH[3] DATA_TO_HASH[4] DATA_TO_HASH[5]
+ DATA_TO_HASH[6] DATA_TO_HASH[7] EXT_RESET_N_fromHost EXT_RESET_N_toClient HASH_ADDR[0]
+ HASH_ADDR[1] HASH_ADDR[2] HASH_ADDR[3] HASH_ADDR[4] HASH_ADDR[5] HASH_EN HASH_LED
+ ID_fromClient ID_toHost IRQ_OUT_fromClient IRQ_OUT_toHost M1_CLK_IN M1_CLK_SELECT
+ MACRO_RD_SELECT[0] MACRO_RD_SELECT[1] MACRO_RD_SELECT[2] MACRO_RD_SELECT[3] MACRO_WR_SELECT[0]
+ MACRO_WR_SELECT[1] MACRO_WR_SELECT[2] MACRO_WR_SELECT[3] MISO_fromClient MISO_toHost
+ MOSI_fromHost MOSI_toClient PLL_INPUT S1_CLK_IN S1_CLK_SELECT SCLK_fromHost SCLK_toClient
+ SCSN_fromHost SCSN_toClient THREAD_COUNT[0] THREAD_COUNT[1] THREAD_COUNT[2] THREAD_COUNT[3]
+ m1_clk_local one zero vccd1 vssd1 vccd2_uq0 vccd2 vssd2 vdda1_uq0 vdda1 vssa1 vdda2_uq0
+ vdda2 vssa2
XFILLER_54_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2037_ _2032_/C _2047_/A _2043_/D _1995_/B vssd1 vssd1 vccd1 vccd1 _2038_/B sky130_fd_sc_hd__nand4_4
X_2106_ _1222_/A SCSN_fromHost vssd1 vssd1 vccd1 vccd1 _2458_/D sky130_fd_sc_hd__or2_4
XFILLER_18_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1270_ _1346_/A vssd1 vssd1 vccd1 vccd1 _2010_/B sky130_fd_sc_hd__buf_2
XFILLER_36_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1606_ _1589_/A _1567_/C vssd1 vssd1 vccd1 vccd1 _1606_/Y sky130_fd_sc_hd__nor2_4
X_1399_ _1231_/A _1397_/Y _1398_/Y vssd1 vssd1 vccd1 vccd1 _1399_/X sky130_fd_sc_hd__a21o_4
X_1468_ _1428_/Y vssd1 vssd1 vccd1 vccd1 _1548_/D sky130_fd_sc_hd__buf_2
X_1537_ _1424_/Y vssd1 vssd1 vccd1 vccd1 _1556_/B sky130_fd_sc_hd__buf_2
X_2586_ _2446_/CLK _2586_/D vssd1 vssd1 vccd1 vccd1 _2127_/C sky130_fd_sc_hd__dfxtp_4
XFILLER_63_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2440_ _2552_/CLK _2143_/Y vssd1 vssd1 vccd1 vccd1 _2440_/Q sky130_fd_sc_hd__dfxtp_4
X_2371_ _2374_/CLK _2370_/Q vssd1 vssd1 vccd1 vccd1 _2372_/D sky130_fd_sc_hd__dfxtp_4
X_1253_ _2364_/D vssd1 vssd1 vccd1 vccd1 _1269_/A sky130_fd_sc_hd__inv_2
X_1322_ _1239_/Y _1321_/X _1316_/D vssd1 vssd1 vccd1 vccd1 _1322_/Y sky130_fd_sc_hd__nand3_4
Xclkbuf_1_0_0_m1_clk_local clkbuf_0_m1_clk_local/X vssd1 vssd1 vccd1 vccd1 clkbuf_1_0_0_m1_clk_local/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_49_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1184_ _1184_/A vssd1 vssd1 vccd1 vccd1 _1185_/A sky130_fd_sc_hd__buf_2
XFILLER_17_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2569_ _2454_/CLK _2569_/D vssd1 vssd1 vccd1 vccd1 _1830_/C sky130_fd_sc_hd__dfxtp_4
X_2638_ _2635_/CLK _1297_/Y vssd1 vssd1 vccd1 vccd1 _1295_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_59_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1871_ _2112_/A DATA_FROM_HASH[7] vssd1 vssd1 vccd1 vccd1 _2566_/D sky130_fd_sc_hd__and2_4
X_1940_ _1938_/A _1746_/Y vssd1 vssd1 vccd1 vccd1 _1940_/Y sky130_fd_sc_hd__nor2_4
XFILLER_9_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2423_ _2404_/CLK _2423_/D vssd1 vssd1 vccd1 vccd1 _2423_/Q sky130_fd_sc_hd__dfxtp_4
X_1236_ _1376_/B _1236_/B vssd1 vssd1 vccd1 vccd1 _1237_/A sky130_fd_sc_hd__nand2_4
X_2354_ _2097_/B _1202_/B _2353_/X vssd1 vssd1 vccd1 vccd1 _2354_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_37_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1305_ _1318_/B _1308_/C _1243_/X _1305_/D vssd1 vssd1 vccd1 vccd1 _1305_/X sky130_fd_sc_hd__and4_4
Xclkbuf_0_m1_clk_local m1_clk_local vssd1 vssd1 vccd1 vccd1 clkbuf_0_m1_clk_local/X
+ sky130_fd_sc_hd__clkbuf_16
X_2285_ _2276_/X _2253_/Y _2278_/X _1924_/B _2280_/X vssd1 vssd1 vccd1 vccd1 _2414_/D
+ sky130_fd_sc_hd__o32ai_4
XFILLER_64_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2070_ _2070_/A vssd1 vssd1 vccd1 vccd1 _2070_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_3_3_0_m1_clk_local clkbuf_3_3_0_m1_clk_local/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_3_0_m1_clk_local/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_61_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1785_ _1783_/Y _1784_/Y _2100_/A vssd1 vssd1 vccd1 vccd1 _2588_/D sky130_fd_sc_hd__a21oi_4
X_1854_ _1854_/A _1854_/B vssd1 vssd1 vccd1 vccd1 _1854_/X sky130_fd_sc_hd__or2_4
X_1923_ _2151_/B vssd1 vssd1 vccd1 vccd1 _1924_/B sky130_fd_sc_hd__inv_2
X_2406_ _2552_/CLK _2406_/D vssd1 vssd1 vccd1 vccd1 HASH_LED sky130_fd_sc_hd__dfxtp_4
XFILLER_55_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2337_ _1574_/Y _2337_/B _1683_/Y vssd1 vssd1 vccd1 vccd1 _2338_/A sky130_fd_sc_hd__nand3_4
X_1219_ _2384_/Q vssd1 vssd1 vccd1 vccd1 _1219_/X sky130_fd_sc_hd__buf_2
XFILLER_29_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2268_ _1477_/X vssd1 vssd1 vccd1 vccd1 _2268_/Y sky130_fd_sc_hd__inv_2
X_2199_ _1623_/Y _2428_/Q vssd1 vssd1 vccd1 vccd1 _2199_/Y sky130_fd_sc_hd__nand2_4
XFILLER_40_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1570_ _1570_/A vssd1 vssd1 vccd1 vccd1 _1571_/A sky130_fd_sc_hd__buf_2
X_2053_ _1992_/A _1990_/Y _2059_/A vssd1 vssd1 vccd1 vccd1 _2053_/Y sky130_fd_sc_hd__nor3_4
X_2122_ _1886_/A _2121_/X _1420_/A vssd1 vssd1 vccd1 vccd1 _2122_/Y sky130_fd_sc_hd__nand3_4
XFILLER_13_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1837_ _1837_/A vssd1 vssd1 vccd1 vccd1 _2570_/D sky130_fd_sc_hd__inv_2
X_1768_ _1438_/B _2401_/Q vssd1 vssd1 vccd1 vccd1 _1768_/X sky130_fd_sc_hd__xor2_4
X_1906_ _2154_/B vssd1 vssd1 vccd1 vccd1 _1906_/Y sky130_fd_sc_hd__inv_2
X_1699_ _1693_/Y _1698_/Y _1454_/X vssd1 vssd1 vccd1 vccd1 _2594_/D sky130_fd_sc_hd__a21oi_4
XFILLER_1_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1622_ _1622_/A vssd1 vssd1 vccd1 vccd1 _1622_/Y sky130_fd_sc_hd__inv_2
XPHY_181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1553_ _1490_/A _1527_/Y _1564_/A _1552_/Y vssd1 vssd1 vccd1 vccd1 _1557_/A sky130_fd_sc_hd__a211o_4
X_1484_ _1484_/A vssd1 vssd1 vccd1 vccd1 _1487_/B sky130_fd_sc_hd__buf_2
X_2036_ _1995_/B _2035_/X _1374_/X vssd1 vssd1 vccd1 vccd1 _2038_/A sky130_fd_sc_hd__o21a_4
X_2105_ _1222_/A _2105_/B vssd1 vssd1 vccd1 vccd1 _2105_/X sky130_fd_sc_hd__or2_4
XFILLER_39_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1605_ _1605_/A vssd1 vssd1 vccd1 vccd1 _1605_/X sky130_fd_sc_hd__buf_2
X_1536_ _1525_/Y _1532_/Y _1535_/X vssd1 vssd1 vccd1 vccd1 _2604_/D sky130_fd_sc_hd__a21oi_4
X_2585_ _2399_/CLK _1796_/X vssd1 vssd1 vccd1 vccd1 _1477_/A sky130_fd_sc_hd__dfxtp_4
X_1398_ _1231_/A _1397_/Y _1374_/X vssd1 vssd1 vccd1 vccd1 _1398_/Y sky130_fd_sc_hd__o21ai_4
X_1467_ _1467_/A vssd1 vssd1 vccd1 vccd1 _1467_/Y sky130_fd_sc_hd__inv_2
X_2019_ _2019_/A _2019_/B _2019_/C vssd1 vssd1 vccd1 vccd1 _2019_/Y sky130_fd_sc_hd__nor3_4
XFILLER_35_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2370_ _2374_/CLK _2369_/Q vssd1 vssd1 vccd1 vccd1 _2370_/Q sky130_fd_sc_hd__dfxtp_4
X_1321_ _1241_/Y vssd1 vssd1 vccd1 vccd1 _1321_/X sky130_fd_sc_hd__buf_2
X_1252_ _1252_/A _1641_/A vssd1 vssd1 vccd1 vccd1 _1263_/A sky130_fd_sc_hd__nand2_4
XFILLER_1_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1183_ _2353_/A _1179_/X _1182_/X vssd1 vssd1 vccd1 vccd1 _1183_/Y sky130_fd_sc_hd__o21ai_4
Xclkbuf_3_4_0_addressalyzerBlock.SPI_CLK clkbuf_3_5_0_addressalyzerBlock.SPI_CLK/A
+ vssd1 vssd1 vccd1 vccd1 clkbuf_4_9_0_addressalyzerBlock.SPI_CLK/A sky130_fd_sc_hd__clkbuf_1
X_2499_ _2511_/CLK _1971_/X vssd1 vssd1 vccd1 vccd1 MACRO_WR_SELECT[0] sky130_fd_sc_hd__dfxtp_4
X_2568_ _2464_/CLK _1863_/Y vssd1 vssd1 vccd1 vccd1 _1862_/B sky130_fd_sc_hd__dfxtp_4
X_2637_ _2635_/CLK _2637_/D vssd1 vssd1 vccd1 vccd1 _1299_/A sky130_fd_sc_hd__dfxtp_4
X_1519_ _1470_/X _1440_/B _1518_/Y vssd1 vssd1 vccd1 vccd1 _1519_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_55_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1870_ _1840_/B vssd1 vssd1 vccd1 vccd1 _2112_/A sky130_fd_sc_hd__buf_2
X_2353_ _2353_/A _1198_/B vssd1 vssd1 vccd1 vccd1 _2353_/X sky130_fd_sc_hd__or2_4
XFILLER_43_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2422_ _2404_/CLK _2422_/D vssd1 vssd1 vccd1 vccd1 _2155_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_56_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1235_ _1234_/Y vssd1 vssd1 vccd1 vccd1 _1365_/D sky130_fd_sc_hd__inv_2
XFILLER_37_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1304_ _2635_/Q vssd1 vssd1 vccd1 vccd1 _1308_/C sky130_fd_sc_hd__buf_2
X_2284_ _2276_/X _2133_/Y _2278_/X _1744_/B _2280_/X vssd1 vssd1 vccd1 vccd1 _2284_/Y
+ sky130_fd_sc_hd__o32ai_4
X_1999_ _1999_/A _1998_/Y _2011_/A _2492_/Q vssd1 vssd1 vccd1 vccd1 _2010_/C sky130_fd_sc_hd__nand4_4
XFILLER_20_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1922_ _1933_/A _2537_/Q vssd1 vssd1 vccd1 vccd1 _2531_/D sky130_fd_sc_hd__and2_4
X_1784_ _1678_/Y _2349_/A vssd1 vssd1 vccd1 vccd1 _1784_/Y sky130_fd_sc_hd__nand2_4
X_1853_ _1850_/X _1852_/X _1472_/A vssd1 vssd1 vccd1 vccd1 _1853_/Y sky130_fd_sc_hd__a21oi_4
X_2336_ _2337_/B _2328_/X _2335_/Y vssd1 vssd1 vccd1 vccd1 _2388_/D sky130_fd_sc_hd__o21ai_4
XFILLER_29_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2405_ _2552_/CLK _2305_/Y vssd1 vssd1 vccd1 vccd1 _1232_/A sky130_fd_sc_hd__dfxtp_4
X_1218_ _1218_/A _1218_/B vssd1 vssd1 vccd1 vccd1 _1218_/Y sky130_fd_sc_hd__nand2_4
X_2267_ _2266_/Y _2262_/X _2258_/X _1937_/Y _2264_/X vssd1 vssd1 vccd1 vccd1 _2425_/D
+ sky130_fd_sc_hd__o32ai_4
X_2198_ _2196_/Y _1708_/X _2198_/C vssd1 vssd1 vccd1 vccd1 _2198_/Y sky130_fd_sc_hd__nand3_4
XFILLER_4_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2052_ _2014_/X _2040_/X _2051_/Y vssd1 vssd1 vccd1 vccd1 _2482_/D sky130_fd_sc_hd__a21oi_4
XFILLER_54_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2121_ _1696_/A vssd1 vssd1 vccd1 vccd1 _2121_/X sky130_fd_sc_hd__buf_2
XFILLER_34_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1905_ _1911_/A _1904_/Y vssd1 vssd1 vccd1 vccd1 _1905_/Y sky130_fd_sc_hd__nor2_4
XFILLER_22_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1836_ _1830_/B _1834_/Y _1835_/Y vssd1 vssd1 vccd1 vccd1 _1837_/A sky130_fd_sc_hd__a21o_4
X_1698_ _1698_/A _1697_/Y _1689_/Y _1687_/Y vssd1 vssd1 vccd1 vccd1 _1698_/Y sky130_fd_sc_hd__nand4_4
XFILLER_30_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1767_ _1483_/B _1767_/B vssd1 vssd1 vccd1 vccd1 _1767_/X sky130_fd_sc_hd__xor2_4
X_2319_ _1771_/Y _2310_/X _1503_/A _2312_/X vssd1 vssd1 vccd1 vccd1 _2319_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_65_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1552_ _1556_/B _1548_/D _1544_/Y vssd1 vssd1 vccd1 vccd1 _1552_/Y sky130_fd_sc_hd__a21oi_4
X_1621_ _2293_/C _2181_/A _1704_/A _1620_/Y vssd1 vssd1 vccd1 vccd1 _1621_/X sky130_fd_sc_hd__a211o_4
X_2104_ _2104_/A _2091_/Y _2103_/Y _2104_/D vssd1 vssd1 vccd1 vccd1 _2460_/D sky130_fd_sc_hd__and4_4
X_1483_ _1482_/Y _1483_/B _2604_/Q _1483_/D vssd1 vssd1 vccd1 vccd1 _1484_/A sky130_fd_sc_hd__and4_4
X_2035_ _2029_/Y _2030_/X _2016_/X _2043_/D vssd1 vssd1 vccd1 vccd1 _2035_/X sky130_fd_sc_hd__and4_4
X_1819_ _2575_/Q _1809_/X _1818_/X vssd1 vssd1 vccd1 vccd1 _2576_/D sky130_fd_sc_hd__o21a_4
XFILLER_45_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1604_ _1604_/A _2600_/Q vssd1 vssd1 vccd1 vccd1 _1605_/A sky130_fd_sc_hd__and2_4
X_2584_ _2399_/CLK _1798_/X vssd1 vssd1 vccd1 vccd1 _1490_/A sky130_fd_sc_hd__dfxtp_4
X_1535_ _1556_/A _1534_/X _1500_/X vssd1 vssd1 vccd1 vccd1 _1535_/X sky130_fd_sc_hd__a21o_4
X_1397_ _1397_/A _1363_/A _1363_/C vssd1 vssd1 vccd1 vccd1 _1397_/Y sky130_fd_sc_hd__nor3_4
XFILLER_27_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1466_ _1466_/A vssd1 vssd1 vccd1 vccd1 _1469_/A sky130_fd_sc_hd__inv_2
X_2018_ _2488_/Q _2017_/X _1984_/A _1999_/A _2011_/A vssd1 vssd1 vccd1 vccd1 _2019_/C
+ sky130_fd_sc_hd__a41oi_4
XFILLER_50_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1320_ _1320_/A vssd1 vssd1 vccd1 vccd1 _1320_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1182_ _2650_/Q _1194_/B vssd1 vssd1 vccd1 vccd1 _1182_/X sky130_fd_sc_hd__or2_4
X_1251_ _1251_/A vssd1 vssd1 vccd1 vccd1 _1641_/A sky130_fd_sc_hd__inv_2
XFILLER_32_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2636_ _2476_/CLK _2636_/D vssd1 vssd1 vccd1 vccd1 _2636_/Q sky130_fd_sc_hd__dfxtp_4
X_2498_ _2508_/CLK _1975_/Y vssd1 vssd1 vccd1 vccd1 _1973_/A sky130_fd_sc_hd__dfxtp_4
X_2567_ _2374_/CLK _2567_/D vssd1 vssd1 vccd1 vccd1 _1868_/A sky130_fd_sc_hd__dfxtp_4
X_1449_ _1441_/Y _1449_/B vssd1 vssd1 vccd1 vccd1 _1449_/Y sky130_fd_sc_hd__nand2_4
X_1518_ _1470_/X _1482_/Y _1473_/C _1466_/A _2340_/C vssd1 vssd1 vccd1 vccd1 _1518_/Y
+ sky130_fd_sc_hd__a41oi_4
XFILLER_23_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2352_ _2543_/Q _2544_/Q _2352_/C vssd1 vssd1 vccd1 vccd1 IRQ_OUT_toHost sky130_fd_sc_hd__or3_4
XFILLER_36_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1303_ _1258_/Y vssd1 vssd1 vccd1 vccd1 _1318_/B sky130_fd_sc_hd__buf_2
X_2283_ _2276_/X _2130_/Y _2278_/X _1845_/B _2280_/X vssd1 vssd1 vccd1 vccd1 _2416_/D
+ sky130_fd_sc_hd__o32ai_4
X_2421_ _2551_/CLK _2273_/Y vssd1 vssd1 vccd1 vccd1 _2421_/Q sky130_fd_sc_hd__dfxtp_4
X_1234_ _2622_/Q _2621_/Q vssd1 vssd1 vccd1 vccd1 _1234_/Y sky130_fd_sc_hd__nand2_4
XFILLER_52_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1998_ _2002_/A _2008_/A vssd1 vssd1 vccd1 vccd1 _1998_/Y sky130_fd_sc_hd__nor2_4
X_2619_ _2619_/CLK _1395_/Y vssd1 vssd1 vccd1 vccd1 _2619_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1921_ _1254_/X vssd1 vssd1 vccd1 vccd1 _1933_/A sky130_fd_sc_hd__buf_2
X_1852_ _2131_/C _1751_/A _1633_/X _1851_/Y vssd1 vssd1 vccd1 vccd1 _1852_/X sky130_fd_sc_hd__a211o_4
X_1783_ _1678_/A _1770_/Y _1783_/C _1777_/X vssd1 vssd1 vccd1 vccd1 _1783_/Y sky130_fd_sc_hd__nand4_4
X_2335_ _2335_/A _2335_/B _1218_/B _2335_/D vssd1 vssd1 vccd1 vccd1 _2335_/Y sky130_fd_sc_hd__nand4_4
XFILLER_29_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2266_ _2266_/A vssd1 vssd1 vccd1 vccd1 _2266_/Y sky130_fd_sc_hd__inv_2
X_2404_ _2404_/CLK _2404_/D vssd1 vssd1 vccd1 vccd1 _2306_/C sky130_fd_sc_hd__dfxtp_4
X_1217_ _1185_/A vssd1 vssd1 vccd1 vccd1 _1218_/B sky130_fd_sc_hd__buf_2
XFILLER_25_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2197_ _2306_/C _1618_/X vssd1 vssd1 vccd1 vccd1 _2198_/C sky130_fd_sc_hd__nand2_4
XFILLER_33_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2120_ _2120_/A vssd1 vssd1 vccd1 vccd1 _2120_/X sky130_fd_sc_hd__buf_2
X_2051_ _2014_/X _2040_/X _1346_/X vssd1 vssd1 vccd1 vccd1 _2051_/Y sky130_fd_sc_hd__o21ai_4
X_1835_ _1830_/B _1834_/Y _1831_/B vssd1 vssd1 vccd1 vccd1 _1835_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_30_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1904_ _2431_/Q vssd1 vssd1 vccd1 vccd1 _1904_/Y sky130_fd_sc_hd__inv_2
XFILLER_15_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1697_ _1697_/A vssd1 vssd1 vccd1 vccd1 _1697_/Y sky130_fd_sc_hd__inv_2
X_1766_ _1438_/C _1766_/B vssd1 vssd1 vccd1 vccd1 _1766_/Y sky130_fd_sc_hd__nor2_4
X_2249_ _2248_/X vssd1 vssd1 vccd1 vccd1 _2249_/X sky130_fd_sc_hd__buf_2
X_2318_ _2158_/B _2311_/X _2136_/A _2313_/X vssd1 vssd1 vccd1 vccd1 _2398_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_31_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1551_ _1546_/X _1550_/Y _1454_/X vssd1 vssd1 vccd1 vccd1 _1551_/Y sky130_fd_sc_hd__a21oi_4
X_1482_ _1467_/Y _1424_/Y _1428_/Y vssd1 vssd1 vccd1 vccd1 _1482_/Y sky130_fd_sc_hd__nor3_4
XFILLER_8_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1620_ _1618_/X _1619_/Y vssd1 vssd1 vccd1 vccd1 _1620_/Y sky130_fd_sc_hd__nor2_4
X_2103_ _2103_/A vssd1 vssd1 vccd1 vccd1 _2103_/Y sky130_fd_sc_hd__inv_2
XFILLER_39_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2034_ _1997_/A _2032_/X _2033_/Y vssd1 vssd1 vccd1 vccd1 _2487_/D sky130_fd_sc_hd__o21a_4
X_1818_ _2576_/Q _1810_/X _1813_/X vssd1 vssd1 vccd1 vccd1 _1818_/X sky130_fd_sc_hd__o21a_4
XFILLER_10_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1749_ _1745_/X _1748_/Y _1628_/X vssd1 vssd1 vccd1 vccd1 _1749_/X sky130_fd_sc_hd__a21o_4
XFILLER_26_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_4_4_0_addressalyzerBlock.SPI_CLK clkbuf_3_2_0_addressalyzerBlock.SPI_CLK/X
+ vssd1 vssd1 vccd1 vccd1 _2555_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_3_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2652_ _2646_/CLK _2356_/Y vssd1 vssd1 vccd1 vccd1 _2097_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_12_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1534_ _1534_/A vssd1 vssd1 vccd1 vccd1 _1534_/X sky130_fd_sc_hd__buf_2
X_1603_ _2117_/A vssd1 vssd1 vccd1 vccd1 _1603_/Y sky130_fd_sc_hd__inv_2
X_2583_ _2446_/CLK _1801_/X vssd1 vssd1 vccd1 vccd1 _2583_/Q sky130_fd_sc_hd__dfxtp_4
X_1465_ _1458_/Y _1463_/Y _1464_/Y vssd1 vssd1 vccd1 vccd1 _2611_/D sky130_fd_sc_hd__a21oi_4
X_2017_ _2047_/A _2016_/X _1997_/A _1997_/D vssd1 vssd1 vccd1 vccd1 _2017_/X sky130_fd_sc_hd__and4_4
X_1396_ _1231_/B vssd1 vssd1 vccd1 vccd1 _1397_/A sky130_fd_sc_hd__inv_2
XFILLER_2_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1181_ _1198_/B vssd1 vssd1 vccd1 vccd1 _1194_/B sky130_fd_sc_hd__buf_2
X_1250_ _1267_/A _1277_/B _1256_/A _1249_/Y vssd1 vssd1 vccd1 vccd1 _1252_/A sky130_fd_sc_hd__nand4_4
XFILLER_32_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_4_8_0_m1_clk_local clkbuf_4_9_0_m1_clk_local/A vssd1 vssd1 vccd1 vccd1 _2476_/CLK
+ sky130_fd_sc_hd__clkbuf_1
X_2635_ _2635_/CLK _1314_/Y vssd1 vssd1 vccd1 vccd1 _2635_/Q sky130_fd_sc_hd__dfxtp_4
X_2497_ _2508_/CLK _2497_/D vssd1 vssd1 vccd1 vccd1 _2497_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_55_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1448_ _1448_/A vssd1 vssd1 vccd1 vccd1 _1449_/B sky130_fd_sc_hd__buf_2
X_2566_ _2551_/CLK _2566_/D vssd1 vssd1 vccd1 vccd1 _2566_/Q sky130_fd_sc_hd__dfxtp_4
X_1517_ _1513_/X _1515_/Y _1516_/X vssd1 vssd1 vccd1 vccd1 _2606_/D sky130_fd_sc_hd__a21oi_4
XFILLER_55_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1379_ _1385_/B vssd1 vssd1 vccd1 vccd1 _1395_/B sky130_fd_sc_hd__buf_2
XFILLER_23_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2420_ _2555_/CLK _2274_/Y vssd1 vssd1 vccd1 vccd1 _1946_/A sky130_fd_sc_hd__dfxtp_4
X_2351_ _2545_/Q _2546_/Q _2351_/C vssd1 vssd1 vccd1 vccd1 _2352_/C sky130_fd_sc_hd__or3_4
X_1233_ _1229_/Y _1363_/A _1231_/Y _1363_/C vssd1 vssd1 vccd1 vccd1 _1385_/B sky130_fd_sc_hd__nor4_4
X_1302_ _1302_/A vssd1 vssd1 vccd1 vccd1 _2637_/D sky130_fd_sc_hd__inv_2
XFILLER_29_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2282_ _2276_/X _2127_/Y _2278_/X _1706_/B _2280_/X vssd1 vssd1 vccd1 vccd1 _2282_/Y
+ sky130_fd_sc_hd__o32ai_4
XFILLER_64_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1997_ _1997_/A _1997_/B _2488_/Q _1997_/D vssd1 vssd1 vccd1 vccd1 _2008_/A sky130_fd_sc_hd__nand4_4
XFILLER_20_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2549_ _2464_/CLK _1893_/X vssd1 vssd1 vccd1 vccd1 _2549_/Q sky130_fd_sc_hd__dfxtp_4
X_2618_ _2619_/CLK _2618_/D vssd1 vssd1 vccd1 vccd1 _1231_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_47_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_0_0_addressalyzerBlock.SPI_CLK clkbuf_0_addressalyzerBlock.SPI_CLK/X vssd1
+ vssd1 vccd1 vccd1 clkbuf_2_1_0_addressalyzerBlock.SPI_CLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_19_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1851_ _1635_/X _1766_/B vssd1 vssd1 vccd1 vccd1 _1851_/Y sky130_fd_sc_hd__nor2_4
X_1920_ _1918_/A _2538_/Q vssd1 vssd1 vccd1 vccd1 _1920_/X sky130_fd_sc_hd__and2_4
X_1782_ _1779_/Y _1780_/Y _2100_/A vssd1 vssd1 vccd1 vccd1 _2589_/D sky130_fd_sc_hd__a21oi_4
X_2403_ _2551_/CLK _2403_/D vssd1 vssd1 vccd1 vccd1 _2089_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_6_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1216_ _1194_/B _1188_/X _2645_/Q vssd1 vssd1 vccd1 vccd1 _1216_/Y sky130_fd_sc_hd__nand3_4
X_2334_ _1530_/C _2333_/Y _2100_/A vssd1 vssd1 vccd1 vccd1 _2389_/D sky130_fd_sc_hd__a21oi_4
X_2265_ _1420_/Y _2262_/X _2258_/X _1622_/Y _2264_/X vssd1 vssd1 vccd1 vccd1 _2426_/D
+ sky130_fd_sc_hd__o32ai_4
X_2196_ _2196_/A _2196_/B vssd1 vssd1 vccd1 vccd1 _2196_/Y sky130_fd_sc_hd__nand2_4
XFILLER_52_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2050_ _2049_/Y vssd1 vssd1 vccd1 vccd1 _2050_/Y sky130_fd_sc_hd__inv_2
XFILLER_62_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1834_ _1833_/Y vssd1 vssd1 vccd1 vccd1 _1834_/Y sky130_fd_sc_hd__inv_2
XFILLER_30_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1765_ _1765_/A vssd1 vssd1 vccd1 vccd1 _1766_/B sky130_fd_sc_hd__inv_2
X_1903_ _1911_/A _1902_/Y vssd1 vssd1 vccd1 vccd1 _2542_/D sky130_fd_sc_hd__nor2_4
X_1696_ _1696_/A vssd1 vssd1 vccd1 vccd1 _1698_/A sky130_fd_sc_hd__buf_2
XFILLER_25_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2248_ _1583_/X _1594_/X _1597_/X _1696_/A _1736_/A vssd1 vssd1 vccd1 vccd1 _2248_/X
+ sky130_fd_sc_hd__a41o_4
X_2317_ _1750_/Y _2311_/X _1490_/A _2313_/X vssd1 vssd1 vccd1 vccd1 _2399_/D sky130_fd_sc_hd__a2bb2o_4
X_2179_ _2177_/Y _2201_/B _2179_/C vssd1 vssd1 vccd1 vccd1 _2179_/Y sky130_fd_sc_hd__nand3_4
XFILLER_25_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1550_ _1547_/X _1548_/Y _1549_/Y vssd1 vssd1 vccd1 vccd1 _1550_/Y sky130_fd_sc_hd__o21ai_4
X_1481_ _1436_/B vssd1 vssd1 vccd1 vccd1 _1487_/A sky130_fd_sc_hd__buf_2
X_2033_ _2032_/C _2047_/A _1997_/A _1997_/D _1275_/X vssd1 vssd1 vccd1 vccd1 _2033_/Y
+ sky130_fd_sc_hd__a41oi_4
X_2102_ _2102_/A _2103_/A _2104_/D _2091_/Y vssd1 vssd1 vccd1 vccd1 _2461_/D sky130_fd_sc_hd__nor4_4
XFILLER_62_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1817_ _2576_/Q _1809_/X _1816_/X vssd1 vssd1 vccd1 vccd1 _2577_/D sky130_fd_sc_hd__o21a_4
X_1748_ _1746_/Y _1624_/X _1747_/Y vssd1 vssd1 vccd1 vccd1 _1748_/Y sky130_fd_sc_hd__o21ai_4
X_1679_ _1566_/X _1683_/A vssd1 vssd1 vccd1 vccd1 _1679_/Y sky130_fd_sc_hd__nor2_4
XFILLER_53_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2651_ _2454_/CLK _1193_/Y vssd1 vssd1 vccd1 vccd1 _2353_/A sky130_fd_sc_hd__dfxtp_4
X_1602_ _1602_/A _1602_/B _1602_/C vssd1 vssd1 vccd1 vccd1 _2117_/A sky130_fd_sc_hd__nand3_4
X_2582_ _2399_/CLK _1803_/X vssd1 vssd1 vccd1 vccd1 _1503_/A sky130_fd_sc_hd__dfxtp_4
X_1395_ _2019_/A _1395_/B _1394_/Y vssd1 vssd1 vccd1 vccd1 _1395_/Y sky130_fd_sc_hd__nor3_4
X_1464_ _1438_/B _1449_/B _1213_/X vssd1 vssd1 vccd1 vccd1 _1464_/Y sky130_fd_sc_hd__o21ai_4
X_1533_ _2604_/Q vssd1 vssd1 vccd1 vccd1 _1534_/A sky130_fd_sc_hd__inv_2
X_2016_ _1987_/A vssd1 vssd1 vccd1 vccd1 _2016_/X sky130_fd_sc_hd__buf_2
XFILLER_35_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1180_ _1833_/A vssd1 vssd1 vccd1 vccd1 _1198_/B sky130_fd_sc_hd__inv_2
XFILLER_32_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2634_ _2476_/CLK _1320_/Y vssd1 vssd1 vccd1 vccd1 _1856_/B sky130_fd_sc_hd__dfxtp_4
X_2565_ _2561_/CLK _2565_/D vssd1 vssd1 vccd1 vccd1 _1883_/B sky130_fd_sc_hd__dfxtp_4
X_1516_ _1450_/X _1512_/Y _1500_/X vssd1 vssd1 vccd1 vccd1 _1516_/X sky130_fd_sc_hd__a21o_4
X_2496_ _2508_/CLK _2496_/D vssd1 vssd1 vccd1 vccd1 _1972_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_55_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1378_ _1378_/A vssd1 vssd1 vccd1 vccd1 _1378_/Y sky130_fd_sc_hd__inv_2
XFILLER_4_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1447_ _1446_/Y vssd1 vssd1 vccd1 vccd1 _1448_/A sky130_fd_sc_hd__inv_2
XFILLER_23_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2350_ _2349_/A _2348_/Y _2349_/Y vssd1 vssd1 vccd1 vccd1 MISO_toHost sky130_fd_sc_hd__a21oi_4
X_1232_ _1232_/A _2615_/Q _2614_/Q _1406_/A vssd1 vssd1 vccd1 vccd1 _1363_/C sky130_fd_sc_hd__nand4_4
X_1301_ _1301_/A _2022_/B _1301_/C vssd1 vssd1 vccd1 vccd1 _1302_/A sky130_fd_sc_hd__nand3_4
X_2281_ _2276_/X _2122_/Y _2278_/X _1619_/Y _2280_/X vssd1 vssd1 vccd1 vccd1 _2281_/Y
+ sky130_fd_sc_hd__o32ai_4
X_1996_ _1995_/Y vssd1 vssd1 vccd1 vccd1 _1997_/D sky130_fd_sc_hd__inv_2
XFILLER_9_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2548_ _2464_/CLK _2548_/D vssd1 vssd1 vccd1 vccd1 _2548_/Q sky130_fd_sc_hd__dfxtp_4
X_2617_ _2619_/CLK _1404_/Y vssd1 vssd1 vccd1 vccd1 _1231_/B sky130_fd_sc_hd__dfxtp_4
X_2479_ _2511_/CLK _2065_/X vssd1 vssd1 vccd1 vccd1 _2479_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_28_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1781_ _1781_/A vssd1 vssd1 vccd1 vccd1 _2100_/A sky130_fd_sc_hd__buf_2
X_1850_ _1846_/X _1849_/Y _1628_/X vssd1 vssd1 vccd1 vccd1 _1850_/X sky130_fd_sc_hd__a21o_4
XFILLER_41_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2333_ _1218_/B _2333_/B vssd1 vssd1 vccd1 vccd1 _2333_/Y sky130_fd_sc_hd__nand2_4
XFILLER_6_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2402_ _2604_/CLK _2402_/D vssd1 vssd1 vccd1 vccd1 _2402_/Q sky130_fd_sc_hd__dfxtp_4
X_1215_ _1211_/Y _2322_/A _1214_/Y vssd1 vssd1 vccd1 vccd1 _1215_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_37_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2195_ _1534_/A _2552_/Q _2148_/X vssd1 vssd1 vccd1 vccd1 _2195_/Y sky130_fd_sc_hd__o21ai_4
X_2264_ _2263_/X vssd1 vssd1 vccd1 vccd1 _2264_/X sky130_fd_sc_hd__buf_2
XFILLER_52_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1979_ _1972_/A _1972_/B vssd1 vssd1 vccd1 vccd1 _1980_/C sky130_fd_sc_hd__or2_4
XFILLER_4_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1902_ _1902_/A vssd1 vssd1 vccd1 vccd1 _1902_/Y sky130_fd_sc_hd__inv_2
X_1833_ _1833_/A _1830_/C vssd1 vssd1 vccd1 vccd1 _1833_/Y sky130_fd_sc_hd__nand2_4
X_1764_ _1764_/A vssd1 vssd1 vccd1 vccd1 _1764_/Y sky130_fd_sc_hd__inv_2
X_1695_ _1694_/X vssd1 vssd1 vccd1 vccd1 _1696_/A sky130_fd_sc_hd__buf_2
X_2316_ _1766_/B _2311_/X _1477_/X _2313_/X vssd1 vssd1 vccd1 vccd1 _2400_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_57_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2247_ _2246_/Y vssd1 vssd1 vccd1 vccd1 _2247_/X sky130_fd_sc_hd__buf_2
X_2178_ _2421_/Q _1634_/X vssd1 vssd1 vccd1 vccd1 _2179_/C sky130_fd_sc_hd__nand2_4
XFILLER_40_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_9_0_addressalyzerBlock.SPI_CLK clkbuf_4_9_0_addressalyzerBlock.SPI_CLK/A
+ vssd1 vssd1 vccd1 vccd1 _2389_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1480_ _1476_/Y _1478_/Y _1479_/Y vssd1 vssd1 vccd1 vccd1 _2610_/D sky130_fd_sc_hd__a21oi_4
X_2032_ _2029_/Y _2030_/X _2032_/C _1997_/D vssd1 vssd1 vccd1 vccd1 _2032_/X sky130_fd_sc_hd__and4_4
X_2101_ _2101_/A vssd1 vssd1 vccd1 vccd1 _2102_/A sky130_fd_sc_hd__buf_2
XFILLER_50_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1678_ _1678_/A vssd1 vssd1 vccd1 vccd1 _1678_/Y sky130_fd_sc_hd__inv_2
X_1816_ _2577_/Q _1810_/X _1813_/X vssd1 vssd1 vccd1 vccd1 _1816_/X sky130_fd_sc_hd__o21a_4
X_1747_ _1625_/X _2431_/Q _1708_/X vssd1 vssd1 vccd1 vccd1 _1747_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_53_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2650_ _2454_/CLK _1197_/Y vssd1 vssd1 vccd1 vccd1 _2650_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_8_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2581_ _2399_/CLK _1805_/X vssd1 vssd1 vccd1 vccd1 _1514_/A sky130_fd_sc_hd__dfxtp_4
X_1601_ _1555_/A vssd1 vssd1 vccd1 vccd1 _1602_/C sky130_fd_sc_hd__buf_2
X_1532_ _1420_/A _1527_/Y _1556_/A vssd1 vssd1 vccd1 vccd1 _1532_/Y sky130_fd_sc_hd__a21oi_4
X_1394_ _2619_/Q _1394_/B vssd1 vssd1 vccd1 vccd1 _1394_/Y sky130_fd_sc_hd__nor2_4
X_1463_ _2266_/A _2333_/B _1462_/X vssd1 vssd1 vccd1 vccd1 _1463_/Y sky130_fd_sc_hd__a21oi_4
X_2015_ _2014_/X _1986_/Y _2015_/C vssd1 vssd1 vccd1 vccd1 _2047_/A sky130_fd_sc_hd__nor3_4
XFILLER_50_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_2_1_0_m1_clk_local clkbuf_1_0_0_m1_clk_local/X vssd1 vssd1 vccd1 vccd1 clkbuf_3_3_0_m1_clk_local/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_53_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_2_0_0_addressalyzerBlock.SPI_CLK clkbuf_2_1_0_addressalyzerBlock.SPI_CLK/A
+ vssd1 vssd1 vccd1 vccd1 clkbuf_3_1_0_addressalyzerBlock.SPI_CLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_20_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2495_ _2508_/CLK _2495_/D vssd1 vssd1 vccd1 vccd1 _1972_/A sky130_fd_sc_hd__dfxtp_4
X_2633_ _2476_/CLK _2633_/D vssd1 vssd1 vccd1 vccd1 _1315_/A sky130_fd_sc_hd__dfxtp_4
X_2564_ _2555_/CLK _2564_/D vssd1 vssd1 vccd1 vccd1 _1884_/B sky130_fd_sc_hd__dfxtp_4
X_1515_ _1514_/X _1460_/X _1462_/X vssd1 vssd1 vccd1 vccd1 _1515_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_55_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1377_ _1375_/X _1376_/Y vssd1 vssd1 vccd1 vccd1 _1378_/A sky130_fd_sc_hd__nand2_4
X_1446_ _1530_/A _1445_/A _1445_/Y vssd1 vssd1 vccd1 vccd1 _1446_/Y sky130_fd_sc_hd__nand3_4
XFILLER_4_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1231_ _1231_/A _1231_/B vssd1 vssd1 vccd1 vccd1 _1231_/Y sky130_fd_sc_hd__nand2_4
XFILLER_37_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1300_ _1300_/A _1299_/Y vssd1 vssd1 vccd1 vccd1 _1301_/C sky130_fd_sc_hd__nand2_4
X_2280_ _2279_/X vssd1 vssd1 vccd1 vccd1 _2280_/X sky130_fd_sc_hd__buf_2
X_1995_ _2043_/D _1995_/B vssd1 vssd1 vccd1 vccd1 _1995_/Y sky130_fd_sc_hd__nand2_4
X_2616_ _2619_/CLK _2616_/D vssd1 vssd1 vccd1 vccd1 _1230_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_20_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2547_ _2464_/CLK _2547_/D vssd1 vssd1 vccd1 vccd1 _2547_/Q sky130_fd_sc_hd__dfxtp_4
X_2478_ _2511_/CLK _2067_/Y vssd1 vssd1 vccd1 vccd1 _2054_/A sky130_fd_sc_hd__dfxtp_4
X_1429_ _1424_/Y _1428_/Y vssd1 vssd1 vccd1 vccd1 _1432_/A sky130_fd_sc_hd__nor2_4
XFILLER_43_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_4_4_0_m1_clk_local clkbuf_3_2_0_m1_clk_local/X vssd1 vssd1 vccd1 vccd1 _2527_/CLK
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_18_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1780_ _1678_/Y _2589_/Q vssd1 vssd1 vccd1 vccd1 _1780_/Y sky130_fd_sc_hd__nand2_4
XFILLER_6_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2332_ _1218_/B _2322_/B _2102_/A _1729_/Y vssd1 vssd1 vccd1 vccd1 _2332_/X sky130_fd_sc_hd__a211o_4
X_2401_ _2399_/CLK _2315_/X vssd1 vssd1 vccd1 vccd1 _2401_/Q sky130_fd_sc_hd__dfxtp_4
X_1214_ _2436_/Q _1187_/A _1213_/X vssd1 vssd1 vccd1 vccd1 _1214_/Y sky130_fd_sc_hd__o21ai_4
X_2194_ _2614_/Q _1571_/A _1568_/A _1660_/A _2146_/Y vssd1 vssd1 vccd1 vccd1 _2194_/Y
+ sky130_fd_sc_hd__o41ai_4
XFILLER_25_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2263_ _1583_/X _1594_/X _1669_/B _1694_/X _1736_/A vssd1 vssd1 vccd1 vccd1 _2263_/X
+ sky130_fd_sc_hd__a41o_4
XFILLER_52_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1978_ _1978_/A _1972_/Y _1977_/X vssd1 vssd1 vccd1 vccd1 _2497_/D sky130_fd_sc_hd__and3_4
XFILLER_29_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1832_ _1829_/Y _1830_/Y _1831_/Y vssd1 vssd1 vccd1 vccd1 _1832_/Y sky130_fd_sc_hd__a21oi_4
X_1901_ _2063_/A vssd1 vssd1 vccd1 vccd1 _1911_/A sky130_fd_sc_hd__buf_2
X_1763_ _1740_/Y _1760_/Y _1762_/Y vssd1 vssd1 vccd1 vccd1 _1763_/Y sky130_fd_sc_hd__o21ai_4
X_1694_ _2594_/Q vssd1 vssd1 vccd1 vccd1 _1694_/X sky130_fd_sc_hd__buf_2
X_2246_ _2245_/Y vssd1 vssd1 vccd1 vccd1 _2246_/Y sky130_fd_sc_hd__inv_2
X_2315_ _1713_/Y _2311_/X _2266_/A _2313_/X vssd1 vssd1 vccd1 vccd1 _2315_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_15_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2177_ _2196_/A _2177_/B vssd1 vssd1 vccd1 vccd1 _2177_/Y sky130_fd_sc_hd__nand2_4
Xclkbuf_4_14_0_addressalyzerBlock.SPI_CLK clkbuf_3_7_0_addressalyzerBlock.SPI_CLK/X
+ vssd1 vssd1 vccd1 vccd1 _2646_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_31_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2100_ _2100_/A _2099_/C _2098_/Y vssd1 vssd1 vccd1 vccd1 _2462_/D sky130_fd_sc_hd__nor3_4
XFILLER_39_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2031_ _2016_/X vssd1 vssd1 vccd1 vccd1 _2032_/C sky130_fd_sc_hd__buf_2
XFILLER_54_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1815_ _2577_/Q _1809_/X _1814_/X vssd1 vssd1 vccd1 vccd1 _1815_/X sky130_fd_sc_hd__o21a_4
X_1677_ _1674_/Y _1677_/B vssd1 vssd1 vccd1 vccd1 _2596_/D sky130_fd_sc_hd__nand2_4
X_1746_ _2423_/Q vssd1 vssd1 vccd1 vccd1 _1746_/Y sky130_fd_sc_hd__inv_2
X_2229_ _1645_/A _1333_/A _1612_/A vssd1 vssd1 vccd1 vccd1 _2229_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_26_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1531_ _1564_/A vssd1 vssd1 vccd1 vccd1 _1556_/A sky130_fd_sc_hd__buf_2
X_1600_ _1541_/X _1597_/X vssd1 vssd1 vccd1 vccd1 _1602_/B sky130_fd_sc_hd__nand2_4
X_2580_ _2611_/CLK _1807_/X vssd1 vssd1 vccd1 vccd1 _2580_/Q sky130_fd_sc_hd__dfxtp_4
X_1462_ _1450_/X vssd1 vssd1 vccd1 vccd1 _1462_/X sky130_fd_sc_hd__buf_2
X_1393_ _1385_/D _1395_/B _1392_/Y vssd1 vssd1 vccd1 vccd1 _2620_/D sky130_fd_sc_hd__o21a_4
X_2014_ _1985_/Y vssd1 vssd1 vccd1 vccd1 _2014_/X sky130_fd_sc_hd__buf_2
XFILLER_35_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1729_ _2386_/Q _1729_/B _1689_/Y vssd1 vssd1 vccd1 vccd1 _1729_/Y sky130_fd_sc_hd__nor3_4
XFILLER_37_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2632_ _2632_/CLK _1337_/Y vssd1 vssd1 vccd1 vccd1 _2632_/Q sky130_fd_sc_hd__dfxtp_4
X_1445_ _1445_/A _1434_/Y _1444_/Y _1445_/D vssd1 vssd1 vccd1 vccd1 _1445_/Y sky130_fd_sc_hd__nand4_4
X_2563_ _2551_/CLK _2563_/D vssd1 vssd1 vccd1 vccd1 _2563_/Q sky130_fd_sc_hd__dfxtp_4
X_2494_ _2588_/CLK _2494_/D vssd1 vssd1 vccd1 vccd1 _1184_/A sky130_fd_sc_hd__dfxtp_4
X_1514_ _1514_/A vssd1 vssd1 vccd1 vccd1 _1514_/X sky130_fd_sc_hd__buf_2
X_1376_ _1366_/X _1376_/B _1376_/C vssd1 vssd1 vccd1 vccd1 _1376_/Y sky130_fd_sc_hd__nand3_4
Xclkbuf_4_12_0_m1_clk_local clkbuf_3_6_0_m1_clk_local/X vssd1 vssd1 vccd1 vccd1 _2619_/CLK
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_23_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1230_ _1230_/A vssd1 vssd1 vccd1 vccd1 _1363_/A sky130_fd_sc_hd__inv_2
XFILLER_49_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1994_ _1985_/Y _1986_/Y _1994_/C _2015_/C vssd1 vssd1 vccd1 vccd1 _1997_/B sky130_fd_sc_hd__nor4_4
XFILLER_20_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2615_ _2619_/CLK _1412_/X vssd1 vssd1 vccd1 vccd1 _2615_/Q sky130_fd_sc_hd__dfxtp_4
X_2546_ _2464_/CLK _1896_/X vssd1 vssd1 vccd1 vccd1 _2546_/Q sky130_fd_sc_hd__dfxtp_4
X_2477_ _2476_/CLK _2070_/Y vssd1 vssd1 vccd1 vccd1 _2477_/Q sky130_fd_sc_hd__dfxtp_4
X_1428_ _1570_/A _1567_/A _1567_/B _1567_/C vssd1 vssd1 vccd1 vccd1 _1428_/Y sky130_fd_sc_hd__nand4_4
XFILLER_28_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1359_ _1359_/A vssd1 vssd1 vccd1 vccd1 _1359_/Y sky130_fd_sc_hd__inv_2
XPHY_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2400_ _2399_/CLK _2400_/D vssd1 vssd1 vccd1 vccd1 _1765_/A sky130_fd_sc_hd__dfxtp_4
X_1213_ _2096_/A vssd1 vssd1 vccd1 vccd1 _1213_/X sky130_fd_sc_hd__buf_2
X_2331_ _2092_/A _2331_/B vssd1 vssd1 vccd1 vccd1 _2331_/Y sky130_fd_sc_hd__nor2_4
X_2262_ _1648_/Y vssd1 vssd1 vccd1 vccd1 _2262_/X sky130_fd_sc_hd__buf_2
XFILLER_65_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2193_ _1676_/A _2191_/Y _2192_/Y vssd1 vssd1 vccd1 vccd1 _2193_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_37_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1977_ _1972_/A _1972_/B _2497_/Q vssd1 vssd1 vccd1 vccd1 _1977_/X sky130_fd_sc_hd__a21o_4
XFILLER_33_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2529_ _2527_/CLK _2529_/D vssd1 vssd1 vccd1 vccd1 _2529_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_20_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1900_ _2093_/A _2547_/Q vssd1 vssd1 vccd1 vccd1 _2543_/D sky130_fd_sc_hd__and2_4
X_1831_ _1831_/A _1831_/B vssd1 vssd1 vccd1 vccd1 _1831_/Y sky130_fd_sc_hd__nand2_4
XFILLER_30_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1762_ _2192_/A _1762_/B vssd1 vssd1 vccd1 vccd1 _1762_/Y sky130_fd_sc_hd__nand2_4
X_1693_ _1688_/Y _1690_/Y _1692_/X vssd1 vssd1 vccd1 vccd1 _1693_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_65_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2245_ _1219_/X _1581_/A _2289_/C vssd1 vssd1 vccd1 vccd1 _2245_/Y sky130_fd_sc_hd__nor3_4
X_2314_ _1636_/Y _2311_/X _1420_/A _2313_/X vssd1 vssd1 vccd1 vccd1 _2402_/D sky130_fd_sc_hd__a2bb2o_4
X_2176_ _2174_/Y _1708_/X _2176_/C vssd1 vssd1 vccd1 vccd1 _2176_/Y sky130_fd_sc_hd__nand3_4
XFILLER_15_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2030_ _2483_/Q vssd1 vssd1 vccd1 vccd1 _2030_/X sky130_fd_sc_hd__buf_2
XFILLER_47_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1814_ _2578_/Q _1810_/X _1813_/X vssd1 vssd1 vccd1 vccd1 _1814_/X sky130_fd_sc_hd__o21a_4
XFILLER_7_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1745_ _2407_/Q _2224_/A _2201_/B _1744_/Y vssd1 vssd1 vccd1 vccd1 _1745_/X sky130_fd_sc_hd__a211o_4
XFILLER_15_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1676_ _1676_/A _1676_/B vssd1 vssd1 vccd1 vccd1 _1677_/B sky130_fd_sc_hd__nand2_4
X_2228_ _2217_/Y _2226_/Y _2227_/Y vssd1 vssd1 vccd1 vccd1 _2228_/Y sky130_fd_sc_hd__o21ai_4
X_2159_ _2442_/Q _1635_/X _1632_/Y _2158_/Y vssd1 vssd1 vccd1 vccd1 _2159_/X sky130_fd_sc_hd__a211o_4
Xclkbuf_3_0_0_addressalyzerBlock.SPI_CLK clkbuf_3_1_0_addressalyzerBlock.SPI_CLK/A
+ vssd1 vssd1 vccd1 vccd1 clkbuf_3_0_0_addressalyzerBlock.SPI_CLK/X sky130_fd_sc_hd__clkbuf_1
XFILLER_13_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1392_ _1395_/B _1385_/D _2063_/A vssd1 vssd1 vccd1 vccd1 _1392_/Y sky130_fd_sc_hd__a21oi_4
X_1530_ _1530_/A _1445_/Y _1530_/C vssd1 vssd1 vccd1 vccd1 _1564_/A sky130_fd_sc_hd__nand3_4
X_1461_ _1460_/X vssd1 vssd1 vccd1 vccd1 _2333_/B sky130_fd_sc_hd__buf_2
X_2013_ _2002_/X _2003_/Y _2013_/C _2013_/D vssd1 vssd1 vccd1 vccd1 _2019_/B sky130_fd_sc_hd__nor4_4
XFILLER_50_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1728_ _1697_/A _2391_/Q _1687_/A vssd1 vssd1 vccd1 vccd1 _1728_/Y sky130_fd_sc_hd__nor3_4
X_1659_ _1659_/A vssd1 vssd1 vccd1 vccd1 _1660_/A sky130_fd_sc_hd__buf_2
XFILLER_26_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2562_ _2561_/CLK _1877_/X vssd1 vssd1 vccd1 vccd1 _2562_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_57_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2631_ _2632_/CLK _2631_/D vssd1 vssd1 vccd1 vccd1 _2631_/Q sky130_fd_sc_hd__dfxtp_4
X_2493_ _2470_/CLK _2493_/D vssd1 vssd1 vccd1 vccd1 CLK_LED sky130_fd_sc_hd__dfxtp_4
X_1375_ _1376_/B _1373_/X _1374_/X vssd1 vssd1 vccd1 vccd1 _1375_/X sky130_fd_sc_hd__o21a_4
X_1444_ _2385_/Q vssd1 vssd1 vccd1 vccd1 _1444_/Y sky130_fd_sc_hd__inv_2
XFILLER_4_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1513_ _1511_/Y _1512_/Y _1508_/X vssd1 vssd1 vccd1 vccd1 _1513_/X sky130_fd_sc_hd__a21o_4
XFILLER_48_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1993_ _2479_/Q _1993_/B _1993_/C _2481_/Q vssd1 vssd1 vccd1 vccd1 _2015_/C sky130_fd_sc_hd__nand4_4
XFILLER_45_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2545_ _2464_/CLK _2545_/D vssd1 vssd1 vccd1 vccd1 _2545_/Q sky130_fd_sc_hd__dfxtp_4
X_2614_ _2623_/CLK _1417_/Y vssd1 vssd1 vccd1 vccd1 _2614_/Q sky130_fd_sc_hd__dfxtp_4
X_2476_ _2476_/CLK _2476_/D vssd1 vssd1 vccd1 vccd1 _2476_/Q sky130_fd_sc_hd__dfxtp_4
X_1358_ _1358_/A _2022_/B _1358_/C vssd1 vssd1 vccd1 vccd1 _1359_/A sky130_fd_sc_hd__nand3_4
X_1427_ _2597_/Q vssd1 vssd1 vccd1 vccd1 _1567_/C sky130_fd_sc_hd__buf_2
XFILLER_18_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1289_ _1289_/A _1289_/B _1289_/C vssd1 vssd1 vccd1 vccd1 _1290_/A sky130_fd_sc_hd__nand3_4
XFILLER_3_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2192_ _2192_/A _2192_/B vssd1 vssd1 vccd1 vccd1 _2192_/Y sky130_fd_sc_hd__nand2_4
X_1212_ _1188_/A vssd1 vssd1 vccd1 vccd1 _2322_/A sky130_fd_sc_hd__buf_2
X_2330_ _1839_/A _2385_/Q _2322_/A _2333_/B vssd1 vssd1 vccd1 vccd1 _2331_/B sky130_fd_sc_hd__a22oi_4
X_2261_ _2243_/Y _2260_/Y _2258_/X _1913_/Y _2248_/X vssd1 vssd1 vccd1 vccd1 _2427_/D
+ sky130_fd_sc_hd__o32ai_4
XFILLER_52_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1976_ _1869_/A _1867_/Y vssd1 vssd1 vccd1 vccd1 _1978_/A sky130_fd_sc_hd__nor2_4
XFILLER_29_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2528_ _2527_/CLK _2528_/D vssd1 vssd1 vccd1 vccd1 _2528_/Q sky130_fd_sc_hd__dfxtp_4
X_2459_ _2646_/CLK _2105_/X vssd1 vssd1 vccd1 vccd1 _2103_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_29_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_4_0_0_m1_clk_local clkbuf_3_0_0_m1_clk_local/X vssd1 vssd1 vccd1 vccd1 _2538_/CLK
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_15_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1830_ _1179_/X _1830_/B _1830_/C vssd1 vssd1 vccd1 vccd1 _1830_/Y sky130_fd_sc_hd__nand3_4
XFILLER_51_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1761_ _1761_/A vssd1 vssd1 vccd1 vccd1 _2192_/A sky130_fd_sc_hd__buf_2
XFILLER_42_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1692_ _2289_/C _1488_/X _2589_/Q _1731_/B vssd1 vssd1 vccd1 vccd1 _1692_/X sky130_fd_sc_hd__a2bb2o_4
X_2313_ _2312_/X vssd1 vssd1 vccd1 vccd1 _2313_/X sky130_fd_sc_hd__buf_2
XFILLER_53_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2244_ _2243_/Y vssd1 vssd1 vccd1 vccd1 _2244_/X sky130_fd_sc_hd__buf_2
X_2175_ _1232_/A _1618_/X vssd1 vssd1 vccd1 vccd1 _2176_/C sky130_fd_sc_hd__nand2_4
XFILLER_40_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1959_ _1969_/A _2515_/Q vssd1 vssd1 vccd1 vccd1 _2507_/D sky130_fd_sc_hd__and2_4
XFILLER_48_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_3_6_0_m1_clk_local clkbuf_3_7_0_m1_clk_local/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_6_0_m1_clk_local/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_21_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1813_ _1789_/X vssd1 vssd1 vccd1 vccd1 _1813_/X sky130_fd_sc_hd__buf_2
XFILLER_7_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1744_ _1630_/X _1744_/B vssd1 vssd1 vccd1 vccd1 _1744_/Y sky130_fd_sc_hd__nor2_4
X_1675_ _1761_/A vssd1 vssd1 vccd1 vccd1 _1676_/A sky130_fd_sc_hd__buf_2
X_2227_ _1299_/Y _1854_/B _1856_/C _1856_/A vssd1 vssd1 vccd1 vccd1 _2227_/Y sky130_fd_sc_hd__a2bb2oi_4
X_2089_ _2089_/A vssd1 vssd1 vccd1 vccd1 _2089_/Y sky130_fd_sc_hd__inv_2
XFILLER_26_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2158_ _2224_/A _2158_/B vssd1 vssd1 vccd1 vccd1 _2158_/Y sky130_fd_sc_hd__nor2_4
XFILLER_32_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1391_ _1274_/X vssd1 vssd1 vccd1 vccd1 _2063_/A sky130_fd_sc_hd__buf_2
X_1460_ _2390_/Q vssd1 vssd1 vccd1 vccd1 _1460_/X sky130_fd_sc_hd__buf_2
X_2012_ _2008_/A vssd1 vssd1 vccd1 vccd1 _2013_/D sky130_fd_sc_hd__buf_2
XFILLER_35_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1727_ _1725_/X _1727_/B vssd1 vssd1 vccd1 vccd1 _1727_/Y sky130_fd_sc_hd__nand2_4
X_1658_ _1612_/X _1653_/Y _1657_/Y vssd1 vssd1 vccd1 vccd1 _1658_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_58_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1589_ _1589_/A vssd1 vssd1 vccd1 vccd1 _1589_/Y sky130_fd_sc_hd__inv_2
XFILLER_41_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2492_ _2492_/CLK _2492_/D vssd1 vssd1 vccd1 vccd1 _2492_/Q sky130_fd_sc_hd__dfxtp_4
X_2561_ _2561_/CLK _2561_/D vssd1 vssd1 vccd1 vccd1 _2561_/Q sky130_fd_sc_hd__dfxtp_4
X_2630_ _2632_/CLK _1343_/X vssd1 vssd1 vccd1 vccd1 _2630_/Q sky130_fd_sc_hd__dfxtp_4
X_1512_ _1486_/A vssd1 vssd1 vccd1 vccd1 _1512_/Y sky130_fd_sc_hd__inv_2
X_1374_ _1269_/A vssd1 vssd1 vccd1 vccd1 _1374_/X sky130_fd_sc_hd__buf_2
X_1443_ _1577_/A vssd1 vssd1 vccd1 vccd1 _1445_/A sky130_fd_sc_hd__inv_2
XFILLER_55_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1992_ _1992_/A _1992_/B _1990_/Y _2059_/A vssd1 vssd1 vccd1 vccd1 _1993_/B sky130_fd_sc_hd__nor4_4
X_2544_ _2464_/CLK _2544_/D vssd1 vssd1 vccd1 vccd1 _2544_/Q sky130_fd_sc_hd__dfxtp_4
X_2475_ _2476_/CLK _2077_/Y vssd1 vssd1 vccd1 vccd1 _2071_/A sky130_fd_sc_hd__dfxtp_4
X_2613_ _2619_/CLK _1419_/X vssd1 vssd1 vccd1 vccd1 _1406_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_55_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1357_ _1351_/B _1361_/B _1351_/A vssd1 vssd1 vccd1 vccd1 _1358_/C sky130_fd_sc_hd__o21ai_4
X_1426_ _1589_/A vssd1 vssd1 vccd1 vccd1 _1567_/B sky130_fd_sc_hd__buf_2
X_1288_ _1265_/A _1300_/A _1225_/X vssd1 vssd1 vccd1 vccd1 _1289_/C sky130_fd_sc_hd__o21ai_4
XPHY_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2191_ _2545_/Q _1739_/B _2190_/Y _2168_/Y vssd1 vssd1 vccd1 vccd1 _2191_/Y sky130_fd_sc_hd__a22oi_4
XFILLER_49_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1211_ _2645_/Q _1194_/B _1210_/X vssd1 vssd1 vccd1 vccd1 _1211_/Y sky130_fd_sc_hd__o21ai_4
X_2260_ _1840_/B _1698_/A _2144_/A vssd1 vssd1 vccd1 vccd1 _2260_/Y sky130_fd_sc_hd__nand3_4
XFILLER_18_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1975_ _1869_/A _1867_/Y _1975_/C vssd1 vssd1 vccd1 vccd1 _1975_/Y sky130_fd_sc_hd__nor3_4
X_2458_ _2646_/CLK _2458_/D vssd1 vssd1 vccd1 vccd1 _2105_/B sky130_fd_sc_hd__dfxtp_4
X_1409_ _1409_/A _2614_/Q _1406_/X vssd1 vssd1 vccd1 vccd1 _1409_/Y sky130_fd_sc_hd__nand3_4
X_2527_ _2527_/CLK _2527_/D vssd1 vssd1 vccd1 vccd1 _2527_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_45_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2389_ _2389_/CLK _2389_/D vssd1 vssd1 vccd1 vccd1 _1577_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_28_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_4_0_0_addressalyzerBlock.SPI_CLK clkbuf_3_0_0_addressalyzerBlock.SPI_CLK/X
+ vssd1 vssd1 vccd1 vccd1 _2418_/CLK sky130_fd_sc_hd__clkbuf_1
X_1760_ _1758_/Y _1759_/Y _2168_/A vssd1 vssd1 vccd1 vccd1 _1760_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_30_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1691_ _2594_/Q vssd1 vssd1 vccd1 vccd1 _2289_/C sky130_fd_sc_hd__inv_2
X_2312_ _1606_/Y _1190_/A _1581_/A _1694_/X vssd1 vssd1 vccd1 vccd1 _2312_/X sky130_fd_sc_hd__and4_4
XFILLER_65_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2174_ _2196_/A _2174_/B vssd1 vssd1 vccd1 vccd1 _2174_/Y sky130_fd_sc_hd__nand2_4
X_2243_ _1606_/Y vssd1 vssd1 vccd1 vccd1 _2243_/Y sky130_fd_sc_hd__inv_2
XFILLER_21_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1889_ _1888_/A _2560_/Q vssd1 vssd1 vccd1 vccd1 _2552_/D sky130_fd_sc_hd__and2_4
X_1958_ _1969_/A _2516_/Q vssd1 vssd1 vccd1 vccd1 _1958_/X sky130_fd_sc_hd__and2_4
Xclkbuf_3_5_0_addressalyzerBlock.SPI_CLK clkbuf_3_5_0_addressalyzerBlock.SPI_CLK/A
+ vssd1 vssd1 vccd1 vccd1 clkbuf_3_5_0_addressalyzerBlock.SPI_CLK/X sky130_fd_sc_hd__clkbuf_1
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1674_ _1658_/Y _1661_/X _1861_/B vssd1 vssd1 vccd1 vccd1 _1674_/Y sky130_fd_sc_hd__nand3_4
X_1812_ _2578_/Q _1809_/X _1811_/X vssd1 vssd1 vccd1 vccd1 _1812_/X sky130_fd_sc_hd__o21a_4
X_1743_ _2415_/Q vssd1 vssd1 vccd1 vccd1 _1744_/B sky130_fd_sc_hd__inv_2
X_2226_ _2222_/X _2225_/X _1472_/A vssd1 vssd1 vccd1 vccd1 _2226_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_53_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2088_ _1289_/B _2469_/Q vssd1 vssd1 vccd1 vccd1 _2088_/X sky130_fd_sc_hd__and2_4
XFILLER_13_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2157_ _2153_/Y _2156_/Y _1628_/X vssd1 vssd1 vccd1 vccd1 _2157_/X sky130_fd_sc_hd__a21o_4
XFILLER_44_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1390_ _2019_/A _1390_/B _1389_/Y vssd1 vssd1 vccd1 vccd1 _1390_/Y sky130_fd_sc_hd__nor3_4
XFILLER_4_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2011_ _2011_/A vssd1 vssd1 vccd1 vccd1 _2013_/C sky130_fd_sc_hd__inv_2
X_1726_ _1676_/A _1726_/B vssd1 vssd1 vccd1 vccd1 _1727_/B sky130_fd_sc_hd__nand2_4
X_1657_ _1612_/X _2628_/Q _1656_/X vssd1 vssd1 vccd1 vccd1 _1657_/Y sky130_fd_sc_hd__a21oi_4
X_1588_ _2335_/D _1460_/X _1514_/X vssd1 vssd1 vccd1 vccd1 _1588_/Y sky130_fd_sc_hd__o21ai_4
X_2209_ _1741_/A _2622_/Q _1655_/A vssd1 vssd1 vccd1 vccd1 _2209_/X sky130_fd_sc_hd__a21o_4
XFILLER_37_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2491_ _2492_/CLK _2019_/Y vssd1 vssd1 vccd1 vccd1 _2011_/A sky130_fd_sc_hd__dfxtp_4
X_1442_ _1434_/Y _1422_/A _1184_/A vssd1 vssd1 vccd1 vccd1 _1530_/A sky130_fd_sc_hd__a21o_4
X_2560_ _2552_/CLK _1879_/X vssd1 vssd1 vccd1 vccd1 _2560_/Q sky130_fd_sc_hd__dfxtp_4
X_1511_ _1487_/B vssd1 vssd1 vccd1 vccd1 _1511_/Y sky130_fd_sc_hd__inv_2
X_1373_ _1385_/B _1376_/C _1383_/C _1365_/D vssd1 vssd1 vccd1 vccd1 _1373_/X sky130_fd_sc_hd__and4_4
XFILLER_31_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1709_ _2433_/Q vssd1 vssd1 vccd1 vccd1 _1710_/B sky130_fd_sc_hd__inv_2
XFILLER_54_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1991_ _1991_/A _1991_/B _2473_/Q _2474_/Q vssd1 vssd1 vccd1 vccd1 _2059_/A sky130_fd_sc_hd__nand4_4
X_2612_ _2588_/CLK _1455_/Y vssd1 vssd1 vccd1 vccd1 _2335_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_9_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2543_ _2464_/CLK _2543_/D vssd1 vssd1 vccd1 vccd1 _2543_/Q sky130_fd_sc_hd__dfxtp_4
X_2474_ _2476_/CLK _2474_/D vssd1 vssd1 vccd1 vccd1 _2474_/Q sky130_fd_sc_hd__dfxtp_4
X_1425_ _2600_/Q vssd1 vssd1 vccd1 vccd1 _1570_/A sky130_fd_sc_hd__buf_2
X_1356_ _1351_/Y vssd1 vssd1 vccd1 vccd1 _1358_/A sky130_fd_sc_hd__inv_2
XFILLER_36_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1287_ _1277_/B vssd1 vssd1 vccd1 vccd1 _1289_/A sky130_fd_sc_hd__inv_2
XPHY_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1210_ _1206_/A _1833_/A vssd1 vssd1 vccd1 vccd1 _1210_/X sky130_fd_sc_hd__or2_4
X_2190_ _2172_/Y _2188_/Y _2189_/Y vssd1 vssd1 vccd1 vccd1 _2190_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_37_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1974_ _1972_/Y _1973_/A _1973_/Y vssd1 vssd1 vccd1 vccd1 _1975_/C sky130_fd_sc_hd__a21oi_4
XFILLER_60_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2457_ _2454_/CLK _2457_/D vssd1 vssd1 vccd1 vccd1 _2457_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_56_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1408_ _2019_/A _1401_/Y _1407_/Y vssd1 vssd1 vccd1 vccd1 _2616_/D sky130_fd_sc_hd__nor3_4
X_2388_ _2646_/CLK _2388_/D vssd1 vssd1 vccd1 vccd1 _1729_/B sky130_fd_sc_hd__dfxtp_4
X_2526_ _2527_/CLK _2526_/D vssd1 vssd1 vccd1 vccd1 MACRO_RD_SELECT[3] sky130_fd_sc_hd__dfxtp_4
XFILLER_43_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1339_ _1274_/X vssd1 vssd1 vccd1 vccd1 _1339_/X sky130_fd_sc_hd__buf_2
XPHY_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1690_ _1697_/A _1687_/A _1689_/Y vssd1 vssd1 vccd1 vccd1 _1690_/Y sky130_fd_sc_hd__nor3_4
X_2242_ _2122_/Y _2241_/A _2241_/Y vssd1 vssd1 vccd1 vccd1 _2434_/D sky130_fd_sc_hd__o21ai_4
X_2311_ _2310_/X vssd1 vssd1 vccd1 vccd1 _2311_/X sky130_fd_sc_hd__buf_2
X_2173_ _1534_/A _2553_/Q _2148_/X vssd1 vssd1 vccd1 vccd1 _2173_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_15_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1957_ _1969_/A _1957_/B vssd1 vssd1 vccd1 vccd1 _2509_/D sky130_fd_sc_hd__and2_4
X_1888_ _1888_/A _2561_/Q vssd1 vssd1 vccd1 vccd1 _2553_/D sky130_fd_sc_hd__and2_4
X_2509_ _2519_/CLK _2509_/D vssd1 vssd1 vccd1 vccd1 DATA_TO_HASH[2] sky130_fd_sc_hd__dfxtp_4
XFILLER_56_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1811_ _2579_/Q _1810_/X _1799_/X vssd1 vssd1 vccd1 vccd1 _1811_/X sky130_fd_sc_hd__o21a_4
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1673_ _1761_/A _1673_/B _2168_/A _1739_/B vssd1 vssd1 vccd1 vccd1 _1861_/B sky130_fd_sc_hd__nor4_4
X_1742_ _1316_/B _1646_/X _1741_/Y vssd1 vssd1 vccd1 vccd1 _1742_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_7_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2225_ _2439_/Q _1751_/A _1633_/X _2224_/Y vssd1 vssd1 vccd1 vccd1 _2225_/X sky130_fd_sc_hd__a211o_4
XFILLER_53_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2087_ _1284_/X _2079_/A vssd1 vssd1 vccd1 vccd1 _2087_/Y sky130_fd_sc_hd__nor2_4
X_2156_ _2154_/Y _2201_/B _2156_/C vssd1 vssd1 vccd1 vccd1 _2156_/Y sky130_fd_sc_hd__nand3_4
XFILLER_21_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2010_ _2009_/X _2010_/B _2010_/C vssd1 vssd1 vccd1 vccd1 _2492_/D sky130_fd_sc_hd__and3_4
XFILLER_35_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_3_2_0_m1_clk_local clkbuf_3_3_0_m1_clk_local/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_2_0_m1_clk_local/X
+ sky130_fd_sc_hd__clkbuf_1
X_1725_ _1722_/Y _1723_/Y _1724_/X vssd1 vssd1 vccd1 vccd1 _1725_/X sky130_fd_sc_hd__a21o_4
X_1656_ _1656_/A vssd1 vssd1 vccd1 vccd1 _1656_/X sky130_fd_sc_hd__buf_2
X_1587_ _1545_/X _1576_/X _1578_/Y _1582_/Y _1586_/X vssd1 vssd1 vccd1 vccd1 _1587_/Y
+ sky130_fd_sc_hd__a41oi_4
XFILLER_7_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2208_ _2630_/Q _1645_/Y _1741_/Y vssd1 vssd1 vccd1 vccd1 _2208_/X sky130_fd_sc_hd__o21a_4
XFILLER_37_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2139_ _1594_/X _1581_/A _1669_/B _2121_/X _2101_/A vssd1 vssd1 vccd1 vccd1 _2139_/X
+ sky130_fd_sc_hd__a41o_4
XFILLER_1_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2490_ _2470_/CLK _2490_/D vssd1 vssd1 vccd1 vccd1 _1999_/A sky130_fd_sc_hd__dfxtp_4
X_1441_ _1420_/Y _1445_/D _1440_/Y vssd1 vssd1 vccd1 vccd1 _1441_/Y sky130_fd_sc_hd__o21ai_4
X_1510_ _1507_/Y _1509_/X _1454_/X vssd1 vssd1 vccd1 vccd1 _1510_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_4_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1372_ _1236_/B vssd1 vssd1 vccd1 vccd1 _1376_/C sky130_fd_sc_hd__buf_2
XFILLER_2_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1708_ _2448_/Q vssd1 vssd1 vccd1 vccd1 _1708_/X sky130_fd_sc_hd__buf_2
X_1639_ _1629_/X _1638_/X _1472_/A vssd1 vssd1 vccd1 vccd1 _1639_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_46_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1990_ _2071_/A _2476_/Q vssd1 vssd1 vccd1 vccd1 _1990_/Y sky130_fd_sc_hd__nand2_4
XFILLER_45_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2542_ _2538_/CLK _2542_/D vssd1 vssd1 vccd1 vccd1 _2542_/Q sky130_fd_sc_hd__dfxtp_4
X_2611_ _2611_/CLK _2611_/D vssd1 vssd1 vccd1 vccd1 _1438_/B sky130_fd_sc_hd__dfxtp_4
X_1355_ _1354_/Y vssd1 vssd1 vccd1 vccd1 _1355_/Y sky130_fd_sc_hd__inv_2
X_2473_ _2476_/CLK _2473_/D vssd1 vssd1 vccd1 vccd1 _2473_/Q sky130_fd_sc_hd__dfxtp_4
X_1424_ _1424_/A vssd1 vssd1 vccd1 vccd1 _1424_/Y sky130_fd_sc_hd__inv_2
XFILLER_63_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1286_ _1284_/X _1261_/Y _1286_/C vssd1 vssd1 vccd1 vccd1 _1286_/Y sky130_fd_sc_hd__nor3_4
XPHY_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_5_0_addressalyzerBlock.SPI_CLK clkbuf_3_2_0_addressalyzerBlock.SPI_CLK/X
+ vssd1 vssd1 vccd1 vccd1 _2551_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_37_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1973_ _1973_/A _1973_/B vssd1 vssd1 vccd1 vccd1 _1973_/Y sky130_fd_sc_hd__nor2_4
XFILLER_60_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2525_ _2521_/CLK _2525_/D vssd1 vssd1 vccd1 vccd1 MACRO_RD_SELECT[2] sky130_fd_sc_hd__dfxtp_4
X_2456_ _2454_/CLK _2456_/D vssd1 vssd1 vccd1 vccd1 _2456_/Q sky130_fd_sc_hd__dfxtp_4
X_1407_ _1409_/A _2615_/Q _2614_/Q _1406_/X _1230_/A vssd1 vssd1 vccd1 vccd1 _1407_/Y
+ sky130_fd_sc_hd__a41oi_4
X_2387_ _2646_/CLK _2327_/Y vssd1 vssd1 vccd1 vccd1 _1683_/A sky130_fd_sc_hd__dfxtp_4
X_1338_ _1353_/A _1335_/D _1329_/X _1321_/X vssd1 vssd1 vccd1 vccd1 _1338_/X sky130_fd_sc_hd__and4_4
X_1269_ _1269_/A vssd1 vssd1 vccd1 vccd1 _1346_/A sky130_fd_sc_hd__buf_2
XFILLER_36_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2172_ _2615_/Q _1571_/A _1568_/A _1660_/A _2146_/Y vssd1 vssd1 vccd1 vccd1 _2172_/Y
+ sky130_fd_sc_hd__o41ai_4
XFILLER_38_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2310_ _1594_/X _1597_/X _1581_/A _1696_/A _1736_/A vssd1 vssd1 vccd1 vccd1 _2310_/X
+ sky130_fd_sc_hd__a41o_4
X_2241_ _2241_/A _2300_/B _2434_/Q vssd1 vssd1 vccd1 vccd1 _2241_/Y sky130_fd_sc_hd__nand3_4
XFILLER_18_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1887_ _1888_/A _2562_/Q vssd1 vssd1 vccd1 vccd1 _2554_/D sky130_fd_sc_hd__and2_4
X_1956_ _1254_/X vssd1 vssd1 vccd1 vccd1 _1969_/A sky130_fd_sc_hd__buf_2
XFILLER_21_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2508_ _2508_/CLK _1958_/X vssd1 vssd1 vccd1 vccd1 DATA_TO_HASH[1] sky130_fd_sc_hd__dfxtp_4
XFILLER_0_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2439_ _2552_/CLK _2145_/Y vssd1 vssd1 vccd1 vccd1 _2439_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1741_ _1741_/A vssd1 vssd1 vccd1 vccd1 _1741_/Y sky130_fd_sc_hd__inv_2
XFILLER_30_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1810_ _2461_/Q vssd1 vssd1 vccd1 vccd1 _1810_/X sky130_fd_sc_hd__buf_2
X_1672_ _2168_/B vssd1 vssd1 vccd1 vccd1 _1739_/B sky130_fd_sc_hd__buf_2
XFILLER_7_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2155_ _2155_/A _1634_/X vssd1 vssd1 vccd1 vccd1 _2156_/C sky130_fd_sc_hd__nand2_4
X_2224_ _2224_/A _2224_/B vssd1 vssd1 vccd1 vccd1 _2224_/Y sky130_fd_sc_hd__nor2_4
X_2086_ _2079_/A _1991_/B _2085_/Y vssd1 vssd1 vccd1 vccd1 _2086_/X sky130_fd_sc_hd__o21a_4
X_1939_ _1938_/A _1847_/Y vssd1 vssd1 vccd1 vccd1 _1939_/Y sky130_fd_sc_hd__nor2_4
XFILLER_44_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0_addressalyzerBlock.SPI_CLK clkbuf_0_addressalyzerBlock.SPI_CLK/X vssd1
+ vssd1 vccd1 vccd1 clkbuf_2_3_0_addressalyzerBlock.SPI_CLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_4_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1724_ _1559_/Y _1856_/A _1663_/A _2168_/B vssd1 vssd1 vccd1 vccd1 _1724_/X sky130_fd_sc_hd__a211o_4
X_1655_ _1655_/A vssd1 vssd1 vccd1 vccd1 _1656_/A sky130_fd_sc_hd__buf_2
X_1586_ _1541_/X _1583_/X _1781_/A vssd1 vssd1 vccd1 vccd1 _1586_/X sky130_fd_sc_hd__a21o_4
X_2069_ _2058_/X _2060_/Y _2068_/Y vssd1 vssd1 vccd1 vccd1 _2070_/A sky130_fd_sc_hd__o21ai_4
X_2207_ _2195_/Y _2205_/Y _2206_/Y vssd1 vssd1 vccd1 vccd1 _2207_/Y sky130_fd_sc_hd__o21ai_4
X_2138_ _2138_/A vssd1 vssd1 vccd1 vccd1 _2138_/Y sky130_fd_sc_hd__inv_2
XFILLER_53_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1371_ _1360_/Y _1361_/B _1370_/Y vssd1 vssd1 vccd1 vccd1 _1371_/Y sky130_fd_sc_hd__a21oi_4
X_1440_ _2326_/B _1440_/B _1488_/A _1439_/X vssd1 vssd1 vccd1 vccd1 _1440_/Y sky130_fd_sc_hd__nand4_4
XFILLER_4_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1707_ _2295_/C _2224_/A _2201_/B _1706_/Y vssd1 vssd1 vccd1 vccd1 _1707_/X sky130_fd_sc_hd__a211o_4
X_1638_ _2125_/C _1751_/A _1633_/X _1637_/Y vssd1 vssd1 vccd1 vccd1 _1638_/X sky130_fd_sc_hd__a211o_4
XFILLER_58_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1569_ _1731_/B _1566_/X _1661_/C vssd1 vssd1 vccd1 vccd1 _1569_/X sky130_fd_sc_hd__o21a_4
XFILLER_66_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2472_ _2476_/CLK _2086_/X vssd1 vssd1 vccd1 vccd1 _1991_/B sky130_fd_sc_hd__dfxtp_4
X_2541_ _2538_/CLK _1905_/Y vssd1 vssd1 vccd1 vccd1 _1917_/B sky130_fd_sc_hd__dfxtp_4
X_2610_ _2611_/CLK _2610_/D vssd1 vssd1 vccd1 vccd1 _1438_/C sky130_fd_sc_hd__dfxtp_4
XFILLER_48_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1354_ _1352_/X _1353_/Y vssd1 vssd1 vccd1 vccd1 _1354_/Y sky130_fd_sc_hd__nand2_4
X_1285_ _1225_/X _1226_/Y _1265_/A _1246_/Y _1256_/Y vssd1 vssd1 vccd1 vccd1 _1286_/C
+ sky130_fd_sc_hd__o41a_4
X_1423_ _2335_/B vssd1 vssd1 vccd1 vccd1 _2326_/B sky130_fd_sc_hd__inv_2
XFILLER_51_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_10_0_addressalyzerBlock.SPI_CLK clkbuf_3_5_0_addressalyzerBlock.SPI_CLK/X
+ vssd1 vssd1 vccd1 vccd1 _2611_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_54_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1972_ _1972_/A _1972_/B _2497_/Q vssd1 vssd1 vccd1 vccd1 _1972_/Y sky130_fd_sc_hd__nand3_4
XFILLER_33_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2455_ _2454_/CLK _2455_/D vssd1 vssd1 vccd1 vccd1 _2455_/Q sky130_fd_sc_hd__dfxtp_4
X_2524_ _2521_/CLK _2524_/D vssd1 vssd1 vccd1 vccd1 MACRO_RD_SELECT[1] sky130_fd_sc_hd__dfxtp_4
X_1406_ _1406_/A vssd1 vssd1 vccd1 vccd1 _1406_/X sky130_fd_sc_hd__buf_2
X_2386_ _2646_/CLK _2329_/Y vssd1 vssd1 vccd1 vccd1 _2386_/Q sky130_fd_sc_hd__dfxtp_4
X_1337_ _1337_/A vssd1 vssd1 vccd1 vccd1 _1337_/Y sky130_fd_sc_hd__inv_2
X_1268_ _1266_/Y _1719_/A vssd1 vssd1 vccd1 vccd1 _1271_/A sky130_fd_sc_hd__nand2_4
X_1199_ _1194_/A _1179_/X _1198_/X vssd1 vssd1 vccd1 vccd1 _1199_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_51_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2171_ _1676_/A _2169_/Y _2170_/Y vssd1 vssd1 vccd1 vccd1 _2171_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_2_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2240_ _1555_/A vssd1 vssd1 vccd1 vccd1 _2300_/B sky130_fd_sc_hd__buf_2
XFILLER_65_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1886_ _1886_/A vssd1 vssd1 vccd1 vccd1 _1888_/A sky130_fd_sc_hd__buf_2
X_1955_ _1954_/A _2518_/Q vssd1 vssd1 vccd1 vccd1 _2510_/D sky130_fd_sc_hd__and2_4
X_2438_ _2464_/CLK _2171_/Y vssd1 vssd1 vccd1 vccd1 _2170_/B sky130_fd_sc_hd__dfxtp_4
X_2507_ _2635_/CLK _2507_/D vssd1 vssd1 vccd1 vccd1 DATA_TO_HASH[0] sky130_fd_sc_hd__dfxtp_4
X_2369_ _2374_/CLK _2369_/D vssd1 vssd1 vccd1 vccd1 _2369_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_56_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1740_ _1739_/Y vssd1 vssd1 vccd1 vccd1 _1740_/Y sky130_fd_sc_hd__inv_2
X_1671_ _1571_/A _1660_/A _2234_/D vssd1 vssd1 vccd1 vccd1 _2168_/B sky130_fd_sc_hd__nor3_4
XFILLER_30_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2085_ _2079_/A _1991_/B _2063_/A vssd1 vssd1 vccd1 vccd1 _2085_/Y sky130_fd_sc_hd__a21oi_4
X_2223_ _1767_/B vssd1 vssd1 vccd1 vccd1 _2224_/B sky130_fd_sc_hd__inv_2
X_2154_ _2196_/A _2154_/B vssd1 vssd1 vccd1 vccd1 _2154_/Y sky130_fd_sc_hd__nand2_4
XFILLER_61_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1869_ _1869_/A _1868_/Y vssd1 vssd1 vccd1 vccd1 _2567_/D sky130_fd_sc_hd__nor2_4
X_1938_ _1938_/A _1937_/Y vssd1 vssd1 vccd1 vccd1 _1938_/Y sky130_fd_sc_hd__nor2_4
XFILLER_29_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1723_ _1656_/X _2619_/Q _1673_/B vssd1 vssd1 vccd1 vccd1 _1723_/Y sky130_fd_sc_hd__a21oi_4
X_1654_ _1570_/A _1568_/A _1659_/A vssd1 vssd1 vccd1 vccd1 _1655_/A sky130_fd_sc_hd__nor3_4
XFILLER_7_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1585_ _1736_/A vssd1 vssd1 vccd1 vccd1 _1781_/A sky130_fd_sc_hd__buf_2
X_2206_ _1293_/Y _1613_/Y _1605_/X _1649_/Y vssd1 vssd1 vccd1 vccd1 _2206_/Y sky130_fd_sc_hd__a2bb2oi_4
XFILLER_66_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2068_ _2060_/Y _2058_/X _1388_/A vssd1 vssd1 vccd1 vccd1 _2068_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_26_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2137_ _2101_/A _2289_/C vssd1 vssd1 vccd1 vccd1 _2138_/A sky130_fd_sc_hd__nor2_4
XFILLER_17_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1370_ _1360_/Y _1361_/B _1346_/X vssd1 vssd1 vccd1 vccd1 _1370_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_4_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1706_ _1630_/X _1706_/B vssd1 vssd1 vccd1 vccd1 _1706_/Y sky130_fd_sc_hd__nor2_4
X_1637_ _1635_/X _1636_/Y vssd1 vssd1 vccd1 vccd1 _1637_/Y sky130_fd_sc_hd__nor2_4
XFILLER_58_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1568_ _1568_/A vssd1 vssd1 vccd1 vccd1 _1661_/C sky130_fd_sc_hd__buf_2
X_1499_ _1487_/A vssd1 vssd1 vccd1 vccd1 _1499_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2471_ _2476_/CLK _2087_/Y vssd1 vssd1 vccd1 vccd1 _1991_/A sky130_fd_sc_hd__dfxtp_4
X_1422_ _1422_/A vssd1 vssd1 vccd1 vccd1 _1445_/D sky130_fd_sc_hd__buf_2
XFILLER_9_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2540_ _2538_/CLK _1907_/Y vssd1 vssd1 vccd1 vccd1 _2540_/Q sky130_fd_sc_hd__dfxtp_4
X_1353_ _1353_/A _2628_/Q _1349_/A vssd1 vssd1 vccd1 vccd1 _1353_/Y sky130_fd_sc_hd__nand3_4
X_1284_ _1388_/A vssd1 vssd1 vccd1 vccd1 _1284_/X sky130_fd_sc_hd__buf_2
XFILLER_63_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1971_ _1289_/B _1971_/B vssd1 vssd1 vccd1 vccd1 _1971_/X sky130_fd_sc_hd__and2_4
X_2454_ _2454_/CLK _2454_/D vssd1 vssd1 vccd1 vccd1 _2454_/Q sky130_fd_sc_hd__dfxtp_4
X_2385_ _2646_/CLK _2339_/X vssd1 vssd1 vccd1 vccd1 _2385_/Q sky130_fd_sc_hd__dfxtp_4
X_1405_ _1232_/A vssd1 vssd1 vccd1 vccd1 _1409_/A sky130_fd_sc_hd__buf_2
X_2523_ _2513_/CLK _1934_/X vssd1 vssd1 vccd1 vccd1 MACRO_RD_SELECT[0] sky130_fd_sc_hd__dfxtp_4
X_1198_ _1202_/A _1198_/B vssd1 vssd1 vccd1 vccd1 _1198_/X sky130_fd_sc_hd__or2_4
X_1336_ _1331_/X _1335_/Y vssd1 vssd1 vccd1 vccd1 _1337_/A sky130_fd_sc_hd__nand2_4
XFILLER_28_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1267_ _1267_/A vssd1 vssd1 vccd1 vccd1 _1719_/A sky130_fd_sc_hd__inv_2
XFILLER_24_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_0_addressalyzerBlock.SPI_CLK _2347_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0_addressalyzerBlock.SPI_CLK/X
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_10_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2170_ _2192_/A _2170_/B vssd1 vssd1 vccd1 vccd1 _2170_/Y sky130_fd_sc_hd__nand2_4
X_1954_ _1954_/A _2519_/Q vssd1 vssd1 vccd1 vccd1 _1954_/X sky130_fd_sc_hd__and2_4
XFILLER_18_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_2_1_0_addressalyzerBlock.SPI_CLK clkbuf_2_1_0_addressalyzerBlock.SPI_CLK/A
+ vssd1 vssd1 vccd1 vccd1 clkbuf_3_3_0_addressalyzerBlock.SPI_CLK/A sky130_fd_sc_hd__clkbuf_1
X_1885_ _1885_/A _2563_/Q vssd1 vssd1 vccd1 vccd1 _2555_/D sky130_fd_sc_hd__and2_4
X_2368_ _2374_/CLK _2367_/Q vssd1 vssd1 vccd1 vccd1 _2369_/D sky130_fd_sc_hd__dfxtp_4
X_2437_ _2437_/CLK _2193_/Y vssd1 vssd1 vccd1 vccd1 _2192_/B sky130_fd_sc_hd__dfxtp_4
Xclkbuf_4_7_0_m1_clk_local clkbuf_3_3_0_m1_clk_local/X vssd1 vssd1 vccd1 vccd1 _2505_/CLK
+ sky130_fd_sc_hd__clkbuf_1
X_2506_ _2505_/CLK _1961_/Y vssd1 vssd1 vccd1 vccd1 _1968_/B sky130_fd_sc_hd__dfxtp_4
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1319_ _1317_/X _1318_/Y vssd1 vssd1 vccd1 vccd1 _1320_/A sky130_fd_sc_hd__nand2_4
XFILLER_44_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2299_ _2268_/Y _2291_/X _2298_/Y vssd1 vssd1 vccd1 vccd1 _2408_/D sky130_fd_sc_hd__o21ai_4
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1670_ _1669_/Y vssd1 vssd1 vccd1 vccd1 _2234_/D sky130_fd_sc_hd__inv_2
XFILLER_7_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2222_ _2219_/Y _2221_/Y _1628_/X vssd1 vssd1 vccd1 vccd1 _2222_/X sky130_fd_sc_hd__a21o_4
X_2084_ _2083_/X _2057_/B _2084_/C vssd1 vssd1 vccd1 vccd1 _2473_/D sky130_fd_sc_hd__and3_4
X_2153_ _2151_/Y _1708_/X _2153_/C vssd1 vssd1 vccd1 vccd1 _2153_/Y sky130_fd_sc_hd__nand3_4
X_1937_ _2425_/Q vssd1 vssd1 vccd1 vccd1 _1937_/Y sky130_fd_sc_hd__inv_2
X_1868_ _1868_/A _1867_/Y vssd1 vssd1 vccd1 vccd1 _1868_/Y sky130_fd_sc_hd__xnor2_4
X_1799_ _1555_/A vssd1 vssd1 vccd1 vccd1 _1799_/X sky130_fd_sc_hd__buf_2
XFILLER_40_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1722_ _1700_/X _1720_/Y _1721_/Y vssd1 vssd1 vccd1 vccd1 _1722_/Y sky130_fd_sc_hd__o21ai_4
X_1584_ _1219_/X vssd1 vssd1 vccd1 vccd1 _1736_/A sky130_fd_sc_hd__buf_2
X_1653_ _1642_/Y _1646_/X _1652_/X vssd1 vssd1 vccd1 vccd1 _1653_/Y sky130_fd_sc_hd__a21oi_4
X_2205_ _2202_/X _2204_/X _1701_/A vssd1 vssd1 vccd1 vccd1 _2205_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_66_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2067_ _2063_/A _1993_/B _2067_/C vssd1 vssd1 vccd1 vccd1 _2067_/Y sky130_fd_sc_hd__nor3_4
XFILLER_34_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2136_ _2136_/A vssd1 vssd1 vccd1 vccd1 _2136_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1705_ _2417_/Q vssd1 vssd1 vccd1 vccd1 _1706_/B sky130_fd_sc_hd__inv_2
X_1567_ _1567_/A _1567_/B _1567_/C vssd1 vssd1 vccd1 vccd1 _1568_/A sky130_fd_sc_hd__nand3_4
X_1636_ _2402_/Q vssd1 vssd1 vccd1 vccd1 _1636_/Y sky130_fd_sc_hd__inv_2
X_1498_ _2136_/A _2333_/B _1462_/X vssd1 vssd1 vccd1 vccd1 _1498_/Y sky130_fd_sc_hd__a21oi_4
X_2119_ _2119_/A vssd1 vssd1 vccd1 vccd1 _2120_/A sky130_fd_sc_hd__inv_2
XFILLER_13_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_4_15_0_addressalyzerBlock.SPI_CLK clkbuf_3_7_0_addressalyzerBlock.SPI_CLK/X
+ vssd1 vssd1 vccd1 vccd1 _2454_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_49_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2470_ _2470_/CLK _2088_/X vssd1 vssd1 vccd1 vccd1 HASH_EN sky130_fd_sc_hd__dfxtp_4
X_1421_ _2390_/Q vssd1 vssd1 vccd1 vccd1 _1422_/A sky130_fd_sc_hd__inv_2
XFILLER_63_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1283_ _2364_/D vssd1 vssd1 vccd1 vccd1 _1388_/A sky130_fd_sc_hd__buf_2
XFILLER_48_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1352_ _2628_/Q _1351_/Y _1306_/X vssd1 vssd1 vccd1 vccd1 _1352_/X sky130_fd_sc_hd__o21a_4
X_2599_ _2437_/CLK _1587_/Y vssd1 vssd1 vccd1 vccd1 _1567_/A sky130_fd_sc_hd__dfxtp_4
X_1619_ _1619_/A vssd1 vssd1 vccd1 vccd1 _1619_/Y sky130_fd_sc_hd__inv_2
XFILLER_54_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1970_ _1289_/B _1970_/B vssd1 vssd1 vccd1 vccd1 _2500_/D sky130_fd_sc_hd__and2_4
X_2522_ _2513_/CLK _2522_/D vssd1 vssd1 vccd1 vccd1 _2522_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_4_15_0_m1_clk_local clkbuf_3_7_0_m1_clk_local/X vssd1 vssd1 vccd1 vccd1 _2508_/CLK
+ sky130_fd_sc_hd__clkbuf_1
X_2384_ _2464_/CLK _2384_/D vssd1 vssd1 vccd1 vccd1 _2384_/Q sky130_fd_sc_hd__dfxtp_4
X_1404_ _1404_/A vssd1 vssd1 vccd1 vccd1 _1404_/Y sky130_fd_sc_hd__inv_2
X_2453_ _2646_/CLK _2111_/Y vssd1 vssd1 vccd1 vccd1 _2099_/C sky130_fd_sc_hd__dfxtp_4
X_1335_ _2632_/Q _1333_/Y _1335_/C _1335_/D vssd1 vssd1 vccd1 vccd1 _1335_/Y sky130_fd_sc_hd__nand4_4
XFILLER_56_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1197_ _1195_/Y _1187_/X _1196_/Y vssd1 vssd1 vccd1 vccd1 _1197_/Y sky130_fd_sc_hd__a21oi_4
X_1266_ _1256_/A _1265_/Y _1224_/A _1249_/Y vssd1 vssd1 vccd1 vccd1 _1266_/Y sky130_fd_sc_hd__nand4_4
XPHY_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1884_ _1885_/A _1884_/B vssd1 vssd1 vccd1 vccd1 _1884_/X sky130_fd_sc_hd__and2_4
X_1953_ _1954_/A _2520_/Q vssd1 vssd1 vccd1 vccd1 _2512_/D sky130_fd_sc_hd__and2_4
XFILLER_21_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2505_ _2505_/CLK _2505_/D vssd1 vssd1 vccd1 vccd1 _2505_/Q sky130_fd_sc_hd__dfxtp_4
X_2367_ _2492_/CLK _2367_/D vssd1 vssd1 vccd1 vccd1 _2367_/Q sky130_fd_sc_hd__dfxtp_4
X_2436_ _2437_/CLK _2436_/D vssd1 vssd1 vccd1 vccd1 _2436_/Q sky130_fd_sc_hd__dfxtp_4
X_1318_ _1856_/B _1318_/B _1316_/B _1316_/D vssd1 vssd1 vccd1 vccd1 _1318_/Y sky130_fd_sc_hd__nand4_4
X_2298_ _2304_/A _2300_/B ID_toHost vssd1 vssd1 vccd1 vccd1 _2298_/Y sky130_fd_sc_hd__nand3_4
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1249_ _1249_/A vssd1 vssd1 vccd1 vccd1 _1249_/Y sky130_fd_sc_hd__inv_2
XFILLER_24_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2221_ _1948_/Y _1624_/X _2220_/Y vssd1 vssd1 vccd1 vccd1 _2221_/Y sky130_fd_sc_hd__o21ai_4
X_2152_ HASH_LED _1618_/X vssd1 vssd1 vccd1 vccd1 _2153_/C sky130_fd_sc_hd__nand2_4
XFILLER_53_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2083_ _2079_/A _1991_/B _2473_/Q vssd1 vssd1 vccd1 vccd1 _2083_/X sky130_fd_sc_hd__a21o_4
XFILLER_38_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1867_ _1973_/A _2497_/Q _1973_/B vssd1 vssd1 vccd1 vccd1 _1867_/Y sky130_fd_sc_hd__nor3_4
X_1936_ _1938_/A _1622_/Y vssd1 vssd1 vccd1 vccd1 _2522_/D sky130_fd_sc_hd__nor2_4
X_1798_ _1983_/B _2576_/Q _1797_/X vssd1 vssd1 vccd1 vccd1 _1798_/X sky130_fd_sc_hd__o21a_4
XFILLER_29_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2419_ _2555_/CLK _2419_/D vssd1 vssd1 vccd1 vccd1 _2419_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_37_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1721_ _1612_/X _1351_/A _1656_/X vssd1 vssd1 vccd1 vccd1 _1721_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_43_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1652_ _1856_/A _2636_/Q _1856_/C vssd1 vssd1 vccd1 vccd1 _1652_/X sky130_fd_sc_hd__and3_4
X_1583_ _1604_/A vssd1 vssd1 vccd1 vccd1 _1583_/X sky130_fd_sc_hd__buf_2
XFILLER_7_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2135_ _2120_/X _2133_/Y _2134_/Y vssd1 vssd1 vccd1 vccd1 _2443_/D sky130_fd_sc_hd__o21ai_4
X_2204_ _2440_/Q _1635_/X _1632_/Y _2203_/Y vssd1 vssd1 vccd1 vccd1 _2204_/X sky130_fd_sc_hd__a211o_4
X_2066_ _2060_/Y _2058_/X _2062_/B vssd1 vssd1 vccd1 vccd1 _2067_/C sky130_fd_sc_hd__a21oi_4
XFILLER_26_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1919_ _1918_/A _1919_/B vssd1 vssd1 vccd1 vccd1 _2533_/D sky130_fd_sc_hd__and2_4
XFILLER_57_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1704_ _1704_/A vssd1 vssd1 vccd1 vccd1 _2201_/B sky130_fd_sc_hd__buf_2
X_1566_ _1729_/B vssd1 vssd1 vccd1 vccd1 _1566_/X sky130_fd_sc_hd__buf_2
X_1497_ _2583_/Q vssd1 vssd1 vccd1 vccd1 _2136_/A sky130_fd_sc_hd__buf_2
X_1635_ _1634_/X vssd1 vssd1 vccd1 vccd1 _1635_/X sky130_fd_sc_hd__buf_2
X_2049_ _2049_/A _2022_/B _2048_/Y vssd1 vssd1 vccd1 vccd1 _2049_/Y sky130_fd_sc_hd__nand3_4
XFILLER_54_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2118_ _1589_/Y _1579_/X _1669_/B _1694_/X vssd1 vssd1 vccd1 vccd1 _2119_/A sky130_fd_sc_hd__and4_4
XFILLER_54_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1351_ _1351_/A _1351_/B _1361_/B vssd1 vssd1 vccd1 vccd1 _1351_/Y sky130_fd_sc_hd__nor3_4
X_1420_ _1420_/A vssd1 vssd1 vccd1 vccd1 _1420_/Y sky130_fd_sc_hd__inv_2
XFILLER_63_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1282_ _1281_/Y _2010_/B _1272_/Y vssd1 vssd1 vccd1 vccd1 _1282_/X sky130_fd_sc_hd__and3_4
XFILLER_0_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1618_ _2447_/Q vssd1 vssd1 vccd1 vccd1 _1618_/X sky130_fd_sc_hd__buf_2
XFILLER_39_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2598_ _2389_/CLK _2598_/D vssd1 vssd1 vccd1 vccd1 _1589_/A sky130_fd_sc_hd__dfxtp_4
X_1549_ _1541_/X vssd1 vssd1 vccd1 vccd1 _1549_/Y sky130_fd_sc_hd__inv_2
XFILLER_54_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_3_1_0_addressalyzerBlock.SPI_CLK clkbuf_3_1_0_addressalyzerBlock.SPI_CLK/A
+ vssd1 vssd1 vccd1 vccd1 clkbuf_4_3_0_addressalyzerBlock.SPI_CLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_49_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2521_ _2521_/CLK _1938_/Y vssd1 vssd1 vccd1 vccd1 _1952_/B sky130_fd_sc_hd__dfxtp_4
X_2383_ _2464_/CLK _2381_/Q vssd1 vssd1 vccd1 vccd1 _2384_/D sky130_fd_sc_hd__dfxtp_4
X_1403_ _1231_/B _1401_/Y _1402_/Y vssd1 vssd1 vccd1 vccd1 _1404_/A sky130_fd_sc_hd__o21ai_4
X_2452_ _2646_/CLK _2452_/D vssd1 vssd1 vccd1 vccd1 _2452_/Q sky130_fd_sc_hd__dfxtp_4
X_1334_ _2630_/Q vssd1 vssd1 vccd1 vccd1 _1335_/D sky130_fd_sc_hd__buf_2
X_1265_ _1265_/A _1300_/A vssd1 vssd1 vccd1 vccd1 _1265_/Y sky130_fd_sc_hd__nor2_4
X_1196_ _1862_/B _1188_/X _1191_/X vssd1 vssd1 vccd1 vccd1 _1196_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_24_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_2_0_0_m1_clk_local clkbuf_1_0_0_m1_clk_local/X vssd1 vssd1 vccd1 vccd1 clkbuf_3_1_0_m1_clk_local/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_42_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1883_ _1885_/A _1883_/B vssd1 vssd1 vccd1 vccd1 _1883_/X sky130_fd_sc_hd__and2_4
X_1952_ _1954_/A _1952_/B vssd1 vssd1 vccd1 vccd1 _1952_/X sky130_fd_sc_hd__and2_4
X_2435_ _2437_/CLK _2237_/Y vssd1 vssd1 vccd1 vccd1 _1218_/A sky130_fd_sc_hd__dfxtp_4
X_2504_ _2635_/CLK _2504_/D vssd1 vssd1 vccd1 vccd1 _1970_/B sky130_fd_sc_hd__dfxtp_4
X_2366_ _2492_/CLK _2366_/D vssd1 vssd1 vccd1 vccd1 _2367_/D sky130_fd_sc_hd__dfxtp_4
XFILLER_56_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1317_ _1856_/B _1316_/X _1306_/X vssd1 vssd1 vccd1 vccd1 _1317_/X sky130_fd_sc_hd__o21a_4
X_1248_ _1273_/A _2641_/Q vssd1 vssd1 vccd1 vccd1 _1249_/A sky130_fd_sc_hd__nand2_4
X_2297_ _2290_/Y vssd1 vssd1 vccd1 vccd1 _2304_/A sky130_fd_sc_hd__buf_2
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1179_ _1202_/B vssd1 vssd1 vccd1 vccd1 _1179_/X sky130_fd_sc_hd__buf_2
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2082_ _2081_/X _2057_/B _2072_/B vssd1 vssd1 vccd1 vccd1 _2474_/D sky130_fd_sc_hd__and3_4
XFILLER_38_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2220_ _1625_/X _1913_/A _2448_/Q vssd1 vssd1 vccd1 vccd1 _2220_/Y sky130_fd_sc_hd__a21oi_4
X_2151_ _2196_/A _2151_/B vssd1 vssd1 vccd1 vccd1 _2151_/Y sky130_fd_sc_hd__nand2_4
XFILLER_61_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1866_ _1972_/A _1972_/B vssd1 vssd1 vccd1 vccd1 _1973_/B sky130_fd_sc_hd__nand2_4
X_1935_ _1339_/X vssd1 vssd1 vccd1 vccd1 _1938_/A sky130_fd_sc_hd__buf_2
X_1797_ _1788_/X _1490_/A _2326_/A vssd1 vssd1 vccd1 vccd1 _1797_/X sky130_fd_sc_hd__o21a_4
X_2418_ _2418_/CLK _2281_/Y vssd1 vssd1 vccd1 vccd1 _1619_/A sky130_fd_sc_hd__dfxtp_4
X_2349_ _2349_/A MISO_fromClient vssd1 vssd1 vccd1 vccd1 _2349_/Y sky130_fd_sc_hd__nor2_4
XFILLER_29_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_4_3_0_m1_clk_local clkbuf_4_3_0_m1_clk_local/A vssd1 vssd1 vccd1 vccd1 _2632_/CLK
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_16_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1651_ _1605_/X vssd1 vssd1 vccd1 vccd1 _1856_/C sky130_fd_sc_hd__buf_2
X_1720_ _1718_/Y _1719_/X _1645_/A vssd1 vssd1 vccd1 vccd1 _1720_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_11_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1582_ _1581_/X _1562_/Y _1569_/X vssd1 vssd1 vccd1 vccd1 _1582_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_3_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2065_ _2055_/X _1993_/B _2064_/Y vssd1 vssd1 vccd1 vccd1 _2065_/X sky130_fd_sc_hd__o21a_4
X_2203_ _2181_/A _1764_/Y vssd1 vssd1 vccd1 vccd1 _2203_/Y sky130_fd_sc_hd__nor2_4
X_2134_ _2120_/A _2335_/A _2443_/Q vssd1 vssd1 vccd1 vccd1 _2134_/Y sky130_fd_sc_hd__nand3_4
XFILLER_1_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1849_ _1847_/Y _1624_/X _1848_/Y vssd1 vssd1 vccd1 vccd1 _1849_/Y sky130_fd_sc_hd__o21ai_4
X_1918_ _1918_/A _2540_/Q vssd1 vssd1 vccd1 vccd1 _1918_/X sky130_fd_sc_hd__and2_4
XFILLER_57_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1703_ _1634_/X vssd1 vssd1 vccd1 vccd1 _2224_/A sky130_fd_sc_hd__buf_2
X_1634_ _2447_/Q vssd1 vssd1 vccd1 vccd1 _1634_/X sky130_fd_sc_hd__buf_2
XPHY_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1565_ _2386_/Q vssd1 vssd1 vccd1 vccd1 _1731_/B sky130_fd_sc_hd__buf_2
X_1496_ _1487_/A _1494_/X _1495_/Y vssd1 vssd1 vccd1 vccd1 _1496_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_66_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2048_ _2014_/X _2040_/X _1986_/Y vssd1 vssd1 vccd1 vccd1 _2048_/Y sky130_fd_sc_hd__o21ai_4
X_2117_ _2117_/A vssd1 vssd1 vccd1 vccd1 _2447_/D sky130_fd_sc_hd__inv_2
XFILLER_57_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1350_ _1238_/Y vssd1 vssd1 vccd1 vccd1 _1361_/B sky130_fd_sc_hd__buf_2
X_1281_ _1256_/Y _1225_/X _1265_/A _1300_/A _1280_/Y vssd1 vssd1 vccd1 vccd1 _1281_/Y
+ sky130_fd_sc_hd__o41ai_4
XFILLER_63_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2597_ _2552_/CLK _1603_/Y vssd1 vssd1 vccd1 vccd1 _2597_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_8_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1617_ _2448_/Q vssd1 vssd1 vccd1 vccd1 _1704_/A sky130_fd_sc_hd__inv_2
XFILLER_54_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1548_ _1467_/A _1556_/B _1451_/X _1548_/D vssd1 vssd1 vccd1 vccd1 _1548_/Y sky130_fd_sc_hd__nor4_4
X_1479_ _1457_/B _1449_/B _1213_/X vssd1 vssd1 vccd1 vccd1 _1479_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_50_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1402_ _1401_/Y _1231_/B _1388_/A vssd1 vssd1 vccd1 vccd1 _1402_/Y sky130_fd_sc_hd__a21oi_4
X_2451_ _2588_/CLK _2113_/X vssd1 vssd1 vccd1 vccd1 _1783_/C sky130_fd_sc_hd__dfxtp_4
X_2520_ _2513_/CLK _1939_/Y vssd1 vssd1 vccd1 vccd1 _2520_/Q sky130_fd_sc_hd__dfxtp_4
X_2382_ _2492_/CLK _2382_/D vssd1 vssd1 vccd1 vccd1 _2382_/Q sky130_fd_sc_hd__dfxtp_4
X_1333_ _1333_/A _1351_/B _1240_/Y _1238_/Y vssd1 vssd1 vccd1 vccd1 _1333_/Y sky130_fd_sc_hd__nor4_4
XFILLER_39_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1264_ _1264_/A vssd1 vssd1 vccd1 vccd1 _1264_/Y sky130_fd_sc_hd__inv_2
X_1195_ _2650_/Q _1179_/X _1194_/X vssd1 vssd1 vccd1 vccd1 _1195_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_51_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2649_ _2454_/CLK _2649_/D vssd1 vssd1 vccd1 vccd1 _1194_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_27_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1882_ _1885_/A _2566_/Q vssd1 vssd1 vccd1 vccd1 _1882_/X sky130_fd_sc_hd__and2_4
X_1951_ _1954_/A _2522_/Q vssd1 vssd1 vccd1 vccd1 _2514_/D sky130_fd_sc_hd__and2_4
XFILLER_14_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2365_ _2492_/CLK _2364_/Q vssd1 vssd1 vccd1 vccd1 _2366_/D sky130_fd_sc_hd__dfxtp_4
X_2503_ _2635_/CLK _1967_/Y vssd1 vssd1 vccd1 vccd1 _1971_/B sky130_fd_sc_hd__dfxtp_4
X_2434_ _2604_/CLK _2434_/D vssd1 vssd1 vccd1 vccd1 _2434_/Q sky130_fd_sc_hd__dfxtp_4
X_1178_ _1833_/A vssd1 vssd1 vccd1 vccd1 _1202_/B sky130_fd_sc_hd__buf_2
X_1316_ _1239_/Y _1316_/B _1241_/Y _1316_/D vssd1 vssd1 vccd1 vccd1 _1316_/X sky130_fd_sc_hd__and4_4
X_1247_ _1225_/X _1226_/Y _1227_/Y _1246_/Y vssd1 vssd1 vccd1 vccd1 _1277_/B sky130_fd_sc_hd__nor4_4
X_2296_ _2266_/Y _2291_/X _2295_/Y vssd1 vssd1 vccd1 vccd1 _2296_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_64_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_4_11_0_m1_clk_local clkbuf_3_5_0_m1_clk_local/X vssd1 vssd1 vccd1 vccd1 _2470_/CLK
+ sky130_fd_sc_hd__clkbuf_1
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2081_ _2474_/Q _2080_/Y vssd1 vssd1 vccd1 vccd1 _2081_/X sky130_fd_sc_hd__or2_4
X_2150_ _1623_/Y vssd1 vssd1 vccd1 vccd1 _2196_/A sky130_fd_sc_hd__buf_2
X_1934_ _1933_/A _2527_/Q vssd1 vssd1 vccd1 vccd1 _1934_/X sky130_fd_sc_hd__and2_4
X_1865_ _2366_/D _2364_/Q _1865_/C vssd1 vssd1 vccd1 vccd1 _1869_/A sky130_fd_sc_hd__nor3_4
X_1796_ _1983_/B _2577_/Q _1795_/X vssd1 vssd1 vccd1 vccd1 _1796_/X sky130_fd_sc_hd__o21a_4
X_2348_ _2464_/Q vssd1 vssd1 vccd1 vccd1 _2348_/Y sky130_fd_sc_hd__inv_2
X_2417_ _2418_/CLK _2282_/Y vssd1 vssd1 vccd1 vccd1 _2417_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_44_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2279_ _1583_/X _1597_/X _1567_/B _1694_/X _1219_/X vssd1 vssd1 vccd1 vccd1 _2279_/X
+ sky130_fd_sc_hd__a41o_4
XFILLER_52_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1650_ _1649_/Y vssd1 vssd1 vccd1 vccd1 _1856_/A sky130_fd_sc_hd__buf_2
X_1581_ _1581_/A vssd1 vssd1 vccd1 vccd1 _1581_/X sky130_fd_sc_hd__buf_2
XFILLER_11_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2202_ _2198_/Y _2201_/Y _2449_/Q vssd1 vssd1 vccd1 vccd1 _2202_/X sky130_fd_sc_hd__a21o_4
XFILLER_21_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2064_ _2058_/X _2060_/Y _2062_/B _2055_/X _1275_/X vssd1 vssd1 vccd1 vccd1 _2064_/Y
+ sky130_fd_sc_hd__a41oi_4
X_2133_ _1886_/A _2121_/X _1490_/A vssd1 vssd1 vccd1 vccd1 _2133_/Y sky130_fd_sc_hd__nand3_4
XFILLER_19_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1917_ _1918_/A _1917_/B vssd1 vssd1 vccd1 vccd1 _1917_/X sky130_fd_sc_hd__and2_4
XFILLER_22_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1779_ _1779_/A _1678_/A _1783_/C vssd1 vssd1 vccd1 vccd1 _1779_/Y sky130_fd_sc_hd__nand3_4
X_1848_ _1625_/X _1902_/A _2448_/Q vssd1 vssd1 vccd1 vccd1 _1848_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_57_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_1_0_addressalyzerBlock.SPI_CLK clkbuf_3_0_0_addressalyzerBlock.SPI_CLK/X
+ vssd1 vssd1 vccd1 vccd1 _2404_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_16_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1564_ _1564_/A _1563_/Y vssd1 vssd1 vccd1 vccd1 _1564_/X sky130_fd_sc_hd__or2_4
X_1702_ _1702_/A vssd1 vssd1 vccd1 vccd1 _1702_/Y sky130_fd_sc_hd__inv_2
X_1633_ _1632_/Y vssd1 vssd1 vccd1 vccd1 _1633_/X sky130_fd_sc_hd__buf_2
XFILLER_66_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1495_ _1487_/A _1487_/B _1504_/A _1486_/X _2340_/C vssd1 vssd1 vccd1 vccd1 _1495_/Y
+ sky130_fd_sc_hd__a41oi_4
X_2047_ _2047_/A vssd1 vssd1 vccd1 vccd1 _2049_/A sky130_fd_sc_hd__inv_2
XFILLER_62_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2116_ _1545_/X _1576_/X _1588_/Y _1593_/Y _1595_/X vssd1 vssd1 vccd1 vccd1 _2448_/D
+ sky130_fd_sc_hd__a41oi_4
XFILLER_22_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_3_6_0_addressalyzerBlock.SPI_CLK clkbuf_3_6_0_addressalyzerBlock.SPI_CLK/A
+ vssd1 vssd1 vccd1 vccd1 clkbuf_3_6_0_addressalyzerBlock.SPI_CLK/X sky130_fd_sc_hd__clkbuf_1
XFILLER_9_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1280_ _2641_/Q vssd1 vssd1 vccd1 vccd1 _1280_/Y sky130_fd_sc_hd__inv_2
X_2596_ _2437_/CLK _2596_/D vssd1 vssd1 vccd1 vccd1 _1676_/B sky130_fd_sc_hd__dfxtp_4
X_1547_ _1577_/A _2390_/Q _1477_/A vssd1 vssd1 vccd1 vccd1 _1547_/X sky130_fd_sc_hd__o21a_4
X_1616_ _2447_/Q vssd1 vssd1 vccd1 vccd1 _2181_/A sky130_fd_sc_hd__buf_2
X_1478_ _1477_/X _2333_/B _1462_/X vssd1 vssd1 vccd1 vccd1 _1478_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_50_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2381_ _2508_/CLK _2381_/D vssd1 vssd1 vccd1 vccd1 _2381_/Q sky130_fd_sc_hd__dfxtp_4
X_1401_ _1363_/A _1363_/C vssd1 vssd1 vccd1 vccd1 _1401_/Y sky130_fd_sc_hd__nor2_4
X_2450_ _2588_/CLK _2114_/X vssd1 vssd1 vccd1 vccd1 _2450_/Q sky130_fd_sc_hd__dfxtp_4
X_1194_ _1194_/A _1194_/B vssd1 vssd1 vccd1 vccd1 _1194_/X sky130_fd_sc_hd__or2_4
X_1332_ _1332_/A vssd1 vssd1 vccd1 vccd1 _1333_/A sky130_fd_sc_hd__inv_2
X_1263_ _1263_/A _1289_/B _1263_/C vssd1 vssd1 vccd1 vccd1 _1264_/A sky130_fd_sc_hd__nand3_4
XFILLER_51_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2648_ _2454_/CLK _1205_/Y vssd1 vssd1 vccd1 vccd1 _1202_/A sky130_fd_sc_hd__dfxtp_4
X_2579_ _2399_/CLK _1812_/X vssd1 vssd1 vccd1 vccd1 _2579_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_42_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1950_ _1254_/X vssd1 vssd1 vccd1 vccd1 _1954_/A sky130_fd_sc_hd__buf_2
XFILLER_14_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1881_ _1885_/A DATA_FROM_HASH[0] vssd1 vssd1 vccd1 vccd1 _1881_/X sky130_fd_sc_hd__and2_4
X_2502_ _2505_/CLK _2502_/D vssd1 vssd1 vccd1 vccd1 MACRO_WR_SELECT[3] sky130_fd_sc_hd__dfxtp_4
X_2364_ _2492_/CLK _2364_/D vssd1 vssd1 vccd1 vccd1 _2364_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_51_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1315_ _1315_/A vssd1 vssd1 vccd1 vccd1 _1316_/B sky130_fd_sc_hd__buf_2
X_2433_ _2418_/CLK _2433_/D vssd1 vssd1 vccd1 vccd1 _2433_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_64_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1246_ _1239_/Y _1241_/Y _1243_/X _1305_/D vssd1 vssd1 vccd1 vccd1 _1246_/Y sky130_fd_sc_hd__nand4_4
X_2295_ _2292_/X _2300_/B _2295_/C vssd1 vssd1 vccd1 vccd1 _2295_/Y sky130_fd_sc_hd__nand3_4
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2080_ _2084_/C vssd1 vssd1 vccd1 vccd1 _2080_/Y sky130_fd_sc_hd__inv_2
XFILLER_34_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1933_ _1933_/A _2528_/Q vssd1 vssd1 vccd1 vccd1 _2524_/D sky130_fd_sc_hd__and2_4
X_1864_ _2367_/D vssd1 vssd1 vccd1 vccd1 _1865_/C sky130_fd_sc_hd__inv_2
X_1795_ _1788_/X _1477_/X _2326_/A vssd1 vssd1 vccd1 vccd1 _1795_/X sky130_fd_sc_hd__o21a_4
X_2347_ _1868_/A S1_CLK_SELECT _2346_/Y vssd1 vssd1 vccd1 vccd1 _2347_/X sky130_fd_sc_hd__o21a_4
XFILLER_29_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2278_ _2277_/Y vssd1 vssd1 vccd1 vccd1 _2278_/X sky130_fd_sc_hd__buf_2
X_2416_ _2404_/CLK _2416_/D vssd1 vssd1 vccd1 vccd1 _2416_/Q sky130_fd_sc_hd__dfxtp_4
X_1229_ _2619_/Q vssd1 vssd1 vccd1 vccd1 _1229_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1580_ _1579_/X vssd1 vssd1 vccd1 vccd1 _1581_/A sky130_fd_sc_hd__buf_2
XFILLER_7_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2132_ _2120_/X _2130_/Y _2131_/Y vssd1 vssd1 vccd1 vccd1 _2444_/D sky130_fd_sc_hd__o21ai_4
X_2201_ _2199_/Y _2201_/B _2201_/C vssd1 vssd1 vccd1 vccd1 _2201_/Y sky130_fd_sc_hd__nand3_4
X_2063_ _2063_/A _2063_/B _2063_/C vssd1 vssd1 vccd1 vccd1 _2063_/Y sky130_fd_sc_hd__nor3_4
X_1847_ _2424_/Q vssd1 vssd1 vccd1 vccd1 _1847_/Y sky130_fd_sc_hd__inv_2
X_1916_ _1918_/A _2542_/Q vssd1 vssd1 vccd1 vccd1 _2536_/D sky130_fd_sc_hd__and2_4
X_1778_ _1770_/Y _1777_/X _1439_/X vssd1 vssd1 vccd1 vccd1 _1779_/A sky130_fd_sc_hd__a21o_4
XFILLER_27_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1701_ _1701_/A _1701_/B vssd1 vssd1 vccd1 vccd1 _1702_/A sky130_fd_sc_hd__nand2_4
XPHY_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1563_ _1488_/A _1559_/Y _1562_/Y _2583_/Q _1527_/Y vssd1 vssd1 vccd1 vccd1 _1563_/Y
+ sky130_fd_sc_hd__a32oi_4
X_1632_ _2449_/Q vssd1 vssd1 vccd1 vccd1 _1632_/Y sky130_fd_sc_hd__inv_2
X_1494_ _1432_/X _1504_/A _1486_/X _1438_/D vssd1 vssd1 vccd1 vccd1 _1494_/X sky130_fd_sc_hd__and4_4
X_2115_ _1545_/X _1576_/X _1578_/Y _1582_/Y _1586_/X vssd1 vssd1 vccd1 vccd1 _2449_/D
+ sky130_fd_sc_hd__a41oi_4
X_2046_ _2019_/A _1997_/B _2045_/Y vssd1 vssd1 vccd1 vccd1 _2046_/Y sky130_fd_sc_hd__nor3_4
XFILLER_22_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_3_5_0_m1_clk_local clkbuf_3_5_0_m1_clk_local/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_5_0_m1_clk_local/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_5_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2595_ _2588_/CLK _2595_/D vssd1 vssd1 vccd1 vccd1 _1678_/A sky130_fd_sc_hd__dfxtp_4
X_1546_ _1544_/Y _1530_/A _1545_/X _1530_/C _1467_/Y vssd1 vssd1 vccd1 vccd1 _1546_/X
+ sky130_fd_sc_hd__a41o_4
X_1615_ _1534_/X _2558_/Q _1614_/X vssd1 vssd1 vccd1 vccd1 _1615_/Y sky130_fd_sc_hd__o21ai_4
X_1477_ _1477_/A vssd1 vssd1 vccd1 vccd1 _1477_/X sky130_fd_sc_hd__buf_2
XFILLER_54_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2029_ _2014_/X _2015_/C vssd1 vssd1 vccd1 vccd1 _2029_/Y sky130_fd_sc_hd__nor2_4
XFILLER_35_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2380_ _2508_/CLK _2379_/Q vssd1 vssd1 vccd1 vccd1 _2381_/D sky130_fd_sc_hd__dfxtp_4
X_1400_ _1399_/X vssd1 vssd1 vccd1 vccd1 _2618_/D sky130_fd_sc_hd__inv_2
X_1331_ _2632_/Q _1330_/X _1306_/X vssd1 vssd1 vccd1 vccd1 _1331_/X sky130_fd_sc_hd__o21a_4
XFILLER_5_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1193_ _1183_/Y _1187_/X _1192_/Y vssd1 vssd1 vccd1 vccd1 _1193_/Y sky130_fd_sc_hd__a21oi_4
X_1262_ _1251_/A _1261_/Y _1267_/A _1249_/Y vssd1 vssd1 vccd1 vccd1 _1263_/C sky130_fd_sc_hd__nand4_4
XFILLER_51_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2647_ _2454_/CLK _1209_/Y vssd1 vssd1 vccd1 vccd1 _2647_/Q sky130_fd_sc_hd__dfxtp_4
X_1529_ _1529_/A vssd1 vssd1 vccd1 vccd1 _1530_/C sky130_fd_sc_hd__inv_2
X_2578_ _2399_/CLK _1815_/X vssd1 vssd1 vccd1 vccd1 _2578_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_27_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1880_ _1886_/A vssd1 vssd1 vccd1 vccd1 _1885_/A sky130_fd_sc_hd__buf_2
XFILLER_14_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2501_ _2508_/CLK _2501_/D vssd1 vssd1 vccd1 vccd1 MACRO_WR_SELECT[2] sky130_fd_sc_hd__dfxtp_4
X_2363_ _2492_/CLK _2382_/Q vssd1 vssd1 vccd1 vccd1 _2364_/D sky130_fd_sc_hd__dfxtp_4
XFILLER_44_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1314_ _1314_/A vssd1 vssd1 vccd1 vccd1 _1314_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2294_ _1420_/Y _2291_/X _2293_/Y vssd1 vssd1 vccd1 vccd1 _2294_/Y sky130_fd_sc_hd__o21ai_4
X_2432_ _2404_/CLK _2432_/D vssd1 vssd1 vccd1 vccd1 _1902_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_64_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1245_ _1245_/A vssd1 vssd1 vccd1 vccd1 _1305_/D sky130_fd_sc_hd__inv_2
XFILLER_32_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1863_ _1861_/Y _1863_/B vssd1 vssd1 vccd1 vccd1 _1863_/Y sky130_fd_sc_hd__nand2_4
X_1932_ _1933_/A _2529_/Q vssd1 vssd1 vccd1 vccd1 _2525_/D sky130_fd_sc_hd__and2_4
XFILLER_21_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1794_ _1983_/B _2578_/Q _1793_/X vssd1 vssd1 vccd1 vccd1 _2586_/D sky130_fd_sc_hd__o21a_4
X_2415_ _2404_/CLK _2284_/Y vssd1 vssd1 vccd1 vccd1 _2415_/Q sky130_fd_sc_hd__dfxtp_4
X_2346_ _2345_/Y S1_CLK_SELECT vssd1 vssd1 vccd1 vccd1 _2346_/Y sky130_fd_sc_hd__nand2_4
X_1228_ _1367_/A _1360_/A vssd1 vssd1 vccd1 vccd1 _1351_/B sky130_fd_sc_hd__nand2_4
XFILLER_37_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2277_ _1590_/Y vssd1 vssd1 vccd1 vccd1 _2277_/Y sky130_fd_sc_hd__inv_2
XFILLER_52_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2062_ _2053_/Y _2062_/B _2055_/X _1993_/C vssd1 vssd1 vccd1 vccd1 _2063_/C sky130_fd_sc_hd__and4_4
X_2131_ _2120_/A _2335_/A _2131_/C vssd1 vssd1 vccd1 vccd1 _2131_/Y sky130_fd_sc_hd__nand3_4
X_2200_ _1946_/A _1634_/X vssd1 vssd1 vccd1 vccd1 _2201_/C sky130_fd_sc_hd__nand2_4
XFILLER_34_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_6_0_addressalyzerBlock.SPI_CLK clkbuf_4_7_0_addressalyzerBlock.SPI_CLK/A
+ vssd1 vssd1 vccd1 vccd1 _2552_/CLK sky130_fd_sc_hd__clkbuf_1
X_1915_ _1254_/X vssd1 vssd1 vccd1 vccd1 _1918_/A sky130_fd_sc_hd__buf_2
XFILLER_8_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1846_ ID_toHost _2181_/A _1704_/A _1845_/Y vssd1 vssd1 vccd1 vccd1 _1846_/X sky130_fd_sc_hd__a211o_4
X_1777_ _1777_/A _1774_/Y _1775_/Y _1776_/Y vssd1 vssd1 vccd1 vccd1 _1777_/X sky130_fd_sc_hd__and4_4
X_2329_ _2102_/A _2322_/A _1683_/Y _1574_/Y _2328_/X vssd1 vssd1 vccd1 vccd1 _2329_/Y
+ sky130_fd_sc_hd__o32ai_4
XFILLER_43_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1700_ _1645_/A _1308_/C _1612_/A vssd1 vssd1 vccd1 vccd1 _1700_/X sky130_fd_sc_hd__a21o_4
XPHY_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1631_ _1630_/X vssd1 vssd1 vccd1 vccd1 _1751_/A sky130_fd_sc_hd__buf_2
XPHY_260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1493_ _2092_/A _1492_/Y vssd1 vssd1 vccd1 vccd1 _1493_/Y sky130_fd_sc_hd__nor2_4
X_1562_ _1561_/Y vssd1 vssd1 vccd1 vccd1 _1562_/Y sky130_fd_sc_hd__inv_2
XFILLER_66_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2045_ _2029_/Y _2030_/X _2032_/C vssd1 vssd1 vccd1 vccd1 _2045_/Y sky130_fd_sc_hd__a21oi_4
X_2114_ _2104_/A ID_fromClient vssd1 vssd1 vccd1 vccd1 _2114_/X sky130_fd_sc_hd__and2_4
X_1829_ _1829_/A vssd1 vssd1 vccd1 vccd1 _1829_/Y sky130_fd_sc_hd__inv_2
XFILLER_57_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2594_ _2389_/CLK _2594_/D vssd1 vssd1 vccd1 vccd1 _2594_/Q sky130_fd_sc_hd__dfxtp_4
X_1614_ _1613_/Y vssd1 vssd1 vccd1 vccd1 _1614_/X sky130_fd_sc_hd__buf_2
XFILLER_8_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1545_ _1445_/Y vssd1 vssd1 vccd1 vccd1 _1545_/X sky130_fd_sc_hd__buf_2
XFILLER_5_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1476_ _1457_/B _1473_/X _1475_/Y vssd1 vssd1 vccd1 vccd1 _1476_/Y sky130_fd_sc_hd__o21ai_4
X_2028_ _2028_/A _2057_/B _2013_/D vssd1 vssd1 vccd1 vccd1 _2028_/X sky130_fd_sc_hd__and3_4
XFILLER_39_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1330_ _1318_/B _1335_/C _2630_/Q _1329_/X vssd1 vssd1 vccd1 vccd1 _1330_/X sky130_fd_sc_hd__and4_4
XFILLER_30_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1261_ _1256_/Y _1225_/X _1265_/A _1300_/A vssd1 vssd1 vccd1 vccd1 _1261_/Y sky130_fd_sc_hd__nor4_4
X_1192_ _1726_/B _1188_/X _1191_/X vssd1 vssd1 vccd1 vccd1 _1192_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_36_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2646_ _2646_/CLK _1215_/Y vssd1 vssd1 vccd1 vccd1 _1206_/A sky130_fd_sc_hd__dfxtp_4
X_2577_ _2399_/CLK _2577_/D vssd1 vssd1 vccd1 vccd1 _2577_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_55_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1528_ _1184_/A _1445_/A vssd1 vssd1 vccd1 vccd1 _1529_/A sky130_fd_sc_hd__nor2_4
X_1459_ _2127_/C vssd1 vssd1 vccd1 vccd1 _2266_/A sky130_fd_sc_hd__buf_2
XFILLER_42_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2500_ _2538_/CLK _2500_/D vssd1 vssd1 vccd1 vccd1 MACRO_WR_SELECT[1] sky130_fd_sc_hd__dfxtp_4
X_2431_ _2404_/CLK _2431_/D vssd1 vssd1 vccd1 vccd1 _2431_/Q sky130_fd_sc_hd__dfxtp_4
X_2362_ SCSN_fromHost vssd1 vssd1 vccd1 vccd1 SCSN_toClient sky130_fd_sc_hd__buf_2
X_1244_ _1856_/B _1315_/A vssd1 vssd1 vccd1 vccd1 _1245_/A sky130_fd_sc_hd__nand2_4
X_1313_ _1308_/C _1308_/A _1312_/Y vssd1 vssd1 vccd1 vccd1 _1314_/A sky130_fd_sc_hd__o21ai_4
XFILLER_37_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2293_ _2292_/X _2300_/B _2293_/C vssd1 vssd1 vccd1 vccd1 _2293_/Y sky130_fd_sc_hd__nand3_4
X_2629_ _2623_/CLK _1348_/Y vssd1 vssd1 vccd1 vccd1 _1332_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_43_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1862_ _2192_/A _1862_/B vssd1 vssd1 vccd1 vccd1 _1863_/B sky130_fd_sc_hd__nand2_4
X_1793_ _1788_/X _2266_/A _2326_/A vssd1 vssd1 vccd1 vccd1 _1793_/X sky130_fd_sc_hd__o21a_4
X_1931_ _1933_/A _2530_/Q vssd1 vssd1 vccd1 vccd1 _2526_/D sky130_fd_sc_hd__and2_4
X_2414_ _2418_/CLK _2414_/D vssd1 vssd1 vccd1 vccd1 _2151_/B sky130_fd_sc_hd__dfxtp_4
X_2345_ S1_CLK_IN vssd1 vssd1 vccd1 vccd1 _2345_/Y sky130_fd_sc_hd__inv_2
X_1227_ _1295_/A _1299_/A vssd1 vssd1 vccd1 vccd1 _1227_/Y sky130_fd_sc_hd__nand2_4
XFILLER_25_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2276_ _1581_/X vssd1 vssd1 vccd1 vccd1 _2276_/X sky130_fd_sc_hd__buf_2
XFILLER_52_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_4_11_0_addressalyzerBlock.SPI_CLK clkbuf_3_5_0_addressalyzerBlock.SPI_CLK/X
+ vssd1 vssd1 vccd1 vccd1 _2588_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_3_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2061_ _2058_/X _2060_/Y _2062_/B _2055_/X _1993_/C vssd1 vssd1 vccd1 vccd1 _2063_/B
+ sky130_fd_sc_hd__a41oi_4
X_2130_ _1840_/B _2121_/X _1477_/X vssd1 vssd1 vccd1 vccd1 _2130_/Y sky130_fd_sc_hd__nand3_4
X_1914_ _1928_/A _1913_/Y vssd1 vssd1 vccd1 vccd1 _2537_/D sky130_fd_sc_hd__nor2_4
X_1845_ _1618_/X _1845_/B vssd1 vssd1 vccd1 vccd1 _1845_/Y sky130_fd_sc_hd__nor2_4
X_1776_ _1512_/Y _1764_/A _1504_/A _1771_/Y vssd1 vssd1 vccd1 vccd1 _1776_/Y sky130_fd_sc_hd__a22oi_4
XFILLER_57_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2328_ _1187_/A _2462_/Q _1781_/A vssd1 vssd1 vccd1 vccd1 _2328_/X sky130_fd_sc_hd__a21o_4
XFILLER_57_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2259_ _2243_/Y _2257_/Y _2258_/X _1910_/Y _2248_/X vssd1 vssd1 vccd1 vccd1 _2259_/Y
+ sky130_fd_sc_hd__o32ai_4
XFILLER_43_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1630_ _2447_/Q vssd1 vssd1 vccd1 vccd1 _1630_/X sky130_fd_sc_hd__buf_2
XPHY_272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1561_ _1567_/B _1669_/B vssd1 vssd1 vccd1 vccd1 _1561_/Y sky130_fd_sc_hd__nand2_4
X_1492_ _2609_/Q _1489_/X _1491_/Y _1449_/B vssd1 vssd1 vccd1 vccd1 _1492_/Y sky130_fd_sc_hd__a22oi_4
XFILLER_66_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2044_ _2044_/A _2057_/B _2044_/C vssd1 vssd1 vccd1 vccd1 _2044_/X sky130_fd_sc_hd__and3_4
XFILLER_54_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2113_ _2104_/A _2450_/Q vssd1 vssd1 vccd1 vccd1 _2113_/X sky130_fd_sc_hd__and2_4
XFILLER_30_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1759_ _1656_/X _1397_/A _1673_/B vssd1 vssd1 vccd1 vccd1 _1759_/Y sky130_fd_sc_hd__a21oi_4
X_1828_ _1809_/A _2455_/Q _1827_/X vssd1 vssd1 vccd1 vccd1 _2572_/D sky130_fd_sc_hd__o21a_4
XFILLER_0_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2593_ _2437_/CLK _1727_/Y vssd1 vssd1 vccd1 vccd1 _1726_/B sky130_fd_sc_hd__dfxtp_4
X_1613_ _1590_/Y _1605_/X _1667_/C _1667_/D vssd1 vssd1 vccd1 vccd1 _1613_/Y sky130_fd_sc_hd__nand4_4
X_1544_ _1556_/B _1548_/D _1488_/A vssd1 vssd1 vccd1 vccd1 _1544_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_5_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1475_ _1457_/B _1440_/B _1470_/X _1438_/A _2340_/C vssd1 vssd1 vccd1 vccd1 _1475_/Y
+ sky130_fd_sc_hd__a41oi_4
XFILLER_54_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2027_ _1346_/A vssd1 vssd1 vccd1 vccd1 _2057_/B sky130_fd_sc_hd__buf_2
XFILLER_35_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1191_ _2096_/A vssd1 vssd1 vccd1 vccd1 _1191_/X sky130_fd_sc_hd__buf_2
XFILLER_39_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1260_ _1258_/Y _1243_/X _1305_/D _1295_/D vssd1 vssd1 vccd1 vccd1 _1300_/A sky130_fd_sc_hd__nand4_4
XFILLER_51_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_3_1_0_m1_clk_local clkbuf_3_1_0_m1_clk_local/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_3_0_m1_clk_local/A
+ sky130_fd_sc_hd__clkbuf_1
X_2645_ _2646_/CLK _1223_/Y vssd1 vssd1 vccd1 vccd1 _2645_/Q sky130_fd_sc_hd__dfxtp_4
X_1527_ _1527_/A vssd1 vssd1 vccd1 vccd1 _1527_/Y sky130_fd_sc_hd__inv_2
X_2576_ _2399_/CLK _2576_/D vssd1 vssd1 vccd1 vccd1 _2576_/Q sky130_fd_sc_hd__dfxtp_4
X_1389_ _1395_/B _1385_/D _2621_/Q vssd1 vssd1 vccd1 vccd1 _1389_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_27_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1458_ _1438_/B _1457_/X _1452_/Y vssd1 vssd1 vccd1 vccd1 _1458_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_50_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2361_ SCLK_fromHost vssd1 vssd1 vccd1 vccd1 SCLK_toClient sky130_fd_sc_hd__buf_2
X_2430_ _2404_/CLK _2254_/Y vssd1 vssd1 vccd1 vccd1 _2154_/B sky130_fd_sc_hd__dfxtp_4
X_1243_ _1243_/A vssd1 vssd1 vccd1 vccd1 _1243_/X sky130_fd_sc_hd__buf_2
X_1312_ _1308_/C _1318_/B _1316_/D _1305_/D _1274_/X vssd1 vssd1 vccd1 vccd1 _1312_/Y
+ sky130_fd_sc_hd__a41oi_4
X_2292_ _2290_/Y vssd1 vssd1 vccd1 vccd1 _2292_/X sky130_fd_sc_hd__buf_2
XFILLER_32_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2628_ _2623_/CLK _1355_/Y vssd1 vssd1 vccd1 vccd1 _2628_/Q sky130_fd_sc_hd__dfxtp_4
X_2559_ _2561_/CLK _1881_/X vssd1 vssd1 vccd1 vccd1 _2559_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_55_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1930_ _1928_/A _1929_/Y vssd1 vssd1 vccd1 vccd1 _2527_/D sky130_fd_sc_hd__nor2_4
XFILLER_14_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1861_ _1859_/Y _1861_/B _1860_/X vssd1 vssd1 vccd1 vccd1 _1861_/Y sky130_fd_sc_hd__nand3_4
X_1792_ _1983_/B _2579_/Q _1791_/X vssd1 vssd1 vccd1 vccd1 _1792_/X sky130_fd_sc_hd__o21a_4
X_2413_ _2418_/CLK _2413_/D vssd1 vssd1 vccd1 vccd1 _2174_/B sky130_fd_sc_hd__dfxtp_4
X_2344_ _2342_/Y M1_CLK_SELECT _2343_/Y vssd1 vssd1 vccd1 vccd1 m1_clk_local sky130_fd_sc_hd__a21oi_4
XFILLER_6_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1226_ _2636_/Q _2635_/Q vssd1 vssd1 vccd1 vccd1 _1226_/Y sky130_fd_sc_hd__nand2_4
X_2275_ _2144_/Y _1648_/Y _2270_/X _1948_/Y _2263_/X vssd1 vssd1 vccd1 vccd1 _2419_/D
+ sky130_fd_sc_hd__o32ai_4
XFILLER_16_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2060_ _1990_/Y _2072_/B vssd1 vssd1 vccd1 vccd1 _2060_/Y sky130_fd_sc_hd__nor2_4
XFILLER_34_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1913_ _1913_/A vssd1 vssd1 vccd1 vccd1 _1913_/Y sky130_fd_sc_hd__inv_2
XFILLER_22_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1844_ _2416_/Q vssd1 vssd1 vccd1 vccd1 _1845_/B sky130_fd_sc_hd__inv_2
X_1775_ _1499_/Y _2398_/Q _1457_/B _1766_/B vssd1 vssd1 vccd1 vccd1 _1775_/Y sky130_fd_sc_hd__a22oi_4
X_2327_ _1222_/A _1218_/B _2462_/Q _1683_/Y _2326_/Y vssd1 vssd1 vccd1 vccd1 _2327_/Y
+ sky130_fd_sc_hd__o41ai_4
XFILLER_27_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2258_ _2246_/Y vssd1 vssd1 vccd1 vccd1 _2258_/X sky130_fd_sc_hd__buf_2
X_1209_ _1207_/Y _1187_/X _1208_/Y vssd1 vssd1 vccd1 vccd1 _1209_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_43_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2189_ _1666_/A THREAD_COUNT[2] vssd1 vssd1 vccd1 vccd1 _2189_/Y sky130_fd_sc_hd__nand2_4
XFILLER_48_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1560_ _1567_/C vssd1 vssd1 vccd1 vccd1 _1669_/B sky130_fd_sc_hd__buf_2
X_2112_ _2112_/A _2103_/Y vssd1 vssd1 vccd1 vccd1 _2452_/D sky130_fd_sc_hd__nand2_4
X_1491_ _2609_/Q _1451_/X _1487_/Y _1490_/Y _1445_/D vssd1 vssd1 vccd1 vccd1 _1491_/Y
+ sky130_fd_sc_hd__o32ai_4
XFILLER_66_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2043_ _2030_/X _2029_/Y _2032_/C _2043_/D vssd1 vssd1 vccd1 vccd1 _2044_/C sky130_fd_sc_hd__nand4_4
X_1827_ _2572_/Q _2461_/Q _2257_/A vssd1 vssd1 vccd1 vccd1 _1827_/X sky130_fd_sc_hd__o21a_4
X_1689_ _2391_/Q vssd1 vssd1 vccd1 vccd1 _1689_/Y sky130_fd_sc_hd__inv_2
X_1758_ _1742_/Y _1756_/Y _1757_/Y vssd1 vssd1 vccd1 vccd1 _1758_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_1_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_2_2_0_addressalyzerBlock.SPI_CLK clkbuf_2_3_0_addressalyzerBlock.SPI_CLK/A
+ vssd1 vssd1 vccd1 vccd1 clkbuf_3_5_0_addressalyzerBlock.SPI_CLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_54_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1612_ _1612_/A vssd1 vssd1 vccd1 vccd1 _1612_/X sky130_fd_sc_hd__buf_2
X_2592_ _2437_/CLK _2592_/D vssd1 vssd1 vccd1 vccd1 _2236_/A sky130_fd_sc_hd__dfxtp_4
X_1474_ _1451_/X vssd1 vssd1 vccd1 vccd1 _2340_/C sky130_fd_sc_hd__buf_2
X_1543_ _1539_/Y _1540_/Y _1542_/X vssd1 vssd1 vccd1 vccd1 _2603_/D sky130_fd_sc_hd__a21oi_4
XFILLER_8_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2026_ _2047_/A _2016_/X _1997_/A _1997_/D _2488_/Q vssd1 vssd1 vccd1 vccd1 _2028_/A
+ sky130_fd_sc_hd__a41o_4
XFILLER_50_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1190_ _1190_/A vssd1 vssd1 vccd1 vccd1 _2096_/A sky130_fd_sc_hd__buf_2
XFILLER_36_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2644_ _2632_/CLK _1264_/Y vssd1 vssd1 vccd1 vccd1 _1251_/A sky130_fd_sc_hd__dfxtp_4
X_1526_ _1577_/A _2390_/Q vssd1 vssd1 vccd1 vccd1 _1527_/A sky130_fd_sc_hd__nor2_4
X_2575_ _2611_/CLK _2575_/D vssd1 vssd1 vccd1 vccd1 _2575_/Q sky130_fd_sc_hd__dfxtp_4
X_1457_ _1440_/B _1457_/B _1438_/D _1438_/A vssd1 vssd1 vccd1 vccd1 _1457_/X sky130_fd_sc_hd__and4_4
X_1388_ _1388_/A vssd1 vssd1 vccd1 vccd1 _2019_/A sky130_fd_sc_hd__buf_2
XFILLER_35_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2009_ _2008_/Y _1984_/A _1999_/A _2011_/A _2492_/Q vssd1 vssd1 vccd1 vccd1 _2009_/X
+ sky130_fd_sc_hd__a41o_4
XFILLER_35_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1311_ _1243_/X vssd1 vssd1 vccd1 vccd1 _1316_/D sky130_fd_sc_hd__buf_2
X_2360_ MOSI_fromHost vssd1 vssd1 vccd1 vccd1 MOSI_toClient sky130_fd_sc_hd__buf_2
X_2291_ _2290_/Y vssd1 vssd1 vccd1 vccd1 _2291_/X sky130_fd_sc_hd__buf_2
XFILLER_49_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1242_ _2632_/Q _2631_/Q _2630_/Q _1332_/A vssd1 vssd1 vccd1 vccd1 _1243_/A sky130_fd_sc_hd__and4_4
XFILLER_2_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2627_ _2623_/CLK _1359_/Y vssd1 vssd1 vccd1 vccd1 _1349_/A sky130_fd_sc_hd__dfxtp_4
X_2489_ _2470_/CLK _2025_/Y vssd1 vssd1 vccd1 vccd1 _1984_/A sky130_fd_sc_hd__dfxtp_4
X_2558_ _2555_/CLK _1882_/X vssd1 vssd1 vccd1 vccd1 _2558_/Q sky130_fd_sc_hd__dfxtp_4
X_1509_ _1508_/X _1448_/A _1504_/Y vssd1 vssd1 vccd1 vccd1 _1509_/X sky130_fd_sc_hd__a21o_4
XFILLER_55_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1860_ _1231_/A _1661_/B _1661_/C _1661_/D vssd1 vssd1 vccd1 vccd1 _1860_/X sky130_fd_sc_hd__or4_4
XFILLER_6_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1791_ _1788_/X _1420_/A _2326_/A vssd1 vssd1 vccd1 vccd1 _1791_/X sky130_fd_sc_hd__o21a_4
X_2412_ _2418_/CLK _2412_/D vssd1 vssd1 vccd1 vccd1 _2196_/B sky130_fd_sc_hd__dfxtp_4
X_2343_ PLL_INPUT M1_CLK_SELECT vssd1 vssd1 vccd1 vccd1 _2343_/Y sky130_fd_sc_hd__nor2_4
X_2274_ _2142_/Y _1648_/Y _2270_/X _1946_/Y _2263_/X vssd1 vssd1 vccd1 vccd1 _2274_/Y
+ sky130_fd_sc_hd__o32ai_4
XFILLER_37_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1225_ _1225_/A vssd1 vssd1 vccd1 vccd1 _1225_/X sky130_fd_sc_hd__buf_2
XFILLER_60_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1989_ _2054_/A vssd1 vssd1 vccd1 vccd1 _1992_/B sky130_fd_sc_hd__inv_2
XFILLER_20_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1843_ _1534_/X _2556_/Q _1614_/X vssd1 vssd1 vccd1 vccd1 _1843_/Y sky130_fd_sc_hd__o21ai_4
X_1912_ _1339_/X vssd1 vssd1 vccd1 vccd1 _1928_/A sky130_fd_sc_hd__buf_2
XFILLER_8_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1774_ _1750_/Y _2609_/Q _1487_/A _2158_/B vssd1 vssd1 vccd1 vccd1 _1774_/Y sky130_fd_sc_hd__a22oi_4
X_1208_ _2192_/B _1187_/A _1191_/X vssd1 vssd1 vccd1 vccd1 _1208_/Y sky130_fd_sc_hd__o21ai_4
X_2326_ _2326_/A _2326_/B _1185_/A _2335_/D vssd1 vssd1 vccd1 vccd1 _2326_/Y sky130_fd_sc_hd__nand4_4
X_2257_ _2257_/A _1698_/A _1514_/X vssd1 vssd1 vccd1 vccd1 _2257_/Y sky130_fd_sc_hd__nand3_4
XFILLER_65_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2188_ _2185_/Y _2186_/X _2187_/X vssd1 vssd1 vccd1 vccd1 _2188_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_25_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1490_ _1490_/A vssd1 vssd1 vccd1 vccd1 _1490_/Y sky130_fd_sc_hd__inv_2
XFILLER_66_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2042_ _2041_/Y _1985_/A _2030_/X _2016_/X _2043_/D vssd1 vssd1 vccd1 vccd1 _2044_/A
+ sky130_fd_sc_hd__a41o_4
X_2111_ _2112_/A _2098_/Y vssd1 vssd1 vccd1 vccd1 _2111_/Y sky130_fd_sc_hd__nand2_4
XFILLER_62_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1826_ _2572_/Q _1809_/A _1825_/X vssd1 vssd1 vccd1 vccd1 _2573_/D sky130_fd_sc_hd__o21a_4
X_1757_ _1612_/A _1360_/A _1656_/A vssd1 vssd1 vccd1 vccd1 _1757_/Y sky130_fd_sc_hd__a21oi_4
X_1688_ _1731_/B _1566_/X _1687_/Y vssd1 vssd1 vccd1 vccd1 _1688_/Y sky130_fd_sc_hd__nor3_4
XFILLER_57_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2309_ _2144_/Y _2292_/X _2308_/Y vssd1 vssd1 vccd1 vccd1 _2403_/D sky130_fd_sc_hd__o21ai_4
XFILLER_48_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1611_ _1741_/A vssd1 vssd1 vccd1 vccd1 _1612_/A sky130_fd_sc_hd__buf_2
XFILLER_8_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1542_ _1541_/X _1469_/A _1500_/X vssd1 vssd1 vccd1 vccd1 _1542_/X sky130_fd_sc_hd__a21o_4
X_2591_ _2611_/CLK _2591_/D vssd1 vssd1 vccd1 vccd1 _2591_/Q sky130_fd_sc_hd__dfxtp_4
X_1473_ _1469_/Y _1470_/X _1473_/C _1438_/A vssd1 vssd1 vccd1 vccd1 _1473_/X sky130_fd_sc_hd__and4_4
X_2025_ _2002_/X _2013_/D _2024_/Y vssd1 vssd1 vccd1 vccd1 _2025_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_54_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1809_ _1809_/A vssd1 vssd1 vccd1 vccd1 _1809_/X sky130_fd_sc_hd__buf_2
XFILLER_53_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2643_ _2632_/CLK _1271_/X vssd1 vssd1 vccd1 vccd1 _1267_/A sky130_fd_sc_hd__dfxtp_4
X_2574_ _2611_/CLK _2574_/D vssd1 vssd1 vccd1 vccd1 _2574_/Q sky130_fd_sc_hd__dfxtp_4
X_1387_ _1386_/Y vssd1 vssd1 vccd1 vccd1 _2622_/D sky130_fd_sc_hd__inv_2
X_1456_ _1438_/C vssd1 vssd1 vccd1 vccd1 _1457_/B sky130_fd_sc_hd__buf_2
X_1525_ _1473_/C _1469_/Y _1524_/Y vssd1 vssd1 vccd1 vccd1 _1525_/Y sky130_fd_sc_hd__o21ai_4
X_2008_ _2008_/A vssd1 vssd1 vccd1 vccd1 _2008_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1241_ _1240_/Y vssd1 vssd1 vccd1 vccd1 _1241_/Y sky130_fd_sc_hd__inv_2
X_1310_ _1309_/Y vssd1 vssd1 vccd1 vccd1 _2636_/D sky130_fd_sc_hd__inv_2
X_2290_ _2289_/Y vssd1 vssd1 vccd1 vccd1 _2290_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2626_ _2623_/CLK _1369_/Y vssd1 vssd1 vccd1 vccd1 _1367_/A sky130_fd_sc_hd__dfxtp_4
X_2557_ _2561_/CLK _1883_/X vssd1 vssd1 vccd1 vccd1 _1701_/B sky130_fd_sc_hd__dfxtp_4
X_2488_ _2470_/CLK _2028_/X vssd1 vssd1 vccd1 vccd1 _2488_/Q sky130_fd_sc_hd__dfxtp_4
X_1439_ _1438_/X vssd1 vssd1 vccd1 vccd1 _1439_/X sky130_fd_sc_hd__buf_2
X_1508_ _1469_/Y _1486_/X _1438_/D _1473_/C _1451_/X vssd1 vssd1 vccd1 vccd1 _1508_/X
+ sky130_fd_sc_hd__a41o_4
XFILLER_62_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1790_ _1789_/X vssd1 vssd1 vccd1 vccd1 _2326_/A sky130_fd_sc_hd__buf_2
X_2411_ _2418_/CLK _2411_/D vssd1 vssd1 vccd1 vccd1 _2411_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_10_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1224_ _1224_/A vssd1 vssd1 vccd1 vccd1 _1225_/A sky130_fd_sc_hd__inv_2
X_2342_ M1_CLK_IN vssd1 vssd1 vccd1 vccd1 _2342_/Y sky130_fd_sc_hd__inv_2
X_2273_ _1503_/Y _1648_/Y _2270_/X _1944_/Y _2263_/X vssd1 vssd1 vccd1 vccd1 _2273_/Y
+ sky130_fd_sc_hd__o32ai_4
X_1988_ _2477_/Q vssd1 vssd1 vccd1 vccd1 _1992_/A sky130_fd_sc_hd__inv_2
Xclkbuf_2_3_0_m1_clk_local clkbuf_2_3_0_m1_clk_local/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_7_0_m1_clk_local/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_57_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2609_ _2588_/CLK _1493_/Y vssd1 vssd1 vccd1 vccd1 _2609_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_16_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_3_2_0_addressalyzerBlock.SPI_CLK clkbuf_3_3_0_addressalyzerBlock.SPI_CLK/A
+ vssd1 vssd1 vccd1 vccd1 clkbuf_3_2_0_addressalyzerBlock.SPI_CLK/X sky130_fd_sc_hd__clkbuf_1
XFILLER_19_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1842_ _1179_/X _1830_/C _1841_/Y vssd1 vssd1 vccd1 vccd1 _2569_/D sky130_fd_sc_hd__o21a_4
XFILLER_8_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1773_ _2398_/Q vssd1 vssd1 vccd1 vccd1 _2158_/B sky130_fd_sc_hd__inv_2
X_1911_ _1911_/A _1910_/Y vssd1 vssd1 vccd1 vccd1 _1911_/Y sky130_fd_sc_hd__nor2_4
X_1207_ _2647_/Q _1202_/B _1206_/X vssd1 vssd1 vccd1 vccd1 _1207_/Y sky130_fd_sc_hd__o21ai_4
X_2325_ _2324_/X _1688_/Y _2112_/A vssd1 vssd1 vccd1 vccd1 _2325_/X sky130_fd_sc_hd__o21a_4
X_2187_ _1741_/A _1376_/C _1656_/A vssd1 vssd1 vccd1 vccd1 _2187_/X sky130_fd_sc_hd__a21o_4
XFILLER_25_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2256_ _2244_/X _2255_/Y _2247_/X _1908_/Y _2249_/X vssd1 vssd1 vccd1 vccd1 _2256_/Y
+ sky130_fd_sc_hd__o32ai_4
XFILLER_4_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2041_ _2040_/X vssd1 vssd1 vccd1 vccd1 _2041_/Y sky130_fd_sc_hd__inv_2
X_2110_ _2107_/A MOSI_fromHost vssd1 vssd1 vccd1 vccd1 _2454_/D sky130_fd_sc_hd__and2_4
XFILLER_39_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1756_ _1753_/X _1754_/X _1755_/Y vssd1 vssd1 vccd1 vccd1 _1756_/Y sky130_fd_sc_hd__a21oi_4
X_1825_ _2573_/Q _2461_/Q _2257_/A vssd1 vssd1 vccd1 vccd1 _1825_/X sky130_fd_sc_hd__o21a_4
X_1687_ _1687_/A vssd1 vssd1 vccd1 vccd1 _1687_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_4_6_0_m1_clk_local clkbuf_3_3_0_m1_clk_local/X vssd1 vssd1 vccd1 vccd1 _2513_/CLK
+ sky130_fd_sc_hd__clkbuf_1
X_2308_ _2290_/Y _1602_/C _2089_/A vssd1 vssd1 vccd1 vccd1 _2308_/Y sky130_fd_sc_hd__nand3_4
XFILLER_38_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2239_ _2239_/A vssd1 vssd1 vccd1 vccd1 _2241_/A sky130_fd_sc_hd__inv_2
XFILLER_13_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2590_ _2437_/CLK _1763_/Y vssd1 vssd1 vccd1 vccd1 _1762_/B sky130_fd_sc_hd__dfxtp_4
X_1610_ _1609_/X vssd1 vssd1 vccd1 vccd1 _1741_/A sky130_fd_sc_hd__buf_2
XFILLER_8_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1541_ _1564_/A vssd1 vssd1 vccd1 vccd1 _1541_/X sky130_fd_sc_hd__buf_2
X_1472_ _1472_/A vssd1 vssd1 vccd1 vccd1 _1473_/C sky130_fd_sc_hd__buf_2
X_2024_ _2002_/X _2013_/D _1346_/X vssd1 vssd1 vccd1 vccd1 _2024_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_35_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1739_ _1761_/A _1739_/B vssd1 vssd1 vccd1 vccd1 _1739_/Y sky130_fd_sc_hd__nor2_4
XFILLER_49_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1808_ _2461_/Q vssd1 vssd1 vccd1 vccd1 _1809_/A sky130_fd_sc_hd__inv_2
XFILLER_65_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2642_ _2632_/CLK _2642_/D vssd1 vssd1 vccd1 vccd1 _1273_/A sky130_fd_sc_hd__dfxtp_4
X_2573_ _2611_/CLK _2573_/D vssd1 vssd1 vccd1 vccd1 _2573_/Q sky130_fd_sc_hd__dfxtp_4
X_1524_ _1473_/C _1432_/A _1466_/A _1467_/A _2340_/C vssd1 vssd1 vccd1 vccd1 _1524_/Y
+ sky130_fd_sc_hd__a41oi_4
X_1386_ _1384_/X _1385_/Y vssd1 vssd1 vccd1 vccd1 _1386_/Y sky130_fd_sc_hd__nand2_4
X_1455_ _1449_/Y _1453_/Y _1454_/X vssd1 vssd1 vccd1 vccd1 _1455_/Y sky130_fd_sc_hd__a21oi_4
X_2007_ _2006_/Y vssd1 vssd1 vccd1 vccd1 _2493_/D sky130_fd_sc_hd__inv_2
XFILLER_35_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1240_ _2628_/Q _1349_/A vssd1 vssd1 vccd1 vccd1 _1240_/Y sky130_fd_sc_hd__nand2_4
XFILLER_64_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2487_ _2470_/CLK _2487_/D vssd1 vssd1 vccd1 vccd1 _1997_/A sky130_fd_sc_hd__dfxtp_4
X_2625_ _2623_/CLK _1371_/Y vssd1 vssd1 vccd1 vccd1 _1360_/A sky130_fd_sc_hd__dfxtp_4
X_2556_ _2555_/CLK _1884_/X vssd1 vssd1 vccd1 vccd1 _2556_/Q sky130_fd_sc_hd__dfxtp_4
X_1507_ _1506_/Y _1449_/B vssd1 vssd1 vccd1 vccd1 _1507_/Y sky130_fd_sc_hd__nand2_4
X_1369_ _1369_/A vssd1 vssd1 vccd1 vccd1 _1369_/Y sky130_fd_sc_hd__inv_2
X_1438_ _1438_/A _1438_/B _1438_/C _1438_/D vssd1 vssd1 vccd1 vccd1 _1438_/X sky130_fd_sc_hd__and4_4
XFILLER_62_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2341_ EXT_RESET_N_fromHost vssd1 vssd1 vccd1 vccd1 _2382_/D sky130_fd_sc_hd__inv_2
X_2410_ _2604_/CLK _2294_/Y vssd1 vssd1 vccd1 vccd1 _2293_/C sky130_fd_sc_hd__dfxtp_4
X_1223_ _1216_/Y _1218_/Y _2092_/A vssd1 vssd1 vccd1 vccd1 _1223_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_28_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2272_ _2136_/Y _2262_/X _2270_/X _1942_/B _2264_/X vssd1 vssd1 vccd1 vccd1 _2422_/D
+ sky130_fd_sc_hd__o32ai_4
XFILLER_52_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1987_ _1987_/A vssd1 vssd1 vccd1 vccd1 _1994_/C sky130_fd_sc_hd__inv_2
XFILLER_9_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2539_ _2519_/CLK _2539_/D vssd1 vssd1 vccd1 vccd1 _1919_/B sky130_fd_sc_hd__dfxtp_4
X_2608_ _2611_/CLK _1502_/Y vssd1 vssd1 vccd1 vccd1 _1436_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_43_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1910_ _2428_/Q vssd1 vssd1 vccd1 vccd1 _1910_/Y sky130_fd_sc_hd__inv_2
XFILLER_19_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1841_ _1840_/Y vssd1 vssd1 vccd1 vccd1 _1841_/Y sky130_fd_sc_hd__inv_2
XFILLER_8_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1772_ _2609_/Q _1750_/Y _2607_/Q _1771_/Y vssd1 vssd1 vccd1 vccd1 _1777_/A sky130_fd_sc_hd__o22a_4
X_2324_ _1731_/B _1566_/X _2391_/Q vssd1 vssd1 vccd1 vccd1 _2324_/X sky130_fd_sc_hd__o21a_4
Xclkbuf_4_14_0_m1_clk_local clkbuf_3_7_0_m1_clk_local/X vssd1 vssd1 vccd1 vccd1 _2374_/CLK
+ sky130_fd_sc_hd__clkbuf_1
X_1206_ _1206_/A _1198_/B vssd1 vssd1 vccd1 vccd1 _1206_/X sky130_fd_sc_hd__or2_4
X_2186_ _1335_/C _1645_/Y _1741_/Y vssd1 vssd1 vccd1 vccd1 _2186_/X sky130_fd_sc_hd__o21a_4
X_2255_ _2257_/A _1698_/A _1503_/A vssd1 vssd1 vccd1 vccd1 _2255_/Y sky130_fd_sc_hd__nand3_4
XFILLER_56_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2040_ _2015_/C vssd1 vssd1 vccd1 vccd1 _2040_/X sky130_fd_sc_hd__buf_2
XFILLER_47_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1686_ _1678_/Y _1682_/Y _1685_/X vssd1 vssd1 vccd1 vccd1 _2595_/D sky130_fd_sc_hd__a21oi_4
X_1755_ _1280_/Y _1614_/X _1646_/X vssd1 vssd1 vccd1 vccd1 _1755_/Y sky130_fd_sc_hd__o21ai_4
X_1824_ _1789_/X vssd1 vssd1 vccd1 vccd1 _2257_/A sky130_fd_sc_hd__buf_2
XFILLER_57_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2238_ _1606_/Y _1190_/A _1583_/X _1696_/A vssd1 vssd1 vccd1 vccd1 _2239_/A sky130_fd_sc_hd__and4_4
X_2307_ _2142_/Y _2292_/X _2306_/Y vssd1 vssd1 vccd1 vccd1 _2404_/D sky130_fd_sc_hd__o21ai_4
XFILLER_65_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2169_ _2546_/Q _1739_/B _2167_/Y _2168_/Y vssd1 vssd1 vccd1 vccd1 _2169_/Y sky130_fd_sc_hd__a22oi_4
XFILLER_13_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1540_ _2266_/A _1527_/Y _1556_/A vssd1 vssd1 vccd1 vccd1 _1540_/Y sky130_fd_sc_hd__a21oi_4
X_1471_ _2604_/Q vssd1 vssd1 vccd1 vccd1 _1472_/A sky130_fd_sc_hd__buf_2
X_2023_ _2022_/Y vssd1 vssd1 vccd1 vccd1 _2490_/D sky130_fd_sc_hd__inv_2
XFILLER_62_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1807_ _1786_/Y _2572_/Q _1806_/X vssd1 vssd1 vccd1 vccd1 _1807_/X sky130_fd_sc_hd__o21a_4
X_1738_ _1831_/A _1738_/B vssd1 vssd1 vccd1 vccd1 _2591_/D sky130_fd_sc_hd__nor2_4
X_1669_ _1579_/X _1669_/B _1589_/Y vssd1 vssd1 vccd1 vccd1 _1669_/Y sky130_fd_sc_hd__nor3_4
XFILLER_65_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1454_ _1222_/A vssd1 vssd1 vccd1 vccd1 _1454_/X sky130_fd_sc_hd__buf_2
X_2641_ _2632_/CLK _1282_/X vssd1 vssd1 vccd1 vccd1 _2641_/Q sky130_fd_sc_hd__dfxtp_4
X_2572_ _2611_/CLK _2572_/D vssd1 vssd1 vccd1 vccd1 _2572_/Q sky130_fd_sc_hd__dfxtp_4
X_1523_ _1519_/Y _1521_/Y _1522_/Y vssd1 vssd1 vccd1 vccd1 _1523_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_55_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1385_ _2622_/Q _1385_/B _2621_/Q _1385_/D vssd1 vssd1 vccd1 vccd1 _1385_/Y sky130_fd_sc_hd__nand4_4
XFILLER_27_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2006_ _2001_/Y _2022_/B _2006_/C vssd1 vssd1 vccd1 vccd1 _2006_/Y sky130_fd_sc_hd__nand3_4
XFILLER_50_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2624_ _2623_/CLK _1378_/Y vssd1 vssd1 vccd1 vccd1 _1376_/B sky130_fd_sc_hd__dfxtp_4
X_2486_ _2511_/CLK _2039_/Y vssd1 vssd1 vccd1 vccd1 _1995_/B sky130_fd_sc_hd__dfxtp_4
X_2555_ _2555_/CLK _2555_/D vssd1 vssd1 vccd1 vccd1 _2555_/Q sky130_fd_sc_hd__dfxtp_4
X_1506_ _1503_/Y _1445_/D _1505_/Y vssd1 vssd1 vccd1 vccd1 _1506_/Y sky130_fd_sc_hd__o21ai_4
Xclkbuf_4_2_0_addressalyzerBlock.SPI_CLK clkbuf_4_3_0_addressalyzerBlock.SPI_CLK/A
+ vssd1 vssd1 vccd1 vccd1 _2446_/CLK sky130_fd_sc_hd__clkbuf_1
X_1437_ _1483_/B vssd1 vssd1 vccd1 vccd1 _1438_/D sky130_fd_sc_hd__buf_2
X_1368_ _1362_/X _1367_/Y vssd1 vssd1 vccd1 vccd1 _1369_/A sky130_fd_sc_hd__nand2_4
X_1299_ _1299_/A vssd1 vssd1 vccd1 vccd1 _1299_/Y sky130_fd_sc_hd__inv_2
XFILLER_23_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_3_7_0_addressalyzerBlock.SPI_CLK clkbuf_3_6_0_addressalyzerBlock.SPI_CLK/A
+ vssd1 vssd1 vccd1 vccd1 clkbuf_3_7_0_addressalyzerBlock.SPI_CLK/X sky130_fd_sc_hd__clkbuf_1
XFILLER_6_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2340_ _2102_/A _1687_/Y _2340_/C vssd1 vssd1 vccd1 vccd1 _2393_/D sky130_fd_sc_hd__nor3_4
X_2271_ _1490_/Y _2262_/X _2270_/X _1746_/Y _2264_/X vssd1 vssd1 vccd1 vccd1 _2423_/D
+ sky130_fd_sc_hd__o32ai_4
X_1222_ _1222_/A vssd1 vssd1 vccd1 vccd1 _2092_/A sky130_fd_sc_hd__buf_2
X_1986_ _2483_/Q vssd1 vssd1 vccd1 vccd1 _1986_/Y sky130_fd_sc_hd__inv_2
XFILLER_52_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2607_ _2588_/CLK _1510_/Y vssd1 vssd1 vccd1 vccd1 _2607_/Q sky130_fd_sc_hd__dfxtp_4
X_2538_ _2538_/CLK _1911_/Y vssd1 vssd1 vccd1 vccd1 _2538_/Q sky130_fd_sc_hd__dfxtp_4
X_2469_ _2635_/CLK _2090_/Y vssd1 vssd1 vccd1 vccd1 _2469_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1840_ _1833_/Y _1840_/B _1840_/C vssd1 vssd1 vccd1 vccd1 _1840_/Y sky130_fd_sc_hd__nand3_4
XFILLER_42_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1771_ _2397_/Q vssd1 vssd1 vccd1 vccd1 _1771_/Y sky130_fd_sc_hd__inv_2
X_2323_ _2322_/Y _1697_/Y _2100_/A vssd1 vssd1 vccd1 vccd1 _2392_/D sky130_fd_sc_hd__a21oi_4
XFILLER_40_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2254_ _2244_/X _2253_/Y _2247_/X _1906_/Y _2249_/X vssd1 vssd1 vccd1 vccd1 _2254_/Y
+ sky130_fd_sc_hd__o32ai_4
X_1205_ _1203_/Y _1187_/X _1204_/Y vssd1 vssd1 vccd1 vccd1 _1205_/Y sky130_fd_sc_hd__a21oi_4
X_2185_ _2173_/Y _2183_/Y _2184_/Y vssd1 vssd1 vccd1 vccd1 _2185_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_25_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1969_ _1969_/A _2505_/Q vssd1 vssd1 vccd1 vccd1 _2501_/D sky130_fd_sc_hd__and2_4
XFILLER_56_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1823_ _2573_/Q _1809_/A _1822_/X vssd1 vssd1 vccd1 vccd1 _2574_/D sky130_fd_sc_hd__o21a_4
XFILLER_22_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1685_ _1681_/X _1684_/Y _1500_/X vssd1 vssd1 vccd1 vccd1 _1685_/X sky130_fd_sc_hd__a21o_4
X_1754_ _1534_/X _2555_/Q _1614_/X vssd1 vssd1 vccd1 vccd1 _1754_/X sky130_fd_sc_hd__o21a_4
X_2237_ _2235_/Y _2236_/A _2236_/Y vssd1 vssd1 vccd1 vccd1 _2237_/Y sky130_fd_sc_hd__a21oi_4
X_2306_ _2304_/A _1602_/C _2306_/C vssd1 vssd1 vccd1 vccd1 _2306_/Y sky130_fd_sc_hd__nand3_4
XFILLER_53_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2168_ _2168_/A _2168_/B vssd1 vssd1 vccd1 vccd1 _2168_/Y sky130_fd_sc_hd__nor2_4
X_2099_ _2104_/A _2098_/Y _2099_/C vssd1 vssd1 vccd1 vccd1 _2463_/D sky130_fd_sc_hd__and3_4
XFILLER_0_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1470_ _1438_/D vssd1 vssd1 vccd1 vccd1 _1470_/X sky130_fd_sc_hd__buf_2
XFILLER_5_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2022_ _2022_/A _2022_/B _2021_/Y vssd1 vssd1 vccd1 vccd1 _2022_/Y sky130_fd_sc_hd__nand3_4
XFILLER_62_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1806_ _2591_/Q _2144_/A _1799_/X vssd1 vssd1 vccd1 vccd1 _1806_/X sky130_fd_sc_hd__o21a_4
X_1737_ _1831_/B vssd1 vssd1 vccd1 vccd1 _1738_/B sky130_fd_sc_hd__inv_2
X_1668_ _1667_/X vssd1 vssd1 vccd1 vccd1 _2168_/A sky130_fd_sc_hd__buf_2
X_1599_ _1597_/X _1488_/X _1598_/X _1564_/A vssd1 vssd1 vccd1 vccd1 _1602_/A sky130_fd_sc_hd__a211o_4
XFILLER_41_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_2_0_m1_clk_local clkbuf_4_3_0_m1_clk_local/A vssd1 vssd1 vccd1 vccd1 _2635_/CLK
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_39_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2640_ _2635_/CLK _1286_/Y vssd1 vssd1 vccd1 vccd1 _1256_/A sky130_fd_sc_hd__dfxtp_4
X_2571_ _2454_/CLK _1832_/Y vssd1 vssd1 vccd1 vccd1 _1829_/A sky130_fd_sc_hd__dfxtp_4
X_1453_ _1450_/X _1452_/Y _2335_/B vssd1 vssd1 vccd1 vccd1 _1453_/Y sky130_fd_sc_hd__o21ai_4
X_1522_ _1470_/X _1448_/A _1213_/X vssd1 vssd1 vccd1 vccd1 _1522_/Y sky130_fd_sc_hd__o21ai_4
X_2005_ _2011_/A _2020_/A _2492_/Q CLK_LED vssd1 vssd1 vccd1 vccd1 _2006_/C sky130_fd_sc_hd__nand4_4
XFILLER_55_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1384_ _2622_/Q _1390_/B _1374_/X vssd1 vssd1 vccd1 vccd1 _1384_/X sky130_fd_sc_hd__o21a_4
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2554_ _2561_/CLK _2554_/D vssd1 vssd1 vccd1 vccd1 _2554_/Q sky130_fd_sc_hd__dfxtp_4
X_2623_ _2623_/CLK _2623_/D vssd1 vssd1 vccd1 vccd1 _1236_/B sky130_fd_sc_hd__dfxtp_4
X_2485_ _2511_/CLK _2044_/X vssd1 vssd1 vccd1 vccd1 _2043_/D sky130_fd_sc_hd__dfxtp_4
X_1367_ _1367_/A _1366_/X _1360_/A _1238_/D vssd1 vssd1 vccd1 vccd1 _1367_/Y sky130_fd_sc_hd__nand4_4
X_1436_ _2609_/Q _1436_/B _2607_/Q _1486_/A vssd1 vssd1 vccd1 vccd1 _1438_/A sky130_fd_sc_hd__and4_4
X_1505_ _1504_/Y _1487_/B _1486_/X _1488_/A vssd1 vssd1 vccd1 vccd1 _1505_/Y sky130_fd_sc_hd__nand4_4
X_1298_ _1346_/A vssd1 vssd1 vccd1 vccd1 _2022_/B sky130_fd_sc_hd__buf_2
XFILLER_28_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1221_ _2101_/A vssd1 vssd1 vccd1 vccd1 _1222_/A sky130_fd_sc_hd__buf_2
XFILLER_6_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2270_ _2246_/Y vssd1 vssd1 vccd1 vccd1 _2270_/X sky130_fd_sc_hd__buf_2
XFILLER_52_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1985_ _1985_/A vssd1 vssd1 vccd1 vccd1 _1985_/Y sky130_fd_sc_hd__inv_2
XFILLER_20_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2537_ _2521_/CLK _2537_/D vssd1 vssd1 vccd1 vccd1 _2537_/Q sky130_fd_sc_hd__dfxtp_4
X_2606_ _2611_/CLK _2606_/D vssd1 vssd1 vccd1 vccd1 _1486_/A sky130_fd_sc_hd__dfxtp_4
X_2468_ _2646_/CLK _2468_/D vssd1 vssd1 vccd1 vccd1 _2104_/D sky130_fd_sc_hd__dfxtp_4
X_1419_ _1419_/A _2010_/B _1419_/C vssd1 vssd1 vccd1 vccd1 _1419_/X sky130_fd_sc_hd__and3_4
X_2399_ _2399_/CLK _2399_/D vssd1 vssd1 vccd1 vccd1 _1750_/A sky130_fd_sc_hd__dfxtp_4
XPHY_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1770_ _1770_/A vssd1 vssd1 vccd1 vccd1 _1770_/Y sky130_fd_sc_hd__inv_2
X_1204_ _2170_/B _1188_/X _1191_/X vssd1 vssd1 vccd1 vccd1 _1204_/Y sky130_fd_sc_hd__o21ai_4
X_2322_ _2322_/A _2322_/B vssd1 vssd1 vccd1 vccd1 _2322_/Y sky130_fd_sc_hd__nand2_4
X_2184_ _1225_/A _2148_/X _1856_/C _1649_/Y vssd1 vssd1 vccd1 vccd1 _2184_/Y sky130_fd_sc_hd__a2bb2oi_4
XFILLER_33_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2253_ _2257_/A _1698_/A _2136_/A vssd1 vssd1 vccd1 vccd1 _2253_/Y sky130_fd_sc_hd__nand3_4
XFILLER_65_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1899_ _2093_/A _2548_/Q vssd1 vssd1 vccd1 vccd1 _2544_/D sky130_fd_sc_hd__and2_4
X_1968_ _1969_/A _1968_/B vssd1 vssd1 vccd1 vccd1 _2502_/D sky130_fd_sc_hd__and2_4
XFILLER_48_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1822_ _2574_/Q _2461_/Q _1813_/X vssd1 vssd1 vccd1 vccd1 _1822_/X sky130_fd_sc_hd__o21a_4
X_1753_ _1749_/X _1752_/X _1472_/A vssd1 vssd1 vccd1 vccd1 _1753_/X sky130_fd_sc_hd__a21o_4
X_1684_ _2337_/B _1683_/Y _1444_/Y vssd1 vssd1 vccd1 vccd1 _1684_/Y sky130_fd_sc_hd__nand3_4
X_2167_ _2147_/Y _2165_/Y _2166_/Y vssd1 vssd1 vccd1 vccd1 _2167_/Y sky130_fd_sc_hd__o21ai_4
X_2236_ _2236_/A _1218_/A vssd1 vssd1 vccd1 vccd1 _2236_/Y sky130_fd_sc_hd__nor2_4
X_2305_ _1503_/Y _2292_/X _2304_/Y vssd1 vssd1 vccd1 vccd1 _2305_/Y sky130_fd_sc_hd__o21ai_4
X_2098_ _2452_/Q vssd1 vssd1 vccd1 vccd1 _2098_/Y sky130_fd_sc_hd__inv_2
XFILLER_21_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_10_0_m1_clk_local clkbuf_3_5_0_m1_clk_local/X vssd1 vssd1 vccd1 vccd1 _2511_/CLK
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_44_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2021_ _2002_/X _2013_/D _2003_/Y vssd1 vssd1 vccd1 vccd1 _2021_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_35_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1736_ _1736_/A _1839_/A vssd1 vssd1 vccd1 vccd1 _1831_/B sky130_fd_sc_hd__nor2_4
X_1805_ _1786_/Y _2573_/Q _1804_/X vssd1 vssd1 vccd1 vccd1 _1805_/X sky130_fd_sc_hd__o21a_4
X_1667_ _1559_/Y _1648_/A _1667_/C _1667_/D vssd1 vssd1 vccd1 vccd1 _1667_/X sky130_fd_sc_hd__and4_4
X_1598_ _1577_/A _2390_/Q _2580_/Q vssd1 vssd1 vccd1 vccd1 _1598_/X sky130_fd_sc_hd__o21a_4
XFILLER_41_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2219_ _2089_/Y _1624_/X _2218_/Y vssd1 vssd1 vccd1 vccd1 _2219_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_14_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2570_ _2646_/CLK _2570_/D vssd1 vssd1 vccd1 vccd1 _1830_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_40_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1383_ _1394_/B _2621_/Q _1383_/C _2619_/Q vssd1 vssd1 vccd1 vccd1 _1390_/B sky130_fd_sc_hd__and4_4
X_1452_ _1440_/B _1439_/X _1451_/X vssd1 vssd1 vccd1 vccd1 _1452_/Y sky130_fd_sc_hd__a21oi_4
X_1521_ _2144_/A _1460_/X _1462_/X vssd1 vssd1 vccd1 vccd1 _1521_/Y sky130_fd_sc_hd__a21oi_4
X_2004_ _2002_/X _2003_/Y _2008_/A vssd1 vssd1 vccd1 vccd1 _2020_/A sky130_fd_sc_hd__nor3_4
Xclkbuf_4_7_0_addressalyzerBlock.SPI_CLK clkbuf_4_7_0_addressalyzerBlock.SPI_CLK/A
+ vssd1 vssd1 vccd1 vccd1 _2561_/CLK sky130_fd_sc_hd__clkbuf_1
X_1719_ _1719_/A _1854_/B vssd1 vssd1 vccd1 vccd1 _1719_/X sky130_fd_sc_hd__or2_4
XFILLER_58_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2553_ _2561_/CLK _2553_/D vssd1 vssd1 vccd1 vccd1 _2553_/Q sky130_fd_sc_hd__dfxtp_4
X_2622_ _2619_/CLK _2622_/D vssd1 vssd1 vccd1 vccd1 _2622_/Q sky130_fd_sc_hd__dfxtp_4
X_1504_ _1504_/A vssd1 vssd1 vccd1 vccd1 _1504_/Y sky130_fd_sc_hd__inv_2
X_2484_ _2470_/CLK _2046_/Y vssd1 vssd1 vccd1 vccd1 _1987_/A sky130_fd_sc_hd__dfxtp_4
X_1366_ _1366_/A vssd1 vssd1 vccd1 vccd1 _1366_/X sky130_fd_sc_hd__buf_2
X_1435_ _1434_/Y vssd1 vssd1 vccd1 vccd1 _1488_/A sky130_fd_sc_hd__inv_2
X_1297_ _1297_/A vssd1 vssd1 vccd1 vccd1 _1297_/Y sky130_fd_sc_hd__inv_2
XFILLER_23_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1220_ _1219_/X vssd1 vssd1 vccd1 vccd1 _2101_/A sky130_fd_sc_hd__buf_2
XFILLER_45_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1984_ _1984_/A vssd1 vssd1 vccd1 vccd1 _2002_/A sky130_fd_sc_hd__inv_2
XFILLER_9_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2467_ _2454_/CLK _2467_/D vssd1 vssd1 vccd1 vccd1 _2091_/A sky130_fd_sc_hd__dfxtp_4
X_2536_ _2538_/CLK _2536_/D vssd1 vssd1 vccd1 vccd1 HASH_ADDR[5] sky130_fd_sc_hd__dfxtp_4
X_2605_ _2389_/CLK _1523_/Y vssd1 vssd1 vccd1 vccd1 _1483_/B sky130_fd_sc_hd__dfxtp_4
X_1349_ _1349_/A vssd1 vssd1 vccd1 vccd1 _1351_/A sky130_fd_sc_hd__inv_2
X_1418_ _1409_/A _1406_/X vssd1 vssd1 vccd1 vccd1 _1419_/A sky130_fd_sc_hd__or2_4
XFILLER_28_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2398_ _2399_/CLK _2398_/D vssd1 vssd1 vccd1 vccd1 _2398_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2321_ _2224_/B _2310_/X _2144_/A _2312_/X vssd1 vssd1 vccd1 vccd1 _2321_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_65_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1203_ _2647_/Q _1194_/B _1202_/X vssd1 vssd1 vccd1 vccd1 _1203_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_26_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2252_ _2244_/X _2133_/Y _2247_/X _1904_/Y _2249_/X vssd1 vssd1 vccd1 vccd1 _2431_/D
+ sky130_fd_sc_hd__o32ai_4
X_2183_ _2180_/X _2182_/X _1701_/A vssd1 vssd1 vccd1 vccd1 _2183_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_65_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1898_ _2096_/A vssd1 vssd1 vccd1 vccd1 _2093_/A sky130_fd_sc_hd__buf_2
X_1967_ _1284_/X _1966_/Y vssd1 vssd1 vccd1 vccd1 _1967_/Y sky130_fd_sc_hd__nor2_4
X_2519_ _2519_/CLK _1940_/Y vssd1 vssd1 vccd1 vccd1 _2519_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1683_ _1683_/A vssd1 vssd1 vccd1 vccd1 _1683_/Y sky130_fd_sc_hd__inv_2
X_1821_ _2574_/Q _1809_/X _1820_/X vssd1 vssd1 vccd1 vccd1 _2575_/D sky130_fd_sc_hd__o21a_4
X_1752_ _2443_/Q _1751_/A _1633_/X _1751_/Y vssd1 vssd1 vccd1 vccd1 _1752_/X sky130_fd_sc_hd__a211o_4
X_2304_ _2304_/A _1602_/C _1409_/A vssd1 vssd1 vccd1 vccd1 _2304_/Y sky130_fd_sc_hd__nand3_4
XFILLER_65_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2097_ _2107_/A _2097_/B vssd1 vssd1 vccd1 vccd1 _2464_/D sky130_fd_sc_hd__and2_4
XFILLER_57_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2166_ _1673_/B THREAD_COUNT[3] vssd1 vssd1 vccd1 vccd1 _2166_/Y sky130_fd_sc_hd__nand2_4
X_2235_ _2233_/Y _2235_/B vssd1 vssd1 vccd1 vccd1 _2235_/Y sky130_fd_sc_hd__nand2_4
XFILLER_21_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2020_ _2020_/A vssd1 vssd1 vccd1 vccd1 _2022_/A sky130_fd_sc_hd__inv_2
XFILLER_47_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1735_ _1829_/A _1202_/B _1830_/B _1830_/C vssd1 vssd1 vccd1 vccd1 _1831_/A sky130_fd_sc_hd__nand4_4
X_1666_ _1666_/A vssd1 vssd1 vccd1 vccd1 _1673_/B sky130_fd_sc_hd__buf_2
X_1804_ _2591_/Q _1514_/X _1799_/X vssd1 vssd1 vccd1 vccd1 _1804_/X sky130_fd_sc_hd__o21a_4
X_1597_ _1664_/A vssd1 vssd1 vccd1 vccd1 _1597_/X sky130_fd_sc_hd__buf_2
XFILLER_38_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2149_ _1534_/A _2554_/Q _2148_/X vssd1 vssd1 vccd1 vccd1 _2149_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_26_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2218_ _1625_/X _2411_/Q _1704_/A vssd1 vssd1 vccd1 vccd1 _2218_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_14_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_1_0_m1_clk_local clkbuf_0_m1_clk_local/X vssd1 vssd1 vccd1 vccd1 clkbuf_2_3_0_m1_clk_local/A
+ sky130_fd_sc_hd__clkbuf_1
X_1520_ _2580_/Q vssd1 vssd1 vccd1 vccd1 _2144_/A sky130_fd_sc_hd__buf_2
X_1382_ _1376_/C _1366_/X _1381_/Y vssd1 vssd1 vccd1 vccd1 _2623_/D sky130_fd_sc_hd__o21a_4
Xclkbuf_4_12_0_addressalyzerBlock.SPI_CLK clkbuf_3_6_0_addressalyzerBlock.SPI_CLK/X
+ vssd1 vssd1 vccd1 vccd1 _2437_/CLK sky130_fd_sc_hd__clkbuf_1
X_1451_ _1434_/Y vssd1 vssd1 vccd1 vccd1 _1451_/X sky130_fd_sc_hd__buf_2
XFILLER_4_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2003_ _1999_/A vssd1 vssd1 vccd1 vccd1 _2003_/Y sky130_fd_sc_hd__inv_2
XFILLER_50_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1649_ _1659_/A _1648_/Y vssd1 vssd1 vccd1 vccd1 _1649_/Y sky130_fd_sc_hd__nor2_4
X_1718_ _1702_/Y _1717_/Y _1614_/X vssd1 vssd1 vccd1 vccd1 _1718_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_58_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2483_ _2511_/CLK _2050_/Y vssd1 vssd1 vccd1 vccd1 _2483_/Q sky130_fd_sc_hd__dfxtp_4
X_2621_ _2619_/CLK _1390_/Y vssd1 vssd1 vccd1 vccd1 _2621_/Q sky130_fd_sc_hd__dfxtp_4
X_2552_ _2552_/CLK _2552_/D vssd1 vssd1 vccd1 vccd1 _2552_/Q sky130_fd_sc_hd__dfxtp_4
X_1503_ _1503_/A vssd1 vssd1 vccd1 vccd1 _1503_/Y sky130_fd_sc_hd__inv_2
X_1365_ _1394_/B _1383_/C _2619_/Q _1365_/D vssd1 vssd1 vccd1 vccd1 _1366_/A sky130_fd_sc_hd__and4_4
X_1434_ _2386_/Q _1729_/B vssd1 vssd1 vccd1 vccd1 _1434_/Y sky130_fd_sc_hd__nor2_4
X_1296_ _1294_/Y _1295_/Y vssd1 vssd1 vccd1 vccd1 _1297_/A sky130_fd_sc_hd__nand2_4
XFILLER_11_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_3_4_0_m1_clk_local clkbuf_3_5_0_m1_clk_local/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_9_0_m1_clk_local/A
+ sky130_fd_sc_hd__clkbuf_1
X_1983_ _2092_/A _1983_/B vssd1 vssd1 vccd1 vccd1 _2494_/D sky130_fd_sc_hd__nor2_4
X_2604_ _2604_/CLK _2604_/D vssd1 vssd1 vccd1 vccd1 _2604_/Q sky130_fd_sc_hd__dfxtp_4
X_2466_ _2464_/CLK _2466_/D vssd1 vssd1 vccd1 vccd1 _2351_/C sky130_fd_sc_hd__dfxtp_4
X_1417_ _1417_/A vssd1 vssd1 vccd1 vccd1 _1417_/Y sky130_fd_sc_hd__inv_2
X_2535_ _2538_/CLK _1917_/X vssd1 vssd1 vccd1 vccd1 HASH_ADDR[4] sky130_fd_sc_hd__dfxtp_4
X_1348_ _1347_/Y vssd1 vssd1 vccd1 vccd1 _1348_/Y sky130_fd_sc_hd__inv_2
XFILLER_36_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1279_ _1278_/Y vssd1 vssd1 vccd1 vccd1 _2642_/D sky130_fd_sc_hd__inv_2
X_2397_ _2604_/CLK _2319_/X vssd1 vssd1 vccd1 vccd1 _2397_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2251_ _2244_/X _2130_/Y _2247_/X _1902_/Y _2249_/X vssd1 vssd1 vccd1 vccd1 _2432_/D
+ sky130_fd_sc_hd__o32ai_4
X_2320_ _1764_/Y _2310_/X _1514_/X _2312_/X vssd1 vssd1 vccd1 vccd1 _2320_/X sky130_fd_sc_hd__a2bb2o_4
X_1202_ _1202_/A _1202_/B vssd1 vssd1 vccd1 vccd1 _1202_/X sky130_fd_sc_hd__or2_4
X_2182_ _2441_/Q _1635_/X _1632_/Y _2181_/Y vssd1 vssd1 vccd1 vccd1 _2182_/X sky130_fd_sc_hd__a211o_4
X_1966_ _2439_/Q vssd1 vssd1 vccd1 vccd1 _1966_/Y sky130_fd_sc_hd__inv_2
X_1897_ _1895_/A _2549_/Q vssd1 vssd1 vccd1 vccd1 _2545_/D sky130_fd_sc_hd__and2_4
X_2449_ _2552_/CLK _2449_/D vssd1 vssd1 vccd1 vccd1 _2449_/Q sky130_fd_sc_hd__dfxtp_4
X_2518_ _2513_/CLK _1942_/Y vssd1 vssd1 vccd1 vccd1 _2518_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_56_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1820_ _2575_/Q _1810_/X _1813_/X vssd1 vssd1 vccd1 vccd1 _1820_/X sky130_fd_sc_hd__o21a_4
XFILLER_15_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1682_ _1566_/X _2335_/D _1683_/A _2385_/Q _1681_/X vssd1 vssd1 vccd1 vccd1 _1682_/Y
+ sky130_fd_sc_hd__o41ai_4
X_1751_ _1751_/A _1750_/Y vssd1 vssd1 vccd1 vccd1 _1751_/Y sky130_fd_sc_hd__nor2_4
X_2234_ _1661_/B _2543_/Q _1661_/D _2234_/D vssd1 vssd1 vccd1 vccd1 _2235_/B sky130_fd_sc_hd__or4_4
X_2303_ _2136_/Y _2291_/X _2302_/Y vssd1 vssd1 vccd1 vccd1 _2406_/D sky130_fd_sc_hd__o21ai_4
X_2096_ _2096_/A vssd1 vssd1 vccd1 vccd1 _2107_/A sky130_fd_sc_hd__buf_2
X_2165_ _2162_/Y _2163_/X _2164_/X vssd1 vssd1 vccd1 vccd1 _2165_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_61_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1949_ _1963_/A _1948_/Y vssd1 vssd1 vccd1 vccd1 _2515_/D sky130_fd_sc_hd__nor2_4
XFILLER_56_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1803_ _1786_/Y _2574_/Q _1802_/X vssd1 vssd1 vccd1 vccd1 _1803_/X sky130_fd_sc_hd__o21a_4
X_1734_ _1733_/Y vssd1 vssd1 vccd1 vccd1 _2592_/D sky130_fd_sc_hd__inv_2
X_1665_ _1570_/A _1664_/Y _1660_/A vssd1 vssd1 vccd1 vccd1 _1666_/A sky130_fd_sc_hd__nor3_4
X_1596_ _1545_/X _1576_/X _1588_/Y _1593_/Y _1595_/X vssd1 vssd1 vccd1 vccd1 _2598_/D
+ sky130_fd_sc_hd__a41oi_4
XFILLER_38_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2217_ _1534_/X _2551_/Q _1854_/B vssd1 vssd1 vccd1 vccd1 _2217_/Y sky130_fd_sc_hd__o21ai_4
X_2079_ _2079_/A _1991_/B _2473_/Q vssd1 vssd1 vccd1 vccd1 _2084_/C sky130_fd_sc_hd__nand3_4
X_2148_ _1613_/Y vssd1 vssd1 vccd1 vccd1 _2148_/X sky130_fd_sc_hd__buf_2
XFILLER_14_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1450_ _1446_/Y vssd1 vssd1 vccd1 vccd1 _1450_/X sky130_fd_sc_hd__buf_2
XFILLER_4_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1381_ _1376_/C _1395_/B _1385_/D _1365_/D _1275_/X vssd1 vssd1 vccd1 vccd1 _1381_/Y
+ sky130_fd_sc_hd__a41oi_4
X_2002_ _2002_/A vssd1 vssd1 vccd1 vccd1 _2002_/X sky130_fd_sc_hd__buf_2
XFILLER_50_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1648_ _1648_/A vssd1 vssd1 vccd1 vccd1 _1648_/Y sky130_fd_sc_hd__inv_2
X_1579_ _1567_/A vssd1 vssd1 vccd1 vccd1 _1579_/X sky130_fd_sc_hd__buf_2
X_1717_ _1712_/Y _1633_/X _1716_/Y vssd1 vssd1 vccd1 vccd1 _1717_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_66_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2620_ _2470_/CLK _2620_/D vssd1 vssd1 vccd1 vccd1 _2620_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_9_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2482_ _2511_/CLK _2482_/D vssd1 vssd1 vccd1 vccd1 _1985_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_49_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2551_ _2551_/CLK _2551_/D vssd1 vssd1 vccd1 vccd1 _2551_/Q sky130_fd_sc_hd__dfxtp_4
X_1502_ _1496_/Y _1498_/Y _1501_/X vssd1 vssd1 vccd1 vccd1 _1502_/Y sky130_fd_sc_hd__a21oi_4
X_1433_ _1432_/X vssd1 vssd1 vccd1 vccd1 _1440_/B sky130_fd_sc_hd__buf_2
X_1364_ _2620_/Q vssd1 vssd1 vccd1 vccd1 _1383_/C sky130_fd_sc_hd__buf_2
X_1295_ _1295_/A _1308_/A _1299_/A _1295_/D vssd1 vssd1 vccd1 vccd1 _1295_/Y sky130_fd_sc_hd__nand4_4
XFILLER_23_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_2_3_0_addressalyzerBlock.SPI_CLK clkbuf_2_3_0_addressalyzerBlock.SPI_CLK/A
+ vssd1 vssd1 vccd1 vccd1 clkbuf_3_6_0_addressalyzerBlock.SPI_CLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_52_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1982_ _1981_/X vssd1 vssd1 vccd1 vccd1 _2495_/D sky130_fd_sc_hd__inv_2
XFILLER_45_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2534_ _2492_/CLK _1918_/X vssd1 vssd1 vccd1 vccd1 HASH_ADDR[3] sky130_fd_sc_hd__dfxtp_4
XFILLER_9_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2603_ _2389_/CLK _2603_/D vssd1 vssd1 vccd1 vccd1 _1483_/D sky130_fd_sc_hd__dfxtp_4
X_2465_ _2464_/CLK _2465_/D vssd1 vssd1 vccd1 vccd1 _2465_/Q sky130_fd_sc_hd__dfxtp_4
X_1416_ _1413_/Y _1419_/C _1415_/Y vssd1 vssd1 vccd1 vccd1 _1417_/A sky130_fd_sc_hd__o21ai_4
X_1347_ _1344_/X _1347_/B _1346_/X vssd1 vssd1 vccd1 vccd1 _1347_/Y sky130_fd_sc_hd__nand3_4
X_2396_ _2389_/CLK _2320_/X vssd1 vssd1 vccd1 vccd1 _1764_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_51_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1278_ _1276_/Y _1277_/Y vssd1 vssd1 vccd1 vccd1 _1278_/Y sky130_fd_sc_hd__nand2_4
XPHY_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1201_ _1199_/Y _1187_/X _1200_/Y vssd1 vssd1 vccd1 vccd1 _2649_/D sky130_fd_sc_hd__a21oi_4
XFILLER_40_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2250_ _2244_/X _2127_/Y _2247_/X _1710_/B _2249_/X vssd1 vssd1 vccd1 vccd1 _2433_/D
+ sky130_fd_sc_hd__o32ai_4
X_2181_ _2181_/A _1771_/Y vssd1 vssd1 vccd1 vccd1 _2181_/Y sky130_fd_sc_hd__nor2_4
XFILLER_18_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1965_ _1284_/X _1965_/B vssd1 vssd1 vccd1 vccd1 _2504_/D sky130_fd_sc_hd__nor2_4
X_1896_ _1895_/A _1896_/B vssd1 vssd1 vccd1 vccd1 _1896_/X sky130_fd_sc_hd__and2_4
X_2517_ _2538_/CLK _2517_/D vssd1 vssd1 vccd1 vccd1 _1957_/B sky130_fd_sc_hd__dfxtp_4
X_2379_ _2508_/CLK _2379_/D vssd1 vssd1 vccd1 vccd1 _2379_/Q sky130_fd_sc_hd__dfxtp_4
X_2448_ _2551_/CLK _2448_/D vssd1 vssd1 vccd1 vccd1 _2448_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1750_ _1750_/A vssd1 vssd1 vccd1 vccd1 _1750_/Y sky130_fd_sc_hd__inv_2
XFILLER_15_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1681_ _1679_/Y _1680_/X _1530_/C vssd1 vssd1 vccd1 vccd1 _1681_/X sky130_fd_sc_hd__o21a_4
X_2233_ _2216_/Y _2231_/Y _2232_/Y vssd1 vssd1 vccd1 vccd1 _2233_/Y sky130_fd_sc_hd__o21ai_4
X_2164_ _1741_/A _1376_/B _1656_/A vssd1 vssd1 vccd1 vccd1 _2164_/X sky130_fd_sc_hd__a21o_4
XFILLER_31_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2302_ _2304_/A _1602_/C HASH_LED vssd1 vssd1 vccd1 vccd1 _2302_/Y sky130_fd_sc_hd__nand3_4
XFILLER_65_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2095_ _2093_/A IRQ_OUT_fromClient vssd1 vssd1 vccd1 vccd1 _2465_/D sky130_fd_sc_hd__and2_4
XFILLER_53_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1879_ _1878_/A DATA_FROM_HASH[1] vssd1 vssd1 vccd1 vccd1 _1879_/X sky130_fd_sc_hd__and2_4
X_1948_ _2419_/Q vssd1 vssd1 vccd1 vccd1 _1948_/Y sky130_fd_sc_hd__inv_2
XFILLER_21_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1733_ _1730_/X _1731_/Y _1732_/Y vssd1 vssd1 vccd1 vccd1 _1733_/Y sky130_fd_sc_hd__o21ai_4
X_1802_ _2591_/Q _1503_/A _1799_/X vssd1 vssd1 vccd1 vccd1 _1802_/X sky130_fd_sc_hd__o21a_4
X_1664_ _1664_/A _1579_/X _1567_/B vssd1 vssd1 vccd1 vccd1 _1664_/Y sky130_fd_sc_hd__nand3_4
X_1595_ _1541_/X _1594_/X _1781_/A vssd1 vssd1 vccd1 vccd1 _1595_/X sky130_fd_sc_hd__a21o_4
X_2147_ _1230_/A _1571_/A _1661_/C _1661_/D _2146_/Y vssd1 vssd1 vccd1 vccd1 _2147_/Y
+ sky130_fd_sc_hd__o41ai_4
X_2216_ _1406_/X _1661_/B _1661_/C _1661_/D _2146_/Y vssd1 vssd1 vccd1 vccd1 _2216_/Y
+ sky130_fd_sc_hd__o41ai_4
XFILLER_53_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2078_ _1991_/A vssd1 vssd1 vccd1 vccd1 _2079_/A sky130_fd_sc_hd__buf_2
XFILLER_39_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1380_ _1383_/C vssd1 vssd1 vccd1 vccd1 _1385_/D sky130_fd_sc_hd__buf_2
XFILLER_4_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2001_ _2010_/C _2001_/B vssd1 vssd1 vccd1 vccd1 _2001_/Y sky130_fd_sc_hd__nand2_4
XFILLER_31_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1716_ _1715_/X _1534_/A vssd1 vssd1 vccd1 vccd1 _1716_/Y sky130_fd_sc_hd__nand2_4
XFILLER_58_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1647_ _1667_/C _1667_/D vssd1 vssd1 vccd1 vccd1 _1659_/A sky130_fd_sc_hd__nand2_4
X_1578_ _2335_/D _1460_/X _1503_/A vssd1 vssd1 vccd1 vccd1 _1578_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_66_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2550_ _2464_/CLK _1891_/X vssd1 vssd1 vccd1 vccd1 _1896_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_9_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2481_ _2511_/CLK _2057_/X vssd1 vssd1 vccd1 vccd1 _2481_/Q sky130_fd_sc_hd__dfxtp_4
X_1363_ _1363_/A _1231_/Y _1363_/C vssd1 vssd1 vccd1 vccd1 _1394_/B sky130_fd_sc_hd__nor3_4
X_1432_ _1432_/A _1701_/A _1466_/A _1467_/A vssd1 vssd1 vccd1 vccd1 _1432_/X sky130_fd_sc_hd__and4_4
X_1501_ _1450_/X _1499_/Y _1500_/X vssd1 vssd1 vccd1 vccd1 _1501_/X sky130_fd_sc_hd__a21o_4
XFILLER_55_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1294_ _1301_/A _1293_/Y _1275_/X vssd1 vssd1 vccd1 vccd1 _1294_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_10_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1981_ _1972_/A _1869_/A _1867_/Y vssd1 vssd1 vccd1 vccd1 _1981_/X sky130_fd_sc_hd__or3_4
XFILLER_60_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2602_ _2389_/CLK _1551_/Y vssd1 vssd1 vccd1 vccd1 _1467_/A sky130_fd_sc_hd__dfxtp_4
X_2533_ _2519_/CLK _2533_/D vssd1 vssd1 vccd1 vccd1 HASH_ADDR[2] sky130_fd_sc_hd__dfxtp_4
X_2464_ _2464_/CLK _2464_/D vssd1 vssd1 vccd1 vccd1 _2464_/Q sky130_fd_sc_hd__dfxtp_4
X_1346_ _1346_/A vssd1 vssd1 vccd1 vccd1 _1346_/X sky130_fd_sc_hd__buf_2
X_1415_ _1419_/C _1413_/Y _1388_/A vssd1 vssd1 vccd1 vccd1 _1415_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_3_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2395_ _2604_/CLK _2321_/X vssd1 vssd1 vccd1 vccd1 _1767_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_51_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1277_ _1273_/A _1277_/B _2641_/Q _1256_/A vssd1 vssd1 vccd1 vccd1 _1277_/Y sky130_fd_sc_hd__nand4_4
XFILLER_11_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1200_ _1762_/B _1188_/X _1191_/X vssd1 vssd1 vccd1 vccd1 _1200_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_33_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2180_ _2176_/Y _2179_/Y _2449_/Q vssd1 vssd1 vccd1 vccd1 _2180_/X sky130_fd_sc_hd__a21o_4
XFILLER_65_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1895_ _1895_/A DATA_AVAILABLE[0] vssd1 vssd1 vccd1 vccd1 _2547_/D sky130_fd_sc_hd__and2_4
Xclkbuf_3_0_0_m1_clk_local clkbuf_3_1_0_m1_clk_local/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_0_0_m1_clk_local/X
+ sky130_fd_sc_hd__clkbuf_1
X_1964_ _2440_/Q vssd1 vssd1 vccd1 vccd1 _1965_/B sky130_fd_sc_hd__inv_2
XFILLER_21_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2447_ _2551_/CLK _2447_/D vssd1 vssd1 vccd1 vccd1 _2447_/Q sky130_fd_sc_hd__dfxtp_4
X_2516_ _2632_/CLK _1947_/Y vssd1 vssd1 vccd1 vccd1 _2516_/Q sky130_fd_sc_hd__dfxtp_4
X_2378_ _2508_/CLK _2377_/Q vssd1 vssd1 vccd1 vccd1 _2379_/D sky130_fd_sc_hd__dfxtp_4
XFILLER_56_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1329_ _1332_/A vssd1 vssd1 vccd1 vccd1 _1329_/X sky130_fd_sc_hd__buf_2
XFILLER_33_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1680_ _1185_/A _2462_/Q vssd1 vssd1 vccd1 vccd1 _1680_/X sky130_fd_sc_hd__or2_4
X_2301_ _1490_/Y _2291_/X _2300_/Y vssd1 vssd1 vccd1 vccd1 _2407_/D sky130_fd_sc_hd__o21ai_4
XFILLER_65_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2232_ THREAD_COUNT[0] _1673_/B _2168_/Y vssd1 vssd1 vccd1 vccd1 _2232_/Y sky130_fd_sc_hd__a21boi_4
X_2163_ _2632_/Q _1646_/X _1741_/Y vssd1 vssd1 vccd1 vccd1 _2163_/X sky130_fd_sc_hd__o21a_4
XFILLER_38_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2094_ _2093_/A _2465_/Q vssd1 vssd1 vccd1 vccd1 _2466_/D sky130_fd_sc_hd__and2_4
XFILLER_0_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1878_ _1878_/A DATA_FROM_HASH[2] vssd1 vssd1 vccd1 vccd1 _2561_/D sky130_fd_sc_hd__and2_4
X_1947_ _1963_/A _1946_/Y vssd1 vssd1 vccd1 vccd1 _1947_/Y sky130_fd_sc_hd__nor2_4
XFILLER_56_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1663_ _1663_/A vssd1 vssd1 vccd1 vccd1 _1761_/A sky130_fd_sc_hd__buf_2
X_1732_ _1730_/X _1761_/A _1781_/A vssd1 vssd1 vccd1 vccd1 _1732_/Y sky130_fd_sc_hd__a21oi_4
X_1801_ _1786_/Y _2575_/Q _1800_/X vssd1 vssd1 vccd1 vccd1 _1801_/X sky130_fd_sc_hd__o21a_4
X_1594_ _1589_/Y vssd1 vssd1 vccd1 vccd1 _1594_/X sky130_fd_sc_hd__buf_2
X_2215_ _1676_/A _2213_/Y _2214_/Y vssd1 vssd1 vccd1 vccd1 _2436_/D sky130_fd_sc_hd__o21ai_4
X_2077_ _2071_/Y _2072_/B _2076_/Y vssd1 vssd1 vccd1 vccd1 _2077_/Y sky130_fd_sc_hd__a21oi_4
X_2146_ _1666_/A vssd1 vssd1 vccd1 vccd1 _2146_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2000_ CLK_LED vssd1 vssd1 vccd1 vccd1 _2001_/B sky130_fd_sc_hd__inv_2
Xclkbuf_3_3_0_addressalyzerBlock.SPI_CLK clkbuf_3_3_0_addressalyzerBlock.SPI_CLK/A
+ vssd1 vssd1 vccd1 vccd1 clkbuf_4_7_0_addressalyzerBlock.SPI_CLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_35_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_9_0_m1_clk_local clkbuf_4_9_0_m1_clk_local/A vssd1 vssd1 vccd1 vccd1 _2623_/CLK
+ sky130_fd_sc_hd__clkbuf_1
X_1646_ _1645_/Y vssd1 vssd1 vccd1 vccd1 _1646_/X sky130_fd_sc_hd__buf_2
X_1715_ _2445_/Q _2224_/A _1632_/Y _1714_/Y vssd1 vssd1 vccd1 vccd1 _1715_/X sky130_fd_sc_hd__a211o_4
X_1577_ _1577_/A vssd1 vssd1 vccd1 vccd1 _2335_/D sky130_fd_sc_hd__buf_2
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2129_ _2120_/X _2127_/Y _2128_/Y vssd1 vssd1 vccd1 vccd1 _2129_/Y sky130_fd_sc_hd__o21ai_4
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2480_ _2511_/CLK _2063_/Y vssd1 vssd1 vccd1 vccd1 _1993_/C sky130_fd_sc_hd__dfxtp_4
XFILLER_40_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1500_ _2101_/A vssd1 vssd1 vccd1 vccd1 _1500_/X sky130_fd_sc_hd__buf_2
XFILLER_9_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1362_ _1367_/A _1361_/Y _1306_/X vssd1 vssd1 vccd1 vccd1 _1362_/X sky130_fd_sc_hd__o21a_4
X_1293_ _1295_/A vssd1 vssd1 vccd1 vccd1 _1293_/Y sky130_fd_sc_hd__inv_2
X_1431_ _1483_/D vssd1 vssd1 vccd1 vccd1 _1466_/A sky130_fd_sc_hd__buf_2
XFILLER_63_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1629_ _1621_/X _1627_/Y _1628_/X vssd1 vssd1 vccd1 vccd1 _1629_/X sky130_fd_sc_hd__a21o_4
XFILLER_54_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1980_ _1978_/A _1973_/B _1980_/C vssd1 vssd1 vccd1 vccd1 _2496_/D sky130_fd_sc_hd__and3_4
XFILLER_26_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2532_ _2492_/CLK _1920_/X vssd1 vssd1 vccd1 vccd1 HASH_ADDR[1] sky130_fd_sc_hd__dfxtp_4
XFILLER_54_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2463_ _2646_/CLK _2463_/D vssd1 vssd1 vccd1 vccd1 _1839_/A sky130_fd_sc_hd__dfxtp_4
X_2601_ _2389_/CLK _1557_/X vssd1 vssd1 vccd1 vccd1 _1424_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_5_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1414_ _1409_/A _1406_/X vssd1 vssd1 vccd1 vccd1 _1419_/C sky130_fd_sc_hd__nand2_4
X_1345_ _1333_/Y vssd1 vssd1 vccd1 vccd1 _1347_/B sky130_fd_sc_hd__inv_2
X_2394_ _2437_/CLK _2325_/X vssd1 vssd1 vccd1 vccd1 _1687_/A sky130_fd_sc_hd__dfxtp_4
X_1276_ _1272_/Y _1854_/A _1275_/X vssd1 vssd1 vccd1 vccd1 _1276_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_28_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1894_ _1895_/A DATA_AVAILABLE[1] vssd1 vssd1 vccd1 vccd1 _2548_/D sky130_fd_sc_hd__and2_4
X_1963_ _1963_/A _1963_/B vssd1 vssd1 vccd1 vccd1 _2505_/D sky130_fd_sc_hd__nor2_4
X_2446_ _2446_/CLK _2446_/D vssd1 vssd1 vccd1 vccd1 _2125_/C sky130_fd_sc_hd__dfxtp_4
X_2515_ _2635_/CLK _2515_/D vssd1 vssd1 vccd1 vccd1 _2515_/Q sky130_fd_sc_hd__dfxtp_4
X_2377_ _2508_/CLK _2377_/D vssd1 vssd1 vccd1 vccd1 _2377_/Q sky130_fd_sc_hd__dfxtp_4
X_1259_ _1226_/Y vssd1 vssd1 vccd1 vccd1 _1295_/D sky130_fd_sc_hd__inv_2
X_1328_ _2631_/Q vssd1 vssd1 vccd1 vccd1 _1335_/C sky130_fd_sc_hd__buf_2
XFILLER_17_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2231_ _2228_/Y _2229_/Y _2230_/X vssd1 vssd1 vccd1 vccd1 _2231_/Y sky130_fd_sc_hd__a21oi_4
X_2300_ _2304_/A _2300_/B _2407_/Q vssd1 vssd1 vccd1 vccd1 _2300_/Y sky130_fd_sc_hd__nand3_4
XFILLER_65_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2093_ _2093_/A _2457_/Q vssd1 vssd1 vccd1 vccd1 _2467_/D sky130_fd_sc_hd__and2_4
XFILLER_38_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2162_ _2149_/Y _2160_/Y _2161_/Y vssd1 vssd1 vccd1 vccd1 _2162_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_0_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1877_ _1878_/A DATA_FROM_HASH[3] vssd1 vssd1 vccd1 vccd1 _1877_/X sky130_fd_sc_hd__and2_4
X_1946_ _1946_/A vssd1 vssd1 vccd1 vccd1 _1946_/Y sky130_fd_sc_hd__inv_2
X_2429_ _2418_/CLK _2256_/Y vssd1 vssd1 vccd1 vccd1 _2177_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_52_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1800_ _1788_/X _2136_/A _1799_/X vssd1 vssd1 vccd1 vccd1 _1800_/X sky130_fd_sc_hd__o21a_4
XPHY_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1662_ _2236_/A vssd1 vssd1 vccd1 vccd1 _1663_/A sky130_fd_sc_hd__inv_2
X_1731_ _1697_/A _1731_/B _2391_/Q vssd1 vssd1 vccd1 vccd1 _1731_/Y sky130_fd_sc_hd__nor3_4
XFILLER_7_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2214_ _2192_/A _2436_/Q vssd1 vssd1 vccd1 vccd1 _2214_/Y sky130_fd_sc_hd__nand2_4
X_1593_ _1590_/Y _1648_/A _1488_/X vssd1 vssd1 vccd1 vccd1 _1593_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_53_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2076_ _2071_/Y _2072_/B _1346_/X vssd1 vssd1 vccd1 vccd1 _2076_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_38_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2145_ _2144_/Y _2138_/Y _2123_/X _1966_/Y _2139_/X vssd1 vssd1 vccd1 vccd1 _2145_/Y
+ sky130_fd_sc_hd__o32ai_4
XFILLER_61_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1929_ _2411_/Q vssd1 vssd1 vccd1 vccd1 _1929_/Y sky130_fd_sc_hd__inv_2
XFILLER_39_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1645_ _1645_/A vssd1 vssd1 vccd1 vccd1 _1645_/Y sky130_fd_sc_hd__inv_2
X_1576_ _1574_/Y _2337_/B _1445_/A _1445_/D _1185_/A vssd1 vssd1 vccd1 vccd1 _1576_/X
+ sky130_fd_sc_hd__a41o_4
X_1714_ _1630_/X _1713_/Y vssd1 vssd1 vccd1 vccd1 _1714_/Y sky130_fd_sc_hd__nor2_4
XFILLER_66_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2059_ _2059_/A vssd1 vssd1 vccd1 vccd1 _2072_/B sky130_fd_sc_hd__buf_2
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2128_ _2123_/X _2335_/A _2445_/Q vssd1 vssd1 vccd1 vccd1 _2128_/Y sky130_fd_sc_hd__nand3_4
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1430_ _2604_/Q vssd1 vssd1 vccd1 vccd1 _1701_/A sky130_fd_sc_hd__buf_2
XFILLER_55_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1361_ _1360_/Y _1361_/B vssd1 vssd1 vccd1 vccd1 _1361_/Y sky130_fd_sc_hd__nor2_4
X_1292_ _1308_/A _1299_/A _1295_/D vssd1 vssd1 vccd1 vccd1 _1301_/A sky130_fd_sc_hd__nand3_4
XFILLER_63_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1559_ _1570_/A _1604_/A vssd1 vssd1 vccd1 vccd1 _1559_/Y sky130_fd_sc_hd__nor2_4
X_1628_ _2449_/Q vssd1 vssd1 vccd1 vccd1 _1628_/X sky130_fd_sc_hd__buf_2
XFILLER_36_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2600_ _2437_/CLK _1573_/Y vssd1 vssd1 vccd1 vccd1 _2600_/Q sky130_fd_sc_hd__dfxtp_4
X_1413_ _2614_/Q vssd1 vssd1 vccd1 vccd1 _1413_/Y sky130_fd_sc_hd__inv_2
XFILLER_47_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2462_ _2646_/CLK _2462_/D vssd1 vssd1 vccd1 vccd1 _2462_/Q sky130_fd_sc_hd__dfxtp_4
X_2393_ _2646_/CLK _2393_/D vssd1 vssd1 vccd1 vccd1 _1697_/A sky130_fd_sc_hd__dfxtp_4
X_2531_ _2513_/CLK _2531_/D vssd1 vssd1 vccd1 vccd1 HASH_ADDR[0] sky130_fd_sc_hd__dfxtp_4
X_1275_ _1274_/X vssd1 vssd1 vccd1 vccd1 _1275_/X sky130_fd_sc_hd__buf_2
X_1344_ _1353_/A _1321_/X _1329_/X vssd1 vssd1 vccd1 vccd1 _1344_/X sky130_fd_sc_hd__a21o_4
XFILLER_51_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1962_ _2441_/Q vssd1 vssd1 vccd1 vccd1 _1963_/B sky130_fd_sc_hd__inv_2
X_1893_ _1895_/A DATA_AVAILABLE[2] vssd1 vssd1 vccd1 vccd1 _1893_/X sky130_fd_sc_hd__and2_4
X_2376_ _2508_/CLK _2376_/D vssd1 vssd1 vccd1 vccd1 _2377_/D sky130_fd_sc_hd__dfxtp_4
X_2514_ _2505_/CLK _2514_/D vssd1 vssd1 vccd1 vccd1 DATA_TO_HASH[7] sky130_fd_sc_hd__dfxtp_4
X_2445_ _2446_/CLK _2129_/Y vssd1 vssd1 vccd1 vccd1 _2445_/Q sky130_fd_sc_hd__dfxtp_4
X_1327_ _1326_/Y vssd1 vssd1 vccd1 vccd1 _2633_/D sky130_fd_sc_hd__inv_2
X_1258_ _1351_/B _1240_/Y _1238_/Y vssd1 vssd1 vccd1 vccd1 _1258_/Y sky130_fd_sc_hd__nor3_4
X_1189_ _2384_/Q vssd1 vssd1 vccd1 vccd1 _1190_/A sky130_fd_sc_hd__inv_2
XPHY_207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2230_ _1612_/A _2621_/Q _1656_/A vssd1 vssd1 vccd1 vccd1 _2230_/X sky130_fd_sc_hd__a21o_4
XFILLER_2_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2092_ _2092_/A _2091_/Y vssd1 vssd1 vccd1 vccd1 _2468_/D sky130_fd_sc_hd__nor2_4
X_2161_ _1256_/Y _2148_/X _1856_/C _1856_/A vssd1 vssd1 vccd1 vccd1 _2161_/Y sky130_fd_sc_hd__a2bb2oi_4
XFILLER_9_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1945_ _1963_/A _1944_/Y vssd1 vssd1 vccd1 vccd1 _2517_/D sky130_fd_sc_hd__nor2_4
X_1876_ _1878_/A DATA_FROM_HASH[4] vssd1 vssd1 vccd1 vccd1 _2563_/D sky130_fd_sc_hd__and2_4
X_2359_ EXT_RESET_N_fromHost vssd1 vssd1 vccd1 vccd1 EXT_RESET_N_toClient sky130_fd_sc_hd__buf_2
X_2428_ _2404_/CLK _2259_/Y vssd1 vssd1 vccd1 vccd1 _2428_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_44_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_3_0_addressalyzerBlock.SPI_CLK clkbuf_4_3_0_addressalyzerBlock.SPI_CLK/A
+ vssd1 vssd1 vccd1 vccd1 _2604_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_12_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1661_ _1383_/C _1661_/B _1661_/C _1661_/D vssd1 vssd1 vccd1 vccd1 _1661_/X sky130_fd_sc_hd__or4_4
X_1730_ _1687_/A _1434_/Y _1728_/Y _1729_/Y vssd1 vssd1 vccd1 vccd1 _1730_/X sky130_fd_sc_hd__a211o_4
X_1592_ _1589_/A _1664_/A vssd1 vssd1 vccd1 vccd1 _1648_/A sky130_fd_sc_hd__nor2_4
XFILLER_7_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2213_ _2544_/Q _1739_/B _2212_/Y _2168_/Y vssd1 vssd1 vccd1 vccd1 _2213_/Y sky130_fd_sc_hd__a22oi_4
X_2144_ _2144_/A vssd1 vssd1 vccd1 vccd1 _2144_/Y sky130_fd_sc_hd__inv_2
X_2075_ _2075_/A vssd1 vssd1 vccd1 vccd1 _2476_/D sky130_fd_sc_hd__inv_2
XFILLER_38_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1859_ _1612_/X _1857_/Y _1858_/Y vssd1 vssd1 vccd1 vccd1 _1859_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_30_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1928_ _1928_/A _1927_/Y vssd1 vssd1 vccd1 vccd1 _2528_/D sky130_fd_sc_hd__nor2_4
Xclkbuf_2_2_0_m1_clk_local clkbuf_2_3_0_m1_clk_local/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_5_0_m1_clk_local/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_57_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1713_ _2401_/Q vssd1 vssd1 vccd1 vccd1 _1713_/Y sky130_fd_sc_hd__inv_2
X_1575_ _1729_/B vssd1 vssd1 vccd1 vccd1 _2337_/B sky130_fd_sc_hd__inv_2
X_1644_ _1644_/A vssd1 vssd1 vccd1 vccd1 _1645_/A sky130_fd_sc_hd__buf_2
XFILLER_6_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2127_ _1840_/B _2121_/X _2127_/C vssd1 vssd1 vccd1 vccd1 _2127_/Y sky130_fd_sc_hd__nand3_4
X_2058_ _2477_/Q vssd1 vssd1 vccd1 vccd1 _2058_/X sky130_fd_sc_hd__buf_2
XFILLER_34_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1360_ _1360_/A vssd1 vssd1 vccd1 vccd1 _1360_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1291_ _1246_/Y vssd1 vssd1 vccd1 vccd1 _1308_/A sky130_fd_sc_hd__inv_2
XFILLER_63_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1558_ _1567_/A vssd1 vssd1 vccd1 vccd1 _1604_/A sky130_fd_sc_hd__inv_2
X_1489_ _1487_/Y _1488_/X _1450_/X vssd1 vssd1 vccd1 vccd1 _1489_/X sky130_fd_sc_hd__a21o_4
X_1627_ _1622_/Y _1624_/X _1626_/Y vssd1 vssd1 vccd1 vccd1 _1627_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_54_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_5_0_m1_clk_local clkbuf_3_2_0_m1_clk_local/X vssd1 vssd1 vccd1 vccd1 _2521_/CLK
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_52_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2530_ _2519_/CLK _2530_/D vssd1 vssd1 vccd1 vccd1 _2530_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_13_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1412_ _1411_/X _2010_/B _1363_/C vssd1 vssd1 vccd1 vccd1 _1412_/X sky130_fd_sc_hd__and3_4
X_2392_ _2646_/CLK _2392_/D vssd1 vssd1 vccd1 vccd1 _2322_/B sky130_fd_sc_hd__dfxtp_4
X_1343_ _1335_/D _1333_/Y _1342_/Y vssd1 vssd1 vccd1 vccd1 _1343_/X sky130_fd_sc_hd__o21a_4
XFILLER_5_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2461_ _2611_/CLK _2461_/D vssd1 vssd1 vccd1 vccd1 _2461_/Q sky130_fd_sc_hd__dfxtp_4
X_1274_ _2364_/D vssd1 vssd1 vccd1 vccd1 _1274_/X sky130_fd_sc_hd__buf_2
XFILLER_36_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1892_ _2096_/A vssd1 vssd1 vccd1 vccd1 _1895_/A sky130_fd_sc_hd__buf_2
X_1961_ _1963_/A _1961_/B vssd1 vssd1 vccd1 vccd1 _1961_/Y sky130_fd_sc_hd__nor2_4
XFILLER_21_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2513_ _2513_/CLK _1952_/X vssd1 vssd1 vccd1 vccd1 DATA_TO_HASH[6] sky130_fd_sc_hd__dfxtp_4
X_2375_ _2374_/CLK _2375_/D vssd1 vssd1 vccd1 vccd1 _2376_/D sky130_fd_sc_hd__dfxtp_4
X_1326_ _1316_/B _1323_/Y _1325_/Y vssd1 vssd1 vccd1 vccd1 _1326_/Y sky130_fd_sc_hd__o21ai_4
X_2444_ _2604_/CLK _2444_/D vssd1 vssd1 vccd1 vccd1 _2131_/C sky130_fd_sc_hd__dfxtp_4
X_1188_ _1188_/A vssd1 vssd1 vccd1 vccd1 _1188_/X sky130_fd_sc_hd__buf_2
X_1257_ _1227_/Y vssd1 vssd1 vccd1 vccd1 _1265_/A sky130_fd_sc_hd__buf_2
XPHY_208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_0 DATA_AVAILABLE[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2160_ _2157_/X _2159_/X _1701_/A vssd1 vssd1 vccd1 vccd1 _2160_/Y sky130_fd_sc_hd__a21oi_4
X_2091_ _2091_/A vssd1 vssd1 vccd1 vccd1 _2091_/Y sky130_fd_sc_hd__inv_2
X_1875_ _1878_/A DATA_FROM_HASH[5] vssd1 vssd1 vccd1 vccd1 _2564_/D sky130_fd_sc_hd__and2_4
XFILLER_14_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1944_ _2421_/Q vssd1 vssd1 vccd1 vccd1 _1944_/Y sky130_fd_sc_hd__inv_2
X_2427_ _2404_/CLK _2427_/D vssd1 vssd1 vccd1 vccd1 _1913_/A sky130_fd_sc_hd__dfxtp_4
X_1309_ _1307_/X _1308_/Y vssd1 vssd1 vccd1 vccd1 _1309_/Y sky130_fd_sc_hd__nand2_4
XFILLER_29_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2289_ _1219_/X _1579_/X _2289_/C _1561_/Y vssd1 vssd1 vccd1 vccd1 _2289_/Y sky130_fd_sc_hd__nor4_4
X_2358_ vssd1 vssd1 vccd1 vccd1 _2358_/HI zero sky130_fd_sc_hd__conb_1
XFILLER_52_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1660_ _1660_/A vssd1 vssd1 vccd1 vccd1 _1661_/D sky130_fd_sc_hd__buf_2
X_1591_ _2597_/Q vssd1 vssd1 vccd1 vccd1 _1664_/A sky130_fd_sc_hd__inv_2
XFILLER_53_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2212_ _2194_/Y _2210_/Y _2211_/Y vssd1 vssd1 vccd1 vccd1 _2212_/Y sky130_fd_sc_hd__o21ai_4
X_2143_ _2142_/Y _2138_/Y _2123_/X _1965_/B _2139_/X vssd1 vssd1 vccd1 vccd1 _2143_/Y
+ sky130_fd_sc_hd__o32ai_4
XFILLER_22_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2074_ _2476_/Q _2072_/Y _2073_/Y vssd1 vssd1 vccd1 vccd1 _2075_/A sky130_fd_sc_hd__a21o_4
X_1858_ _1612_/X _1367_/A _1656_/X vssd1 vssd1 vccd1 vccd1 _1858_/Y sky130_fd_sc_hd__a21oi_4
X_1927_ _2196_/B vssd1 vssd1 vccd1 vccd1 _1927_/Y sky130_fd_sc_hd__inv_2
X_1789_ _1190_/A vssd1 vssd1 vccd1 vccd1 _1789_/X sky130_fd_sc_hd__buf_2
XFILLER_29_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1643_ _1605_/X _1648_/A _1667_/C _1667_/D vssd1 vssd1 vccd1 vccd1 _1644_/A sky130_fd_sc_hd__and4_4
XFILLER_31_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1712_ _1707_/X _1712_/B vssd1 vssd1 vccd1 vccd1 _1712_/Y sky130_fd_sc_hd__nand2_4
X_1574_ _2386_/Q vssd1 vssd1 vccd1 vccd1 _1574_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_4_13_0_m1_clk_local clkbuf_3_6_0_m1_clk_local/X vssd1 vssd1 vccd1 vccd1 _2492_/CLK
+ sky130_fd_sc_hd__clkbuf_1
X_2057_ _2056_/X _2057_/B _2040_/X vssd1 vssd1 vccd1 vccd1 _2057_/X sky130_fd_sc_hd__and3_4
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2126_ _2120_/X _2122_/Y _2125_/Y vssd1 vssd1 vccd1 vccd1 _2446_/D sky130_fd_sc_hd__o21ai_4
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1290_ _1290_/A vssd1 vssd1 vccd1 vccd1 _1290_/Y sky130_fd_sc_hd__inv_2
XFILLER_8_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1626_ _1625_/X _2434_/Q _2448_/Q vssd1 vssd1 vccd1 vccd1 _1626_/Y sky130_fd_sc_hd__a21oi_4
X_1488_ _1488_/A vssd1 vssd1 vccd1 vccd1 _1488_/X sky130_fd_sc_hd__buf_2
X_1557_ _1557_/A _2104_/A _1557_/C vssd1 vssd1 vccd1 vccd1 _1557_/X sky130_fd_sc_hd__and3_4
X_2109_ _2107_/A _2454_/Q vssd1 vssd1 vccd1 vccd1 _2455_/D sky130_fd_sc_hd__and2_4
XFILLER_39_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2460_ _2646_/CLK _2460_/D vssd1 vssd1 vccd1 vccd1 _1833_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_9_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2391_ _2437_/CLK _2332_/X vssd1 vssd1 vccd1 vccd1 _2391_/Q sky130_fd_sc_hd__dfxtp_4
X_1411_ _2615_/Q _1411_/B vssd1 vssd1 vccd1 vccd1 _1411_/X sky130_fd_sc_hd__or2_4
X_1342_ _1335_/D _1353_/A _1329_/X _1321_/X _1339_/X vssd1 vssd1 vccd1 vccd1 _1342_/Y
+ sky130_fd_sc_hd__a41oi_4
X_1273_ _1273_/A vssd1 vssd1 vccd1 vccd1 _1854_/A sky130_fd_sc_hd__inv_2
XFILLER_51_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1609_ _1605_/X _1606_/Y _1667_/C _1667_/D vssd1 vssd1 vccd1 vccd1 _1609_/X sky130_fd_sc_hd__and4_4
X_2589_ _2588_/CLK _2589_/D vssd1 vssd1 vccd1 vccd1 _2589_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_59_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1891_ _1888_/A DATA_AVAILABLE[3] vssd1 vssd1 vccd1 vccd1 _1891_/X sky130_fd_sc_hd__and2_4
XFILLER_41_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1960_ _2442_/Q vssd1 vssd1 vccd1 vccd1 _1961_/B sky130_fd_sc_hd__inv_2
XFILLER_52_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2512_ _2513_/CLK _2512_/D vssd1 vssd1 vccd1 vccd1 DATA_TO_HASH[5] sky130_fd_sc_hd__dfxtp_4
X_2443_ _2604_/CLK _2443_/D vssd1 vssd1 vccd1 vccd1 _2443_/Q sky130_fd_sc_hd__dfxtp_4
X_2374_ _2374_/CLK _2373_/Q vssd1 vssd1 vccd1 vccd1 _2375_/D sky130_fd_sc_hd__dfxtp_4
XFILLER_49_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1325_ _1316_/B _1353_/A _1321_/X _1316_/D _1274_/X vssd1 vssd1 vccd1 vccd1 _1325_/Y
+ sky130_fd_sc_hd__a41oi_4
X_1256_ _1256_/A vssd1 vssd1 vccd1 vccd1 _1256_/Y sky130_fd_sc_hd__inv_2
XFILLER_64_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1187_ _1187_/A vssd1 vssd1 vccd1 vccd1 _1187_/X sky130_fd_sc_hd__buf_2
XFILLER_24_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XINSDIODE2_1 SCLK_fromHost vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_4_8_0_addressalyzerBlock.SPI_CLK clkbuf_4_9_0_addressalyzerBlock.SPI_CLK/A
+ vssd1 vssd1 vccd1 vccd1 _2399_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_47_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2090_ _1284_/X _2089_/Y vssd1 vssd1 vccd1 vccd1 _2090_/Y sky130_fd_sc_hd__nor2_4
XFILLER_61_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1874_ _1886_/A vssd1 vssd1 vccd1 vccd1 _1878_/A sky130_fd_sc_hd__buf_2
XFILLER_14_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1943_ _1339_/X vssd1 vssd1 vccd1 vccd1 _1963_/A sky130_fd_sc_hd__buf_2
X_2426_ _2446_/CLK _2426_/D vssd1 vssd1 vccd1 vccd1 _1622_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_44_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1239_ _1351_/B _1238_/Y vssd1 vssd1 vccd1 vccd1 _1239_/Y sky130_fd_sc_hd__nor2_4
XFILLER_37_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1308_ _1308_/A _2636_/Q _1308_/C vssd1 vssd1 vccd1 vccd1 _1308_/Y sky130_fd_sc_hd__nand3_4
XFILLER_29_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2288_ _1581_/X _2260_/Y _2277_/Y _1929_/Y _2279_/X vssd1 vssd1 vccd1 vccd1 _2411_/D
+ sky130_fd_sc_hd__o32ai_4
X_2357_ vssd1 vssd1 vccd1 vccd1 one _2357_/LO sky130_fd_sc_hd__conb_1
XFILLER_20_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1590_ _1567_/C _1589_/Y vssd1 vssd1 vccd1 vccd1 _1590_/Y sky130_fd_sc_hd__nor2_4
XFILLER_59_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2073_ _2476_/Q _2072_/Y _1374_/X vssd1 vssd1 vccd1 vccd1 _2073_/Y sky130_fd_sc_hd__o21ai_4
X_2211_ _1666_/A THREAD_COUNT[1] vssd1 vssd1 vccd1 vccd1 _2211_/Y sky130_fd_sc_hd__nand2_4
X_2142_ _1514_/A vssd1 vssd1 vccd1 vccd1 _2142_/Y sky130_fd_sc_hd__inv_2
XFILLER_15_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1857_ _1855_/Y _1646_/X _1856_/X vssd1 vssd1 vccd1 vccd1 _1857_/Y sky130_fd_sc_hd__a21oi_4
X_1926_ _1928_/A _1926_/B vssd1 vssd1 vccd1 vccd1 _2529_/D sky130_fd_sc_hd__nor2_4
X_1788_ _2591_/Q vssd1 vssd1 vccd1 vccd1 _1788_/X sky130_fd_sc_hd__buf_2
X_2409_ _2446_/CLK _2296_/Y vssd1 vssd1 vccd1 vccd1 _2295_/C sky130_fd_sc_hd__dfxtp_4
XFILLER_29_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1642_ _1615_/Y _1639_/Y _1641_/X vssd1 vssd1 vccd1 vccd1 _1642_/Y sky130_fd_sc_hd__o21ai_4
X_1711_ _2425_/Q _2181_/A _1708_/X _1710_/Y vssd1 vssd1 vccd1 vccd1 _1712_/B sky130_fd_sc_hd__a211o_4
X_1573_ _1564_/X _1572_/Y _1454_/X vssd1 vssd1 vccd1 vccd1 _1573_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_66_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2056_ _2053_/Y _2062_/B _2055_/X _1993_/C _2481_/Q vssd1 vssd1 vccd1 vccd1 _2056_/X
+ sky130_fd_sc_hd__a41o_4
XFILLER_26_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2125_ _2123_/X _2335_/A _2125_/C vssd1 vssd1 vccd1 vccd1 _2125_/Y sky130_fd_sc_hd__nand3_4
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1909_ _1911_/A _1908_/Y vssd1 vssd1 vccd1 vccd1 _2539_/D sky130_fd_sc_hd__nor2_4
XFILLER_57_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1556_ _1556_/A _1556_/B vssd1 vssd1 vccd1 vccd1 _1557_/C sky130_fd_sc_hd__nand2_4
XFILLER_8_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1625_ _1623_/Y vssd1 vssd1 vccd1 vccd1 _1625_/X sky130_fd_sc_hd__buf_2
XFILLER_39_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1487_ _1487_/A _1487_/B _1504_/A _1486_/X vssd1 vssd1 vccd1 vccd1 _1487_/Y sky130_fd_sc_hd__nand4_4
X_2108_ _2107_/A SCLK_fromHost vssd1 vssd1 vccd1 vccd1 _2456_/D sky130_fd_sc_hd__and2_4
X_2039_ _2039_/A vssd1 vssd1 vccd1 vccd1 _2039_/Y sky130_fd_sc_hd__inv_2
XFILLER_52_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1410_ _1409_/Y vssd1 vssd1 vccd1 vccd1 _1411_/B sky130_fd_sc_hd__inv_2
XFILLER_42_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2390_ _2588_/CLK _2331_/Y vssd1 vssd1 vccd1 vccd1 _2390_/Q sky130_fd_sc_hd__dfxtp_4
X_1341_ _1335_/C _1338_/X _1340_/Y vssd1 vssd1 vccd1 vccd1 _2631_/D sky130_fd_sc_hd__o21a_4
X_1272_ _2641_/Q _1265_/Y _1256_/A _1224_/A vssd1 vssd1 vccd1 vccd1 _1272_/Y sky130_fd_sc_hd__nand4_4
XFILLER_36_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2588_ _2588_/CLK _2588_/D vssd1 vssd1 vccd1 vccd1 _2349_/A sky130_fd_sc_hd__dfxtp_4
X_1608_ _1467_/A _1424_/A vssd1 vssd1 vccd1 vccd1 _1667_/D sky130_fd_sc_hd__nor2_4
X_1539_ _1466_/A _1482_/Y _1538_/X vssd1 vssd1 vccd1 vccd1 _1539_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_63_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_1_0_m1_clk_local clkbuf_3_0_0_m1_clk_local/X vssd1 vssd1 vccd1 vccd1 _2519_/CLK
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_2_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1890_ _1888_/A _2559_/Q vssd1 vssd1 vccd1 vccd1 _2551_/D sky130_fd_sc_hd__and2_4
X_2511_ _2511_/CLK _1954_/X vssd1 vssd1 vccd1 vccd1 DATA_TO_HASH[4] sky130_fd_sc_hd__dfxtp_4
X_2373_ _2374_/CLK _2373_/D vssd1 vssd1 vccd1 vccd1 _2373_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_45_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2442_ _2604_/CLK _2140_/Y vssd1 vssd1 vccd1 vccd1 _2442_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_4_13_0_addressalyzerBlock.SPI_CLK clkbuf_3_6_0_addressalyzerBlock.SPI_CLK/X
+ vssd1 vssd1 vccd1 vccd1 _2464_/CLK sky130_fd_sc_hd__clkbuf_1
X_1186_ _1188_/A vssd1 vssd1 vccd1 vccd1 _1187_/A sky130_fd_sc_hd__buf_2
X_1324_ _1239_/Y vssd1 vssd1 vccd1 vccd1 _1353_/A sky130_fd_sc_hd__buf_2
X_1255_ _1254_/X vssd1 vssd1 vccd1 vccd1 _1289_/B sky130_fd_sc_hd__buf_2
XFILLER_64_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_2 _2501_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_3_7_0_m1_clk_local clkbuf_3_7_0_m1_clk_local/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_7_0_m1_clk_local/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_7_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1942_ _1938_/A _1942_/B vssd1 vssd1 vccd1 vccd1 _1942_/Y sky130_fd_sc_hd__nor2_4
XFILLER_9_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1873_ _1789_/X vssd1 vssd1 vccd1 vccd1 _1886_/A sky130_fd_sc_hd__buf_2
X_2356_ _2354_/Y _2322_/A _2355_/Y vssd1 vssd1 vccd1 vccd1 _2356_/Y sky130_fd_sc_hd__a21oi_4
X_2425_ _2446_/CLK _2425_/D vssd1 vssd1 vccd1 vccd1 _2425_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_52_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1238_ _2620_/Q _1385_/B _1365_/D _1238_/D vssd1 vssd1 vccd1 vccd1 _1238_/Y sky130_fd_sc_hd__nand4_4
X_1307_ _2636_/Q _1305_/X _1306_/X vssd1 vssd1 vccd1 vccd1 _1307_/X sky130_fd_sc_hd__o21a_4
X_2287_ _1581_/X _2257_/Y _2277_/Y _1927_/Y _2279_/X vssd1 vssd1 vccd1 vccd1 _2412_/D
+ sky130_fd_sc_hd__o32ai_4
XFILLER_20_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2210_ _2207_/Y _2208_/X _2209_/X vssd1 vssd1 vccd1 vccd1 _2210_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_53_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2072_ _2071_/Y _2072_/B vssd1 vssd1 vccd1 vccd1 _2072_/Y sky130_fd_sc_hd__nor2_4
XFILLER_38_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2141_ _1503_/Y _2138_/Y _2123_/X _1963_/B _2139_/X vssd1 vssd1 vccd1 vccd1 _2141_/Y
+ sky130_fd_sc_hd__o32ai_4
XFILLER_61_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1925_ _2174_/B vssd1 vssd1 vccd1 vccd1 _1926_/B sky130_fd_sc_hd__inv_2
X_1856_ _1856_/A _1856_/B _1856_/C vssd1 vssd1 vccd1 vccd1 _1856_/X sky130_fd_sc_hd__and3_4
X_1787_ _1786_/Y vssd1 vssd1 vccd1 vccd1 _1983_/B sky130_fd_sc_hd__buf_2
X_2339_ _1840_/C _2385_/Q _2102_/A _2338_/X vssd1 vssd1 vccd1 vccd1 _2339_/X sky130_fd_sc_hd__a211o_4
X_2408_ _2604_/CLK _2408_/D vssd1 vssd1 vccd1 vccd1 ID_toHost sky130_fd_sc_hd__dfxtp_4
XFILLER_52_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1572_ _1569_/X _1556_/A _1661_/B vssd1 vssd1 vccd1 vccd1 _1572_/Y sky130_fd_sc_hd__o21ai_4
X_1641_ _1641_/A _1854_/B vssd1 vssd1 vccd1 vccd1 _1641_/X sky130_fd_sc_hd__or2_4
X_1710_ _1630_/X _1710_/B vssd1 vssd1 vccd1 vccd1 _1710_/Y sky130_fd_sc_hd__nor2_4
X_2124_ _1555_/A vssd1 vssd1 vccd1 vccd1 _2335_/A sky130_fd_sc_hd__buf_2
X_2055_ _2479_/Q vssd1 vssd1 vccd1 vccd1 _2055_/X sky130_fd_sc_hd__buf_2
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1839_ _1839_/A vssd1 vssd1 vccd1 vccd1 _1840_/C sky130_fd_sc_hd__inv_2
X_1908_ _2177_/B vssd1 vssd1 vccd1 vccd1 _1908_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1624_ _1623_/Y vssd1 vssd1 vccd1 vccd1 _1624_/X sky130_fd_sc_hd__buf_2
X_1555_ _1555_/A vssd1 vssd1 vccd1 vccd1 _2104_/A sky130_fd_sc_hd__buf_2
X_2107_ _2107_/A _2456_/Q vssd1 vssd1 vccd1 vccd1 _2457_/D sky130_fd_sc_hd__and2_4
XFILLER_54_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1486_ _1486_/A vssd1 vssd1 vccd1 vccd1 _1486_/X sky130_fd_sc_hd__buf_2
X_2038_ _2038_/A _2038_/B vssd1 vssd1 vccd1 vccd1 _2039_/A sky130_fd_sc_hd__nand2_4
XFILLER_10_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1340_ _1335_/C _1318_/B _1335_/D _1329_/X _1339_/X vssd1 vssd1 vccd1 vccd1 _1340_/Y
+ sky130_fd_sc_hd__a41oi_4
X_1271_ _1271_/A _2010_/B _1252_/A vssd1 vssd1 vccd1 vccd1 _1271_/X sky130_fd_sc_hd__and3_4
X_1538_ _1469_/A _1467_/Y _1556_/B _1548_/D _1488_/X vssd1 vssd1 vccd1 vccd1 _1538_/X
+ sky130_fd_sc_hd__o41a_4
X_1469_ _1469_/A _1467_/Y _1424_/Y _1548_/D vssd1 vssd1 vccd1 vccd1 _1469_/Y sky130_fd_sc_hd__nor4_4
X_2587_ _2399_/CLK _1792_/X vssd1 vssd1 vccd1 vccd1 _1420_/A sky130_fd_sc_hd__dfxtp_4
X_1607_ _2604_/Q _1483_/D vssd1 vssd1 vccd1 vccd1 _1667_/C sky130_fd_sc_hd__nor2_4
XFILLER_63_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2510_ _2505_/CLK _2510_/D vssd1 vssd1 vccd1 vccd1 DATA_TO_HASH[3] sky130_fd_sc_hd__dfxtp_4
X_2372_ _2374_/CLK _2372_/D vssd1 vssd1 vccd1 vccd1 _2373_/D sky130_fd_sc_hd__dfxtp_4
X_1323_ _1322_/Y vssd1 vssd1 vccd1 vccd1 _1323_/Y sky130_fd_sc_hd__inv_2
X_2441_ _2552_/CLK _2141_/Y vssd1 vssd1 vccd1 vccd1 _2441_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_64_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1185_ _1185_/A vssd1 vssd1 vccd1 vccd1 _1188_/A sky130_fd_sc_hd__inv_2
X_1254_ _1269_/A vssd1 vssd1 vccd1 vccd1 _1254_/X sky130_fd_sc_hd__buf_2
XFILLER_64_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2639_ _2632_/CLK _1290_/Y vssd1 vssd1 vccd1 vccd1 _1224_/A sky130_fd_sc_hd__dfxtp_4
XINSDIODE2_3 _1920_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1872_ _2112_/A DATA_FROM_HASH[6] vssd1 vssd1 vccd1 vccd1 _2565_/D sky130_fd_sc_hd__and2_4
XFILLER_0_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1941_ _2155_/A vssd1 vssd1 vccd1 vccd1 _1942_/B sky130_fd_sc_hd__inv_2
XFILLER_21_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1306_ _1346_/A vssd1 vssd1 vccd1 vccd1 _1306_/X sky130_fd_sc_hd__buf_2
X_2355_ _1676_/B _1187_/A _1213_/X vssd1 vssd1 vccd1 vccd1 _2355_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_29_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2424_ _2446_/CLK _2269_/Y vssd1 vssd1 vccd1 vccd1 _2424_/Q sky130_fd_sc_hd__dfxtp_4
X_2286_ _1581_/X _2255_/Y _2277_/Y _1926_/B _2279_/X vssd1 vssd1 vccd1 vccd1 _2413_/D
+ sky130_fd_sc_hd__o32ai_4
XFILLER_56_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1237_ _1237_/A vssd1 vssd1 vccd1 vccd1 _1238_/D sky130_fd_sc_hd__inv_2
XFILLER_44_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2140_ _2136_/Y _2138_/Y _2120_/X _1961_/B _2139_/X vssd1 vssd1 vccd1 vccd1 _2140_/Y
+ sky130_fd_sc_hd__o32ai_4
X_2071_ _2071_/A vssd1 vssd1 vccd1 vccd1 _2071_/Y sky130_fd_sc_hd__inv_2
XFILLER_46_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1855_ _1843_/Y _1853_/Y _1854_/X vssd1 vssd1 vccd1 vccd1 _1855_/Y sky130_fd_sc_hd__o21ai_4
X_1924_ _1928_/A _1924_/B vssd1 vssd1 vccd1 vccd1 _2530_/D sky130_fd_sc_hd__nor2_4
X_1786_ _2591_/Q vssd1 vssd1 vccd1 vccd1 _1786_/Y sky130_fd_sc_hd__inv_2
X_2338_ _2338_/A _1188_/A _2462_/Q vssd1 vssd1 vccd1 vccd1 _2338_/X sky130_fd_sc_hd__and3_4
XFILLER_37_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2269_ _2268_/Y _2262_/X _2258_/X _1847_/Y _2264_/X vssd1 vssd1 vccd1 vccd1 _2269_/Y
+ sky130_fd_sc_hd__o32ai_4
X_2407_ _2604_/CLK _2407_/D vssd1 vssd1 vccd1 vccd1 _2407_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_37_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1571_ _1571_/A vssd1 vssd1 vccd1 vccd1 _1661_/B sky130_fd_sc_hd__buf_2
X_1640_ _1613_/Y vssd1 vssd1 vccd1 vccd1 _1854_/B sky130_fd_sc_hd__buf_2
XFILLER_6_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2123_ _2120_/A vssd1 vssd1 vccd1 vccd1 _2123_/X sky130_fd_sc_hd__buf_2
XFILLER_20_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2054_ _2054_/A vssd1 vssd1 vccd1 vccd1 _2062_/B sky130_fd_sc_hd__buf_2
X_1838_ _1789_/X vssd1 vssd1 vccd1 vccd1 _1840_/B sky130_fd_sc_hd__buf_2
X_1907_ _1911_/A _1906_/Y vssd1 vssd1 vccd1 vccd1 _1907_/Y sky130_fd_sc_hd__nor2_4
XFILLER_66_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1769_ _1486_/A _1764_/Y _1766_/Y _1767_/X _1768_/X vssd1 vssd1 vccd1 vccd1 _1770_/A
+ sky130_fd_sc_hd__a2111o_4
XFILLER_40_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1554_ _1190_/A vssd1 vssd1 vccd1 vccd1 _1555_/A sky130_fd_sc_hd__buf_2
X_1623_ _2447_/Q vssd1 vssd1 vccd1 vccd1 _1623_/Y sky130_fd_sc_hd__inv_2
X_1485_ _2607_/Q vssd1 vssd1 vccd1 vccd1 _1504_/A sky130_fd_sc_hd__buf_2
.ends


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO decred_controller
  CLASS BLOCK ;
  FOREIGN decred_controller ;
  ORIGIN 0.000 0.000 ;
  SIZE 205.000 BY 205.000 ;
  PIN CLK_LED
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.730 201.000 62.010 205.000 ;
    END
  END CLK_LED
  PIN DATA_AVAILABLE[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.130 201.000 149.410 205.000 ;
    END
  END DATA_AVAILABLE[0]
  PIN DATA_AVAILABLE[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.810 201.000 130.090 205.000 ;
    END
  END DATA_AVAILABLE[1]
  PIN DATA_AVAILABLE[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 145.560 4.000 146.160 ;
    END
  END DATA_AVAILABLE[2]
  PIN DATA_AVAILABLE[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 201.000 193.160 205.000 193.760 ;
    END
  END DATA_AVAILABLE[3]
  PIN DATA_AVAILABLE[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.330 0.000 89.610 4.000 ;
    END
  END DATA_AVAILABLE[4]
  PIN DATA_AVAILABLE[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.650 0.000 108.930 4.000 ;
    END
  END DATA_AVAILABLE[5]
  PIN DATA_FROM_HASH[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 187.770 201.000 188.050 205.000 ;
    END
  END DATA_FROM_HASH[0]
  PIN DATA_FROM_HASH[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.850 201.000 72.130 205.000 ;
    END
  END DATA_FROM_HASH[1]
  PIN DATA_FROM_HASH[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 174.120 4.000 174.720 ;
    END
  END DATA_FROM_HASH[2]
  PIN DATA_FROM_HASH[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 201.000 21.800 205.000 22.400 ;
    END
  END DATA_FROM_HASH[3]
  PIN DATA_FROM_HASH[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.690 201.000 119.970 205.000 ;
    END
  END DATA_FROM_HASH[4]
  PIN DATA_FROM_HASH[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.850 0.000 118.130 4.000 ;
    END
  END DATA_FROM_HASH[5]
  PIN DATA_FROM_HASH[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.890 201.000 14.170 205.000 ;
    END
  END DATA_FROM_HASH[6]
  PIN DATA_FROM_HASH[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 201.000 179.560 205.000 180.160 ;
    END
  END DATA_FROM_HASH[7]
  PIN DATA_TO_HASH[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.250 0.000 21.530 4.000 ;
    END
  END DATA_TO_HASH[0]
  PIN DATA_TO_HASH[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 166.610 0.000 166.890 4.000 ;
    END
  END DATA_TO_HASH[1]
  PIN DATA_TO_HASH[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.050 201.000 81.330 205.000 ;
    END
  END DATA_TO_HASH[2]
  PIN DATA_TO_HASH[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.930 0.000 186.210 4.000 ;
    END
  END DATA_TO_HASH[3]
  PIN DATA_TO_HASH[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 201.000 65.320 205.000 65.920 ;
    END
  END DATA_TO_HASH[4]
  PIN DATA_TO_HASH[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.490 0.000 156.770 4.000 ;
    END
  END DATA_TO_HASH[5]
  PIN DATA_TO_HASH[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 158.330 201.000 158.610 205.000 ;
    END
  END DATA_TO_HASH[6]
  PIN DATA_TO_HASH[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.090 201.000 23.370 205.000 ;
    END
  END DATA_TO_HASH[7]
  PIN EXT_RESET_N_fromHost
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.290 0.000 147.570 4.000 ;
    END
  END EXT_RESET_N_fromHost
  PIN EXT_RESET_N_toClient
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.970 201.000 197.250 205.000 ;
    END
  END EXT_RESET_N_toClient
  PIN HASH_ADDR[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.690 0.000 50.970 4.000 ;
    END
  END HASH_ADDR[0]
  PIN HASH_ADDR[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.650 201.000 177.930 205.000 ;
    END
  END HASH_ADDR[1]
  PIN HASH_ADDR[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 117.000 4.000 117.600 ;
    END
  END HASH_ADDR[2]
  PIN HASH_ADDR[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 131.960 4.000 132.560 ;
    END
  END HASH_ADDR[3]
  PIN HASH_ADDR[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.490 201.000 110.770 205.000 ;
    END
  END HASH_ADDR[4]
  PIN HASH_ADDR[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 160.520 4.000 161.120 ;
    END
  END HASH_ADDR[5]
  PIN HASH_EN
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 201.000 36.760 205.000 37.360 ;
    END
  END HASH_EN
  PIN HASH_LED
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 46.280 4.000 46.880 ;
    END
  END HASH_LED
  PIN ID_fromClient
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 201.000 78.920 205.000 79.520 ;
    END
  END ID_fromClient
  PIN ID_toHost
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 103.400 4.000 104.000 ;
    END
  END ID_toHost
  PIN IRQ_OUT_fromClient
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.570 0.000 40.850 4.000 ;
    END
  END IRQ_OUT_fromClient
  PIN IRQ_OUT_toHost
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.370 0.000 31.650 4.000 ;
    END
  END IRQ_OUT_toHost
  PIN M1_CLK_IN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.970 0.000 128.250 4.000 ;
    END
  END M1_CLK_IN
  PIN M1_CLK_SELECT
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.530 0.000 98.810 4.000 ;
    END
  END M1_CLK_SELECT
  PIN MACRO_RD_SELECT[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.210 0.000 79.490 4.000 ;
    END
  END MACRO_RD_SELECT[0]
  PIN MACRO_RD_SELECT[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.890 0.000 60.170 4.000 ;
    END
  END MACRO_RD_SELECT[1]
  PIN MACRO_RD_SELECT[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.170 201.000 91.450 205.000 ;
    END
  END MACRO_RD_SELECT[2]
  PIN MACRO_RD_SELECT[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.050 0.000 12.330 4.000 ;
    END
  END MACRO_RD_SELECT[3]
  PIN MACRO_RD_SELECT[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 201.000 164.600 205.000 165.200 ;
    END
  END MACRO_RD_SELECT[4]
  PIN MACRO_RD_SELECT[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 201.000 8.200 205.000 8.800 ;
    END
  END MACRO_RD_SELECT[5]
  PIN MACRO_WR_SELECT[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.530 201.000 52.810 205.000 ;
    END
  END MACRO_WR_SELECT[0]
  PIN MACRO_WR_SELECT[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 168.450 201.000 168.730 205.000 ;
    END
  END MACRO_WR_SELECT[1]
  PIN MACRO_WR_SELECT[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 201.000 151.000 205.000 151.600 ;
    END
  END MACRO_WR_SELECT[2]
  PIN MACRO_WR_SELECT[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 201.000 50.360 205.000 50.960 ;
    END
  END MACRO_WR_SELECT[3]
  PIN MACRO_WR_SELECT[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 195.130 0.000 195.410 4.000 ;
    END
  END MACRO_WR_SELECT[4]
  PIN MACRO_WR_SELECT[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 189.080 4.000 189.680 ;
    END
  END MACRO_WR_SELECT[5]
  PIN MISO_fromClient
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 201.000 136.040 205.000 136.640 ;
    END
  END MISO_fromClient
  PIN MISO_toHost
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 201.000 122.440 205.000 123.040 ;
    END
  END MISO_toHost
  PIN MOSI_fromHost
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.410 201.000 42.690 205.000 ;
    END
  END MOSI_fromHost
  PIN MOSI_toClient
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.010 201.000 139.290 205.000 ;
    END
  END MOSI_toClient
  PIN PLL_INPUT
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.720 4.000 18.320 ;
    END
  END PLL_INPUT
  PIN S1_CLK_IN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.850 0.000 3.130 4.000 ;
    END
  END S1_CLK_IN
  PIN S1_CLK_SELECT
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 59.880 4.000 60.480 ;
    END
  END S1_CLK_SELECT
  PIN SCLK_fromHost
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.010 0.000 70.290 4.000 ;
    END
  END SCLK_fromHost
  PIN SCLK_toClient
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.440 4.000 89.040 ;
    END
  END SCLK_toClient
  PIN SCSN_fromHost
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 4.000 75.440 ;
    END
  END SCSN_fromHost
  PIN SCSN_toClient
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.170 0.000 137.450 4.000 ;
    END
  END SCSN_toClient
  PIN THREAD_COUNT[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.810 0.000 176.090 4.000 ;
    END
  END THREAD_COUNT[0]
  PIN THREAD_COUNT[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.370 201.000 100.650 205.000 ;
    END
  END THREAD_COUNT[1]
  PIN THREAD_COUNT[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.770 201.000 4.050 205.000 ;
    END
  END THREAD_COUNT[2]
  PIN THREAD_COUNT[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 201.000 93.880 205.000 94.480 ;
    END
  END THREAD_COUNT[3]
  PIN m1_clk_local
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 31.320 4.000 31.920 ;
    END
  END m1_clk_local
  PIN one
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.210 201.000 33.490 205.000 ;
    END
  END one
  PIN zero
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 201.000 107.480 205.000 108.080 ;
    END
  END zero
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 193.360 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 193.360 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 193.360 ;
    END
  END vssd1
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 177.940 10.880 179.540 193.120 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 24.340 10.880 25.940 193.120 ;
    END
  END vccd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 101.140 10.880 102.740 193.120 ;
    END
  END vssd2
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 181.240 10.880 182.840 193.120 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 27.640 10.880 29.240 193.120 ;
    END
  END vdda1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 104.440 10.880 106.040 193.120 ;
    END
  END vssa1
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 184.540 10.880 186.140 193.120 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 30.940 10.880 32.540 193.120 ;
    END
  END vdda2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 107.740 10.880 109.340 193.120 ;
    END
  END vssa2
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 199.955 193.205 ;
      LAYER met1 ;
        RECT 0.070 5.480 200.030 193.360 ;
      LAYER met2 ;
        RECT 0.090 200.720 3.490 201.000 ;
        RECT 4.330 200.720 13.610 201.000 ;
        RECT 14.450 200.720 22.810 201.000 ;
        RECT 23.650 200.720 32.930 201.000 ;
        RECT 33.770 200.720 42.130 201.000 ;
        RECT 42.970 200.720 52.250 201.000 ;
        RECT 53.090 200.720 61.450 201.000 ;
        RECT 62.290 200.720 71.570 201.000 ;
        RECT 72.410 200.720 80.770 201.000 ;
        RECT 81.610 200.720 90.890 201.000 ;
        RECT 91.730 200.720 100.090 201.000 ;
        RECT 100.930 200.720 110.210 201.000 ;
        RECT 111.050 200.720 119.410 201.000 ;
        RECT 120.250 200.720 129.530 201.000 ;
        RECT 130.370 200.720 138.730 201.000 ;
        RECT 139.570 200.720 148.850 201.000 ;
        RECT 149.690 200.720 158.050 201.000 ;
        RECT 158.890 200.720 168.170 201.000 ;
        RECT 169.010 200.720 177.370 201.000 ;
        RECT 178.210 200.720 187.490 201.000 ;
        RECT 188.330 200.720 196.690 201.000 ;
        RECT 197.530 200.720 200.010 201.000 ;
        RECT 0.090 4.280 200.010 200.720 ;
        RECT 0.090 4.000 2.570 4.280 ;
        RECT 3.410 4.000 11.770 4.280 ;
        RECT 12.610 4.000 20.970 4.280 ;
        RECT 21.810 4.000 31.090 4.280 ;
        RECT 31.930 4.000 40.290 4.280 ;
        RECT 41.130 4.000 50.410 4.280 ;
        RECT 51.250 4.000 59.610 4.280 ;
        RECT 60.450 4.000 69.730 4.280 ;
        RECT 70.570 4.000 78.930 4.280 ;
        RECT 79.770 4.000 89.050 4.280 ;
        RECT 89.890 4.000 98.250 4.280 ;
        RECT 99.090 4.000 108.370 4.280 ;
        RECT 109.210 4.000 117.570 4.280 ;
        RECT 118.410 4.000 127.690 4.280 ;
        RECT 128.530 4.000 136.890 4.280 ;
        RECT 137.730 4.000 147.010 4.280 ;
        RECT 147.850 4.000 156.210 4.280 ;
        RECT 157.050 4.000 166.330 4.280 ;
        RECT 167.170 4.000 175.530 4.280 ;
        RECT 176.370 4.000 185.650 4.280 ;
        RECT 186.490 4.000 194.850 4.280 ;
        RECT 195.690 4.000 200.010 4.280 ;
      LAYER met3 ;
        RECT 0.065 192.760 200.600 193.625 ;
        RECT 0.065 190.080 201.000 192.760 ;
        RECT 4.400 188.680 201.000 190.080 ;
        RECT 0.065 180.560 201.000 188.680 ;
        RECT 0.065 179.160 200.600 180.560 ;
        RECT 0.065 175.120 201.000 179.160 ;
        RECT 4.400 173.720 201.000 175.120 ;
        RECT 0.065 165.600 201.000 173.720 ;
        RECT 0.065 164.200 200.600 165.600 ;
        RECT 0.065 161.520 201.000 164.200 ;
        RECT 4.400 160.120 201.000 161.520 ;
        RECT 0.065 152.000 201.000 160.120 ;
        RECT 0.065 150.600 200.600 152.000 ;
        RECT 0.065 146.560 201.000 150.600 ;
        RECT 4.400 145.160 201.000 146.560 ;
        RECT 0.065 137.040 201.000 145.160 ;
        RECT 0.065 135.640 200.600 137.040 ;
        RECT 0.065 132.960 201.000 135.640 ;
        RECT 4.400 131.560 201.000 132.960 ;
        RECT 0.065 123.440 201.000 131.560 ;
        RECT 0.065 122.040 200.600 123.440 ;
        RECT 0.065 118.000 201.000 122.040 ;
        RECT 4.400 116.600 201.000 118.000 ;
        RECT 0.065 108.480 201.000 116.600 ;
        RECT 0.065 107.080 200.600 108.480 ;
        RECT 0.065 104.400 201.000 107.080 ;
        RECT 4.400 103.000 201.000 104.400 ;
        RECT 0.065 94.880 201.000 103.000 ;
        RECT 0.065 93.480 200.600 94.880 ;
        RECT 0.065 89.440 201.000 93.480 ;
        RECT 4.400 88.040 201.000 89.440 ;
        RECT 0.065 79.920 201.000 88.040 ;
        RECT 0.065 78.520 200.600 79.920 ;
        RECT 0.065 75.840 201.000 78.520 ;
        RECT 4.400 74.440 201.000 75.840 ;
        RECT 0.065 66.320 201.000 74.440 ;
        RECT 0.065 64.920 200.600 66.320 ;
        RECT 0.065 60.880 201.000 64.920 ;
        RECT 4.400 59.480 201.000 60.880 ;
        RECT 0.065 51.360 201.000 59.480 ;
        RECT 0.065 49.960 200.600 51.360 ;
        RECT 0.065 47.280 201.000 49.960 ;
        RECT 4.400 45.880 201.000 47.280 ;
        RECT 0.065 37.760 201.000 45.880 ;
        RECT 0.065 36.360 200.600 37.760 ;
        RECT 0.065 32.320 201.000 36.360 ;
        RECT 4.400 30.920 201.000 32.320 ;
        RECT 0.065 22.800 201.000 30.920 ;
        RECT 0.065 21.400 200.600 22.800 ;
        RECT 0.065 18.720 201.000 21.400 ;
        RECT 4.400 17.320 201.000 18.720 ;
        RECT 0.065 9.200 201.000 17.320 ;
        RECT 0.065 8.335 200.600 9.200 ;
      LAYER met4 ;
        RECT 96.895 17.855 97.440 160.305 ;
        RECT 99.840 17.855 100.740 160.305 ;
        RECT 103.140 17.855 104.040 160.305 ;
        RECT 106.440 17.855 107.340 160.305 ;
        RECT 109.740 17.855 174.240 160.305 ;
        RECT 176.640 17.855 177.540 160.305 ;
        RECT 179.940 17.855 180.840 160.305 ;
        RECT 183.240 17.855 184.140 160.305 ;
        RECT 186.540 17.855 189.225 160.305 ;
  END
END decred_controller
END LIBRARY


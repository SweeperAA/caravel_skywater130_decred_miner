magic
tech sky130A
magscale 1 2
timestamp 1608308602
<< locali >>
rect 24593 37179 24627 37417
rect 6101 36227 6135 36329
rect 6653 34527 6687 34629
rect 28089 32283 28123 32453
rect 19533 20791 19567 20893
rect 4077 19907 4111 20009
rect 14013 18683 14047 18785
rect 20729 12087 20763 12393
rect 32781 11679 32815 11781
rect 34897 8347 34931 8585
rect 9505 7735 9539 8041
rect 15761 6103 15795 6205
rect 12817 5015 12851 5253
rect 9781 2975 9815 3077
<< viali >>
rect 24593 37417 24627 37451
rect 4997 37349 5031 37383
rect 9229 37349 9263 37383
rect 4261 37281 4295 37315
rect 4905 37281 4939 37315
rect 5549 37281 5583 37315
rect 7573 37281 7607 37315
rect 7849 37281 7883 37315
rect 9781 37281 9815 37315
rect 11713 37281 11747 37315
rect 15485 37213 15519 37247
rect 15761 37213 15795 37247
rect 31677 37349 31711 37383
rect 34437 37349 34471 37383
rect 24685 37281 24719 37315
rect 24961 37281 24995 37315
rect 29837 37281 29871 37315
rect 30297 37281 30331 37315
rect 33701 37281 33735 37315
rect 34161 37281 34195 37315
rect 35909 37281 35943 37315
rect 36277 37281 36311 37315
rect 36921 37281 36955 37315
rect 37105 37281 37139 37315
rect 37197 37281 37231 37315
rect 30021 37213 30055 37247
rect 36369 37213 36403 37247
rect 24593 37145 24627 37179
rect 35725 37145 35759 37179
rect 4353 37077 4387 37111
rect 5733 37077 5767 37111
rect 9873 37077 9907 37111
rect 11805 37077 11839 37111
rect 16865 37077 16899 37111
rect 26249 37077 26283 37111
rect 37381 37077 37415 37111
rect 2697 36873 2731 36907
rect 35265 36873 35299 36907
rect 2421 36805 2455 36839
rect 7021 36805 7055 36839
rect 13829 36805 13863 36839
rect 15025 36805 15059 36839
rect 37381 36805 37415 36839
rect 16037 36737 16071 36771
rect 30573 36737 30607 36771
rect 32689 36737 32723 36771
rect 36277 36737 36311 36771
rect 1777 36669 1811 36703
rect 2513 36669 2547 36703
rect 3341 36669 3375 36703
rect 3985 36669 4019 36703
rect 4261 36669 4295 36703
rect 6101 36669 6135 36703
rect 6837 36669 6871 36703
rect 8677 36669 8711 36703
rect 8953 36669 8987 36703
rect 11069 36669 11103 36703
rect 11713 36669 11747 36703
rect 12449 36669 12483 36703
rect 12725 36669 12759 36703
rect 14933 36669 14967 36703
rect 15761 36669 15795 36703
rect 18061 36669 18095 36703
rect 18337 36669 18371 36703
rect 20545 36669 20579 36703
rect 21281 36669 21315 36703
rect 21557 36669 21591 36703
rect 23673 36669 23707 36703
rect 23949 36669 23983 36703
rect 26893 36669 26927 36703
rect 27169 36669 27203 36703
rect 29561 36669 29595 36703
rect 29745 36669 29779 36703
rect 30849 36669 30883 36703
rect 32965 36669 32999 36703
rect 35173 36669 35207 36703
rect 36001 36669 36035 36703
rect 3433 36601 3467 36635
rect 5641 36601 5675 36635
rect 22937 36601 22971 36635
rect 28549 36601 28583 36635
rect 32229 36601 32263 36635
rect 34989 36601 35023 36635
rect 1961 36533 1995 36567
rect 6193 36533 6227 36567
rect 10057 36533 10091 36567
rect 11161 36533 11195 36567
rect 11805 36533 11839 36567
rect 17141 36533 17175 36567
rect 19441 36533 19475 36567
rect 20637 36533 20671 36567
rect 25053 36533 25087 36567
rect 29377 36533 29411 36567
rect 34253 36533 34287 36567
rect 6101 36329 6135 36363
rect 7665 36329 7699 36363
rect 22293 36329 22327 36363
rect 24409 36329 24443 36363
rect 27905 36329 27939 36363
rect 18521 36261 18555 36295
rect 37197 36261 37231 36295
rect 2697 36193 2731 36227
rect 3157 36193 3191 36227
rect 4353 36193 4387 36227
rect 4629 36193 4663 36227
rect 4813 36193 4847 36227
rect 6101 36193 6135 36227
rect 6285 36193 6319 36227
rect 8401 36193 8435 36227
rect 9965 36193 9999 36227
rect 10149 36193 10183 36227
rect 10425 36193 10459 36227
rect 11345 36193 11379 36227
rect 12265 36193 12299 36227
rect 14105 36193 14139 36227
rect 15485 36193 15519 36227
rect 15577 36193 15611 36227
rect 16865 36193 16899 36227
rect 19441 36193 19475 36227
rect 19717 36193 19751 36227
rect 20085 36193 20119 36227
rect 21189 36193 21223 36227
rect 23305 36193 23339 36227
rect 26801 36193 26835 36227
rect 28917 36193 28951 36227
rect 31125 36193 31159 36227
rect 32873 36193 32907 36227
rect 33425 36193 33459 36227
rect 35081 36193 35115 36227
rect 35357 36193 35391 36227
rect 35541 36193 35575 36227
rect 36001 36193 36035 36227
rect 36645 36193 36679 36227
rect 36737 36193 36771 36227
rect 37749 36193 37783 36227
rect 2421 36125 2455 36159
rect 4169 36125 4203 36159
rect 6561 36125 6595 36159
rect 9781 36125 9815 36159
rect 11989 36125 12023 36159
rect 13645 36125 13679 36159
rect 17141 36125 17175 36159
rect 20913 36125 20947 36159
rect 23029 36125 23063 36159
rect 26525 36125 26559 36159
rect 28641 36125 28675 36159
rect 33517 36125 33551 36159
rect 36461 36125 36495 36159
rect 3065 36057 3099 36091
rect 33425 36057 33459 36091
rect 8493 35989 8527 36023
rect 11437 35989 11471 36023
rect 14197 35989 14231 36023
rect 15301 35989 15335 36023
rect 15761 35989 15795 36023
rect 20361 35989 20395 36023
rect 30021 35989 30055 36023
rect 31217 35989 31251 36023
rect 37841 35989 37875 36023
rect 20821 35785 20855 35819
rect 21373 35785 21407 35819
rect 25329 35785 25363 35819
rect 27629 35785 27663 35819
rect 28917 35785 28951 35819
rect 32965 35785 32999 35819
rect 34989 35717 35023 35751
rect 2145 35649 2179 35683
rect 5733 35649 5767 35683
rect 9413 35649 9447 35683
rect 11161 35649 11195 35683
rect 14565 35649 14599 35683
rect 16405 35649 16439 35683
rect 19533 35649 19567 35683
rect 23949 35649 23983 35683
rect 24225 35649 24259 35683
rect 26065 35649 26099 35683
rect 29285 35649 29319 35683
rect 29561 35649 29595 35683
rect 35725 35649 35759 35683
rect 36461 35649 36495 35683
rect 36737 35649 36771 35683
rect 2421 35581 2455 35615
rect 5089 35581 5123 35615
rect 5641 35581 5675 35615
rect 6929 35581 6963 35615
rect 7297 35581 7331 35615
rect 7849 35581 7883 35615
rect 8033 35581 8067 35615
rect 9321 35581 9355 35615
rect 9781 35581 9815 35615
rect 10241 35581 10275 35615
rect 10885 35581 10919 35615
rect 11069 35581 11103 35615
rect 11529 35581 11563 35615
rect 12449 35581 12483 35615
rect 12541 35581 12575 35615
rect 13093 35581 13127 35615
rect 13553 35581 13587 35615
rect 14289 35581 14323 35615
rect 16497 35581 16531 35615
rect 18245 35581 18279 35615
rect 18337 35581 18371 35615
rect 19257 35581 19291 35615
rect 21557 35581 21591 35615
rect 22109 35581 22143 35615
rect 22201 35581 22235 35615
rect 26341 35581 26375 35615
rect 29101 35581 29135 35615
rect 31401 35581 31435 35615
rect 31677 35581 31711 35615
rect 33885 35581 33919 35615
rect 34161 35581 34195 35615
rect 34345 35581 34379 35615
rect 34897 35581 34931 35615
rect 35633 35581 35667 35615
rect 3801 35513 3835 35547
rect 13829 35513 13863 35547
rect 16957 35513 16991 35547
rect 18797 35513 18831 35547
rect 22661 35513 22695 35547
rect 4905 35445 4939 35479
rect 8033 35445 8067 35479
rect 15669 35445 15703 35479
rect 30665 35445 30699 35479
rect 31217 35445 31251 35479
rect 37841 35445 37875 35479
rect 2237 35241 2271 35275
rect 8677 35241 8711 35275
rect 20361 35241 20395 35275
rect 22109 35241 22143 35275
rect 25513 35241 25547 35275
rect 28641 35241 28675 35275
rect 33793 35241 33827 35275
rect 14105 35173 14139 35207
rect 1409 35105 1443 35139
rect 2329 35105 2363 35139
rect 2881 35105 2915 35139
rect 4629 35105 4663 35139
rect 4997 35105 5031 35139
rect 5917 35105 5951 35139
rect 6469 35105 6503 35139
rect 7297 35105 7331 35139
rect 9689 35105 9723 35139
rect 10701 35105 10735 35139
rect 11069 35105 11103 35139
rect 11437 35105 11471 35139
rect 13185 35105 13219 35139
rect 13277 35105 13311 35139
rect 13829 35105 13863 35139
rect 14197 35105 14231 35139
rect 16129 35105 16163 35139
rect 17233 35105 17267 35139
rect 19441 35105 19475 35139
rect 20545 35105 20579 35139
rect 21005 35105 21039 35139
rect 22293 35105 22327 35139
rect 22661 35105 22695 35139
rect 24041 35105 24075 35139
rect 24593 35105 24627 35139
rect 25697 35105 25731 35139
rect 26801 35105 26835 35139
rect 28825 35105 28859 35139
rect 29377 35105 29411 35139
rect 29929 35105 29963 35139
rect 30205 35105 30239 35139
rect 30941 35105 30975 35139
rect 31125 35105 31159 35139
rect 32505 35105 32539 35139
rect 34345 35105 34379 35139
rect 35173 35105 35207 35139
rect 35357 35105 35391 35139
rect 36093 35105 36127 35139
rect 36461 35105 36495 35139
rect 3157 35037 3191 35071
rect 4261 35037 4295 35071
rect 6653 35037 6687 35071
rect 7573 35037 7607 35071
rect 11713 35037 11747 35071
rect 15301 35037 15335 35071
rect 15853 35037 15887 35071
rect 16313 35037 16347 35071
rect 17509 35037 17543 35071
rect 19349 35037 19383 35071
rect 20913 35037 20947 35071
rect 22385 35037 22419 35071
rect 24501 35037 24535 35071
rect 26525 35037 26559 35071
rect 31033 35037 31067 35071
rect 31585 35037 31619 35071
rect 32229 35037 32263 35071
rect 36277 35037 36311 35071
rect 4905 34969 4939 35003
rect 29285 34969 29319 35003
rect 30757 34969 30791 35003
rect 1593 34901 1627 34935
rect 9873 34901 9907 34935
rect 18797 34901 18831 34935
rect 19625 34901 19659 34935
rect 21189 34901 21223 34935
rect 24777 34901 24811 34935
rect 27905 34901 27939 34935
rect 35449 34901 35483 34935
rect 15209 34697 15243 34731
rect 17417 34697 17451 34731
rect 32781 34697 32815 34731
rect 6653 34629 6687 34663
rect 12633 34629 12667 34663
rect 18153 34629 18187 34663
rect 33701 34629 33735 34663
rect 1409 34561 1443 34595
rect 2145 34561 2179 34595
rect 4721 34561 4755 34595
rect 7941 34561 7975 34595
rect 9413 34561 9447 34595
rect 10333 34561 10367 34595
rect 11713 34561 11747 34595
rect 13185 34561 13219 34595
rect 15853 34561 15887 34595
rect 16129 34561 16163 34595
rect 19349 34561 19383 34595
rect 19625 34561 19659 34595
rect 21465 34561 21499 34595
rect 24409 34561 24443 34595
rect 25513 34561 25547 34595
rect 27353 34561 27387 34595
rect 34345 34561 34379 34595
rect 37289 34561 37323 34595
rect 1685 34493 1719 34527
rect 2697 34493 2731 34527
rect 3249 34493 3283 34527
rect 3617 34493 3651 34527
rect 3801 34493 3835 34527
rect 4077 34493 4111 34527
rect 5273 34493 5307 34527
rect 5457 34493 5491 34527
rect 5641 34493 5675 34527
rect 5825 34493 5859 34527
rect 6101 34493 6135 34527
rect 6653 34493 6687 34527
rect 7297 34493 7331 34527
rect 7665 34493 7699 34527
rect 9781 34493 9815 34527
rect 10149 34493 10183 34527
rect 10793 34493 10827 34527
rect 11621 34493 11655 34527
rect 12449 34493 12483 34527
rect 13645 34493 13679 34527
rect 13829 34493 13863 34527
rect 14013 34493 14047 34527
rect 14197 34493 14231 34527
rect 14473 34493 14507 34527
rect 15117 34493 15151 34527
rect 18061 34493 18095 34527
rect 18613 34493 18647 34527
rect 21005 34493 21039 34527
rect 21741 34493 21775 34527
rect 23121 34493 23155 34527
rect 24133 34493 24167 34527
rect 27077 34493 27111 34527
rect 29285 34493 29319 34527
rect 29561 34493 29595 34527
rect 31401 34493 31435 34527
rect 31677 34493 31711 34527
rect 33609 34493 33643 34527
rect 33885 34493 33919 34527
rect 35633 34493 35667 34527
rect 36553 34493 36587 34527
rect 1593 34425 1627 34459
rect 7205 34357 7239 34391
rect 11069 34357 11103 34391
rect 28457 34357 28491 34391
rect 30665 34357 30699 34391
rect 2789 34153 2823 34187
rect 6009 34153 6043 34187
rect 8861 34153 8895 34187
rect 9873 34153 9907 34187
rect 11161 34153 11195 34187
rect 14381 34153 14415 34187
rect 29561 34153 29595 34187
rect 9965 34085 9999 34119
rect 10057 34085 10091 34119
rect 20361 34085 20395 34119
rect 21741 34085 21775 34119
rect 31585 34085 31619 34119
rect 4905 34017 4939 34051
rect 6745 34017 6779 34051
rect 7297 34017 7331 34051
rect 7481 34017 7515 34051
rect 8033 34017 8067 34051
rect 8677 34017 8711 34051
rect 11069 34017 11103 34051
rect 11529 34017 11563 34051
rect 11805 34017 11839 34051
rect 12081 34017 12115 34051
rect 15577 34017 15611 34051
rect 18705 34017 18739 34051
rect 18981 34017 19015 34051
rect 21281 34017 21315 34051
rect 23857 34017 23891 34051
rect 26617 34017 26651 34051
rect 28457 34017 28491 34051
rect 30297 34017 30331 34051
rect 31125 34017 31159 34051
rect 32137 34017 32171 34051
rect 32965 34017 32999 34051
rect 33425 34017 33459 34051
rect 34161 34017 34195 34051
rect 37013 34017 37047 34051
rect 1409 33949 1443 33983
rect 1685 33949 1719 33983
rect 4629 33949 4663 33983
rect 6929 33949 6963 33983
rect 9689 33949 9723 33983
rect 10425 33949 10459 33983
rect 13001 33949 13035 33983
rect 13277 33949 13311 33983
rect 16221 33949 16255 33983
rect 16497 33949 16531 33983
rect 21189 33949 21223 33983
rect 22201 33949 22235 33983
rect 22477 33949 22511 33983
rect 24317 33949 24351 33983
rect 24593 33949 24627 33983
rect 26525 33949 26559 33983
rect 28181 33949 28215 33983
rect 31033 33949 31067 33983
rect 32873 33949 32907 33983
rect 33885 33949 33919 33983
rect 36185 33949 36219 33983
rect 36737 33949 36771 33983
rect 37197 33949 37231 33983
rect 32321 33881 32355 33915
rect 15669 33813 15703 33847
rect 17785 33813 17819 33847
rect 25881 33813 25915 33847
rect 26801 33813 26835 33847
rect 30481 33813 30515 33847
rect 35265 33813 35299 33847
rect 1869 33609 1903 33643
rect 4169 33609 4203 33643
rect 9781 33609 9815 33643
rect 11897 33609 11931 33643
rect 15945 33609 15979 33643
rect 18153 33609 18187 33643
rect 22477 33609 22511 33643
rect 23949 33609 23983 33643
rect 24961 33609 24995 33643
rect 33517 33609 33551 33643
rect 37841 33609 37875 33643
rect 7573 33541 7607 33575
rect 12541 33541 12575 33575
rect 16497 33541 16531 33575
rect 2605 33473 2639 33507
rect 15761 33473 15795 33507
rect 17233 33473 17267 33507
rect 29837 33473 29871 33507
rect 32413 33473 32447 33507
rect 35633 33473 35667 33507
rect 1501 33405 1535 33439
rect 1685 33405 1719 33439
rect 2881 33405 2915 33439
rect 4721 33405 4755 33439
rect 5733 33405 5767 33439
rect 7021 33405 7055 33439
rect 7481 33405 7515 33439
rect 7665 33405 7699 33439
rect 8585 33405 8619 33439
rect 8953 33405 8987 33439
rect 9137 33405 9171 33439
rect 9781 33405 9815 33439
rect 11069 33405 11103 33439
rect 11253 33405 11287 33439
rect 11621 33405 11655 33439
rect 12541 33405 12575 33439
rect 13001 33405 13035 33439
rect 13369 33405 13403 33439
rect 13921 33405 13955 33439
rect 14197 33405 14231 33439
rect 15117 33405 15151 33439
rect 15669 33405 15703 33439
rect 16589 33405 16623 33439
rect 17141 33405 17175 33439
rect 18061 33405 18095 33439
rect 18429 33405 18463 33439
rect 19073 33405 19107 33439
rect 19349 33405 19383 33439
rect 20085 33405 20119 33439
rect 20361 33405 20395 33439
rect 22201 33405 22235 33439
rect 22293 33405 22327 33439
rect 23673 33405 23707 33439
rect 23765 33405 23799 33439
rect 24685 33405 24719 33439
rect 24777 33405 24811 33439
rect 25789 33405 25823 33439
rect 26065 33405 26099 33439
rect 28181 33405 28215 33439
rect 28365 33405 28399 33439
rect 28549 33405 28583 33439
rect 29561 33405 29595 33439
rect 32137 33405 32171 33439
rect 35541 33405 35575 33439
rect 35909 33405 35943 33439
rect 36461 33405 36495 33439
rect 36737 33405 36771 33439
rect 1593 33337 1627 33371
rect 5549 33337 5583 33371
rect 5917 33337 5951 33371
rect 6285 33337 6319 33371
rect 22109 33337 22143 33371
rect 4905 33269 4939 33303
rect 5825 33269 5859 33303
rect 21465 33269 21499 33303
rect 27169 33269 27203 33303
rect 30941 33269 30975 33303
rect 5641 33065 5675 33099
rect 11253 33065 11287 33099
rect 36645 33065 36679 33099
rect 2053 32997 2087 33031
rect 4077 32997 4111 33031
rect 13645 32997 13679 33031
rect 2605 32929 2639 32963
rect 2789 32929 2823 32963
rect 2973 32929 3007 32963
rect 3157 32929 3191 32963
rect 3341 32929 3375 32963
rect 4905 32929 4939 32963
rect 5549 32929 5583 32963
rect 7021 32929 7055 32963
rect 8217 32929 8251 32963
rect 8401 32929 8435 32963
rect 8585 32929 8619 32963
rect 8769 32929 8803 32963
rect 8953 32929 8987 32963
rect 9689 32929 9723 32963
rect 11989 32929 12023 32963
rect 14473 32929 14507 32963
rect 15577 32929 15611 32963
rect 17417 32929 17451 32963
rect 18160 32929 18194 32963
rect 20913 32929 20947 32963
rect 21649 32929 21683 32963
rect 21925 32929 21959 32963
rect 24317 32929 24351 32963
rect 26801 32929 26835 32963
rect 28641 32929 28675 32963
rect 29377 32929 29411 32963
rect 30573 32929 30607 32963
rect 31217 32929 31251 32963
rect 33241 32929 33275 32963
rect 33609 32929 33643 32963
rect 34253 32929 34287 32963
rect 34345 32929 34379 32963
rect 35357 32929 35391 32963
rect 36369 32929 36403 32963
rect 36921 32929 36955 32963
rect 4629 32861 4663 32895
rect 5089 32861 5123 32895
rect 6193 32861 6227 32895
rect 6745 32861 6779 32895
rect 7205 32861 7239 32895
rect 7665 32861 7699 32895
rect 9965 32861 9999 32895
rect 12265 32861 12299 32895
rect 15301 32861 15335 32895
rect 18429 32861 18463 32895
rect 24041 32861 24075 32895
rect 26525 32861 26559 32895
rect 31493 32861 31527 32895
rect 32781 32861 32815 32895
rect 33517 32861 33551 32895
rect 34805 32861 34839 32895
rect 35265 32861 35299 32895
rect 17601 32793 17635 32827
rect 30757 32793 30791 32827
rect 14657 32725 14691 32759
rect 16865 32725 16899 32759
rect 19533 32725 19567 32759
rect 21097 32725 21131 32759
rect 23213 32725 23247 32759
rect 25421 32725 25455 32759
rect 27905 32725 27939 32759
rect 28733 32725 28767 32759
rect 35541 32725 35575 32759
rect 28457 32521 28491 32555
rect 32781 32521 32815 32555
rect 34069 32521 34103 32555
rect 7757 32453 7791 32487
rect 12541 32453 12575 32487
rect 14381 32453 14415 32487
rect 20361 32453 20395 32487
rect 21833 32453 21867 32487
rect 24869 32453 24903 32487
rect 28089 32453 28123 32487
rect 30573 32453 30607 32487
rect 3341 32385 3375 32419
rect 5549 32385 5583 32419
rect 6285 32385 6319 32419
rect 13277 32385 13311 32419
rect 17509 32385 17543 32419
rect 18061 32385 18095 32419
rect 19073 32385 19107 32419
rect 20453 32385 20487 32419
rect 23673 32385 23707 32419
rect 27353 32385 27387 32419
rect 1685 32317 1719 32351
rect 2237 32317 2271 32351
rect 2421 32317 2455 32351
rect 3249 32317 3283 32351
rect 3709 32317 3743 32351
rect 3893 32317 3927 32351
rect 4261 32317 4295 32351
rect 4629 32317 4663 32351
rect 5733 32317 5767 32351
rect 5825 32317 5859 32351
rect 7021 32317 7055 32351
rect 8217 32317 8251 32351
rect 8677 32317 8711 32351
rect 9229 32317 9263 32351
rect 9413 32317 9447 32351
rect 10701 32317 10735 32351
rect 10885 32317 10919 32351
rect 11345 32317 11379 32351
rect 11621 32317 11655 32351
rect 12449 32317 12483 32351
rect 13001 32317 13035 32351
rect 14289 32317 14323 32351
rect 14933 32317 14967 32351
rect 15485 32317 15519 32351
rect 15761 32317 15795 32351
rect 16221 32317 16255 32351
rect 17049 32317 17083 32351
rect 18613 32317 18647 32351
rect 18889 32317 18923 32351
rect 19809 32317 19843 32351
rect 20361 32317 20395 32351
rect 22017 32317 22051 32351
rect 22201 32317 22235 32351
rect 22385 32317 22419 32351
rect 23765 32317 23799 32351
rect 24777 32317 24811 32351
rect 25053 32317 25087 32351
rect 25973 32317 26007 32351
rect 26249 32317 26283 32351
rect 31493 32385 31527 32419
rect 35817 32385 35851 32419
rect 28181 32317 28215 32351
rect 28273 32317 28307 32351
rect 29653 32317 29687 32351
rect 30205 32317 30239 32351
rect 30481 32317 30515 32351
rect 31217 32317 31251 32351
rect 33977 32317 34011 32351
rect 35541 32317 35575 32351
rect 37657 32317 37691 32351
rect 5917 32249 5951 32283
rect 8125 32249 8159 32283
rect 16773 32249 16807 32283
rect 17141 32249 17175 32283
rect 24225 32249 24259 32283
rect 28089 32249 28123 32283
rect 33793 32249 33827 32283
rect 1685 32181 1719 32215
rect 7205 32181 7239 32215
rect 16957 32181 16991 32215
rect 25237 32181 25271 32215
rect 36921 32181 36955 32215
rect 37749 32181 37783 32215
rect 9229 31977 9263 32011
rect 15393 31977 15427 32011
rect 23213 31977 23247 32011
rect 29469 31977 29503 32011
rect 34989 31977 35023 32011
rect 3065 31909 3099 31943
rect 6837 31909 6871 31943
rect 17969 31909 18003 31943
rect 18337 31909 18371 31943
rect 18705 31909 18739 31943
rect 20361 31909 20395 31943
rect 22385 31909 22419 31943
rect 32597 31909 32631 31943
rect 36277 31909 36311 31943
rect 1685 31841 1719 31875
rect 4629 31841 4663 31875
rect 7297 31841 7331 31875
rect 7665 31841 7699 31875
rect 8125 31841 8159 31875
rect 8585 31841 8619 31875
rect 9413 31841 9447 31875
rect 9689 31841 9723 31875
rect 9873 31841 9907 31875
rect 9965 31841 9999 31875
rect 11253 31841 11287 31875
rect 11805 31841 11839 31875
rect 12633 31841 12667 31875
rect 14289 31841 14323 31875
rect 14565 31841 14599 31875
rect 15485 31841 15519 31875
rect 15853 31841 15887 31875
rect 16865 31841 16899 31875
rect 18153 31841 18187 31875
rect 18245 31841 18279 31875
rect 19901 31841 19935 31875
rect 20085 31841 20119 31875
rect 21833 31841 21867 31875
rect 22201 31841 22235 31875
rect 23029 31841 23063 31875
rect 23765 31841 23799 31875
rect 24041 31841 24075 31875
rect 26893 31841 26927 31875
rect 27445 31841 27479 31875
rect 28365 31841 28399 31875
rect 30665 31841 30699 31875
rect 31217 31841 31251 31875
rect 32781 31841 32815 31875
rect 33609 31841 33643 31875
rect 35817 31841 35851 31875
rect 36737 31841 36771 31875
rect 37749 31841 37783 31875
rect 1409 31773 1443 31807
rect 5181 31773 5215 31807
rect 5457 31773 5491 31807
rect 12081 31773 12115 31807
rect 13737 31773 13771 31807
rect 14749 31773 14783 31807
rect 16221 31773 16255 31807
rect 21465 31773 21499 31807
rect 25329 31773 25363 31807
rect 26617 31773 26651 31807
rect 28089 31773 28123 31807
rect 31493 31773 31527 31807
rect 33149 31773 33183 31807
rect 33885 31773 33919 31807
rect 35725 31773 35759 31807
rect 37841 31773 37875 31807
rect 11345 31705 11379 31739
rect 27353 31705 27387 31739
rect 30757 31705 30791 31739
rect 4445 31637 4479 31671
rect 7389 31637 7423 31671
rect 10149 31637 10183 31671
rect 12725 31637 12759 31671
rect 17049 31637 17083 31671
rect 36829 31637 36863 31671
rect 7297 31433 7331 31467
rect 9413 31433 9447 31467
rect 15761 31433 15795 31467
rect 23029 31433 23063 31467
rect 26433 31433 26467 31467
rect 2881 31365 2915 31399
rect 5641 31365 5675 31399
rect 11437 31365 11471 31399
rect 22017 31365 22051 31399
rect 33977 31365 34011 31399
rect 1593 31297 1627 31331
rect 2329 31297 2363 31331
rect 7849 31297 7883 31331
rect 10793 31297 10827 31331
rect 13829 31297 13863 31331
rect 18429 31297 18463 31331
rect 24133 31297 24167 31331
rect 27261 31297 27295 31331
rect 31309 31297 31343 31331
rect 35817 31297 35851 31331
rect 36737 31297 36771 31331
rect 1777 31229 1811 31263
rect 1869 31229 1903 31263
rect 3065 31229 3099 31263
rect 3525 31229 3559 31263
rect 3893 31229 3927 31263
rect 4169 31229 4203 31263
rect 4445 31229 4479 31263
rect 5825 31229 5859 31263
rect 6193 31229 6227 31263
rect 7205 31229 7239 31263
rect 8125 31229 8159 31263
rect 9965 31229 9999 31263
rect 11161 31229 11195 31263
rect 11437 31229 11471 31263
rect 12449 31229 12483 31263
rect 13553 31229 13587 31263
rect 15669 31229 15703 31263
rect 16313 31229 16347 31263
rect 16681 31229 16715 31263
rect 16957 31229 16991 31263
rect 18337 31229 18371 31263
rect 18797 31229 18831 31263
rect 19625 31229 19659 31263
rect 20085 31229 20119 31263
rect 20361 31229 20395 31263
rect 20637 31229 20671 31263
rect 21557 31229 21591 31263
rect 21741 31229 21775 31263
rect 22109 31229 22143 31263
rect 22845 31229 22879 31263
rect 24041 31229 24075 31263
rect 24317 31229 24351 31263
rect 25421 31229 25455 31263
rect 25605 31229 25639 31263
rect 25789 31229 25823 31263
rect 26617 31229 26651 31263
rect 26985 31229 27019 31263
rect 28641 31229 28675 31263
rect 29469 31229 29503 31263
rect 30021 31229 30055 31263
rect 30389 31229 30423 31263
rect 31033 31229 31067 31263
rect 32689 31229 32723 31263
rect 33149 31229 33183 31263
rect 33517 31229 33551 31263
rect 33977 31229 34011 31263
rect 34897 31229 34931 31263
rect 35265 31229 35299 31263
rect 35725 31229 35759 31263
rect 36461 31229 36495 31263
rect 1961 31161 1995 31195
rect 15209 31161 15243 31195
rect 30573 31161 30607 31195
rect 10057 31093 10091 31127
rect 12633 31093 12667 31127
rect 20545 31093 20579 31127
rect 24501 31093 24535 31127
rect 37841 31093 37875 31127
rect 5733 30889 5767 30923
rect 14657 30889 14691 30923
rect 21005 30889 21039 30923
rect 23397 30889 23431 30923
rect 24225 30889 24259 30923
rect 25881 30889 25915 30923
rect 33609 30889 33643 30923
rect 36737 30889 36771 30923
rect 7849 30821 7883 30855
rect 16773 30821 16807 30855
rect 17141 30821 17175 30855
rect 2605 30753 2639 30787
rect 2973 30753 3007 30787
rect 3157 30753 3191 30787
rect 4997 30753 5031 30787
rect 5641 30753 5675 30787
rect 6837 30753 6871 30787
rect 7021 30753 7055 30787
rect 7389 30753 7423 30787
rect 8401 30753 8435 30787
rect 8677 30753 8711 30787
rect 9689 30753 9723 30787
rect 10333 30753 10367 30787
rect 11161 30753 11195 30787
rect 13553 30753 13587 30787
rect 13829 30753 13863 30787
rect 14565 30753 14599 30787
rect 15393 30753 15427 30787
rect 16129 30753 16163 30787
rect 16957 30753 16991 30787
rect 17049 30753 17083 30787
rect 17969 30753 18003 30787
rect 18521 30753 18555 30787
rect 19625 30753 19659 30787
rect 20361 30753 20395 30787
rect 20913 30753 20947 30787
rect 24317 30753 24351 30787
rect 24685 30753 24719 30787
rect 25789 30753 25823 30787
rect 26801 30753 26835 30787
rect 27169 30753 27203 30787
rect 27721 30753 27755 30787
rect 29837 30753 29871 30787
rect 30297 30753 30331 30787
rect 30665 30753 30699 30787
rect 32597 30753 32631 30787
rect 33517 30753 33551 30787
rect 34253 30753 34287 30787
rect 35357 30753 35391 30787
rect 35633 30753 35667 30787
rect 37749 30753 37783 30787
rect 8861 30685 8895 30719
rect 11437 30685 11471 30719
rect 13645 30685 13679 30719
rect 17509 30685 17543 30719
rect 19993 30685 20027 30719
rect 22017 30685 22051 30719
rect 22293 30685 22327 30719
rect 24961 30685 24995 30719
rect 27997 30685 28031 30719
rect 32505 30685 32539 30719
rect 33057 30685 33091 30719
rect 34345 30685 34379 30719
rect 3157 30617 3191 30651
rect 15485 30617 15519 30651
rect 26617 30617 26651 30651
rect 30665 30617 30699 30651
rect 5089 30549 5123 30583
rect 9781 30549 9815 30583
rect 10425 30549 10459 30583
rect 12725 30549 12759 30583
rect 18061 30549 18095 30583
rect 29285 30549 29319 30583
rect 37841 30549 37875 30583
rect 6193 30345 6227 30379
rect 13737 30345 13771 30379
rect 26709 30345 26743 30379
rect 32689 30345 32723 30379
rect 3617 30277 3651 30311
rect 9137 30277 9171 30311
rect 23949 30277 23983 30311
rect 28273 30277 28307 30311
rect 29377 30277 29411 30311
rect 1685 30209 1719 30243
rect 4353 30209 4387 30243
rect 9689 30209 9723 30243
rect 16497 30209 16531 30243
rect 20821 30209 20855 30243
rect 22017 30209 22051 30243
rect 24501 30209 24535 30243
rect 25605 30209 25639 30243
rect 36461 30209 36495 30243
rect 1409 30141 1443 30175
rect 3525 30141 3559 30175
rect 4077 30141 4111 30175
rect 5273 30141 5307 30175
rect 5365 30141 5399 30175
rect 6009 30141 6043 30175
rect 7021 30141 7055 30175
rect 7389 30141 7423 30175
rect 7665 30141 7699 30175
rect 8401 30141 8435 30175
rect 9321 30141 9355 30175
rect 9413 30141 9447 30175
rect 11529 30141 11563 30175
rect 12541 30141 12575 30175
rect 12909 30141 12943 30175
rect 13737 30141 13771 30175
rect 14289 30141 14323 30175
rect 14473 30141 14507 30175
rect 14933 30141 14967 30175
rect 15577 30141 15611 30175
rect 17049 30141 17083 30175
rect 17325 30141 17359 30175
rect 17509 30141 17543 30175
rect 18245 30141 18279 30175
rect 18981 30141 19015 30175
rect 19257 30141 19291 30175
rect 19993 30141 20027 30175
rect 20729 30141 20763 30175
rect 22385 30141 22419 30175
rect 22661 30141 22695 30175
rect 23857 30141 23891 30175
rect 24225 30141 24259 30175
rect 25329 30141 25363 30175
rect 27445 30141 27479 30175
rect 27813 30141 27847 30175
rect 28365 30141 28399 30175
rect 29469 30141 29503 30175
rect 29837 30141 29871 30175
rect 31125 30141 31159 30175
rect 31861 30141 31895 30175
rect 32045 30141 32079 30175
rect 32873 30141 32907 30175
rect 33241 30141 33275 30175
rect 33609 30141 33643 30175
rect 34161 30141 34195 30175
rect 35449 30141 35483 30175
rect 35633 30141 35667 30175
rect 36001 30141 36035 30175
rect 36737 30141 36771 30175
rect 7941 30073 7975 30107
rect 11069 30073 11103 30107
rect 22937 30073 22971 30107
rect 34345 30073 34379 30107
rect 2973 30005 3007 30039
rect 5089 30005 5123 30039
rect 5457 30005 5491 30039
rect 8585 30005 8619 30039
rect 11621 30005 11655 30039
rect 12541 30005 12575 30039
rect 15761 30005 15795 30039
rect 18337 30005 18371 30039
rect 19993 30005 20027 30039
rect 31217 30005 31251 30039
rect 37841 30005 37875 30039
rect 3065 29801 3099 29835
rect 4169 29801 4203 29835
rect 14565 29801 14599 29835
rect 29193 29801 29227 29835
rect 31493 29801 31527 29835
rect 11529 29733 11563 29767
rect 17141 29733 17175 29767
rect 20269 29733 20303 29767
rect 21281 29733 21315 29767
rect 33425 29733 33459 29767
rect 2237 29665 2271 29699
rect 2881 29665 2915 29699
rect 4077 29665 4111 29699
rect 4629 29665 4663 29699
rect 5365 29665 5399 29699
rect 5641 29665 5675 29699
rect 7481 29665 7515 29699
rect 7941 29665 7975 29699
rect 8125 29665 8159 29699
rect 8309 29665 8343 29699
rect 8953 29665 8987 29699
rect 9689 29665 9723 29699
rect 10425 29665 10459 29699
rect 12357 29665 12391 29699
rect 13001 29665 13035 29699
rect 15301 29665 15335 29699
rect 15945 29665 15979 29699
rect 16313 29665 16347 29699
rect 16957 29665 16991 29699
rect 20177 29665 20211 29699
rect 21741 29665 21775 29699
rect 22109 29665 22143 29699
rect 22937 29665 22971 29699
rect 23305 29665 23339 29699
rect 23581 29665 23615 29699
rect 24777 29665 24811 29699
rect 25053 29665 25087 29699
rect 25513 29665 25547 29699
rect 25973 29665 26007 29699
rect 26893 29665 26927 29699
rect 27353 29665 27387 29699
rect 29929 29665 29963 29699
rect 30297 29665 30331 29699
rect 30757 29665 30791 29699
rect 31677 29665 31711 29699
rect 32873 29665 32907 29699
rect 33149 29665 33183 29699
rect 33885 29665 33919 29699
rect 36093 29665 36127 29699
rect 36829 29665 36863 29699
rect 37749 29665 37783 29699
rect 7021 29597 7055 29631
rect 12081 29597 12115 29631
rect 12541 29597 12575 29631
rect 13277 29597 13311 29631
rect 15393 29597 15427 29631
rect 18061 29597 18095 29631
rect 18337 29597 18371 29631
rect 22201 29597 22235 29631
rect 24961 29597 24995 29631
rect 26985 29597 27019 29631
rect 27813 29597 27847 29631
rect 28089 29597 28123 29631
rect 32505 29597 32539 29631
rect 34161 29597 34195 29631
rect 37105 29597 37139 29631
rect 10609 29529 10643 29563
rect 22845 29529 22879 29563
rect 30849 29529 30883 29563
rect 36369 29529 36403 29563
rect 2329 29461 2363 29495
rect 9045 29461 9079 29495
rect 9873 29461 9907 29495
rect 19625 29461 19659 29495
rect 35265 29461 35299 29495
rect 37933 29461 37967 29495
rect 6929 29257 6963 29291
rect 10333 29257 10367 29291
rect 26893 29257 26927 29291
rect 28917 29257 28951 29291
rect 32965 29257 32999 29291
rect 37841 29257 37875 29291
rect 6193 29189 6227 29223
rect 14473 29189 14507 29223
rect 28089 29189 28123 29223
rect 5273 29121 5307 29155
rect 8401 29121 8435 29155
rect 15025 29121 15059 29155
rect 17233 29121 17267 29155
rect 18337 29121 18371 29155
rect 22661 29121 22695 29155
rect 25053 29121 25087 29155
rect 29929 29121 29963 29155
rect 30941 29121 30975 29155
rect 31401 29121 31435 29155
rect 31677 29121 31711 29155
rect 34345 29121 34379 29155
rect 35449 29121 35483 29155
rect 36461 29121 36495 29155
rect 36737 29121 36771 29155
rect 1869 29053 1903 29087
rect 1961 29053 1995 29087
rect 2697 29053 2731 29087
rect 2973 29053 3007 29087
rect 3525 29053 3559 29087
rect 3893 29053 3927 29087
rect 4537 29053 4571 29087
rect 4997 29053 5031 29087
rect 6009 29053 6043 29087
rect 7021 29053 7055 29087
rect 7389 29053 7423 29087
rect 8125 29053 8159 29087
rect 10517 29053 10551 29087
rect 10609 29053 10643 29087
rect 11253 29053 11287 29087
rect 12633 29053 12667 29087
rect 12817 29053 12851 29087
rect 13185 29053 13219 29087
rect 14381 29053 14415 29087
rect 14933 29053 14967 29087
rect 15853 29053 15887 29087
rect 16129 29053 16163 29087
rect 18705 29053 18739 29087
rect 18981 29053 19015 29087
rect 20177 29053 20211 29087
rect 20453 29053 20487 29087
rect 22385 29053 22419 29087
rect 23029 29053 23063 29087
rect 23673 29053 23707 29087
rect 24777 29053 24811 29087
rect 25237 29053 25271 29087
rect 25421 29053 25455 29087
rect 26065 29053 26099 29087
rect 27077 29053 27111 29087
rect 27169 29053 27203 29087
rect 27537 29053 27571 29087
rect 27997 29053 28031 29087
rect 29101 29053 29135 29087
rect 30389 29053 30423 29087
rect 30665 29053 30699 29087
rect 33977 29053 34011 29087
rect 35725 29053 35759 29087
rect 35909 29053 35943 29087
rect 19257 28985 19291 29019
rect 23765 28985 23799 29019
rect 33793 28985 33827 29019
rect 34897 28985 34931 29019
rect 2789 28917 2823 28951
rect 4537 28917 4571 28951
rect 9689 28917 9723 28951
rect 21557 28917 21591 28951
rect 7481 28713 7515 28747
rect 14289 28713 14323 28747
rect 17049 28713 17083 28747
rect 20361 28713 20395 28747
rect 21005 28713 21039 28747
rect 21649 28713 21683 28747
rect 22293 28713 22327 28747
rect 33609 28713 33643 28747
rect 37933 28713 37967 28747
rect 12173 28645 12207 28679
rect 16497 28645 16531 28679
rect 32505 28645 32539 28679
rect 33057 28645 33091 28679
rect 35173 28645 35207 28679
rect 4629 28577 4663 28611
rect 4905 28577 4939 28611
rect 5825 28577 5859 28611
rect 6193 28577 6227 28611
rect 7205 28577 7239 28611
rect 7665 28577 7699 28611
rect 8401 28577 8435 28611
rect 9965 28577 9999 28611
rect 10057 28577 10091 28611
rect 10425 28577 10459 28611
rect 11345 28577 11379 28611
rect 11897 28577 11931 28611
rect 12081 28577 12115 28611
rect 12725 28577 12759 28611
rect 13001 28577 13035 28611
rect 13553 28577 13587 28611
rect 14197 28577 14231 28611
rect 15393 28577 15427 28611
rect 15761 28577 15795 28611
rect 16221 28577 16255 28611
rect 16957 28577 16991 28611
rect 17693 28577 17727 28611
rect 18245 28577 18279 28611
rect 18521 28577 18555 28611
rect 19533 28577 19567 28611
rect 20085 28577 20119 28611
rect 20913 28577 20947 28611
rect 21557 28577 21591 28611
rect 22201 28577 22235 28611
rect 23029 28577 23063 28611
rect 23581 28577 23615 28611
rect 23673 28577 23707 28611
rect 24869 28577 24903 28611
rect 24961 28577 24995 28611
rect 25329 28577 25363 28611
rect 26525 28577 26559 28611
rect 27077 28577 27111 28611
rect 27721 28577 27755 28611
rect 28181 28577 28215 28611
rect 29193 28577 29227 28611
rect 29653 28577 29687 28611
rect 30665 28577 30699 28611
rect 31217 28577 31251 28611
rect 32689 28577 32723 28611
rect 33517 28577 33551 28611
rect 34253 28577 34287 28611
rect 35081 28577 35115 28611
rect 35725 28577 35759 28611
rect 36369 28577 36403 28611
rect 36461 28577 36495 28611
rect 37197 28577 37231 28611
rect 37749 28577 37783 28611
rect 1409 28509 1443 28543
rect 1685 28509 1719 28543
rect 4261 28509 4295 28543
rect 6653 28509 6687 28543
rect 18797 28509 18831 28543
rect 20177 28509 20211 28543
rect 23489 28509 23523 28543
rect 25789 28509 25823 28543
rect 26893 28509 26927 28543
rect 28273 28509 28307 28543
rect 31493 28509 31527 28543
rect 34345 28509 34379 28543
rect 4905 28441 4939 28475
rect 5733 28441 5767 28475
rect 13461 28441 13495 28475
rect 29009 28441 29043 28475
rect 30573 28441 30607 28475
rect 2973 28373 3007 28407
rect 8585 28373 8619 28407
rect 37105 28373 37139 28407
rect 1869 28169 1903 28203
rect 4353 28169 4387 28203
rect 17049 28169 17083 28203
rect 23029 28169 23063 28203
rect 31861 28169 31895 28203
rect 34161 28169 34195 28203
rect 35173 28169 35207 28203
rect 37933 28169 37967 28203
rect 3341 28101 3375 28135
rect 5825 28101 5859 28135
rect 7941 28101 7975 28135
rect 8677 28101 8711 28135
rect 12541 28101 12575 28135
rect 15577 28101 15611 28135
rect 18337 28101 18371 28135
rect 22661 28101 22695 28135
rect 25513 28101 25547 28135
rect 33241 28101 33275 28135
rect 5181 28033 5215 28067
rect 9965 28033 9999 28067
rect 10609 28033 10643 28067
rect 11161 28033 11195 28067
rect 11621 28033 11655 28067
rect 14565 28033 14599 28067
rect 16129 28033 16163 28067
rect 18889 28033 18923 28067
rect 22753 28033 22787 28067
rect 26893 28033 26927 28067
rect 32505 28033 32539 28067
rect 37105 28033 37139 28067
rect 1777 27965 1811 27999
rect 2789 27965 2823 27999
rect 3249 27965 3283 27999
rect 3433 27965 3467 27999
rect 4169 27965 4203 27999
rect 5365 27965 5399 27999
rect 5917 27965 5951 27999
rect 7021 27965 7055 27999
rect 7757 27965 7791 27999
rect 8861 27965 8895 27999
rect 9229 27965 9263 27999
rect 9321 27965 9355 27999
rect 9781 27965 9815 27999
rect 11437 27965 11471 27999
rect 12541 27965 12575 27999
rect 13185 27965 13219 27999
rect 13737 27965 13771 27999
rect 14473 27965 14507 27999
rect 15485 27965 15519 27999
rect 15945 27965 15979 27999
rect 16865 27965 16899 27999
rect 18061 27965 18095 27999
rect 18613 27965 18647 27999
rect 20269 27965 20303 27999
rect 20545 27965 20579 27999
rect 21189 27965 21223 27999
rect 22532 27965 22566 27999
rect 24409 27965 24443 27999
rect 24685 27965 24719 27999
rect 25145 27965 25179 27999
rect 25513 27965 25547 27999
rect 26525 27965 26559 27999
rect 26617 27965 26651 27999
rect 29285 27965 29319 27999
rect 29469 27965 29503 27999
rect 30297 27965 30331 27999
rect 30573 27965 30607 27999
rect 32873 27965 32907 27999
rect 33241 27965 33275 27999
rect 33977 27965 34011 27999
rect 34897 27965 34931 27999
rect 35081 27965 35115 27999
rect 36001 27965 36035 27999
rect 36645 27965 36679 27999
rect 36737 27965 36771 27999
rect 37749 27965 37783 27999
rect 22385 27897 22419 27931
rect 28273 27897 28307 27931
rect 29837 27897 29871 27931
rect 7205 27829 7239 27863
rect 13829 27829 13863 27863
rect 20269 27829 20303 27863
rect 21281 27829 21315 27863
rect 26341 27829 26375 27863
rect 4261 27625 4295 27659
rect 11437 27625 11471 27659
rect 6837 27557 6871 27591
rect 8953 27557 8987 27591
rect 20085 27557 20119 27591
rect 21281 27557 21315 27591
rect 37105 27557 37139 27591
rect 2697 27489 2731 27523
rect 3065 27489 3099 27523
rect 4077 27489 4111 27523
rect 4997 27489 5031 27523
rect 5457 27489 5491 27523
rect 7481 27489 7515 27523
rect 7757 27489 7791 27523
rect 8125 27489 8159 27523
rect 8493 27489 8527 27523
rect 9689 27489 9723 27523
rect 10425 27489 10459 27523
rect 11621 27489 11655 27523
rect 11805 27489 11839 27523
rect 12357 27489 12391 27523
rect 12725 27489 12759 27523
rect 13829 27489 13863 27523
rect 14013 27489 14047 27523
rect 14473 27489 14507 27523
rect 15669 27489 15703 27523
rect 16129 27489 16163 27523
rect 16865 27489 16899 27523
rect 17877 27489 17911 27523
rect 19533 27489 19567 27523
rect 19993 27489 20027 27523
rect 21373 27489 21407 27523
rect 22017 27489 22051 27523
rect 22385 27489 22419 27523
rect 22845 27489 22879 27523
rect 23397 27489 23431 27523
rect 23857 27489 23891 27523
rect 24133 27489 24167 27523
rect 24593 27489 24627 27523
rect 24961 27489 24995 27523
rect 25697 27489 25731 27523
rect 27261 27489 27295 27523
rect 27629 27489 27663 27523
rect 30297 27489 30331 27523
rect 30665 27489 30699 27523
rect 31217 27489 31251 27523
rect 32965 27489 32999 27523
rect 33333 27489 33367 27523
rect 34713 27489 34747 27523
rect 36553 27489 36587 27523
rect 36737 27489 36771 27523
rect 37749 27489 37783 27523
rect 2237 27421 2271 27455
rect 3157 27421 3191 27455
rect 5181 27421 5215 27455
rect 14749 27421 14783 27455
rect 15485 27421 15519 27455
rect 18153 27421 18187 27455
rect 23489 27421 23523 27455
rect 28181 27421 28215 27455
rect 28457 27421 28491 27455
rect 32505 27421 32539 27455
rect 34437 27421 34471 27455
rect 7297 27353 7331 27387
rect 10609 27353 10643 27387
rect 16221 27353 16255 27387
rect 20913 27353 20947 27387
rect 25881 27353 25915 27387
rect 27077 27353 27111 27387
rect 31125 27353 31159 27387
rect 33241 27353 33275 27387
rect 4813 27285 4847 27319
rect 9873 27285 9907 27319
rect 17049 27285 17083 27319
rect 29745 27285 29779 27319
rect 36001 27285 36035 27319
rect 37841 27285 37875 27319
rect 1501 27081 1535 27115
rect 1961 27081 1995 27115
rect 4077 27081 4111 27115
rect 5089 27081 5123 27115
rect 6193 27081 6227 27115
rect 22937 27081 22971 27115
rect 24501 27081 24535 27115
rect 31861 27081 31895 27115
rect 33793 27081 33827 27115
rect 17417 27013 17451 27047
rect 23995 27013 24029 27047
rect 28457 27013 28491 27047
rect 34529 27013 34563 27047
rect 8953 26945 8987 26979
rect 9229 26945 9263 26979
rect 20269 26945 20303 26979
rect 24225 26945 24259 26979
rect 25513 26945 25547 26979
rect 32413 26945 32447 26979
rect 35081 26945 35115 26979
rect 36737 26945 36771 26979
rect 1777 26877 1811 26911
rect 2697 26877 2731 26911
rect 3065 26877 3099 26911
rect 3433 26877 3467 26911
rect 4077 26877 4111 26911
rect 4629 26877 4663 26911
rect 4905 26877 4939 26911
rect 6101 26877 6135 26911
rect 7205 26877 7239 26911
rect 7941 26877 7975 26911
rect 10609 26877 10643 26911
rect 11437 26877 11471 26911
rect 11713 26877 11747 26911
rect 12449 26877 12483 26911
rect 12909 26877 12943 26911
rect 13277 26877 13311 26911
rect 14197 26877 14231 26911
rect 14749 26877 14783 26911
rect 15025 26877 15059 26911
rect 15945 26877 15979 26911
rect 16405 26877 16439 26911
rect 16589 26877 16623 26911
rect 17325 26877 17359 26911
rect 18061 26877 18095 26911
rect 18245 26877 18279 26911
rect 19257 26877 19291 26911
rect 19717 26877 19751 26911
rect 20085 26877 20119 26911
rect 20729 26877 20763 26911
rect 21005 26877 21039 26911
rect 22845 26877 22879 26911
rect 24087 26877 24121 26911
rect 25053 26877 25087 26911
rect 25605 26877 25639 26911
rect 25881 26877 25915 26911
rect 26249 26877 26283 26911
rect 27629 26877 27663 26911
rect 27905 26877 27939 26911
rect 28457 26877 28491 26911
rect 29285 26877 29319 26911
rect 29929 26877 29963 26911
rect 30389 26877 30423 26911
rect 30849 26877 30883 26911
rect 31677 26877 31711 26911
rect 32689 26877 32723 26911
rect 34713 26877 34747 26911
rect 35449 26877 35483 26911
rect 35725 26877 35759 26911
rect 36461 26877 36495 26911
rect 1685 26809 1719 26843
rect 4813 26809 4847 26843
rect 23857 26809 23891 26843
rect 31033 26809 31067 26843
rect 36001 26809 36035 26843
rect 7389 26741 7423 26775
rect 8125 26741 8159 26775
rect 11253 26741 11287 26775
rect 12541 26741 12575 26775
rect 14105 26741 14139 26775
rect 15853 26741 15887 26775
rect 18337 26741 18371 26775
rect 22109 26741 22143 26775
rect 29377 26741 29411 26775
rect 37841 26741 37875 26775
rect 15669 26537 15703 26571
rect 25881 26537 25915 26571
rect 26985 26537 27019 26571
rect 32321 26537 32355 26571
rect 19809 26469 19843 26503
rect 1409 26401 1443 26435
rect 1685 26401 1719 26435
rect 4813 26401 4847 26435
rect 7205 26401 7239 26435
rect 8585 26401 8619 26435
rect 8769 26401 8803 26435
rect 8953 26401 8987 26435
rect 10149 26401 10183 26435
rect 10609 26401 10643 26435
rect 11069 26401 11103 26435
rect 11713 26401 11747 26435
rect 11805 26401 11839 26435
rect 12541 26401 12575 26435
rect 13001 26401 13035 26435
rect 13737 26401 13771 26435
rect 14565 26401 14599 26435
rect 14749 26401 14783 26435
rect 15761 26401 15795 26435
rect 16129 26401 16163 26435
rect 16405 26401 16439 26435
rect 17601 26401 17635 26435
rect 17785 26401 17819 26435
rect 17969 26401 18003 26435
rect 18889 26401 18923 26435
rect 19257 26401 19291 26435
rect 19993 26401 20027 26435
rect 21097 26401 21131 26435
rect 21230 26401 21264 26435
rect 22293 26401 22327 26435
rect 22753 26401 22787 26435
rect 23213 26401 23247 26435
rect 23581 26401 23615 26435
rect 23765 26401 23799 26435
rect 24501 26401 24535 26435
rect 25053 26401 25087 26435
rect 25697 26401 25731 26435
rect 26801 26401 26835 26435
rect 27537 26401 27571 26435
rect 28089 26401 28123 26435
rect 29377 26401 29411 26435
rect 29653 26401 29687 26435
rect 30573 26401 30607 26435
rect 31125 26401 31159 26435
rect 32229 26401 32263 26435
rect 32965 26401 32999 26435
rect 33793 26401 33827 26435
rect 34621 26401 34655 26435
rect 34897 26401 34931 26435
rect 35541 26401 35575 26435
rect 36645 26401 36679 26435
rect 36829 26401 36863 26435
rect 37013 26401 37047 26435
rect 37749 26401 37783 26435
rect 4537 26333 4571 26367
rect 5917 26333 5951 26367
rect 10241 26333 10275 26367
rect 11161 26333 11195 26367
rect 13093 26333 13127 26367
rect 14289 26333 14323 26367
rect 17141 26333 17175 26367
rect 20361 26333 20395 26367
rect 20913 26333 20947 26367
rect 24961 26333 24995 26367
rect 28549 26333 28583 26367
rect 31217 26333 31251 26367
rect 33057 26333 33091 26367
rect 37841 26333 37875 26367
rect 2789 26265 2823 26299
rect 8401 26265 8435 26299
rect 18705 26265 18739 26299
rect 27813 26265 27847 26299
rect 29193 26265 29227 26299
rect 30665 26265 30699 26299
rect 36461 26265 36495 26299
rect 7389 26197 7423 26231
rect 21373 26197 21407 26231
rect 22201 26197 22235 26231
rect 33977 26197 34011 26231
rect 34621 26197 34655 26231
rect 1961 25993 1995 26027
rect 12541 25993 12575 26027
rect 16773 25993 16807 26027
rect 21005 25993 21039 26027
rect 28641 25993 28675 26027
rect 32597 25993 32631 26027
rect 34253 25993 34287 26027
rect 35357 25993 35391 26027
rect 5365 25925 5399 25959
rect 7757 25925 7791 25959
rect 15393 25925 15427 25959
rect 23949 25925 23983 25959
rect 2605 25857 2639 25891
rect 4629 25857 4663 25891
rect 10885 25857 10919 25891
rect 14657 25857 14691 25891
rect 18061 25857 18095 25891
rect 22201 25857 22235 25891
rect 23121 25857 23155 25891
rect 26709 25857 26743 25891
rect 30389 25857 30423 25891
rect 30665 25857 30699 25891
rect 1869 25789 1903 25823
rect 2697 25789 2731 25823
rect 3157 25789 3191 25823
rect 3249 25789 3283 25823
rect 4169 25789 4203 25823
rect 4353 25789 4387 25823
rect 5181 25789 5215 25823
rect 5917 25789 5951 25823
rect 6929 25789 6963 25823
rect 7941 25789 7975 25823
rect 8401 25789 8435 25823
rect 8861 25789 8895 25823
rect 8953 25789 8987 25823
rect 9321 25789 9355 25823
rect 10057 25789 10091 25823
rect 12449 25789 12483 25823
rect 13737 25789 13771 25823
rect 13921 25789 13955 25823
rect 14381 25789 14415 25823
rect 15577 25789 15611 25823
rect 15761 25789 15795 25823
rect 15945 25789 15979 25823
rect 17049 25789 17083 25823
rect 18521 25789 18555 25823
rect 18705 25789 18739 25823
rect 18889 25789 18923 25823
rect 19901 25789 19935 25823
rect 20269 25789 20303 25823
rect 20637 25789 20671 25823
rect 20913 25789 20947 25823
rect 21925 25789 21959 25823
rect 22385 25789 22419 25823
rect 22937 25789 22971 25823
rect 23673 25789 23707 25823
rect 24409 25789 24443 25823
rect 24685 25789 24719 25823
rect 25421 25789 25455 25823
rect 26433 25789 26467 25823
rect 28089 25789 28123 25823
rect 28549 25789 28583 25823
rect 29653 25789 29687 25823
rect 32045 25789 32079 25823
rect 32505 25789 32539 25823
rect 32873 25789 32907 25823
rect 33425 25789 33459 25823
rect 34161 25789 34195 25823
rect 35541 25789 35575 25823
rect 36001 25789 36035 25823
rect 36461 25789 36495 25823
rect 36737 25789 36771 25823
rect 11253 25721 11287 25755
rect 11621 25721 11655 25755
rect 16957 25721 16991 25755
rect 17509 25721 17543 25755
rect 6009 25653 6043 25687
rect 7113 25653 7147 25687
rect 10241 25653 10275 25687
rect 11069 25653 11103 25687
rect 11161 25653 11195 25687
rect 21741 25653 21775 25687
rect 25605 25653 25639 25687
rect 29837 25653 29871 25687
rect 37841 25653 37875 25687
rect 4261 25449 4295 25483
rect 8033 25449 8067 25483
rect 15853 25449 15887 25483
rect 1409 25313 1443 25347
rect 4077 25313 4111 25347
rect 5457 25313 5491 25347
rect 5641 25313 5675 25347
rect 6009 25313 6043 25347
rect 8585 25313 8619 25347
rect 11805 25313 11839 25347
rect 12633 25313 12667 25347
rect 15669 25313 15703 25347
rect 16865 25313 16899 25347
rect 17049 25313 17083 25347
rect 17233 25313 17267 25347
rect 17877 25313 17911 25347
rect 18797 25313 18831 25347
rect 21741 25313 21775 25347
rect 22017 25313 22051 25347
rect 22293 25313 22327 25347
rect 22937 25313 22971 25347
rect 23121 25313 23155 25347
rect 24041 25313 24075 25347
rect 24188 25313 24222 25347
rect 25513 25313 25547 25347
rect 25973 25313 26007 25347
rect 26525 25313 26559 25347
rect 27077 25313 27111 25347
rect 28181 25313 28215 25347
rect 30573 25313 30607 25347
rect 30757 25313 30791 25347
rect 30941 25313 30975 25347
rect 32137 25313 32171 25347
rect 32781 25313 32815 25347
rect 37749 25313 37783 25347
rect 1685 25245 1719 25279
rect 6469 25245 6503 25279
rect 6745 25245 6779 25279
rect 9689 25245 9723 25279
rect 9965 25245 9999 25279
rect 12909 25245 12943 25279
rect 18521 25245 18555 25279
rect 19901 25245 19935 25279
rect 22109 25245 22143 25279
rect 24409 25245 24443 25279
rect 24777 25245 24811 25279
rect 26893 25245 26927 25279
rect 27905 25245 27939 25279
rect 29561 25245 29595 25279
rect 33057 25245 33091 25279
rect 35357 25245 35391 25279
rect 35633 25245 35667 25279
rect 16681 25177 16715 25211
rect 17969 25177 18003 25211
rect 24317 25177 24351 25211
rect 37933 25177 37967 25211
rect 2973 25109 3007 25143
rect 8769 25109 8803 25143
rect 11253 25109 11287 25143
rect 11989 25109 12023 25143
rect 14197 25109 14231 25143
rect 25329 25109 25363 25143
rect 32229 25109 32263 25143
rect 34161 25109 34195 25143
rect 36737 25109 36771 25143
rect 36461 24905 36495 24939
rect 20085 24837 20119 24871
rect 25513 24837 25547 24871
rect 28181 24837 28215 24871
rect 2329 24769 2363 24803
rect 3065 24769 3099 24803
rect 4169 24769 4203 24803
rect 5549 24769 5583 24803
rect 7205 24769 7239 24803
rect 7757 24769 7791 24803
rect 8217 24769 8251 24803
rect 12449 24769 12483 24803
rect 13461 24769 13495 24803
rect 13921 24769 13955 24803
rect 17233 24769 17267 24803
rect 21097 24769 21131 24803
rect 24685 24769 24719 24803
rect 27445 24769 27479 24803
rect 32137 24769 32171 24803
rect 34345 24769 34379 24803
rect 35173 24769 35207 24803
rect 1869 24701 1903 24735
rect 2145 24701 2179 24735
rect 2789 24701 2823 24735
rect 5273 24701 5307 24735
rect 5365 24701 5399 24735
rect 5733 24701 5767 24735
rect 8033 24701 8067 24735
rect 9229 24701 9263 24735
rect 9873 24701 9907 24735
rect 10149 24701 10183 24735
rect 10609 24701 10643 24735
rect 10885 24701 10919 24735
rect 11621 24701 11655 24735
rect 13001 24701 13035 24735
rect 13277 24701 13311 24735
rect 14473 24701 14507 24735
rect 14749 24701 14783 24735
rect 14933 24701 14967 24735
rect 15669 24701 15703 24735
rect 16497 24701 16531 24735
rect 17141 24701 17175 24735
rect 18613 24701 18647 24735
rect 18797 24701 18831 24735
rect 18981 24701 19015 24735
rect 19901 24701 19935 24735
rect 21281 24701 21315 24735
rect 21649 24701 21683 24735
rect 21833 24701 21867 24735
rect 22477 24701 22511 24735
rect 22661 24701 22695 24735
rect 23673 24701 23707 24735
rect 24961 24701 24995 24735
rect 25421 24701 25455 24735
rect 26157 24701 26191 24735
rect 27721 24701 27755 24735
rect 28089 24701 28123 24735
rect 29285 24701 29319 24735
rect 29837 24701 29871 24735
rect 30481 24701 30515 24735
rect 31401 24701 31435 24735
rect 32045 24701 32079 24735
rect 32873 24701 32907 24735
rect 33885 24701 33919 24735
rect 34897 24701 34931 24735
rect 37197 24701 37231 24735
rect 37565 24701 37599 24735
rect 9597 24633 9631 24667
rect 18153 24633 18187 24667
rect 33609 24633 33643 24667
rect 33977 24633 34011 24667
rect 37749 24633 37783 24667
rect 11805 24565 11839 24599
rect 15853 24565 15887 24599
rect 16497 24565 16531 24599
rect 23857 24565 23891 24599
rect 26341 24565 26375 24599
rect 29377 24565 29411 24599
rect 30573 24565 30607 24599
rect 31401 24565 31435 24599
rect 33057 24565 33091 24599
rect 33793 24565 33827 24599
rect 1777 24361 1811 24395
rect 16313 24361 16347 24395
rect 27629 24361 27663 24395
rect 37841 24361 37875 24395
rect 6929 24293 6963 24327
rect 8585 24293 8619 24327
rect 8769 24293 8803 24327
rect 9689 24293 9723 24327
rect 22017 24293 22051 24327
rect 1685 24225 1719 24259
rect 2329 24225 2363 24259
rect 3065 24225 3099 24259
rect 5089 24225 5123 24259
rect 6469 24225 6503 24259
rect 7757 24225 7791 24259
rect 8677 24225 8711 24259
rect 9137 24225 9171 24259
rect 10241 24225 10275 24259
rect 10517 24225 10551 24259
rect 10701 24225 10735 24259
rect 12357 24225 12391 24259
rect 13277 24225 13311 24259
rect 13829 24225 13863 24259
rect 14197 24225 14231 24259
rect 15301 24225 15335 24259
rect 16405 24225 16439 24259
rect 16957 24225 16991 24259
rect 18153 24225 18187 24259
rect 18613 24225 18647 24259
rect 20085 24225 20119 24259
rect 21097 24225 21131 24259
rect 21281 24225 21315 24259
rect 21741 24225 21775 24259
rect 22753 24225 22787 24259
rect 23673 24225 23707 24259
rect 24317 24225 24351 24259
rect 24501 24225 24535 24259
rect 25053 24225 25087 24259
rect 25697 24225 25731 24259
rect 26525 24225 26559 24259
rect 27537 24225 27571 24259
rect 28273 24225 28307 24259
rect 29101 24225 29135 24259
rect 31309 24225 31343 24259
rect 32137 24225 32171 24259
rect 32689 24225 32723 24259
rect 34161 24225 34195 24259
rect 34529 24225 34563 24259
rect 34713 24225 34747 24259
rect 35541 24225 35575 24259
rect 36277 24225 36311 24259
rect 36553 24225 36587 24259
rect 36829 24225 36863 24259
rect 37749 24225 37783 24259
rect 3157 24157 3191 24191
rect 4813 24157 4847 24191
rect 7481 24157 7515 24191
rect 7941 24157 7975 24191
rect 8401 24157 8435 24191
rect 11529 24157 11563 24191
rect 12081 24157 12115 24191
rect 12219 24157 12253 24191
rect 17049 24157 17083 24191
rect 18889 24157 18923 24191
rect 28365 24157 28399 24191
rect 29377 24157 29411 24191
rect 34253 24157 34287 24191
rect 2421 24089 2455 24123
rect 14105 24089 14139 24123
rect 18337 24089 18371 24123
rect 22937 24089 22971 24123
rect 25881 24089 25915 24123
rect 31493 24089 31527 24123
rect 32229 24089 32263 24123
rect 36921 24089 36955 24123
rect 15485 24021 15519 24055
rect 20269 24021 20303 24055
rect 24593 24021 24627 24055
rect 25145 24021 25179 24055
rect 26709 24021 26743 24055
rect 30481 24021 30515 24055
rect 33609 24021 33643 24055
rect 7389 23817 7423 23851
rect 23029 23817 23063 23851
rect 23949 23817 23983 23851
rect 29653 23817 29687 23851
rect 32597 23817 32631 23851
rect 14289 23749 14323 23783
rect 17141 23749 17175 23783
rect 1869 23681 1903 23715
rect 2421 23681 2455 23715
rect 5825 23681 5859 23715
rect 8033 23681 8067 23715
rect 10701 23681 10735 23715
rect 11529 23681 11563 23715
rect 13093 23681 13127 23715
rect 13553 23681 13587 23715
rect 19349 23681 19383 23715
rect 20453 23681 20487 23715
rect 22201 23681 22235 23715
rect 24961 23681 24995 23715
rect 26525 23681 26559 23715
rect 30113 23681 30147 23715
rect 30665 23681 30699 23715
rect 31493 23681 31527 23715
rect 35725 23681 35759 23715
rect 36461 23681 36495 23715
rect 2697 23613 2731 23647
rect 2881 23613 2915 23647
rect 3341 23613 3375 23647
rect 4353 23613 4387 23647
rect 5181 23613 5215 23647
rect 5457 23613 5491 23647
rect 5917 23613 5951 23647
rect 7205 23613 7239 23647
rect 8125 23613 8159 23647
rect 8585 23613 8619 23647
rect 8953 23613 8987 23647
rect 9413 23613 9447 23647
rect 10149 23613 10183 23647
rect 11161 23613 11195 23647
rect 11713 23613 11747 23647
rect 12541 23613 12575 23647
rect 13369 23613 13403 23647
rect 14197 23613 14231 23647
rect 14749 23613 14783 23647
rect 14933 23613 14967 23647
rect 15577 23613 15611 23647
rect 16405 23613 16439 23647
rect 16773 23613 16807 23647
rect 17141 23613 17175 23647
rect 18521 23613 18555 23647
rect 18981 23613 19015 23647
rect 19257 23613 19291 23647
rect 20361 23613 20395 23647
rect 20821 23613 20855 23647
rect 21557 23613 21591 23647
rect 22109 23613 22143 23647
rect 22845 23613 22879 23647
rect 24501 23613 24535 23647
rect 24593 23613 24627 23647
rect 24869 23613 24903 23647
rect 26801 23613 26835 23647
rect 26985 23613 27019 23647
rect 27721 23613 27755 23647
rect 28273 23613 28307 23647
rect 28457 23613 28491 23647
rect 30205 23613 30239 23647
rect 30573 23613 30607 23647
rect 31217 23613 31251 23647
rect 33885 23613 33919 23647
rect 34161 23613 34195 23647
rect 35449 23613 35483 23647
rect 35633 23613 35667 23647
rect 36737 23613 36771 23647
rect 3433 23545 3467 23579
rect 9965 23545 9999 23579
rect 10333 23545 10367 23579
rect 25973 23545 26007 23579
rect 34345 23545 34379 23579
rect 4445 23477 4479 23511
rect 10241 23477 10275 23511
rect 15669 23477 15703 23511
rect 21557 23477 21591 23511
rect 27721 23477 27755 23511
rect 37841 23477 37875 23511
rect 17141 23273 17175 23307
rect 21005 23273 21039 23307
rect 28089 23273 28123 23307
rect 31493 23273 31527 23307
rect 37841 23273 37875 23307
rect 24317 23205 24351 23239
rect 29285 23205 29319 23239
rect 32413 23205 32447 23239
rect 32965 23205 32999 23239
rect 1685 23137 1719 23171
rect 2605 23137 2639 23171
rect 2973 23137 3007 23171
rect 3341 23137 3375 23171
rect 4537 23137 4571 23171
rect 6745 23137 6779 23171
rect 6929 23137 6963 23171
rect 7389 23137 7423 23171
rect 7941 23137 7975 23171
rect 8125 23137 8159 23171
rect 8861 23137 8895 23171
rect 10701 23137 10735 23171
rect 11345 23137 11379 23171
rect 11437 23137 11471 23171
rect 12173 23137 12207 23171
rect 12633 23137 12667 23171
rect 13829 23137 13863 23171
rect 14381 23137 14415 23171
rect 15485 23137 15519 23171
rect 16221 23137 16255 23171
rect 16773 23137 16807 23171
rect 17417 23137 17451 23171
rect 17877 23137 17911 23171
rect 18521 23137 18555 23171
rect 19073 23137 19107 23171
rect 19349 23137 19383 23171
rect 20085 23137 20119 23171
rect 21189 23137 21223 23171
rect 21741 23137 21775 23171
rect 22477 23137 22511 23171
rect 23213 23137 23247 23171
rect 24133 23137 24167 23171
rect 24225 23137 24259 23171
rect 24685 23137 24719 23171
rect 25145 23137 25179 23171
rect 26801 23137 26835 23171
rect 28641 23137 28675 23171
rect 29929 23137 29963 23171
rect 30297 23137 30331 23171
rect 30481 23137 30515 23171
rect 31309 23137 31343 23171
rect 32597 23137 32631 23171
rect 33425 23137 33459 23171
rect 33701 23137 33735 23171
rect 36001 23137 36035 23171
rect 36461 23137 36495 23171
rect 37749 23137 37783 23171
rect 2421 23069 2455 23103
rect 4261 23069 4295 23103
rect 11161 23069 11195 23103
rect 14473 23069 14507 23103
rect 21649 23069 21683 23103
rect 23949 23069 23983 23103
rect 26525 23069 26559 23103
rect 30021 23069 30055 23103
rect 36553 23069 36587 23103
rect 6561 23001 6595 23035
rect 9045 23001 9079 23035
rect 13921 23001 13955 23035
rect 15669 23001 15703 23035
rect 19349 23001 19383 23035
rect 25329 23001 25363 23035
rect 1777 22933 1811 22967
rect 5641 22933 5675 22967
rect 12725 22933 12759 22967
rect 20269 22933 20303 22967
rect 22661 22933 22695 22967
rect 23397 22933 23431 22967
rect 28733 22933 28767 22967
rect 34989 22933 35023 22967
rect 3617 22729 3651 22763
rect 22753 22729 22787 22763
rect 37473 22729 37507 22763
rect 8677 22661 8711 22695
rect 11253 22661 11287 22695
rect 17141 22661 17175 22695
rect 20269 22661 20303 22695
rect 30021 22661 30055 22695
rect 31033 22661 31067 22695
rect 1409 22593 1443 22627
rect 1685 22593 1719 22627
rect 7389 22593 7423 22627
rect 8125 22593 8159 22627
rect 13185 22593 13219 22627
rect 16497 22593 16531 22627
rect 24409 22593 24443 22627
rect 27353 22593 27387 22627
rect 27905 22593 27939 22627
rect 28365 22593 28399 22627
rect 31585 22593 31619 22627
rect 34345 22593 34379 22627
rect 35265 22593 35299 22627
rect 36369 22593 36403 22627
rect 3709 22525 3743 22559
rect 3893 22525 3927 22559
rect 4537 22525 4571 22559
rect 5457 22525 5491 22559
rect 5733 22525 5767 22559
rect 6101 22525 6135 22559
rect 7573 22525 7607 22559
rect 7665 22525 7699 22559
rect 9413 22525 9447 22559
rect 9597 22525 9631 22559
rect 10057 22525 10091 22559
rect 10333 22525 10367 22559
rect 11345 22525 11379 22559
rect 11897 22525 11931 22559
rect 12633 22525 12667 22559
rect 14381 22525 14415 22559
rect 14473 22525 14507 22559
rect 15025 22525 15059 22559
rect 15485 22525 15519 22559
rect 16681 22525 16715 22559
rect 17233 22525 17267 22559
rect 18061 22525 18095 22559
rect 19257 22525 19291 22559
rect 19441 22525 19475 22559
rect 20361 22525 20395 22559
rect 20913 22525 20947 22559
rect 21833 22525 21867 22559
rect 22569 22525 22603 22559
rect 23673 22525 23707 22559
rect 24133 22525 24167 22559
rect 25881 22525 25915 22559
rect 26157 22525 26191 22559
rect 26341 22525 26375 22559
rect 28181 22525 28215 22559
rect 29561 22525 29595 22559
rect 29745 22525 29779 22559
rect 30113 22525 30147 22559
rect 30849 22525 30883 22559
rect 31861 22525 31895 22559
rect 33793 22525 33827 22559
rect 33977 22525 34011 22559
rect 34897 22525 34931 22559
rect 35449 22525 35483 22559
rect 36093 22525 36127 22559
rect 7757 22457 7791 22491
rect 9045 22457 9079 22491
rect 12449 22457 12483 22491
rect 12817 22457 12851 22491
rect 19717 22457 19751 22491
rect 25329 22457 25363 22491
rect 2973 22389 3007 22423
rect 12725 22389 12759 22423
rect 14749 22389 14783 22423
rect 18245 22389 18279 22423
rect 22017 22389 22051 22423
rect 33149 22389 33183 22423
rect 5733 22185 5767 22219
rect 13277 22185 13311 22219
rect 17509 22185 17543 22219
rect 19625 22185 19659 22219
rect 24133 22185 24167 22219
rect 26801 22185 26835 22219
rect 28365 22185 28399 22219
rect 30113 22185 30147 22219
rect 14013 22117 14047 22151
rect 15485 22117 15519 22151
rect 19809 22117 19843 22151
rect 20177 22117 20211 22151
rect 36645 22117 36679 22151
rect 1777 22049 1811 22083
rect 2605 22049 2639 22083
rect 3157 22049 3191 22083
rect 4353 22049 4387 22083
rect 4813 22049 4847 22083
rect 5549 22049 5583 22083
rect 6653 22049 6687 22083
rect 7205 22049 7239 22083
rect 7665 22049 7699 22083
rect 8125 22049 8159 22083
rect 8585 22049 8619 22083
rect 9505 22049 9539 22083
rect 9689 22049 9723 22083
rect 10057 22049 10091 22083
rect 10425 22049 10459 22083
rect 14105 22049 14139 22083
rect 15577 22049 15611 22083
rect 16589 22049 16623 22083
rect 16957 22049 16991 22083
rect 17785 22049 17819 22083
rect 18245 22049 18279 22083
rect 19073 22049 19107 22083
rect 19717 22049 19751 22083
rect 20913 22049 20947 22083
rect 22017 22049 22051 22083
rect 22385 22049 22419 22083
rect 22753 22049 22787 22083
rect 23397 22049 23431 22083
rect 23949 22049 23983 22083
rect 25421 22049 25455 22083
rect 25697 22049 25731 22083
rect 26893 22049 26927 22083
rect 27353 22049 27387 22083
rect 27537 22049 27571 22083
rect 28549 22049 28583 22083
rect 29101 22049 29135 22083
rect 29837 22049 29871 22083
rect 30665 22049 30699 22083
rect 30849 22049 30883 22083
rect 31401 22049 31435 22083
rect 32137 22049 32171 22083
rect 32689 22049 32723 22083
rect 33149 22049 33183 22083
rect 33333 22049 33367 22083
rect 33793 22049 33827 22083
rect 34529 22049 34563 22083
rect 35081 22049 35115 22083
rect 35541 22049 35575 22083
rect 35817 22049 35851 22083
rect 36737 22049 36771 22083
rect 37749 22049 37783 22083
rect 3433 21981 3467 22015
rect 7297 21981 7331 22015
rect 10609 21981 10643 22015
rect 11713 21981 11747 22015
rect 11989 21981 12023 22015
rect 19441 21981 19475 22015
rect 24961 21981 24995 22015
rect 25973 21981 26007 22015
rect 29009 21981 29043 22015
rect 32229 21981 32263 22015
rect 34805 21981 34839 22015
rect 2513 21913 2547 21947
rect 4169 21913 4203 21947
rect 8769 21913 8803 21947
rect 13829 21913 13863 21947
rect 15301 21913 15335 21947
rect 18889 21913 18923 21947
rect 21097 21913 21131 21947
rect 23397 21913 23431 21947
rect 1869 21845 1903 21879
rect 9321 21845 9355 21879
rect 14289 21845 14323 21879
rect 15761 21845 15795 21879
rect 31493 21845 31527 21879
rect 36461 21845 36495 21879
rect 36921 21845 36955 21879
rect 37841 21845 37875 21879
rect 8493 21641 8527 21675
rect 17601 21641 17635 21675
rect 21649 21641 21683 21675
rect 23949 21641 23983 21675
rect 28641 21641 28675 21675
rect 33977 21641 34011 21675
rect 11529 21573 11563 21607
rect 23213 21573 23247 21607
rect 26893 21573 26927 21607
rect 2237 21505 2271 21539
rect 9229 21505 9263 21539
rect 10149 21505 10183 21539
rect 16405 21505 16439 21539
rect 17325 21505 17359 21539
rect 23673 21505 23707 21539
rect 24961 21505 24995 21539
rect 27629 21505 27663 21539
rect 32781 21505 32815 21539
rect 35173 21505 35207 21539
rect 1501 21437 1535 21471
rect 2421 21437 2455 21471
rect 2789 21437 2823 21471
rect 3157 21437 3191 21471
rect 3433 21437 3467 21471
rect 4905 21437 4939 21471
rect 5089 21437 5123 21471
rect 5181 21437 5215 21471
rect 5457 21437 5491 21471
rect 5825 21437 5859 21471
rect 7389 21437 7423 21471
rect 8401 21437 8435 21471
rect 9597 21437 9631 21471
rect 9873 21437 9907 21471
rect 10609 21437 10643 21471
rect 11345 21437 11379 21471
rect 12449 21437 12483 21471
rect 13737 21437 13771 21471
rect 14013 21437 14047 21471
rect 14197 21437 14231 21471
rect 14657 21437 14691 21471
rect 15485 21437 15519 21471
rect 15761 21437 15795 21471
rect 16129 21437 16163 21471
rect 16865 21437 16899 21471
rect 17417 21437 17451 21471
rect 18245 21437 18279 21471
rect 18613 21437 18647 21471
rect 18981 21437 19015 21471
rect 19533 21437 19567 21471
rect 19809 21437 19843 21471
rect 19993 21437 20027 21471
rect 20545 21437 20579 21471
rect 21833 21437 21867 21471
rect 22201 21437 22235 21471
rect 22569 21437 22603 21471
rect 23397 21437 23431 21471
rect 23765 21437 23799 21471
rect 24685 21437 24719 21471
rect 26893 21437 26927 21471
rect 27353 21437 27387 21471
rect 28457 21437 28491 21471
rect 29561 21437 29595 21471
rect 29745 21437 29779 21471
rect 30113 21437 30147 21471
rect 30849 21437 30883 21471
rect 31309 21437 31343 21471
rect 32505 21437 32539 21471
rect 32873 21437 32907 21471
rect 32965 21437 32999 21471
rect 33885 21437 33919 21471
rect 34897 21437 34931 21471
rect 37013 21437 37047 21471
rect 37657 21437 37691 21471
rect 37841 21437 37875 21471
rect 10701 21369 10735 21403
rect 13185 21369 13219 21403
rect 19165 21369 19199 21403
rect 20453 21369 20487 21403
rect 31585 21369 31619 21403
rect 1593 21301 1627 21335
rect 4445 21301 4479 21335
rect 7573 21301 7607 21335
rect 12541 21301 12575 21335
rect 14749 21301 14783 21335
rect 17049 21301 17083 21335
rect 26065 21301 26099 21335
rect 29377 21301 29411 21335
rect 36277 21301 36311 21335
rect 37289 21301 37323 21335
rect 4261 21097 4295 21131
rect 8401 21097 8435 21131
rect 11345 21097 11379 21131
rect 14657 21097 14691 21131
rect 19809 21097 19843 21131
rect 30297 21097 30331 21131
rect 37841 21097 37875 21131
rect 16773 21029 16807 21063
rect 19993 21029 20027 21063
rect 20361 21029 20395 21063
rect 32137 21029 32171 21063
rect 1869 20961 1903 20995
rect 2329 20961 2363 20995
rect 2973 20961 3007 20995
rect 3433 20961 3467 20995
rect 4169 20961 4203 20995
rect 5089 20961 5123 20995
rect 5457 20961 5491 20995
rect 5641 20961 5675 20995
rect 6193 20961 6227 20995
rect 7297 20961 7331 20995
rect 7389 20961 7423 20995
rect 8309 20961 8343 20995
rect 8953 20961 8987 20995
rect 9781 20961 9815 20995
rect 10057 20961 10091 20995
rect 13369 20961 13403 20995
rect 13737 20961 13771 20995
rect 14565 20961 14599 20995
rect 15853 20961 15887 20995
rect 16037 20961 16071 20995
rect 16497 20961 16531 20995
rect 17233 20961 17267 20995
rect 17785 20961 17819 20995
rect 18429 20961 18463 20995
rect 18889 20961 18923 20995
rect 19901 20961 19935 20995
rect 21649 20961 21683 20995
rect 21741 20961 21775 20995
rect 22109 20961 22143 20995
rect 23029 20961 23063 20995
rect 25145 20961 25179 20995
rect 27261 20961 27295 20995
rect 27629 20961 27663 20995
rect 27997 20961 28031 20995
rect 28273 20961 28307 20995
rect 28917 20961 28951 20995
rect 29193 20961 29227 20995
rect 31309 20961 31343 20995
rect 32597 20961 32631 20995
rect 32965 20961 32999 20995
rect 33057 20961 33091 20995
rect 33885 20961 33919 20995
rect 34345 20961 34379 20995
rect 34713 20961 34747 20995
rect 34897 20961 34931 20995
rect 35541 20961 35575 20995
rect 36645 20961 36679 20995
rect 37013 20961 37047 20995
rect 37749 20961 37783 20995
rect 3157 20893 3191 20927
rect 6285 20893 6319 20927
rect 7849 20893 7883 20927
rect 12909 20893 12943 20927
rect 19533 20893 19567 20927
rect 19625 20893 19659 20927
rect 23305 20893 23339 20927
rect 24409 20893 24443 20927
rect 34161 20893 34195 20927
rect 36829 20893 36863 20927
rect 1685 20825 1719 20859
rect 9045 20825 9079 20859
rect 13645 20825 13679 20859
rect 18153 20825 18187 20859
rect 31493 20825 31527 20859
rect 7113 20757 7147 20791
rect 19533 20757 19567 20791
rect 21465 20757 21499 20791
rect 25329 20757 25363 20791
rect 28181 20757 28215 20791
rect 3617 20553 3651 20587
rect 10609 20553 10643 20587
rect 14013 20553 14047 20587
rect 14565 20553 14599 20587
rect 20085 20553 20119 20587
rect 20637 20553 20671 20587
rect 23305 20553 23339 20587
rect 24501 20553 24535 20587
rect 29469 20553 29503 20587
rect 31401 20553 31435 20587
rect 37657 20553 37691 20587
rect 5181 20485 5215 20519
rect 15761 20485 15795 20519
rect 23857 20485 23891 20519
rect 28457 20485 28491 20519
rect 1685 20417 1719 20451
rect 7113 20417 7147 20451
rect 9229 20417 9263 20451
rect 9505 20417 9539 20451
rect 11897 20417 11931 20451
rect 12725 20417 12759 20451
rect 14933 20417 14967 20451
rect 25513 20417 25547 20451
rect 30297 20417 30331 20451
rect 33057 20417 33091 20451
rect 35449 20417 35483 20451
rect 36553 20417 36587 20451
rect 1409 20349 1443 20383
rect 3065 20349 3099 20383
rect 3525 20349 3559 20383
rect 4537 20349 4571 20383
rect 4905 20349 4939 20383
rect 5273 20349 5307 20383
rect 5917 20349 5951 20383
rect 7021 20349 7055 20383
rect 7297 20349 7331 20383
rect 7665 20349 7699 20383
rect 8125 20349 8159 20383
rect 8769 20349 8803 20383
rect 11345 20349 11379 20383
rect 11437 20349 11471 20383
rect 12449 20349 12483 20383
rect 14749 20349 14783 20383
rect 14841 20349 14875 20383
rect 15485 20349 15519 20383
rect 16129 20349 16163 20383
rect 16313 20349 16347 20383
rect 17049 20349 17083 20383
rect 18613 20349 18647 20383
rect 18705 20349 18739 20383
rect 18981 20349 19015 20383
rect 20453 20349 20487 20383
rect 20821 20349 20855 20383
rect 21649 20349 21683 20383
rect 21833 20349 21867 20383
rect 22569 20349 22603 20383
rect 23489 20349 23523 20383
rect 23673 20349 23707 20383
rect 24409 20349 24443 20383
rect 25789 20349 25823 20383
rect 27629 20349 27663 20383
rect 28181 20349 28215 20383
rect 28457 20349 28491 20383
rect 29285 20349 29319 20383
rect 30021 20349 30055 20383
rect 32321 20349 32355 20383
rect 32505 20349 32539 20383
rect 32965 20349 32999 20383
rect 33977 20349 34011 20383
rect 35357 20349 35391 20383
rect 35725 20349 35759 20383
rect 36277 20349 36311 20383
rect 33793 20281 33827 20315
rect 34345 20281 34379 20315
rect 6101 20213 6135 20247
rect 17233 20213 17267 20247
rect 18429 20213 18463 20247
rect 21005 20213 21039 20247
rect 21465 20213 21499 20247
rect 22753 20213 22787 20247
rect 26893 20213 26927 20247
rect 4077 20009 4111 20043
rect 4261 20009 4295 20043
rect 11529 20009 11563 20043
rect 13461 20009 13495 20043
rect 21465 20009 21499 20043
rect 23765 20009 23799 20043
rect 25881 20009 25915 20043
rect 27169 20009 27203 20043
rect 28641 20009 28675 20043
rect 29929 20009 29963 20043
rect 30665 20009 30699 20043
rect 15301 19941 15335 19975
rect 15853 19941 15887 19975
rect 25145 19941 25179 19975
rect 32873 19941 32907 19975
rect 33425 19941 33459 19975
rect 35541 19941 35575 19975
rect 2421 19873 2455 19907
rect 3249 19873 3283 19907
rect 3433 19873 3467 19907
rect 4077 19873 4111 19907
rect 4445 19873 4479 19907
rect 4629 19873 4663 19907
rect 5181 19873 5215 19907
rect 5457 19873 5491 19907
rect 6377 19873 6411 19907
rect 6929 19873 6963 19907
rect 7573 19873 7607 19907
rect 8217 19873 8251 19907
rect 8309 19873 8343 19907
rect 9045 19873 9079 19907
rect 10149 19873 10183 19907
rect 12357 19873 12391 19907
rect 13553 19873 13587 19907
rect 14013 19873 14047 19907
rect 14197 19873 14231 19907
rect 15117 19873 15151 19907
rect 15485 19873 15519 19907
rect 16589 19873 16623 19907
rect 18981 19873 19015 19907
rect 21373 19873 21407 19907
rect 21925 19873 21959 19907
rect 22569 19873 22603 19907
rect 23029 19873 23063 19907
rect 23949 19873 23983 19907
rect 24133 19873 24167 19907
rect 24409 19873 24443 19907
rect 24961 19873 24995 19907
rect 25789 19873 25823 19907
rect 27261 19873 27295 19907
rect 27813 19873 27847 19907
rect 28089 19873 28123 19907
rect 28825 19873 28859 19907
rect 29101 19873 29135 19907
rect 29745 19873 29779 19907
rect 30481 19873 30515 19907
rect 31217 19873 31251 19907
rect 32781 19873 32815 19907
rect 32965 19873 32999 19907
rect 34161 19873 34195 19907
rect 36093 19873 36127 19907
rect 36737 19873 36771 19907
rect 36921 19873 36955 19907
rect 37749 19873 37783 19907
rect 7113 19805 7147 19839
rect 10425 19805 10459 19839
rect 12265 19805 12299 19839
rect 16313 19805 16347 19839
rect 23121 19805 23155 19839
rect 33885 19805 33919 19839
rect 3249 19737 3283 19771
rect 20269 19737 20303 19771
rect 36369 19737 36403 19771
rect 8953 19669 8987 19703
rect 12541 19669 12575 19703
rect 14933 19669 14967 19703
rect 17693 19669 17727 19703
rect 29193 19669 29227 19703
rect 31401 19669 31435 19703
rect 37841 19669 37875 19703
rect 4629 19465 4663 19499
rect 10885 19465 10919 19499
rect 27997 19465 28031 19499
rect 3985 19397 4019 19431
rect 22385 19397 22419 19431
rect 23765 19397 23799 19431
rect 30849 19397 30883 19431
rect 7389 19329 7423 19363
rect 13461 19329 13495 19363
rect 15945 19329 15979 19363
rect 20913 19329 20947 19363
rect 26801 19329 26835 19363
rect 33333 19329 33367 19363
rect 36461 19329 36495 19363
rect 2421 19261 2455 19295
rect 2697 19261 2731 19295
rect 4537 19261 4571 19295
rect 5273 19261 5307 19295
rect 5457 19261 5491 19295
rect 7021 19261 7055 19295
rect 7297 19261 7331 19295
rect 7573 19261 7607 19295
rect 8309 19261 8343 19295
rect 9045 19261 9079 19295
rect 9689 19261 9723 19295
rect 10057 19261 10091 19295
rect 10609 19261 10643 19295
rect 10701 19261 10735 19295
rect 11621 19261 11655 19295
rect 13645 19261 13679 19295
rect 14197 19261 14231 19295
rect 14381 19261 14415 19295
rect 14841 19261 14875 19295
rect 15209 19261 15243 19295
rect 15669 19261 15703 19295
rect 16405 19261 16439 19295
rect 16497 19261 16531 19295
rect 17877 19261 17911 19295
rect 18061 19261 18095 19295
rect 18153 19261 18187 19295
rect 21005 19261 21039 19295
rect 21281 19261 21315 19295
rect 22753 19261 22787 19295
rect 23673 19261 23707 19295
rect 24409 19261 24443 19295
rect 24869 19261 24903 19295
rect 25053 19261 25087 19295
rect 25329 19261 25363 19295
rect 26157 19261 26191 19295
rect 26985 19261 27019 19295
rect 27537 19261 27571 19295
rect 27721 19261 27755 19295
rect 29285 19261 29319 19295
rect 29745 19261 29779 19295
rect 31033 19261 31067 19295
rect 31401 19261 31435 19295
rect 31493 19261 31527 19295
rect 32045 19261 32079 19295
rect 32965 19261 32999 19295
rect 33149 19261 33183 19295
rect 33425 19261 33459 19295
rect 34897 19261 34931 19295
rect 35449 19261 35483 19295
rect 36737 19261 36771 19295
rect 5365 19193 5399 19227
rect 5917 19193 5951 19227
rect 16957 19193 16991 19227
rect 18613 19193 18647 19227
rect 19165 19193 19199 19227
rect 9137 19125 9171 19159
rect 11713 19125 11747 19159
rect 17693 19125 17727 19159
rect 22937 19125 22971 19159
rect 26249 19125 26283 19159
rect 29377 19125 29411 19159
rect 34989 19125 35023 19159
rect 37841 19125 37875 19159
rect 18245 18921 18279 18955
rect 37841 18921 37875 18955
rect 13553 18853 13587 18887
rect 14657 18853 14691 18887
rect 21005 18853 21039 18887
rect 28825 18853 28859 18887
rect 2329 18785 2363 18819
rect 2697 18785 2731 18819
rect 3065 18785 3099 18819
rect 3433 18785 3467 18819
rect 4077 18785 4111 18819
rect 5089 18785 5123 18819
rect 5273 18785 5307 18819
rect 5641 18785 5675 18819
rect 6101 18785 6135 18819
rect 6745 18785 6779 18819
rect 7113 18785 7147 18819
rect 7389 18785 7423 18819
rect 8401 18785 8435 18819
rect 8953 18785 8987 18819
rect 9689 18785 9723 18819
rect 10241 18785 10275 18819
rect 10793 18785 10827 18819
rect 10977 18785 11011 18819
rect 11897 18785 11931 18819
rect 12173 18785 12207 18819
rect 14013 18785 14047 18819
rect 14105 18785 14139 18819
rect 14289 18785 14323 18819
rect 15485 18785 15519 18819
rect 15853 18785 15887 18819
rect 16129 18785 16163 18819
rect 17141 18785 17175 18819
rect 19073 18785 19107 18819
rect 19717 18785 19751 18819
rect 20269 18785 20303 18819
rect 20913 18785 20947 18819
rect 21557 18785 21591 18819
rect 22385 18785 22419 18819
rect 24041 18785 24075 18819
rect 24501 18785 24535 18819
rect 24777 18785 24811 18819
rect 25145 18785 25179 18819
rect 25697 18785 25731 18819
rect 26525 18785 26559 18819
rect 29285 18785 29319 18819
rect 31401 18785 31435 18819
rect 32873 18785 32907 18819
rect 33241 18785 33275 18819
rect 33333 18785 33367 18819
rect 33885 18785 33919 18819
rect 34437 18785 34471 18819
rect 34989 18785 35023 18819
rect 35357 18785 35391 18819
rect 35541 18785 35575 18819
rect 36461 18785 36495 18819
rect 37013 18785 37047 18819
rect 37749 18785 37783 18819
rect 2881 18717 2915 18751
rect 10885 18717 10919 18751
rect 16865 18717 16899 18751
rect 18981 18717 19015 18751
rect 19625 18717 19659 18751
rect 22293 18717 22327 18751
rect 22661 18717 22695 18751
rect 27169 18717 27203 18751
rect 27445 18717 27479 18751
rect 29561 18717 29595 18751
rect 34529 18717 34563 18751
rect 4169 18649 4203 18683
rect 14013 18649 14047 18683
rect 16129 18649 16163 18683
rect 20453 18649 20487 18683
rect 23305 18649 23339 18683
rect 23397 18649 23431 18683
rect 31493 18649 31527 18683
rect 32689 18649 32723 18683
rect 6193 18581 6227 18615
rect 8309 18581 8343 18615
rect 9781 18581 9815 18615
rect 11161 18581 11195 18615
rect 19257 18581 19291 18615
rect 19901 18581 19935 18615
rect 25881 18581 25915 18615
rect 26617 18581 26651 18615
rect 30665 18581 30699 18615
rect 36553 18581 36587 18615
rect 2789 18377 2823 18411
rect 5457 18377 5491 18411
rect 6101 18377 6135 18411
rect 7573 18377 7607 18411
rect 9689 18377 9723 18411
rect 11805 18377 11839 18411
rect 12725 18377 12759 18411
rect 19717 18377 19751 18411
rect 26985 18377 27019 18411
rect 29561 18309 29595 18343
rect 37841 18309 37875 18343
rect 10517 18241 10551 18275
rect 14473 18241 14507 18275
rect 18613 18241 18647 18275
rect 20913 18241 20947 18275
rect 22109 18241 22143 18275
rect 31493 18241 31527 18275
rect 33977 18241 34011 18275
rect 35725 18241 35759 18275
rect 36737 18241 36771 18275
rect 1409 18173 1443 18207
rect 1685 18173 1719 18207
rect 4077 18173 4111 18207
rect 4721 18173 4755 18207
rect 5089 18173 5123 18207
rect 5365 18173 5399 18207
rect 6009 18173 6043 18207
rect 6837 18173 6871 18207
rect 7481 18173 7515 18207
rect 8125 18173 8159 18207
rect 8401 18173 8435 18207
rect 10241 18173 10275 18207
rect 12449 18173 12483 18207
rect 12582 18173 12616 18207
rect 13829 18173 13863 18207
rect 13921 18173 13955 18207
rect 14105 18173 14139 18207
rect 14933 18173 14967 18207
rect 15209 18173 15243 18207
rect 17233 18173 17267 18207
rect 18337 18173 18371 18207
rect 20637 18173 20671 18207
rect 21649 18173 21683 18207
rect 22569 18173 22603 18207
rect 22937 18173 22971 18207
rect 23029 18173 23063 18207
rect 23673 18173 23707 18207
rect 24409 18173 24443 18207
rect 25513 18173 25547 18207
rect 25697 18173 25731 18207
rect 25881 18173 25915 18207
rect 27169 18173 27203 18207
rect 27445 18173 27479 18207
rect 28089 18173 28123 18207
rect 29469 18173 29503 18207
rect 29837 18173 29871 18207
rect 30205 18173 30239 18207
rect 30849 18173 30883 18207
rect 32045 18173 32079 18207
rect 32229 18173 32263 18207
rect 32321 18173 32355 18207
rect 32505 18173 32539 18207
rect 32781 18173 32815 18207
rect 33425 18173 33459 18207
rect 33885 18173 33919 18207
rect 34897 18173 34931 18207
rect 35633 18173 35667 18207
rect 36461 18173 36495 18207
rect 16589 18105 16623 18139
rect 21281 18105 21315 18139
rect 25053 18105 25087 18139
rect 30941 18105 30975 18139
rect 6929 18037 6963 18071
rect 13645 18037 13679 18071
rect 17417 18037 17451 18071
rect 20453 18037 20487 18071
rect 21097 18037 21131 18071
rect 21189 18037 21223 18071
rect 23857 18037 23891 18071
rect 24501 18037 24535 18071
rect 28273 18037 28307 18071
rect 34989 18037 35023 18071
rect 3433 17833 3467 17867
rect 8769 17833 8803 17867
rect 11713 17833 11747 17867
rect 19625 17833 19659 17867
rect 21189 17833 21223 17867
rect 29837 17833 29871 17867
rect 7021 17765 7055 17799
rect 14657 17765 14691 17799
rect 23581 17765 23615 17799
rect 27077 17765 27111 17799
rect 33793 17765 33827 17799
rect 37197 17765 37231 17799
rect 4353 17697 4387 17731
rect 4813 17697 4847 17731
rect 7665 17697 7699 17731
rect 8677 17697 8711 17731
rect 10425 17697 10459 17731
rect 12541 17697 12575 17731
rect 14565 17697 14599 17731
rect 15669 17697 15703 17731
rect 16129 17697 16163 17731
rect 16865 17697 16899 17731
rect 17233 17697 17267 17731
rect 17693 17697 17727 17731
rect 18521 17697 18555 17731
rect 19441 17697 19475 17731
rect 20177 17697 20211 17731
rect 21005 17697 21039 17731
rect 22201 17697 22235 17731
rect 22569 17697 22603 17731
rect 23213 17697 23247 17731
rect 23949 17697 23983 17731
rect 24409 17697 24443 17731
rect 24685 17697 24719 17731
rect 24869 17697 24903 17731
rect 25697 17697 25731 17731
rect 26525 17697 26559 17731
rect 26709 17697 26743 17731
rect 28273 17697 28307 17731
rect 28365 17697 28399 17731
rect 28641 17697 28675 17731
rect 29653 17697 29687 17731
rect 30481 17697 30515 17731
rect 31033 17697 31067 17731
rect 31217 17697 31251 17731
rect 32137 17697 32171 17731
rect 32597 17697 32631 17731
rect 32781 17697 32815 17731
rect 32965 17697 32999 17731
rect 34621 17697 34655 17731
rect 34805 17697 34839 17731
rect 35817 17697 35851 17731
rect 37749 17697 37783 17731
rect 1869 17629 1903 17663
rect 2145 17629 2179 17663
rect 5365 17629 5399 17663
rect 5641 17629 5675 17663
rect 7573 17629 7607 17663
rect 10149 17629 10183 17663
rect 12265 17629 12299 17663
rect 15393 17629 15427 17663
rect 18429 17629 18463 17663
rect 22661 17629 22695 17663
rect 28733 17629 28767 17663
rect 30573 17629 30607 17663
rect 34345 17629 34379 17663
rect 35541 17629 35575 17663
rect 16129 17561 16163 17595
rect 17693 17561 17727 17595
rect 22017 17561 22051 17595
rect 4169 17493 4203 17527
rect 7849 17493 7883 17527
rect 13829 17493 13863 17527
rect 18705 17493 18739 17527
rect 20269 17493 20303 17527
rect 25881 17493 25915 17527
rect 27721 17493 27755 17527
rect 37841 17493 37875 17527
rect 2145 17289 2179 17323
rect 27905 17289 27939 17323
rect 28365 17289 28399 17323
rect 20453 17221 20487 17255
rect 24869 17221 24903 17255
rect 25881 17221 25915 17255
rect 35173 17221 35207 17255
rect 2789 17153 2823 17187
rect 10701 17153 10735 17187
rect 14565 17153 14599 17187
rect 15117 17153 15151 17187
rect 15393 17153 15427 17187
rect 18613 17153 18647 17187
rect 29469 17153 29503 17187
rect 34069 17153 34103 17187
rect 36737 17153 36771 17187
rect 37841 17153 37875 17187
rect 2053 17085 2087 17119
rect 2881 17085 2915 17119
rect 3341 17085 3375 17119
rect 3709 17085 3743 17119
rect 4997 17085 5031 17119
rect 5365 17085 5399 17119
rect 5733 17085 5767 17119
rect 7021 17085 7055 17119
rect 7757 17085 7791 17119
rect 8033 17085 8067 17119
rect 9873 17085 9907 17119
rect 10425 17085 10459 17119
rect 10793 17085 10827 17119
rect 12817 17085 12851 17119
rect 13645 17085 13679 17119
rect 13829 17085 13863 17119
rect 14289 17085 14323 17119
rect 17233 17085 17267 17119
rect 18061 17085 18095 17119
rect 18153 17085 18187 17119
rect 19073 17085 19107 17119
rect 19349 17085 19383 17119
rect 21189 17085 21223 17119
rect 21925 17085 21959 17119
rect 22017 17085 22051 17119
rect 22569 17085 22603 17119
rect 23489 17085 23523 17119
rect 23949 17085 23983 17119
rect 24501 17085 24535 17119
rect 24869 17085 24903 17119
rect 25789 17085 25823 17119
rect 26157 17085 26191 17119
rect 26525 17085 26559 17119
rect 26709 17085 26743 17119
rect 27169 17085 27203 17119
rect 28181 17085 28215 17119
rect 29929 17085 29963 17119
rect 30113 17085 30147 17119
rect 30389 17085 30423 17119
rect 30481 17085 30515 17119
rect 30757 17085 30791 17119
rect 31401 17085 31435 17119
rect 31769 17085 31803 17119
rect 32137 17085 32171 17119
rect 33425 17085 33459 17119
rect 33793 17085 33827 17119
rect 35081 17085 35115 17119
rect 35633 17085 35667 17119
rect 35817 17085 35851 17119
rect 36461 17085 36495 17119
rect 5917 17017 5951 17051
rect 28089 17017 28123 17051
rect 32597 17017 32631 17051
rect 7205 16949 7239 16983
rect 9321 16949 9355 16983
rect 12909 16949 12943 16983
rect 16497 16949 16531 16983
rect 17417 16949 17451 16983
rect 21281 16949 21315 16983
rect 23305 16949 23339 16983
rect 33333 16949 33367 16983
rect 2973 16745 3007 16779
rect 7941 16745 7975 16779
rect 8953 16745 8987 16779
rect 25789 16745 25823 16779
rect 35909 16745 35943 16779
rect 36829 16745 36863 16779
rect 10241 16677 10275 16711
rect 29837 16677 29871 16711
rect 1685 16609 1719 16643
rect 4169 16609 4203 16643
rect 5549 16609 5583 16643
rect 6009 16609 6043 16643
rect 6469 16609 6503 16643
rect 7021 16609 7055 16643
rect 7665 16609 7699 16643
rect 8217 16609 8251 16643
rect 8861 16609 8895 16643
rect 9781 16609 9815 16643
rect 10977 16609 11011 16643
rect 11437 16609 11471 16643
rect 11805 16609 11839 16643
rect 12725 16609 12759 16643
rect 13001 16609 13035 16643
rect 14381 16609 14415 16643
rect 16129 16609 16163 16643
rect 16405 16609 16439 16643
rect 17325 16609 17359 16643
rect 19165 16609 19199 16643
rect 19809 16609 19843 16643
rect 20177 16609 20211 16643
rect 21097 16609 21131 16643
rect 21557 16609 21591 16643
rect 21833 16609 21867 16643
rect 21925 16609 21959 16643
rect 22201 16609 22235 16643
rect 22477 16609 22511 16643
rect 23213 16609 23247 16643
rect 23673 16609 23707 16643
rect 24133 16609 24167 16643
rect 24685 16609 24719 16643
rect 24869 16609 24903 16643
rect 25605 16609 25639 16643
rect 26525 16609 26559 16643
rect 27353 16609 27387 16643
rect 27813 16609 27847 16643
rect 29285 16609 29319 16643
rect 29653 16609 29687 16643
rect 31125 16609 31159 16643
rect 31585 16609 31619 16643
rect 32321 16609 32355 16643
rect 32873 16609 32907 16643
rect 33149 16609 33183 16643
rect 33793 16609 33827 16643
rect 34529 16609 34563 16643
rect 34805 16609 34839 16643
rect 36645 16609 36679 16643
rect 37749 16609 37783 16643
rect 1409 16541 1443 16575
rect 4077 16541 4111 16575
rect 5457 16541 5491 16575
rect 7113 16541 7147 16575
rect 9689 16541 9723 16575
rect 11069 16541 11103 16575
rect 17049 16541 17083 16575
rect 28181 16541 28215 16575
rect 28917 16541 28951 16575
rect 31217 16541 31251 16575
rect 33333 16541 33367 16575
rect 15945 16473 15979 16507
rect 23305 16473 23339 16507
rect 27445 16473 27479 16507
rect 33977 16473 34011 16507
rect 4353 16405 4387 16439
rect 18613 16405 18647 16439
rect 19257 16405 19291 16439
rect 26617 16405 26651 16439
rect 37933 16405 37967 16439
rect 3525 16201 3559 16235
rect 5641 16201 5675 16235
rect 8401 16201 8435 16235
rect 11161 16201 11195 16235
rect 11805 16201 11839 16235
rect 15209 16201 15243 16235
rect 18245 16201 18279 16235
rect 24133 16201 24167 16235
rect 25881 16201 25915 16235
rect 32689 16201 32723 16235
rect 36553 16201 36587 16235
rect 30205 16133 30239 16167
rect 4261 16065 4295 16099
rect 7113 16065 7147 16099
rect 9873 16065 9907 16099
rect 18797 16065 18831 16099
rect 22293 16065 22327 16099
rect 24777 16065 24811 16099
rect 25145 16065 25179 16099
rect 29469 16065 29503 16099
rect 33977 16065 34011 16099
rect 34989 16065 35023 16099
rect 36001 16065 36035 16099
rect 1961 15997 1995 16031
rect 2237 15997 2271 16031
rect 4537 15997 4571 16031
rect 6837 15997 6871 16031
rect 9597 15997 9631 16031
rect 11713 15997 11747 16031
rect 12725 15997 12759 16031
rect 13645 15997 13679 16031
rect 13921 15997 13955 16031
rect 15761 15997 15795 16031
rect 16037 15997 16071 16031
rect 18061 15997 18095 16031
rect 19073 15997 19107 16031
rect 20913 15997 20947 16031
rect 21005 15997 21039 16031
rect 21465 15997 21499 16031
rect 22017 15997 22051 16031
rect 22477 15997 22511 16031
rect 24685 15997 24719 16031
rect 25053 15997 25087 16031
rect 25789 15997 25823 16031
rect 26433 15997 26467 16031
rect 27445 15997 27479 16031
rect 27629 15997 27663 16031
rect 28457 15997 28491 16031
rect 29745 15997 29779 16031
rect 30113 15997 30147 16031
rect 31125 15997 31159 16031
rect 31401 15997 31435 16031
rect 33333 15997 33367 16031
rect 33793 15997 33827 16031
rect 35541 15997 35575 16031
rect 35817 15997 35851 16031
rect 36737 15997 36771 16031
rect 37013 15997 37047 16031
rect 37197 15997 37231 16031
rect 20453 15929 20487 15963
rect 12909 15861 12943 15895
rect 17141 15861 17175 15895
rect 26617 15861 26651 15895
rect 27261 15861 27295 15895
rect 28641 15861 28675 15895
rect 2697 15657 2731 15691
rect 4445 15657 4479 15691
rect 5549 15657 5583 15691
rect 7665 15657 7699 15691
rect 15945 15657 15979 15691
rect 19073 15657 19107 15691
rect 29745 15657 29779 15691
rect 32229 15657 32263 15691
rect 36921 15589 36955 15623
rect 2881 15521 2915 15555
rect 3157 15521 3191 15555
rect 4169 15521 4203 15555
rect 4721 15521 4755 15555
rect 5365 15521 5399 15555
rect 11161 15521 11195 15555
rect 13645 15521 13679 15555
rect 13921 15521 13955 15555
rect 14197 15521 14231 15555
rect 15853 15521 15887 15555
rect 16681 15521 16715 15555
rect 16957 15521 16991 15555
rect 17509 15521 17543 15555
rect 17877 15521 17911 15555
rect 18153 15521 18187 15555
rect 18981 15521 19015 15555
rect 19901 15521 19935 15555
rect 20085 15521 20119 15555
rect 21189 15521 21223 15555
rect 21741 15521 21775 15555
rect 23213 15521 23247 15555
rect 23581 15521 23615 15555
rect 24133 15521 24167 15555
rect 25421 15521 25455 15555
rect 25789 15521 25823 15555
rect 25881 15521 25915 15555
rect 27077 15521 27111 15555
rect 27261 15521 27295 15555
rect 27445 15521 27479 15555
rect 27629 15521 27663 15555
rect 27813 15521 27847 15555
rect 28549 15521 28583 15555
rect 29009 15521 29043 15555
rect 29377 15521 29411 15555
rect 29745 15521 29779 15555
rect 30849 15521 30883 15555
rect 31309 15521 31343 15555
rect 32137 15521 32171 15555
rect 33057 15521 33091 15555
rect 33149 15521 33183 15555
rect 33701 15521 33735 15555
rect 34069 15521 34103 15555
rect 34713 15521 34747 15555
rect 35725 15521 35759 15555
rect 36369 15521 36403 15555
rect 36645 15521 36679 15555
rect 37197 15521 37231 15555
rect 37749 15521 37783 15555
rect 6285 15453 6319 15487
rect 6561 15453 6595 15487
rect 11437 15453 11471 15487
rect 14013 15453 14047 15487
rect 20177 15453 20211 15487
rect 21833 15453 21867 15487
rect 24961 15453 24995 15487
rect 31401 15453 31435 15487
rect 33333 15453 33367 15487
rect 16589 15385 16623 15419
rect 21649 15385 21683 15419
rect 23029 15385 23063 15419
rect 34897 15385 34931 15419
rect 12541 15317 12575 15351
rect 24317 15317 24351 15351
rect 26617 15317 26651 15351
rect 37933 15317 37967 15351
rect 2421 15113 2455 15147
rect 6193 15113 6227 15147
rect 18153 15113 18187 15147
rect 20545 15113 20579 15147
rect 37841 15113 37875 15147
rect 11805 15045 11839 15079
rect 13277 15045 13311 15079
rect 29745 15045 29779 15079
rect 35725 15045 35759 15079
rect 3893 14977 3927 15011
rect 5457 14977 5491 15011
rect 10517 14977 10551 15011
rect 15301 14977 15335 15011
rect 16129 14977 16163 15011
rect 19257 14977 19291 15011
rect 25973 14977 26007 15011
rect 30297 14977 30331 15011
rect 33885 14977 33919 15011
rect 35081 14977 35115 15011
rect 36737 14977 36771 15011
rect 2145 14909 2179 14943
rect 2237 14909 2271 14943
rect 3249 14909 3283 14943
rect 4169 14909 4203 14943
rect 6009 14909 6043 14943
rect 6837 14909 6871 14943
rect 7757 14909 7791 14943
rect 8033 14909 8067 14943
rect 9873 14909 9907 14943
rect 10241 14909 10275 14943
rect 10885 14909 10919 14943
rect 11621 14909 11655 14943
rect 12541 14909 12575 14943
rect 12817 14909 12851 14943
rect 13277 14909 13311 14943
rect 14013 14909 14047 14943
rect 15209 14909 15243 14943
rect 15853 14909 15887 14943
rect 18061 14909 18095 14943
rect 18705 14909 18739 14943
rect 19165 14909 19199 14943
rect 20361 14909 20395 14943
rect 21557 14909 21591 14943
rect 21741 14909 21775 14943
rect 22017 14909 22051 14943
rect 22109 14909 22143 14943
rect 22477 14909 22511 14943
rect 23673 14909 23707 14943
rect 24501 14909 24535 14943
rect 25329 14909 25363 14943
rect 25697 14909 25731 14943
rect 26065 14909 26099 14943
rect 26985 14909 27019 14943
rect 27445 14909 27479 14943
rect 27813 14909 27847 14943
rect 28181 14909 28215 14943
rect 29561 14909 29595 14943
rect 30573 14909 30607 14943
rect 33149 14909 33183 14943
rect 33517 14909 33551 14943
rect 33793 14909 33827 14943
rect 34161 14909 34195 14943
rect 35449 14909 35483 14943
rect 35725 14909 35759 14943
rect 36461 14909 36495 14943
rect 3341 14841 3375 14875
rect 9413 14841 9447 14875
rect 17509 14841 17543 14875
rect 21097 14841 21131 14875
rect 24593 14841 24627 14875
rect 7021 14773 7055 14807
rect 14197 14773 14231 14807
rect 23857 14773 23891 14807
rect 28181 14773 28215 14807
rect 31677 14773 31711 14807
rect 2789 14569 2823 14603
rect 26985 14569 27019 14603
rect 28733 14569 28767 14603
rect 30573 14569 30607 14603
rect 32873 14569 32907 14603
rect 37841 14569 37875 14603
rect 12449 14501 12483 14535
rect 20913 14501 20947 14535
rect 3893 14433 3927 14467
rect 4537 14433 4571 14467
rect 4813 14433 4847 14467
rect 5365 14433 5399 14467
rect 5733 14433 5767 14467
rect 6285 14433 6319 14467
rect 7297 14433 7331 14467
rect 8585 14433 8619 14467
rect 8953 14433 8987 14467
rect 9137 14433 9171 14467
rect 10241 14433 10275 14467
rect 10517 14433 10551 14467
rect 11345 14433 11379 14467
rect 11897 14433 11931 14467
rect 11989 14433 12023 14467
rect 13461 14433 13495 14467
rect 14013 14433 14047 14467
rect 15761 14433 15795 14467
rect 16129 14433 16163 14467
rect 16865 14433 16899 14467
rect 17517 14433 17551 14467
rect 18429 14433 18463 14467
rect 19073 14433 19107 14467
rect 19165 14433 19199 14467
rect 19809 14433 19843 14467
rect 20085 14433 20119 14467
rect 21465 14433 21499 14467
rect 21649 14433 21683 14467
rect 21833 14433 21867 14467
rect 22017 14433 22051 14467
rect 22293 14433 22327 14467
rect 23305 14433 23339 14467
rect 23489 14433 23523 14467
rect 23673 14433 23707 14467
rect 23857 14433 23891 14467
rect 24133 14433 24167 14467
rect 24777 14433 24811 14467
rect 25513 14433 25547 14467
rect 27169 14433 27203 14467
rect 27353 14433 27387 14467
rect 27721 14433 27755 14467
rect 28917 14433 28951 14467
rect 29469 14433 29503 14467
rect 29653 14433 29687 14467
rect 29837 14433 29871 14467
rect 30757 14433 30791 14467
rect 30941 14433 30975 14467
rect 32689 14433 32723 14467
rect 33425 14433 33459 14467
rect 34437 14433 34471 14467
rect 34621 14433 34655 14467
rect 35081 14433 35115 14467
rect 36277 14433 36311 14467
rect 36461 14433 36495 14467
rect 36645 14433 36679 14467
rect 37749 14433 37783 14467
rect 1409 14365 1443 14399
rect 1685 14365 1719 14399
rect 4445 14365 4479 14399
rect 8217 14365 8251 14399
rect 9873 14365 9907 14399
rect 13185 14365 13219 14399
rect 15485 14365 15519 14399
rect 19441 14365 19475 14399
rect 22845 14365 22879 14399
rect 25789 14365 25823 14399
rect 10517 14297 10551 14331
rect 13921 14297 13955 14331
rect 16129 14297 16163 14331
rect 17601 14297 17635 14331
rect 24869 14297 24903 14331
rect 29285 14297 29319 14331
rect 35081 14297 35115 14331
rect 36093 14297 36127 14331
rect 3709 14229 3743 14263
rect 7481 14229 7515 14263
rect 16957 14229 16991 14263
rect 33609 14229 33643 14263
rect 10517 14025 10551 14059
rect 16313 14025 16347 14059
rect 21557 14025 21591 14059
rect 28641 14025 28675 14059
rect 34345 14025 34379 14059
rect 8033 13957 8067 13991
rect 13277 13957 13311 13991
rect 17049 13957 17083 13991
rect 19441 13957 19475 13991
rect 26801 13957 26835 13991
rect 1869 13889 1903 13923
rect 2145 13889 2179 13923
rect 4077 13889 4111 13923
rect 8861 13889 8895 13923
rect 12633 13889 12667 13923
rect 14289 13889 14323 13923
rect 15393 13889 15427 13923
rect 18061 13889 18095 13923
rect 20453 13889 20487 13923
rect 22385 13889 22419 13923
rect 23673 13889 23707 13923
rect 24409 13889 24443 13923
rect 27537 13889 27571 13923
rect 29745 13889 29779 13923
rect 33241 13889 33275 13923
rect 35449 13889 35483 13923
rect 37841 13889 37875 13923
rect 3985 13821 4019 13855
rect 4629 13821 4663 13855
rect 4997 13821 5031 13855
rect 5365 13821 5399 13855
rect 5917 13821 5951 13855
rect 7389 13821 7423 13855
rect 7757 13821 7791 13855
rect 8125 13821 8159 13855
rect 9045 13821 9079 13855
rect 9413 13821 9447 13855
rect 9689 13821 9723 13855
rect 10701 13821 10735 13855
rect 11069 13821 11103 13855
rect 11161 13821 11195 13855
rect 12817 13821 12851 13855
rect 13369 13821 13403 13855
rect 14013 13821 14047 13855
rect 16129 13821 16163 13855
rect 16865 13821 16899 13855
rect 18337 13821 18371 13855
rect 20177 13821 20211 13855
rect 23121 13821 23155 13855
rect 23949 13821 23983 13855
rect 25053 13821 25087 13855
rect 25237 13821 25271 13855
rect 25697 13821 25731 13855
rect 26157 13821 26191 13855
rect 26709 13821 26743 13855
rect 27261 13821 27295 13855
rect 28457 13821 28491 13855
rect 29561 13821 29595 13855
rect 29837 13821 29871 13855
rect 30205 13821 30239 13855
rect 30481 13821 30515 13855
rect 31217 13821 31251 13855
rect 32137 13821 32171 13855
rect 32597 13821 32631 13855
rect 32781 13821 32815 13855
rect 33333 13821 33367 13855
rect 33885 13821 33919 13855
rect 34529 13821 34563 13855
rect 35541 13821 35575 13855
rect 36001 13821 36035 13855
rect 36461 13821 36495 13855
rect 36737 13821 36771 13855
rect 22661 13753 22695 13787
rect 22753 13753 22787 13787
rect 24041 13753 24075 13787
rect 3433 13685 3467 13719
rect 22569 13685 22603 13719
rect 23857 13685 23891 13719
rect 24869 13685 24903 13719
rect 25237 13685 25271 13719
rect 31401 13685 31435 13719
rect 31953 13685 31987 13719
rect 1685 13481 1719 13515
rect 11069 13481 11103 13515
rect 14657 13481 14691 13515
rect 19073 13481 19107 13515
rect 23489 13481 23523 13515
rect 24225 13481 24259 13515
rect 28365 13481 28399 13515
rect 35449 13481 35483 13515
rect 1777 13345 1811 13379
rect 2145 13345 2179 13379
rect 3341 13345 3375 13379
rect 4077 13345 4111 13379
rect 4721 13345 4755 13379
rect 5365 13345 5399 13379
rect 6101 13345 6135 13379
rect 8677 13345 8711 13379
rect 9689 13345 9723 13379
rect 9965 13345 9999 13379
rect 12449 13345 12483 13379
rect 14473 13345 14507 13379
rect 14565 13345 14599 13379
rect 15301 13345 15335 13379
rect 16037 13345 16071 13379
rect 16773 13345 16807 13379
rect 17233 13345 17267 13379
rect 17417 13345 17451 13379
rect 17877 13345 17911 13379
rect 18245 13345 18279 13379
rect 18981 13345 19015 13379
rect 19625 13345 19659 13379
rect 20085 13345 20119 13379
rect 21925 13345 21959 13379
rect 22109 13345 22143 13379
rect 22201 13345 22235 13379
rect 22477 13345 22511 13379
rect 22753 13345 22787 13379
rect 23305 13345 23339 13379
rect 24041 13345 24075 13379
rect 25053 13345 25087 13379
rect 25513 13345 25547 13379
rect 25697 13345 25731 13379
rect 27077 13345 27111 13379
rect 27353 13345 27387 13379
rect 28181 13345 28215 13379
rect 29101 13345 29135 13379
rect 29377 13345 29411 13379
rect 29929 13345 29963 13379
rect 30205 13345 30239 13379
rect 30665 13345 30699 13379
rect 31309 13345 31343 13379
rect 32229 13345 32263 13379
rect 32597 13345 32631 13379
rect 33057 13345 33091 13379
rect 33977 13345 34011 13379
rect 37013 13345 37047 13379
rect 37749 13345 37783 13379
rect 3433 13277 3467 13311
rect 6377 13277 6411 13311
rect 7481 13277 7515 13311
rect 12173 13277 12207 13311
rect 17601 13277 17635 13311
rect 20361 13277 20395 13311
rect 21373 13277 21407 13311
rect 26709 13277 26743 13311
rect 29837 13277 29871 13311
rect 34069 13277 34103 13311
rect 34345 13277 34379 13311
rect 36185 13277 36219 13311
rect 36737 13277 36771 13311
rect 37197 13277 37231 13311
rect 4813 13209 4847 13243
rect 14289 13209 14323 13243
rect 24961 13209 24995 13243
rect 27353 13209 27387 13243
rect 33057 13209 33091 13243
rect 4169 13141 4203 13175
rect 5549 13141 5583 13175
rect 8861 13141 8895 13175
rect 13737 13141 13771 13175
rect 15393 13141 15427 13175
rect 31493 13141 31527 13175
rect 33793 13141 33827 13175
rect 37933 13141 37967 13175
rect 22293 12937 22327 12971
rect 6929 12869 6963 12903
rect 16681 12869 16715 12903
rect 30941 12869 30975 12903
rect 33517 12869 33551 12903
rect 1685 12801 1719 12835
rect 1961 12801 1995 12835
rect 3893 12801 3927 12835
rect 9597 12801 9631 12835
rect 11161 12801 11195 12835
rect 13461 12801 13495 12835
rect 15853 12801 15887 12835
rect 18797 12801 18831 12835
rect 19901 12801 19935 12835
rect 23949 12801 23983 12835
rect 26709 12801 26743 12835
rect 32413 12801 32447 12835
rect 35173 12801 35207 12835
rect 35725 12801 35759 12835
rect 3985 12733 4019 12767
rect 4445 12733 4479 12767
rect 4813 12733 4847 12767
rect 5181 12733 5215 12767
rect 5733 12733 5767 12767
rect 6653 12733 6687 12767
rect 7021 12733 7055 12767
rect 7297 12733 7331 12767
rect 7573 12733 7607 12767
rect 8033 12733 8067 12767
rect 8769 12733 8803 12767
rect 9413 12733 9447 12767
rect 9781 12733 9815 12767
rect 10609 12733 10643 12767
rect 10977 12733 11011 12767
rect 11253 12733 11287 12767
rect 11437 12733 11471 12767
rect 12909 12733 12943 12767
rect 13185 12733 13219 12767
rect 13369 12733 13403 12767
rect 14933 12733 14967 12767
rect 15209 12733 15243 12767
rect 15669 12733 15703 12767
rect 16405 12733 16439 12767
rect 16957 12733 16991 12767
rect 17417 12733 17451 12767
rect 18061 12733 18095 12767
rect 18705 12733 18739 12767
rect 19349 12733 19383 12767
rect 19993 12733 20027 12767
rect 20361 12733 20395 12767
rect 20545 12733 20579 12767
rect 21005 12733 21039 12767
rect 22109 12733 22143 12767
rect 22845 12733 22879 12767
rect 23673 12733 23707 12767
rect 26065 12733 26099 12767
rect 26617 12733 26651 12767
rect 27077 12733 27111 12767
rect 27261 12733 27295 12767
rect 27813 12733 27847 12767
rect 28273 12733 28307 12767
rect 29377 12733 29411 12767
rect 29929 12733 29963 12767
rect 30113 12733 30147 12767
rect 31125 12733 31159 12767
rect 31401 12733 31435 12767
rect 32229 12733 32263 12767
rect 32781 12733 32815 12767
rect 33241 12733 33275 12767
rect 33793 12733 33827 12767
rect 34253 12733 34287 12767
rect 35265 12733 35299 12767
rect 36185 12733 36219 12767
rect 36461 12733 36495 12767
rect 3341 12665 3375 12699
rect 25329 12665 25363 12699
rect 6469 12597 6503 12631
rect 10425 12597 10459 12631
rect 18153 12597 18187 12631
rect 23029 12597 23063 12631
rect 25881 12597 25915 12631
rect 29377 12597 29411 12631
rect 37565 12597 37599 12631
rect 15577 12393 15611 12427
rect 20729 12393 20763 12427
rect 23213 12393 23247 12427
rect 1409 12257 1443 12291
rect 4353 12257 4387 12291
rect 4721 12257 4755 12291
rect 5273 12257 5307 12291
rect 6101 12257 6135 12291
rect 6561 12257 6595 12291
rect 6837 12257 6871 12291
rect 7297 12257 7331 12291
rect 7849 12257 7883 12291
rect 8585 12257 8619 12291
rect 9045 12257 9079 12291
rect 9965 12257 9999 12291
rect 12081 12257 12115 12291
rect 12725 12257 12759 12291
rect 13185 12257 13219 12291
rect 13737 12257 13771 12291
rect 14381 12257 14415 12291
rect 15669 12257 15703 12291
rect 16221 12257 16255 12291
rect 17693 12257 17727 12291
rect 18061 12257 18095 12291
rect 18245 12257 18279 12291
rect 19349 12257 19383 12291
rect 19717 12257 19751 12291
rect 19809 12257 19843 12291
rect 1685 12189 1719 12223
rect 4445 12189 4479 12223
rect 5365 12189 5399 12223
rect 10241 12189 10275 12223
rect 13369 12189 13403 12223
rect 16497 12189 16531 12223
rect 17049 12189 17083 12223
rect 17785 12189 17819 12223
rect 19257 12189 19291 12223
rect 6009 12121 6043 12155
rect 27077 12325 27111 12359
rect 27445 12325 27479 12359
rect 29377 12325 29411 12359
rect 32321 12325 32355 12359
rect 32505 12325 32539 12359
rect 21189 12257 21223 12291
rect 23029 12257 23063 12291
rect 24041 12257 24075 12291
rect 27261 12257 27295 12291
rect 27353 12257 27387 12291
rect 28825 12257 28859 12291
rect 29101 12257 29135 12291
rect 29837 12257 29871 12291
rect 30849 12257 30883 12291
rect 31309 12257 31343 12291
rect 32413 12257 32447 12291
rect 33977 12257 34011 12291
rect 34345 12257 34379 12291
rect 36829 12257 36863 12291
rect 37749 12257 37783 12291
rect 20913 12189 20947 12223
rect 23765 12189 23799 12223
rect 27813 12189 27847 12223
rect 28365 12189 28399 12223
rect 30573 12189 30607 12223
rect 31585 12189 31619 12223
rect 32137 12189 32171 12223
rect 32873 12189 32907 12223
rect 33517 12189 33551 12223
rect 35173 12189 35207 12223
rect 35449 12189 35483 12223
rect 37841 12189 37875 12223
rect 34253 12121 34287 12155
rect 2789 12053 2823 12087
rect 8401 12053 8435 12087
rect 11345 12053 11379 12087
rect 12173 12053 12207 12087
rect 14565 12053 14599 12087
rect 18797 12053 18831 12087
rect 20729 12053 20763 12087
rect 22293 12053 22327 12087
rect 25329 12053 25363 12087
rect 29929 12053 29963 12087
rect 4261 11849 4295 11883
rect 8125 11849 8159 11883
rect 18889 11849 18923 11883
rect 20913 11849 20947 11883
rect 37841 11849 37875 11883
rect 6929 11781 6963 11815
rect 10885 11781 10919 11815
rect 12817 11781 12851 11815
rect 16589 11781 16623 11815
rect 32781 11781 32815 11815
rect 33149 11781 33183 11815
rect 2973 11713 3007 11747
rect 8953 11713 8987 11747
rect 14473 11713 14507 11747
rect 17325 11713 17359 11747
rect 19809 11713 19843 11747
rect 22017 11713 22051 11747
rect 24593 11713 24627 11747
rect 25237 11713 25271 11747
rect 33793 11713 33827 11747
rect 35725 11713 35759 11747
rect 1777 11645 1811 11679
rect 2053 11645 2087 11679
rect 2697 11645 2731 11679
rect 4813 11645 4847 11679
rect 5273 11645 5307 11679
rect 5549 11645 5583 11679
rect 7113 11645 7147 11679
rect 7389 11645 7423 11679
rect 8309 11645 8343 11679
rect 8401 11645 8435 11679
rect 8769 11645 8803 11679
rect 9137 11645 9171 11679
rect 10057 11645 10091 11679
rect 10425 11645 10459 11679
rect 10977 11645 11011 11679
rect 11621 11645 11655 11679
rect 13001 11645 13035 11679
rect 13185 11645 13219 11679
rect 13369 11645 13403 11679
rect 14289 11645 14323 11679
rect 14657 11645 14691 11679
rect 15117 11645 15151 11679
rect 16405 11645 16439 11679
rect 16865 11645 16899 11679
rect 18061 11645 18095 11679
rect 18797 11645 18831 11679
rect 19533 11645 19567 11679
rect 22109 11645 22143 11679
rect 24133 11645 24167 11679
rect 24409 11645 24443 11679
rect 26709 11645 26743 11679
rect 27169 11645 27203 11679
rect 27353 11645 27387 11679
rect 27721 11645 27755 11679
rect 28089 11645 28123 11679
rect 29101 11645 29135 11679
rect 29837 11645 29871 11679
rect 30021 11645 30055 11679
rect 30205 11645 30239 11679
rect 30389 11645 30423 11679
rect 30665 11645 30699 11679
rect 31217 11645 31251 11679
rect 31585 11645 31619 11679
rect 31999 11645 32033 11679
rect 32781 11645 32815 11679
rect 32873 11645 32907 11679
rect 33425 11645 33459 11679
rect 34897 11645 34931 11679
rect 35633 11645 35667 11679
rect 36461 11645 36495 11679
rect 36737 11645 36771 11679
rect 6009 11577 6043 11611
rect 22569 11577 22603 11611
rect 25605 11577 25639 11611
rect 25973 11577 26007 11611
rect 26801 11577 26835 11611
rect 29285 11577 29319 11611
rect 32321 11577 32355 11611
rect 1593 11509 1627 11543
rect 11805 11509 11839 11543
rect 18245 11509 18279 11543
rect 25421 11509 25455 11543
rect 25513 11509 25547 11543
rect 28917 11509 28951 11543
rect 34989 11509 35023 11543
rect 5273 11305 5307 11339
rect 7573 11305 7607 11339
rect 15485 11305 15519 11339
rect 19533 11305 19567 11339
rect 22661 11305 22695 11339
rect 23581 11305 23615 11339
rect 25605 11305 25639 11339
rect 37013 11305 37047 11339
rect 17785 11237 17819 11271
rect 2421 11169 2455 11203
rect 4353 11169 4387 11203
rect 4629 11169 4663 11203
rect 5457 11169 5491 11203
rect 5825 11169 5859 11203
rect 6101 11169 6135 11203
rect 6561 11169 6595 11203
rect 7389 11169 7423 11203
rect 8585 11169 8619 11203
rect 8769 11169 8803 11203
rect 8953 11169 8987 11203
rect 10609 11169 10643 11203
rect 10977 11169 11011 11203
rect 11069 11169 11103 11203
rect 12725 11169 12759 11203
rect 13093 11169 13127 11203
rect 14197 11169 14231 11203
rect 14381 11169 14415 11203
rect 14565 11169 14599 11203
rect 15577 11169 15611 11203
rect 16037 11169 16071 11203
rect 17049 11169 17083 11203
rect 18429 11169 18463 11203
rect 18521 11169 18555 11203
rect 18797 11169 18831 11203
rect 19441 11169 19475 11203
rect 19993 11169 20027 11203
rect 21189 11169 21223 11203
rect 21833 11169 21867 11203
rect 22477 11169 22511 11203
rect 23397 11169 23431 11203
rect 24317 11169 24351 11203
rect 24685 11169 24719 11203
rect 25421 11169 25455 11203
rect 26525 11169 26559 11203
rect 28641 11169 28675 11203
rect 29193 11169 29227 11203
rect 29377 11169 29411 11203
rect 29929 11169 29963 11203
rect 31447 11169 31481 11203
rect 31585 11169 31619 11203
rect 32137 11169 32171 11203
rect 32689 11169 32723 11203
rect 33057 11169 33091 11203
rect 34069 11169 34103 11203
rect 34437 11169 34471 11203
rect 2329 11101 2363 11135
rect 2881 11101 2915 11135
rect 4445 11101 4479 11135
rect 10701 11101 10735 11135
rect 12265 11101 12299 11135
rect 16405 11101 16439 11135
rect 18889 11101 18923 11135
rect 26801 11101 26835 11135
rect 29101 11101 29135 11135
rect 30573 11101 30607 11135
rect 31125 11101 31159 11135
rect 34713 11101 34747 11135
rect 35449 11101 35483 11135
rect 35725 11101 35759 11135
rect 8401 11033 8435 11067
rect 13093 11033 13127 11067
rect 14013 11033 14047 11067
rect 17233 11033 17267 11067
rect 21281 11033 21315 11067
rect 24133 11033 24167 11067
rect 24869 11033 24903 11067
rect 27905 11033 27939 11067
rect 32229 11033 32263 11067
rect 34161 11033 34195 11067
rect 5641 10965 5675 10999
rect 10057 10965 10091 10999
rect 21925 10965 21959 10999
rect 15853 10761 15887 10795
rect 16681 10693 16715 10727
rect 18153 10693 18187 10727
rect 21189 10693 21223 10727
rect 23765 10693 23799 10727
rect 29653 10693 29687 10727
rect 31217 10693 31251 10727
rect 5273 10625 5307 10659
rect 6285 10625 6319 10659
rect 9505 10625 9539 10659
rect 14197 10625 14231 10659
rect 26801 10625 26835 10659
rect 27997 10625 28031 10659
rect 31769 10625 31803 10659
rect 35909 10625 35943 10659
rect 36461 10625 36495 10659
rect 2145 10557 2179 10591
rect 3065 10557 3099 10591
rect 3157 10557 3191 10591
rect 4353 10557 4387 10591
rect 4537 10557 4571 10591
rect 4813 10557 4847 10591
rect 5733 10557 5767 10591
rect 5825 10557 5859 10591
rect 7481 10557 7515 10591
rect 8033 10557 8067 10591
rect 8309 10557 8343 10591
rect 9413 10557 9447 10591
rect 9873 10557 9907 10591
rect 10333 10557 10367 10591
rect 10977 10557 11011 10591
rect 11069 10557 11103 10591
rect 11345 10557 11379 10591
rect 11529 10557 11563 10591
rect 12449 10557 12483 10591
rect 13001 10557 13035 10591
rect 13277 10557 13311 10591
rect 14657 10557 14691 10591
rect 15025 10557 15059 10591
rect 15117 10557 15151 10591
rect 15669 10557 15703 10591
rect 16497 10557 16531 10591
rect 16957 10557 16991 10591
rect 17417 10557 17451 10591
rect 18337 10557 18371 10591
rect 18613 10557 18647 10591
rect 19441 10557 19475 10591
rect 19993 10557 20027 10591
rect 21097 10557 21131 10591
rect 21879 10557 21913 10591
rect 22017 10557 22051 10591
rect 22385 10557 22419 10591
rect 22477 10557 22511 10591
rect 23673 10557 23707 10591
rect 24961 10557 24995 10591
rect 25697 10557 25731 10591
rect 28181 10557 28215 10591
rect 28273 10557 28307 10591
rect 29837 10557 29871 10591
rect 30021 10557 30055 10591
rect 30205 10557 30239 10591
rect 31033 10557 31067 10591
rect 32275 10557 32309 10591
rect 32597 10557 32631 10591
rect 32781 10557 32815 10591
rect 33241 10557 33275 10591
rect 33609 10557 33643 10591
rect 34069 10557 34103 10591
rect 34897 10557 34931 10591
rect 35449 10557 35483 10591
rect 36737 10557 36771 10591
rect 3617 10489 3651 10523
rect 8585 10489 8619 10523
rect 13553 10489 13587 10523
rect 23029 10489 23063 10523
rect 26249 10489 26283 10523
rect 27077 10489 27111 10523
rect 27169 10489 27203 10523
rect 27537 10489 27571 10523
rect 28365 10489 28399 10523
rect 28733 10489 28767 10523
rect 34345 10489 34379 10523
rect 38117 10489 38151 10523
rect 2329 10421 2363 10455
rect 19533 10421 19567 10455
rect 26985 10421 27019 10455
rect 34989 10421 35023 10455
rect 3157 10217 3191 10251
rect 6929 10217 6963 10251
rect 7849 10217 7883 10251
rect 37841 10217 37875 10251
rect 4813 10149 4847 10183
rect 16681 10149 16715 10183
rect 18337 10149 18371 10183
rect 33701 10149 33735 10183
rect 4261 10081 4295 10115
rect 4353 10081 4387 10115
rect 5457 10081 5491 10115
rect 7941 10081 7975 10115
rect 8493 10081 8527 10115
rect 9505 10081 9539 10115
rect 9689 10081 9723 10115
rect 10149 10081 10183 10115
rect 10333 10081 10367 10115
rect 10517 10081 10551 10115
rect 12173 10081 12207 10115
rect 12541 10081 12575 10115
rect 12725 10081 12759 10115
rect 13645 10081 13679 10115
rect 13829 10081 13863 10115
rect 14013 10081 14047 10115
rect 15761 10081 15795 10115
rect 16221 10081 16255 10115
rect 17325 10081 17359 10115
rect 17417 10081 17451 10115
rect 17693 10081 17727 10115
rect 18981 10081 19015 10115
rect 19349 10081 19383 10115
rect 19441 10081 19475 10115
rect 19993 10081 20027 10115
rect 20913 10081 20947 10115
rect 21281 10081 21315 10115
rect 21649 10081 21683 10115
rect 23305 10081 23339 10115
rect 25513 10081 25547 10115
rect 25697 10081 25731 10115
rect 26709 10081 26743 10115
rect 27629 10081 27663 10115
rect 27905 10081 27939 10115
rect 28365 10081 28399 10115
rect 28917 10081 28951 10115
rect 29193 10081 29227 10115
rect 30021 10081 30055 10115
rect 30665 10081 30699 10115
rect 31125 10081 31159 10115
rect 32965 10081 32999 10115
rect 33425 10081 33459 10115
rect 34345 10081 34379 10115
rect 34713 10081 34747 10115
rect 36553 10081 36587 10115
rect 37749 10081 37783 10115
rect 1777 10013 1811 10047
rect 2053 10013 2087 10047
rect 5549 10013 5583 10047
rect 5825 10013 5859 10047
rect 8677 10013 8711 10047
rect 12081 10013 12115 10047
rect 15669 10013 15703 10047
rect 17785 10013 17819 10047
rect 19073 10013 19107 10047
rect 21741 10013 21775 10047
rect 23029 10013 23063 10047
rect 25973 10013 26007 10047
rect 27813 10013 27847 10047
rect 30481 10013 30515 10047
rect 32781 10013 32815 10047
rect 34437 10013 34471 10047
rect 13461 9945 13495 9979
rect 31217 9945 31251 9979
rect 34161 9945 34195 9979
rect 36737 9945 36771 9979
rect 5273 9877 5307 9911
rect 9321 9877 9355 9911
rect 11621 9877 11655 9911
rect 20177 9877 20211 9911
rect 24409 9877 24443 9911
rect 26893 9877 26927 9911
rect 29837 9877 29871 9911
rect 35817 9877 35851 9911
rect 2789 9673 2823 9707
rect 15761 9673 15795 9707
rect 22017 9673 22051 9707
rect 11161 9605 11195 9639
rect 13093 9605 13127 9639
rect 20085 9605 20119 9639
rect 22937 9605 22971 9639
rect 34253 9605 34287 9639
rect 1409 9537 1443 9571
rect 9045 9537 9079 9571
rect 17509 9537 17543 9571
rect 30481 9537 30515 9571
rect 37841 9537 37875 9571
rect 1685 9469 1719 9503
rect 3525 9469 3559 9503
rect 4077 9469 4111 9503
rect 4905 9469 4939 9503
rect 5825 9469 5859 9503
rect 6101 9469 6135 9503
rect 6837 9469 6871 9503
rect 7297 9469 7331 9503
rect 8033 9469 8067 9503
rect 8677 9469 8711 9503
rect 8861 9469 8895 9503
rect 9229 9469 9263 9503
rect 9965 9469 9999 9503
rect 11345 9469 11379 9503
rect 11529 9469 11563 9503
rect 11713 9469 11747 9503
rect 12817 9469 12851 9503
rect 13553 9469 13587 9503
rect 13829 9469 13863 9503
rect 14381 9469 14415 9503
rect 14657 9469 14691 9503
rect 16773 9469 16807 9503
rect 17325 9469 17359 9503
rect 18061 9469 18095 9503
rect 18797 9469 18831 9503
rect 19349 9469 19383 9503
rect 19993 9469 20027 9503
rect 20637 9469 20671 9503
rect 20913 9469 20947 9503
rect 22753 9469 22787 9503
rect 23949 9469 23983 9503
rect 25513 9469 25547 9503
rect 25973 9469 26007 9503
rect 26525 9469 26559 9503
rect 26985 9469 27019 9503
rect 27169 9469 27203 9503
rect 27537 9469 27571 9503
rect 27721 9469 27755 9503
rect 27905 9469 27939 9503
rect 28457 9469 28491 9503
rect 29377 9469 29411 9503
rect 30113 9469 30147 9503
rect 30849 9469 30883 9503
rect 31217 9469 31251 9503
rect 31493 9469 31527 9503
rect 32045 9469 32079 9503
rect 32505 9469 32539 9503
rect 32965 9469 32999 9503
rect 33425 9469 33459 9503
rect 34069 9469 34103 9503
rect 35541 9469 35575 9503
rect 35679 9469 35713 9503
rect 35817 9469 35851 9503
rect 36461 9469 36495 9503
rect 36737 9469 36771 9503
rect 33609 9401 33643 9435
rect 34989 9401 35023 9435
rect 3617 9333 3651 9367
rect 4997 9333 5031 9367
rect 5825 9333 5859 9367
rect 7113 9333 7147 9367
rect 18245 9333 18279 9367
rect 18889 9333 18923 9367
rect 24041 9333 24075 9367
rect 29561 9333 29595 9367
rect 8033 9129 8067 9163
rect 15393 9129 15427 9163
rect 17049 9129 17083 9163
rect 24593 9129 24627 9163
rect 25881 9129 25915 9163
rect 34161 9129 34195 9163
rect 3525 9061 3559 9095
rect 9965 9061 9999 9095
rect 12357 9061 12391 9095
rect 19165 9061 19199 9095
rect 30573 9061 30607 9095
rect 35357 9061 35391 9095
rect 1869 8993 1903 9027
rect 4813 8993 4847 9027
rect 5457 8993 5491 9027
rect 5917 8993 5951 9027
rect 6469 8993 6503 9027
rect 6837 8993 6871 9027
rect 7113 8993 7147 9027
rect 8217 8993 8251 9027
rect 8677 8993 8711 9027
rect 9045 8993 9079 9027
rect 10609 8993 10643 9027
rect 10977 8993 11011 9027
rect 11621 8993 11655 9027
rect 12081 8993 12115 9027
rect 13553 8993 13587 9027
rect 13921 8993 13955 9027
rect 14013 8993 14047 9027
rect 14565 8993 14599 9027
rect 15485 8993 15519 9027
rect 15853 8993 15887 9027
rect 16313 8993 16347 9027
rect 16865 8993 16899 9027
rect 17785 8993 17819 9027
rect 18337 8993 18371 9027
rect 19809 8993 19843 9027
rect 20177 8993 20211 9027
rect 21465 8993 21499 9027
rect 21741 8993 21775 9027
rect 22477 8993 22511 9027
rect 25697 8993 25731 9027
rect 27537 8993 27571 9027
rect 27905 8993 27939 9027
rect 28641 8993 28675 9027
rect 29193 8993 29227 9027
rect 29653 8993 29687 9027
rect 29929 8993 29963 9027
rect 31401 8993 31435 9027
rect 32137 8993 32171 9027
rect 33057 8993 33091 9027
rect 36185 8993 36219 9027
rect 36829 8993 36863 9027
rect 2145 8925 2179 8959
rect 8769 8925 8803 8959
rect 10517 8925 10551 8959
rect 11069 8925 11103 8959
rect 13461 8925 13495 8959
rect 18429 8925 18463 8959
rect 19717 8925 19751 8959
rect 20269 8925 20303 8959
rect 21005 8925 21039 8959
rect 23213 8925 23247 8959
rect 23489 8925 23523 8959
rect 27261 8925 27295 8959
rect 28181 8925 28215 8959
rect 30021 8925 30055 8959
rect 31125 8925 31159 8959
rect 31585 8925 31619 8959
rect 32781 8925 32815 8959
rect 35909 8925 35943 8959
rect 36369 8925 36403 8959
rect 5549 8857 5583 8891
rect 14657 8857 14691 8891
rect 21741 8857 21775 8891
rect 32229 8857 32263 8891
rect 4905 8789 4939 8823
rect 13001 8789 13035 8823
rect 22661 8789 22695 8823
rect 37013 8789 37047 8823
rect 1777 8585 1811 8619
rect 5825 8585 5859 8619
rect 6929 8585 6963 8619
rect 10149 8585 10183 8619
rect 14013 8585 14047 8619
rect 16221 8585 16255 8619
rect 34897 8585 34931 8619
rect 37841 8585 37875 8619
rect 8309 8517 8343 8551
rect 12725 8517 12759 8551
rect 14841 8517 14875 8551
rect 19625 8517 19659 8551
rect 28641 8517 28675 8551
rect 29837 8517 29871 8551
rect 32873 8517 32907 8551
rect 1501 8449 1535 8483
rect 3065 8449 3099 8483
rect 4721 8449 4755 8483
rect 8861 8449 8895 8483
rect 11897 8449 11931 8483
rect 19073 8449 19107 8483
rect 20085 8449 20119 8483
rect 23029 8449 23063 8483
rect 24409 8449 24443 8483
rect 26801 8449 26835 8483
rect 1593 8381 1627 8415
rect 2513 8381 2547 8415
rect 2973 8381 3007 8415
rect 3801 8381 3835 8415
rect 4445 8381 4479 8415
rect 6837 8381 6871 8415
rect 7389 8381 7423 8415
rect 8493 8381 8527 8415
rect 8585 8381 8619 8415
rect 11345 8381 11379 8415
rect 11713 8381 11747 8415
rect 12909 8381 12943 8415
rect 13277 8381 13311 8415
rect 13369 8381 13403 8415
rect 13921 8381 13955 8415
rect 14749 8381 14783 8415
rect 15117 8381 15151 8415
rect 15577 8381 15611 8415
rect 16221 8381 16255 8415
rect 16681 8381 16715 8415
rect 17325 8381 17359 8415
rect 18613 8381 18647 8415
rect 18889 8381 18923 8415
rect 20177 8381 20211 8415
rect 20545 8381 20579 8415
rect 20729 8381 20763 8415
rect 21925 8381 21959 8415
rect 22017 8381 22051 8415
rect 22385 8381 22419 8415
rect 22477 8381 22511 8415
rect 24133 8381 24167 8415
rect 27077 8381 27111 8415
rect 27261 8381 27295 8415
rect 27629 8381 27663 8415
rect 27813 8381 27847 8415
rect 28457 8381 28491 8415
rect 30021 8381 30055 8415
rect 30389 8381 30423 8415
rect 30481 8381 30515 8415
rect 31033 8381 31067 8415
rect 31585 8381 31619 8415
rect 32045 8381 32079 8415
rect 32781 8381 32815 8415
rect 33149 8381 33183 8415
rect 33425 8381 33459 8415
rect 34161 8381 34195 8415
rect 34989 8449 35023 8483
rect 36737 8449 36771 8483
rect 35541 8381 35575 8415
rect 35679 8381 35713 8415
rect 35817 8381 35851 8415
rect 36461 8381 36495 8415
rect 3893 8313 3927 8347
rect 25789 8313 25823 8347
rect 34253 8313 34287 8347
rect 34897 8313 34931 8347
rect 17417 8245 17451 8279
rect 31125 8245 31159 8279
rect 2789 8041 2823 8075
rect 8953 8041 8987 8075
rect 9505 8041 9539 8075
rect 11713 8041 11747 8075
rect 14105 8041 14139 8075
rect 20085 8041 20119 8075
rect 21005 8041 21039 8075
rect 23489 8041 23523 8075
rect 30113 8041 30147 8075
rect 31033 8041 31067 8075
rect 31125 8041 31159 8075
rect 32321 8041 32355 8075
rect 34897 8041 34931 8075
rect 1409 7905 1443 7939
rect 4537 7905 4571 7939
rect 4997 7905 5031 7939
rect 5641 7905 5675 7939
rect 6561 7905 6595 7939
rect 6929 7905 6963 7939
rect 7297 7905 7331 7939
rect 7757 7905 7791 7939
rect 8309 7905 8343 7939
rect 8769 7905 8803 7939
rect 1685 7837 1719 7871
rect 6745 7837 6779 7871
rect 4353 7769 4387 7803
rect 5825 7769 5859 7803
rect 18245 7973 18279 8007
rect 30849 7973 30883 8007
rect 31217 7973 31251 8007
rect 31585 7973 31619 8007
rect 10517 7905 10551 7939
rect 10701 7905 10735 7939
rect 10977 7905 11011 7939
rect 11529 7905 11563 7939
rect 13001 7905 13035 7939
rect 13277 7905 13311 7939
rect 14197 7905 14231 7939
rect 14473 7905 14507 7939
rect 15853 7905 15887 7939
rect 16313 7905 16347 7939
rect 16497 7905 16531 7939
rect 16865 7905 16899 7939
rect 17601 7905 17635 7939
rect 18889 7905 18923 7939
rect 18981 7905 19015 7939
rect 19257 7905 19291 7939
rect 19901 7905 19935 7939
rect 20913 7905 20947 7939
rect 21465 7905 21499 7939
rect 22477 7905 22511 7939
rect 23029 7905 23063 7939
rect 23213 7905 23247 7939
rect 24409 7905 24443 7939
rect 24501 7905 24535 7939
rect 25145 7905 25179 7939
rect 25789 7905 25823 7939
rect 26801 7905 26835 7939
rect 27445 7905 27479 7939
rect 27813 7905 27847 7939
rect 27997 7905 28031 7939
rect 29009 7905 29043 7939
rect 32137 7905 32171 7939
rect 33425 7905 33459 7939
rect 33885 7905 33919 7939
rect 34253 7905 34287 7939
rect 34805 7905 34839 7939
rect 35357 7905 35391 7939
rect 36369 7905 36403 7939
rect 12541 7837 12575 7871
rect 13369 7837 13403 7871
rect 19349 7837 19383 7871
rect 22293 7837 22327 7871
rect 27169 7837 27203 7871
rect 28733 7837 28767 7871
rect 35633 7837 35667 7871
rect 15761 7769 15795 7803
rect 33333 7769 33367 7803
rect 9505 7701 9539 7735
rect 24225 7701 24259 7735
rect 25881 7701 25915 7735
rect 36461 7701 36495 7735
rect 4169 7497 4203 7531
rect 7297 7497 7331 7531
rect 16865 7497 16899 7531
rect 25881 7497 25915 7531
rect 32505 7497 32539 7531
rect 37841 7497 37875 7531
rect 10425 7429 10459 7463
rect 13645 7429 13679 7463
rect 33425 7429 33459 7463
rect 5089 7361 5123 7395
rect 7941 7361 7975 7395
rect 10885 7361 10919 7395
rect 11805 7361 11839 7395
rect 14565 7361 14599 7395
rect 15301 7361 15335 7395
rect 15577 7361 15611 7395
rect 19165 7361 19199 7395
rect 19901 7361 19935 7395
rect 22201 7361 22235 7395
rect 26893 7361 26927 7395
rect 30941 7361 30975 7395
rect 31217 7361 31251 7395
rect 34161 7361 34195 7395
rect 35541 7361 35575 7395
rect 36001 7361 36035 7395
rect 36737 7361 36771 7395
rect 2605 7293 2639 7327
rect 2881 7293 2915 7327
rect 4813 7293 4847 7327
rect 5457 7293 5491 7327
rect 6009 7293 6043 7327
rect 7113 7293 7147 7327
rect 7849 7293 7883 7327
rect 8493 7293 8527 7327
rect 8861 7293 8895 7327
rect 9045 7293 9079 7327
rect 9597 7293 9631 7327
rect 10609 7293 10643 7327
rect 11345 7293 11379 7327
rect 11713 7293 11747 7327
rect 12909 7293 12943 7327
rect 13737 7293 13771 7327
rect 14105 7293 14139 7327
rect 18429 7293 18463 7327
rect 18981 7293 19015 7327
rect 19625 7293 19659 7327
rect 20269 7293 20303 7327
rect 20545 7293 20579 7327
rect 21925 7293 21959 7327
rect 22385 7293 22419 7327
rect 22753 7293 22787 7327
rect 23857 7293 23891 7327
rect 23949 7293 23983 7327
rect 24409 7293 24443 7327
rect 24593 7293 24627 7327
rect 25697 7293 25731 7327
rect 26709 7293 26743 7327
rect 26985 7293 27019 7327
rect 27261 7293 27295 7327
rect 27905 7293 27939 7327
rect 28365 7293 28399 7327
rect 29745 7293 29779 7327
rect 29929 7293 29963 7327
rect 30113 7293 30147 7327
rect 33149 7293 33183 7327
rect 33701 7293 33735 7327
rect 34989 7293 35023 7327
rect 35817 7293 35851 7327
rect 36461 7293 36495 7327
rect 29285 7225 29319 7259
rect 6193 7157 6227 7191
rect 13001 7157 13035 7191
rect 24869 7157 24903 7191
rect 28549 7157 28583 7191
rect 11805 6953 11839 6987
rect 16497 6953 16531 6987
rect 36461 6953 36495 6987
rect 10885 6885 10919 6919
rect 32505 6885 32539 6919
rect 1869 6817 1903 6851
rect 4261 6817 4295 6851
rect 4721 6817 4755 6851
rect 5089 6817 5123 6851
rect 5457 6817 5491 6851
rect 5917 6817 5951 6851
rect 6745 6817 6779 6851
rect 8591 6817 8625 6851
rect 10149 6817 10183 6851
rect 10609 6817 10643 6851
rect 11897 6817 11931 6851
rect 12265 6817 12299 6851
rect 13645 6817 13679 6851
rect 14013 6817 14047 6851
rect 15485 6817 15519 6851
rect 15853 6817 15887 6851
rect 16681 6817 16715 6851
rect 16865 6817 16899 6851
rect 17325 6817 17359 6851
rect 17509 6817 17543 6851
rect 18153 6817 18187 6851
rect 18429 6817 18463 6851
rect 19441 6817 19475 6851
rect 19809 6817 19843 6851
rect 20177 6817 20211 6851
rect 20913 6817 20947 6851
rect 21741 6817 21775 6851
rect 22569 6817 22603 6851
rect 22845 6817 22879 6851
rect 23213 6817 23247 6851
rect 24225 6817 24259 6851
rect 24501 6817 24535 6851
rect 26617 6817 26651 6851
rect 27261 6817 27295 6851
rect 27537 6817 27571 6851
rect 27905 6817 27939 6851
rect 28825 6817 28859 6851
rect 29193 6817 29227 6851
rect 29469 6817 29503 6851
rect 31033 6817 31067 6851
rect 31401 6817 31435 6851
rect 31493 6817 31527 6851
rect 32137 6817 32171 6851
rect 32321 6817 32355 6851
rect 32413 6817 32447 6851
rect 32873 6817 32907 6851
rect 34253 6817 34287 6851
rect 35725 6817 35759 6851
rect 35909 6817 35943 6851
rect 36369 6817 36403 6851
rect 2145 6749 2179 6783
rect 4169 6749 4203 6783
rect 6469 6749 6503 6783
rect 12541 6749 12575 6783
rect 14473 6749 14507 6783
rect 19257 6749 19291 6783
rect 25605 6749 25639 6783
rect 27077 6749 27111 6783
rect 33425 6749 33459 6783
rect 33977 6749 34011 6783
rect 34437 6749 34471 6783
rect 34897 6749 34931 6783
rect 35449 6749 35483 6783
rect 8769 6681 8803 6715
rect 13553 6681 13587 6715
rect 15393 6681 15427 6715
rect 16865 6681 16899 6715
rect 21925 6681 21959 6715
rect 28917 6681 28951 6715
rect 30849 6681 30883 6715
rect 3433 6613 3467 6647
rect 7849 6613 7883 6647
rect 21097 6613 21131 6647
rect 22569 6613 22603 6647
rect 21465 6409 21499 6443
rect 24685 6409 24719 6443
rect 30849 6409 30883 6443
rect 38025 6409 38059 6443
rect 3525 6341 3559 6375
rect 20177 6341 20211 6375
rect 7849 6273 7883 6307
rect 13369 6273 13403 6307
rect 16129 6273 16163 6307
rect 17233 6273 17267 6307
rect 28733 6273 28767 6307
rect 29561 6273 29595 6307
rect 31861 6273 31895 6307
rect 32413 6273 32447 6307
rect 32873 6273 32907 6307
rect 34345 6273 34379 6307
rect 34989 6273 35023 6307
rect 36001 6273 36035 6307
rect 1869 6205 1903 6239
rect 2329 6205 2363 6239
rect 3617 6205 3651 6239
rect 3893 6205 3927 6239
rect 4445 6205 4479 6239
rect 4813 6205 4847 6239
rect 5365 6205 5399 6239
rect 5825 6205 5859 6239
rect 6837 6205 6871 6239
rect 7573 6205 7607 6239
rect 10149 6205 10183 6239
rect 10425 6205 10459 6239
rect 11161 6205 11195 6239
rect 11713 6205 11747 6239
rect 12449 6205 12483 6239
rect 13277 6205 13311 6239
rect 13645 6205 13679 6239
rect 15669 6205 15703 6239
rect 15761 6205 15795 6239
rect 15853 6205 15887 6239
rect 18061 6205 18095 6239
rect 18797 6205 18831 6239
rect 19073 6205 19107 6239
rect 21373 6205 21407 6239
rect 22017 6205 22051 6239
rect 22385 6205 22419 6239
rect 23673 6205 23707 6239
rect 24501 6205 24535 6239
rect 25237 6205 25271 6239
rect 25513 6205 25547 6239
rect 26893 6205 26927 6239
rect 28273 6205 28307 6239
rect 28549 6205 28583 6239
rect 29285 6205 29319 6239
rect 32689 6205 32723 6239
rect 33885 6205 33919 6239
rect 34161 6205 34195 6239
rect 35541 6205 35575 6239
rect 35817 6205 35851 6239
rect 37013 6205 37047 6239
rect 37289 6205 37323 6239
rect 37473 6205 37507 6239
rect 37933 6205 37967 6239
rect 10701 6137 10735 6171
rect 11897 6137 11931 6171
rect 27721 6137 27755 6171
rect 33333 6137 33367 6171
rect 36461 6137 36495 6171
rect 1869 6069 1903 6103
rect 6009 6069 6043 6103
rect 7021 6069 7055 6103
rect 9137 6069 9171 6103
rect 12541 6069 12575 6103
rect 13093 6069 13127 6103
rect 14749 6069 14783 6103
rect 15485 6069 15519 6103
rect 15761 6069 15795 6103
rect 18153 6069 18187 6103
rect 23857 6069 23891 6103
rect 2789 5865 2823 5899
rect 4261 5865 4295 5899
rect 9781 5865 9815 5899
rect 27077 5865 27111 5899
rect 11345 5797 11379 5831
rect 25329 5797 25363 5831
rect 26801 5797 26835 5831
rect 26985 5797 27019 5831
rect 27169 5797 27203 5831
rect 27537 5797 27571 5831
rect 27997 5797 28031 5831
rect 36093 5797 36127 5831
rect 4169 5729 4203 5763
rect 5089 5729 5123 5763
rect 5917 5729 5951 5763
rect 6377 5729 6411 5763
rect 6469 5729 6503 5763
rect 7113 5729 7147 5763
rect 7389 5729 7423 5763
rect 8309 5729 8343 5763
rect 8401 5729 8435 5763
rect 9689 5729 9723 5763
rect 10609 5729 10643 5763
rect 11069 5729 11103 5763
rect 11989 5729 12023 5763
rect 12357 5729 12391 5763
rect 12817 5729 12851 5763
rect 13185 5729 13219 5763
rect 13737 5729 13771 5763
rect 14473 5729 14507 5763
rect 15485 5729 15519 5763
rect 15853 5729 15887 5763
rect 16313 5729 16347 5763
rect 16681 5729 16715 5763
rect 17233 5729 17267 5763
rect 17693 5729 17727 5763
rect 19349 5729 19383 5763
rect 19901 5729 19935 5763
rect 20913 5729 20947 5763
rect 21005 5729 21039 5763
rect 21557 5729 21591 5763
rect 22477 5729 22511 5763
rect 22661 5729 22695 5763
rect 23121 5729 23155 5763
rect 24225 5729 24259 5763
rect 24777 5729 24811 5763
rect 24961 5729 24995 5763
rect 28825 5729 28859 5763
rect 29469 5729 29503 5763
rect 30297 5729 30331 5763
rect 31309 5729 31343 5763
rect 34713 5729 34747 5763
rect 36553 5729 36587 5763
rect 37749 5729 37783 5763
rect 1409 5661 1443 5695
rect 1685 5661 1719 5695
rect 6745 5661 6779 5695
rect 12725 5661 12759 5695
rect 19073 5661 19107 5695
rect 19809 5661 19843 5695
rect 22293 5661 22327 5695
rect 24041 5661 24075 5695
rect 28549 5661 28583 5695
rect 29009 5661 29043 5695
rect 30021 5661 30055 5695
rect 30481 5661 30515 5695
rect 32137 5661 32171 5695
rect 32413 5661 32447 5695
rect 33517 5661 33551 5695
rect 34437 5661 34471 5695
rect 8585 5593 8619 5627
rect 15393 5593 15427 5627
rect 36737 5593 36771 5627
rect 37933 5593 37967 5627
rect 5181 5525 5215 5559
rect 8125 5525 8159 5559
rect 14657 5525 14691 5559
rect 17877 5525 17911 5559
rect 21649 5525 21683 5559
rect 31493 5525 31527 5559
rect 2237 5321 2271 5355
rect 21373 5321 21407 5355
rect 23857 5321 23891 5355
rect 28457 5321 28491 5355
rect 33609 5321 33643 5355
rect 37749 5321 37783 5355
rect 6193 5253 6227 5287
rect 6929 5253 6963 5287
rect 9045 5253 9079 5287
rect 12817 5253 12851 5287
rect 13093 5253 13127 5287
rect 13921 5253 13955 5287
rect 22017 5253 22051 5287
rect 3433 5185 3467 5219
rect 7757 5185 7791 5219
rect 9689 5185 9723 5219
rect 1961 5117 1995 5151
rect 2053 5117 2087 5151
rect 3525 5117 3559 5151
rect 3801 5117 3835 5151
rect 4353 5117 4387 5151
rect 4721 5117 4755 5151
rect 5273 5117 5307 5151
rect 6009 5117 6043 5151
rect 6837 5117 6871 5151
rect 7481 5117 7515 5151
rect 9781 5117 9815 5151
rect 10241 5117 10275 5151
rect 10609 5117 10643 5151
rect 10977 5117 11011 5151
rect 11529 5117 11563 5151
rect 24961 5185 24995 5219
rect 27077 5185 27111 5219
rect 29837 5185 29871 5219
rect 32505 5185 32539 5219
rect 34897 5185 34931 5219
rect 35909 5185 35943 5219
rect 36645 5185 36679 5219
rect 12909 5117 12943 5151
rect 13645 5117 13679 5151
rect 14289 5117 14323 5151
rect 14657 5117 14691 5151
rect 15025 5117 15059 5151
rect 15577 5117 15611 5151
rect 16497 5117 16531 5151
rect 16957 5117 16991 5151
rect 18061 5117 18095 5151
rect 18613 5117 18647 5151
rect 19533 5117 19567 5151
rect 20085 5117 20119 5151
rect 20545 5117 20579 5151
rect 21189 5117 21223 5151
rect 22201 5117 22235 5151
rect 22569 5117 22603 5151
rect 22937 5117 22971 5151
rect 23673 5117 23707 5151
rect 25237 5117 25271 5151
rect 27353 5117 27387 5151
rect 30389 5117 30423 5151
rect 30665 5117 30699 5151
rect 30849 5117 30883 5151
rect 32781 5117 32815 5151
rect 32965 5117 32999 5151
rect 33425 5117 33459 5151
rect 35449 5117 35483 5151
rect 35725 5117 35759 5151
rect 36369 5117 36403 5151
rect 17233 5049 17267 5083
rect 18797 5049 18831 5083
rect 20729 5049 20763 5083
rect 26617 5049 26651 5083
rect 31953 5049 31987 5083
rect 12817 4981 12851 5015
rect 2789 4777 2823 4811
rect 14657 4777 14691 4811
rect 21005 4777 21039 4811
rect 23397 4777 23431 4811
rect 31125 4777 31159 4811
rect 9137 4709 9171 4743
rect 25237 4709 25271 4743
rect 25881 4709 25915 4743
rect 32137 4709 32171 4743
rect 33609 4709 33643 4743
rect 4445 4641 4479 4675
rect 5273 4641 5307 4675
rect 5549 4641 5583 4675
rect 6101 4641 6135 4675
rect 6469 4641 6503 4675
rect 6837 4641 6871 4675
rect 7481 4641 7515 4675
rect 10241 4641 10275 4675
rect 10701 4641 10735 4675
rect 10885 4641 10919 4675
rect 11253 4641 11287 4675
rect 11713 4641 11747 4675
rect 12725 4641 12759 4675
rect 14565 4641 14599 4675
rect 15761 4641 15795 4675
rect 16865 4641 16899 4675
rect 17509 4641 17543 4675
rect 17877 4641 17911 4675
rect 18245 4641 18279 4675
rect 18521 4641 18555 4675
rect 19809 4641 19843 4675
rect 20177 4641 20211 4675
rect 20913 4641 20947 4675
rect 21925 4641 21959 4675
rect 22293 4641 22327 4675
rect 22569 4641 22603 4675
rect 23305 4641 23339 4675
rect 24133 4641 24167 4675
rect 24225 4641 24259 4675
rect 24685 4641 24719 4675
rect 24869 4641 24903 4675
rect 25789 4641 25823 4675
rect 26801 4641 26835 4675
rect 27077 4641 27111 4675
rect 30021 4641 30055 4675
rect 30297 4641 30331 4675
rect 30481 4641 30515 4675
rect 30941 4641 30975 4675
rect 32689 4641 32723 4675
rect 32827 4641 32861 4675
rect 32965 4641 32999 4675
rect 34437 4641 34471 4675
rect 34621 4641 34655 4675
rect 35633 4641 35667 4675
rect 35909 4641 35943 4675
rect 36553 4641 36587 4675
rect 37749 4641 37783 4675
rect 1409 4573 1443 4607
rect 1685 4573 1719 4607
rect 5457 4573 5491 4607
rect 7757 4573 7791 4607
rect 12449 4573 12483 4607
rect 15669 4573 15703 4607
rect 19441 4573 19475 4607
rect 21741 4573 21775 4607
rect 28181 4573 28215 4607
rect 29469 4573 29503 4607
rect 34161 4573 34195 4607
rect 35081 4573 35115 4607
rect 36093 4573 36127 4607
rect 10149 4505 10183 4539
rect 16957 4505 16991 4539
rect 20085 4505 20119 4539
rect 4537 4437 4571 4471
rect 13829 4437 13863 4471
rect 15945 4437 15979 4471
rect 36737 4437 36771 4471
rect 37933 4437 37967 4471
rect 8217 4233 8251 4267
rect 19441 4233 19475 4267
rect 21557 4233 21591 4267
rect 27169 4233 27203 4267
rect 9505 4165 9539 4199
rect 30665 4165 30699 4199
rect 3249 4097 3283 4131
rect 7113 4097 7147 4131
rect 12541 4097 12575 4131
rect 15025 4097 15059 4131
rect 16129 4097 16163 4131
rect 18337 4097 18371 4131
rect 23673 4097 23707 4131
rect 24869 4097 24903 4131
rect 28733 4097 28767 4131
rect 29285 4097 29319 4131
rect 32229 4097 32263 4131
rect 32689 4097 32723 4131
rect 33701 4097 33735 4131
rect 34161 4097 34195 4131
rect 37473 4097 37507 4131
rect 1961 4029 1995 4063
rect 2237 4029 2271 4063
rect 2973 4029 3007 4063
rect 5089 4029 5123 4063
rect 5549 4029 5583 4063
rect 6837 4029 6871 4063
rect 9597 4029 9631 4063
rect 9873 4029 9907 4063
rect 10425 4029 10459 4063
rect 10609 4029 10643 4063
rect 11345 4029 11379 4063
rect 12449 4029 12483 4063
rect 13093 4029 13127 4063
rect 13737 4029 13771 4063
rect 13870 4029 13904 4063
rect 14749 4029 14783 4063
rect 16957 4029 16991 4063
rect 17049 4029 17083 4063
rect 18061 4029 18095 4063
rect 20177 4029 20211 4063
rect 20453 4029 20487 4063
rect 22293 4029 22327 4063
rect 22385 4029 22419 4063
rect 23765 4029 23799 4063
rect 25145 4029 25179 4063
rect 26985 4029 27019 4063
rect 28273 4029 28307 4063
rect 28549 4029 28583 4063
rect 29561 4029 29595 4063
rect 32505 4029 32539 4063
rect 33977 4029 34011 4063
rect 34989 4029 35023 4063
rect 36093 4029 36127 4063
rect 36369 4029 36403 4063
rect 14289 3961 14323 3995
rect 17509 3961 17543 3995
rect 22845 3961 22879 3995
rect 24225 3961 24259 3995
rect 26525 3961 26559 3995
rect 27721 3961 27755 3995
rect 31677 3961 31711 3995
rect 33149 3961 33183 3995
rect 1777 3893 1811 3927
rect 4537 3893 4571 3927
rect 5181 3893 5215 3927
rect 13185 3893 13219 3927
rect 35173 3893 35207 3927
rect 6561 3689 6595 3723
rect 11989 3689 12023 3723
rect 15393 3689 15427 3723
rect 25789 3689 25823 3723
rect 26617 3689 26651 3723
rect 36277 3689 36311 3723
rect 37933 3689 37967 3723
rect 20361 3621 20395 3655
rect 29469 3621 29503 3655
rect 29929 3621 29963 3655
rect 34437 3621 34471 3655
rect 2145 3553 2179 3587
rect 3525 3553 3559 3587
rect 4261 3553 4295 3587
rect 5457 3553 5491 3587
rect 7481 3553 7515 3587
rect 8677 3553 8711 3587
rect 8953 3553 8987 3587
rect 9137 3553 9171 3587
rect 9965 3553 9999 3587
rect 11805 3553 11839 3587
rect 12817 3553 12851 3587
rect 15301 3553 15335 3587
rect 15853 3553 15887 3587
rect 16865 3553 16899 3587
rect 19625 3553 19659 3587
rect 20177 3553 20211 3587
rect 21189 3553 21223 3587
rect 21281 3553 21315 3587
rect 21649 3553 21683 3587
rect 22753 3553 22787 3587
rect 22937 3553 22971 3587
rect 23397 3553 23431 3587
rect 23489 3553 23523 3587
rect 24777 3553 24811 3587
rect 25329 3553 25363 3587
rect 25513 3553 25547 3587
rect 26525 3553 26559 3587
rect 27169 3553 27203 3587
rect 28089 3553 28123 3587
rect 30481 3553 30515 3587
rect 30757 3553 30791 3587
rect 35173 3553 35207 3587
rect 37749 3553 37783 3587
rect 1869 3485 1903 3519
rect 4169 3485 4203 3519
rect 4721 3485 4755 3519
rect 5181 3485 5215 3519
rect 7389 3485 7423 3519
rect 7941 3485 7975 3519
rect 9689 3485 9723 3519
rect 11345 3485 11379 3519
rect 12541 3485 12575 3519
rect 16589 3485 16623 3519
rect 19349 3485 19383 3519
rect 21005 3485 21039 3519
rect 24593 3485 24627 3519
rect 27813 3485 27847 3519
rect 30941 3485 30975 3519
rect 32781 3485 32815 3519
rect 33057 3485 33091 3519
rect 34897 3485 34931 3519
rect 17969 3417 18003 3451
rect 14105 3349 14139 3383
rect 23949 3349 23983 3383
rect 27261 3349 27295 3383
rect 2053 3145 2087 3179
rect 4905 3145 4939 3179
rect 8217 3145 8251 3179
rect 9229 3145 9263 3179
rect 11437 3145 11471 3179
rect 14013 3145 14047 3179
rect 15945 3145 15979 3179
rect 19441 3145 19475 3179
rect 9781 3077 9815 3111
rect 22201 3077 22235 3111
rect 23029 3077 23063 3111
rect 27537 3077 27571 3111
rect 32597 3077 32631 3111
rect 2881 3009 2915 3043
rect 6285 3009 6319 3043
rect 12449 3009 12483 3043
rect 14841 3009 14875 3043
rect 23673 3009 23707 3043
rect 23949 3009 23983 3043
rect 25053 3009 25087 3043
rect 25973 3009 26007 3043
rect 29285 3009 29319 3043
rect 29837 3009 29871 3043
rect 30297 3009 30331 3043
rect 34345 3009 34379 3043
rect 34897 3009 34931 3043
rect 35449 3009 35483 3043
rect 36737 3009 36771 3043
rect 1961 2941 1995 2975
rect 2605 2941 2639 2975
rect 4721 2941 4755 2975
rect 5825 2941 5859 2975
rect 6101 2941 6135 2975
rect 6837 2941 6871 2975
rect 7113 2941 7147 2975
rect 9045 2941 9079 2975
rect 9781 2941 9815 2975
rect 9873 2941 9907 2975
rect 10149 2941 10183 2975
rect 12725 2941 12759 2975
rect 14565 2941 14599 2975
rect 16773 2941 16807 2975
rect 17325 2941 17359 2975
rect 18061 2941 18095 2975
rect 18337 2941 18371 2975
rect 20637 2941 20671 2975
rect 20913 2941 20947 2975
rect 22937 2941 22971 2975
rect 26249 2941 26283 2975
rect 28089 2941 28123 2975
rect 30113 2941 30147 2975
rect 31217 2941 31251 2975
rect 31493 2941 31527 2975
rect 33885 2941 33919 2975
rect 34161 2941 34195 2975
rect 35587 2941 35621 2975
rect 35725 2941 35759 2975
rect 36461 2941 36495 2975
rect 4261 2873 4295 2907
rect 17509 2873 17543 2907
rect 28181 2873 28215 2907
rect 33333 2873 33367 2907
rect 38117 2873 38151 2907
rect 9873 2601 9907 2635
rect 22569 2601 22603 2635
rect 6285 2533 6319 2567
rect 12081 2533 12115 2567
rect 14933 2533 14967 2567
rect 32045 2533 32079 2567
rect 35449 2533 35483 2567
rect 1685 2465 1719 2499
rect 4629 2465 4663 2499
rect 4905 2465 4939 2499
rect 6929 2465 6963 2499
rect 7573 2465 7607 2499
rect 8125 2465 8159 2499
rect 8401 2465 8435 2499
rect 9781 2465 9815 2499
rect 10701 2465 10735 2499
rect 12725 2465 12759 2499
rect 13737 2465 13771 2499
rect 14473 2465 14507 2499
rect 15669 2465 15703 2499
rect 15945 2465 15979 2499
rect 18337 2465 18371 2499
rect 21465 2465 21499 2499
rect 24869 2465 24903 2499
rect 27169 2465 27203 2499
rect 30389 2465 30423 2499
rect 30665 2465 30699 2499
rect 33517 2465 33551 2499
rect 36001 2465 36035 2499
rect 36277 2465 36311 2499
rect 36461 2465 36495 2499
rect 1409 2397 1443 2431
rect 7021 2397 7055 2431
rect 10425 2397 10459 2431
rect 12633 2397 12667 2431
rect 14381 2397 14415 2431
rect 18981 2397 19015 2431
rect 19257 2397 19291 2431
rect 21189 2397 21223 2431
rect 24593 2397 24627 2431
rect 26893 2397 26927 2431
rect 29745 2397 29779 2431
rect 33241 2397 33275 2431
rect 7757 2329 7791 2363
rect 13829 2329 13863 2363
rect 2789 2261 2823 2295
rect 12909 2261 12943 2295
rect 17049 2261 17083 2295
rect 18429 2261 18463 2295
rect 20545 2261 20579 2295
rect 26157 2261 26191 2295
rect 28457 2261 28491 2295
rect 33149 2261 33183 2295
rect 34805 2261 34839 2295
rect 37565 2261 37599 2295
<< metal1 >>
rect 21910 39108 21916 39160
rect 21968 39148 21974 39160
rect 23750 39148 23756 39160
rect 21968 39120 23756 39148
rect 21968 39108 21974 39120
rect 23750 39108 23756 39120
rect 23808 39108 23814 39160
rect 1104 37562 38824 37584
rect 1104 37510 19606 37562
rect 19658 37510 19670 37562
rect 19722 37510 19734 37562
rect 19786 37510 19798 37562
rect 19850 37510 38824 37562
rect 1104 37488 38824 37510
rect 24581 37451 24639 37457
rect 24581 37417 24593 37451
rect 24627 37448 24639 37451
rect 24627 37420 25820 37448
rect 24627 37417 24639 37420
rect 24581 37411 24639 37417
rect 4985 37383 5043 37389
rect 4985 37349 4997 37383
rect 5031 37380 5043 37383
rect 5442 37380 5448 37392
rect 5031 37352 5448 37380
rect 5031 37349 5043 37352
rect 4985 37343 5043 37349
rect 5442 37340 5448 37352
rect 5500 37340 5506 37392
rect 9217 37383 9275 37389
rect 9217 37349 9229 37383
rect 9263 37380 9275 37383
rect 9398 37380 9404 37392
rect 9263 37352 9404 37380
rect 9263 37349 9275 37352
rect 9217 37343 9275 37349
rect 9398 37340 9404 37352
rect 9456 37340 9462 37392
rect 4249 37315 4307 37321
rect 4249 37281 4261 37315
rect 4295 37312 4307 37315
rect 4706 37312 4712 37324
rect 4295 37284 4712 37312
rect 4295 37281 4307 37284
rect 4249 37275 4307 37281
rect 4706 37272 4712 37284
rect 4764 37272 4770 37324
rect 4893 37315 4951 37321
rect 4893 37281 4905 37315
rect 4939 37312 4951 37315
rect 5537 37315 5595 37321
rect 4939 37284 5488 37312
rect 4939 37281 4951 37284
rect 4893 37275 4951 37281
rect 5460 37244 5488 37284
rect 5537 37281 5549 37315
rect 5583 37312 5595 37315
rect 6914 37312 6920 37324
rect 5583 37284 6920 37312
rect 5583 37281 5595 37284
rect 5537 37275 5595 37281
rect 6914 37272 6920 37284
rect 6972 37272 6978 37324
rect 7558 37312 7564 37324
rect 7519 37284 7564 37312
rect 7558 37272 7564 37284
rect 7616 37272 7622 37324
rect 7834 37312 7840 37324
rect 7795 37284 7840 37312
rect 7834 37272 7840 37284
rect 7892 37272 7898 37324
rect 7926 37272 7932 37324
rect 7984 37312 7990 37324
rect 9674 37312 9680 37324
rect 7984 37284 9680 37312
rect 7984 37272 7990 37284
rect 9674 37272 9680 37284
rect 9732 37272 9738 37324
rect 9769 37315 9827 37321
rect 9769 37281 9781 37315
rect 9815 37312 9827 37315
rect 9858 37312 9864 37324
rect 9815 37284 9864 37312
rect 9815 37281 9827 37284
rect 9769 37275 9827 37281
rect 9858 37272 9864 37284
rect 9916 37272 9922 37324
rect 11698 37312 11704 37324
rect 11659 37284 11704 37312
rect 11698 37272 11704 37284
rect 11756 37272 11762 37324
rect 21266 37272 21272 37324
rect 21324 37312 21330 37324
rect 24673 37315 24731 37321
rect 24673 37312 24685 37315
rect 21324 37284 24685 37312
rect 21324 37272 21330 37284
rect 24673 37281 24685 37284
rect 24719 37281 24731 37315
rect 24946 37312 24952 37324
rect 24907 37284 24952 37312
rect 24673 37275 24731 37281
rect 24946 37272 24952 37284
rect 25004 37272 25010 37324
rect 5626 37244 5632 37256
rect 5460 37216 5632 37244
rect 5626 37204 5632 37216
rect 5684 37204 5690 37256
rect 15470 37244 15476 37256
rect 15431 37216 15476 37244
rect 15470 37204 15476 37216
rect 15528 37204 15534 37256
rect 15746 37244 15752 37256
rect 15707 37216 15752 37244
rect 15746 37204 15752 37216
rect 15804 37204 15810 37256
rect 1302 37136 1308 37188
rect 1360 37176 1366 37188
rect 7466 37176 7472 37188
rect 1360 37148 7472 37176
rect 1360 37136 1366 37148
rect 7466 37136 7472 37148
rect 7524 37136 7530 37188
rect 9674 37136 9680 37188
rect 9732 37176 9738 37188
rect 24581 37179 24639 37185
rect 24581 37176 24593 37179
rect 9732 37148 12388 37176
rect 9732 37136 9738 37148
rect 4341 37111 4399 37117
rect 4341 37077 4353 37111
rect 4387 37108 4399 37111
rect 4798 37108 4804 37120
rect 4387 37080 4804 37108
rect 4387 37077 4399 37080
rect 4341 37071 4399 37077
rect 4798 37068 4804 37080
rect 4856 37068 4862 37120
rect 5718 37108 5724 37120
rect 5679 37080 5724 37108
rect 5718 37068 5724 37080
rect 5776 37068 5782 37120
rect 9858 37108 9864 37120
rect 9819 37080 9864 37108
rect 9858 37068 9864 37080
rect 9916 37068 9922 37120
rect 11793 37111 11851 37117
rect 11793 37077 11805 37111
rect 11839 37108 11851 37111
rect 12250 37108 12256 37120
rect 11839 37080 12256 37108
rect 11839 37077 11851 37080
rect 11793 37071 11851 37077
rect 12250 37068 12256 37080
rect 12308 37068 12314 37120
rect 12360 37108 12388 37148
rect 16408 37148 24593 37176
rect 16408 37108 16436 37148
rect 24581 37145 24593 37148
rect 24627 37145 24639 37179
rect 25792 37176 25820 37420
rect 31665 37383 31723 37389
rect 31665 37349 31677 37383
rect 31711 37380 31723 37383
rect 32030 37380 32036 37392
rect 31711 37352 32036 37380
rect 31711 37349 31723 37352
rect 31665 37343 31723 37349
rect 32030 37340 32036 37352
rect 32088 37340 32094 37392
rect 34425 37383 34483 37389
rect 34425 37349 34437 37383
rect 34471 37380 34483 37383
rect 36446 37380 36452 37392
rect 34471 37352 36452 37380
rect 34471 37349 34483 37352
rect 34425 37343 34483 37349
rect 36446 37340 36452 37352
rect 36504 37380 36510 37392
rect 36504 37352 36952 37380
rect 36504 37340 36510 37352
rect 29178 37272 29184 37324
rect 29236 37312 29242 37324
rect 29825 37315 29883 37321
rect 29825 37312 29837 37315
rect 29236 37284 29837 37312
rect 29236 37272 29242 37284
rect 29825 37281 29837 37284
rect 29871 37312 29883 37315
rect 30285 37315 30343 37321
rect 30285 37312 30297 37315
rect 29871 37284 30297 37312
rect 29871 37281 29883 37284
rect 29825 37275 29883 37281
rect 30285 37281 30297 37284
rect 30331 37281 30343 37315
rect 30285 37275 30343 37281
rect 33134 37272 33140 37324
rect 33192 37312 33198 37324
rect 33689 37315 33747 37321
rect 33689 37312 33701 37315
rect 33192 37284 33701 37312
rect 33192 37272 33198 37284
rect 33689 37281 33701 37284
rect 33735 37281 33747 37315
rect 33689 37275 33747 37281
rect 34149 37315 34207 37321
rect 34149 37281 34161 37315
rect 34195 37281 34207 37315
rect 35894 37312 35900 37324
rect 35855 37284 35900 37312
rect 34149 37275 34207 37281
rect 28994 37204 29000 37256
rect 29052 37244 29058 37256
rect 30006 37244 30012 37256
rect 29052 37216 30012 37244
rect 29052 37204 29058 37216
rect 30006 37204 30012 37216
rect 30064 37204 30070 37256
rect 33502 37204 33508 37256
rect 33560 37244 33566 37256
rect 34164 37244 34192 37275
rect 35894 37272 35900 37284
rect 35952 37272 35958 37324
rect 36924 37321 36952 37352
rect 36265 37315 36323 37321
rect 36265 37312 36277 37315
rect 36004 37284 36277 37312
rect 33560 37216 34192 37244
rect 33560 37204 33566 37216
rect 35526 37204 35532 37256
rect 35584 37244 35590 37256
rect 36004 37244 36032 37284
rect 36265 37281 36277 37284
rect 36311 37281 36323 37315
rect 36265 37275 36323 37281
rect 36909 37315 36967 37321
rect 36909 37281 36921 37315
rect 36955 37281 36967 37315
rect 36909 37275 36967 37281
rect 36998 37272 37004 37324
rect 37056 37312 37062 37324
rect 37093 37315 37151 37321
rect 37093 37312 37105 37315
rect 37056 37284 37105 37312
rect 37056 37272 37062 37284
rect 37093 37281 37105 37284
rect 37139 37281 37151 37315
rect 37093 37275 37151 37281
rect 37182 37272 37188 37324
rect 37240 37312 37246 37324
rect 37240 37284 37285 37312
rect 37240 37272 37246 37284
rect 35584 37216 36032 37244
rect 36357 37247 36415 37253
rect 35584 37204 35590 37216
rect 36357 37213 36369 37247
rect 36403 37244 36415 37247
rect 36403 37216 37136 37244
rect 36403 37213 36415 37216
rect 36357 37207 36415 37213
rect 37108 37188 37136 37216
rect 35713 37179 35771 37185
rect 25792 37148 30052 37176
rect 24581 37139 24639 37145
rect 16850 37108 16856 37120
rect 12360 37080 16436 37108
rect 16811 37080 16856 37108
rect 16850 37068 16856 37080
rect 16908 37068 16914 37120
rect 26234 37108 26240 37120
rect 26195 37080 26240 37108
rect 26234 37068 26240 37080
rect 26292 37068 26298 37120
rect 30024 37108 30052 37148
rect 35713 37145 35725 37179
rect 35759 37176 35771 37179
rect 36722 37176 36728 37188
rect 35759 37148 36728 37176
rect 35759 37145 35771 37148
rect 35713 37139 35771 37145
rect 36722 37136 36728 37148
rect 36780 37136 36786 37188
rect 37090 37136 37096 37188
rect 37148 37136 37154 37188
rect 31018 37108 31024 37120
rect 30024 37080 31024 37108
rect 31018 37068 31024 37080
rect 31076 37068 31082 37120
rect 36998 37068 37004 37120
rect 37056 37108 37062 37120
rect 37369 37111 37427 37117
rect 37369 37108 37381 37111
rect 37056 37080 37381 37108
rect 37056 37068 37062 37080
rect 37369 37077 37381 37080
rect 37415 37077 37427 37111
rect 37369 37071 37427 37077
rect 1104 37018 38824 37040
rect 1104 36966 4246 37018
rect 4298 36966 4310 37018
rect 4362 36966 4374 37018
rect 4426 36966 4438 37018
rect 4490 36966 34966 37018
rect 35018 36966 35030 37018
rect 35082 36966 35094 37018
rect 35146 36966 35158 37018
rect 35210 36966 38824 37018
rect 1104 36944 38824 36966
rect 2685 36907 2743 36913
rect 2685 36873 2697 36907
rect 2731 36904 2743 36907
rect 2774 36904 2780 36916
rect 2731 36876 2780 36904
rect 2731 36873 2743 36876
rect 2685 36867 2743 36873
rect 2774 36864 2780 36876
rect 2832 36864 2838 36916
rect 3988 36876 7144 36904
rect 2409 36839 2467 36845
rect 2409 36805 2421 36839
rect 2455 36836 2467 36839
rect 2498 36836 2504 36848
rect 2455 36808 2504 36836
rect 2455 36805 2467 36808
rect 2409 36799 2467 36805
rect 2498 36796 2504 36808
rect 2556 36836 2562 36848
rect 3988 36836 4016 36876
rect 2556 36808 4016 36836
rect 2556 36796 2562 36808
rect 6822 36796 6828 36848
rect 6880 36836 6886 36848
rect 7009 36839 7067 36845
rect 7009 36836 7021 36839
rect 6880 36808 7021 36836
rect 6880 36796 6886 36808
rect 7009 36805 7021 36808
rect 7055 36805 7067 36839
rect 7116 36836 7144 36876
rect 7466 36864 7472 36916
rect 7524 36904 7530 36916
rect 35253 36907 35311 36913
rect 7524 36876 29776 36904
rect 7524 36864 7530 36876
rect 7926 36836 7932 36848
rect 7116 36808 7932 36836
rect 7009 36799 7067 36805
rect 7926 36796 7932 36808
rect 7984 36796 7990 36848
rect 13814 36836 13820 36848
rect 13775 36808 13820 36836
rect 13814 36796 13820 36808
rect 13872 36796 13878 36848
rect 15013 36839 15071 36845
rect 15013 36805 15025 36839
rect 15059 36836 15071 36839
rect 15746 36836 15752 36848
rect 15059 36808 15752 36836
rect 15059 36805 15071 36808
rect 15013 36799 15071 36805
rect 15746 36796 15752 36808
rect 15804 36796 15810 36848
rect 16025 36771 16083 36777
rect 1780 36740 2728 36768
rect 1780 36709 1808 36740
rect 1765 36703 1823 36709
rect 1765 36669 1777 36703
rect 1811 36669 1823 36703
rect 2498 36700 2504 36712
rect 2459 36672 2504 36700
rect 1765 36663 1823 36669
rect 2498 36660 2504 36672
rect 2556 36660 2562 36712
rect 2700 36700 2728 36740
rect 3160 36740 14964 36768
rect 3160 36700 3188 36740
rect 3326 36700 3332 36712
rect 2700 36672 3188 36700
rect 3287 36672 3332 36700
rect 3326 36660 3332 36672
rect 3384 36660 3390 36712
rect 3970 36700 3976 36712
rect 3931 36672 3976 36700
rect 3970 36660 3976 36672
rect 4028 36660 4034 36712
rect 4249 36703 4307 36709
rect 4249 36700 4261 36703
rect 4080 36672 4261 36700
rect 3421 36635 3479 36641
rect 3421 36601 3433 36635
rect 3467 36632 3479 36635
rect 4080 36632 4108 36672
rect 4249 36669 4261 36672
rect 4295 36669 4307 36703
rect 4249 36663 4307 36669
rect 5810 36660 5816 36712
rect 5868 36700 5874 36712
rect 6089 36703 6147 36709
rect 6089 36700 6101 36703
rect 5868 36672 6101 36700
rect 5868 36660 5874 36672
rect 6089 36669 6101 36672
rect 6135 36669 6147 36703
rect 6089 36663 6147 36669
rect 6825 36703 6883 36709
rect 6825 36669 6837 36703
rect 6871 36669 6883 36703
rect 6825 36663 6883 36669
rect 5626 36632 5632 36644
rect 3467 36604 4108 36632
rect 5539 36604 5632 36632
rect 3467 36601 3479 36604
rect 3421 36595 3479 36601
rect 5626 36592 5632 36604
rect 5684 36632 5690 36644
rect 6840 36632 6868 36663
rect 7466 36660 7472 36712
rect 7524 36700 7530 36712
rect 8202 36700 8208 36712
rect 7524 36672 8208 36700
rect 7524 36660 7530 36672
rect 8202 36660 8208 36672
rect 8260 36700 8266 36712
rect 8665 36703 8723 36709
rect 8665 36700 8677 36703
rect 8260 36672 8677 36700
rect 8260 36660 8266 36672
rect 8665 36669 8677 36672
rect 8711 36669 8723 36703
rect 8665 36663 8723 36669
rect 8941 36703 8999 36709
rect 8941 36669 8953 36703
rect 8987 36700 8999 36703
rect 9858 36700 9864 36712
rect 8987 36672 9864 36700
rect 8987 36669 8999 36672
rect 8941 36663 8999 36669
rect 9858 36660 9864 36672
rect 9916 36660 9922 36712
rect 11054 36700 11060 36712
rect 11015 36672 11060 36700
rect 11054 36660 11060 36672
rect 11112 36660 11118 36712
rect 11514 36660 11520 36712
rect 11572 36700 11578 36712
rect 11701 36703 11759 36709
rect 11701 36700 11713 36703
rect 11572 36672 11713 36700
rect 11572 36660 11578 36672
rect 11701 36669 11713 36672
rect 11747 36669 11759 36703
rect 12434 36700 12440 36712
rect 12395 36672 12440 36700
rect 11701 36663 11759 36669
rect 12434 36660 12440 36672
rect 12492 36660 12498 36712
rect 12713 36703 12771 36709
rect 12713 36669 12725 36703
rect 12759 36700 12771 36703
rect 12802 36700 12808 36712
rect 12759 36672 12808 36700
rect 12759 36669 12771 36672
rect 12713 36663 12771 36669
rect 12802 36660 12808 36672
rect 12860 36660 12866 36712
rect 14936 36709 14964 36740
rect 16025 36737 16037 36771
rect 16071 36768 16083 36771
rect 16850 36768 16856 36780
rect 16071 36740 16856 36768
rect 16071 36737 16083 36740
rect 16025 36731 16083 36737
rect 16850 36728 16856 36740
rect 16908 36728 16914 36780
rect 23842 36768 23848 36780
rect 16960 36740 23848 36768
rect 14921 36703 14979 36709
rect 14921 36669 14933 36703
rect 14967 36669 14979 36703
rect 14921 36663 14979 36669
rect 5684 36604 6868 36632
rect 14936 36632 14964 36663
rect 15470 36660 15476 36712
rect 15528 36700 15534 36712
rect 15746 36700 15752 36712
rect 15528 36672 15752 36700
rect 15528 36660 15534 36672
rect 15746 36660 15752 36672
rect 15804 36660 15810 36712
rect 16960 36700 16988 36740
rect 23842 36728 23848 36740
rect 23900 36728 23906 36780
rect 15856 36672 16988 36700
rect 18049 36703 18107 36709
rect 15856 36632 15884 36672
rect 18049 36669 18061 36703
rect 18095 36669 18107 36703
rect 18322 36700 18328 36712
rect 18283 36672 18328 36700
rect 18049 36663 18107 36669
rect 14936 36604 15884 36632
rect 5684 36592 5690 36604
rect 18064 36576 18092 36663
rect 18322 36660 18328 36672
rect 18380 36660 18386 36712
rect 20533 36703 20591 36709
rect 20533 36669 20545 36703
rect 20579 36700 20591 36703
rect 20806 36700 20812 36712
rect 20579 36672 20812 36700
rect 20579 36669 20591 36672
rect 20533 36663 20591 36669
rect 20806 36660 20812 36672
rect 20864 36660 20870 36712
rect 21266 36700 21272 36712
rect 21227 36672 21272 36700
rect 21266 36660 21272 36672
rect 21324 36660 21330 36712
rect 21542 36700 21548 36712
rect 21503 36672 21548 36700
rect 21542 36660 21548 36672
rect 21600 36660 21606 36712
rect 23014 36660 23020 36712
rect 23072 36700 23078 36712
rect 23661 36703 23719 36709
rect 23661 36700 23673 36703
rect 23072 36672 23673 36700
rect 23072 36660 23078 36672
rect 23661 36669 23673 36672
rect 23707 36669 23719 36703
rect 23934 36700 23940 36712
rect 23895 36672 23940 36700
rect 23661 36663 23719 36669
rect 23934 36660 23940 36672
rect 23992 36660 23998 36712
rect 26510 36660 26516 36712
rect 26568 36700 26574 36712
rect 26881 36703 26939 36709
rect 26881 36700 26893 36703
rect 26568 36672 26893 36700
rect 26568 36660 26574 36672
rect 26881 36669 26893 36672
rect 26927 36669 26939 36703
rect 27154 36700 27160 36712
rect 27115 36672 27160 36700
rect 26881 36663 26939 36669
rect 27154 36660 27160 36672
rect 27212 36660 27218 36712
rect 29748 36709 29776 36876
rect 32692 36876 33640 36904
rect 30006 36728 30012 36780
rect 30064 36768 30070 36780
rect 30282 36768 30288 36780
rect 30064 36740 30288 36768
rect 30064 36728 30070 36740
rect 30282 36728 30288 36740
rect 30340 36768 30346 36780
rect 32692 36777 32720 36876
rect 33612 36836 33640 36876
rect 35253 36873 35265 36907
rect 35299 36904 35311 36907
rect 37182 36904 37188 36916
rect 35299 36876 37188 36904
rect 35299 36873 35311 36876
rect 35253 36867 35311 36873
rect 37182 36864 37188 36876
rect 37240 36864 37246 36916
rect 35986 36836 35992 36848
rect 33612 36808 35992 36836
rect 35986 36796 35992 36808
rect 36044 36796 36050 36848
rect 37090 36796 37096 36848
rect 37148 36836 37154 36848
rect 37369 36839 37427 36845
rect 37369 36836 37381 36839
rect 37148 36808 37381 36836
rect 37148 36796 37154 36808
rect 37369 36805 37381 36808
rect 37415 36805 37427 36839
rect 37369 36799 37427 36805
rect 30561 36771 30619 36777
rect 30561 36768 30573 36771
rect 30340 36740 30573 36768
rect 30340 36728 30346 36740
rect 30561 36737 30573 36740
rect 30607 36768 30619 36771
rect 32677 36771 32735 36777
rect 32677 36768 32689 36771
rect 30607 36740 32689 36768
rect 30607 36737 30619 36740
rect 30561 36731 30619 36737
rect 32677 36737 32689 36740
rect 32723 36737 32735 36771
rect 36170 36768 36176 36780
rect 32677 36731 32735 36737
rect 32784 36740 36176 36768
rect 29549 36703 29607 36709
rect 29549 36669 29561 36703
rect 29595 36669 29607 36703
rect 29549 36663 29607 36669
rect 29733 36703 29791 36709
rect 29733 36669 29745 36703
rect 29779 36669 29791 36703
rect 30834 36700 30840 36712
rect 30795 36672 30840 36700
rect 29733 36663 29791 36669
rect 21284 36632 21312 36660
rect 18984 36604 21312 36632
rect 22925 36635 22983 36641
rect 1946 36564 1952 36576
rect 1907 36536 1952 36564
rect 1946 36524 1952 36536
rect 2004 36524 2010 36576
rect 6181 36567 6239 36573
rect 6181 36533 6193 36567
rect 6227 36564 6239 36567
rect 6914 36564 6920 36576
rect 6227 36536 6920 36564
rect 6227 36533 6239 36536
rect 6181 36527 6239 36533
rect 6914 36524 6920 36536
rect 6972 36524 6978 36576
rect 10042 36564 10048 36576
rect 10003 36536 10048 36564
rect 10042 36524 10048 36536
rect 10100 36524 10106 36576
rect 11149 36567 11207 36573
rect 11149 36533 11161 36567
rect 11195 36564 11207 36567
rect 11422 36564 11428 36576
rect 11195 36536 11428 36564
rect 11195 36533 11207 36536
rect 11149 36527 11207 36533
rect 11422 36524 11428 36536
rect 11480 36524 11486 36576
rect 11790 36564 11796 36576
rect 11751 36536 11796 36564
rect 11790 36524 11796 36536
rect 11848 36524 11854 36576
rect 17034 36524 17040 36576
rect 17092 36564 17098 36576
rect 17129 36567 17187 36573
rect 17129 36564 17141 36567
rect 17092 36536 17141 36564
rect 17092 36524 17098 36536
rect 17129 36533 17141 36536
rect 17175 36533 17187 36567
rect 18046 36564 18052 36576
rect 17959 36536 18052 36564
rect 17129 36527 17187 36533
rect 18046 36524 18052 36536
rect 18104 36564 18110 36576
rect 18984 36564 19012 36604
rect 22925 36601 22937 36635
rect 22971 36632 22983 36635
rect 23290 36632 23296 36644
rect 22971 36604 23296 36632
rect 22971 36601 22983 36604
rect 22925 36595 22983 36601
rect 23290 36592 23296 36604
rect 23348 36592 23354 36644
rect 28537 36635 28595 36641
rect 28537 36601 28549 36635
rect 28583 36632 28595 36635
rect 28902 36632 28908 36644
rect 28583 36604 28908 36632
rect 28583 36601 28595 36604
rect 28537 36595 28595 36601
rect 28902 36592 28908 36604
rect 28960 36592 28966 36644
rect 29564 36632 29592 36663
rect 30834 36660 30840 36672
rect 30892 36660 30898 36712
rect 30098 36632 30104 36644
rect 29564 36604 30104 36632
rect 30098 36592 30104 36604
rect 30156 36592 30162 36644
rect 32217 36635 32275 36641
rect 32217 36601 32229 36635
rect 32263 36632 32275 36635
rect 32784 36632 32812 36740
rect 36170 36728 36176 36740
rect 36228 36728 36234 36780
rect 36265 36771 36323 36777
rect 36265 36737 36277 36771
rect 36311 36768 36323 36771
rect 36998 36768 37004 36780
rect 36311 36740 37004 36768
rect 36311 36737 36323 36740
rect 36265 36731 36323 36737
rect 36998 36728 37004 36740
rect 37056 36728 37062 36780
rect 32950 36700 32956 36712
rect 32911 36672 32956 36700
rect 32950 36660 32956 36672
rect 33008 36660 33014 36712
rect 35161 36703 35219 36709
rect 35161 36669 35173 36703
rect 35207 36700 35219 36703
rect 35526 36700 35532 36712
rect 35207 36672 35532 36700
rect 35207 36669 35219 36672
rect 35161 36663 35219 36669
rect 35526 36660 35532 36672
rect 35584 36660 35590 36712
rect 35986 36700 35992 36712
rect 35947 36672 35992 36700
rect 35986 36660 35992 36672
rect 36044 36660 36050 36712
rect 37108 36700 37136 36796
rect 36096 36672 37136 36700
rect 36096 36644 36124 36672
rect 32263 36604 32812 36632
rect 34977 36635 35035 36641
rect 32263 36601 32275 36604
rect 32217 36595 32275 36601
rect 34977 36601 34989 36635
rect 35023 36632 35035 36635
rect 35342 36632 35348 36644
rect 35023 36604 35348 36632
rect 35023 36601 35035 36604
rect 34977 36595 35035 36601
rect 35342 36592 35348 36604
rect 35400 36632 35406 36644
rect 36078 36632 36084 36644
rect 35400 36604 36084 36632
rect 35400 36592 35406 36604
rect 36078 36592 36084 36604
rect 36136 36592 36142 36644
rect 19426 36564 19432 36576
rect 18104 36536 19012 36564
rect 19387 36536 19432 36564
rect 18104 36524 18110 36536
rect 19426 36524 19432 36536
rect 19484 36524 19490 36576
rect 20070 36524 20076 36576
rect 20128 36564 20134 36576
rect 20625 36567 20683 36573
rect 20625 36564 20637 36567
rect 20128 36536 20637 36564
rect 20128 36524 20134 36536
rect 20625 36533 20637 36536
rect 20671 36533 20683 36567
rect 25038 36564 25044 36576
rect 24999 36536 25044 36564
rect 20625 36527 20683 36533
rect 25038 36524 25044 36536
rect 25096 36524 25102 36576
rect 29362 36564 29368 36576
rect 29323 36536 29368 36564
rect 29362 36524 29368 36536
rect 29420 36524 29426 36576
rect 34241 36567 34299 36573
rect 34241 36533 34253 36567
rect 34287 36564 34299 36567
rect 35894 36564 35900 36576
rect 34287 36536 35900 36564
rect 34287 36533 34299 36536
rect 34241 36527 34299 36533
rect 35894 36524 35900 36536
rect 35952 36524 35958 36576
rect 1104 36474 38824 36496
rect 1104 36422 19606 36474
rect 19658 36422 19670 36474
rect 19722 36422 19734 36474
rect 19786 36422 19798 36474
rect 19850 36422 38824 36474
rect 1104 36400 38824 36422
rect 3970 36320 3976 36372
rect 4028 36360 4034 36372
rect 6089 36363 6147 36369
rect 6089 36360 6101 36363
rect 4028 36332 6101 36360
rect 4028 36320 4034 36332
rect 6089 36329 6101 36332
rect 6135 36329 6147 36363
rect 6089 36323 6147 36329
rect 7374 36320 7380 36372
rect 7432 36360 7438 36372
rect 7653 36363 7711 36369
rect 7653 36360 7665 36363
rect 7432 36332 7665 36360
rect 7432 36320 7438 36332
rect 7653 36329 7665 36332
rect 7699 36329 7711 36363
rect 10134 36360 10140 36372
rect 7653 36323 7711 36329
rect 8128 36332 10140 36360
rect 4632 36264 6408 36292
rect 2682 36224 2688 36236
rect 2643 36196 2688 36224
rect 2682 36184 2688 36196
rect 2740 36184 2746 36236
rect 4632 36233 4660 36264
rect 3145 36227 3203 36233
rect 3145 36193 3157 36227
rect 3191 36193 3203 36227
rect 3145 36187 3203 36193
rect 4341 36227 4399 36233
rect 4341 36193 4353 36227
rect 4387 36193 4399 36227
rect 4341 36187 4399 36193
rect 4617 36227 4675 36233
rect 4617 36193 4629 36227
rect 4663 36193 4675 36227
rect 4798 36224 4804 36236
rect 4759 36196 4804 36224
rect 4617 36187 4675 36193
rect 2409 36159 2467 36165
rect 2409 36125 2421 36159
rect 2455 36156 2467 36159
rect 2866 36156 2872 36168
rect 2455 36128 2872 36156
rect 2455 36125 2467 36128
rect 2409 36119 2467 36125
rect 2866 36116 2872 36128
rect 2924 36116 2930 36168
rect 3050 36088 3056 36100
rect 3011 36060 3056 36088
rect 3050 36048 3056 36060
rect 3108 36048 3114 36100
rect 3160 36088 3188 36187
rect 3326 36116 3332 36168
rect 3384 36156 3390 36168
rect 4157 36159 4215 36165
rect 4157 36156 4169 36159
rect 3384 36128 4169 36156
rect 3384 36116 3390 36128
rect 4157 36125 4169 36128
rect 4203 36125 4215 36159
rect 4356 36156 4384 36187
rect 4798 36184 4804 36196
rect 4856 36184 4862 36236
rect 6089 36227 6147 36233
rect 6089 36193 6101 36227
rect 6135 36224 6147 36227
rect 6273 36227 6331 36233
rect 6273 36224 6285 36227
rect 6135 36196 6285 36224
rect 6135 36193 6147 36196
rect 6089 36187 6147 36193
rect 6273 36193 6285 36196
rect 6319 36193 6331 36227
rect 6380 36224 6408 36264
rect 8128 36224 8156 36332
rect 10134 36320 10140 36332
rect 10192 36320 10198 36372
rect 21542 36320 21548 36372
rect 21600 36360 21606 36372
rect 22281 36363 22339 36369
rect 22281 36360 22293 36363
rect 21600 36332 22293 36360
rect 21600 36320 21606 36332
rect 22281 36329 22293 36332
rect 22327 36329 22339 36363
rect 22281 36323 22339 36329
rect 23934 36320 23940 36372
rect 23992 36360 23998 36372
rect 24397 36363 24455 36369
rect 24397 36360 24409 36363
rect 23992 36332 24409 36360
rect 23992 36320 23998 36332
rect 24397 36329 24409 36332
rect 24443 36329 24455 36363
rect 24397 36323 24455 36329
rect 27154 36320 27160 36372
rect 27212 36360 27218 36372
rect 27893 36363 27951 36369
rect 27893 36360 27905 36363
rect 27212 36332 27905 36360
rect 27212 36320 27218 36332
rect 27893 36329 27905 36332
rect 27939 36329 27951 36363
rect 27893 36323 27951 36329
rect 8202 36252 8208 36304
rect 8260 36292 8266 36304
rect 8260 36264 11468 36292
rect 8260 36252 8266 36264
rect 8386 36224 8392 36236
rect 6380 36196 8156 36224
rect 8347 36196 8392 36224
rect 6273 36187 6331 36193
rect 8386 36184 8392 36196
rect 8444 36184 8450 36236
rect 9953 36227 10011 36233
rect 9953 36193 9965 36227
rect 9999 36193 10011 36227
rect 10134 36224 10140 36236
rect 10095 36196 10140 36224
rect 9953 36187 10011 36193
rect 4890 36156 4896 36168
rect 4356 36128 4896 36156
rect 4157 36119 4215 36125
rect 4890 36116 4896 36128
rect 4948 36116 4954 36168
rect 6549 36159 6607 36165
rect 6549 36125 6561 36159
rect 6595 36156 6607 36159
rect 6730 36156 6736 36168
rect 6595 36128 6736 36156
rect 6595 36125 6607 36128
rect 6549 36119 6607 36125
rect 6730 36116 6736 36128
rect 6788 36116 6794 36168
rect 9766 36156 9772 36168
rect 9727 36128 9772 36156
rect 9766 36116 9772 36128
rect 9824 36116 9830 36168
rect 9968 36156 9996 36187
rect 10134 36184 10140 36196
rect 10192 36184 10198 36236
rect 10410 36224 10416 36236
rect 10371 36196 10416 36224
rect 10410 36184 10416 36196
rect 10468 36184 10474 36236
rect 11333 36227 11391 36233
rect 11333 36193 11345 36227
rect 11379 36193 11391 36227
rect 11333 36187 11391 36193
rect 11146 36156 11152 36168
rect 9968 36128 11152 36156
rect 11146 36116 11152 36128
rect 11204 36116 11210 36168
rect 6270 36088 6276 36100
rect 3160 36060 6276 36088
rect 6270 36048 6276 36060
rect 6328 36048 6334 36100
rect 10042 36048 10048 36100
rect 10100 36088 10106 36100
rect 11348 36088 11376 36187
rect 11440 36156 11468 36264
rect 18322 36252 18328 36304
rect 18380 36292 18386 36304
rect 18509 36295 18567 36301
rect 18509 36292 18521 36295
rect 18380 36264 18521 36292
rect 18380 36252 18386 36264
rect 18509 36261 18521 36264
rect 18555 36292 18567 36295
rect 18555 36264 19748 36292
rect 18555 36261 18567 36264
rect 18509 36255 18567 36261
rect 12250 36224 12256 36236
rect 12211 36196 12256 36224
rect 12250 36184 12256 36196
rect 12308 36184 12314 36236
rect 13538 36184 13544 36236
rect 13596 36224 13602 36236
rect 14093 36227 14151 36233
rect 14093 36224 14105 36227
rect 13596 36196 14105 36224
rect 13596 36184 13602 36196
rect 14093 36193 14105 36196
rect 14139 36193 14151 36227
rect 15470 36224 15476 36236
rect 15431 36196 15476 36224
rect 14093 36187 14151 36193
rect 15470 36184 15476 36196
rect 15528 36184 15534 36236
rect 15562 36184 15568 36236
rect 15620 36224 15626 36236
rect 15620 36196 15665 36224
rect 15620 36184 15626 36196
rect 15746 36184 15752 36236
rect 15804 36224 15810 36236
rect 16853 36227 16911 36233
rect 16853 36224 16865 36227
rect 15804 36196 16865 36224
rect 15804 36184 15810 36196
rect 16853 36193 16865 36196
rect 16899 36224 16911 36227
rect 18046 36224 18052 36236
rect 16899 36196 18052 36224
rect 16899 36193 16911 36196
rect 16853 36187 16911 36193
rect 18046 36184 18052 36196
rect 18104 36184 18110 36236
rect 19426 36224 19432 36236
rect 19387 36196 19432 36224
rect 19426 36184 19432 36196
rect 19484 36184 19490 36236
rect 19720 36233 19748 36264
rect 29564 36264 32904 36292
rect 19705 36227 19763 36233
rect 19705 36193 19717 36227
rect 19751 36193 19763 36227
rect 20070 36224 20076 36236
rect 20031 36196 20076 36224
rect 19705 36187 19763 36193
rect 20070 36184 20076 36196
rect 20128 36184 20134 36236
rect 20806 36184 20812 36236
rect 20864 36224 20870 36236
rect 21177 36227 21235 36233
rect 21177 36224 21189 36227
rect 20864 36196 21189 36224
rect 20864 36184 20870 36196
rect 21177 36193 21189 36196
rect 21223 36193 21235 36227
rect 23290 36224 23296 36236
rect 23251 36196 23296 36224
rect 21177 36187 21235 36193
rect 23290 36184 23296 36196
rect 23348 36184 23354 36236
rect 26234 36184 26240 36236
rect 26292 36224 26298 36236
rect 26789 36227 26847 36233
rect 26789 36224 26801 36227
rect 26292 36196 26801 36224
rect 26292 36184 26298 36196
rect 26789 36193 26801 36196
rect 26835 36193 26847 36227
rect 28902 36224 28908 36236
rect 28863 36196 28908 36224
rect 26789 36187 26847 36193
rect 28902 36184 28908 36196
rect 28960 36184 28966 36236
rect 11977 36159 12035 36165
rect 11977 36156 11989 36159
rect 11440 36128 11989 36156
rect 11977 36125 11989 36128
rect 12023 36156 12035 36159
rect 12434 36156 12440 36168
rect 12023 36128 12440 36156
rect 12023 36125 12035 36128
rect 11977 36119 12035 36125
rect 12434 36116 12440 36128
rect 12492 36116 12498 36168
rect 13633 36159 13691 36165
rect 13633 36125 13645 36159
rect 13679 36156 13691 36159
rect 14182 36156 14188 36168
rect 13679 36128 14188 36156
rect 13679 36125 13691 36128
rect 13633 36119 13691 36125
rect 14182 36116 14188 36128
rect 14240 36116 14246 36168
rect 17034 36116 17040 36168
rect 17092 36156 17098 36168
rect 17129 36159 17187 36165
rect 17129 36156 17141 36159
rect 17092 36128 17141 36156
rect 17092 36116 17098 36128
rect 17129 36125 17141 36128
rect 17175 36125 17187 36159
rect 17129 36119 17187 36125
rect 19150 36116 19156 36168
rect 19208 36156 19214 36168
rect 20901 36159 20959 36165
rect 20901 36156 20913 36159
rect 19208 36128 20913 36156
rect 19208 36116 19214 36128
rect 20901 36125 20913 36128
rect 20947 36125 20959 36159
rect 23014 36156 23020 36168
rect 22975 36128 23020 36156
rect 20901 36119 20959 36125
rect 23014 36116 23020 36128
rect 23072 36116 23078 36168
rect 26510 36156 26516 36168
rect 26471 36128 26516 36156
rect 26510 36116 26516 36128
rect 26568 36156 26574 36168
rect 28629 36159 28687 36165
rect 28629 36156 28641 36159
rect 26568 36128 28641 36156
rect 26568 36116 26574 36128
rect 28629 36125 28641 36128
rect 28675 36156 28687 36159
rect 28994 36156 29000 36168
rect 28675 36128 29000 36156
rect 28675 36125 28687 36128
rect 28629 36119 28687 36125
rect 28994 36116 29000 36128
rect 29052 36116 29058 36168
rect 10100 36060 11376 36088
rect 10100 36048 10106 36060
rect 8478 36020 8484 36032
rect 8439 35992 8484 36020
rect 8478 35980 8484 35992
rect 8536 35980 8542 36032
rect 9674 35980 9680 36032
rect 9732 36020 9738 36032
rect 11425 36023 11483 36029
rect 11425 36020 11437 36023
rect 9732 35992 11437 36020
rect 9732 35980 9738 35992
rect 11425 35989 11437 35992
rect 11471 35989 11483 36023
rect 11425 35983 11483 35989
rect 13906 35980 13912 36032
rect 13964 36020 13970 36032
rect 14185 36023 14243 36029
rect 14185 36020 14197 36023
rect 13964 35992 14197 36020
rect 13964 35980 13970 35992
rect 14185 35989 14197 35992
rect 14231 35989 14243 36023
rect 14185 35983 14243 35989
rect 14274 35980 14280 36032
rect 14332 36020 14338 36032
rect 15289 36023 15347 36029
rect 15289 36020 15301 36023
rect 14332 35992 15301 36020
rect 14332 35980 14338 35992
rect 15289 35989 15301 35992
rect 15335 35989 15347 36023
rect 15746 36020 15752 36032
rect 15707 35992 15752 36020
rect 15289 35983 15347 35989
rect 15746 35980 15752 35992
rect 15804 35980 15810 36032
rect 20349 36023 20407 36029
rect 20349 35989 20361 36023
rect 20395 36020 20407 36023
rect 29564 36020 29592 36264
rect 31113 36227 31171 36233
rect 31113 36193 31125 36227
rect 31159 36224 31171 36227
rect 32306 36224 32312 36236
rect 31159 36196 32312 36224
rect 31159 36193 31171 36196
rect 31113 36187 31171 36193
rect 32306 36184 32312 36196
rect 32364 36184 32370 36236
rect 32876 36233 32904 36264
rect 32950 36252 32956 36304
rect 33008 36292 33014 36304
rect 37185 36295 37243 36301
rect 37185 36292 37197 36295
rect 33008 36264 37197 36292
rect 33008 36252 33014 36264
rect 37185 36261 37197 36264
rect 37231 36261 37243 36295
rect 37185 36255 37243 36261
rect 32861 36227 32919 36233
rect 32861 36193 32873 36227
rect 32907 36224 32919 36227
rect 33134 36224 33140 36236
rect 32907 36196 33140 36224
rect 32907 36193 32919 36196
rect 32861 36187 32919 36193
rect 33134 36184 33140 36196
rect 33192 36184 33198 36236
rect 33413 36227 33471 36233
rect 33413 36193 33425 36227
rect 33459 36224 33471 36227
rect 34698 36224 34704 36236
rect 33459 36196 34704 36224
rect 33459 36193 33471 36196
rect 33413 36187 33471 36193
rect 34698 36184 34704 36196
rect 34756 36184 34762 36236
rect 35069 36227 35127 36233
rect 35069 36193 35081 36227
rect 35115 36193 35127 36227
rect 35342 36224 35348 36236
rect 35303 36196 35348 36224
rect 35069 36187 35127 36193
rect 33502 36156 33508 36168
rect 33463 36128 33508 36156
rect 33502 36116 33508 36128
rect 33560 36116 33566 36168
rect 35084 36156 35112 36187
rect 35342 36184 35348 36196
rect 35400 36184 35406 36236
rect 35526 36224 35532 36236
rect 35487 36196 35532 36224
rect 35526 36184 35532 36196
rect 35584 36184 35590 36236
rect 35618 36184 35624 36236
rect 35676 36224 35682 36236
rect 35989 36227 36047 36233
rect 35989 36224 36001 36227
rect 35676 36196 36001 36224
rect 35676 36184 35682 36196
rect 35989 36193 36001 36196
rect 36035 36224 36047 36227
rect 36633 36227 36691 36233
rect 36633 36224 36645 36227
rect 36035 36196 36645 36224
rect 36035 36193 36047 36196
rect 35989 36187 36047 36193
rect 36633 36193 36645 36196
rect 36679 36193 36691 36227
rect 36633 36187 36691 36193
rect 36722 36184 36728 36236
rect 36780 36224 36786 36236
rect 37737 36227 37795 36233
rect 36780 36196 36825 36224
rect 36780 36184 36786 36196
rect 37737 36193 37749 36227
rect 37783 36193 37795 36227
rect 37737 36187 37795 36193
rect 35894 36156 35900 36168
rect 35084 36128 35900 36156
rect 35894 36116 35900 36128
rect 35952 36116 35958 36168
rect 36446 36156 36452 36168
rect 36407 36128 36452 36156
rect 36446 36116 36452 36128
rect 36504 36116 36510 36168
rect 33410 36088 33416 36100
rect 33371 36060 33416 36088
rect 33410 36048 33416 36060
rect 33468 36048 33474 36100
rect 34514 36048 34520 36100
rect 34572 36088 34578 36100
rect 37752 36088 37780 36187
rect 34572 36060 37780 36088
rect 34572 36048 34578 36060
rect 30006 36020 30012 36032
rect 20395 35992 29592 36020
rect 29967 35992 30012 36020
rect 20395 35989 20407 35992
rect 20349 35983 20407 35989
rect 30006 35980 30012 35992
rect 30064 35980 30070 36032
rect 30374 35980 30380 36032
rect 30432 36020 30438 36032
rect 31205 36023 31263 36029
rect 31205 36020 31217 36023
rect 30432 35992 31217 36020
rect 30432 35980 30438 35992
rect 31205 35989 31217 35992
rect 31251 35989 31263 36023
rect 31205 35983 31263 35989
rect 37090 35980 37096 36032
rect 37148 36020 37154 36032
rect 37829 36023 37887 36029
rect 37829 36020 37841 36023
rect 37148 35992 37841 36020
rect 37148 35980 37154 35992
rect 37829 35989 37841 35992
rect 37875 35989 37887 36023
rect 37829 35983 37887 35989
rect 1104 35930 38824 35952
rect 1104 35878 4246 35930
rect 4298 35878 4310 35930
rect 4362 35878 4374 35930
rect 4426 35878 4438 35930
rect 4490 35878 34966 35930
rect 35018 35878 35030 35930
rect 35082 35878 35094 35930
rect 35146 35878 35158 35930
rect 35210 35878 38824 35930
rect 1104 35856 38824 35878
rect 20806 35816 20812 35828
rect 20767 35788 20812 35816
rect 20806 35776 20812 35788
rect 20864 35776 20870 35828
rect 21266 35776 21272 35828
rect 21324 35816 21330 35828
rect 21361 35819 21419 35825
rect 21361 35816 21373 35819
rect 21324 35788 21373 35816
rect 21324 35776 21330 35788
rect 21361 35785 21373 35788
rect 21407 35785 21419 35819
rect 21361 35779 21419 35785
rect 24946 35776 24952 35828
rect 25004 35816 25010 35828
rect 25317 35819 25375 35825
rect 25317 35816 25329 35819
rect 25004 35788 25329 35816
rect 25004 35776 25010 35788
rect 25317 35785 25329 35788
rect 25363 35785 25375 35819
rect 27617 35819 27675 35825
rect 25317 35779 25375 35785
rect 25976 35788 27016 35816
rect 5626 35748 5632 35760
rect 5368 35720 5632 35748
rect 2133 35683 2191 35689
rect 2133 35649 2145 35683
rect 2179 35680 2191 35683
rect 3970 35680 3976 35692
rect 2179 35652 3976 35680
rect 2179 35649 2191 35652
rect 2133 35643 2191 35649
rect 3970 35640 3976 35652
rect 4028 35640 4034 35692
rect 2222 35572 2228 35624
rect 2280 35612 2286 35624
rect 2409 35615 2467 35621
rect 2409 35612 2421 35615
rect 2280 35584 2421 35612
rect 2280 35572 2286 35584
rect 2409 35581 2421 35584
rect 2455 35581 2467 35615
rect 2409 35575 2467 35581
rect 5077 35615 5135 35621
rect 5077 35581 5089 35615
rect 5123 35612 5135 35615
rect 5368 35612 5396 35720
rect 5626 35708 5632 35720
rect 5684 35708 5690 35760
rect 23014 35708 23020 35760
rect 23072 35748 23078 35760
rect 23072 35720 23980 35748
rect 23072 35708 23078 35720
rect 5442 35640 5448 35692
rect 5500 35680 5506 35692
rect 5721 35683 5779 35689
rect 5721 35680 5733 35683
rect 5500 35652 5733 35680
rect 5500 35640 5506 35652
rect 5721 35649 5733 35652
rect 5767 35680 5779 35683
rect 8478 35680 8484 35692
rect 5767 35652 7328 35680
rect 5767 35649 5779 35652
rect 5721 35643 5779 35649
rect 5123 35584 5396 35612
rect 5629 35615 5687 35621
rect 5123 35581 5135 35584
rect 5077 35575 5135 35581
rect 5629 35581 5641 35615
rect 5675 35581 5687 35615
rect 6914 35612 6920 35624
rect 6875 35584 6920 35612
rect 5629 35575 5687 35581
rect 3789 35547 3847 35553
rect 3789 35513 3801 35547
rect 3835 35544 3847 35547
rect 5534 35544 5540 35556
rect 3835 35516 5540 35544
rect 3835 35513 3847 35516
rect 3789 35507 3847 35513
rect 5534 35504 5540 35516
rect 5592 35504 5598 35556
rect 5644 35544 5672 35575
rect 6914 35572 6920 35584
rect 6972 35572 6978 35624
rect 7300 35621 7328 35652
rect 7852 35652 8484 35680
rect 7852 35621 7880 35652
rect 8478 35640 8484 35652
rect 8536 35640 8542 35692
rect 9401 35683 9459 35689
rect 9401 35649 9413 35683
rect 9447 35680 9459 35683
rect 10410 35680 10416 35692
rect 9447 35652 10416 35680
rect 9447 35649 9459 35652
rect 9401 35643 9459 35649
rect 10410 35640 10416 35652
rect 10468 35640 10474 35692
rect 11146 35680 11152 35692
rect 11107 35652 11152 35680
rect 11146 35640 11152 35652
rect 11204 35640 11210 35692
rect 14553 35683 14611 35689
rect 14553 35649 14565 35683
rect 14599 35680 14611 35683
rect 15746 35680 15752 35692
rect 14599 35652 15752 35680
rect 14599 35649 14611 35652
rect 14553 35643 14611 35649
rect 15746 35640 15752 35652
rect 15804 35640 15810 35692
rect 16393 35683 16451 35689
rect 16393 35649 16405 35683
rect 16439 35680 16451 35683
rect 16439 35652 17908 35680
rect 16439 35649 16451 35652
rect 16393 35643 16451 35649
rect 17880 35624 17908 35652
rect 18340 35652 19380 35680
rect 7285 35615 7343 35621
rect 7285 35581 7297 35615
rect 7331 35581 7343 35615
rect 7285 35575 7343 35581
rect 7837 35615 7895 35621
rect 7837 35581 7849 35615
rect 7883 35581 7895 35615
rect 7837 35575 7895 35581
rect 8021 35615 8079 35621
rect 8021 35581 8033 35615
rect 8067 35581 8079 35615
rect 8021 35575 8079 35581
rect 9309 35615 9367 35621
rect 9309 35581 9321 35615
rect 9355 35581 9367 35615
rect 9309 35575 9367 35581
rect 9769 35615 9827 35621
rect 9769 35581 9781 35615
rect 9815 35612 9827 35615
rect 9950 35612 9956 35624
rect 9815 35584 9956 35612
rect 9815 35581 9827 35584
rect 9769 35575 9827 35581
rect 6454 35544 6460 35556
rect 5644 35516 6460 35544
rect 6454 35504 6460 35516
rect 6512 35544 6518 35556
rect 8036 35544 8064 35575
rect 6512 35516 8064 35544
rect 9324 35544 9352 35575
rect 9950 35572 9956 35584
rect 10008 35572 10014 35624
rect 10042 35572 10048 35624
rect 10100 35612 10106 35624
rect 10229 35615 10287 35621
rect 10229 35612 10241 35615
rect 10100 35584 10241 35612
rect 10100 35572 10106 35584
rect 10229 35581 10241 35584
rect 10275 35581 10287 35615
rect 10870 35612 10876 35624
rect 10831 35584 10876 35612
rect 10229 35575 10287 35581
rect 10870 35572 10876 35584
rect 10928 35572 10934 35624
rect 11054 35612 11060 35624
rect 11015 35584 11060 35612
rect 11054 35572 11060 35584
rect 11112 35572 11118 35624
rect 11514 35612 11520 35624
rect 11475 35584 11520 35612
rect 11514 35572 11520 35584
rect 11572 35572 11578 35624
rect 12437 35615 12495 35621
rect 12437 35581 12449 35615
rect 12483 35581 12495 35615
rect 12437 35575 12495 35581
rect 9674 35544 9680 35556
rect 9324 35516 9680 35544
rect 6512 35504 6518 35516
rect 9674 35504 9680 35516
rect 9732 35504 9738 35556
rect 12452 35544 12480 35575
rect 12526 35572 12532 35624
rect 12584 35612 12590 35624
rect 13081 35615 13139 35621
rect 13081 35612 13093 35615
rect 12584 35584 13093 35612
rect 12584 35572 12590 35584
rect 13081 35581 13093 35584
rect 13127 35581 13139 35615
rect 13538 35612 13544 35624
rect 13499 35584 13544 35612
rect 13081 35575 13139 35581
rect 13538 35572 13544 35584
rect 13596 35572 13602 35624
rect 13998 35612 14004 35624
rect 13648 35584 14004 35612
rect 13648 35544 13676 35584
rect 13998 35572 14004 35584
rect 14056 35572 14062 35624
rect 14277 35615 14335 35621
rect 14277 35581 14289 35615
rect 14323 35612 14335 35615
rect 15838 35612 15844 35624
rect 14323 35584 15844 35612
rect 14323 35581 14335 35584
rect 14277 35575 14335 35581
rect 15838 35572 15844 35584
rect 15896 35572 15902 35624
rect 16482 35572 16488 35624
rect 16540 35612 16546 35624
rect 16540 35584 16585 35612
rect 16540 35572 16546 35584
rect 17862 35572 17868 35624
rect 17920 35612 17926 35624
rect 18340 35621 18368 35652
rect 18233 35615 18291 35621
rect 18233 35612 18245 35615
rect 17920 35584 18245 35612
rect 17920 35572 17926 35584
rect 18233 35581 18245 35584
rect 18279 35581 18291 35615
rect 18233 35575 18291 35581
rect 18325 35615 18383 35621
rect 18325 35581 18337 35615
rect 18371 35581 18383 35615
rect 18325 35575 18383 35581
rect 19150 35572 19156 35624
rect 19208 35612 19214 35624
rect 19245 35615 19303 35621
rect 19245 35612 19257 35615
rect 19208 35584 19257 35612
rect 19208 35572 19214 35584
rect 19245 35581 19257 35584
rect 19291 35581 19303 35615
rect 19352 35612 19380 35652
rect 19426 35640 19432 35692
rect 19484 35680 19490 35692
rect 23952 35689 23980 35720
rect 19521 35683 19579 35689
rect 19521 35680 19533 35683
rect 19484 35652 19533 35680
rect 19484 35640 19490 35652
rect 19521 35649 19533 35652
rect 19567 35649 19579 35683
rect 23937 35683 23995 35689
rect 19521 35643 19579 35649
rect 20180 35652 23428 35680
rect 20180 35612 20208 35652
rect 21542 35612 21548 35624
rect 19352 35584 20208 35612
rect 21503 35584 21548 35612
rect 19245 35575 19303 35581
rect 21542 35572 21548 35584
rect 21600 35572 21606 35624
rect 22097 35615 22155 35621
rect 22097 35581 22109 35615
rect 22143 35581 22155 35615
rect 22097 35575 22155 35581
rect 22189 35615 22247 35621
rect 22189 35581 22201 35615
rect 22235 35581 22247 35615
rect 23400 35612 23428 35652
rect 23937 35649 23949 35683
rect 23983 35649 23995 35683
rect 23937 35643 23995 35649
rect 24213 35683 24271 35689
rect 24213 35649 24225 35683
rect 24259 35680 24271 35683
rect 25038 35680 25044 35692
rect 24259 35652 25044 35680
rect 24259 35649 24271 35652
rect 24213 35643 24271 35649
rect 25038 35640 25044 35652
rect 25096 35640 25102 35692
rect 25976 35612 26004 35788
rect 26988 35748 27016 35788
rect 27617 35785 27629 35819
rect 27663 35816 27675 35819
rect 27982 35816 27988 35828
rect 27663 35788 27988 35816
rect 27663 35785 27675 35788
rect 27617 35779 27675 35785
rect 27982 35776 27988 35788
rect 28040 35776 28046 35828
rect 28905 35819 28963 35825
rect 28905 35785 28917 35819
rect 28951 35816 28963 35819
rect 28994 35816 29000 35828
rect 28951 35788 29000 35816
rect 28951 35785 28963 35788
rect 28905 35779 28963 35785
rect 28994 35776 29000 35788
rect 29052 35776 29058 35828
rect 29914 35816 29920 35828
rect 29104 35788 29920 35816
rect 29104 35748 29132 35788
rect 29914 35776 29920 35788
rect 29972 35776 29978 35828
rect 32953 35819 33011 35825
rect 32953 35785 32965 35819
rect 32999 35816 33011 35819
rect 38286 35816 38292 35828
rect 32999 35788 38292 35816
rect 32999 35785 33011 35788
rect 32953 35779 33011 35785
rect 38286 35776 38292 35788
rect 38344 35776 38350 35828
rect 34238 35748 34244 35760
rect 26988 35720 29132 35748
rect 32968 35720 34244 35748
rect 26053 35683 26111 35689
rect 26053 35649 26065 35683
rect 26099 35680 26111 35683
rect 26510 35680 26516 35692
rect 26099 35652 26516 35680
rect 26099 35649 26111 35652
rect 26053 35643 26111 35649
rect 26510 35640 26516 35652
rect 26568 35640 26574 35692
rect 28902 35640 28908 35692
rect 28960 35680 28966 35692
rect 29273 35683 29331 35689
rect 29273 35680 29285 35683
rect 28960 35652 29285 35680
rect 28960 35640 28966 35652
rect 29273 35649 29285 35652
rect 29319 35649 29331 35683
rect 29273 35643 29331 35649
rect 29549 35683 29607 35689
rect 29549 35649 29561 35683
rect 29595 35680 29607 35683
rect 30006 35680 30012 35692
rect 29595 35652 30012 35680
rect 29595 35649 29607 35652
rect 29549 35643 29607 35649
rect 30006 35640 30012 35652
rect 30064 35640 30070 35692
rect 32968 35680 32996 35720
rect 34238 35708 34244 35720
rect 34296 35708 34302 35760
rect 34698 35708 34704 35760
rect 34756 35748 34762 35760
rect 34977 35751 35035 35757
rect 34977 35748 34989 35751
rect 34756 35720 34989 35748
rect 34756 35708 34762 35720
rect 34977 35717 34989 35720
rect 35023 35717 35035 35751
rect 34977 35711 35035 35717
rect 35713 35683 35771 35689
rect 35713 35680 35725 35683
rect 30116 35652 32996 35680
rect 33888 35652 35725 35680
rect 26326 35612 26332 35624
rect 23400 35584 26004 35612
rect 26287 35584 26332 35612
rect 22189 35575 22247 35581
rect 13814 35544 13820 35556
rect 12452 35516 13676 35544
rect 13775 35516 13820 35544
rect 13814 35504 13820 35516
rect 13872 35504 13878 35556
rect 16114 35504 16120 35556
rect 16172 35544 16178 35556
rect 16945 35547 17003 35553
rect 16945 35544 16957 35547
rect 16172 35516 16957 35544
rect 16172 35504 16178 35516
rect 16945 35513 16957 35516
rect 16991 35513 17003 35547
rect 16945 35507 17003 35513
rect 18785 35547 18843 35553
rect 18785 35513 18797 35547
rect 18831 35544 18843 35547
rect 18966 35544 18972 35556
rect 18831 35516 18972 35544
rect 18831 35513 18843 35516
rect 18785 35507 18843 35513
rect 18966 35504 18972 35516
rect 19024 35504 19030 35556
rect 20806 35504 20812 35556
rect 20864 35544 20870 35556
rect 22112 35544 22140 35575
rect 20864 35516 22140 35544
rect 20864 35504 20870 35516
rect 4706 35436 4712 35488
rect 4764 35476 4770 35488
rect 4893 35479 4951 35485
rect 4893 35476 4905 35479
rect 4764 35448 4905 35476
rect 4764 35436 4770 35448
rect 4893 35445 4905 35448
rect 4939 35476 4951 35479
rect 5258 35476 5264 35488
rect 4939 35448 5264 35476
rect 4939 35445 4951 35448
rect 4893 35439 4951 35445
rect 5258 35436 5264 35448
rect 5316 35436 5322 35488
rect 5350 35436 5356 35488
rect 5408 35476 5414 35488
rect 7742 35476 7748 35488
rect 5408 35448 7748 35476
rect 5408 35436 5414 35448
rect 7742 35436 7748 35448
rect 7800 35436 7806 35488
rect 8018 35476 8024 35488
rect 7979 35448 8024 35476
rect 8018 35436 8024 35448
rect 8076 35436 8082 35488
rect 13354 35436 13360 35488
rect 13412 35476 13418 35488
rect 15657 35479 15715 35485
rect 15657 35476 15669 35479
rect 13412 35448 15669 35476
rect 13412 35436 13418 35448
rect 15657 35445 15669 35448
rect 15703 35445 15715 35479
rect 22204 35476 22232 35575
rect 26326 35572 26332 35584
rect 26384 35572 26390 35624
rect 29086 35612 29092 35624
rect 29047 35584 29092 35612
rect 29086 35572 29092 35584
rect 29144 35572 29150 35624
rect 30116 35612 30144 35652
rect 29380 35584 30144 35612
rect 22646 35544 22652 35556
rect 22607 35516 22652 35544
rect 22646 35504 22652 35516
rect 22704 35504 22710 35556
rect 29380 35544 29408 35584
rect 30282 35572 30288 35624
rect 30340 35612 30346 35624
rect 31389 35615 31447 35621
rect 31389 35612 31401 35615
rect 30340 35584 31401 35612
rect 30340 35572 30346 35584
rect 31389 35581 31401 35584
rect 31435 35581 31447 35615
rect 31665 35615 31723 35621
rect 31665 35612 31677 35615
rect 31389 35575 31447 35581
rect 31496 35584 31677 35612
rect 26988 35516 29408 35544
rect 26988 35476 27016 35516
rect 30650 35476 30656 35488
rect 22204 35448 27016 35476
rect 30611 35448 30656 35476
rect 15657 35439 15715 35445
rect 30650 35436 30656 35448
rect 30708 35436 30714 35488
rect 31110 35436 31116 35488
rect 31168 35476 31174 35488
rect 31205 35479 31263 35485
rect 31205 35476 31217 35479
rect 31168 35448 31217 35476
rect 31168 35436 31174 35448
rect 31205 35445 31217 35448
rect 31251 35476 31263 35479
rect 31496 35476 31524 35584
rect 31665 35581 31677 35584
rect 31711 35581 31723 35615
rect 31665 35575 31723 35581
rect 33778 35572 33784 35624
rect 33836 35612 33842 35624
rect 33888 35621 33916 35652
rect 35713 35649 35725 35652
rect 35759 35649 35771 35683
rect 35713 35643 35771 35649
rect 35986 35640 35992 35692
rect 36044 35680 36050 35692
rect 36449 35683 36507 35689
rect 36449 35680 36461 35683
rect 36044 35652 36461 35680
rect 36044 35640 36050 35652
rect 36449 35649 36461 35652
rect 36495 35649 36507 35683
rect 36449 35643 36507 35649
rect 36725 35683 36783 35689
rect 36725 35649 36737 35683
rect 36771 35680 36783 35683
rect 37090 35680 37096 35692
rect 36771 35652 37096 35680
rect 36771 35649 36783 35652
rect 36725 35643 36783 35649
rect 37090 35640 37096 35652
rect 37148 35640 37154 35692
rect 33873 35615 33931 35621
rect 33873 35612 33885 35615
rect 33836 35584 33885 35612
rect 33836 35572 33842 35584
rect 33873 35581 33885 35584
rect 33919 35581 33931 35615
rect 34146 35612 34152 35624
rect 34107 35584 34152 35612
rect 33873 35575 33931 35581
rect 34146 35572 34152 35584
rect 34204 35572 34210 35624
rect 34333 35615 34391 35621
rect 34333 35581 34345 35615
rect 34379 35612 34391 35615
rect 34885 35615 34943 35621
rect 34885 35612 34897 35615
rect 34379 35584 34897 35612
rect 34379 35581 34391 35584
rect 34333 35575 34391 35581
rect 34885 35581 34897 35584
rect 34931 35581 34943 35615
rect 35618 35612 35624 35624
rect 35579 35584 35624 35612
rect 34885 35575 34943 35581
rect 35618 35572 35624 35584
rect 35676 35572 35682 35624
rect 31251 35448 31524 35476
rect 31251 35445 31263 35448
rect 31205 35439 31263 35445
rect 35802 35436 35808 35488
rect 35860 35476 35866 35488
rect 37829 35479 37887 35485
rect 37829 35476 37841 35479
rect 35860 35448 37841 35476
rect 35860 35436 35866 35448
rect 37829 35445 37841 35448
rect 37875 35445 37887 35479
rect 37829 35439 37887 35445
rect 1104 35386 38824 35408
rect 1104 35334 19606 35386
rect 19658 35334 19670 35386
rect 19722 35334 19734 35386
rect 19786 35334 19798 35386
rect 19850 35334 38824 35386
rect 1104 35312 38824 35334
rect 2222 35272 2228 35284
rect 2183 35244 2228 35272
rect 2222 35232 2228 35244
rect 2280 35232 2286 35284
rect 3418 35232 3424 35284
rect 3476 35272 3482 35284
rect 3476 35244 8340 35272
rect 3476 35232 3482 35244
rect 3050 35204 3056 35216
rect 2332 35176 3056 35204
rect 2332 35145 2360 35176
rect 3050 35164 3056 35176
rect 3108 35164 3114 35216
rect 5258 35164 5264 35216
rect 5316 35204 5322 35216
rect 8312 35204 8340 35244
rect 8386 35232 8392 35284
rect 8444 35272 8450 35284
rect 8665 35275 8723 35281
rect 8665 35272 8677 35275
rect 8444 35244 8677 35272
rect 8444 35232 8450 35244
rect 8665 35241 8677 35244
rect 8711 35241 8723 35275
rect 16482 35272 16488 35284
rect 8665 35235 8723 35241
rect 10152 35244 16488 35272
rect 10042 35204 10048 35216
rect 5316 35176 7236 35204
rect 8312 35176 10048 35204
rect 5316 35164 5322 35176
rect 1397 35139 1455 35145
rect 1397 35105 1409 35139
rect 1443 35105 1455 35139
rect 1397 35099 1455 35105
rect 2317 35139 2375 35145
rect 2317 35105 2329 35139
rect 2363 35105 2375 35139
rect 2866 35136 2872 35148
rect 2779 35108 2872 35136
rect 2317 35099 2375 35105
rect 1412 35000 1440 35099
rect 2866 35096 2872 35108
rect 2924 35136 2930 35148
rect 4617 35139 4675 35145
rect 2924 35108 4292 35136
rect 2924 35096 2930 35108
rect 2682 35028 2688 35080
rect 2740 35068 2746 35080
rect 4264 35077 4292 35108
rect 4617 35105 4629 35139
rect 4663 35136 4675 35139
rect 4706 35136 4712 35148
rect 4663 35108 4712 35136
rect 4663 35105 4675 35108
rect 4617 35099 4675 35105
rect 4706 35096 4712 35108
rect 4764 35096 4770 35148
rect 4985 35139 5043 35145
rect 4985 35105 4997 35139
rect 5031 35136 5043 35139
rect 5442 35136 5448 35148
rect 5031 35108 5448 35136
rect 5031 35105 5043 35108
rect 4985 35099 5043 35105
rect 5442 35096 5448 35108
rect 5500 35096 5506 35148
rect 5626 35096 5632 35148
rect 5684 35136 5690 35148
rect 5905 35139 5963 35145
rect 5905 35136 5917 35139
rect 5684 35108 5917 35136
rect 5684 35096 5690 35108
rect 5905 35105 5917 35108
rect 5951 35105 5963 35139
rect 6454 35136 6460 35148
rect 6415 35108 6460 35136
rect 5905 35099 5963 35105
rect 6454 35096 6460 35108
rect 6512 35096 6518 35148
rect 3145 35071 3203 35077
rect 3145 35068 3157 35071
rect 2740 35040 3157 35068
rect 2740 35028 2746 35040
rect 3145 35037 3157 35040
rect 3191 35037 3203 35071
rect 3145 35031 3203 35037
rect 4249 35071 4307 35077
rect 4249 35037 4261 35071
rect 4295 35068 4307 35071
rect 5644 35068 5672 35096
rect 4295 35040 5672 35068
rect 4295 35037 4307 35040
rect 4249 35031 4307 35037
rect 3160 35000 3188 35031
rect 4706 35000 4712 35012
rect 1412 34972 2912 35000
rect 3160 34972 4712 35000
rect 1581 34935 1639 34941
rect 1581 34901 1593 34935
rect 1627 34932 1639 34935
rect 1670 34932 1676 34944
rect 1627 34904 1676 34932
rect 1627 34901 1639 34904
rect 1581 34895 1639 34901
rect 1670 34892 1676 34904
rect 1728 34932 1734 34944
rect 2682 34932 2688 34944
rect 1728 34904 2688 34932
rect 1728 34892 1734 34904
rect 2682 34892 2688 34904
rect 2740 34892 2746 34944
rect 2884 34932 2912 34972
rect 4706 34960 4712 34972
rect 4764 34960 4770 35012
rect 4890 35000 4896 35012
rect 4851 34972 4896 35000
rect 4890 34960 4896 34972
rect 4948 34960 4954 35012
rect 3786 34932 3792 34944
rect 2884 34904 3792 34932
rect 3786 34892 3792 34904
rect 3844 34932 3850 34944
rect 6472 34932 6500 35096
rect 6641 35071 6699 35077
rect 6641 35037 6653 35071
rect 6687 35068 6699 35071
rect 7006 35068 7012 35080
rect 6687 35040 7012 35068
rect 6687 35037 6699 35040
rect 6641 35031 6699 35037
rect 7006 35028 7012 35040
rect 7064 35028 7070 35080
rect 3844 34904 6500 34932
rect 7208 34932 7236 35176
rect 10042 35164 10048 35176
rect 10100 35164 10106 35216
rect 7285 35139 7343 35145
rect 7285 35105 7297 35139
rect 7331 35136 7343 35139
rect 7374 35136 7380 35148
rect 7331 35108 7380 35136
rect 7331 35105 7343 35108
rect 7285 35099 7343 35105
rect 7374 35096 7380 35108
rect 7432 35096 7438 35148
rect 9674 35096 9680 35148
rect 9732 35136 9738 35148
rect 9732 35108 9777 35136
rect 9732 35096 9738 35108
rect 7558 35068 7564 35080
rect 7519 35040 7564 35068
rect 7558 35028 7564 35040
rect 7616 35028 7622 35080
rect 7742 35028 7748 35080
rect 7800 35068 7806 35080
rect 10152 35068 10180 35244
rect 16482 35232 16488 35244
rect 16540 35232 16546 35284
rect 18874 35272 18880 35284
rect 17236 35244 18880 35272
rect 10226 35164 10232 35216
rect 10284 35204 10290 35216
rect 10284 35176 10824 35204
rect 10284 35164 10290 35176
rect 10796 35148 10824 35176
rect 10870 35164 10876 35216
rect 10928 35204 10934 35216
rect 13354 35204 13360 35216
rect 10928 35176 13360 35204
rect 10928 35164 10934 35176
rect 10318 35096 10324 35148
rect 10376 35136 10382 35148
rect 10689 35139 10747 35145
rect 10689 35136 10701 35139
rect 10376 35108 10701 35136
rect 10376 35096 10382 35108
rect 10689 35105 10701 35108
rect 10735 35105 10747 35139
rect 10689 35099 10747 35105
rect 10778 35096 10784 35148
rect 10836 35136 10842 35148
rect 11057 35139 11115 35145
rect 11057 35136 11069 35139
rect 10836 35108 11069 35136
rect 10836 35096 10842 35108
rect 11057 35105 11069 35108
rect 11103 35105 11115 35139
rect 11422 35136 11428 35148
rect 11383 35108 11428 35136
rect 11057 35099 11115 35105
rect 11422 35096 11428 35108
rect 11480 35096 11486 35148
rect 11514 35096 11520 35148
rect 11572 35136 11578 35148
rect 12618 35136 12624 35148
rect 11572 35108 12624 35136
rect 11572 35096 11578 35108
rect 12618 35096 12624 35108
rect 12676 35136 12682 35148
rect 13188 35145 13216 35176
rect 13354 35164 13360 35176
rect 13412 35164 13418 35216
rect 14093 35207 14151 35213
rect 14093 35204 14105 35207
rect 13648 35176 14105 35204
rect 13173 35139 13231 35145
rect 12676 35108 13124 35136
rect 12676 35096 12682 35108
rect 11698 35068 11704 35080
rect 7800 35040 10180 35068
rect 11659 35040 11704 35068
rect 7800 35028 7806 35040
rect 11698 35028 11704 35040
rect 11756 35028 11762 35080
rect 13096 35068 13124 35108
rect 13173 35105 13185 35139
rect 13219 35105 13231 35139
rect 13173 35099 13231 35105
rect 13265 35139 13323 35145
rect 13265 35105 13277 35139
rect 13311 35105 13323 35139
rect 13265 35099 13323 35105
rect 13280 35068 13308 35099
rect 13096 35040 13308 35068
rect 9674 34960 9680 35012
rect 9732 35000 9738 35012
rect 11882 35000 11888 35012
rect 9732 34972 11888 35000
rect 9732 34960 9738 34972
rect 11882 34960 11888 34972
rect 11940 35000 11946 35012
rect 13538 35000 13544 35012
rect 11940 34972 13544 35000
rect 11940 34960 11946 34972
rect 13538 34960 13544 34972
rect 13596 34960 13602 35012
rect 8294 34932 8300 34944
rect 7208 34904 8300 34932
rect 3844 34892 3850 34904
rect 8294 34892 8300 34904
rect 8352 34892 8358 34944
rect 9858 34932 9864 34944
rect 9819 34904 9864 34932
rect 9858 34892 9864 34904
rect 9916 34892 9922 34944
rect 9950 34892 9956 34944
rect 10008 34932 10014 34944
rect 13648 34932 13676 35176
rect 14093 35173 14105 35176
rect 14139 35204 14151 35207
rect 15562 35204 15568 35216
rect 14139 35176 15568 35204
rect 14139 35173 14151 35176
rect 14093 35167 14151 35173
rect 15562 35164 15568 35176
rect 15620 35164 15626 35216
rect 13814 35136 13820 35148
rect 13775 35108 13820 35136
rect 13814 35096 13820 35108
rect 13872 35096 13878 35148
rect 14182 35136 14188 35148
rect 14143 35108 14188 35136
rect 14182 35096 14188 35108
rect 14240 35096 14246 35148
rect 16117 35139 16175 35145
rect 16117 35105 16129 35139
rect 16163 35136 16175 35139
rect 17126 35136 17132 35148
rect 16163 35108 17132 35136
rect 16163 35105 16175 35108
rect 16117 35099 16175 35105
rect 17126 35096 17132 35108
rect 17184 35096 17190 35148
rect 17236 35145 17264 35244
rect 18874 35232 18880 35244
rect 18932 35232 18938 35284
rect 19150 35232 19156 35284
rect 19208 35272 19214 35284
rect 20349 35275 20407 35281
rect 20349 35272 20361 35275
rect 19208 35244 20361 35272
rect 19208 35232 19214 35244
rect 20349 35241 20361 35244
rect 20395 35241 20407 35275
rect 21542 35272 21548 35284
rect 20349 35235 20407 35241
rect 20548 35244 21548 35272
rect 17221 35139 17279 35145
rect 17221 35105 17233 35139
rect 17267 35105 17279 35139
rect 17221 35099 17279 35105
rect 17586 35096 17592 35148
rect 17644 35136 17650 35148
rect 20548 35145 20576 35244
rect 21542 35232 21548 35244
rect 21600 35272 21606 35284
rect 22097 35275 22155 35281
rect 22097 35272 22109 35275
rect 21600 35244 22109 35272
rect 21600 35232 21606 35244
rect 22097 35241 22109 35244
rect 22143 35241 22155 35275
rect 25501 35275 25559 35281
rect 25501 35272 25513 35275
rect 22097 35235 22155 35241
rect 22296 35244 25513 35272
rect 19429 35139 19487 35145
rect 19429 35136 19441 35139
rect 17644 35108 19441 35136
rect 17644 35096 17650 35108
rect 19429 35105 19441 35108
rect 19475 35105 19487 35139
rect 19429 35099 19487 35105
rect 20533 35139 20591 35145
rect 20533 35105 20545 35139
rect 20579 35105 20591 35139
rect 20990 35136 20996 35148
rect 20951 35108 20996 35136
rect 20533 35099 20591 35105
rect 20990 35096 20996 35108
rect 21048 35096 21054 35148
rect 22296 35145 22324 35244
rect 25501 35241 25513 35244
rect 25547 35272 25559 35275
rect 28629 35275 28687 35281
rect 25547 35244 26648 35272
rect 25547 35241 25559 35244
rect 25501 35235 25559 35241
rect 22281 35139 22339 35145
rect 22281 35105 22293 35139
rect 22327 35105 22339 35139
rect 22646 35136 22652 35148
rect 22607 35108 22652 35136
rect 22281 35099 22339 35105
rect 22646 35096 22652 35108
rect 22704 35096 22710 35148
rect 24029 35139 24087 35145
rect 24029 35105 24041 35139
rect 24075 35136 24087 35139
rect 24581 35139 24639 35145
rect 24581 35136 24593 35139
rect 24075 35108 24593 35136
rect 24075 35105 24087 35108
rect 24029 35099 24087 35105
rect 24581 35105 24593 35108
rect 24627 35105 24639 35139
rect 24581 35099 24639 35105
rect 24762 35096 24768 35148
rect 24820 35136 24826 35148
rect 25685 35139 25743 35145
rect 25685 35136 25697 35139
rect 24820 35108 25697 35136
rect 24820 35096 24826 35108
rect 25685 35105 25697 35108
rect 25731 35105 25743 35139
rect 25685 35099 25743 35105
rect 15289 35071 15347 35077
rect 15289 35037 15301 35071
rect 15335 35068 15347 35071
rect 15562 35068 15568 35080
rect 15335 35040 15568 35068
rect 15335 35037 15347 35040
rect 15289 35031 15347 35037
rect 15562 35028 15568 35040
rect 15620 35028 15626 35080
rect 15838 35068 15844 35080
rect 15799 35040 15844 35068
rect 15838 35028 15844 35040
rect 15896 35028 15902 35080
rect 16301 35071 16359 35077
rect 16301 35037 16313 35071
rect 16347 35068 16359 35071
rect 16482 35068 16488 35080
rect 16347 35040 16488 35068
rect 16347 35037 16359 35040
rect 16301 35031 16359 35037
rect 16482 35028 16488 35040
rect 16540 35028 16546 35080
rect 17497 35071 17555 35077
rect 17497 35037 17509 35071
rect 17543 35068 17555 35071
rect 19337 35071 19395 35077
rect 17543 35040 18552 35068
rect 17543 35037 17555 35040
rect 17497 35031 17555 35037
rect 18524 35000 18552 35040
rect 19337 35037 19349 35071
rect 19383 35068 19395 35071
rect 20806 35068 20812 35080
rect 19383 35040 20812 35068
rect 19383 35037 19395 35040
rect 19337 35031 19395 35037
rect 20806 35028 20812 35040
rect 20864 35068 20870 35080
rect 20901 35071 20959 35077
rect 20901 35068 20913 35071
rect 20864 35040 20913 35068
rect 20864 35028 20870 35040
rect 20901 35037 20913 35040
rect 20947 35037 20959 35071
rect 22370 35068 22376 35080
rect 22331 35040 22376 35068
rect 20901 35031 20959 35037
rect 22370 35028 22376 35040
rect 22428 35028 22434 35080
rect 23382 35028 23388 35080
rect 23440 35068 23446 35080
rect 24489 35071 24547 35077
rect 24489 35068 24501 35071
rect 23440 35040 24501 35068
rect 23440 35028 23446 35040
rect 24489 35037 24501 35040
rect 24535 35037 24547 35071
rect 26510 35068 26516 35080
rect 26471 35040 26516 35068
rect 24489 35031 24547 35037
rect 26510 35028 26516 35040
rect 26568 35028 26574 35080
rect 26620 35068 26648 35244
rect 28629 35241 28641 35275
rect 28675 35272 28687 35275
rect 29086 35272 29092 35284
rect 28675 35244 29092 35272
rect 28675 35241 28687 35244
rect 28629 35235 28687 35241
rect 29086 35232 29092 35244
rect 29144 35272 29150 35284
rect 33778 35272 33784 35284
rect 29144 35244 30972 35272
rect 33739 35244 33784 35272
rect 29144 35232 29150 35244
rect 30650 35204 30656 35216
rect 28736 35176 30656 35204
rect 26789 35139 26847 35145
rect 26789 35105 26801 35139
rect 26835 35136 26847 35139
rect 28736 35136 28764 35176
rect 30650 35164 30656 35176
rect 30708 35164 30714 35216
rect 26835 35108 28764 35136
rect 28813 35139 28871 35145
rect 26835 35105 26847 35108
rect 26789 35099 26847 35105
rect 28813 35105 28825 35139
rect 28859 35105 28871 35139
rect 29362 35136 29368 35148
rect 29323 35108 29368 35136
rect 28813 35099 28871 35105
rect 28828 35068 28856 35099
rect 29362 35096 29368 35108
rect 29420 35096 29426 35148
rect 29917 35139 29975 35145
rect 29917 35105 29929 35139
rect 29963 35136 29975 35139
rect 30098 35136 30104 35148
rect 29963 35108 30104 35136
rect 29963 35105 29975 35108
rect 29917 35099 29975 35105
rect 30098 35096 30104 35108
rect 30156 35096 30162 35148
rect 30193 35139 30251 35145
rect 30193 35105 30205 35139
rect 30239 35136 30251 35139
rect 30374 35136 30380 35148
rect 30239 35108 30380 35136
rect 30239 35105 30251 35108
rect 30193 35099 30251 35105
rect 30374 35096 30380 35108
rect 30432 35096 30438 35148
rect 30944 35145 30972 35244
rect 33778 35232 33784 35244
rect 33836 35232 33842 35284
rect 35894 35272 35900 35284
rect 35360 35244 35900 35272
rect 31018 35164 31024 35216
rect 31076 35204 31082 35216
rect 31076 35176 31156 35204
rect 31076 35164 31082 35176
rect 31128 35145 31156 35176
rect 30929 35139 30987 35145
rect 30929 35105 30941 35139
rect 30975 35105 30987 35139
rect 30929 35099 30987 35105
rect 31113 35139 31171 35145
rect 31113 35105 31125 35139
rect 31159 35136 31171 35139
rect 32493 35139 32551 35145
rect 31159 35108 32444 35136
rect 31159 35105 31171 35108
rect 31113 35099 31171 35105
rect 31018 35068 31024 35080
rect 26620 35040 28856 35068
rect 30979 35040 31024 35068
rect 31018 35028 31024 35040
rect 31076 35028 31082 35080
rect 31573 35071 31631 35077
rect 31573 35037 31585 35071
rect 31619 35068 31631 35071
rect 31846 35068 31852 35080
rect 31619 35040 31852 35068
rect 31619 35037 31631 35040
rect 31573 35031 31631 35037
rect 31846 35028 31852 35040
rect 31904 35028 31910 35080
rect 32214 35068 32220 35080
rect 32175 35040 32220 35068
rect 32214 35028 32220 35040
rect 32272 35028 32278 35080
rect 32416 35068 32444 35108
rect 32493 35105 32505 35139
rect 32539 35136 32551 35139
rect 33410 35136 33416 35148
rect 32539 35108 33416 35136
rect 32539 35105 32551 35108
rect 32493 35099 32551 35105
rect 33410 35096 33416 35108
rect 33468 35096 33474 35148
rect 33796 35136 33824 35232
rect 34146 35164 34152 35216
rect 34204 35204 34210 35216
rect 34204 35176 35204 35204
rect 34204 35164 34210 35176
rect 35176 35145 35204 35176
rect 35360 35145 35388 35244
rect 35894 35232 35900 35244
rect 35952 35232 35958 35284
rect 35526 35164 35532 35216
rect 35584 35204 35590 35216
rect 35802 35204 35808 35216
rect 35584 35176 35808 35204
rect 35584 35164 35590 35176
rect 35802 35164 35808 35176
rect 35860 35204 35866 35216
rect 35860 35176 36492 35204
rect 35860 35164 35866 35176
rect 34333 35139 34391 35145
rect 34333 35136 34345 35139
rect 33796 35108 34345 35136
rect 34333 35105 34345 35108
rect 34379 35105 34391 35139
rect 34333 35099 34391 35105
rect 35161 35139 35219 35145
rect 35161 35105 35173 35139
rect 35207 35105 35219 35139
rect 35161 35099 35219 35105
rect 35345 35139 35403 35145
rect 35345 35105 35357 35139
rect 35391 35105 35403 35139
rect 36078 35136 36084 35148
rect 36039 35108 36084 35136
rect 35345 35099 35403 35105
rect 35176 35068 35204 35099
rect 36078 35096 36084 35108
rect 36136 35096 36142 35148
rect 36464 35145 36492 35176
rect 36449 35139 36507 35145
rect 36449 35105 36461 35139
rect 36495 35105 36507 35139
rect 36449 35099 36507 35105
rect 36265 35071 36323 35077
rect 36265 35068 36277 35071
rect 32416 35040 34928 35068
rect 35176 35040 36277 35068
rect 29273 35003 29331 35009
rect 29273 35000 29285 35003
rect 18524 34972 19656 35000
rect 10008 34904 13676 34932
rect 18785 34935 18843 34941
rect 10008 34892 10014 34904
rect 18785 34901 18797 34935
rect 18831 34932 18843 34935
rect 19058 34932 19064 34944
rect 18831 34904 19064 34932
rect 18831 34901 18843 34904
rect 18785 34895 18843 34901
rect 19058 34892 19064 34904
rect 19116 34892 19122 34944
rect 19628 34941 19656 34972
rect 27448 34972 29285 35000
rect 19613 34935 19671 34941
rect 19613 34901 19625 34935
rect 19659 34901 19671 34935
rect 21174 34932 21180 34944
rect 21135 34904 21180 34932
rect 19613 34895 19671 34901
rect 21174 34892 21180 34904
rect 21232 34892 21238 34944
rect 24394 34892 24400 34944
rect 24452 34932 24458 34944
rect 24765 34935 24823 34941
rect 24765 34932 24777 34935
rect 24452 34904 24777 34932
rect 24452 34892 24458 34904
rect 24765 34901 24777 34904
rect 24811 34901 24823 34935
rect 24765 34895 24823 34901
rect 25958 34892 25964 34944
rect 26016 34932 26022 34944
rect 27448 34932 27476 34972
rect 29273 34969 29285 34972
rect 29319 34969 29331 35003
rect 30742 35000 30748 35012
rect 30655 34972 30748 35000
rect 29273 34963 29331 34969
rect 30742 34960 30748 34972
rect 30800 35000 30806 35012
rect 32232 35000 32260 35028
rect 30800 34972 32260 35000
rect 34900 35000 34928 35040
rect 36265 35037 36277 35040
rect 36311 35068 36323 35071
rect 36906 35068 36912 35080
rect 36311 35040 36912 35068
rect 36311 35037 36323 35040
rect 36265 35031 36323 35037
rect 36906 35028 36912 35040
rect 36964 35028 36970 35080
rect 35250 35000 35256 35012
rect 34900 34972 35256 35000
rect 30800 34960 30806 34972
rect 35250 34960 35256 34972
rect 35308 34960 35314 35012
rect 26016 34904 27476 34932
rect 26016 34892 26022 34904
rect 27522 34892 27528 34944
rect 27580 34932 27586 34944
rect 27893 34935 27951 34941
rect 27893 34932 27905 34935
rect 27580 34904 27905 34932
rect 27580 34892 27586 34904
rect 27893 34901 27905 34904
rect 27939 34901 27951 34935
rect 27893 34895 27951 34901
rect 35434 34892 35440 34944
rect 35492 34932 35498 34944
rect 35492 34904 35537 34932
rect 35492 34892 35498 34904
rect 1104 34842 38824 34864
rect 1104 34790 4246 34842
rect 4298 34790 4310 34842
rect 4362 34790 4374 34842
rect 4426 34790 4438 34842
rect 4490 34790 34966 34842
rect 35018 34790 35030 34842
rect 35082 34790 35094 34842
rect 35146 34790 35158 34842
rect 35210 34790 38824 34842
rect 1104 34768 38824 34790
rect 2222 34688 2228 34740
rect 2280 34728 2286 34740
rect 6914 34728 6920 34740
rect 2280 34700 6920 34728
rect 2280 34688 2286 34700
rect 6914 34688 6920 34700
rect 6972 34688 6978 34740
rect 15197 34731 15255 34737
rect 15197 34728 15209 34731
rect 11900 34700 15209 34728
rect 5534 34660 5540 34672
rect 2056 34632 4752 34660
rect 1397 34595 1455 34601
rect 1397 34561 1409 34595
rect 1443 34592 1455 34595
rect 2056 34592 2084 34632
rect 1443 34564 2084 34592
rect 2133 34595 2191 34601
rect 1443 34561 1455 34564
rect 1397 34555 1455 34561
rect 2133 34561 2145 34595
rect 2179 34592 2191 34595
rect 4154 34592 4160 34604
rect 2179 34564 4160 34592
rect 2179 34561 2191 34564
rect 2133 34555 2191 34561
rect 4154 34552 4160 34564
rect 4212 34552 4218 34604
rect 4724 34601 4752 34632
rect 5460 34632 5540 34660
rect 4709 34595 4767 34601
rect 4709 34561 4721 34595
rect 4755 34561 4767 34595
rect 4709 34555 4767 34561
rect 1673 34527 1731 34533
rect 1673 34493 1685 34527
rect 1719 34524 1731 34527
rect 2222 34524 2228 34536
rect 1719 34496 2228 34524
rect 1719 34493 1731 34496
rect 1673 34487 1731 34493
rect 2222 34484 2228 34496
rect 2280 34484 2286 34536
rect 2682 34524 2688 34536
rect 2643 34496 2688 34524
rect 2682 34484 2688 34496
rect 2740 34484 2746 34536
rect 3234 34524 3240 34536
rect 3195 34496 3240 34524
rect 3234 34484 3240 34496
rect 3292 34484 3298 34536
rect 3602 34524 3608 34536
rect 3563 34496 3608 34524
rect 3602 34484 3608 34496
rect 3660 34484 3666 34536
rect 3786 34524 3792 34536
rect 3747 34496 3792 34524
rect 3786 34484 3792 34496
rect 3844 34484 3850 34536
rect 4065 34527 4123 34533
rect 4065 34493 4077 34527
rect 4111 34524 4123 34527
rect 4614 34524 4620 34536
rect 4111 34496 4620 34524
rect 4111 34493 4123 34496
rect 4065 34487 4123 34493
rect 4614 34484 4620 34496
rect 4672 34484 4678 34536
rect 5460 34533 5488 34632
rect 5534 34620 5540 34632
rect 5592 34620 5598 34672
rect 6641 34663 6699 34669
rect 6641 34629 6653 34663
rect 6687 34660 6699 34663
rect 8570 34660 8576 34672
rect 6687 34632 8576 34660
rect 6687 34629 6699 34632
rect 6641 34623 6699 34629
rect 8570 34620 8576 34632
rect 8628 34620 8634 34672
rect 10778 34660 10784 34672
rect 9416 34632 10784 34660
rect 6822 34592 6828 34604
rect 5828 34564 6828 34592
rect 5261 34527 5319 34533
rect 5261 34493 5273 34527
rect 5307 34524 5319 34527
rect 5445 34527 5503 34533
rect 5307 34496 5396 34524
rect 5307 34493 5319 34496
rect 5261 34487 5319 34493
rect 1578 34456 1584 34468
rect 1539 34428 1584 34456
rect 1578 34416 1584 34428
rect 1636 34416 1642 34468
rect 5368 34456 5396 34496
rect 5445 34493 5457 34527
rect 5491 34493 5503 34527
rect 5626 34524 5632 34536
rect 5587 34496 5632 34524
rect 5445 34487 5503 34493
rect 5626 34484 5632 34496
rect 5684 34484 5690 34536
rect 5718 34484 5724 34536
rect 5776 34524 5782 34536
rect 5828 34533 5856 34564
rect 6822 34552 6828 34564
rect 6880 34592 6886 34604
rect 7926 34592 7932 34604
rect 6880 34564 7932 34592
rect 6880 34552 6886 34564
rect 7926 34552 7932 34564
rect 7984 34552 7990 34604
rect 9416 34601 9444 34632
rect 10778 34620 10784 34632
rect 10836 34620 10842 34672
rect 9401 34595 9459 34601
rect 9401 34561 9413 34595
rect 9447 34561 9459 34595
rect 10318 34592 10324 34604
rect 10279 34564 10324 34592
rect 9401 34555 9459 34561
rect 10318 34552 10324 34564
rect 10376 34552 10382 34604
rect 11514 34592 11520 34604
rect 10704 34564 11520 34592
rect 5813 34527 5871 34533
rect 5813 34524 5825 34527
rect 5776 34496 5825 34524
rect 5776 34484 5782 34496
rect 5813 34493 5825 34496
rect 5859 34493 5871 34527
rect 5813 34487 5871 34493
rect 6089 34527 6147 34533
rect 6089 34493 6101 34527
rect 6135 34524 6147 34527
rect 6641 34527 6699 34533
rect 6641 34524 6653 34527
rect 6135 34496 6653 34524
rect 6135 34493 6147 34496
rect 6089 34487 6147 34493
rect 6641 34493 6653 34496
rect 6687 34493 6699 34527
rect 7282 34524 7288 34536
rect 7243 34496 7288 34524
rect 6641 34487 6699 34493
rect 7282 34484 7288 34496
rect 7340 34484 7346 34536
rect 7653 34527 7711 34533
rect 7653 34493 7665 34527
rect 7699 34493 7711 34527
rect 7653 34487 7711 34493
rect 9769 34527 9827 34533
rect 9769 34493 9781 34527
rect 9815 34524 9827 34527
rect 9858 34524 9864 34536
rect 9815 34496 9864 34524
rect 9815 34493 9827 34496
rect 9769 34487 9827 34493
rect 5994 34456 6000 34468
rect 5368 34428 6000 34456
rect 5994 34416 6000 34428
rect 6052 34416 6058 34468
rect 7006 34416 7012 34468
rect 7064 34456 7070 34468
rect 7668 34456 7696 34487
rect 9858 34484 9864 34496
rect 9916 34484 9922 34536
rect 10137 34527 10195 34533
rect 10137 34493 10149 34527
rect 10183 34524 10195 34527
rect 10704 34524 10732 34564
rect 11514 34552 11520 34564
rect 11572 34592 11578 34604
rect 11701 34595 11759 34601
rect 11701 34592 11713 34595
rect 11572 34564 11713 34592
rect 11572 34552 11578 34564
rect 11701 34561 11713 34564
rect 11747 34592 11759 34595
rect 11900 34592 11928 34700
rect 15197 34697 15209 34700
rect 15243 34697 15255 34731
rect 15197 34691 15255 34697
rect 17405 34731 17463 34737
rect 17405 34697 17417 34731
rect 17451 34728 17463 34731
rect 17586 34728 17592 34740
rect 17451 34700 17592 34728
rect 17451 34697 17463 34700
rect 17405 34691 17463 34697
rect 17586 34688 17592 34700
rect 17644 34688 17650 34740
rect 19352 34700 21496 34728
rect 12621 34663 12679 34669
rect 12621 34660 12633 34663
rect 11747 34564 11928 34592
rect 11992 34632 12633 34660
rect 11747 34561 11759 34564
rect 11701 34555 11759 34561
rect 10183 34496 10732 34524
rect 10183 34493 10195 34496
rect 10137 34487 10195 34493
rect 10778 34484 10784 34536
rect 10836 34524 10842 34536
rect 11609 34527 11667 34533
rect 10836 34496 10881 34524
rect 10836 34484 10842 34496
rect 11609 34493 11621 34527
rect 11655 34524 11667 34527
rect 11882 34524 11888 34536
rect 11655 34496 11888 34524
rect 11655 34493 11667 34496
rect 11609 34487 11667 34493
rect 11882 34484 11888 34496
rect 11940 34484 11946 34536
rect 7064 34428 7696 34456
rect 7064 34416 7070 34428
rect 11146 34416 11152 34468
rect 11204 34456 11210 34468
rect 11992 34456 12020 34632
rect 12621 34629 12633 34632
rect 12667 34629 12679 34663
rect 12621 34623 12679 34629
rect 16850 34620 16856 34672
rect 16908 34660 16914 34672
rect 18141 34663 18199 34669
rect 18141 34660 18153 34663
rect 16908 34632 18153 34660
rect 16908 34620 16914 34632
rect 18141 34629 18153 34632
rect 18187 34629 18199 34663
rect 18141 34623 18199 34629
rect 13173 34595 13231 34601
rect 13173 34561 13185 34595
rect 13219 34592 13231 34595
rect 14274 34592 14280 34604
rect 13219 34564 14280 34592
rect 13219 34561 13231 34564
rect 13173 34555 13231 34561
rect 14274 34552 14280 34564
rect 14332 34552 14338 34604
rect 15010 34552 15016 34604
rect 15068 34592 15074 34604
rect 15841 34595 15899 34601
rect 15841 34592 15853 34595
rect 15068 34564 15853 34592
rect 15068 34552 15074 34564
rect 15841 34561 15853 34564
rect 15887 34561 15899 34595
rect 16114 34592 16120 34604
rect 16075 34564 16120 34592
rect 15841 34555 15899 34561
rect 16114 34552 16120 34564
rect 16172 34552 16178 34604
rect 17678 34552 17684 34604
rect 17736 34592 17742 34604
rect 19242 34592 19248 34604
rect 17736 34564 19248 34592
rect 17736 34552 17742 34564
rect 19242 34552 19248 34564
rect 19300 34552 19306 34604
rect 19352 34601 19380 34700
rect 19337 34595 19395 34601
rect 19337 34561 19349 34595
rect 19383 34561 19395 34595
rect 19337 34555 19395 34561
rect 19613 34595 19671 34601
rect 19613 34561 19625 34595
rect 19659 34592 19671 34595
rect 21174 34592 21180 34604
rect 19659 34564 21180 34592
rect 19659 34561 19671 34564
rect 19613 34555 19671 34561
rect 12437 34527 12495 34533
rect 12437 34493 12449 34527
rect 12483 34524 12495 34527
rect 12526 34524 12532 34536
rect 12483 34496 12532 34524
rect 12483 34493 12495 34496
rect 12437 34487 12495 34493
rect 12526 34484 12532 34496
rect 12584 34484 12590 34536
rect 13354 34484 13360 34536
rect 13412 34524 13418 34536
rect 13633 34527 13691 34533
rect 13633 34524 13645 34527
rect 13412 34496 13645 34524
rect 13412 34484 13418 34496
rect 13633 34493 13645 34496
rect 13679 34493 13691 34527
rect 13814 34524 13820 34536
rect 13775 34496 13820 34524
rect 13633 34487 13691 34493
rect 13814 34484 13820 34496
rect 13872 34484 13878 34536
rect 13998 34524 14004 34536
rect 13959 34496 14004 34524
rect 13998 34484 14004 34496
rect 14056 34484 14062 34536
rect 14182 34524 14188 34536
rect 14143 34496 14188 34524
rect 14182 34484 14188 34496
rect 14240 34484 14246 34536
rect 14458 34524 14464 34536
rect 14419 34496 14464 34524
rect 14458 34484 14464 34496
rect 14516 34484 14522 34536
rect 15105 34527 15163 34533
rect 15105 34493 15117 34527
rect 15151 34493 15163 34527
rect 18046 34524 18052 34536
rect 18007 34496 18052 34524
rect 15105 34487 15163 34493
rect 11204 34428 12020 34456
rect 14200 34456 14228 34484
rect 15120 34456 15148 34487
rect 18046 34484 18052 34496
rect 18104 34484 18110 34536
rect 18138 34484 18144 34536
rect 18196 34524 18202 34536
rect 18601 34527 18659 34533
rect 18601 34524 18613 34527
rect 18196 34496 18613 34524
rect 18196 34484 18202 34496
rect 18601 34493 18613 34496
rect 18647 34493 18659 34527
rect 18601 34487 18659 34493
rect 14200 34428 15148 34456
rect 11204 34416 11210 34428
rect 18690 34416 18696 34468
rect 18748 34456 18754 34468
rect 19352 34456 19380 34555
rect 21174 34552 21180 34564
rect 21232 34552 21238 34604
rect 21468 34601 21496 34700
rect 32306 34688 32312 34740
rect 32364 34728 32370 34740
rect 32769 34731 32827 34737
rect 32769 34728 32781 34731
rect 32364 34700 32781 34728
rect 32364 34688 32370 34700
rect 32769 34697 32781 34700
rect 32815 34697 32827 34731
rect 32769 34691 32827 34697
rect 33134 34688 33140 34740
rect 33192 34728 33198 34740
rect 36354 34728 36360 34740
rect 33192 34700 36360 34728
rect 33192 34688 33198 34700
rect 33704 34669 33732 34700
rect 36354 34688 36360 34700
rect 36412 34688 36418 34740
rect 33689 34663 33747 34669
rect 33689 34629 33701 34663
rect 33735 34629 33747 34663
rect 35802 34660 35808 34672
rect 33689 34623 33747 34629
rect 33888 34632 35808 34660
rect 21453 34595 21511 34601
rect 21453 34561 21465 34595
rect 21499 34592 21511 34595
rect 22370 34592 22376 34604
rect 21499 34564 22376 34592
rect 21499 34561 21511 34564
rect 21453 34555 21511 34561
rect 22370 34552 22376 34564
rect 22428 34552 22434 34604
rect 24394 34592 24400 34604
rect 24355 34564 24400 34592
rect 24394 34552 24400 34564
rect 24452 34552 24458 34604
rect 25498 34592 25504 34604
rect 25459 34564 25504 34592
rect 25498 34552 25504 34564
rect 25556 34552 25562 34604
rect 27341 34595 27399 34601
rect 27341 34561 27353 34595
rect 27387 34592 27399 34595
rect 27522 34592 27528 34604
rect 27387 34564 27528 34592
rect 27387 34561 27399 34564
rect 27341 34555 27399 34561
rect 27522 34552 27528 34564
rect 27580 34552 27586 34604
rect 20993 34527 21051 34533
rect 20993 34493 21005 34527
rect 21039 34524 21051 34527
rect 21358 34524 21364 34536
rect 21039 34496 21364 34524
rect 21039 34493 21051 34496
rect 20993 34487 21051 34493
rect 21358 34484 21364 34496
rect 21416 34484 21422 34536
rect 21726 34524 21732 34536
rect 21687 34496 21732 34524
rect 21726 34484 21732 34496
rect 21784 34484 21790 34536
rect 23109 34527 23167 34533
rect 23109 34493 23121 34527
rect 23155 34524 23167 34527
rect 23842 34524 23848 34536
rect 23155 34496 23848 34524
rect 23155 34493 23167 34496
rect 23109 34487 23167 34493
rect 23842 34484 23848 34496
rect 23900 34484 23906 34536
rect 24121 34527 24179 34533
rect 24121 34493 24133 34527
rect 24167 34524 24179 34527
rect 24210 34524 24216 34536
rect 24167 34496 24216 34524
rect 24167 34493 24179 34496
rect 24121 34487 24179 34493
rect 24210 34484 24216 34496
rect 24268 34484 24274 34536
rect 26510 34484 26516 34536
rect 26568 34524 26574 34536
rect 27065 34527 27123 34533
rect 27065 34524 27077 34527
rect 26568 34496 27077 34524
rect 26568 34484 26574 34496
rect 27065 34493 27077 34496
rect 27111 34524 27123 34527
rect 28902 34524 28908 34536
rect 27111 34496 28908 34524
rect 27111 34493 27123 34496
rect 27065 34487 27123 34493
rect 28902 34484 28908 34496
rect 28960 34524 28966 34536
rect 29273 34527 29331 34533
rect 29273 34524 29285 34527
rect 28960 34496 29285 34524
rect 28960 34484 28966 34496
rect 29273 34493 29285 34496
rect 29319 34493 29331 34527
rect 29546 34524 29552 34536
rect 29507 34496 29552 34524
rect 29273 34487 29331 34493
rect 29546 34484 29552 34496
rect 29604 34484 29610 34536
rect 31386 34524 31392 34536
rect 31347 34496 31392 34524
rect 31386 34484 31392 34496
rect 31444 34484 31450 34536
rect 31662 34524 31668 34536
rect 31623 34496 31668 34524
rect 31662 34484 31668 34496
rect 31720 34484 31726 34536
rect 33502 34484 33508 34536
rect 33560 34524 33566 34536
rect 33888 34533 33916 34632
rect 35802 34620 35808 34632
rect 35860 34620 35866 34672
rect 34333 34595 34391 34601
rect 34333 34561 34345 34595
rect 34379 34592 34391 34595
rect 34514 34592 34520 34604
rect 34379 34564 34520 34592
rect 34379 34561 34391 34564
rect 34333 34555 34391 34561
rect 34514 34552 34520 34564
rect 34572 34552 34578 34604
rect 37274 34592 37280 34604
rect 37235 34564 37280 34592
rect 37274 34552 37280 34564
rect 37332 34552 37338 34604
rect 33597 34527 33655 34533
rect 33597 34524 33609 34527
rect 33560 34496 33609 34524
rect 33560 34484 33566 34496
rect 33597 34493 33609 34496
rect 33643 34524 33655 34527
rect 33873 34527 33931 34533
rect 33643 34496 33824 34524
rect 33643 34493 33655 34496
rect 33597 34487 33655 34493
rect 18748 34428 19380 34456
rect 33796 34456 33824 34496
rect 33873 34493 33885 34527
rect 33919 34493 33931 34527
rect 35434 34524 35440 34536
rect 33873 34487 33931 34493
rect 33980 34496 35440 34524
rect 33980 34456 34008 34496
rect 35434 34484 35440 34496
rect 35492 34524 35498 34536
rect 35621 34527 35679 34533
rect 35621 34524 35633 34527
rect 35492 34496 35633 34524
rect 35492 34484 35498 34496
rect 35621 34493 35633 34496
rect 35667 34493 35679 34527
rect 35621 34487 35679 34493
rect 36541 34527 36599 34533
rect 36541 34493 36553 34527
rect 36587 34524 36599 34527
rect 37182 34524 37188 34536
rect 36587 34496 37188 34524
rect 36587 34493 36599 34496
rect 36541 34487 36599 34493
rect 37182 34484 37188 34496
rect 37240 34484 37246 34536
rect 33796 34428 34008 34456
rect 18748 34416 18754 34428
rect 7193 34391 7251 34397
rect 7193 34357 7205 34391
rect 7239 34388 7251 34391
rect 7650 34388 7656 34400
rect 7239 34360 7656 34388
rect 7239 34357 7251 34360
rect 7193 34351 7251 34357
rect 7650 34348 7656 34360
rect 7708 34348 7714 34400
rect 11054 34388 11060 34400
rect 11015 34360 11060 34388
rect 11054 34348 11060 34360
rect 11112 34348 11118 34400
rect 28442 34388 28448 34400
rect 28403 34360 28448 34388
rect 28442 34348 28448 34360
rect 28500 34348 28506 34400
rect 30650 34388 30656 34400
rect 30611 34360 30656 34388
rect 30650 34348 30656 34360
rect 30708 34348 30714 34400
rect 1104 34298 38824 34320
rect 1104 34246 19606 34298
rect 19658 34246 19670 34298
rect 19722 34246 19734 34298
rect 19786 34246 19798 34298
rect 19850 34246 38824 34298
rect 1104 34224 38824 34246
rect 2682 34144 2688 34196
rect 2740 34184 2746 34196
rect 2777 34187 2835 34193
rect 2777 34184 2789 34187
rect 2740 34156 2789 34184
rect 2740 34144 2746 34156
rect 2777 34153 2789 34156
rect 2823 34153 2835 34187
rect 5994 34184 6000 34196
rect 5955 34156 6000 34184
rect 2777 34147 2835 34153
rect 5994 34144 6000 34156
rect 6052 34184 6058 34196
rect 6052 34156 6776 34184
rect 6052 34144 6058 34156
rect 4154 34008 4160 34060
rect 4212 34048 4218 34060
rect 6748 34057 6776 34156
rect 8570 34144 8576 34196
rect 8628 34184 8634 34196
rect 8849 34187 8907 34193
rect 8849 34184 8861 34187
rect 8628 34156 8861 34184
rect 8628 34144 8634 34156
rect 8849 34153 8861 34156
rect 8895 34184 8907 34187
rect 9861 34187 9919 34193
rect 9861 34184 9873 34187
rect 8895 34156 9873 34184
rect 8895 34153 8907 34156
rect 8849 34147 8907 34153
rect 9861 34153 9873 34156
rect 9907 34153 9919 34187
rect 9861 34147 9919 34153
rect 11149 34187 11207 34193
rect 11149 34153 11161 34187
rect 11195 34184 11207 34187
rect 11238 34184 11244 34196
rect 11195 34156 11244 34184
rect 11195 34153 11207 34156
rect 11149 34147 11207 34153
rect 11238 34144 11244 34156
rect 11296 34144 11302 34196
rect 12618 34144 12624 34196
rect 12676 34184 12682 34196
rect 14369 34187 14427 34193
rect 14369 34184 14381 34187
rect 12676 34156 14381 34184
rect 12676 34144 12682 34156
rect 14369 34153 14381 34156
rect 14415 34184 14427 34187
rect 14458 34184 14464 34196
rect 14415 34156 14464 34184
rect 14415 34153 14427 34156
rect 14369 34147 14427 34153
rect 14458 34144 14464 34156
rect 14516 34144 14522 34196
rect 29546 34184 29552 34196
rect 29507 34156 29552 34184
rect 29546 34144 29552 34156
rect 29604 34144 29610 34196
rect 30300 34156 32168 34184
rect 7006 34076 7012 34128
rect 7064 34116 7070 34128
rect 7064 34088 7512 34116
rect 7064 34076 7070 34088
rect 4893 34051 4951 34057
rect 4893 34048 4905 34051
rect 4212 34020 4905 34048
rect 4212 34008 4218 34020
rect 4893 34017 4905 34020
rect 4939 34017 4951 34051
rect 4893 34011 4951 34017
rect 6733 34051 6791 34057
rect 6733 34017 6745 34051
rect 6779 34017 6791 34051
rect 7282 34048 7288 34060
rect 7243 34020 7288 34048
rect 6733 34011 6791 34017
rect 7282 34008 7288 34020
rect 7340 34008 7346 34060
rect 7484 34057 7512 34088
rect 9766 34076 9772 34128
rect 9824 34116 9830 34128
rect 9953 34119 10011 34125
rect 9953 34116 9965 34119
rect 9824 34088 9965 34116
rect 9824 34076 9830 34088
rect 9953 34085 9965 34088
rect 9999 34085 10011 34119
rect 9953 34079 10011 34085
rect 10045 34119 10103 34125
rect 10045 34085 10057 34119
rect 10091 34085 10103 34119
rect 10045 34079 10103 34085
rect 7469 34051 7527 34057
rect 7469 34017 7481 34051
rect 7515 34017 7527 34051
rect 7469 34011 7527 34017
rect 7926 34008 7932 34060
rect 7984 34048 7990 34060
rect 8021 34051 8079 34057
rect 8021 34048 8033 34051
rect 7984 34020 8033 34048
rect 7984 34008 7990 34020
rect 8021 34017 8033 34020
rect 8067 34017 8079 34051
rect 8021 34011 8079 34017
rect 8386 34008 8392 34060
rect 8444 34048 8450 34060
rect 8665 34051 8723 34057
rect 8665 34048 8677 34051
rect 8444 34020 8677 34048
rect 8444 34008 8450 34020
rect 8665 34017 8677 34020
rect 8711 34017 8723 34051
rect 8665 34011 8723 34017
rect 8754 34008 8760 34060
rect 8812 34048 8818 34060
rect 10060 34048 10088 34079
rect 10134 34076 10140 34128
rect 10192 34116 10198 34128
rect 10870 34116 10876 34128
rect 10192 34088 10876 34116
rect 10192 34076 10198 34088
rect 10870 34076 10876 34088
rect 10928 34116 10934 34128
rect 20349 34119 20407 34125
rect 10928 34088 12112 34116
rect 10928 34076 10934 34088
rect 11054 34048 11060 34060
rect 8812 34020 10088 34048
rect 11015 34020 11060 34048
rect 8812 34008 8818 34020
rect 11054 34008 11060 34020
rect 11112 34008 11118 34060
rect 11514 34048 11520 34060
rect 11475 34020 11520 34048
rect 11514 34008 11520 34020
rect 11572 34008 11578 34060
rect 11790 34048 11796 34060
rect 11751 34020 11796 34048
rect 11790 34008 11796 34020
rect 11848 34008 11854 34060
rect 12084 34057 12112 34088
rect 20349 34085 20361 34119
rect 20395 34116 20407 34119
rect 20990 34116 20996 34128
rect 20395 34088 20996 34116
rect 20395 34085 20407 34088
rect 20349 34079 20407 34085
rect 20990 34076 20996 34088
rect 21048 34076 21054 34128
rect 21726 34116 21732 34128
rect 21687 34088 21732 34116
rect 21726 34076 21732 34088
rect 21784 34076 21790 34128
rect 12069 34051 12127 34057
rect 12069 34017 12081 34051
rect 12115 34017 12127 34051
rect 13354 34048 13360 34060
rect 12069 34011 12127 34017
rect 12820 34020 13360 34048
rect 1394 33980 1400 33992
rect 1355 33952 1400 33980
rect 1394 33940 1400 33952
rect 1452 33940 1458 33992
rect 1673 33983 1731 33989
rect 1673 33949 1685 33983
rect 1719 33980 1731 33983
rect 1854 33980 1860 33992
rect 1719 33952 1860 33980
rect 1719 33949 1731 33952
rect 1673 33943 1731 33949
rect 1854 33940 1860 33952
rect 1912 33940 1918 33992
rect 3970 33940 3976 33992
rect 4028 33980 4034 33992
rect 4617 33983 4675 33989
rect 4617 33980 4629 33983
rect 4028 33952 4629 33980
rect 4028 33940 4034 33952
rect 4617 33949 4629 33952
rect 4663 33980 4675 33983
rect 5074 33980 5080 33992
rect 4663 33952 5080 33980
rect 4663 33949 4675 33952
rect 4617 33943 4675 33949
rect 5074 33940 5080 33952
rect 5132 33940 5138 33992
rect 6914 33980 6920 33992
rect 6875 33952 6920 33980
rect 6914 33940 6920 33952
rect 6972 33940 6978 33992
rect 8294 33940 8300 33992
rect 8352 33980 8358 33992
rect 9677 33983 9735 33989
rect 9677 33980 9689 33983
rect 8352 33952 9689 33980
rect 8352 33940 8358 33952
rect 9677 33949 9689 33952
rect 9723 33949 9735 33983
rect 9677 33943 9735 33949
rect 10413 33983 10471 33989
rect 10413 33949 10425 33983
rect 10459 33980 10471 33983
rect 12820 33980 12848 34020
rect 13354 34008 13360 34020
rect 13412 34008 13418 34060
rect 15565 34051 15623 34057
rect 15565 34017 15577 34051
rect 15611 34048 15623 34051
rect 16850 34048 16856 34060
rect 15611 34020 16856 34048
rect 15611 34017 15623 34020
rect 15565 34011 15623 34017
rect 16850 34008 16856 34020
rect 16908 34008 16914 34060
rect 18690 34048 18696 34060
rect 18651 34020 18696 34048
rect 18690 34008 18696 34020
rect 18748 34008 18754 34060
rect 18966 34048 18972 34060
rect 18927 34020 18972 34048
rect 18966 34008 18972 34020
rect 19024 34008 19030 34060
rect 19242 34008 19248 34060
rect 19300 34048 19306 34060
rect 21269 34051 21327 34057
rect 21269 34048 21281 34051
rect 19300 34020 21281 34048
rect 19300 34008 19306 34020
rect 21269 34017 21281 34020
rect 21315 34017 21327 34051
rect 23382 34048 23388 34060
rect 21269 34011 21327 34017
rect 22112 34020 23388 34048
rect 10459 33952 12848 33980
rect 12989 33983 13047 33989
rect 10459 33949 10471 33952
rect 10413 33943 10471 33949
rect 12989 33949 13001 33983
rect 13035 33949 13047 33983
rect 13262 33980 13268 33992
rect 13223 33952 13268 33980
rect 12989 33943 13047 33949
rect 12434 33872 12440 33924
rect 12492 33912 12498 33924
rect 13004 33912 13032 33943
rect 13262 33940 13268 33952
rect 13320 33940 13326 33992
rect 15286 33940 15292 33992
rect 15344 33980 15350 33992
rect 16209 33983 16267 33989
rect 16209 33980 16221 33983
rect 15344 33952 16221 33980
rect 15344 33940 15350 33952
rect 16209 33949 16221 33952
rect 16255 33949 16267 33983
rect 16209 33943 16267 33949
rect 16390 33940 16396 33992
rect 16448 33980 16454 33992
rect 16485 33983 16543 33989
rect 16485 33980 16497 33983
rect 16448 33952 16497 33980
rect 16448 33940 16454 33952
rect 16485 33949 16497 33952
rect 16531 33949 16543 33983
rect 16485 33943 16543 33949
rect 21177 33983 21235 33989
rect 21177 33949 21189 33983
rect 21223 33980 21235 33983
rect 22112 33980 22140 34020
rect 23382 34008 23388 34020
rect 23440 34008 23446 34060
rect 23845 34051 23903 34057
rect 23845 34017 23857 34051
rect 23891 34048 23903 34051
rect 26605 34051 26663 34057
rect 26605 34048 26617 34051
rect 23891 34020 26617 34048
rect 23891 34017 23903 34020
rect 23845 34011 23903 34017
rect 26605 34017 26617 34020
rect 26651 34017 26663 34051
rect 28442 34048 28448 34060
rect 28403 34020 28448 34048
rect 26605 34011 26663 34017
rect 28442 34008 28448 34020
rect 28500 34008 28506 34060
rect 29270 34008 29276 34060
rect 29328 34048 29334 34060
rect 30300 34057 30328 34156
rect 31573 34119 31631 34125
rect 31573 34085 31585 34119
rect 31619 34116 31631 34119
rect 31662 34116 31668 34128
rect 31619 34088 31668 34116
rect 31619 34085 31631 34088
rect 31573 34079 31631 34085
rect 31662 34076 31668 34088
rect 31720 34076 31726 34128
rect 30285 34051 30343 34057
rect 30285 34048 30297 34051
rect 29328 34020 30297 34048
rect 29328 34008 29334 34020
rect 30285 34017 30297 34020
rect 30331 34017 30343 34051
rect 30285 34011 30343 34017
rect 31113 34051 31171 34057
rect 31113 34017 31125 34051
rect 31159 34048 31171 34051
rect 31938 34048 31944 34060
rect 31159 34020 31944 34048
rect 31159 34017 31171 34020
rect 31113 34011 31171 34017
rect 31938 34008 31944 34020
rect 31996 34008 32002 34060
rect 32140 34057 32168 34156
rect 32214 34144 32220 34196
rect 32272 34184 32278 34196
rect 36446 34184 36452 34196
rect 32272 34156 36452 34184
rect 32272 34144 32278 34156
rect 36446 34144 36452 34156
rect 36504 34144 36510 34196
rect 32125 34051 32183 34057
rect 32125 34017 32137 34051
rect 32171 34017 32183 34051
rect 32125 34011 32183 34017
rect 32953 34051 33011 34057
rect 32953 34017 32965 34051
rect 32999 34048 33011 34051
rect 33042 34048 33048 34060
rect 32999 34020 33048 34048
rect 32999 34017 33011 34020
rect 32953 34011 33011 34017
rect 33042 34008 33048 34020
rect 33100 34008 33106 34060
rect 33413 34051 33471 34057
rect 33413 34017 33425 34051
rect 33459 34048 33471 34051
rect 34149 34051 34207 34057
rect 34149 34048 34161 34051
rect 33459 34020 34161 34048
rect 33459 34017 33471 34020
rect 33413 34011 33471 34017
rect 34149 34017 34161 34020
rect 34195 34017 34207 34051
rect 34149 34011 34207 34017
rect 35526 34008 35532 34060
rect 35584 34048 35590 34060
rect 36998 34048 37004 34060
rect 35584 34020 37004 34048
rect 35584 34008 35590 34020
rect 36998 34008 37004 34020
rect 37056 34008 37062 34060
rect 21223 33952 22140 33980
rect 22189 33983 22247 33989
rect 21223 33949 21235 33952
rect 21177 33943 21235 33949
rect 22189 33949 22201 33983
rect 22235 33949 22247 33983
rect 22189 33943 22247 33949
rect 22465 33983 22523 33989
rect 22465 33949 22477 33983
rect 22511 33980 22523 33983
rect 23934 33980 23940 33992
rect 22511 33952 23940 33980
rect 22511 33949 22523 33952
rect 22465 33943 22523 33949
rect 12492 33884 13032 33912
rect 12492 33872 12498 33884
rect 15657 33847 15715 33853
rect 15657 33813 15669 33847
rect 15703 33844 15715 33847
rect 17586 33844 17592 33856
rect 15703 33816 17592 33844
rect 15703 33813 15715 33816
rect 15657 33807 15715 33813
rect 17586 33804 17592 33816
rect 17644 33804 17650 33856
rect 17773 33847 17831 33853
rect 17773 33813 17785 33847
rect 17819 33844 17831 33847
rect 18414 33844 18420 33856
rect 17819 33816 18420 33844
rect 17819 33813 17831 33816
rect 17773 33807 17831 33813
rect 18414 33804 18420 33816
rect 18472 33804 18478 33856
rect 21634 33804 21640 33856
rect 21692 33844 21698 33856
rect 22204 33844 22232 33943
rect 23934 33940 23940 33952
rect 23992 33940 23998 33992
rect 24210 33940 24216 33992
rect 24268 33980 24274 33992
rect 24305 33983 24363 33989
rect 24305 33980 24317 33983
rect 24268 33952 24317 33980
rect 24268 33940 24274 33952
rect 24305 33949 24317 33952
rect 24351 33949 24363 33983
rect 24305 33943 24363 33949
rect 24581 33983 24639 33989
rect 24581 33949 24593 33983
rect 24627 33980 24639 33983
rect 24946 33980 24952 33992
rect 24627 33952 24952 33980
rect 24627 33949 24639 33952
rect 24581 33943 24639 33949
rect 24946 33940 24952 33952
rect 25004 33940 25010 33992
rect 26513 33983 26571 33989
rect 26513 33980 26525 33983
rect 25240 33952 26525 33980
rect 22370 33844 22376 33856
rect 21692 33816 22376 33844
rect 21692 33804 21698 33816
rect 22370 33804 22376 33816
rect 22428 33844 22434 33856
rect 24210 33844 24216 33856
rect 22428 33816 24216 33844
rect 22428 33804 22434 33816
rect 24210 33804 24216 33816
rect 24268 33804 24274 33856
rect 24670 33804 24676 33856
rect 24728 33844 24734 33856
rect 25240 33844 25268 33952
rect 26513 33949 26525 33952
rect 26559 33980 26571 33983
rect 28169 33983 28227 33989
rect 26559 33952 26924 33980
rect 26559 33949 26571 33952
rect 26513 33943 26571 33949
rect 25866 33844 25872 33856
rect 24728 33816 25268 33844
rect 25827 33816 25872 33844
rect 24728 33804 24734 33816
rect 25866 33804 25872 33816
rect 25924 33804 25930 33856
rect 25958 33804 25964 33856
rect 26016 33844 26022 33856
rect 26789 33847 26847 33853
rect 26789 33844 26801 33847
rect 26016 33816 26801 33844
rect 26016 33804 26022 33816
rect 26789 33813 26801 33816
rect 26835 33813 26847 33847
rect 26896 33844 26924 33952
rect 28169 33949 28181 33983
rect 28215 33980 28227 33983
rect 28902 33980 28908 33992
rect 28215 33952 28908 33980
rect 28215 33949 28227 33952
rect 28169 33943 28227 33949
rect 28902 33940 28908 33952
rect 28960 33940 28966 33992
rect 31018 33980 31024 33992
rect 30979 33952 31024 33980
rect 31018 33940 31024 33952
rect 31076 33980 31082 33992
rect 32861 33983 32919 33989
rect 32861 33980 32873 33983
rect 31076 33952 32873 33980
rect 31076 33940 31082 33952
rect 32324 33921 32352 33952
rect 32861 33949 32873 33952
rect 32907 33949 32919 33983
rect 32861 33943 32919 33949
rect 33686 33940 33692 33992
rect 33744 33980 33750 33992
rect 33873 33983 33931 33989
rect 33873 33980 33885 33983
rect 33744 33952 33885 33980
rect 33744 33940 33750 33952
rect 33873 33949 33885 33952
rect 33919 33949 33931 33983
rect 36170 33980 36176 33992
rect 36131 33952 36176 33980
rect 33873 33943 33931 33949
rect 36170 33940 36176 33952
rect 36228 33940 36234 33992
rect 36630 33940 36636 33992
rect 36688 33980 36694 33992
rect 36725 33983 36783 33989
rect 36725 33980 36737 33983
rect 36688 33952 36737 33980
rect 36688 33940 36694 33952
rect 36725 33949 36737 33952
rect 36771 33949 36783 33983
rect 37182 33980 37188 33992
rect 37143 33952 37188 33980
rect 36725 33943 36783 33949
rect 37182 33940 37188 33952
rect 37240 33940 37246 33992
rect 32309 33915 32367 33921
rect 32309 33881 32321 33915
rect 32355 33881 32367 33915
rect 32309 33875 32367 33881
rect 29086 33844 29092 33856
rect 26896 33816 29092 33844
rect 26789 33807 26847 33813
rect 29086 33804 29092 33816
rect 29144 33804 29150 33856
rect 30466 33844 30472 33856
rect 30427 33816 30472 33844
rect 30466 33804 30472 33816
rect 30524 33804 30530 33856
rect 35253 33847 35311 33853
rect 35253 33813 35265 33847
rect 35299 33844 35311 33847
rect 35342 33844 35348 33856
rect 35299 33816 35348 33844
rect 35299 33813 35311 33816
rect 35253 33807 35311 33813
rect 35342 33804 35348 33816
rect 35400 33804 35406 33856
rect 1104 33754 38824 33776
rect 1104 33702 4246 33754
rect 4298 33702 4310 33754
rect 4362 33702 4374 33754
rect 4426 33702 4438 33754
rect 4490 33702 34966 33754
rect 35018 33702 35030 33754
rect 35082 33702 35094 33754
rect 35146 33702 35158 33754
rect 35210 33702 38824 33754
rect 1104 33680 38824 33702
rect 1854 33640 1860 33652
rect 1815 33612 1860 33640
rect 1854 33600 1860 33612
rect 1912 33600 1918 33652
rect 4157 33643 4215 33649
rect 4157 33609 4169 33643
rect 4203 33640 4215 33643
rect 4614 33640 4620 33652
rect 4203 33612 4620 33640
rect 4203 33609 4215 33612
rect 4157 33603 4215 33609
rect 4614 33600 4620 33612
rect 4672 33600 4678 33652
rect 7006 33640 7012 33652
rect 6196 33612 7012 33640
rect 6086 33572 6092 33584
rect 4540 33544 6092 33572
rect 1394 33464 1400 33516
rect 1452 33504 1458 33516
rect 2593 33507 2651 33513
rect 2593 33504 2605 33507
rect 1452 33476 2605 33504
rect 1452 33464 1458 33476
rect 2593 33473 2605 33476
rect 2639 33504 2651 33507
rect 3970 33504 3976 33516
rect 2639 33476 3976 33504
rect 2639 33473 2651 33476
rect 2593 33467 2651 33473
rect 3970 33464 3976 33476
rect 4028 33464 4034 33516
rect 1486 33436 1492 33448
rect 1447 33408 1492 33436
rect 1486 33396 1492 33408
rect 1544 33396 1550 33448
rect 1670 33436 1676 33448
rect 1631 33408 1676 33436
rect 1670 33396 1676 33408
rect 1728 33396 1734 33448
rect 2869 33439 2927 33445
rect 2869 33405 2881 33439
rect 2915 33436 2927 33439
rect 4154 33436 4160 33448
rect 2915 33408 4160 33436
rect 2915 33405 2927 33408
rect 2869 33399 2927 33405
rect 4154 33396 4160 33408
rect 4212 33396 4218 33448
rect 1578 33368 1584 33380
rect 1539 33340 1584 33368
rect 1578 33328 1584 33340
rect 1636 33328 1642 33380
rect 1596 33300 1624 33328
rect 4540 33300 4568 33544
rect 6086 33532 6092 33544
rect 6144 33532 6150 33584
rect 6196 33504 6224 33612
rect 7006 33600 7012 33612
rect 7064 33600 7070 33652
rect 9674 33600 9680 33652
rect 9732 33640 9738 33652
rect 9769 33643 9827 33649
rect 9769 33640 9781 33643
rect 9732 33612 9781 33640
rect 9732 33600 9738 33612
rect 9769 33609 9781 33612
rect 9815 33609 9827 33643
rect 9769 33603 9827 33609
rect 11885 33643 11943 33649
rect 11885 33609 11897 33643
rect 11931 33640 11943 33643
rect 13262 33640 13268 33652
rect 11931 33612 13268 33640
rect 11931 33609 11943 33612
rect 11885 33603 11943 33609
rect 13262 33600 13268 33612
rect 13320 33600 13326 33652
rect 15933 33643 15991 33649
rect 15933 33609 15945 33643
rect 15979 33640 15991 33643
rect 16390 33640 16396 33652
rect 15979 33612 16396 33640
rect 15979 33609 15991 33612
rect 15933 33603 15991 33609
rect 16390 33600 16396 33612
rect 16448 33600 16454 33652
rect 16574 33600 16580 33652
rect 16632 33600 16638 33652
rect 18046 33600 18052 33652
rect 18104 33640 18110 33652
rect 18141 33643 18199 33649
rect 18141 33640 18153 33643
rect 18104 33612 18153 33640
rect 18104 33600 18110 33612
rect 18141 33609 18153 33612
rect 18187 33609 18199 33643
rect 18141 33603 18199 33609
rect 22370 33600 22376 33652
rect 22428 33640 22434 33652
rect 22465 33643 22523 33649
rect 22465 33640 22477 33643
rect 22428 33612 22477 33640
rect 22428 33600 22434 33612
rect 22465 33609 22477 33612
rect 22511 33609 22523 33643
rect 23934 33640 23940 33652
rect 23895 33612 23940 33640
rect 22465 33603 22523 33609
rect 23934 33600 23940 33612
rect 23992 33600 23998 33652
rect 24946 33640 24952 33652
rect 24907 33612 24952 33640
rect 24946 33600 24952 33612
rect 25004 33600 25010 33652
rect 33042 33600 33048 33652
rect 33100 33640 33106 33652
rect 33505 33643 33563 33649
rect 33505 33640 33517 33643
rect 33100 33612 33517 33640
rect 33100 33600 33106 33612
rect 33505 33609 33517 33612
rect 33551 33609 33563 33643
rect 33505 33603 33563 33609
rect 37182 33600 37188 33652
rect 37240 33640 37246 33652
rect 37829 33643 37887 33649
rect 37829 33640 37841 33643
rect 37240 33612 37841 33640
rect 37240 33600 37246 33612
rect 37829 33609 37841 33612
rect 37875 33609 37887 33643
rect 37829 33603 37887 33609
rect 7558 33572 7564 33584
rect 7519 33544 7564 33572
rect 7558 33532 7564 33544
rect 7616 33532 7622 33584
rect 7926 33532 7932 33584
rect 7984 33572 7990 33584
rect 12529 33575 12587 33581
rect 7984 33544 11100 33572
rect 7984 33532 7990 33544
rect 5552 33476 6224 33504
rect 4614 33396 4620 33448
rect 4672 33436 4678 33448
rect 4709 33439 4767 33445
rect 4709 33436 4721 33439
rect 4672 33408 4721 33436
rect 4672 33396 4678 33408
rect 4709 33405 4721 33408
rect 4755 33405 4767 33439
rect 4709 33399 4767 33405
rect 5552 33380 5580 33476
rect 6638 33464 6644 33516
rect 6696 33504 6702 33516
rect 6696 33476 7788 33504
rect 6696 33464 6702 33476
rect 5718 33436 5724 33448
rect 5679 33408 5724 33436
rect 5718 33396 5724 33408
rect 5776 33396 5782 33448
rect 6914 33436 6920 33448
rect 5920 33408 6920 33436
rect 5534 33368 5540 33380
rect 5495 33340 5540 33368
rect 5534 33328 5540 33340
rect 5592 33328 5598 33380
rect 5920 33377 5948 33408
rect 6914 33396 6920 33408
rect 6972 33396 6978 33448
rect 7024 33445 7052 33476
rect 7009 33439 7067 33445
rect 7009 33405 7021 33439
rect 7055 33405 7067 33439
rect 7466 33436 7472 33448
rect 7427 33408 7472 33436
rect 7009 33399 7067 33405
rect 7466 33396 7472 33408
rect 7524 33396 7530 33448
rect 7650 33436 7656 33448
rect 7611 33408 7656 33436
rect 7650 33396 7656 33408
rect 7708 33396 7714 33448
rect 7760 33436 7788 33476
rect 7926 33436 7932 33448
rect 7760 33408 7932 33436
rect 7926 33396 7932 33408
rect 7984 33396 7990 33448
rect 8573 33439 8631 33445
rect 8573 33405 8585 33439
rect 8619 33436 8631 33439
rect 8754 33436 8760 33448
rect 8619 33408 8760 33436
rect 8619 33405 8631 33408
rect 8573 33399 8631 33405
rect 8754 33396 8760 33408
rect 8812 33396 8818 33448
rect 8941 33439 8999 33445
rect 8941 33405 8953 33439
rect 8987 33405 8999 33439
rect 9122 33436 9128 33448
rect 9083 33408 9128 33436
rect 8941 33399 8999 33405
rect 5905 33371 5963 33377
rect 5905 33337 5917 33371
rect 5951 33337 5963 33371
rect 5905 33331 5963 33337
rect 6273 33371 6331 33377
rect 6273 33337 6285 33371
rect 6319 33368 6331 33371
rect 8662 33368 8668 33380
rect 6319 33340 8668 33368
rect 6319 33337 6331 33340
rect 6273 33331 6331 33337
rect 8662 33328 8668 33340
rect 8720 33328 8726 33380
rect 1596 33272 4568 33300
rect 4614 33260 4620 33312
rect 4672 33300 4678 33312
rect 4893 33303 4951 33309
rect 4893 33300 4905 33303
rect 4672 33272 4905 33300
rect 4672 33260 4678 33272
rect 4893 33269 4905 33272
rect 4939 33269 4951 33303
rect 4893 33263 4951 33269
rect 5813 33303 5871 33309
rect 5813 33269 5825 33303
rect 5859 33300 5871 33303
rect 7282 33300 7288 33312
rect 5859 33272 7288 33300
rect 5859 33269 5871 33272
rect 5813 33263 5871 33269
rect 7282 33260 7288 33272
rect 7340 33260 7346 33312
rect 8478 33260 8484 33312
rect 8536 33300 8542 33312
rect 8956 33300 8984 33399
rect 9122 33396 9128 33408
rect 9180 33396 9186 33448
rect 9766 33436 9772 33448
rect 9727 33408 9772 33436
rect 9766 33396 9772 33408
rect 9824 33396 9830 33448
rect 11072 33445 11100 33544
rect 12529 33541 12541 33575
rect 12575 33541 12587 33575
rect 12529 33535 12587 33541
rect 16485 33575 16543 33581
rect 16485 33541 16497 33575
rect 16531 33541 16543 33575
rect 16485 33535 16543 33541
rect 12544 33504 12572 33535
rect 11624 33476 12572 33504
rect 11057 33439 11115 33445
rect 11057 33405 11069 33439
rect 11103 33405 11115 33439
rect 11238 33436 11244 33448
rect 11199 33408 11244 33436
rect 11057 33399 11115 33405
rect 11072 33368 11100 33399
rect 11238 33396 11244 33408
rect 11296 33396 11302 33448
rect 11624 33445 11652 33476
rect 12618 33464 12624 33516
rect 12676 33464 12682 33516
rect 15749 33507 15807 33513
rect 12728 33476 15148 33504
rect 11609 33439 11667 33445
rect 11609 33405 11621 33439
rect 11655 33405 11667 33439
rect 11609 33399 11667 33405
rect 12529 33439 12587 33445
rect 12529 33405 12541 33439
rect 12575 33436 12587 33439
rect 12636 33436 12664 33464
rect 12575 33408 12664 33436
rect 12575 33405 12587 33408
rect 12529 33399 12587 33405
rect 12728 33368 12756 33476
rect 12986 33436 12992 33448
rect 12947 33408 12992 33436
rect 12986 33396 12992 33408
rect 13044 33396 13050 33448
rect 13354 33396 13360 33448
rect 13412 33436 13418 33448
rect 13909 33439 13967 33445
rect 13412 33408 13457 33436
rect 13412 33396 13418 33408
rect 13909 33405 13921 33439
rect 13955 33436 13967 33439
rect 13998 33436 14004 33448
rect 13955 33408 14004 33436
rect 13955 33405 13967 33408
rect 13909 33399 13967 33405
rect 13998 33396 14004 33408
rect 14056 33396 14062 33448
rect 14182 33436 14188 33448
rect 14143 33408 14188 33436
rect 14182 33396 14188 33408
rect 14240 33396 14246 33448
rect 15120 33445 15148 33476
rect 15749 33473 15761 33507
rect 15795 33504 15807 33507
rect 16390 33504 16396 33516
rect 15795 33476 16396 33504
rect 15795 33473 15807 33476
rect 15749 33467 15807 33473
rect 16390 33464 16396 33476
rect 16448 33464 16454 33516
rect 15105 33439 15163 33445
rect 15105 33405 15117 33439
rect 15151 33436 15163 33439
rect 15657 33439 15715 33445
rect 15151 33408 15240 33436
rect 15151 33405 15163 33408
rect 15105 33399 15163 33405
rect 11072 33340 12756 33368
rect 11238 33300 11244 33312
rect 8536 33272 11244 33300
rect 8536 33260 8542 33272
rect 11238 33260 11244 33272
rect 11296 33260 11302 33312
rect 15212 33300 15240 33408
rect 15657 33405 15669 33439
rect 15703 33436 15715 33439
rect 16500 33436 16528 33535
rect 16592 33504 16620 33600
rect 17221 33507 17279 33513
rect 17221 33504 17233 33507
rect 16592 33476 17233 33504
rect 17221 33473 17233 33476
rect 17267 33473 17279 33507
rect 23014 33504 23020 33516
rect 17221 33467 17279 33473
rect 20088 33476 23020 33504
rect 15703 33408 16528 33436
rect 16577 33439 16635 33445
rect 15703 33405 15715 33408
rect 15657 33399 15715 33405
rect 16577 33405 16589 33439
rect 16623 33436 16635 33439
rect 17126 33436 17132 33448
rect 16623 33408 16988 33436
rect 17087 33408 17132 33436
rect 16623 33405 16635 33408
rect 16577 33399 16635 33405
rect 16960 33368 16988 33408
rect 17126 33396 17132 33408
rect 17184 33396 17190 33448
rect 17236 33436 17264 33467
rect 18049 33439 18107 33445
rect 18049 33436 18061 33439
rect 17236 33408 18061 33436
rect 18049 33405 18061 33408
rect 18095 33405 18107 33439
rect 18414 33436 18420 33448
rect 18375 33408 18420 33436
rect 18049 33399 18107 33405
rect 18414 33396 18420 33408
rect 18472 33396 18478 33448
rect 19061 33439 19119 33445
rect 19061 33405 19073 33439
rect 19107 33405 19119 33439
rect 19334 33436 19340 33448
rect 19295 33408 19340 33436
rect 19061 33399 19119 33405
rect 17218 33368 17224 33380
rect 16960 33340 17224 33368
rect 17218 33328 17224 33340
rect 17276 33328 17282 33380
rect 19076 33368 19104 33399
rect 19334 33396 19340 33408
rect 19392 33396 19398 33448
rect 19426 33396 19432 33448
rect 19484 33436 19490 33448
rect 20088 33445 20116 33476
rect 23014 33464 23020 33476
rect 23072 33464 23078 33516
rect 23842 33464 23848 33516
rect 23900 33504 23906 33516
rect 29825 33507 29883 33513
rect 23900 33476 24808 33504
rect 23900 33464 23906 33476
rect 20073 33439 20131 33445
rect 20073 33436 20085 33439
rect 19484 33408 20085 33436
rect 19484 33396 19490 33408
rect 20073 33405 20085 33408
rect 20119 33405 20131 33439
rect 20346 33436 20352 33448
rect 20307 33408 20352 33436
rect 20073 33399 20131 33405
rect 20346 33396 20352 33408
rect 20404 33396 20410 33448
rect 22189 33439 22247 33445
rect 22189 33436 22201 33439
rect 22020 33408 22201 33436
rect 19978 33368 19984 33380
rect 19076 33340 19984 33368
rect 19978 33328 19984 33340
rect 20036 33328 20042 33380
rect 20070 33300 20076 33312
rect 15212 33272 20076 33300
rect 20070 33260 20076 33272
rect 20128 33260 20134 33312
rect 20622 33260 20628 33312
rect 20680 33300 20686 33312
rect 21453 33303 21511 33309
rect 21453 33300 21465 33303
rect 20680 33272 21465 33300
rect 20680 33260 20686 33272
rect 21453 33269 21465 33272
rect 21499 33269 21511 33303
rect 22020 33300 22048 33408
rect 22189 33405 22201 33408
rect 22235 33405 22247 33439
rect 22189 33399 22247 33405
rect 22281 33439 22339 33445
rect 22281 33405 22293 33439
rect 22327 33436 22339 33439
rect 22646 33436 22652 33448
rect 22327 33408 22652 33436
rect 22327 33405 22339 33408
rect 22281 33399 22339 33405
rect 22097 33371 22155 33377
rect 22097 33337 22109 33371
rect 22143 33368 22155 33371
rect 22296 33368 22324 33399
rect 22646 33396 22652 33408
rect 22704 33396 22710 33448
rect 23382 33396 23388 33448
rect 23440 33436 23446 33448
rect 23661 33439 23719 33445
rect 23661 33436 23673 33439
rect 23440 33408 23673 33436
rect 23440 33396 23446 33408
rect 23661 33405 23673 33408
rect 23707 33405 23719 33439
rect 23661 33399 23719 33405
rect 23750 33396 23756 33448
rect 23808 33436 23814 33448
rect 24670 33436 24676 33448
rect 23808 33408 23853 33436
rect 24631 33408 24676 33436
rect 23808 33396 23814 33408
rect 24670 33396 24676 33408
rect 24728 33396 24734 33448
rect 24780 33445 24808 33476
rect 29825 33473 29837 33507
rect 29871 33504 29883 33507
rect 30650 33504 30656 33516
rect 29871 33476 30656 33504
rect 29871 33473 29883 33476
rect 29825 33467 29883 33473
rect 30650 33464 30656 33476
rect 30708 33464 30714 33516
rect 31846 33464 31852 33516
rect 31904 33504 31910 33516
rect 32401 33507 32459 33513
rect 32401 33504 32413 33507
rect 31904 33476 32413 33504
rect 31904 33464 31910 33476
rect 32401 33473 32413 33476
rect 32447 33473 32459 33507
rect 32401 33467 32459 33473
rect 35621 33507 35679 33513
rect 35621 33473 35633 33507
rect 35667 33504 35679 33507
rect 36630 33504 36636 33516
rect 35667 33476 36636 33504
rect 35667 33473 35679 33476
rect 35621 33467 35679 33473
rect 36630 33464 36636 33476
rect 36688 33464 36694 33516
rect 24765 33439 24823 33445
rect 24765 33405 24777 33439
rect 24811 33405 24823 33439
rect 25774 33436 25780 33448
rect 25735 33408 25780 33436
rect 24765 33399 24823 33405
rect 25774 33396 25780 33408
rect 25832 33396 25838 33448
rect 26053 33439 26111 33445
rect 26053 33405 26065 33439
rect 26099 33436 26111 33439
rect 28169 33439 28227 33445
rect 26099 33408 27384 33436
rect 26099 33405 26111 33408
rect 26053 33399 26111 33405
rect 22143 33340 22324 33368
rect 22143 33337 22155 33340
rect 22097 33331 22155 33337
rect 23014 33328 23020 33380
rect 23072 33368 23078 33380
rect 24688 33368 24716 33396
rect 23072 33340 24716 33368
rect 23072 33328 23078 33340
rect 23382 33300 23388 33312
rect 22020 33272 23388 33300
rect 21453 33263 21511 33269
rect 23382 33260 23388 33272
rect 23440 33260 23446 33312
rect 27154 33300 27160 33312
rect 27115 33272 27160 33300
rect 27154 33260 27160 33272
rect 27212 33260 27218 33312
rect 27356 33300 27384 33408
rect 28169 33405 28181 33439
rect 28215 33405 28227 33439
rect 28350 33436 28356 33448
rect 28311 33408 28356 33436
rect 28169 33399 28227 33405
rect 28184 33368 28212 33399
rect 28350 33396 28356 33408
rect 28408 33396 28414 33448
rect 28534 33436 28540 33448
rect 28495 33408 28540 33436
rect 28534 33396 28540 33408
rect 28592 33396 28598 33448
rect 28902 33396 28908 33448
rect 28960 33436 28966 33448
rect 29549 33439 29607 33445
rect 29549 33436 29561 33439
rect 28960 33408 29561 33436
rect 28960 33396 28966 33408
rect 29549 33405 29561 33408
rect 29595 33436 29607 33439
rect 30742 33436 30748 33448
rect 29595 33408 30748 33436
rect 29595 33405 29607 33408
rect 29549 33399 29607 33405
rect 30742 33396 30748 33408
rect 30800 33396 30806 33448
rect 31386 33396 31392 33448
rect 31444 33436 31450 33448
rect 32125 33439 32183 33445
rect 32125 33436 32137 33439
rect 31444 33408 32137 33436
rect 31444 33396 31450 33408
rect 32125 33405 32137 33408
rect 32171 33405 32183 33439
rect 35526 33436 35532 33448
rect 35487 33408 35532 33436
rect 32125 33399 32183 33405
rect 35526 33396 35532 33408
rect 35584 33396 35590 33448
rect 35897 33439 35955 33445
rect 35897 33405 35909 33439
rect 35943 33405 35955 33439
rect 36446 33436 36452 33448
rect 36407 33408 36452 33436
rect 35897 33399 35955 33405
rect 29362 33368 29368 33380
rect 28184 33340 29368 33368
rect 29362 33328 29368 33340
rect 29420 33328 29426 33380
rect 30929 33303 30987 33309
rect 30929 33300 30941 33303
rect 27356 33272 30941 33300
rect 30929 33269 30941 33272
rect 30975 33269 30987 33303
rect 35912 33300 35940 33399
rect 36446 33396 36452 33408
rect 36504 33396 36510 33448
rect 36722 33436 36728 33448
rect 36683 33408 36728 33436
rect 36722 33396 36728 33408
rect 36780 33396 36786 33448
rect 36262 33300 36268 33312
rect 35912 33272 36268 33300
rect 30929 33263 30987 33269
rect 36262 33260 36268 33272
rect 36320 33260 36326 33312
rect 1104 33210 38824 33232
rect 1104 33158 19606 33210
rect 19658 33158 19670 33210
rect 19722 33158 19734 33210
rect 19786 33158 19798 33210
rect 19850 33158 38824 33210
rect 1104 33136 38824 33158
rect 5626 33096 5632 33108
rect 5587 33068 5632 33096
rect 5626 33056 5632 33068
rect 5684 33056 5690 33108
rect 6362 33056 6368 33108
rect 6420 33096 6426 33108
rect 11238 33096 11244 33108
rect 6420 33068 10916 33096
rect 11151 33068 11244 33096
rect 6420 33056 6426 33068
rect 1486 32988 1492 33040
rect 1544 33028 1550 33040
rect 2041 33031 2099 33037
rect 2041 33028 2053 33031
rect 1544 33000 2053 33028
rect 1544 32988 1550 33000
rect 2041 32997 2053 33000
rect 2087 32997 2099 33031
rect 2041 32991 2099 32997
rect 4065 33031 4123 33037
rect 4065 32997 4077 33031
rect 4111 33028 4123 33031
rect 4154 33028 4160 33040
rect 4111 33000 4160 33028
rect 4111 32997 4123 33000
rect 4065 32991 4123 32997
rect 4154 32988 4160 33000
rect 4212 32988 4218 33040
rect 4706 32988 4712 33040
rect 4764 33028 4770 33040
rect 8478 33028 8484 33040
rect 4764 33000 5580 33028
rect 4764 32988 4770 33000
rect 2590 32960 2596 32972
rect 2551 32932 2596 32960
rect 2590 32920 2596 32932
rect 2648 32920 2654 32972
rect 2774 32920 2780 32972
rect 2832 32960 2838 32972
rect 2958 32960 2964 32972
rect 2832 32932 2877 32960
rect 2919 32932 2964 32960
rect 2832 32920 2838 32932
rect 2958 32920 2964 32932
rect 3016 32920 3022 32972
rect 3142 32960 3148 32972
rect 3103 32932 3148 32960
rect 3142 32920 3148 32932
rect 3200 32920 3206 32972
rect 3234 32920 3240 32972
rect 3292 32960 3298 32972
rect 3329 32963 3387 32969
rect 3329 32960 3341 32963
rect 3292 32932 3341 32960
rect 3292 32920 3298 32932
rect 3329 32929 3341 32932
rect 3375 32929 3387 32963
rect 3329 32923 3387 32929
rect 3602 32920 3608 32972
rect 3660 32960 3666 32972
rect 5552 32969 5580 33000
rect 8220 33000 8484 33028
rect 4893 32963 4951 32969
rect 4893 32960 4905 32963
rect 3660 32932 4905 32960
rect 3660 32920 3666 32932
rect 4893 32929 4905 32932
rect 4939 32929 4951 32963
rect 4893 32923 4951 32929
rect 5537 32963 5595 32969
rect 5537 32929 5549 32963
rect 5583 32929 5595 32963
rect 5537 32923 5595 32929
rect 6270 32920 6276 32972
rect 6328 32960 6334 32972
rect 8220 32969 8248 33000
rect 8478 32988 8484 33000
rect 8536 32988 8542 33040
rect 10888 33028 10916 33068
rect 11238 33056 11244 33068
rect 11296 33096 11302 33108
rect 12986 33096 12992 33108
rect 11296 33068 12992 33096
rect 11296 33056 11302 33068
rect 12986 33056 12992 33068
rect 13044 33056 13050 33108
rect 15286 33056 15292 33108
rect 15344 33096 15350 33108
rect 19150 33096 19156 33108
rect 15344 33068 19156 33096
rect 15344 33056 15350 33068
rect 11330 33028 11336 33040
rect 10888 33000 11336 33028
rect 11330 32988 11336 33000
rect 11388 32988 11394 33040
rect 13633 33031 13691 33037
rect 13633 32997 13645 33031
rect 13679 33028 13691 33031
rect 13998 33028 14004 33040
rect 13679 33000 14004 33028
rect 13679 32997 13691 33000
rect 13633 32991 13691 32997
rect 13998 32988 14004 33000
rect 14056 32988 14062 33040
rect 7009 32963 7067 32969
rect 7009 32960 7021 32963
rect 6328 32932 7021 32960
rect 6328 32920 6334 32932
rect 7009 32929 7021 32932
rect 7055 32929 7067 32963
rect 7009 32923 7067 32929
rect 8205 32963 8263 32969
rect 8205 32929 8217 32963
rect 8251 32929 8263 32963
rect 8386 32960 8392 32972
rect 8347 32932 8392 32960
rect 8205 32923 8263 32929
rect 8386 32920 8392 32932
rect 8444 32920 8450 32972
rect 8570 32960 8576 32972
rect 8531 32932 8576 32960
rect 8570 32920 8576 32932
rect 8628 32920 8634 32972
rect 8754 32960 8760 32972
rect 8715 32932 8760 32960
rect 8754 32920 8760 32932
rect 8812 32920 8818 32972
rect 8846 32920 8852 32972
rect 8904 32960 8910 32972
rect 8941 32963 8999 32969
rect 8941 32960 8953 32963
rect 8904 32932 8953 32960
rect 8904 32920 8910 32932
rect 8941 32929 8953 32932
rect 8987 32929 8999 32963
rect 8941 32923 8999 32929
rect 9677 32963 9735 32969
rect 9677 32929 9689 32963
rect 9723 32960 9735 32963
rect 11146 32960 11152 32972
rect 9723 32932 11152 32960
rect 9723 32929 9735 32932
rect 9677 32923 9735 32929
rect 11146 32920 11152 32932
rect 11204 32960 11210 32972
rect 11977 32963 12035 32969
rect 11977 32960 11989 32963
rect 11204 32932 11989 32960
rect 11204 32920 11210 32932
rect 11977 32929 11989 32932
rect 12023 32960 12035 32963
rect 12342 32960 12348 32972
rect 12023 32932 12348 32960
rect 12023 32929 12035 32932
rect 11977 32923 12035 32929
rect 12342 32920 12348 32932
rect 12400 32920 12406 32972
rect 14461 32963 14519 32969
rect 14461 32929 14473 32963
rect 14507 32960 14519 32963
rect 15562 32960 15568 32972
rect 14507 32932 15424 32960
rect 15523 32932 15568 32960
rect 14507 32929 14519 32932
rect 14461 32923 14519 32929
rect 4062 32852 4068 32904
rect 4120 32892 4126 32904
rect 4617 32895 4675 32901
rect 4617 32892 4629 32895
rect 4120 32864 4629 32892
rect 4120 32852 4126 32864
rect 4617 32861 4629 32864
rect 4663 32861 4675 32895
rect 4617 32855 4675 32861
rect 4706 32852 4712 32904
rect 4764 32892 4770 32904
rect 5077 32895 5135 32901
rect 5077 32892 5089 32895
rect 4764 32864 5089 32892
rect 4764 32852 4770 32864
rect 5077 32861 5089 32864
rect 5123 32861 5135 32895
rect 6178 32892 6184 32904
rect 6139 32864 6184 32892
rect 5077 32855 5135 32861
rect 6178 32852 6184 32864
rect 6236 32852 6242 32904
rect 6733 32895 6791 32901
rect 6733 32861 6745 32895
rect 6779 32861 6791 32895
rect 6733 32855 6791 32861
rect 6748 32824 6776 32855
rect 6822 32852 6828 32904
rect 6880 32892 6886 32904
rect 7193 32895 7251 32901
rect 7193 32892 7205 32895
rect 6880 32864 7205 32892
rect 6880 32852 6886 32864
rect 7193 32861 7205 32864
rect 7239 32861 7251 32895
rect 7193 32855 7251 32861
rect 7653 32895 7711 32901
rect 7653 32861 7665 32895
rect 7699 32892 7711 32895
rect 9582 32892 9588 32904
rect 7699 32864 9588 32892
rect 7699 32861 7711 32864
rect 7653 32855 7711 32861
rect 9582 32852 9588 32864
rect 9640 32852 9646 32904
rect 9950 32892 9956 32904
rect 9911 32864 9956 32892
rect 9950 32852 9956 32864
rect 10008 32852 10014 32904
rect 12250 32892 12256 32904
rect 12211 32864 12256 32892
rect 12250 32852 12256 32864
rect 12308 32852 12314 32904
rect 15286 32892 15292 32904
rect 15247 32864 15292 32892
rect 15286 32852 15292 32864
rect 15344 32852 15350 32904
rect 15396 32892 15424 32932
rect 15562 32920 15568 32932
rect 15620 32920 15626 32972
rect 18156 32969 18184 33068
rect 19150 33056 19156 33068
rect 19208 33056 19214 33108
rect 36633 33099 36691 33105
rect 36633 33065 36645 33099
rect 36679 33096 36691 33099
rect 36722 33096 36728 33108
rect 36679 33068 36728 33096
rect 36679 33065 36691 33068
rect 36633 33059 36691 33065
rect 36722 33056 36728 33068
rect 36780 33056 36786 33108
rect 29086 32988 29092 33040
rect 29144 33028 29150 33040
rect 29144 33000 34468 33028
rect 29144 32988 29150 33000
rect 17405 32963 17463 32969
rect 17405 32929 17417 32963
rect 17451 32929 17463 32963
rect 17405 32923 17463 32929
rect 18148 32963 18206 32969
rect 18148 32929 18160 32963
rect 18194 32929 18206 32963
rect 18148 32923 18206 32929
rect 16942 32892 16948 32904
rect 15396 32864 16948 32892
rect 16942 32852 16948 32864
rect 17000 32852 17006 32904
rect 7558 32824 7564 32836
rect 6748 32796 7564 32824
rect 7558 32784 7564 32796
rect 7616 32784 7622 32836
rect 7374 32716 7380 32768
rect 7432 32756 7438 32768
rect 9214 32756 9220 32768
rect 7432 32728 9220 32756
rect 7432 32716 7438 32728
rect 9214 32716 9220 32728
rect 9272 32716 9278 32768
rect 14645 32759 14703 32765
rect 14645 32725 14657 32759
rect 14691 32756 14703 32759
rect 16298 32756 16304 32768
rect 14691 32728 16304 32756
rect 14691 32725 14703 32728
rect 14645 32719 14703 32725
rect 16298 32716 16304 32728
rect 16356 32716 16362 32768
rect 16850 32756 16856 32768
rect 16811 32728 16856 32756
rect 16850 32716 16856 32728
rect 16908 32716 16914 32768
rect 17420 32756 17448 32923
rect 19978 32920 19984 32972
rect 20036 32960 20042 32972
rect 20530 32960 20536 32972
rect 20036 32932 20536 32960
rect 20036 32920 20042 32932
rect 20530 32920 20536 32932
rect 20588 32960 20594 32972
rect 20901 32963 20959 32969
rect 20901 32960 20913 32963
rect 20588 32932 20913 32960
rect 20588 32920 20594 32932
rect 20901 32929 20913 32932
rect 20947 32929 20959 32963
rect 21634 32960 21640 32972
rect 21595 32932 21640 32960
rect 20901 32923 20959 32929
rect 21634 32920 21640 32932
rect 21692 32920 21698 32972
rect 21913 32963 21971 32969
rect 21913 32929 21925 32963
rect 21959 32960 21971 32963
rect 22370 32960 22376 32972
rect 21959 32932 22376 32960
rect 21959 32929 21971 32932
rect 21913 32923 21971 32929
rect 22370 32920 22376 32932
rect 22428 32920 22434 32972
rect 24305 32963 24363 32969
rect 24305 32929 24317 32963
rect 24351 32960 24363 32963
rect 25958 32960 25964 32972
rect 24351 32932 25964 32960
rect 24351 32929 24363 32932
rect 24305 32923 24363 32929
rect 25958 32920 25964 32932
rect 26016 32920 26022 32972
rect 26789 32963 26847 32969
rect 26789 32929 26801 32963
rect 26835 32960 26847 32963
rect 27154 32960 27160 32972
rect 26835 32932 27160 32960
rect 26835 32929 26847 32932
rect 26789 32923 26847 32929
rect 27154 32920 27160 32932
rect 27212 32920 27218 32972
rect 28626 32960 28632 32972
rect 28587 32932 28632 32960
rect 28626 32920 28632 32932
rect 28684 32920 28690 32972
rect 29365 32963 29423 32969
rect 29365 32929 29377 32963
rect 29411 32960 29423 32963
rect 29822 32960 29828 32972
rect 29411 32932 29828 32960
rect 29411 32929 29423 32932
rect 29365 32923 29423 32929
rect 29822 32920 29828 32932
rect 29880 32920 29886 32972
rect 30558 32960 30564 32972
rect 30519 32932 30564 32960
rect 30558 32920 30564 32932
rect 30616 32920 30622 32972
rect 31205 32963 31263 32969
rect 31205 32929 31217 32963
rect 31251 32960 31263 32963
rect 33226 32960 33232 32972
rect 31251 32932 32904 32960
rect 33187 32932 33232 32960
rect 31251 32929 31263 32932
rect 31205 32923 31263 32929
rect 17678 32852 17684 32904
rect 17736 32892 17742 32904
rect 18417 32895 18475 32901
rect 18417 32892 18429 32895
rect 17736 32864 18429 32892
rect 17736 32852 17742 32864
rect 18417 32861 18429 32864
rect 18463 32861 18475 32895
rect 18417 32855 18475 32861
rect 23842 32852 23848 32904
rect 23900 32892 23906 32904
rect 24029 32895 24087 32901
rect 24029 32892 24041 32895
rect 23900 32864 24041 32892
rect 23900 32852 23906 32864
rect 24029 32861 24041 32864
rect 24075 32892 24087 32895
rect 24210 32892 24216 32904
rect 24075 32864 24216 32892
rect 24075 32861 24087 32864
rect 24029 32855 24087 32861
rect 24210 32852 24216 32864
rect 24268 32892 24274 32904
rect 26513 32895 26571 32901
rect 24268 32864 25820 32892
rect 24268 32852 24274 32864
rect 25792 32836 25820 32864
rect 26513 32861 26525 32895
rect 26559 32861 26571 32895
rect 26513 32855 26571 32861
rect 31481 32895 31539 32901
rect 31481 32861 31493 32895
rect 31527 32892 31539 32895
rect 31754 32892 31760 32904
rect 31527 32864 31760 32892
rect 31527 32861 31539 32864
rect 31481 32855 31539 32861
rect 17494 32784 17500 32836
rect 17552 32824 17558 32836
rect 17589 32827 17647 32833
rect 17589 32824 17601 32827
rect 17552 32796 17601 32824
rect 17552 32784 17558 32796
rect 17589 32793 17601 32796
rect 17635 32793 17647 32827
rect 17589 32787 17647 32793
rect 25774 32784 25780 32836
rect 25832 32824 25838 32836
rect 25958 32824 25964 32836
rect 25832 32796 25964 32824
rect 25832 32784 25838 32796
rect 25958 32784 25964 32796
rect 26016 32824 26022 32836
rect 26528 32824 26556 32855
rect 31754 32852 31760 32864
rect 31812 32852 31818 32904
rect 32766 32892 32772 32904
rect 32727 32864 32772 32892
rect 32766 32852 32772 32864
rect 32824 32852 32830 32904
rect 32876 32892 32904 32932
rect 33226 32920 33232 32932
rect 33284 32920 33290 32972
rect 33594 32960 33600 32972
rect 33555 32932 33600 32960
rect 33594 32920 33600 32932
rect 33652 32920 33658 32972
rect 34256 32969 34284 33000
rect 34241 32963 34299 32969
rect 34241 32929 34253 32963
rect 34287 32929 34299 32963
rect 34241 32923 34299 32929
rect 34333 32963 34391 32969
rect 34333 32929 34345 32963
rect 34379 32929 34391 32963
rect 34440 32960 34468 33000
rect 35342 32960 35348 32972
rect 34440 32932 34928 32960
rect 35303 32932 35348 32960
rect 34333 32923 34391 32929
rect 33505 32895 33563 32901
rect 33505 32892 33517 32895
rect 32876 32864 33517 32892
rect 33505 32861 33517 32864
rect 33551 32861 33563 32895
rect 33505 32855 33563 32861
rect 30742 32824 30748 32836
rect 26016 32796 26556 32824
rect 30703 32796 30748 32824
rect 26016 32784 26022 32796
rect 30742 32784 30748 32796
rect 30800 32784 30806 32836
rect 34348 32824 34376 32923
rect 34790 32892 34796 32904
rect 34751 32864 34796 32892
rect 34790 32852 34796 32864
rect 34848 32852 34854 32904
rect 34900 32892 34928 32932
rect 35342 32920 35348 32932
rect 35400 32920 35406 32972
rect 36354 32960 36360 32972
rect 36315 32932 36360 32960
rect 36354 32920 36360 32932
rect 36412 32920 36418 32972
rect 36909 32963 36967 32969
rect 36909 32929 36921 32963
rect 36955 32960 36967 32963
rect 37274 32960 37280 32972
rect 36955 32932 37280 32960
rect 36955 32929 36967 32932
rect 36909 32923 36967 32929
rect 37274 32920 37280 32932
rect 37332 32920 37338 32972
rect 35253 32895 35311 32901
rect 35253 32892 35265 32895
rect 34900 32864 35265 32892
rect 35253 32861 35265 32864
rect 35299 32892 35311 32895
rect 35710 32892 35716 32904
rect 35299 32864 35716 32892
rect 35299 32861 35311 32864
rect 35253 32855 35311 32861
rect 35710 32852 35716 32864
rect 35768 32852 35774 32904
rect 35434 32824 35440 32836
rect 34348 32796 35440 32824
rect 35434 32784 35440 32796
rect 35492 32784 35498 32836
rect 18506 32756 18512 32768
rect 17420 32728 18512 32756
rect 18506 32716 18512 32728
rect 18564 32716 18570 32768
rect 18782 32716 18788 32768
rect 18840 32756 18846 32768
rect 19334 32756 19340 32768
rect 18840 32728 19340 32756
rect 18840 32716 18846 32728
rect 19334 32716 19340 32728
rect 19392 32756 19398 32768
rect 19521 32759 19579 32765
rect 19521 32756 19533 32759
rect 19392 32728 19533 32756
rect 19392 32716 19398 32728
rect 19521 32725 19533 32728
rect 19567 32725 19579 32759
rect 21082 32756 21088 32768
rect 21043 32728 21088 32756
rect 19521 32719 19579 32725
rect 21082 32716 21088 32728
rect 21140 32716 21146 32768
rect 23201 32759 23259 32765
rect 23201 32725 23213 32759
rect 23247 32756 23259 32759
rect 23750 32756 23756 32768
rect 23247 32728 23756 32756
rect 23247 32725 23259 32728
rect 23201 32719 23259 32725
rect 23750 32716 23756 32728
rect 23808 32716 23814 32768
rect 24302 32716 24308 32768
rect 24360 32756 24366 32768
rect 25409 32759 25467 32765
rect 25409 32756 25421 32759
rect 24360 32728 25421 32756
rect 24360 32716 24366 32728
rect 25409 32725 25421 32728
rect 25455 32725 25467 32759
rect 25409 32719 25467 32725
rect 27798 32716 27804 32768
rect 27856 32756 27862 32768
rect 27893 32759 27951 32765
rect 27893 32756 27905 32759
rect 27856 32728 27905 32756
rect 27856 32716 27862 32728
rect 27893 32725 27905 32728
rect 27939 32725 27951 32759
rect 27893 32719 27951 32725
rect 27982 32716 27988 32768
rect 28040 32756 28046 32768
rect 28721 32759 28779 32765
rect 28721 32756 28733 32759
rect 28040 32728 28733 32756
rect 28040 32716 28046 32728
rect 28721 32725 28733 32728
rect 28767 32725 28779 32759
rect 28721 32719 28779 32725
rect 35529 32759 35587 32765
rect 35529 32725 35541 32759
rect 35575 32756 35587 32759
rect 35618 32756 35624 32768
rect 35575 32728 35624 32756
rect 35575 32725 35587 32728
rect 35529 32719 35587 32725
rect 35618 32716 35624 32728
rect 35676 32716 35682 32768
rect 1104 32666 38824 32688
rect 1104 32614 4246 32666
rect 4298 32614 4310 32666
rect 4362 32614 4374 32666
rect 4426 32614 4438 32666
rect 4490 32614 34966 32666
rect 35018 32614 35030 32666
rect 35082 32614 35094 32666
rect 35146 32614 35158 32666
rect 35210 32614 38824 32666
rect 1104 32592 38824 32614
rect 6086 32512 6092 32564
rect 6144 32552 6150 32564
rect 7926 32552 7932 32564
rect 6144 32524 7932 32552
rect 6144 32512 6150 32524
rect 7926 32512 7932 32524
rect 7984 32512 7990 32564
rect 8036 32524 13400 32552
rect 8036 32496 8064 32524
rect 2958 32444 2964 32496
rect 3016 32484 3022 32496
rect 3970 32484 3976 32496
rect 3016 32456 3976 32484
rect 3016 32444 3022 32456
rect 3970 32444 3976 32456
rect 4028 32484 4034 32496
rect 7745 32487 7803 32493
rect 7745 32484 7757 32487
rect 4028 32456 4200 32484
rect 4028 32444 4034 32456
rect 3329 32419 3387 32425
rect 3329 32385 3341 32419
rect 3375 32416 3387 32419
rect 4062 32416 4068 32428
rect 3375 32388 4068 32416
rect 3375 32385 3387 32388
rect 3329 32379 3387 32385
rect 4062 32376 4068 32388
rect 4120 32376 4126 32428
rect 4172 32416 4200 32456
rect 5368 32456 7757 32484
rect 4172 32388 4292 32416
rect 1673 32351 1731 32357
rect 1673 32317 1685 32351
rect 1719 32348 1731 32351
rect 1854 32348 1860 32360
rect 1719 32320 1860 32348
rect 1719 32317 1731 32320
rect 1673 32311 1731 32317
rect 1854 32308 1860 32320
rect 1912 32308 1918 32360
rect 2222 32348 2228 32360
rect 2183 32320 2228 32348
rect 2222 32308 2228 32320
rect 2280 32308 2286 32360
rect 2409 32351 2467 32357
rect 2409 32317 2421 32351
rect 2455 32348 2467 32351
rect 2866 32348 2872 32360
rect 2455 32320 2872 32348
rect 2455 32317 2467 32320
rect 2409 32311 2467 32317
rect 2866 32308 2872 32320
rect 2924 32308 2930 32360
rect 3237 32351 3295 32357
rect 3237 32317 3249 32351
rect 3283 32317 3295 32351
rect 3694 32348 3700 32360
rect 3655 32320 3700 32348
rect 3237 32311 3295 32317
rect 3252 32280 3280 32311
rect 3694 32308 3700 32320
rect 3752 32308 3758 32360
rect 3878 32348 3884 32360
rect 3839 32320 3884 32348
rect 3878 32308 3884 32320
rect 3936 32308 3942 32360
rect 4264 32357 4292 32388
rect 4249 32351 4307 32357
rect 4249 32317 4261 32351
rect 4295 32317 4307 32351
rect 4614 32348 4620 32360
rect 4575 32320 4620 32348
rect 4249 32311 4307 32317
rect 4614 32308 4620 32320
rect 4672 32308 4678 32360
rect 5368 32280 5396 32456
rect 7745 32453 7757 32456
rect 7791 32484 7803 32487
rect 8018 32484 8024 32496
rect 7791 32456 8024 32484
rect 7791 32453 7803 32456
rect 7745 32447 7803 32453
rect 8018 32444 8024 32456
rect 8076 32444 8082 32496
rect 12250 32444 12256 32496
rect 12308 32484 12314 32496
rect 12529 32487 12587 32493
rect 12529 32484 12541 32487
rect 12308 32456 12541 32484
rect 12308 32444 12314 32456
rect 12529 32453 12541 32456
rect 12575 32453 12587 32487
rect 12529 32447 12587 32453
rect 5534 32416 5540 32428
rect 5495 32388 5540 32416
rect 5534 32376 5540 32388
rect 5592 32376 5598 32428
rect 6270 32416 6276 32428
rect 6231 32388 6276 32416
rect 6270 32376 6276 32388
rect 6328 32376 6334 32428
rect 8570 32416 8576 32428
rect 7024 32388 8576 32416
rect 5718 32348 5724 32360
rect 5679 32320 5724 32348
rect 5718 32308 5724 32320
rect 5776 32308 5782 32360
rect 7024 32357 7052 32388
rect 8570 32376 8576 32388
rect 8628 32376 8634 32428
rect 8846 32376 8852 32428
rect 8904 32416 8910 32428
rect 13265 32419 13323 32425
rect 13265 32416 13277 32419
rect 8904 32388 9444 32416
rect 8904 32376 8910 32388
rect 5813 32351 5871 32357
rect 5813 32317 5825 32351
rect 5859 32348 5871 32351
rect 7009 32351 7067 32357
rect 7009 32348 7021 32351
rect 5859 32320 7021 32348
rect 5859 32317 5871 32320
rect 5813 32311 5871 32317
rect 7009 32317 7021 32320
rect 7055 32317 7067 32351
rect 8202 32348 8208 32360
rect 8163 32320 8208 32348
rect 7009 32311 7067 32317
rect 8202 32308 8208 32320
rect 8260 32308 8266 32360
rect 8294 32308 8300 32360
rect 8352 32348 8358 32360
rect 8665 32351 8723 32357
rect 8665 32348 8677 32351
rect 8352 32320 8677 32348
rect 8352 32308 8358 32320
rect 8665 32317 8677 32320
rect 8711 32317 8723 32351
rect 8665 32311 8723 32317
rect 8754 32308 8760 32360
rect 8812 32348 8818 32360
rect 9416 32357 9444 32388
rect 10888 32388 13277 32416
rect 10888 32360 10916 32388
rect 13265 32385 13277 32388
rect 13311 32385 13323 32419
rect 13265 32379 13323 32385
rect 9217 32351 9275 32357
rect 9217 32348 9229 32351
rect 8812 32320 9229 32348
rect 8812 32308 8818 32320
rect 9217 32317 9229 32320
rect 9263 32317 9275 32351
rect 9217 32311 9275 32317
rect 9401 32351 9459 32357
rect 9401 32317 9413 32351
rect 9447 32317 9459 32351
rect 9401 32311 9459 32317
rect 10689 32351 10747 32357
rect 10689 32317 10701 32351
rect 10735 32317 10747 32351
rect 10870 32348 10876 32360
rect 10831 32320 10876 32348
rect 10689 32311 10747 32317
rect 3252 32252 5396 32280
rect 5905 32283 5963 32289
rect 5905 32249 5917 32283
rect 5951 32280 5963 32283
rect 5994 32280 6000 32292
rect 5951 32252 6000 32280
rect 5951 32249 5963 32252
rect 5905 32243 5963 32249
rect 5994 32240 6000 32252
rect 6052 32280 6058 32292
rect 7650 32280 7656 32292
rect 6052 32252 7656 32280
rect 6052 32240 6058 32252
rect 7650 32240 7656 32252
rect 7708 32240 7714 32292
rect 8113 32283 8171 32289
rect 8113 32249 8125 32283
rect 8159 32280 8171 32283
rect 8386 32280 8392 32292
rect 8159 32252 8392 32280
rect 8159 32249 8171 32252
rect 8113 32243 8171 32249
rect 8386 32240 8392 32252
rect 8444 32240 8450 32292
rect 9232 32280 9260 32311
rect 9766 32280 9772 32292
rect 9232 32252 9772 32280
rect 9766 32240 9772 32252
rect 9824 32240 9830 32292
rect 10704 32280 10732 32311
rect 10870 32308 10876 32320
rect 10928 32308 10934 32360
rect 11330 32348 11336 32360
rect 11291 32320 11336 32348
rect 11330 32308 11336 32320
rect 11388 32308 11394 32360
rect 11609 32351 11667 32357
rect 11609 32317 11621 32351
rect 11655 32348 11667 32351
rect 12437 32351 12495 32357
rect 12437 32348 12449 32351
rect 11655 32320 12449 32348
rect 11655 32317 11667 32320
rect 11609 32311 11667 32317
rect 12437 32317 12449 32320
rect 12483 32317 12495 32351
rect 12437 32311 12495 32317
rect 12989 32351 13047 32357
rect 12989 32317 13001 32351
rect 13035 32317 13047 32351
rect 13372 32348 13400 32524
rect 15488 32524 17172 32552
rect 14274 32444 14280 32496
rect 14332 32484 14338 32496
rect 14369 32487 14427 32493
rect 14369 32484 14381 32487
rect 14332 32456 14381 32484
rect 14332 32444 14338 32456
rect 14369 32453 14381 32456
rect 14415 32453 14427 32487
rect 14369 32447 14427 32453
rect 14277 32351 14335 32357
rect 14277 32348 14289 32351
rect 13372 32320 14289 32348
rect 12989 32311 13047 32317
rect 14277 32317 14289 32320
rect 14323 32317 14335 32351
rect 14918 32348 14924 32360
rect 14879 32320 14924 32348
rect 14277 32311 14335 32317
rect 11054 32280 11060 32292
rect 10704 32252 11060 32280
rect 11054 32240 11060 32252
rect 11112 32280 11118 32292
rect 13004 32280 13032 32311
rect 14918 32308 14924 32320
rect 14976 32308 14982 32360
rect 15488 32357 15516 32524
rect 17144 32496 17172 32524
rect 17218 32512 17224 32564
rect 17276 32552 17282 32564
rect 18414 32552 18420 32564
rect 17276 32524 18420 32552
rect 17276 32512 17282 32524
rect 18414 32512 18420 32524
rect 18472 32512 18478 32564
rect 28445 32555 28503 32561
rect 28445 32521 28457 32555
rect 28491 32552 28503 32555
rect 32766 32552 32772 32564
rect 28491 32524 32628 32552
rect 32727 32524 32772 32552
rect 28491 32521 28503 32524
rect 28445 32515 28503 32521
rect 16298 32444 16304 32496
rect 16356 32444 16362 32496
rect 17126 32444 17132 32496
rect 17184 32484 17190 32496
rect 20346 32484 20352 32496
rect 17184 32456 19196 32484
rect 20307 32456 20352 32484
rect 17184 32444 17190 32456
rect 16316 32416 16344 32444
rect 15764 32388 16344 32416
rect 15473 32351 15531 32357
rect 15473 32317 15485 32351
rect 15519 32348 15531 32351
rect 15562 32348 15568 32360
rect 15519 32320 15568 32348
rect 15519 32317 15531 32320
rect 15473 32311 15531 32317
rect 15562 32308 15568 32320
rect 15620 32308 15626 32360
rect 15764 32357 15792 32388
rect 16574 32376 16580 32428
rect 16632 32416 16638 32428
rect 17497 32419 17555 32425
rect 17497 32416 17509 32419
rect 16632 32388 17509 32416
rect 16632 32376 16638 32388
rect 17497 32385 17509 32388
rect 17543 32385 17555 32419
rect 17497 32379 17555 32385
rect 18049 32419 18107 32425
rect 18049 32385 18061 32419
rect 18095 32416 18107 32419
rect 18138 32416 18144 32428
rect 18095 32388 18144 32416
rect 18095 32385 18107 32388
rect 18049 32379 18107 32385
rect 15749 32351 15807 32357
rect 15749 32317 15761 32351
rect 15795 32317 15807 32351
rect 15749 32311 15807 32317
rect 16209 32351 16267 32357
rect 16209 32317 16221 32351
rect 16255 32348 16267 32351
rect 16298 32348 16304 32360
rect 16255 32320 16304 32348
rect 16255 32317 16267 32320
rect 16209 32311 16267 32317
rect 16298 32308 16304 32320
rect 16356 32308 16362 32360
rect 16666 32308 16672 32360
rect 16724 32348 16730 32360
rect 16942 32348 16948 32360
rect 16724 32320 16948 32348
rect 16724 32308 16730 32320
rect 16942 32308 16948 32320
rect 17000 32348 17006 32360
rect 17037 32351 17095 32357
rect 17037 32348 17049 32351
rect 17000 32320 17049 32348
rect 17000 32308 17006 32320
rect 17037 32317 17049 32320
rect 17083 32317 17095 32351
rect 17037 32311 17095 32317
rect 16758 32280 16764 32292
rect 11112 32252 13032 32280
rect 16719 32252 16764 32280
rect 11112 32240 11118 32252
rect 16758 32240 16764 32252
rect 16816 32240 16822 32292
rect 17129 32283 17187 32289
rect 17129 32249 17141 32283
rect 17175 32280 17187 32283
rect 17512 32280 17540 32379
rect 18138 32376 18144 32388
rect 18196 32376 18202 32428
rect 18782 32376 18788 32428
rect 18840 32416 18846 32428
rect 19061 32419 19119 32425
rect 19061 32416 19073 32419
rect 18840 32388 19073 32416
rect 18840 32376 18846 32388
rect 19061 32385 19073 32388
rect 19107 32385 19119 32419
rect 19168 32416 19196 32456
rect 20346 32444 20352 32456
rect 20404 32444 20410 32496
rect 21821 32487 21879 32493
rect 21821 32453 21833 32487
rect 21867 32484 21879 32487
rect 22186 32484 22192 32496
rect 21867 32456 22192 32484
rect 21867 32453 21879 32456
rect 21821 32447 21879 32453
rect 22186 32444 22192 32456
rect 22244 32444 22250 32496
rect 24857 32487 24915 32493
rect 24857 32453 24869 32487
rect 24903 32484 24915 32487
rect 25498 32484 25504 32496
rect 24903 32456 25504 32484
rect 24903 32453 24915 32456
rect 24857 32447 24915 32453
rect 25498 32444 25504 32456
rect 25556 32444 25562 32496
rect 28077 32487 28135 32493
rect 28077 32453 28089 32487
rect 28123 32484 28135 32487
rect 30558 32484 30564 32496
rect 28123 32456 30420 32484
rect 30519 32456 30564 32484
rect 28123 32453 28135 32456
rect 28077 32447 28135 32453
rect 20441 32419 20499 32425
rect 20441 32416 20453 32419
rect 19168 32388 20453 32416
rect 19061 32379 19119 32385
rect 20441 32385 20453 32388
rect 20487 32416 20499 32419
rect 21082 32416 21088 32428
rect 20487 32388 21088 32416
rect 20487 32385 20499 32388
rect 20441 32379 20499 32385
rect 21082 32376 21088 32388
rect 21140 32376 21146 32428
rect 23382 32376 23388 32428
rect 23440 32416 23446 32428
rect 23661 32419 23719 32425
rect 23661 32416 23673 32419
rect 23440 32388 23673 32416
rect 23440 32376 23446 32388
rect 23661 32385 23673 32388
rect 23707 32385 23719 32419
rect 27341 32419 27399 32425
rect 27341 32416 27353 32419
rect 23661 32379 23719 32385
rect 24780 32388 27353 32416
rect 17770 32308 17776 32360
rect 17828 32348 17834 32360
rect 18598 32348 18604 32360
rect 17828 32320 18604 32348
rect 17828 32308 17834 32320
rect 18598 32308 18604 32320
rect 18656 32308 18662 32360
rect 18877 32351 18935 32357
rect 18877 32317 18889 32351
rect 18923 32317 18935 32351
rect 18877 32311 18935 32317
rect 19797 32351 19855 32357
rect 19797 32317 19809 32351
rect 19843 32348 19855 32351
rect 19886 32348 19892 32360
rect 19843 32320 19892 32348
rect 19843 32317 19855 32320
rect 19797 32311 19855 32317
rect 18892 32280 18920 32311
rect 19886 32308 19892 32320
rect 19944 32348 19950 32360
rect 20070 32348 20076 32360
rect 19944 32320 20076 32348
rect 19944 32308 19950 32320
rect 20070 32308 20076 32320
rect 20128 32308 20134 32360
rect 20346 32348 20352 32360
rect 20307 32320 20352 32348
rect 20346 32308 20352 32320
rect 20404 32308 20410 32360
rect 22002 32348 22008 32360
rect 21963 32320 22008 32348
rect 22002 32308 22008 32320
rect 22060 32308 22066 32360
rect 22189 32351 22247 32357
rect 22189 32317 22201 32351
rect 22235 32317 22247 32351
rect 22370 32348 22376 32360
rect 22331 32320 22376 32348
rect 22189 32311 22247 32317
rect 17175 32252 17448 32280
rect 17512 32252 18920 32280
rect 17175 32249 17187 32252
rect 17129 32243 17187 32249
rect 1670 32212 1676 32224
rect 1631 32184 1676 32212
rect 1670 32172 1676 32184
rect 1728 32172 1734 32224
rect 7193 32215 7251 32221
rect 7193 32181 7205 32215
rect 7239 32212 7251 32215
rect 7282 32212 7288 32224
rect 7239 32184 7288 32212
rect 7239 32181 7251 32184
rect 7193 32175 7251 32181
rect 7282 32172 7288 32184
rect 7340 32212 7346 32224
rect 8202 32212 8208 32224
rect 7340 32184 8208 32212
rect 7340 32172 7346 32184
rect 8202 32172 8208 32184
rect 8260 32172 8266 32224
rect 16945 32215 17003 32221
rect 16945 32181 16957 32215
rect 16991 32212 17003 32215
rect 17218 32212 17224 32224
rect 16991 32184 17224 32212
rect 16991 32181 17003 32184
rect 16945 32175 17003 32181
rect 17218 32172 17224 32184
rect 17276 32172 17282 32224
rect 17420 32212 17448 32252
rect 21818 32240 21824 32292
rect 21876 32280 21882 32292
rect 22204 32280 22232 32311
rect 22370 32308 22376 32320
rect 22428 32308 22434 32360
rect 23750 32348 23756 32360
rect 23711 32320 23756 32348
rect 23750 32308 23756 32320
rect 23808 32308 23814 32360
rect 24780 32357 24808 32388
rect 27341 32385 27353 32388
rect 27387 32385 27399 32419
rect 29730 32416 29736 32428
rect 27341 32379 27399 32385
rect 28092 32388 29736 32416
rect 24765 32351 24823 32357
rect 24765 32317 24777 32351
rect 24811 32317 24823 32351
rect 24765 32311 24823 32317
rect 25041 32351 25099 32357
rect 25041 32317 25053 32351
rect 25087 32348 25099 32351
rect 25314 32348 25320 32360
rect 25087 32320 25320 32348
rect 25087 32317 25099 32320
rect 25041 32311 25099 32317
rect 25314 32308 25320 32320
rect 25372 32308 25378 32360
rect 25958 32348 25964 32360
rect 25919 32320 25964 32348
rect 25958 32308 25964 32320
rect 26016 32308 26022 32360
rect 26237 32351 26295 32357
rect 26237 32317 26249 32351
rect 26283 32348 26295 32351
rect 28092 32348 28120 32388
rect 29730 32376 29736 32388
rect 29788 32376 29794 32428
rect 30392 32416 30420 32456
rect 30558 32444 30564 32456
rect 30616 32444 30622 32496
rect 32600 32484 32628 32524
rect 32766 32512 32772 32524
rect 32824 32512 32830 32564
rect 33594 32512 33600 32564
rect 33652 32552 33658 32564
rect 34057 32555 34115 32561
rect 34057 32552 34069 32555
rect 33652 32524 34069 32552
rect 33652 32512 33658 32524
rect 34057 32521 34069 32524
rect 34103 32521 34115 32555
rect 36630 32552 36636 32564
rect 34057 32515 34115 32521
rect 34164 32524 36636 32552
rect 34164 32484 34192 32524
rect 36630 32512 36636 32524
rect 36688 32512 36694 32564
rect 32600 32456 34192 32484
rect 30392 32388 30696 32416
rect 26283 32320 28120 32348
rect 28169 32351 28227 32357
rect 26283 32317 26295 32320
rect 26237 32311 26295 32317
rect 28169 32317 28181 32351
rect 28215 32317 28227 32351
rect 28169 32311 28227 32317
rect 28261 32351 28319 32357
rect 28261 32317 28273 32351
rect 28307 32317 28319 32351
rect 28261 32311 28319 32317
rect 21876 32252 22232 32280
rect 21876 32240 21882 32252
rect 24026 32240 24032 32292
rect 24084 32280 24090 32292
rect 24213 32283 24271 32289
rect 24213 32280 24225 32283
rect 24084 32252 24225 32280
rect 24084 32240 24090 32252
rect 24213 32249 24225 32252
rect 24259 32249 24271 32283
rect 24213 32243 24271 32249
rect 28077 32283 28135 32289
rect 28077 32249 28089 32283
rect 28123 32280 28135 32283
rect 28184 32280 28212 32311
rect 28123 32252 28212 32280
rect 28123 32249 28135 32252
rect 28077 32243 28135 32249
rect 18230 32212 18236 32224
rect 17420 32184 18236 32212
rect 18230 32172 18236 32184
rect 18288 32172 18294 32224
rect 25222 32212 25228 32224
rect 25183 32184 25228 32212
rect 25222 32172 25228 32184
rect 25280 32172 25286 32224
rect 28276 32212 28304 32311
rect 29454 32308 29460 32360
rect 29512 32348 29518 32360
rect 29641 32351 29699 32357
rect 29641 32348 29653 32351
rect 29512 32320 29653 32348
rect 29512 32308 29518 32320
rect 29641 32317 29653 32320
rect 29687 32317 29699 32351
rect 29641 32311 29699 32317
rect 30193 32351 30251 32357
rect 30193 32317 30205 32351
rect 30239 32348 30251 32351
rect 30282 32348 30288 32360
rect 30239 32320 30288 32348
rect 30239 32317 30251 32320
rect 30193 32311 30251 32317
rect 30282 32308 30288 32320
rect 30340 32308 30346 32360
rect 30466 32308 30472 32360
rect 30524 32348 30530 32360
rect 30668 32348 30696 32388
rect 30742 32376 30748 32428
rect 30800 32416 30806 32428
rect 31481 32419 31539 32425
rect 31481 32416 31493 32419
rect 30800 32388 31493 32416
rect 30800 32376 30806 32388
rect 31481 32385 31493 32388
rect 31527 32385 31539 32419
rect 31481 32379 31539 32385
rect 34790 32376 34796 32428
rect 34848 32416 34854 32428
rect 35805 32419 35863 32425
rect 35805 32416 35817 32419
rect 34848 32388 35817 32416
rect 34848 32376 34854 32388
rect 35805 32385 35817 32388
rect 35851 32385 35863 32419
rect 38102 32416 38108 32428
rect 35805 32379 35863 32385
rect 35912 32388 38108 32416
rect 31018 32348 31024 32360
rect 30524 32320 30569 32348
rect 30668 32320 31024 32348
rect 30524 32308 30530 32320
rect 31018 32308 31024 32320
rect 31076 32308 31082 32360
rect 31202 32348 31208 32360
rect 31163 32320 31208 32348
rect 31202 32308 31208 32320
rect 31260 32308 31266 32360
rect 33965 32351 34023 32357
rect 33965 32317 33977 32351
rect 34011 32348 34023 32351
rect 34882 32348 34888 32360
rect 34011 32320 34888 32348
rect 34011 32317 34023 32320
rect 33965 32311 34023 32317
rect 34882 32308 34888 32320
rect 34940 32308 34946 32360
rect 35250 32308 35256 32360
rect 35308 32348 35314 32360
rect 35529 32351 35587 32357
rect 35529 32348 35541 32351
rect 35308 32320 35541 32348
rect 35308 32308 35314 32320
rect 35529 32317 35541 32320
rect 35575 32317 35587 32351
rect 35912 32348 35940 32388
rect 38102 32376 38108 32388
rect 38160 32376 38166 32428
rect 35529 32311 35587 32317
rect 35636 32320 35940 32348
rect 37645 32351 37703 32357
rect 30926 32240 30932 32292
rect 30984 32280 30990 32292
rect 31220 32280 31248 32308
rect 30984 32252 31248 32280
rect 30984 32240 30990 32252
rect 33410 32240 33416 32292
rect 33468 32280 33474 32292
rect 33781 32283 33839 32289
rect 33781 32280 33793 32283
rect 33468 32252 33793 32280
rect 33468 32240 33474 32252
rect 33781 32249 33793 32252
rect 33827 32249 33839 32283
rect 33781 32243 33839 32249
rect 35636 32212 35664 32320
rect 37645 32317 37657 32351
rect 37691 32348 37703 32351
rect 37918 32348 37924 32360
rect 37691 32320 37924 32348
rect 37691 32317 37703 32320
rect 37645 32311 37703 32317
rect 37918 32308 37924 32320
rect 37976 32308 37982 32360
rect 28276 32184 35664 32212
rect 35802 32172 35808 32224
rect 35860 32212 35866 32224
rect 36909 32215 36967 32221
rect 36909 32212 36921 32215
rect 35860 32184 36921 32212
rect 35860 32172 35866 32184
rect 36909 32181 36921 32184
rect 36955 32181 36967 32215
rect 36909 32175 36967 32181
rect 37550 32172 37556 32224
rect 37608 32212 37614 32224
rect 37737 32215 37795 32221
rect 37737 32212 37749 32215
rect 37608 32184 37749 32212
rect 37608 32172 37614 32184
rect 37737 32181 37749 32184
rect 37783 32181 37795 32215
rect 37737 32175 37795 32181
rect 1104 32122 38824 32144
rect 1104 32070 19606 32122
rect 19658 32070 19670 32122
rect 19722 32070 19734 32122
rect 19786 32070 19798 32122
rect 19850 32070 38824 32122
rect 1104 32048 38824 32070
rect 7098 31968 7104 32020
rect 7156 32008 7162 32020
rect 8846 32008 8852 32020
rect 7156 31980 8852 32008
rect 7156 31968 7162 31980
rect 8846 31968 8852 31980
rect 8904 31968 8910 32020
rect 9214 32008 9220 32020
rect 9175 31980 9220 32008
rect 9214 31968 9220 31980
rect 9272 31968 9278 32020
rect 15381 32011 15439 32017
rect 15381 31977 15393 32011
rect 15427 32008 15439 32011
rect 15838 32008 15844 32020
rect 15427 31980 15844 32008
rect 15427 31977 15439 31980
rect 15381 31971 15439 31977
rect 15838 31968 15844 31980
rect 15896 31968 15902 32020
rect 20070 32008 20076 32020
rect 17972 31980 20076 32008
rect 3053 31943 3111 31949
rect 3053 31909 3065 31943
rect 3099 31940 3111 31943
rect 3234 31940 3240 31952
rect 3099 31912 3240 31940
rect 3099 31909 3111 31912
rect 3053 31903 3111 31909
rect 3234 31900 3240 31912
rect 3292 31900 3298 31952
rect 4430 31900 4436 31952
rect 4488 31940 4494 31952
rect 5074 31940 5080 31952
rect 4488 31912 5080 31940
rect 4488 31900 4494 31912
rect 5074 31900 5080 31912
rect 5132 31900 5138 31952
rect 6822 31940 6828 31952
rect 6783 31912 6828 31940
rect 6822 31900 6828 31912
rect 6880 31900 6886 31952
rect 7484 31912 15516 31940
rect 1670 31872 1676 31884
rect 1631 31844 1676 31872
rect 1670 31832 1676 31844
rect 1728 31832 1734 31884
rect 4617 31875 4675 31881
rect 4617 31841 4629 31875
rect 4663 31872 4675 31875
rect 4982 31872 4988 31884
rect 4663 31844 4988 31872
rect 4663 31841 4675 31844
rect 4617 31835 4675 31841
rect 4982 31832 4988 31844
rect 5040 31832 5046 31884
rect 6840 31872 6868 31900
rect 7285 31875 7343 31881
rect 7285 31872 7297 31875
rect 6840 31844 7297 31872
rect 7285 31841 7297 31844
rect 7331 31841 7343 31875
rect 7285 31835 7343 31841
rect 1394 31804 1400 31816
rect 1355 31776 1400 31804
rect 1394 31764 1400 31776
rect 1452 31764 1458 31816
rect 4430 31764 4436 31816
rect 4488 31764 4494 31816
rect 5166 31764 5172 31816
rect 5224 31804 5230 31816
rect 5445 31807 5503 31813
rect 5224 31776 5269 31804
rect 5224 31764 5230 31776
rect 5445 31773 5457 31807
rect 5491 31804 5503 31807
rect 5534 31804 5540 31816
rect 5491 31776 5540 31804
rect 5491 31773 5503 31776
rect 5445 31767 5503 31773
rect 5534 31764 5540 31776
rect 5592 31764 5598 31816
rect 4448 31677 4476 31764
rect 6454 31696 6460 31748
rect 6512 31736 6518 31748
rect 7484 31736 7512 31912
rect 7650 31872 7656 31884
rect 7611 31844 7656 31872
rect 7650 31832 7656 31844
rect 7708 31832 7714 31884
rect 8110 31872 8116 31884
rect 8071 31844 8116 31872
rect 8110 31832 8116 31844
rect 8168 31832 8174 31884
rect 8202 31832 8208 31884
rect 8260 31872 8266 31884
rect 8573 31875 8631 31881
rect 8573 31872 8585 31875
rect 8260 31844 8585 31872
rect 8260 31832 8266 31844
rect 8573 31841 8585 31844
rect 8619 31841 8631 31875
rect 8573 31835 8631 31841
rect 8846 31832 8852 31884
rect 8904 31872 8910 31884
rect 9401 31875 9459 31881
rect 9401 31872 9413 31875
rect 8904 31844 9413 31872
rect 8904 31832 8910 31844
rect 9401 31841 9413 31844
rect 9447 31841 9459 31875
rect 9401 31835 9459 31841
rect 9582 31832 9588 31884
rect 9640 31872 9646 31884
rect 9677 31875 9735 31881
rect 9677 31872 9689 31875
rect 9640 31844 9689 31872
rect 9640 31832 9646 31844
rect 9677 31841 9689 31844
rect 9723 31841 9735 31875
rect 9677 31835 9735 31841
rect 9861 31875 9919 31881
rect 9861 31841 9873 31875
rect 9907 31841 9919 31875
rect 9861 31835 9919 31841
rect 9953 31875 10011 31881
rect 9953 31841 9965 31875
rect 9999 31872 10011 31875
rect 10870 31872 10876 31884
rect 9999 31844 10876 31872
rect 9999 31841 10011 31844
rect 9953 31835 10011 31841
rect 7926 31764 7932 31816
rect 7984 31804 7990 31816
rect 9876 31804 9904 31835
rect 10870 31832 10876 31844
rect 10928 31832 10934 31884
rect 11238 31872 11244 31884
rect 11199 31844 11244 31872
rect 11238 31832 11244 31844
rect 11296 31832 11302 31884
rect 11793 31875 11851 31881
rect 11793 31841 11805 31875
rect 11839 31841 11851 31875
rect 11793 31835 11851 31841
rect 12621 31875 12679 31881
rect 12621 31841 12633 31875
rect 12667 31872 12679 31875
rect 14274 31872 14280 31884
rect 12667 31844 12756 31872
rect 14235 31844 14280 31872
rect 12667 31841 12679 31844
rect 12621 31835 12679 31841
rect 7984 31776 9904 31804
rect 7984 31764 7990 31776
rect 6512 31708 7512 31736
rect 11333 31739 11391 31745
rect 6512 31696 6518 31708
rect 11333 31705 11345 31739
rect 11379 31736 11391 31739
rect 11422 31736 11428 31748
rect 11379 31708 11428 31736
rect 11379 31705 11391 31708
rect 11333 31699 11391 31705
rect 11422 31696 11428 31708
rect 11480 31696 11486 31748
rect 4433 31671 4491 31677
rect 4433 31637 4445 31671
rect 4479 31637 4491 31671
rect 4433 31631 4491 31637
rect 5810 31628 5816 31680
rect 5868 31668 5874 31680
rect 7377 31671 7435 31677
rect 7377 31668 7389 31671
rect 5868 31640 7389 31668
rect 5868 31628 5874 31640
rect 7377 31637 7389 31640
rect 7423 31637 7435 31671
rect 7377 31631 7435 31637
rect 9950 31628 9956 31680
rect 10008 31668 10014 31680
rect 10137 31671 10195 31677
rect 10137 31668 10149 31671
rect 10008 31640 10149 31668
rect 10008 31628 10014 31640
rect 10137 31637 10149 31640
rect 10183 31637 10195 31671
rect 10137 31631 10195 31637
rect 10778 31628 10784 31680
rect 10836 31668 10842 31680
rect 11808 31668 11836 31835
rect 12728 31816 12756 31844
rect 14274 31832 14280 31844
rect 14332 31832 14338 31884
rect 14366 31832 14372 31884
rect 14424 31872 14430 31884
rect 15488 31881 15516 31912
rect 16758 31900 16764 31952
rect 16816 31940 16822 31952
rect 17972 31949 18000 31980
rect 20070 31968 20076 31980
rect 20128 31968 20134 32020
rect 20622 32008 20628 32020
rect 20180 31980 20628 32008
rect 17957 31943 18015 31949
rect 17957 31940 17969 31943
rect 16816 31912 17969 31940
rect 16816 31900 16822 31912
rect 17957 31909 17969 31912
rect 18003 31909 18015 31943
rect 18322 31940 18328 31952
rect 18283 31912 18328 31940
rect 17957 31903 18015 31909
rect 18322 31900 18328 31912
rect 18380 31900 18386 31952
rect 18506 31900 18512 31952
rect 18564 31940 18570 31952
rect 18693 31943 18751 31949
rect 18693 31940 18705 31943
rect 18564 31912 18705 31940
rect 18564 31900 18570 31912
rect 18693 31909 18705 31912
rect 18739 31909 18751 31943
rect 20180 31940 20208 31980
rect 20622 31968 20628 31980
rect 20680 31968 20686 32020
rect 23201 32011 23259 32017
rect 23201 31977 23213 32011
rect 23247 32008 23259 32011
rect 23382 32008 23388 32020
rect 23247 31980 23388 32008
rect 23247 31977 23259 31980
rect 23201 31971 23259 31977
rect 23382 31968 23388 31980
rect 23440 31968 23446 32020
rect 29270 32008 29276 32020
rect 23676 31980 29276 32008
rect 20346 31940 20352 31952
rect 18693 31903 18751 31909
rect 19904 31912 20208 31940
rect 20307 31912 20352 31940
rect 14553 31875 14611 31881
rect 14553 31872 14565 31875
rect 14424 31844 14565 31872
rect 14424 31832 14430 31844
rect 14553 31841 14565 31844
rect 14599 31841 14611 31875
rect 14553 31835 14611 31841
rect 15473 31875 15531 31881
rect 15473 31841 15485 31875
rect 15519 31841 15531 31875
rect 15473 31835 15531 31841
rect 15562 31832 15568 31884
rect 15620 31872 15626 31884
rect 15841 31875 15899 31881
rect 15841 31872 15853 31875
rect 15620 31844 15853 31872
rect 15620 31832 15626 31844
rect 15841 31841 15853 31844
rect 15887 31841 15899 31875
rect 16574 31872 16580 31884
rect 15841 31835 15899 31841
rect 15948 31844 16580 31872
rect 12066 31804 12072 31816
rect 12027 31776 12072 31804
rect 12066 31764 12072 31776
rect 12124 31764 12130 31816
rect 12710 31764 12716 31816
rect 12768 31764 12774 31816
rect 13725 31807 13783 31813
rect 13725 31773 13737 31807
rect 13771 31804 13783 31807
rect 13814 31804 13820 31816
rect 13771 31776 13820 31804
rect 13771 31773 13783 31776
rect 13725 31767 13783 31773
rect 13814 31764 13820 31776
rect 13872 31764 13878 31816
rect 14737 31807 14795 31813
rect 14737 31773 14749 31807
rect 14783 31804 14795 31807
rect 14918 31804 14924 31816
rect 14783 31776 14924 31804
rect 14783 31773 14795 31776
rect 14737 31767 14795 31773
rect 14918 31764 14924 31776
rect 14976 31804 14982 31816
rect 15948 31804 15976 31844
rect 16574 31832 16580 31844
rect 16632 31832 16638 31884
rect 16850 31872 16856 31884
rect 16811 31844 16856 31872
rect 16850 31832 16856 31844
rect 16908 31832 16914 31884
rect 17586 31832 17592 31884
rect 17644 31872 17650 31884
rect 18141 31875 18199 31881
rect 18141 31872 18153 31875
rect 17644 31844 18153 31872
rect 17644 31832 17650 31844
rect 18141 31841 18153 31844
rect 18187 31841 18199 31875
rect 18141 31835 18199 31841
rect 18230 31832 18236 31884
rect 18288 31872 18294 31884
rect 19904 31881 19932 31912
rect 20346 31900 20352 31912
rect 20404 31900 20410 31952
rect 20456 31912 21956 31940
rect 19889 31875 19947 31881
rect 19889 31872 19901 31875
rect 18288 31844 19901 31872
rect 18288 31832 18294 31844
rect 19889 31841 19901 31844
rect 19935 31841 19947 31875
rect 20070 31872 20076 31884
rect 20031 31844 20076 31872
rect 19889 31835 19947 31841
rect 20070 31832 20076 31844
rect 20128 31832 20134 31884
rect 16206 31804 16212 31816
rect 14976 31776 15976 31804
rect 16167 31776 16212 31804
rect 14976 31764 14982 31776
rect 16206 31764 16212 31776
rect 16264 31764 16270 31816
rect 18322 31764 18328 31816
rect 18380 31764 18386 31816
rect 18598 31764 18604 31816
rect 18656 31804 18662 31816
rect 20456 31804 20484 31912
rect 21818 31872 21824 31884
rect 21779 31844 21824 31872
rect 21818 31832 21824 31844
rect 21876 31832 21882 31884
rect 21928 31872 21956 31912
rect 22002 31900 22008 31952
rect 22060 31940 22066 31952
rect 22373 31943 22431 31949
rect 22373 31940 22385 31943
rect 22060 31912 22385 31940
rect 22060 31900 22066 31912
rect 22373 31909 22385 31912
rect 22419 31909 22431 31943
rect 22373 31903 22431 31909
rect 22189 31875 22247 31881
rect 22189 31872 22201 31875
rect 21928 31844 22201 31872
rect 22189 31841 22201 31844
rect 22235 31841 22247 31875
rect 22189 31835 22247 31841
rect 23017 31875 23075 31881
rect 23017 31841 23029 31875
rect 23063 31872 23075 31875
rect 23198 31872 23204 31884
rect 23063 31844 23204 31872
rect 23063 31841 23075 31844
rect 23017 31835 23075 31841
rect 23198 31832 23204 31844
rect 23256 31872 23262 31884
rect 23676 31872 23704 31980
rect 29270 31968 29276 31980
rect 29328 31968 29334 32020
rect 29454 32008 29460 32020
rect 29415 31980 29460 32008
rect 29454 31968 29460 31980
rect 29512 31968 29518 32020
rect 29730 31968 29736 32020
rect 29788 32008 29794 32020
rect 29788 31980 34560 32008
rect 29788 31968 29794 31980
rect 32585 31943 32643 31949
rect 32585 31909 32597 31943
rect 32631 31940 32643 31943
rect 33410 31940 33416 31952
rect 32631 31912 33416 31940
rect 32631 31909 32643 31912
rect 32585 31903 32643 31909
rect 33410 31900 33416 31912
rect 33468 31900 33474 31952
rect 34532 31940 34560 31980
rect 34882 31968 34888 32020
rect 34940 32008 34946 32020
rect 34977 32011 35035 32017
rect 34977 32008 34989 32011
rect 34940 31980 34989 32008
rect 34940 31968 34946 31980
rect 34977 31977 34989 31980
rect 35023 31977 35035 32011
rect 34977 31971 35035 31977
rect 36265 31943 36323 31949
rect 36265 31940 36277 31943
rect 34532 31912 36277 31940
rect 36265 31909 36277 31912
rect 36311 31909 36323 31943
rect 36265 31903 36323 31909
rect 23256 31844 23704 31872
rect 23753 31875 23811 31881
rect 23256 31832 23262 31844
rect 23753 31841 23765 31875
rect 23799 31872 23811 31875
rect 23842 31872 23848 31884
rect 23799 31844 23848 31872
rect 23799 31841 23811 31844
rect 23753 31835 23811 31841
rect 23842 31832 23848 31844
rect 23900 31832 23906 31884
rect 24026 31872 24032 31884
rect 23987 31844 24032 31872
rect 24026 31832 24032 31844
rect 24084 31832 24090 31884
rect 24854 31832 24860 31884
rect 24912 31872 24918 31884
rect 26881 31875 26939 31881
rect 26881 31872 26893 31875
rect 24912 31844 26893 31872
rect 24912 31832 24918 31844
rect 26881 31841 26893 31844
rect 26927 31841 26939 31875
rect 26881 31835 26939 31841
rect 27433 31875 27491 31881
rect 27433 31841 27445 31875
rect 27479 31872 27491 31875
rect 27982 31872 27988 31884
rect 27479 31844 27988 31872
rect 27479 31841 27491 31844
rect 27433 31835 27491 31841
rect 27982 31832 27988 31844
rect 28040 31832 28046 31884
rect 28350 31872 28356 31884
rect 28311 31844 28356 31872
rect 28350 31832 28356 31844
rect 28408 31832 28414 31884
rect 30650 31872 30656 31884
rect 30611 31844 30656 31872
rect 30650 31832 30656 31844
rect 30708 31832 30714 31884
rect 31205 31875 31263 31881
rect 31205 31841 31217 31875
rect 31251 31872 31263 31875
rect 32490 31872 32496 31884
rect 31251 31844 32496 31872
rect 31251 31841 31263 31844
rect 31205 31835 31263 31841
rect 32490 31832 32496 31844
rect 32548 31832 32554 31884
rect 32766 31872 32772 31884
rect 32727 31844 32772 31872
rect 32766 31832 32772 31844
rect 32824 31832 32830 31884
rect 33594 31872 33600 31884
rect 33555 31844 33600 31872
rect 33594 31832 33600 31844
rect 33652 31832 33658 31884
rect 33962 31872 33968 31884
rect 33704 31844 33968 31872
rect 18656 31776 20484 31804
rect 21453 31807 21511 31813
rect 18656 31764 18662 31776
rect 21453 31773 21465 31807
rect 21499 31804 21511 31807
rect 22370 31804 22376 31816
rect 21499 31776 22376 31804
rect 21499 31773 21511 31776
rect 21453 31767 21511 31773
rect 22370 31764 22376 31776
rect 22428 31764 22434 31816
rect 25314 31804 25320 31816
rect 25275 31776 25320 31804
rect 25314 31764 25320 31776
rect 25372 31764 25378 31816
rect 26602 31804 26608 31816
rect 26563 31776 26608 31804
rect 26602 31764 26608 31776
rect 26660 31764 26666 31816
rect 27706 31764 27712 31816
rect 27764 31804 27770 31816
rect 28077 31807 28135 31813
rect 28077 31804 28089 31807
rect 27764 31776 28089 31804
rect 27764 31764 27770 31776
rect 28077 31773 28089 31776
rect 28123 31773 28135 31807
rect 28077 31767 28135 31773
rect 31481 31807 31539 31813
rect 31481 31773 31493 31807
rect 31527 31804 31539 31807
rect 31754 31804 31760 31816
rect 31527 31776 31760 31804
rect 31527 31773 31539 31776
rect 31481 31767 31539 31773
rect 31754 31764 31760 31776
rect 31812 31804 31818 31816
rect 32030 31804 32036 31816
rect 31812 31776 32036 31804
rect 31812 31764 31818 31776
rect 32030 31764 32036 31776
rect 32088 31764 32094 31816
rect 33137 31807 33195 31813
rect 33137 31773 33149 31807
rect 33183 31804 33195 31807
rect 33704 31804 33732 31844
rect 33962 31832 33968 31844
rect 34020 31832 34026 31884
rect 35802 31872 35808 31884
rect 35763 31844 35808 31872
rect 35802 31832 35808 31844
rect 35860 31832 35866 31884
rect 36722 31872 36728 31884
rect 36683 31844 36728 31872
rect 36722 31832 36728 31844
rect 36780 31832 36786 31884
rect 37458 31832 37464 31884
rect 37516 31872 37522 31884
rect 37737 31875 37795 31881
rect 37737 31872 37749 31875
rect 37516 31844 37749 31872
rect 37516 31832 37522 31844
rect 37737 31841 37749 31844
rect 37783 31841 37795 31875
rect 37737 31835 37795 31841
rect 33870 31804 33876 31816
rect 33183 31776 33732 31804
rect 33831 31776 33876 31804
rect 33183 31773 33195 31776
rect 33137 31767 33195 31773
rect 33870 31764 33876 31776
rect 33928 31764 33934 31816
rect 35710 31804 35716 31816
rect 35671 31776 35716 31804
rect 35710 31764 35716 31776
rect 35768 31764 35774 31816
rect 37274 31764 37280 31816
rect 37332 31804 37338 31816
rect 37829 31807 37887 31813
rect 37829 31804 37841 31807
rect 37332 31776 37841 31804
rect 37332 31764 37338 31776
rect 37829 31773 37841 31776
rect 37875 31773 37887 31807
rect 37829 31767 37887 31773
rect 18340 31736 18368 31764
rect 19150 31736 19156 31748
rect 18340 31708 19156 31736
rect 19150 31696 19156 31708
rect 19208 31696 19214 31748
rect 20346 31696 20352 31748
rect 20404 31736 20410 31748
rect 20806 31736 20812 31748
rect 20404 31708 20812 31736
rect 20404 31696 20410 31708
rect 20806 31696 20812 31708
rect 20864 31696 20870 31748
rect 27246 31696 27252 31748
rect 27304 31736 27310 31748
rect 27341 31739 27399 31745
rect 27341 31736 27353 31739
rect 27304 31708 27353 31736
rect 27304 31696 27310 31708
rect 27341 31705 27353 31708
rect 27387 31705 27399 31739
rect 30742 31736 30748 31748
rect 30703 31708 30748 31736
rect 27341 31699 27399 31705
rect 30742 31696 30748 31708
rect 30800 31696 30806 31748
rect 12526 31668 12532 31680
rect 10836 31640 12532 31668
rect 10836 31628 10842 31640
rect 12526 31628 12532 31640
rect 12584 31668 12590 31680
rect 12713 31671 12771 31677
rect 12713 31668 12725 31671
rect 12584 31640 12725 31668
rect 12584 31628 12590 31640
rect 12713 31637 12725 31640
rect 12759 31637 12771 31671
rect 12713 31631 12771 31637
rect 16666 31628 16672 31680
rect 16724 31668 16730 31680
rect 17037 31671 17095 31677
rect 17037 31668 17049 31671
rect 16724 31640 17049 31668
rect 16724 31628 16730 31640
rect 17037 31637 17049 31640
rect 17083 31668 17095 31671
rect 17586 31668 17592 31680
rect 17083 31640 17592 31668
rect 17083 31637 17095 31640
rect 17037 31631 17095 31637
rect 17586 31628 17592 31640
rect 17644 31628 17650 31680
rect 36817 31671 36875 31677
rect 36817 31637 36829 31671
rect 36863 31668 36875 31671
rect 36906 31668 36912 31680
rect 36863 31640 36912 31668
rect 36863 31637 36875 31640
rect 36817 31631 36875 31637
rect 36906 31628 36912 31640
rect 36964 31628 36970 31680
rect 1104 31578 38824 31600
rect 1104 31526 4246 31578
rect 4298 31526 4310 31578
rect 4362 31526 4374 31578
rect 4426 31526 4438 31578
rect 4490 31526 34966 31578
rect 35018 31526 35030 31578
rect 35082 31526 35094 31578
rect 35146 31526 35158 31578
rect 35210 31526 38824 31578
rect 1104 31504 38824 31526
rect 3510 31464 3516 31476
rect 1504 31436 3516 31464
rect 1504 31260 1532 31436
rect 3510 31424 3516 31436
rect 3568 31464 3574 31476
rect 3970 31464 3976 31476
rect 3568 31436 3976 31464
rect 3568 31424 3574 31436
rect 3970 31424 3976 31436
rect 4028 31464 4034 31476
rect 4028 31436 4200 31464
rect 4028 31424 4034 31436
rect 2866 31396 2872 31408
rect 1596 31368 2452 31396
rect 2827 31368 2872 31396
rect 1596 31337 1624 31368
rect 1581 31331 1639 31337
rect 1581 31297 1593 31331
rect 1627 31297 1639 31331
rect 1581 31291 1639 31297
rect 2222 31288 2228 31340
rect 2280 31328 2286 31340
rect 2317 31331 2375 31337
rect 2317 31328 2329 31331
rect 2280 31300 2329 31328
rect 2280 31288 2286 31300
rect 2317 31297 2329 31300
rect 2363 31297 2375 31331
rect 2424 31328 2452 31368
rect 2866 31356 2872 31368
rect 2924 31356 2930 31408
rect 2774 31328 2780 31340
rect 2424 31300 2780 31328
rect 2317 31291 2375 31297
rect 2774 31288 2780 31300
rect 2832 31328 2838 31340
rect 3326 31328 3332 31340
rect 2832 31300 3332 31328
rect 2832 31288 2838 31300
rect 3326 31288 3332 31300
rect 3384 31288 3390 31340
rect 1765 31263 1823 31269
rect 1765 31260 1777 31263
rect 1504 31232 1777 31260
rect 1765 31229 1777 31232
rect 1811 31229 1823 31263
rect 1765 31223 1823 31229
rect 1857 31263 1915 31269
rect 1857 31229 1869 31263
rect 1903 31260 1915 31263
rect 2130 31260 2136 31272
rect 1903 31232 2136 31260
rect 1903 31229 1915 31232
rect 1857 31223 1915 31229
rect 2130 31220 2136 31232
rect 2188 31220 2194 31272
rect 3053 31263 3111 31269
rect 3053 31260 3065 31263
rect 2240 31232 3065 31260
rect 1949 31195 2007 31201
rect 1949 31161 1961 31195
rect 1995 31192 2007 31195
rect 2240 31192 2268 31232
rect 3053 31229 3065 31232
rect 3099 31260 3111 31263
rect 3234 31260 3240 31272
rect 3099 31232 3240 31260
rect 3099 31229 3111 31232
rect 3053 31223 3111 31229
rect 3234 31220 3240 31232
rect 3292 31220 3298 31272
rect 3513 31263 3571 31269
rect 3513 31229 3525 31263
rect 3559 31260 3571 31263
rect 3694 31260 3700 31272
rect 3559 31232 3700 31260
rect 3559 31229 3571 31232
rect 3513 31223 3571 31229
rect 3694 31220 3700 31232
rect 3752 31220 3758 31272
rect 3878 31260 3884 31272
rect 3839 31232 3884 31260
rect 3878 31220 3884 31232
rect 3936 31220 3942 31272
rect 4172 31269 4200 31436
rect 7098 31424 7104 31476
rect 7156 31464 7162 31476
rect 7285 31467 7343 31473
rect 7285 31464 7297 31467
rect 7156 31436 7297 31464
rect 7156 31424 7162 31436
rect 7285 31433 7297 31436
rect 7331 31433 7343 31467
rect 7285 31427 7343 31433
rect 9401 31467 9459 31473
rect 9401 31433 9413 31467
rect 9447 31464 9459 31467
rect 9766 31464 9772 31476
rect 9447 31436 9772 31464
rect 9447 31433 9459 31436
rect 9401 31427 9459 31433
rect 9766 31424 9772 31436
rect 9824 31424 9830 31476
rect 15749 31467 15807 31473
rect 15749 31464 15761 31467
rect 13464 31436 15761 31464
rect 5626 31396 5632 31408
rect 5587 31368 5632 31396
rect 5626 31356 5632 31368
rect 5684 31356 5690 31408
rect 11238 31356 11244 31408
rect 11296 31396 11302 31408
rect 11425 31399 11483 31405
rect 11425 31396 11437 31399
rect 11296 31368 11437 31396
rect 11296 31356 11302 31368
rect 11425 31365 11437 31368
rect 11471 31365 11483 31399
rect 11425 31359 11483 31365
rect 7374 31288 7380 31340
rect 7432 31328 7438 31340
rect 7837 31331 7895 31337
rect 7837 31328 7849 31331
rect 7432 31300 7849 31328
rect 7432 31288 7438 31300
rect 7837 31297 7849 31300
rect 7883 31297 7895 31331
rect 10778 31328 10784 31340
rect 10739 31300 10784 31328
rect 7837 31291 7895 31297
rect 10778 31288 10784 31300
rect 10836 31288 10842 31340
rect 4157 31263 4215 31269
rect 4157 31229 4169 31263
rect 4203 31229 4215 31263
rect 4430 31260 4436 31272
rect 4391 31232 4436 31260
rect 4157 31223 4215 31229
rect 4430 31220 4436 31232
rect 4488 31220 4494 31272
rect 5810 31260 5816 31272
rect 5771 31232 5816 31260
rect 5810 31220 5816 31232
rect 5868 31220 5874 31272
rect 6178 31260 6184 31272
rect 6139 31232 6184 31260
rect 6178 31220 6184 31232
rect 6236 31220 6242 31272
rect 7006 31220 7012 31272
rect 7064 31260 7070 31272
rect 7193 31263 7251 31269
rect 7193 31260 7205 31263
rect 7064 31232 7205 31260
rect 7064 31220 7070 31232
rect 7193 31229 7205 31232
rect 7239 31229 7251 31263
rect 8110 31260 8116 31272
rect 8071 31232 8116 31260
rect 7193 31223 7251 31229
rect 8110 31220 8116 31232
rect 8168 31220 8174 31272
rect 9950 31260 9956 31272
rect 9911 31232 9956 31260
rect 9950 31220 9956 31232
rect 10008 31220 10014 31272
rect 11149 31263 11207 31269
rect 11149 31229 11161 31263
rect 11195 31229 11207 31263
rect 11149 31223 11207 31229
rect 1995 31164 2268 31192
rect 1995 31161 2007 31164
rect 1949 31155 2007 31161
rect 10042 31124 10048 31136
rect 10003 31096 10048 31124
rect 10042 31084 10048 31096
rect 10100 31084 10106 31136
rect 11164 31124 11192 31223
rect 11330 31220 11336 31272
rect 11388 31260 11394 31272
rect 11425 31263 11483 31269
rect 11425 31260 11437 31263
rect 11388 31232 11437 31260
rect 11388 31220 11394 31232
rect 11425 31229 11437 31232
rect 11471 31229 11483 31263
rect 11425 31223 11483 31229
rect 12437 31263 12495 31269
rect 12437 31229 12449 31263
rect 12483 31260 12495 31263
rect 13078 31260 13084 31272
rect 12483 31232 13084 31260
rect 12483 31229 12495 31232
rect 12437 31223 12495 31229
rect 13078 31220 13084 31232
rect 13136 31260 13142 31272
rect 13464 31260 13492 31436
rect 15749 31433 15761 31436
rect 15795 31433 15807 31467
rect 23014 31464 23020 31476
rect 22975 31436 23020 31464
rect 15749 31427 15807 31433
rect 23014 31424 23020 31436
rect 23072 31424 23078 31476
rect 25958 31424 25964 31476
rect 26016 31464 26022 31476
rect 26421 31467 26479 31473
rect 26421 31464 26433 31467
rect 26016 31436 26433 31464
rect 26016 31424 26022 31436
rect 26421 31433 26433 31436
rect 26467 31464 26479 31467
rect 27706 31464 27712 31476
rect 26467 31436 27712 31464
rect 26467 31433 26479 31436
rect 26421 31427 26479 31433
rect 27706 31424 27712 31436
rect 27764 31424 27770 31476
rect 20254 31356 20260 31408
rect 20312 31396 20318 31408
rect 20438 31396 20444 31408
rect 20312 31368 20444 31396
rect 20312 31356 20318 31368
rect 20438 31356 20444 31368
rect 20496 31356 20502 31408
rect 21818 31356 21824 31408
rect 21876 31396 21882 31408
rect 22005 31399 22063 31405
rect 22005 31396 22017 31399
rect 21876 31368 22017 31396
rect 21876 31356 21882 31368
rect 22005 31365 22017 31368
rect 22051 31365 22063 31399
rect 25222 31396 25228 31408
rect 22005 31359 22063 31365
rect 24044 31368 25228 31396
rect 13814 31328 13820 31340
rect 13775 31300 13820 31328
rect 13814 31288 13820 31300
rect 13872 31288 13878 31340
rect 16850 31288 16856 31340
rect 16908 31288 16914 31340
rect 18417 31331 18475 31337
rect 18417 31297 18429 31331
rect 18463 31328 18475 31331
rect 20162 31328 20168 31340
rect 18463 31300 20168 31328
rect 18463 31297 18475 31300
rect 18417 31291 18475 31297
rect 20162 31288 20168 31300
rect 20220 31288 20226 31340
rect 20272 31300 21772 31328
rect 13136 31232 13492 31260
rect 13541 31263 13599 31269
rect 13136 31220 13142 31232
rect 13541 31229 13553 31263
rect 13587 31260 13599 31263
rect 15286 31260 15292 31272
rect 13587 31232 15292 31260
rect 13587 31229 13599 31232
rect 13541 31223 13599 31229
rect 15286 31220 15292 31232
rect 15344 31220 15350 31272
rect 15657 31263 15715 31269
rect 15657 31229 15669 31263
rect 15703 31229 15715 31263
rect 16298 31260 16304 31272
rect 16259 31232 16304 31260
rect 15657 31223 15715 31229
rect 15194 31192 15200 31204
rect 15155 31164 15200 31192
rect 15194 31152 15200 31164
rect 15252 31152 15258 31204
rect 12066 31124 12072 31136
rect 11164 31096 12072 31124
rect 12066 31084 12072 31096
rect 12124 31124 12130 31136
rect 12621 31127 12679 31133
rect 12621 31124 12633 31127
rect 12124 31096 12633 31124
rect 12124 31084 12130 31096
rect 12621 31093 12633 31096
rect 12667 31124 12679 31127
rect 12894 31124 12900 31136
rect 12667 31096 12900 31124
rect 12667 31093 12679 31096
rect 12621 31087 12679 31093
rect 12894 31084 12900 31096
rect 12952 31084 12958 31136
rect 14642 31084 14648 31136
rect 14700 31124 14706 31136
rect 15672 31124 15700 31223
rect 16298 31220 16304 31232
rect 16356 31220 16362 31272
rect 16669 31263 16727 31269
rect 16669 31229 16681 31263
rect 16715 31260 16727 31263
rect 16868 31260 16896 31288
rect 16945 31263 17003 31269
rect 16945 31260 16957 31263
rect 16715 31232 16804 31260
rect 16868 31232 16957 31260
rect 16715 31229 16727 31232
rect 16669 31223 16727 31229
rect 16776 31136 16804 31232
rect 16945 31229 16957 31232
rect 16991 31229 17003 31263
rect 16945 31223 17003 31229
rect 18325 31263 18383 31269
rect 18325 31229 18337 31263
rect 18371 31260 18383 31263
rect 18598 31260 18604 31272
rect 18371 31232 18604 31260
rect 18371 31229 18383 31232
rect 18325 31223 18383 31229
rect 18598 31220 18604 31232
rect 18656 31220 18662 31272
rect 18782 31260 18788 31272
rect 18743 31232 18788 31260
rect 18782 31220 18788 31232
rect 18840 31220 18846 31272
rect 19613 31263 19671 31269
rect 19613 31229 19625 31263
rect 19659 31229 19671 31263
rect 19613 31223 19671 31229
rect 19628 31192 19656 31223
rect 19978 31220 19984 31272
rect 20036 31260 20042 31272
rect 20073 31263 20131 31269
rect 20073 31260 20085 31263
rect 20036 31232 20085 31260
rect 20036 31220 20042 31232
rect 20073 31229 20085 31232
rect 20119 31260 20131 31263
rect 20272 31260 20300 31300
rect 20119 31232 20300 31260
rect 20349 31263 20407 31269
rect 20119 31229 20131 31232
rect 20073 31223 20131 31229
rect 20349 31229 20361 31263
rect 20395 31229 20407 31263
rect 20349 31223 20407 31229
rect 20625 31263 20683 31269
rect 20625 31229 20637 31263
rect 20671 31260 20683 31263
rect 20990 31260 20996 31272
rect 20671 31232 20996 31260
rect 20671 31229 20683 31232
rect 20625 31223 20683 31229
rect 20254 31192 20260 31204
rect 19628 31164 20260 31192
rect 20254 31152 20260 31164
rect 20312 31152 20318 31204
rect 20364 31192 20392 31223
rect 20990 31220 20996 31232
rect 21048 31220 21054 31272
rect 21542 31260 21548 31272
rect 21503 31232 21548 31260
rect 21542 31220 21548 31232
rect 21600 31220 21606 31272
rect 21744 31269 21772 31300
rect 21729 31263 21787 31269
rect 21729 31229 21741 31263
rect 21775 31229 21787 31263
rect 21729 31223 21787 31229
rect 22097 31263 22155 31269
rect 22097 31229 22109 31263
rect 22143 31229 22155 31263
rect 22830 31260 22836 31272
rect 22791 31232 22836 31260
rect 22097 31223 22155 31229
rect 20806 31192 20812 31204
rect 20364 31164 20812 31192
rect 20806 31152 20812 31164
rect 20864 31152 20870 31204
rect 21008 31192 21036 31220
rect 22112 31192 22140 31223
rect 22830 31220 22836 31232
rect 22888 31260 22894 31272
rect 23198 31260 23204 31272
rect 22888 31232 23204 31260
rect 22888 31220 22894 31232
rect 23198 31220 23204 31232
rect 23256 31220 23262 31272
rect 24044 31269 24072 31368
rect 25222 31356 25228 31368
rect 25280 31356 25286 31408
rect 32490 31356 32496 31408
rect 32548 31396 32554 31408
rect 33965 31399 34023 31405
rect 33965 31396 33977 31399
rect 32548 31368 33977 31396
rect 32548 31356 32554 31368
rect 33965 31365 33977 31368
rect 34011 31365 34023 31399
rect 33965 31359 34023 31365
rect 24121 31331 24179 31337
rect 24121 31297 24133 31331
rect 24167 31328 24179 31331
rect 25866 31328 25872 31340
rect 24167 31300 25872 31328
rect 24167 31297 24179 31300
rect 24121 31291 24179 31297
rect 25866 31288 25872 31300
rect 25924 31288 25930 31340
rect 27246 31328 27252 31340
rect 27207 31300 27252 31328
rect 27246 31288 27252 31300
rect 27304 31288 27310 31340
rect 30742 31288 30748 31340
rect 30800 31328 30806 31340
rect 31297 31331 31355 31337
rect 31297 31328 31309 31331
rect 30800 31300 31309 31328
rect 30800 31288 30806 31300
rect 31297 31297 31309 31300
rect 31343 31297 31355 31331
rect 31297 31291 31355 31297
rect 34238 31288 34244 31340
rect 34296 31328 34302 31340
rect 35805 31331 35863 31337
rect 35805 31328 35817 31331
rect 34296 31300 35817 31328
rect 34296 31288 34302 31300
rect 35805 31297 35817 31300
rect 35851 31297 35863 31331
rect 35805 31291 35863 31297
rect 36630 31288 36636 31340
rect 36688 31328 36694 31340
rect 36725 31331 36783 31337
rect 36725 31328 36737 31331
rect 36688 31300 36737 31328
rect 36688 31288 36694 31300
rect 36725 31297 36737 31300
rect 36771 31297 36783 31331
rect 36725 31291 36783 31297
rect 24029 31263 24087 31269
rect 24029 31229 24041 31263
rect 24075 31229 24087 31263
rect 24302 31260 24308 31272
rect 24263 31232 24308 31260
rect 24029 31223 24087 31229
rect 24302 31220 24308 31232
rect 24360 31220 24366 31272
rect 25406 31260 25412 31272
rect 25367 31232 25412 31260
rect 25406 31220 25412 31232
rect 25464 31220 25470 31272
rect 25590 31260 25596 31272
rect 25551 31232 25596 31260
rect 25590 31220 25596 31232
rect 25648 31220 25654 31272
rect 25774 31260 25780 31272
rect 25735 31232 25780 31260
rect 25774 31220 25780 31232
rect 25832 31220 25838 31272
rect 26605 31263 26663 31269
rect 26605 31229 26617 31263
rect 26651 31260 26663 31263
rect 26878 31260 26884 31272
rect 26651 31232 26884 31260
rect 26651 31229 26663 31232
rect 26605 31223 26663 31229
rect 26878 31220 26884 31232
rect 26936 31220 26942 31272
rect 26970 31220 26976 31272
rect 27028 31260 27034 31272
rect 28626 31260 28632 31272
rect 27028 31232 27073 31260
rect 28539 31232 28632 31260
rect 27028 31220 27034 31232
rect 28626 31220 28632 31232
rect 28684 31260 28690 31272
rect 29457 31263 29515 31269
rect 29457 31260 29469 31263
rect 28684 31232 29469 31260
rect 28684 31220 28690 31232
rect 29457 31229 29469 31232
rect 29503 31229 29515 31263
rect 29457 31223 29515 31229
rect 30009 31263 30067 31269
rect 30009 31229 30021 31263
rect 30055 31260 30067 31263
rect 30282 31260 30288 31272
rect 30055 31232 30288 31260
rect 30055 31229 30067 31232
rect 30009 31223 30067 31229
rect 30282 31220 30288 31232
rect 30340 31220 30346 31272
rect 30377 31263 30435 31269
rect 30377 31229 30389 31263
rect 30423 31260 30435 31263
rect 30466 31260 30472 31272
rect 30423 31232 30472 31260
rect 30423 31229 30435 31232
rect 30377 31223 30435 31229
rect 30466 31220 30472 31232
rect 30524 31220 30530 31272
rect 30926 31220 30932 31272
rect 30984 31260 30990 31272
rect 31021 31263 31079 31269
rect 31021 31260 31033 31263
rect 30984 31232 31033 31260
rect 30984 31220 30990 31232
rect 31021 31229 31033 31232
rect 31067 31229 31079 31263
rect 31021 31223 31079 31229
rect 32677 31263 32735 31269
rect 32677 31229 32689 31263
rect 32723 31260 32735 31263
rect 33137 31263 33195 31269
rect 33137 31260 33149 31263
rect 32723 31232 33149 31260
rect 32723 31229 32735 31232
rect 32677 31223 32735 31229
rect 33137 31229 33149 31232
rect 33183 31229 33195 31263
rect 33137 31223 33195 31229
rect 30558 31192 30564 31204
rect 21008 31164 22140 31192
rect 30519 31164 30564 31192
rect 30558 31152 30564 31164
rect 30616 31152 30622 31204
rect 16758 31124 16764 31136
rect 14700 31096 15700 31124
rect 16671 31096 16764 31124
rect 14700 31084 14706 31096
rect 16758 31084 16764 31096
rect 16816 31124 16822 31136
rect 20530 31124 20536 31136
rect 16816 31096 20536 31124
rect 16816 31084 16822 31096
rect 20530 31084 20536 31096
rect 20588 31084 20594 31136
rect 24486 31124 24492 31136
rect 24447 31096 24492 31124
rect 24486 31084 24492 31096
rect 24544 31084 24550 31136
rect 30190 31084 30196 31136
rect 30248 31124 30254 31136
rect 32692 31124 32720 31223
rect 33226 31220 33232 31272
rect 33284 31260 33290 31272
rect 33505 31263 33563 31269
rect 33505 31260 33517 31263
rect 33284 31232 33517 31260
rect 33284 31220 33290 31232
rect 33505 31229 33517 31232
rect 33551 31229 33563 31263
rect 33962 31260 33968 31272
rect 33923 31232 33968 31260
rect 33505 31223 33563 31229
rect 33520 31192 33548 31223
rect 33962 31220 33968 31232
rect 34020 31220 34026 31272
rect 34790 31220 34796 31272
rect 34848 31260 34854 31272
rect 34885 31263 34943 31269
rect 34885 31260 34897 31263
rect 34848 31232 34897 31260
rect 34848 31220 34854 31232
rect 34885 31229 34897 31232
rect 34931 31229 34943 31263
rect 34885 31223 34943 31229
rect 35253 31263 35311 31269
rect 35253 31229 35265 31263
rect 35299 31229 35311 31263
rect 35253 31223 35311 31229
rect 35268 31192 35296 31223
rect 35342 31220 35348 31272
rect 35400 31260 35406 31272
rect 35713 31263 35771 31269
rect 35713 31260 35725 31263
rect 35400 31232 35725 31260
rect 35400 31220 35406 31232
rect 35713 31229 35725 31232
rect 35759 31229 35771 31263
rect 36446 31260 36452 31272
rect 36407 31232 36452 31260
rect 35713 31223 35771 31229
rect 36446 31220 36452 31232
rect 36504 31220 36510 31272
rect 35434 31192 35440 31204
rect 33520 31164 35440 31192
rect 35434 31152 35440 31164
rect 35492 31152 35498 31204
rect 30248 31096 32720 31124
rect 30248 31084 30254 31096
rect 32766 31084 32772 31136
rect 32824 31124 32830 31136
rect 37829 31127 37887 31133
rect 37829 31124 37841 31127
rect 32824 31096 37841 31124
rect 32824 31084 32830 31096
rect 37829 31093 37841 31096
rect 37875 31093 37887 31127
rect 37829 31087 37887 31093
rect 1104 31034 38824 31056
rect 1104 30982 19606 31034
rect 19658 30982 19670 31034
rect 19722 30982 19734 31034
rect 19786 30982 19798 31034
rect 19850 30982 38824 31034
rect 1104 30960 38824 30982
rect 3602 30920 3608 30932
rect 2976 30892 3608 30920
rect 2976 30796 3004 30892
rect 3602 30880 3608 30892
rect 3660 30880 3666 30932
rect 5534 30880 5540 30932
rect 5592 30920 5598 30932
rect 5721 30923 5779 30929
rect 5721 30920 5733 30923
rect 5592 30892 5733 30920
rect 5592 30880 5598 30892
rect 5721 30889 5733 30892
rect 5767 30889 5779 30923
rect 14642 30920 14648 30932
rect 14603 30892 14648 30920
rect 5721 30883 5779 30889
rect 14642 30880 14648 30892
rect 14700 30880 14706 30932
rect 16298 30880 16304 30932
rect 16356 30920 16362 30932
rect 16356 30892 17172 30920
rect 16356 30880 16362 30892
rect 7837 30855 7895 30861
rect 7837 30821 7849 30855
rect 7883 30852 7895 30855
rect 8110 30852 8116 30864
rect 7883 30824 8116 30852
rect 7883 30821 7895 30824
rect 7837 30815 7895 30821
rect 8110 30812 8116 30824
rect 8168 30812 8174 30864
rect 16758 30852 16764 30864
rect 16719 30824 16764 30852
rect 16758 30812 16764 30824
rect 16816 30812 16822 30864
rect 17144 30861 17172 30892
rect 20254 30880 20260 30932
rect 20312 30920 20318 30932
rect 20993 30923 21051 30929
rect 20993 30920 21005 30923
rect 20312 30892 21005 30920
rect 20312 30880 20318 30892
rect 20993 30889 21005 30892
rect 21039 30889 21051 30923
rect 20993 30883 21051 30889
rect 22002 30880 22008 30932
rect 22060 30920 22066 30932
rect 22370 30920 22376 30932
rect 22060 30892 22376 30920
rect 22060 30880 22066 30892
rect 22370 30880 22376 30892
rect 22428 30920 22434 30932
rect 23385 30923 23443 30929
rect 23385 30920 23397 30923
rect 22428 30892 23397 30920
rect 22428 30880 22434 30892
rect 23385 30889 23397 30892
rect 23431 30889 23443 30923
rect 23385 30883 23443 30889
rect 24213 30923 24271 30929
rect 24213 30889 24225 30923
rect 24259 30920 24271 30923
rect 24854 30920 24860 30932
rect 24259 30892 24860 30920
rect 24259 30889 24271 30892
rect 24213 30883 24271 30889
rect 24854 30880 24860 30892
rect 24912 30880 24918 30932
rect 25869 30923 25927 30929
rect 25869 30889 25881 30923
rect 25915 30920 25927 30923
rect 26602 30920 26608 30932
rect 25915 30892 26608 30920
rect 25915 30889 25927 30892
rect 25869 30883 25927 30889
rect 26602 30880 26608 30892
rect 26660 30880 26666 30932
rect 33597 30923 33655 30929
rect 33597 30889 33609 30923
rect 33643 30920 33655 30923
rect 33870 30920 33876 30932
rect 33643 30892 33876 30920
rect 33643 30889 33655 30892
rect 33597 30883 33655 30889
rect 33870 30880 33876 30892
rect 33928 30880 33934 30932
rect 36722 30920 36728 30932
rect 36683 30892 36728 30920
rect 36722 30880 36728 30892
rect 36780 30880 36786 30932
rect 17129 30855 17187 30861
rect 17129 30821 17141 30855
rect 17175 30852 17187 30855
rect 19150 30852 19156 30864
rect 17175 30824 19156 30852
rect 17175 30821 17187 30824
rect 17129 30815 17187 30821
rect 19150 30812 19156 30824
rect 19208 30812 19214 30864
rect 22020 30852 22048 30880
rect 25130 30852 25136 30864
rect 20364 30824 22048 30852
rect 24320 30824 25136 30852
rect 1854 30744 1860 30796
rect 1912 30784 1918 30796
rect 2593 30787 2651 30793
rect 2593 30784 2605 30787
rect 1912 30756 2605 30784
rect 1912 30744 1918 30756
rect 2593 30753 2605 30756
rect 2639 30753 2651 30787
rect 2958 30784 2964 30796
rect 2919 30756 2964 30784
rect 2593 30747 2651 30753
rect 2608 30716 2636 30747
rect 2958 30744 2964 30756
rect 3016 30744 3022 30796
rect 3145 30787 3203 30793
rect 3145 30753 3157 30787
rect 3191 30784 3203 30787
rect 3602 30784 3608 30796
rect 3191 30756 3608 30784
rect 3191 30753 3203 30756
rect 3145 30747 3203 30753
rect 3602 30744 3608 30756
rect 3660 30744 3666 30796
rect 4985 30787 5043 30793
rect 4985 30753 4997 30787
rect 5031 30753 5043 30787
rect 5626 30784 5632 30796
rect 5587 30756 5632 30784
rect 4985 30747 5043 30753
rect 5000 30716 5028 30747
rect 5626 30744 5632 30756
rect 5684 30744 5690 30796
rect 6822 30784 6828 30796
rect 6783 30756 6828 30784
rect 6822 30744 6828 30756
rect 6880 30744 6886 30796
rect 7006 30784 7012 30796
rect 6967 30756 7012 30784
rect 7006 30744 7012 30756
rect 7064 30744 7070 30796
rect 7377 30787 7435 30793
rect 7377 30753 7389 30787
rect 7423 30784 7435 30787
rect 7650 30784 7656 30796
rect 7423 30756 7656 30784
rect 7423 30753 7435 30756
rect 7377 30747 7435 30753
rect 7650 30744 7656 30756
rect 7708 30744 7714 30796
rect 8386 30784 8392 30796
rect 8347 30756 8392 30784
rect 8386 30744 8392 30756
rect 8444 30744 8450 30796
rect 8662 30784 8668 30796
rect 8623 30756 8668 30784
rect 8662 30744 8668 30756
rect 8720 30744 8726 30796
rect 8938 30744 8944 30796
rect 8996 30784 9002 30796
rect 9677 30787 9735 30793
rect 9677 30784 9689 30787
rect 8996 30756 9689 30784
rect 8996 30744 9002 30756
rect 9677 30753 9689 30756
rect 9723 30753 9735 30787
rect 10318 30784 10324 30796
rect 10279 30756 10324 30784
rect 9677 30747 9735 30753
rect 10318 30744 10324 30756
rect 10376 30744 10382 30796
rect 11146 30784 11152 30796
rect 11107 30756 11152 30784
rect 11146 30744 11152 30756
rect 11204 30744 11210 30796
rect 13541 30787 13599 30793
rect 13541 30753 13553 30787
rect 13587 30753 13599 30787
rect 13541 30747 13599 30753
rect 6546 30716 6552 30728
rect 2608 30688 3464 30716
rect 5000 30688 6552 30716
rect 3142 30648 3148 30660
rect 3103 30620 3148 30648
rect 3142 30608 3148 30620
rect 3200 30608 3206 30660
rect 3436 30648 3464 30688
rect 6546 30676 6552 30688
rect 6604 30676 6610 30728
rect 8849 30719 8907 30725
rect 8849 30685 8861 30719
rect 8895 30716 8907 30719
rect 9766 30716 9772 30728
rect 8895 30688 9772 30716
rect 8895 30685 8907 30688
rect 8849 30679 8907 30685
rect 9766 30676 9772 30688
rect 9824 30676 9830 30728
rect 11422 30716 11428 30728
rect 11383 30688 11428 30716
rect 11422 30676 11428 30688
rect 11480 30676 11486 30728
rect 6454 30648 6460 30660
rect 3436 30620 6460 30648
rect 6454 30608 6460 30620
rect 6512 30608 6518 30660
rect 13556 30648 13584 30747
rect 13722 30744 13728 30796
rect 13780 30784 13786 30796
rect 13817 30787 13875 30793
rect 13817 30784 13829 30787
rect 13780 30756 13829 30784
rect 13780 30744 13786 30756
rect 13817 30753 13829 30756
rect 13863 30753 13875 30787
rect 13817 30747 13875 30753
rect 14553 30787 14611 30793
rect 14553 30753 14565 30787
rect 14599 30753 14611 30787
rect 14553 30747 14611 30753
rect 13633 30719 13691 30725
rect 13633 30685 13645 30719
rect 13679 30716 13691 30719
rect 14458 30716 14464 30728
rect 13679 30688 14464 30716
rect 13679 30685 13691 30688
rect 13633 30679 13691 30685
rect 14458 30676 14464 30688
rect 14516 30676 14522 30728
rect 14568 30716 14596 30747
rect 15194 30744 15200 30796
rect 15252 30784 15258 30796
rect 15381 30787 15439 30793
rect 15381 30784 15393 30787
rect 15252 30756 15393 30784
rect 15252 30744 15258 30756
rect 15381 30753 15393 30756
rect 15427 30753 15439 30787
rect 15381 30747 15439 30753
rect 16117 30787 16175 30793
rect 16117 30753 16129 30787
rect 16163 30784 16175 30787
rect 16390 30784 16396 30796
rect 16163 30756 16396 30784
rect 16163 30753 16175 30756
rect 16117 30747 16175 30753
rect 16390 30744 16396 30756
rect 16448 30744 16454 30796
rect 16945 30787 17003 30793
rect 16945 30753 16957 30787
rect 16991 30753 17003 30787
rect 16945 30747 17003 30753
rect 17037 30787 17095 30793
rect 17037 30753 17049 30787
rect 17083 30784 17095 30787
rect 17586 30784 17592 30796
rect 17083 30756 17592 30784
rect 17083 30753 17095 30756
rect 17037 30747 17095 30753
rect 14568 30688 15516 30716
rect 13814 30648 13820 30660
rect 13556 30620 13820 30648
rect 13814 30608 13820 30620
rect 13872 30608 13878 30660
rect 15488 30657 15516 30688
rect 16758 30676 16764 30728
rect 16816 30716 16822 30728
rect 16960 30716 16988 30747
rect 17586 30744 17592 30756
rect 17644 30744 17650 30796
rect 17954 30784 17960 30796
rect 17915 30756 17960 30784
rect 17954 30744 17960 30756
rect 18012 30744 18018 30796
rect 18506 30784 18512 30796
rect 18467 30756 18512 30784
rect 18506 30744 18512 30756
rect 18564 30744 18570 30796
rect 19426 30744 19432 30796
rect 19484 30784 19490 30796
rect 20364 30793 20392 30824
rect 19613 30787 19671 30793
rect 19613 30784 19625 30787
rect 19484 30756 19625 30784
rect 19484 30744 19490 30756
rect 19613 30753 19625 30756
rect 19659 30753 19671 30787
rect 19613 30747 19671 30753
rect 20349 30787 20407 30793
rect 20349 30753 20361 30787
rect 20395 30753 20407 30787
rect 20349 30747 20407 30753
rect 20622 30744 20628 30796
rect 20680 30784 20686 30796
rect 20901 30787 20959 30793
rect 20901 30784 20913 30787
rect 20680 30756 20913 30784
rect 20680 30744 20686 30756
rect 20901 30753 20913 30756
rect 20947 30784 20959 30787
rect 23566 30784 23572 30796
rect 20947 30756 23572 30784
rect 20947 30753 20959 30756
rect 20901 30747 20959 30753
rect 23566 30744 23572 30756
rect 23624 30744 23630 30796
rect 24320 30793 24348 30824
rect 25130 30812 25136 30824
rect 25188 30812 25194 30864
rect 26804 30824 27844 30852
rect 24305 30787 24363 30793
rect 24305 30753 24317 30787
rect 24351 30753 24363 30787
rect 24305 30747 24363 30753
rect 24673 30787 24731 30793
rect 24673 30753 24685 30787
rect 24719 30753 24731 30787
rect 24673 30747 24731 30753
rect 25777 30787 25835 30793
rect 25777 30753 25789 30787
rect 25823 30753 25835 30787
rect 25777 30747 25835 30753
rect 16816 30688 16988 30716
rect 16816 30676 16822 30688
rect 17310 30676 17316 30728
rect 17368 30716 17374 30728
rect 17497 30719 17555 30725
rect 17497 30716 17509 30719
rect 17368 30688 17509 30716
rect 17368 30676 17374 30688
rect 17497 30685 17509 30688
rect 17543 30685 17555 30719
rect 17497 30679 17555 30685
rect 19981 30719 20039 30725
rect 19981 30685 19993 30719
rect 20027 30716 20039 30719
rect 20806 30716 20812 30728
rect 20027 30688 20812 30716
rect 20027 30685 20039 30688
rect 19981 30679 20039 30685
rect 20806 30676 20812 30688
rect 20864 30676 20870 30728
rect 21082 30676 21088 30728
rect 21140 30716 21146 30728
rect 22005 30719 22063 30725
rect 22005 30716 22017 30719
rect 21140 30688 22017 30716
rect 21140 30676 21146 30688
rect 22005 30685 22017 30688
rect 22051 30685 22063 30719
rect 22278 30716 22284 30728
rect 22239 30688 22284 30716
rect 22005 30679 22063 30685
rect 22278 30676 22284 30688
rect 22336 30676 22342 30728
rect 15473 30651 15531 30657
rect 15473 30617 15485 30651
rect 15519 30617 15531 30651
rect 15473 30611 15531 30617
rect 16868 30620 18368 30648
rect 5077 30583 5135 30589
rect 5077 30549 5089 30583
rect 5123 30580 5135 30583
rect 5626 30580 5632 30592
rect 5123 30552 5632 30580
rect 5123 30549 5135 30552
rect 5077 30543 5135 30549
rect 5626 30540 5632 30552
rect 5684 30540 5690 30592
rect 9214 30540 9220 30592
rect 9272 30580 9278 30592
rect 9769 30583 9827 30589
rect 9769 30580 9781 30583
rect 9272 30552 9781 30580
rect 9272 30540 9278 30552
rect 9769 30549 9781 30552
rect 9815 30549 9827 30583
rect 10410 30580 10416 30592
rect 10371 30552 10416 30580
rect 9769 30543 9827 30549
rect 10410 30540 10416 30552
rect 10468 30540 10474 30592
rect 12710 30580 12716 30592
rect 12671 30552 12716 30580
rect 12710 30540 12716 30552
rect 12768 30540 12774 30592
rect 14734 30540 14740 30592
rect 14792 30580 14798 30592
rect 16868 30580 16896 30620
rect 14792 30552 16896 30580
rect 14792 30540 14798 30552
rect 16942 30540 16948 30592
rect 17000 30580 17006 30592
rect 18049 30583 18107 30589
rect 18049 30580 18061 30583
rect 17000 30552 18061 30580
rect 17000 30540 17006 30552
rect 18049 30549 18061 30552
rect 18095 30549 18107 30583
rect 18340 30580 18368 30620
rect 24688 30580 24716 30747
rect 24946 30716 24952 30728
rect 24907 30688 24952 30716
rect 24946 30676 24952 30688
rect 25004 30676 25010 30728
rect 25792 30716 25820 30747
rect 26694 30744 26700 30796
rect 26752 30784 26758 30796
rect 26804 30793 26832 30824
rect 26789 30787 26847 30793
rect 26789 30784 26801 30787
rect 26752 30756 26801 30784
rect 26752 30744 26758 30756
rect 26789 30753 26801 30756
rect 26835 30753 26847 30787
rect 27154 30784 27160 30796
rect 27115 30756 27160 30784
rect 26789 30747 26847 30753
rect 27154 30744 27160 30756
rect 27212 30744 27218 30796
rect 27706 30784 27712 30796
rect 27667 30756 27712 30784
rect 27706 30744 27712 30756
rect 27764 30744 27770 30796
rect 27816 30784 27844 30824
rect 30558 30812 30564 30864
rect 30616 30852 30622 30864
rect 30616 30824 33548 30852
rect 30616 30812 30622 30824
rect 29825 30787 29883 30793
rect 29825 30784 29837 30787
rect 27816 30756 29837 30784
rect 29825 30753 29837 30756
rect 29871 30753 29883 30787
rect 30282 30784 30288 30796
rect 30243 30756 30288 30784
rect 29825 30747 29883 30753
rect 30282 30744 30288 30756
rect 30340 30744 30346 30796
rect 30466 30744 30472 30796
rect 30524 30784 30530 30796
rect 30653 30787 30711 30793
rect 30653 30784 30665 30787
rect 30524 30756 30665 30784
rect 30524 30744 30530 30756
rect 30653 30753 30665 30756
rect 30699 30753 30711 30787
rect 30653 30747 30711 30753
rect 32585 30787 32643 30793
rect 32585 30753 32597 30787
rect 32631 30784 32643 30787
rect 32766 30784 32772 30796
rect 32631 30756 32772 30784
rect 32631 30753 32643 30756
rect 32585 30747 32643 30753
rect 32766 30744 32772 30756
rect 32824 30744 32830 30796
rect 33520 30793 33548 30824
rect 33686 30812 33692 30864
rect 33744 30852 33750 30864
rect 35250 30852 35256 30864
rect 33744 30824 35256 30852
rect 33744 30812 33750 30824
rect 35250 30812 35256 30824
rect 35308 30852 35314 30864
rect 35308 30824 35388 30852
rect 35308 30812 35314 30824
rect 33505 30787 33563 30793
rect 33505 30753 33517 30787
rect 33551 30753 33563 30787
rect 34238 30784 34244 30796
rect 34199 30756 34244 30784
rect 33505 30747 33563 30753
rect 34238 30744 34244 30756
rect 34296 30744 34302 30796
rect 35360 30793 35388 30824
rect 35345 30787 35403 30793
rect 35345 30753 35357 30787
rect 35391 30753 35403 30787
rect 35618 30784 35624 30796
rect 35579 30756 35624 30784
rect 35345 30747 35403 30753
rect 35618 30744 35624 30756
rect 35676 30744 35682 30796
rect 37734 30784 37740 30796
rect 37695 30756 37740 30784
rect 37734 30744 37740 30756
rect 37792 30744 37798 30796
rect 27982 30716 27988 30728
rect 25792 30688 27752 30716
rect 27943 30688 27988 30716
rect 25406 30608 25412 30660
rect 25464 30648 25470 30660
rect 26605 30651 26663 30657
rect 26605 30648 26617 30651
rect 25464 30620 26617 30648
rect 25464 30608 25470 30620
rect 26605 30617 26617 30620
rect 26651 30617 26663 30651
rect 26605 30611 26663 30617
rect 18340 30552 24716 30580
rect 27724 30580 27752 30688
rect 27982 30676 27988 30688
rect 28040 30676 28046 30728
rect 31018 30676 31024 30728
rect 31076 30716 31082 30728
rect 32493 30719 32551 30725
rect 32493 30716 32505 30719
rect 31076 30688 32505 30716
rect 31076 30676 31082 30688
rect 32493 30685 32505 30688
rect 32539 30685 32551 30719
rect 32493 30679 32551 30685
rect 33045 30719 33103 30725
rect 33045 30685 33057 30719
rect 33091 30716 33103 30719
rect 33134 30716 33140 30728
rect 33091 30688 33140 30716
rect 33091 30685 33103 30688
rect 33045 30679 33103 30685
rect 33134 30676 33140 30688
rect 33192 30676 33198 30728
rect 34333 30719 34391 30725
rect 34333 30685 34345 30719
rect 34379 30685 34391 30719
rect 34333 30679 34391 30685
rect 30650 30648 30656 30660
rect 30611 30620 30656 30648
rect 30650 30608 30656 30620
rect 30708 30608 30714 30660
rect 32030 30608 32036 30660
rect 32088 30648 32094 30660
rect 34348 30648 34376 30679
rect 32088 30620 34376 30648
rect 32088 30608 32094 30620
rect 27890 30580 27896 30592
rect 27724 30552 27896 30580
rect 18049 30543 18107 30549
rect 27890 30540 27896 30552
rect 27948 30540 27954 30592
rect 29270 30580 29276 30592
rect 29231 30552 29276 30580
rect 29270 30540 29276 30552
rect 29328 30540 29334 30592
rect 36814 30540 36820 30592
rect 36872 30580 36878 30592
rect 37829 30583 37887 30589
rect 37829 30580 37841 30583
rect 36872 30552 37841 30580
rect 36872 30540 36878 30552
rect 37829 30549 37841 30552
rect 37875 30549 37887 30583
rect 37829 30543 37887 30549
rect 1104 30490 38824 30512
rect 1104 30438 4246 30490
rect 4298 30438 4310 30490
rect 4362 30438 4374 30490
rect 4426 30438 4438 30490
rect 4490 30438 34966 30490
rect 35018 30438 35030 30490
rect 35082 30438 35094 30490
rect 35146 30438 35158 30490
rect 35210 30438 38824 30490
rect 1104 30416 38824 30438
rect 6181 30379 6239 30385
rect 6181 30345 6193 30379
rect 6227 30376 6239 30379
rect 6638 30376 6644 30388
rect 6227 30348 6644 30376
rect 6227 30345 6239 30348
rect 6181 30339 6239 30345
rect 6638 30336 6644 30348
rect 6696 30336 6702 30388
rect 13725 30379 13783 30385
rect 13725 30345 13737 30379
rect 13771 30376 13783 30379
rect 13814 30376 13820 30388
rect 13771 30348 13820 30376
rect 13771 30345 13783 30348
rect 13725 30339 13783 30345
rect 13814 30336 13820 30348
rect 13872 30336 13878 30388
rect 26694 30376 26700 30388
rect 26655 30348 26700 30376
rect 26694 30336 26700 30348
rect 26752 30336 26758 30388
rect 30926 30336 30932 30388
rect 30984 30376 30990 30388
rect 31386 30376 31392 30388
rect 30984 30348 31392 30376
rect 30984 30336 30990 30348
rect 31386 30336 31392 30348
rect 31444 30376 31450 30388
rect 32677 30379 32735 30385
rect 32677 30376 32689 30379
rect 31444 30348 32689 30376
rect 31444 30336 31450 30348
rect 32677 30345 32689 30348
rect 32723 30376 32735 30379
rect 33594 30376 33600 30388
rect 32723 30348 33600 30376
rect 32723 30345 32735 30348
rect 32677 30339 32735 30345
rect 33594 30336 33600 30348
rect 33652 30336 33658 30388
rect 3602 30308 3608 30320
rect 3563 30280 3608 30308
rect 3602 30268 3608 30280
rect 3660 30268 3666 30320
rect 8846 30268 8852 30320
rect 8904 30308 8910 30320
rect 9125 30311 9183 30317
rect 9125 30308 9137 30311
rect 8904 30280 9137 30308
rect 8904 30268 8910 30280
rect 9125 30277 9137 30280
rect 9171 30277 9183 30311
rect 9125 30271 9183 30277
rect 12618 30268 12624 30320
rect 12676 30308 12682 30320
rect 17034 30308 17040 30320
rect 12676 30280 17040 30308
rect 12676 30268 12682 30280
rect 17034 30268 17040 30280
rect 17092 30268 17098 30320
rect 21542 30268 21548 30320
rect 21600 30308 21606 30320
rect 23937 30311 23995 30317
rect 21600 30280 23336 30308
rect 21600 30268 21606 30280
rect 1673 30243 1731 30249
rect 1673 30209 1685 30243
rect 1719 30240 1731 30243
rect 3142 30240 3148 30252
rect 1719 30212 3148 30240
rect 1719 30209 1731 30212
rect 1673 30203 1731 30209
rect 3142 30200 3148 30212
rect 3200 30200 3206 30252
rect 3694 30200 3700 30252
rect 3752 30240 3758 30252
rect 4341 30243 4399 30249
rect 4341 30240 4353 30243
rect 3752 30212 4353 30240
rect 3752 30200 3758 30212
rect 4341 30209 4353 30212
rect 4387 30240 4399 30243
rect 4706 30240 4712 30252
rect 4387 30212 4712 30240
rect 4387 30209 4399 30212
rect 4341 30203 4399 30209
rect 4706 30200 4712 30212
rect 4764 30200 4770 30252
rect 7282 30240 7288 30252
rect 5276 30212 7288 30240
rect 1394 30172 1400 30184
rect 1307 30144 1400 30172
rect 1394 30132 1400 30144
rect 1452 30172 1458 30184
rect 3510 30172 3516 30184
rect 1452 30144 3372 30172
rect 3471 30144 3516 30172
rect 1452 30132 1458 30144
rect 3344 30104 3372 30144
rect 3510 30132 3516 30144
rect 3568 30132 3574 30184
rect 3878 30132 3884 30184
rect 3936 30172 3942 30184
rect 5276 30181 5304 30212
rect 7282 30200 7288 30212
rect 7340 30240 7346 30252
rect 9677 30243 9735 30249
rect 7340 30212 9352 30240
rect 7340 30200 7346 30212
rect 4065 30175 4123 30181
rect 4065 30172 4077 30175
rect 3936 30144 4077 30172
rect 3936 30132 3942 30144
rect 4065 30141 4077 30144
rect 4111 30141 4123 30175
rect 4065 30135 4123 30141
rect 5261 30175 5319 30181
rect 5261 30141 5273 30175
rect 5307 30141 5319 30175
rect 5261 30135 5319 30141
rect 5353 30175 5411 30181
rect 5353 30141 5365 30175
rect 5399 30172 5411 30175
rect 5902 30172 5908 30184
rect 5399 30144 5908 30172
rect 5399 30141 5411 30144
rect 5353 30135 5411 30141
rect 5902 30132 5908 30144
rect 5960 30132 5966 30184
rect 5997 30175 6055 30181
rect 5997 30141 6009 30175
rect 6043 30141 6055 30175
rect 7006 30172 7012 30184
rect 6967 30144 7012 30172
rect 5997 30135 6055 30141
rect 5166 30104 5172 30116
rect 3344 30076 5172 30104
rect 5166 30064 5172 30076
rect 5224 30064 5230 30116
rect 6012 30104 6040 30135
rect 7006 30132 7012 30144
rect 7064 30132 7070 30184
rect 7374 30172 7380 30184
rect 7335 30144 7380 30172
rect 7374 30132 7380 30144
rect 7432 30132 7438 30184
rect 7558 30132 7564 30184
rect 7616 30172 7622 30184
rect 7653 30175 7711 30181
rect 7653 30172 7665 30175
rect 7616 30144 7665 30172
rect 7616 30132 7622 30144
rect 7653 30141 7665 30144
rect 7699 30141 7711 30175
rect 8386 30172 8392 30184
rect 7653 30135 7711 30141
rect 7760 30144 8064 30172
rect 8347 30144 8392 30172
rect 7760 30104 7788 30144
rect 7926 30104 7932 30116
rect 5276 30076 7788 30104
rect 7887 30076 7932 30104
rect 5276 30048 5304 30076
rect 7926 30064 7932 30076
rect 7984 30064 7990 30116
rect 8036 30104 8064 30144
rect 8386 30132 8392 30144
rect 8444 30132 8450 30184
rect 9324 30181 9352 30212
rect 9677 30209 9689 30243
rect 9723 30240 9735 30243
rect 10042 30240 10048 30252
rect 9723 30212 10048 30240
rect 9723 30209 9735 30212
rect 9677 30203 9735 30209
rect 10042 30200 10048 30212
rect 10100 30200 10106 30252
rect 12986 30240 12992 30252
rect 10152 30212 12992 30240
rect 9309 30175 9367 30181
rect 9309 30141 9321 30175
rect 9355 30141 9367 30175
rect 9309 30135 9367 30141
rect 9398 30132 9404 30184
rect 9456 30172 9462 30184
rect 10152 30172 10180 30212
rect 12986 30200 12992 30212
rect 13044 30200 13050 30252
rect 14642 30240 14648 30252
rect 13740 30212 14648 30240
rect 11517 30175 11575 30181
rect 11517 30172 11529 30175
rect 9456 30144 10180 30172
rect 11072 30144 11529 30172
rect 9456 30132 9462 30144
rect 11072 30116 11100 30144
rect 11517 30141 11529 30144
rect 11563 30141 11575 30175
rect 11517 30135 11575 30141
rect 11606 30132 11612 30184
rect 11664 30132 11670 30184
rect 12526 30172 12532 30184
rect 12487 30144 12532 30172
rect 12526 30132 12532 30144
rect 12584 30132 12590 30184
rect 12894 30172 12900 30184
rect 12855 30144 12900 30172
rect 12894 30132 12900 30144
rect 12952 30132 12958 30184
rect 13740 30181 13768 30212
rect 14642 30200 14648 30212
rect 14700 30200 14706 30252
rect 16485 30243 16543 30249
rect 16485 30209 16497 30243
rect 16531 30240 16543 30243
rect 18506 30240 18512 30252
rect 16531 30212 18512 30240
rect 16531 30209 16543 30212
rect 16485 30203 16543 30209
rect 18506 30200 18512 30212
rect 18564 30200 18570 30252
rect 20806 30240 20812 30252
rect 20767 30212 20812 30240
rect 20806 30200 20812 30212
rect 20864 30200 20870 30252
rect 22005 30243 22063 30249
rect 22005 30209 22017 30243
rect 22051 30240 22063 30243
rect 23308 30240 23336 30280
rect 23937 30277 23949 30311
rect 23983 30308 23995 30311
rect 24946 30308 24952 30320
rect 23983 30280 24952 30308
rect 23983 30277 23995 30280
rect 23937 30271 23995 30277
rect 24946 30268 24952 30280
rect 25004 30268 25010 30320
rect 27982 30268 27988 30320
rect 28040 30308 28046 30320
rect 28261 30311 28319 30317
rect 28261 30308 28273 30311
rect 28040 30280 28273 30308
rect 28040 30268 28046 30280
rect 28261 30277 28273 30280
rect 28307 30277 28319 30311
rect 29362 30308 29368 30320
rect 29323 30280 29368 30308
rect 28261 30271 28319 30277
rect 29362 30268 29368 30280
rect 29420 30268 29426 30320
rect 35250 30268 35256 30320
rect 35308 30308 35314 30320
rect 35308 30280 36492 30308
rect 35308 30268 35314 30280
rect 36464 30252 36492 30280
rect 24489 30243 24547 30249
rect 24489 30240 24501 30243
rect 22051 30212 22784 30240
rect 23308 30212 24501 30240
rect 22051 30209 22063 30212
rect 22005 30203 22063 30209
rect 13725 30175 13783 30181
rect 13725 30141 13737 30175
rect 13771 30141 13783 30175
rect 14274 30172 14280 30184
rect 14235 30144 14280 30172
rect 13725 30135 13783 30141
rect 14274 30132 14280 30144
rect 14332 30132 14338 30184
rect 14366 30132 14372 30184
rect 14424 30172 14430 30184
rect 14461 30175 14519 30181
rect 14461 30172 14473 30175
rect 14424 30144 14473 30172
rect 14424 30132 14430 30144
rect 14461 30141 14473 30144
rect 14507 30141 14519 30175
rect 14461 30135 14519 30141
rect 9122 30104 9128 30116
rect 8036 30076 9128 30104
rect 9122 30064 9128 30076
rect 9180 30064 9186 30116
rect 11054 30104 11060 30116
rect 11015 30076 11060 30104
rect 11054 30064 11060 30076
rect 11112 30064 11118 30116
rect 11624 30104 11652 30132
rect 14476 30104 14504 30135
rect 14550 30132 14556 30184
rect 14608 30172 14614 30184
rect 14921 30175 14979 30181
rect 14921 30172 14933 30175
rect 14608 30144 14933 30172
rect 14608 30132 14614 30144
rect 14921 30141 14933 30144
rect 14967 30141 14979 30175
rect 14921 30135 14979 30141
rect 15194 30132 15200 30184
rect 15252 30172 15258 30184
rect 15565 30175 15623 30181
rect 15565 30172 15577 30175
rect 15252 30144 15577 30172
rect 15252 30132 15258 30144
rect 15565 30141 15577 30144
rect 15611 30141 15623 30175
rect 17034 30172 17040 30184
rect 16995 30144 17040 30172
rect 15565 30135 15623 30141
rect 17034 30132 17040 30144
rect 17092 30132 17098 30184
rect 17310 30172 17316 30184
rect 17271 30144 17316 30172
rect 17310 30132 17316 30144
rect 17368 30132 17374 30184
rect 17497 30175 17555 30181
rect 17497 30141 17509 30175
rect 17543 30141 17555 30175
rect 17497 30135 17555 30141
rect 17402 30104 17408 30116
rect 11624 30076 14412 30104
rect 14476 30076 17408 30104
rect 2866 29996 2872 30048
rect 2924 30036 2930 30048
rect 2961 30039 3019 30045
rect 2961 30036 2973 30039
rect 2924 30008 2973 30036
rect 2924 29996 2930 30008
rect 2961 30005 2973 30008
rect 3007 30005 3019 30039
rect 2961 29999 3019 30005
rect 4982 29996 4988 30048
rect 5040 30036 5046 30048
rect 5077 30039 5135 30045
rect 5077 30036 5089 30039
rect 5040 30008 5089 30036
rect 5040 29996 5046 30008
rect 5077 30005 5089 30008
rect 5123 30005 5135 30039
rect 5077 29999 5135 30005
rect 5258 29996 5264 30048
rect 5316 29996 5322 30048
rect 5442 30036 5448 30048
rect 5403 30008 5448 30036
rect 5442 29996 5448 30008
rect 5500 29996 5506 30048
rect 7190 29996 7196 30048
rect 7248 30036 7254 30048
rect 8573 30039 8631 30045
rect 8573 30036 8585 30039
rect 7248 30008 8585 30036
rect 7248 29996 7254 30008
rect 8573 30005 8585 30008
rect 8619 30005 8631 30039
rect 11606 30036 11612 30048
rect 11567 30008 11612 30036
rect 8573 29999 8631 30005
rect 11606 29996 11612 30008
rect 11664 29996 11670 30048
rect 12342 29996 12348 30048
rect 12400 30036 12406 30048
rect 12529 30039 12587 30045
rect 12529 30036 12541 30039
rect 12400 30008 12541 30036
rect 12400 29996 12406 30008
rect 12529 30005 12541 30008
rect 12575 30005 12587 30039
rect 14384 30036 14412 30076
rect 17402 30064 17408 30076
rect 17460 30064 17466 30116
rect 15654 30036 15660 30048
rect 14384 30008 15660 30036
rect 12529 29999 12587 30005
rect 15654 29996 15660 30008
rect 15712 29996 15718 30048
rect 15746 29996 15752 30048
rect 15804 30036 15810 30048
rect 15804 30008 15849 30036
rect 15804 29996 15810 30008
rect 16022 29996 16028 30048
rect 16080 30036 16086 30048
rect 16390 30036 16396 30048
rect 16080 30008 16396 30036
rect 16080 29996 16086 30008
rect 16390 29996 16396 30008
rect 16448 30036 16454 30048
rect 17512 30036 17540 30135
rect 18046 30132 18052 30184
rect 18104 30172 18110 30184
rect 18233 30175 18291 30181
rect 18233 30172 18245 30175
rect 18104 30144 18245 30172
rect 18104 30132 18110 30144
rect 18233 30141 18245 30144
rect 18279 30141 18291 30175
rect 18233 30135 18291 30141
rect 18969 30175 19027 30181
rect 18969 30141 18981 30175
rect 19015 30141 19027 30175
rect 18969 30135 19027 30141
rect 19245 30175 19303 30181
rect 19245 30141 19257 30175
rect 19291 30172 19303 30175
rect 19426 30172 19432 30184
rect 19291 30144 19432 30172
rect 19291 30141 19303 30144
rect 19245 30135 19303 30141
rect 18984 30104 19012 30135
rect 19426 30132 19432 30144
rect 19484 30132 19490 30184
rect 19978 30172 19984 30184
rect 19939 30144 19984 30172
rect 19978 30132 19984 30144
rect 20036 30172 20042 30184
rect 20622 30172 20628 30184
rect 20036 30144 20628 30172
rect 20036 30132 20042 30144
rect 20622 30132 20628 30144
rect 20680 30132 20686 30184
rect 20717 30175 20775 30181
rect 20717 30141 20729 30175
rect 20763 30172 20775 30175
rect 20990 30172 20996 30184
rect 20763 30144 20996 30172
rect 20763 30141 20775 30144
rect 20717 30135 20775 30141
rect 20990 30132 20996 30144
rect 21048 30132 21054 30184
rect 22373 30175 22431 30181
rect 22373 30141 22385 30175
rect 22419 30172 22431 30175
rect 22462 30172 22468 30184
rect 22419 30144 22468 30172
rect 22419 30141 22431 30144
rect 22373 30135 22431 30141
rect 22462 30132 22468 30144
rect 22520 30132 22526 30184
rect 22646 30172 22652 30184
rect 22607 30144 22652 30172
rect 22646 30132 22652 30144
rect 22704 30132 22710 30184
rect 22756 30172 22784 30212
rect 24489 30209 24501 30212
rect 24535 30209 24547 30243
rect 25590 30240 25596 30252
rect 25551 30212 25596 30240
rect 24489 30203 24547 30209
rect 25590 30200 25596 30212
rect 25648 30200 25654 30252
rect 33134 30200 33140 30252
rect 33192 30240 33198 30252
rect 36446 30240 36452 30252
rect 33192 30212 36308 30240
rect 36359 30212 36452 30240
rect 33192 30200 33198 30212
rect 23474 30172 23480 30184
rect 22756 30144 23480 30172
rect 23474 30132 23480 30144
rect 23532 30132 23538 30184
rect 23842 30172 23848 30184
rect 23803 30144 23848 30172
rect 23842 30132 23848 30144
rect 23900 30132 23906 30184
rect 24210 30172 24216 30184
rect 24171 30144 24216 30172
rect 24210 30132 24216 30144
rect 24268 30132 24274 30184
rect 25317 30175 25375 30181
rect 25317 30141 25329 30175
rect 25363 30141 25375 30175
rect 25317 30135 25375 30141
rect 19334 30104 19340 30116
rect 18984 30076 19340 30104
rect 19334 30064 19340 30076
rect 19392 30064 19398 30116
rect 22925 30107 22983 30113
rect 22925 30073 22937 30107
rect 22971 30104 22983 30107
rect 25038 30104 25044 30116
rect 22971 30076 25044 30104
rect 22971 30073 22983 30076
rect 22925 30067 22983 30073
rect 25038 30064 25044 30076
rect 25096 30064 25102 30116
rect 16448 30008 17540 30036
rect 18325 30039 18383 30045
rect 16448 29996 16454 30008
rect 18325 30005 18337 30039
rect 18371 30036 18383 30039
rect 18966 30036 18972 30048
rect 18371 30008 18972 30036
rect 18371 30005 18383 30008
rect 18325 29999 18383 30005
rect 18966 29996 18972 30008
rect 19024 29996 19030 30048
rect 19981 30039 20039 30045
rect 19981 30005 19993 30039
rect 20027 30036 20039 30039
rect 20070 30036 20076 30048
rect 20027 30008 20076 30036
rect 20027 30005 20039 30008
rect 19981 29999 20039 30005
rect 20070 29996 20076 30008
rect 20128 29996 20134 30048
rect 25332 30036 25360 30135
rect 27154 30132 27160 30184
rect 27212 30172 27218 30184
rect 27433 30175 27491 30181
rect 27433 30172 27445 30175
rect 27212 30144 27445 30172
rect 27212 30132 27218 30144
rect 27433 30141 27445 30144
rect 27479 30141 27491 30175
rect 27433 30135 27491 30141
rect 27801 30175 27859 30181
rect 27801 30141 27813 30175
rect 27847 30141 27859 30175
rect 27801 30135 27859 30141
rect 28353 30175 28411 30181
rect 28353 30141 28365 30175
rect 28399 30172 28411 30175
rect 28994 30172 29000 30184
rect 28399 30144 29000 30172
rect 28399 30141 28411 30144
rect 28353 30135 28411 30141
rect 26418 30064 26424 30116
rect 26476 30104 26482 30116
rect 27816 30104 27844 30135
rect 28994 30132 29000 30144
rect 29052 30132 29058 30184
rect 29454 30172 29460 30184
rect 29415 30144 29460 30172
rect 29454 30132 29460 30144
rect 29512 30132 29518 30184
rect 29638 30132 29644 30184
rect 29696 30172 29702 30184
rect 29822 30172 29828 30184
rect 29696 30144 29828 30172
rect 29696 30132 29702 30144
rect 29822 30132 29828 30144
rect 29880 30132 29886 30184
rect 30926 30132 30932 30184
rect 30984 30172 30990 30184
rect 31113 30175 31171 30181
rect 31113 30172 31125 30175
rect 30984 30144 31125 30172
rect 30984 30132 30990 30144
rect 31113 30141 31125 30144
rect 31159 30141 31171 30175
rect 31846 30172 31852 30184
rect 31807 30144 31852 30172
rect 31113 30135 31171 30141
rect 31846 30132 31852 30144
rect 31904 30132 31910 30184
rect 32030 30172 32036 30184
rect 31991 30144 32036 30172
rect 32030 30132 32036 30144
rect 32088 30132 32094 30184
rect 32861 30175 32919 30181
rect 32861 30172 32873 30175
rect 32784 30144 32873 30172
rect 26476 30076 27844 30104
rect 26476 30064 26482 30076
rect 32784 30048 32812 30144
rect 32861 30141 32873 30144
rect 32907 30141 32919 30175
rect 32861 30135 32919 30141
rect 32950 30132 32956 30184
rect 33008 30172 33014 30184
rect 33229 30175 33287 30181
rect 33229 30172 33241 30175
rect 33008 30144 33241 30172
rect 33008 30132 33014 30144
rect 33229 30141 33241 30144
rect 33275 30141 33287 30175
rect 33229 30135 33287 30141
rect 33410 30132 33416 30184
rect 33468 30172 33474 30184
rect 33597 30175 33655 30181
rect 33597 30172 33609 30175
rect 33468 30144 33609 30172
rect 33468 30132 33474 30144
rect 33597 30141 33609 30144
rect 33643 30141 33655 30175
rect 33597 30135 33655 30141
rect 34149 30175 34207 30181
rect 34149 30141 34161 30175
rect 34195 30172 34207 30175
rect 34514 30172 34520 30184
rect 34195 30144 34520 30172
rect 34195 30141 34207 30144
rect 34149 30135 34207 30141
rect 34514 30132 34520 30144
rect 34572 30132 34578 30184
rect 35437 30175 35495 30181
rect 35437 30141 35449 30175
rect 35483 30141 35495 30175
rect 35618 30172 35624 30184
rect 35579 30144 35624 30172
rect 35437 30135 35495 30141
rect 34238 30064 34244 30116
rect 34296 30104 34302 30116
rect 34333 30107 34391 30113
rect 34333 30104 34345 30107
rect 34296 30076 34345 30104
rect 34296 30064 34302 30076
rect 34333 30073 34345 30076
rect 34379 30073 34391 30107
rect 35452 30104 35480 30135
rect 35618 30132 35624 30144
rect 35676 30132 35682 30184
rect 35989 30175 36047 30181
rect 35989 30141 36001 30175
rect 36035 30172 36047 30175
rect 36035 30144 36216 30172
rect 36035 30141 36047 30144
rect 35989 30135 36047 30141
rect 35894 30104 35900 30116
rect 35452 30076 35900 30104
rect 34333 30067 34391 30073
rect 35894 30064 35900 30076
rect 35952 30064 35958 30116
rect 26970 30036 26976 30048
rect 25332 30008 26976 30036
rect 26970 29996 26976 30008
rect 27028 30036 27034 30048
rect 27430 30036 27436 30048
rect 27028 30008 27436 30036
rect 27028 29996 27034 30008
rect 27430 29996 27436 30008
rect 27488 29996 27494 30048
rect 31205 30039 31263 30045
rect 31205 30005 31217 30039
rect 31251 30036 31263 30039
rect 31662 30036 31668 30048
rect 31251 30008 31668 30036
rect 31251 30005 31263 30008
rect 31205 29999 31263 30005
rect 31662 29996 31668 30008
rect 31720 29996 31726 30048
rect 32766 30036 32772 30048
rect 32679 30008 32772 30036
rect 32766 29996 32772 30008
rect 32824 30036 32830 30048
rect 34606 30036 34612 30048
rect 32824 30008 34612 30036
rect 32824 29996 32830 30008
rect 34606 29996 34612 30008
rect 34664 29996 34670 30048
rect 36188 30036 36216 30144
rect 36280 30104 36308 30212
rect 36446 30200 36452 30212
rect 36504 30200 36510 30252
rect 36725 30175 36783 30181
rect 36725 30172 36737 30175
rect 36556 30144 36737 30172
rect 36556 30104 36584 30144
rect 36725 30141 36737 30144
rect 36771 30141 36783 30175
rect 36725 30135 36783 30141
rect 37366 30132 37372 30184
rect 37424 30172 37430 30184
rect 37550 30172 37556 30184
rect 37424 30144 37556 30172
rect 37424 30132 37430 30144
rect 37550 30132 37556 30144
rect 37608 30132 37614 30184
rect 36280 30076 36584 30104
rect 37182 30036 37188 30048
rect 36188 30008 37188 30036
rect 37182 29996 37188 30008
rect 37240 29996 37246 30048
rect 37550 29996 37556 30048
rect 37608 30036 37614 30048
rect 37829 30039 37887 30045
rect 37829 30036 37841 30039
rect 37608 30008 37841 30036
rect 37608 29996 37614 30008
rect 37829 30005 37841 30008
rect 37875 30005 37887 30039
rect 37829 29999 37887 30005
rect 1104 29946 38824 29968
rect 1104 29894 19606 29946
rect 19658 29894 19670 29946
rect 19722 29894 19734 29946
rect 19786 29894 19798 29946
rect 19850 29894 38824 29946
rect 1104 29872 38824 29894
rect 3053 29835 3111 29841
rect 3053 29801 3065 29835
rect 3099 29832 3111 29835
rect 3510 29832 3516 29844
rect 3099 29804 3516 29832
rect 3099 29801 3111 29804
rect 3053 29795 3111 29801
rect 3510 29792 3516 29804
rect 3568 29792 3574 29844
rect 3878 29792 3884 29844
rect 3936 29832 3942 29844
rect 4157 29835 4215 29841
rect 4157 29832 4169 29835
rect 3936 29804 4169 29832
rect 3936 29792 3942 29804
rect 4157 29801 4169 29804
rect 4203 29832 4215 29835
rect 4614 29832 4620 29844
rect 4203 29804 4620 29832
rect 4203 29801 4215 29804
rect 4157 29795 4215 29801
rect 4614 29792 4620 29804
rect 4672 29792 4678 29844
rect 4798 29792 4804 29844
rect 4856 29832 4862 29844
rect 5258 29832 5264 29844
rect 4856 29804 5264 29832
rect 4856 29792 4862 29804
rect 5258 29792 5264 29804
rect 5316 29792 5322 29844
rect 12618 29832 12624 29844
rect 9692 29804 12624 29832
rect 5166 29724 5172 29776
rect 5224 29764 5230 29776
rect 5224 29736 5396 29764
rect 5224 29724 5230 29736
rect 2225 29699 2283 29705
rect 2225 29665 2237 29699
rect 2271 29696 2283 29699
rect 2866 29696 2872 29708
rect 2271 29668 2872 29696
rect 2271 29665 2283 29668
rect 2225 29659 2283 29665
rect 2866 29656 2872 29668
rect 2924 29656 2930 29708
rect 4062 29696 4068 29708
rect 4023 29668 4068 29696
rect 4062 29656 4068 29668
rect 4120 29656 4126 29708
rect 4617 29699 4675 29705
rect 4617 29665 4629 29699
rect 4663 29696 4675 29699
rect 5258 29696 5264 29708
rect 4663 29668 5264 29696
rect 4663 29665 4675 29668
rect 4617 29659 4675 29665
rect 5258 29656 5264 29668
rect 5316 29656 5322 29708
rect 5368 29705 5396 29736
rect 7374 29724 7380 29776
rect 7432 29764 7438 29776
rect 7432 29736 8156 29764
rect 7432 29724 7438 29736
rect 5353 29699 5411 29705
rect 5353 29665 5365 29699
rect 5399 29665 5411 29699
rect 5626 29696 5632 29708
rect 5587 29668 5632 29696
rect 5353 29659 5411 29665
rect 5626 29656 5632 29668
rect 5684 29656 5690 29708
rect 6546 29656 6552 29708
rect 6604 29696 6610 29708
rect 7469 29699 7527 29705
rect 7469 29696 7481 29699
rect 6604 29668 7481 29696
rect 6604 29656 6610 29668
rect 7469 29665 7481 29668
rect 7515 29665 7527 29699
rect 7926 29696 7932 29708
rect 7887 29668 7932 29696
rect 7469 29659 7527 29665
rect 7926 29656 7932 29668
rect 7984 29656 7990 29708
rect 8128 29705 8156 29736
rect 8113 29699 8171 29705
rect 8113 29665 8125 29699
rect 8159 29665 8171 29699
rect 8113 29659 8171 29665
rect 8297 29699 8355 29705
rect 8297 29665 8309 29699
rect 8343 29665 8355 29699
rect 8297 29659 8355 29665
rect 7006 29628 7012 29640
rect 6919 29600 7012 29628
rect 7006 29588 7012 29600
rect 7064 29628 7070 29640
rect 8312 29628 8340 29659
rect 8386 29656 8392 29708
rect 8444 29696 8450 29708
rect 9692 29705 9720 29804
rect 12618 29792 12624 29804
rect 12676 29792 12682 29844
rect 13722 29832 13728 29844
rect 13096 29804 13728 29832
rect 11517 29767 11575 29773
rect 11517 29733 11529 29767
rect 11563 29764 11575 29767
rect 13096 29764 13124 29804
rect 13722 29792 13728 29804
rect 13780 29792 13786 29844
rect 14550 29832 14556 29844
rect 13924 29804 14556 29832
rect 11563 29736 13124 29764
rect 11563 29733 11575 29736
rect 11517 29727 11575 29733
rect 8941 29699 8999 29705
rect 8941 29696 8953 29699
rect 8444 29668 8953 29696
rect 8444 29656 8450 29668
rect 8941 29665 8953 29668
rect 8987 29696 8999 29699
rect 9677 29699 9735 29705
rect 9677 29696 9689 29699
rect 8987 29668 9689 29696
rect 8987 29665 8999 29668
rect 8941 29659 8999 29665
rect 9677 29665 9689 29668
rect 9723 29665 9735 29699
rect 9677 29659 9735 29665
rect 10413 29699 10471 29705
rect 10413 29665 10425 29699
rect 10459 29665 10471 29699
rect 12342 29696 12348 29708
rect 12303 29668 12348 29696
rect 10413 29659 10471 29665
rect 7064 29600 8340 29628
rect 7064 29588 7070 29600
rect 9030 29588 9036 29640
rect 9088 29628 9094 29640
rect 10428 29628 10456 29659
rect 12342 29656 12348 29668
rect 12400 29656 12406 29708
rect 12986 29696 12992 29708
rect 12947 29668 12992 29696
rect 12986 29656 12992 29668
rect 13044 29656 13050 29708
rect 13924 29696 13952 29804
rect 14550 29792 14556 29804
rect 14608 29792 14614 29844
rect 15654 29792 15660 29844
rect 15712 29832 15718 29844
rect 21174 29832 21180 29844
rect 15712 29804 21180 29832
rect 15712 29792 15718 29804
rect 21174 29792 21180 29804
rect 21232 29792 21238 29844
rect 25774 29832 25780 29844
rect 21284 29804 25780 29832
rect 17129 29767 17187 29773
rect 17129 29733 17141 29767
rect 17175 29764 17187 29767
rect 17954 29764 17960 29776
rect 17175 29736 17960 29764
rect 17175 29733 17187 29736
rect 17129 29727 17187 29733
rect 17954 29724 17960 29736
rect 18012 29724 18018 29776
rect 19150 29724 19156 29776
rect 19208 29764 19214 29776
rect 21284 29773 21312 29804
rect 25774 29792 25780 29804
rect 25832 29792 25838 29844
rect 29181 29835 29239 29841
rect 29181 29832 29193 29835
rect 26896 29804 29193 29832
rect 20257 29767 20315 29773
rect 20257 29764 20269 29767
rect 19208 29736 20269 29764
rect 19208 29724 19214 29736
rect 20257 29733 20269 29736
rect 20303 29733 20315 29767
rect 20257 29727 20315 29733
rect 21269 29767 21327 29773
rect 21269 29733 21281 29767
rect 21315 29733 21327 29767
rect 23198 29764 23204 29776
rect 21269 29727 21327 29733
rect 21744 29736 23204 29764
rect 13188 29668 13952 29696
rect 9088 29600 10456 29628
rect 9088 29588 9094 29600
rect 11330 29588 11336 29640
rect 11388 29628 11394 29640
rect 12069 29631 12127 29637
rect 12069 29628 12081 29631
rect 11388 29600 12081 29628
rect 11388 29588 11394 29600
rect 12069 29597 12081 29600
rect 12115 29597 12127 29631
rect 12069 29591 12127 29597
rect 12529 29631 12587 29637
rect 12529 29597 12541 29631
rect 12575 29628 12587 29631
rect 13188 29628 13216 29668
rect 14458 29656 14464 29708
rect 14516 29696 14522 29708
rect 15289 29699 15347 29705
rect 15289 29696 15301 29699
rect 14516 29668 15301 29696
rect 14516 29656 14522 29668
rect 15289 29665 15301 29668
rect 15335 29665 15347 29699
rect 15289 29659 15347 29665
rect 15746 29656 15752 29708
rect 15804 29696 15810 29708
rect 15933 29699 15991 29705
rect 15933 29696 15945 29699
rect 15804 29668 15945 29696
rect 15804 29656 15810 29668
rect 15933 29665 15945 29668
rect 15979 29665 15991 29699
rect 15933 29659 15991 29665
rect 12575 29600 13216 29628
rect 13265 29631 13323 29637
rect 12575 29597 12587 29600
rect 12529 29591 12587 29597
rect 13265 29597 13277 29631
rect 13311 29628 13323 29631
rect 15381 29631 15439 29637
rect 15381 29628 15393 29631
rect 13311 29600 15393 29628
rect 13311 29597 13323 29600
rect 13265 29591 13323 29597
rect 15381 29597 15393 29600
rect 15427 29597 15439 29631
rect 15948 29628 15976 29659
rect 16022 29656 16028 29708
rect 16080 29696 16086 29708
rect 16301 29699 16359 29705
rect 16301 29696 16313 29699
rect 16080 29668 16313 29696
rect 16080 29656 16086 29668
rect 16301 29665 16313 29668
rect 16347 29665 16359 29699
rect 16301 29659 16359 29665
rect 16945 29699 17003 29705
rect 16945 29665 16957 29699
rect 16991 29696 17003 29699
rect 17494 29696 17500 29708
rect 16991 29668 17500 29696
rect 16991 29665 17003 29668
rect 16945 29659 17003 29665
rect 17494 29656 17500 29668
rect 17552 29656 17558 29708
rect 20162 29696 20168 29708
rect 20123 29668 20168 29696
rect 20162 29656 20168 29668
rect 20220 29656 20226 29708
rect 21744 29705 21772 29736
rect 23198 29724 23204 29736
rect 23256 29724 23262 29776
rect 24210 29764 24216 29776
rect 23308 29736 24216 29764
rect 23308 29708 23336 29736
rect 24210 29724 24216 29736
rect 24268 29724 24274 29776
rect 21729 29699 21787 29705
rect 21729 29665 21741 29699
rect 21775 29665 21787 29699
rect 21729 29659 21787 29665
rect 22097 29699 22155 29705
rect 22097 29665 22109 29699
rect 22143 29665 22155 29699
rect 22922 29696 22928 29708
rect 22883 29668 22928 29696
rect 22097 29659 22155 29665
rect 16758 29628 16764 29640
rect 15948 29600 16764 29628
rect 15381 29591 15439 29597
rect 16758 29588 16764 29600
rect 16816 29588 16822 29640
rect 18049 29631 18107 29637
rect 18049 29597 18061 29631
rect 18095 29628 18107 29631
rect 18230 29628 18236 29640
rect 18095 29600 18236 29628
rect 18095 29597 18107 29600
rect 18049 29591 18107 29597
rect 18230 29588 18236 29600
rect 18288 29588 18294 29640
rect 18325 29631 18383 29637
rect 18325 29597 18337 29631
rect 18371 29628 18383 29631
rect 20070 29628 20076 29640
rect 18371 29600 20076 29628
rect 18371 29597 18383 29600
rect 18325 29591 18383 29597
rect 20070 29588 20076 29600
rect 20128 29588 20134 29640
rect 20530 29588 20536 29640
rect 20588 29628 20594 29640
rect 22112 29628 22140 29659
rect 22922 29656 22928 29668
rect 22980 29656 22986 29708
rect 23290 29696 23296 29708
rect 23251 29668 23296 29696
rect 23290 29656 23296 29668
rect 23348 29656 23354 29708
rect 23566 29696 23572 29708
rect 23527 29668 23572 29696
rect 23566 29656 23572 29668
rect 23624 29656 23630 29708
rect 24762 29696 24768 29708
rect 24723 29668 24768 29696
rect 24762 29656 24768 29668
rect 24820 29656 24826 29708
rect 25038 29696 25044 29708
rect 24999 29668 25044 29696
rect 25038 29656 25044 29668
rect 25096 29656 25102 29708
rect 25498 29696 25504 29708
rect 25459 29668 25504 29696
rect 25498 29656 25504 29668
rect 25556 29656 25562 29708
rect 25961 29699 26019 29705
rect 25961 29665 25973 29699
rect 26007 29696 26019 29699
rect 26050 29696 26056 29708
rect 26007 29668 26056 29696
rect 26007 29665 26019 29668
rect 25961 29659 26019 29665
rect 26050 29656 26056 29668
rect 26108 29656 26114 29708
rect 26896 29705 26924 29804
rect 29181 29801 29193 29804
rect 29227 29832 29239 29835
rect 29914 29832 29920 29844
rect 29227 29804 29920 29832
rect 29227 29801 29239 29804
rect 29181 29795 29239 29801
rect 29914 29792 29920 29804
rect 29972 29792 29978 29844
rect 31481 29835 31539 29841
rect 31481 29801 31493 29835
rect 31527 29832 31539 29835
rect 32766 29832 32772 29844
rect 31527 29804 32772 29832
rect 31527 29801 31539 29804
rect 31481 29795 31539 29801
rect 32766 29792 32772 29804
rect 32824 29792 32830 29844
rect 31846 29724 31852 29776
rect 31904 29764 31910 29776
rect 33413 29767 33471 29773
rect 33413 29764 33425 29767
rect 31904 29736 33425 29764
rect 31904 29724 31910 29736
rect 33413 29733 33425 29736
rect 33459 29733 33471 29767
rect 33413 29727 33471 29733
rect 26881 29699 26939 29705
rect 26881 29665 26893 29699
rect 26927 29665 26939 29699
rect 26881 29659 26939 29665
rect 27341 29699 27399 29705
rect 27341 29665 27353 29699
rect 27387 29696 27399 29699
rect 27387 29668 28856 29696
rect 27387 29665 27399 29668
rect 27341 29659 27399 29665
rect 20588 29600 22140 29628
rect 22189 29631 22247 29637
rect 20588 29588 20594 29600
rect 22189 29597 22201 29631
rect 22235 29628 22247 29631
rect 24949 29631 25007 29637
rect 22235 29600 22876 29628
rect 22235 29597 22247 29600
rect 22189 29591 22247 29597
rect 7558 29520 7564 29572
rect 7616 29560 7622 29572
rect 10594 29560 10600 29572
rect 7616 29532 10600 29560
rect 7616 29520 7622 29532
rect 10594 29520 10600 29532
rect 10652 29520 10658 29572
rect 17954 29560 17960 29572
rect 17052 29532 17960 29560
rect 2317 29495 2375 29501
rect 2317 29461 2329 29495
rect 2363 29492 2375 29495
rect 2958 29492 2964 29504
rect 2363 29464 2964 29492
rect 2363 29461 2375 29464
rect 2317 29455 2375 29461
rect 2958 29452 2964 29464
rect 3016 29452 3022 29504
rect 8478 29452 8484 29504
rect 8536 29492 8542 29504
rect 9030 29492 9036 29504
rect 8536 29464 9036 29492
rect 8536 29452 8542 29464
rect 9030 29452 9036 29464
rect 9088 29452 9094 29504
rect 9122 29452 9128 29504
rect 9180 29492 9186 29504
rect 9861 29495 9919 29501
rect 9861 29492 9873 29495
rect 9180 29464 9873 29492
rect 9180 29452 9186 29464
rect 9861 29461 9873 29464
rect 9907 29492 9919 29495
rect 17052 29492 17080 29532
rect 17954 29520 17960 29532
rect 18012 29520 18018 29572
rect 19702 29560 19708 29572
rect 18984 29532 19708 29560
rect 9907 29464 17080 29492
rect 9907 29461 9919 29464
rect 9861 29455 9919 29461
rect 17126 29452 17132 29504
rect 17184 29492 17190 29504
rect 18984 29492 19012 29532
rect 19702 29520 19708 29532
rect 19760 29520 19766 29572
rect 19794 29520 19800 29572
rect 19852 29560 19858 29572
rect 21082 29560 21088 29572
rect 19852 29532 21088 29560
rect 19852 29520 19858 29532
rect 21082 29520 21088 29532
rect 21140 29520 21146 29572
rect 22848 29569 22876 29600
rect 24949 29597 24961 29631
rect 24995 29628 25007 29631
rect 26418 29628 26424 29640
rect 24995 29600 26424 29628
rect 24995 29597 25007 29600
rect 24949 29591 25007 29597
rect 26418 29588 26424 29600
rect 26476 29588 26482 29640
rect 26973 29631 27031 29637
rect 26973 29597 26985 29631
rect 27019 29628 27031 29631
rect 27614 29628 27620 29640
rect 27019 29600 27620 29628
rect 27019 29597 27031 29600
rect 26973 29591 27031 29597
rect 27614 29588 27620 29600
rect 27672 29588 27678 29640
rect 27801 29631 27859 29637
rect 27801 29597 27813 29631
rect 27847 29597 27859 29631
rect 28074 29628 28080 29640
rect 28035 29600 28080 29628
rect 27801 29591 27859 29597
rect 22833 29563 22891 29569
rect 22833 29529 22845 29563
rect 22879 29529 22891 29563
rect 22833 29523 22891 29529
rect 27430 29520 27436 29572
rect 27488 29560 27494 29572
rect 27816 29560 27844 29591
rect 28074 29588 28080 29600
rect 28132 29588 28138 29640
rect 28828 29628 28856 29668
rect 29270 29656 29276 29708
rect 29328 29696 29334 29708
rect 29917 29699 29975 29705
rect 29917 29696 29929 29699
rect 29328 29668 29929 29696
rect 29328 29656 29334 29668
rect 29917 29665 29929 29668
rect 29963 29665 29975 29699
rect 30282 29696 30288 29708
rect 30195 29668 30288 29696
rect 29917 29659 29975 29665
rect 30282 29656 30288 29668
rect 30340 29656 30346 29708
rect 30466 29656 30472 29708
rect 30524 29696 30530 29708
rect 30745 29699 30803 29705
rect 30745 29696 30757 29699
rect 30524 29668 30757 29696
rect 30524 29656 30530 29668
rect 30745 29665 30757 29668
rect 30791 29665 30803 29699
rect 30745 29659 30803 29665
rect 31018 29656 31024 29708
rect 31076 29696 31082 29708
rect 31665 29699 31723 29705
rect 31665 29696 31677 29699
rect 31076 29668 31677 29696
rect 31076 29656 31082 29668
rect 31665 29665 31677 29668
rect 31711 29665 31723 29699
rect 32858 29696 32864 29708
rect 32819 29668 32864 29696
rect 31665 29659 31723 29665
rect 32858 29656 32864 29668
rect 32916 29656 32922 29708
rect 33134 29696 33140 29708
rect 33095 29668 33140 29696
rect 33134 29656 33140 29668
rect 33192 29656 33198 29708
rect 33594 29656 33600 29708
rect 33652 29696 33658 29708
rect 33873 29699 33931 29705
rect 33873 29696 33885 29699
rect 33652 29668 33885 29696
rect 33652 29656 33658 29668
rect 33873 29665 33885 29668
rect 33919 29665 33931 29699
rect 33873 29659 33931 29665
rect 35618 29656 35624 29708
rect 35676 29696 35682 29708
rect 36081 29699 36139 29705
rect 36081 29696 36093 29699
rect 35676 29668 36093 29696
rect 35676 29656 35682 29668
rect 36081 29665 36093 29668
rect 36127 29665 36139 29699
rect 36814 29696 36820 29708
rect 36775 29668 36820 29696
rect 36081 29659 36139 29665
rect 36814 29656 36820 29668
rect 36872 29656 36878 29708
rect 37642 29656 37648 29708
rect 37700 29696 37706 29708
rect 37737 29699 37795 29705
rect 37737 29696 37749 29699
rect 37700 29668 37749 29696
rect 37700 29656 37706 29668
rect 37737 29665 37749 29668
rect 37783 29665 37795 29699
rect 37737 29659 37795 29665
rect 29638 29628 29644 29640
rect 28828 29600 29644 29628
rect 29638 29588 29644 29600
rect 29696 29588 29702 29640
rect 30300 29628 30328 29656
rect 31754 29628 31760 29640
rect 30300 29600 31760 29628
rect 31754 29588 31760 29600
rect 31812 29588 31818 29640
rect 32493 29631 32551 29637
rect 32493 29597 32505 29631
rect 32539 29628 32551 29631
rect 32950 29628 32956 29640
rect 32539 29600 32956 29628
rect 32539 29597 32551 29600
rect 32493 29591 32551 29597
rect 32950 29588 32956 29600
rect 33008 29588 33014 29640
rect 34146 29628 34152 29640
rect 34107 29600 34152 29628
rect 34146 29588 34152 29600
rect 34204 29588 34210 29640
rect 37090 29628 37096 29640
rect 37051 29600 37096 29628
rect 37090 29588 37096 29600
rect 37148 29588 37154 29640
rect 27488 29532 27844 29560
rect 30837 29563 30895 29569
rect 27488 29520 27494 29532
rect 30837 29529 30849 29563
rect 30883 29560 30895 29563
rect 32766 29560 32772 29572
rect 30883 29532 32772 29560
rect 30883 29529 30895 29532
rect 30837 29523 30895 29529
rect 32766 29520 32772 29532
rect 32824 29520 32830 29572
rect 36357 29563 36415 29569
rect 36357 29529 36369 29563
rect 36403 29560 36415 29563
rect 36722 29560 36728 29572
rect 36403 29532 36728 29560
rect 36403 29529 36415 29532
rect 36357 29523 36415 29529
rect 36722 29520 36728 29532
rect 36780 29520 36786 29572
rect 17184 29464 19012 29492
rect 17184 29452 17190 29464
rect 19426 29452 19432 29504
rect 19484 29492 19490 29504
rect 19613 29495 19671 29501
rect 19613 29492 19625 29495
rect 19484 29464 19625 29492
rect 19484 29452 19490 29464
rect 19613 29461 19625 29464
rect 19659 29492 19671 29495
rect 20162 29492 20168 29504
rect 19659 29464 20168 29492
rect 19659 29461 19671 29464
rect 19613 29455 19671 29461
rect 20162 29452 20168 29464
rect 20220 29452 20226 29504
rect 35250 29492 35256 29504
rect 35211 29464 35256 29492
rect 35250 29452 35256 29464
rect 35308 29452 35314 29504
rect 36814 29452 36820 29504
rect 36872 29492 36878 29504
rect 37921 29495 37979 29501
rect 37921 29492 37933 29495
rect 36872 29464 37933 29492
rect 36872 29452 36878 29464
rect 37921 29461 37933 29464
rect 37967 29461 37979 29495
rect 37921 29455 37979 29461
rect 1104 29402 38824 29424
rect 1104 29350 4246 29402
rect 4298 29350 4310 29402
rect 4362 29350 4374 29402
rect 4426 29350 4438 29402
rect 4490 29350 34966 29402
rect 35018 29350 35030 29402
rect 35082 29350 35094 29402
rect 35146 29350 35158 29402
rect 35210 29350 38824 29402
rect 1104 29328 38824 29350
rect 4062 29248 4068 29300
rect 4120 29288 4126 29300
rect 6917 29291 6975 29297
rect 6917 29288 6929 29291
rect 4120 29260 6929 29288
rect 4120 29248 4126 29260
rect 6917 29257 6929 29260
rect 6963 29257 6975 29291
rect 6917 29251 6975 29257
rect 9950 29248 9956 29300
rect 10008 29288 10014 29300
rect 10321 29291 10379 29297
rect 10321 29288 10333 29291
rect 10008 29260 10333 29288
rect 10008 29248 10014 29260
rect 10321 29257 10333 29260
rect 10367 29257 10379 29291
rect 10321 29251 10379 29257
rect 18230 29248 18236 29300
rect 18288 29288 18294 29300
rect 19794 29288 19800 29300
rect 18288 29260 19800 29288
rect 18288 29248 18294 29260
rect 19794 29248 19800 29260
rect 19852 29248 19858 29300
rect 20438 29248 20444 29300
rect 20496 29288 20502 29300
rect 21726 29288 21732 29300
rect 20496 29260 21732 29288
rect 20496 29248 20502 29260
rect 21726 29248 21732 29260
rect 21784 29248 21790 29300
rect 26418 29248 26424 29300
rect 26476 29288 26482 29300
rect 26878 29288 26884 29300
rect 26476 29260 26884 29288
rect 26476 29248 26482 29260
rect 26878 29248 26884 29260
rect 26936 29248 26942 29300
rect 28905 29291 28963 29297
rect 28905 29257 28917 29291
rect 28951 29288 28963 29291
rect 31018 29288 31024 29300
rect 28951 29260 31024 29288
rect 28951 29257 28963 29260
rect 28905 29251 28963 29257
rect 4080 29152 4108 29248
rect 6086 29180 6092 29232
rect 6144 29220 6150 29232
rect 6181 29223 6239 29229
rect 6181 29220 6193 29223
rect 6144 29192 6193 29220
rect 6144 29180 6150 29192
rect 6181 29189 6193 29192
rect 6227 29189 6239 29223
rect 12710 29220 12716 29232
rect 12623 29192 12716 29220
rect 6181 29183 6239 29189
rect 3528 29124 4108 29152
rect 1857 29087 1915 29093
rect 1857 29053 1869 29087
rect 1903 29053 1915 29087
rect 1857 29047 1915 29053
rect 1949 29087 2007 29093
rect 1949 29053 1961 29087
rect 1995 29084 2007 29087
rect 2685 29087 2743 29093
rect 2685 29084 2697 29087
rect 1995 29056 2697 29084
rect 1995 29053 2007 29056
rect 1949 29047 2007 29053
rect 2685 29053 2697 29056
rect 2731 29084 2743 29087
rect 2774 29084 2780 29096
rect 2731 29056 2780 29084
rect 2731 29053 2743 29056
rect 2685 29047 2743 29053
rect 1872 29016 1900 29047
rect 2774 29044 2780 29056
rect 2832 29044 2838 29096
rect 2958 29084 2964 29096
rect 2919 29056 2964 29084
rect 2958 29044 2964 29056
rect 3016 29044 3022 29096
rect 3234 29044 3240 29096
rect 3292 29084 3298 29096
rect 3528 29093 3556 29124
rect 4706 29112 4712 29164
rect 4764 29152 4770 29164
rect 5261 29155 5319 29161
rect 5261 29152 5273 29155
rect 4764 29124 5273 29152
rect 4764 29112 4770 29124
rect 5261 29121 5273 29124
rect 5307 29121 5319 29155
rect 5261 29115 5319 29121
rect 5902 29112 5908 29164
rect 5960 29152 5966 29164
rect 6822 29152 6828 29164
rect 5960 29124 6828 29152
rect 5960 29112 5966 29124
rect 6822 29112 6828 29124
rect 6880 29152 6886 29164
rect 8389 29155 8447 29161
rect 6880 29124 7420 29152
rect 6880 29112 6886 29124
rect 3513 29087 3571 29093
rect 3513 29084 3525 29087
rect 3292 29056 3525 29084
rect 3292 29044 3298 29056
rect 3513 29053 3525 29056
rect 3559 29053 3571 29087
rect 3513 29047 3571 29053
rect 3881 29087 3939 29093
rect 3881 29053 3893 29087
rect 3927 29084 3939 29087
rect 4062 29084 4068 29096
rect 3927 29056 4068 29084
rect 3927 29053 3939 29056
rect 3881 29047 3939 29053
rect 4062 29044 4068 29056
rect 4120 29044 4126 29096
rect 4525 29087 4583 29093
rect 4525 29053 4537 29087
rect 4571 29053 4583 29087
rect 4525 29047 4583 29053
rect 4540 29016 4568 29047
rect 4614 29044 4620 29096
rect 4672 29084 4678 29096
rect 4985 29087 5043 29093
rect 4985 29084 4997 29087
rect 4672 29056 4997 29084
rect 4672 29044 4678 29056
rect 4985 29053 4997 29056
rect 5031 29053 5043 29087
rect 4985 29047 5043 29053
rect 5997 29087 6055 29093
rect 5997 29053 6009 29087
rect 6043 29053 6055 29087
rect 7006 29084 7012 29096
rect 6967 29056 7012 29084
rect 5997 29047 6055 29053
rect 4798 29016 4804 29028
rect 1872 28988 3004 29016
rect 4540 28988 4804 29016
rect 2976 28960 3004 28988
rect 4798 28976 4804 28988
rect 4856 29016 4862 29028
rect 5166 29016 5172 29028
rect 4856 28988 5172 29016
rect 4856 28976 4862 28988
rect 5166 28976 5172 28988
rect 5224 28976 5230 29028
rect 6012 29016 6040 29047
rect 7006 29044 7012 29056
rect 7064 29044 7070 29096
rect 7392 29093 7420 29124
rect 8389 29121 8401 29155
rect 8435 29152 8447 29155
rect 10410 29152 10416 29164
rect 8435 29124 10416 29152
rect 8435 29121 8447 29124
rect 8389 29115 8447 29121
rect 10410 29112 10416 29124
rect 10468 29112 10474 29164
rect 12158 29152 12164 29164
rect 10520 29124 12164 29152
rect 7377 29087 7435 29093
rect 7377 29053 7389 29087
rect 7423 29053 7435 29087
rect 7377 29047 7435 29053
rect 8113 29087 8171 29093
rect 8113 29053 8125 29087
rect 8159 29084 8171 29087
rect 8662 29084 8668 29096
rect 8159 29056 8668 29084
rect 8159 29053 8171 29056
rect 8113 29047 8171 29053
rect 8662 29044 8668 29056
rect 8720 29084 8726 29096
rect 9398 29084 9404 29096
rect 8720 29056 9404 29084
rect 8720 29044 8726 29056
rect 9398 29044 9404 29056
rect 9456 29044 9462 29096
rect 10520 29093 10548 29124
rect 12158 29112 12164 29124
rect 12216 29112 12222 29164
rect 10505 29087 10563 29093
rect 10505 29053 10517 29087
rect 10551 29053 10563 29087
rect 10505 29047 10563 29053
rect 10597 29087 10655 29093
rect 10597 29053 10609 29087
rect 10643 29084 10655 29087
rect 10686 29084 10692 29096
rect 10643 29056 10692 29084
rect 10643 29053 10655 29056
rect 10597 29047 10655 29053
rect 6914 29016 6920 29028
rect 6012 28988 6920 29016
rect 6914 28976 6920 28988
rect 6972 28976 6978 29028
rect 10612 29016 10640 29047
rect 10686 29044 10692 29056
rect 10744 29044 10750 29096
rect 12636 29093 12664 29192
rect 12710 29180 12716 29192
rect 12768 29220 12774 29232
rect 14274 29220 14280 29232
rect 12768 29192 14280 29220
rect 12768 29180 12774 29192
rect 14274 29180 14280 29192
rect 14332 29180 14338 29232
rect 14461 29223 14519 29229
rect 14461 29189 14473 29223
rect 14507 29220 14519 29223
rect 15838 29220 15844 29232
rect 14507 29192 15844 29220
rect 14507 29189 14519 29192
rect 14461 29183 14519 29189
rect 15838 29180 15844 29192
rect 15896 29180 15902 29232
rect 19426 29220 19432 29232
rect 18340 29192 19432 29220
rect 14550 29152 14556 29164
rect 13188 29124 14556 29152
rect 11241 29087 11299 29093
rect 11241 29053 11253 29087
rect 11287 29053 11299 29087
rect 11241 29047 11299 29053
rect 12621 29087 12679 29093
rect 12621 29053 12633 29087
rect 12667 29053 12679 29087
rect 12621 29047 12679 29053
rect 9508 28988 10640 29016
rect 11256 29016 11284 29047
rect 12710 29044 12716 29096
rect 12768 29084 12774 29096
rect 13188 29093 13216 29124
rect 14550 29112 14556 29124
rect 14608 29152 14614 29164
rect 15013 29155 15071 29161
rect 15013 29152 15025 29155
rect 14608 29124 15025 29152
rect 14608 29112 14614 29124
rect 15013 29121 15025 29124
rect 15059 29121 15071 29155
rect 15013 29115 15071 29121
rect 16022 29112 16028 29164
rect 16080 29152 16086 29164
rect 18340 29161 18368 29192
rect 19426 29180 19432 29192
rect 19484 29180 19490 29232
rect 21174 29180 21180 29232
rect 21232 29220 21238 29232
rect 28074 29220 28080 29232
rect 21232 29192 22416 29220
rect 28035 29192 28080 29220
rect 21232 29180 21238 29192
rect 17221 29155 17279 29161
rect 17221 29152 17233 29155
rect 16080 29124 17233 29152
rect 16080 29112 16086 29124
rect 17221 29121 17233 29124
rect 17267 29121 17279 29155
rect 17221 29115 17279 29121
rect 18325 29155 18383 29161
rect 18325 29121 18337 29155
rect 18371 29121 18383 29155
rect 19334 29152 19340 29164
rect 18325 29115 18383 29121
rect 18708 29124 19340 29152
rect 12805 29087 12863 29093
rect 12805 29084 12817 29087
rect 12768 29056 12817 29084
rect 12768 29044 12774 29056
rect 12805 29053 12817 29056
rect 12851 29053 12863 29087
rect 12805 29047 12863 29053
rect 13173 29087 13231 29093
rect 13173 29053 13185 29087
rect 13219 29053 13231 29087
rect 14366 29084 14372 29096
rect 14327 29056 14372 29084
rect 13173 29047 13231 29053
rect 14366 29044 14372 29056
rect 14424 29044 14430 29096
rect 14918 29084 14924 29096
rect 14879 29056 14924 29084
rect 14918 29044 14924 29056
rect 14976 29044 14982 29096
rect 15841 29087 15899 29093
rect 15841 29053 15853 29087
rect 15887 29084 15899 29087
rect 16117 29087 16175 29093
rect 15887 29056 15976 29084
rect 15887 29053 15899 29056
rect 15841 29047 15899 29053
rect 13354 29016 13360 29028
rect 11256 28988 13360 29016
rect 2777 28951 2835 28957
rect 2777 28917 2789 28951
rect 2823 28948 2835 28951
rect 2866 28948 2872 28960
rect 2823 28920 2872 28948
rect 2823 28917 2835 28920
rect 2777 28911 2835 28917
rect 2866 28908 2872 28920
rect 2924 28908 2930 28960
rect 2958 28908 2964 28960
rect 3016 28908 3022 28960
rect 4525 28951 4583 28957
rect 4525 28917 4537 28951
rect 4571 28948 4583 28951
rect 4890 28948 4896 28960
rect 4571 28920 4896 28948
rect 4571 28917 4583 28920
rect 4525 28911 4583 28917
rect 4890 28908 4896 28920
rect 4948 28908 4954 28960
rect 7558 28908 7564 28960
rect 7616 28948 7622 28960
rect 9508 28948 9536 28988
rect 13354 28976 13360 28988
rect 13412 28976 13418 29028
rect 7616 28920 9536 28948
rect 7616 28908 7622 28920
rect 9674 28908 9680 28960
rect 9732 28948 9738 28960
rect 15948 28948 15976 29056
rect 16117 29053 16129 29087
rect 16163 29084 16175 29087
rect 17034 29084 17040 29096
rect 16163 29056 17040 29084
rect 16163 29053 16175 29056
rect 16117 29047 16175 29053
rect 17034 29044 17040 29056
rect 17092 29044 17098 29096
rect 18708 29093 18736 29124
rect 19334 29112 19340 29124
rect 19392 29152 19398 29164
rect 19392 29124 20300 29152
rect 19392 29112 19398 29124
rect 20272 29096 20300 29124
rect 18693 29087 18751 29093
rect 18693 29053 18705 29087
rect 18739 29053 18751 29087
rect 18966 29084 18972 29096
rect 18927 29056 18972 29084
rect 18693 29047 18751 29053
rect 18966 29044 18972 29056
rect 19024 29044 19030 29096
rect 19794 29044 19800 29096
rect 19852 29084 19858 29096
rect 20165 29087 20223 29093
rect 20165 29084 20177 29087
rect 19852 29056 20177 29084
rect 19852 29044 19858 29056
rect 20165 29053 20177 29056
rect 20211 29053 20223 29087
rect 20165 29047 20223 29053
rect 20254 29044 20260 29096
rect 20312 29044 20318 29096
rect 20438 29084 20444 29096
rect 20399 29056 20444 29084
rect 20438 29044 20444 29056
rect 20496 29044 20502 29096
rect 22388 29093 22416 29192
rect 28074 29180 28080 29192
rect 28132 29180 28138 29232
rect 22646 29152 22652 29164
rect 22607 29124 22652 29152
rect 22646 29112 22652 29124
rect 22704 29112 22710 29164
rect 22922 29112 22928 29164
rect 22980 29152 22986 29164
rect 23842 29152 23848 29164
rect 22980 29124 23848 29152
rect 22980 29112 22986 29124
rect 23032 29093 23060 29124
rect 23842 29112 23848 29124
rect 23900 29152 23906 29164
rect 24670 29152 24676 29164
rect 23900 29124 24676 29152
rect 23900 29112 23906 29124
rect 24670 29112 24676 29124
rect 24728 29112 24734 29164
rect 25041 29155 25099 29161
rect 25041 29121 25053 29155
rect 25087 29152 25099 29155
rect 25087 29124 27568 29152
rect 25087 29121 25099 29124
rect 25041 29115 25099 29121
rect 22373 29087 22431 29093
rect 22373 29053 22385 29087
rect 22419 29053 22431 29087
rect 22373 29047 22431 29053
rect 23017 29087 23075 29093
rect 23017 29053 23029 29087
rect 23063 29053 23075 29087
rect 23017 29047 23075 29053
rect 23661 29087 23719 29093
rect 23661 29053 23673 29087
rect 23707 29084 23719 29087
rect 24762 29084 24768 29096
rect 23707 29056 24440 29084
rect 24723 29056 24768 29084
rect 23707 29053 23719 29056
rect 23661 29047 23719 29053
rect 19150 29016 19156 29028
rect 16776 28988 19156 29016
rect 16776 28948 16804 28988
rect 19150 28976 19156 28988
rect 19208 28976 19214 29028
rect 19245 29019 19303 29025
rect 19245 28985 19257 29019
rect 19291 29016 19303 29019
rect 19978 29016 19984 29028
rect 19291 28988 19984 29016
rect 19291 28985 19303 28988
rect 19245 28979 19303 28985
rect 19978 28976 19984 28988
rect 20036 28976 20042 29028
rect 23382 28976 23388 29028
rect 23440 29016 23446 29028
rect 23753 29019 23811 29025
rect 23753 29016 23765 29019
rect 23440 28988 23765 29016
rect 23440 28976 23446 28988
rect 23753 28985 23765 28988
rect 23799 28985 23811 29019
rect 24412 29016 24440 29056
rect 24762 29044 24768 29056
rect 24820 29044 24826 29096
rect 25222 29084 25228 29096
rect 25183 29056 25228 29084
rect 25222 29044 25228 29056
rect 25280 29044 25286 29096
rect 25314 29044 25320 29096
rect 25372 29084 25378 29096
rect 25409 29087 25467 29093
rect 25409 29084 25421 29087
rect 25372 29056 25421 29084
rect 25372 29044 25378 29056
rect 25409 29053 25421 29056
rect 25455 29053 25467 29087
rect 26050 29084 26056 29096
rect 26011 29056 26056 29084
rect 25409 29047 25467 29053
rect 26050 29044 26056 29056
rect 26108 29044 26114 29096
rect 27065 29087 27123 29093
rect 27065 29053 27077 29087
rect 27111 29053 27123 29087
rect 27065 29047 27123 29053
rect 26142 29016 26148 29028
rect 24412 28988 26148 29016
rect 23753 28979 23811 28985
rect 26142 28976 26148 28988
rect 26200 28976 26206 29028
rect 27080 29016 27108 29047
rect 27154 29044 27160 29096
rect 27212 29084 27218 29096
rect 27540 29093 27568 29124
rect 27525 29087 27583 29093
rect 27212 29056 27257 29084
rect 27212 29044 27218 29056
rect 27525 29053 27537 29087
rect 27571 29053 27583 29087
rect 27525 29047 27583 29053
rect 27614 29044 27620 29096
rect 27672 29084 27678 29096
rect 27985 29087 28043 29093
rect 27985 29084 27997 29087
rect 27672 29056 27997 29084
rect 27672 29044 27678 29056
rect 27985 29053 27997 29056
rect 28031 29053 28043 29087
rect 27985 29047 28043 29053
rect 28920 29016 28948 29251
rect 31018 29248 31024 29260
rect 31076 29248 31082 29300
rect 32950 29288 32956 29300
rect 32911 29260 32956 29288
rect 32950 29248 32956 29260
rect 33008 29248 33014 29300
rect 37734 29248 37740 29300
rect 37792 29288 37798 29300
rect 37829 29291 37887 29297
rect 37829 29288 37841 29291
rect 37792 29260 37841 29288
rect 37792 29248 37798 29260
rect 37829 29257 37841 29260
rect 37875 29257 37887 29291
rect 37829 29251 37887 29257
rect 34422 29180 34428 29232
rect 34480 29220 34486 29232
rect 34480 29192 35480 29220
rect 34480 29180 34486 29192
rect 29914 29152 29920 29164
rect 29875 29124 29920 29152
rect 29914 29112 29920 29124
rect 29972 29112 29978 29164
rect 30926 29152 30932 29164
rect 30887 29124 30932 29152
rect 30926 29112 30932 29124
rect 30984 29112 30990 29164
rect 31386 29152 31392 29164
rect 31347 29124 31392 29152
rect 31386 29112 31392 29124
rect 31444 29112 31450 29164
rect 31662 29152 31668 29164
rect 31623 29124 31668 29152
rect 31662 29112 31668 29124
rect 31720 29112 31726 29164
rect 34333 29155 34391 29161
rect 34333 29121 34345 29155
rect 34379 29152 34391 29155
rect 35342 29152 35348 29164
rect 34379 29124 35348 29152
rect 34379 29121 34391 29124
rect 34333 29115 34391 29121
rect 35342 29112 35348 29124
rect 35400 29112 35406 29164
rect 35452 29161 35480 29192
rect 35437 29155 35495 29161
rect 35437 29121 35449 29155
rect 35483 29121 35495 29155
rect 36446 29152 36452 29164
rect 36407 29124 36452 29152
rect 35437 29115 35495 29121
rect 36446 29112 36452 29124
rect 36504 29112 36510 29164
rect 36722 29152 36728 29164
rect 36683 29124 36728 29152
rect 36722 29112 36728 29124
rect 36780 29112 36786 29164
rect 29089 29087 29147 29093
rect 29089 29053 29101 29087
rect 29135 29084 29147 29087
rect 29454 29084 29460 29096
rect 29135 29056 29460 29084
rect 29135 29053 29147 29056
rect 29089 29047 29147 29053
rect 29454 29044 29460 29056
rect 29512 29044 29518 29096
rect 30374 29084 30380 29096
rect 30335 29056 30380 29084
rect 30374 29044 30380 29056
rect 30432 29044 30438 29096
rect 30466 29044 30472 29096
rect 30524 29084 30530 29096
rect 30653 29087 30711 29093
rect 30653 29084 30665 29087
rect 30524 29056 30665 29084
rect 30524 29044 30530 29056
rect 30653 29053 30665 29056
rect 30699 29053 30711 29087
rect 30653 29047 30711 29053
rect 33965 29087 34023 29093
rect 33965 29053 33977 29087
rect 34011 29084 34023 29087
rect 35250 29084 35256 29096
rect 34011 29056 35256 29084
rect 34011 29053 34023 29056
rect 33965 29047 34023 29053
rect 35250 29044 35256 29056
rect 35308 29044 35314 29096
rect 35526 29044 35532 29096
rect 35584 29084 35590 29096
rect 35713 29087 35771 29093
rect 35713 29084 35725 29087
rect 35584 29056 35725 29084
rect 35584 29044 35590 29056
rect 35713 29053 35725 29056
rect 35759 29053 35771 29087
rect 35713 29047 35771 29053
rect 35897 29087 35955 29093
rect 35897 29053 35909 29087
rect 35943 29053 35955 29087
rect 35897 29047 35955 29053
rect 27080 28988 28948 29016
rect 33502 28976 33508 29028
rect 33560 29016 33566 29028
rect 33781 29019 33839 29025
rect 33781 29016 33793 29019
rect 33560 28988 33793 29016
rect 33560 28976 33566 28988
rect 33781 28985 33793 28988
rect 33827 28985 33839 29019
rect 33781 28979 33839 28985
rect 34698 28976 34704 29028
rect 34756 29016 34762 29028
rect 34885 29019 34943 29025
rect 34885 29016 34897 29019
rect 34756 28988 34897 29016
rect 34756 28976 34762 28988
rect 34885 28985 34897 28988
rect 34931 28985 34943 29019
rect 34885 28979 34943 28985
rect 35434 28976 35440 29028
rect 35492 29016 35498 29028
rect 35912 29016 35940 29047
rect 37918 29016 37924 29028
rect 35492 28988 35940 29016
rect 35492 28976 35498 28988
rect 9732 28920 9777 28948
rect 15948 28920 16804 28948
rect 9732 28908 9738 28920
rect 20162 28908 20168 28960
rect 20220 28948 20226 28960
rect 20806 28948 20812 28960
rect 20220 28920 20812 28948
rect 20220 28908 20226 28920
rect 20806 28908 20812 28920
rect 20864 28908 20870 28960
rect 21082 28908 21088 28960
rect 21140 28948 21146 28960
rect 21545 28951 21603 28957
rect 21545 28948 21557 28951
rect 21140 28920 21557 28948
rect 21140 28908 21146 28920
rect 21545 28917 21557 28920
rect 21591 28917 21603 28951
rect 35912 28948 35940 28988
rect 37844 28988 37924 29016
rect 36722 28948 36728 28960
rect 35912 28920 36728 28948
rect 21545 28911 21603 28917
rect 36722 28908 36728 28920
rect 36780 28908 36786 28960
rect 37844 28948 37872 28988
rect 37918 28976 37924 28988
rect 37976 28976 37982 29028
rect 38010 28948 38016 28960
rect 37844 28920 38016 28948
rect 38010 28908 38016 28920
rect 38068 28908 38074 28960
rect 1104 28858 38824 28880
rect 1104 28806 19606 28858
rect 19658 28806 19670 28858
rect 19722 28806 19734 28858
rect 19786 28806 19798 28858
rect 19850 28806 38824 28858
rect 1104 28784 38824 28806
rect 7374 28704 7380 28756
rect 7432 28744 7438 28756
rect 7469 28747 7527 28753
rect 7469 28744 7481 28747
rect 7432 28716 7481 28744
rect 7432 28704 7438 28716
rect 7469 28713 7481 28716
rect 7515 28713 7527 28747
rect 7469 28707 7527 28713
rect 11606 28704 11612 28756
rect 11664 28744 11670 28756
rect 13262 28744 13268 28756
rect 11664 28716 13268 28744
rect 11664 28704 11670 28716
rect 13262 28704 13268 28716
rect 13320 28704 13326 28756
rect 13354 28704 13360 28756
rect 13412 28744 13418 28756
rect 14277 28747 14335 28753
rect 14277 28744 14289 28747
rect 13412 28716 14289 28744
rect 13412 28704 13418 28716
rect 14277 28713 14289 28716
rect 14323 28713 14335 28747
rect 17034 28744 17040 28756
rect 16995 28716 17040 28744
rect 14277 28707 14335 28713
rect 17034 28704 17040 28716
rect 17092 28704 17098 28756
rect 20349 28747 20407 28753
rect 20349 28713 20361 28747
rect 20395 28744 20407 28747
rect 20438 28744 20444 28756
rect 20395 28716 20444 28744
rect 20395 28713 20407 28716
rect 20349 28707 20407 28713
rect 20438 28704 20444 28716
rect 20496 28704 20502 28756
rect 20622 28704 20628 28756
rect 20680 28744 20686 28756
rect 20993 28747 21051 28753
rect 20993 28744 21005 28747
rect 20680 28716 21005 28744
rect 20680 28704 20686 28716
rect 20993 28713 21005 28716
rect 21039 28713 21051 28747
rect 20993 28707 21051 28713
rect 21542 28704 21548 28756
rect 21600 28744 21606 28756
rect 21637 28747 21695 28753
rect 21637 28744 21649 28747
rect 21600 28716 21649 28744
rect 21600 28704 21606 28716
rect 21637 28713 21649 28716
rect 21683 28713 21695 28747
rect 22278 28744 22284 28756
rect 22239 28716 22284 28744
rect 21637 28707 21695 28713
rect 22278 28704 22284 28716
rect 22336 28704 22342 28756
rect 32306 28744 32312 28756
rect 25792 28716 32312 28744
rect 5442 28636 5448 28688
rect 5500 28676 5506 28688
rect 5500 28648 6224 28676
rect 5500 28636 5506 28648
rect 4614 28608 4620 28620
rect 4575 28580 4620 28608
rect 4614 28568 4620 28580
rect 4672 28568 4678 28620
rect 4890 28608 4896 28620
rect 4851 28580 4896 28608
rect 4890 28568 4896 28580
rect 4948 28568 4954 28620
rect 5810 28608 5816 28620
rect 5771 28580 5816 28608
rect 5810 28568 5816 28580
rect 5868 28568 5874 28620
rect 6196 28617 6224 28648
rect 11422 28636 11428 28688
rect 11480 28676 11486 28688
rect 12161 28679 12219 28685
rect 12161 28676 12173 28679
rect 11480 28648 12173 28676
rect 11480 28636 11486 28648
rect 12161 28645 12173 28648
rect 12207 28676 12219 28679
rect 16485 28679 16543 28685
rect 12207 28648 13216 28676
rect 12207 28645 12219 28648
rect 12161 28639 12219 28645
rect 6181 28611 6239 28617
rect 6181 28577 6193 28611
rect 6227 28608 6239 28611
rect 7193 28611 7251 28617
rect 7193 28608 7205 28611
rect 6227 28580 7205 28608
rect 6227 28577 6239 28580
rect 6181 28571 6239 28577
rect 7193 28577 7205 28580
rect 7239 28577 7251 28611
rect 7193 28571 7251 28577
rect 7653 28611 7711 28617
rect 7653 28577 7665 28611
rect 7699 28577 7711 28611
rect 7653 28571 7711 28577
rect 1394 28540 1400 28552
rect 1355 28512 1400 28540
rect 1394 28500 1400 28512
rect 1452 28500 1458 28552
rect 1673 28543 1731 28549
rect 1673 28509 1685 28543
rect 1719 28540 1731 28543
rect 1854 28540 1860 28552
rect 1719 28512 1860 28540
rect 1719 28509 1731 28512
rect 1673 28503 1731 28509
rect 1854 28500 1860 28512
rect 1912 28500 1918 28552
rect 4249 28543 4307 28549
rect 4249 28509 4261 28543
rect 4295 28540 4307 28543
rect 4706 28540 4712 28552
rect 4295 28512 4712 28540
rect 4295 28509 4307 28512
rect 4249 28503 4307 28509
rect 4706 28500 4712 28512
rect 4764 28500 4770 28552
rect 5350 28500 5356 28552
rect 5408 28540 5414 28552
rect 6641 28543 6699 28549
rect 6641 28540 6653 28543
rect 5408 28512 6653 28540
rect 5408 28500 5414 28512
rect 6641 28509 6653 28512
rect 6687 28540 6699 28543
rect 7668 28540 7696 28571
rect 7926 28568 7932 28620
rect 7984 28608 7990 28620
rect 8389 28611 8447 28617
rect 8389 28608 8401 28611
rect 7984 28580 8401 28608
rect 7984 28568 7990 28580
rect 8389 28577 8401 28580
rect 8435 28577 8447 28611
rect 9950 28608 9956 28620
rect 9911 28580 9956 28608
rect 8389 28571 8447 28577
rect 9950 28568 9956 28580
rect 10008 28568 10014 28620
rect 10045 28611 10103 28617
rect 10045 28577 10057 28611
rect 10091 28608 10103 28611
rect 10318 28608 10324 28620
rect 10091 28580 10324 28608
rect 10091 28577 10103 28580
rect 10045 28571 10103 28577
rect 10318 28568 10324 28580
rect 10376 28568 10382 28620
rect 10413 28611 10471 28617
rect 10413 28577 10425 28611
rect 10459 28608 10471 28611
rect 10594 28608 10600 28620
rect 10459 28580 10600 28608
rect 10459 28577 10471 28580
rect 10413 28571 10471 28577
rect 10594 28568 10600 28580
rect 10652 28568 10658 28620
rect 11333 28611 11391 28617
rect 11333 28577 11345 28611
rect 11379 28608 11391 28611
rect 11606 28608 11612 28620
rect 11379 28580 11612 28608
rect 11379 28577 11391 28580
rect 11333 28571 11391 28577
rect 11606 28568 11612 28580
rect 11664 28568 11670 28620
rect 11885 28611 11943 28617
rect 11885 28577 11897 28611
rect 11931 28577 11943 28611
rect 11885 28571 11943 28577
rect 12069 28611 12127 28617
rect 12069 28577 12081 28611
rect 12115 28608 12127 28611
rect 12710 28608 12716 28620
rect 12115 28580 12716 28608
rect 12115 28577 12127 28580
rect 12069 28571 12127 28577
rect 6687 28512 7696 28540
rect 11900 28540 11928 28571
rect 12710 28568 12716 28580
rect 12768 28568 12774 28620
rect 12989 28611 13047 28617
rect 12989 28577 13001 28611
rect 13035 28577 13047 28611
rect 12989 28571 13047 28577
rect 12894 28540 12900 28552
rect 11900 28512 12900 28540
rect 6687 28509 6699 28512
rect 6641 28503 6699 28509
rect 12894 28500 12900 28512
rect 12952 28540 12958 28552
rect 13004 28540 13032 28571
rect 12952 28512 13032 28540
rect 13188 28540 13216 28648
rect 13372 28648 14228 28676
rect 13372 28540 13400 28648
rect 13446 28568 13452 28620
rect 13504 28608 13510 28620
rect 14200 28617 14228 28648
rect 16485 28645 16497 28679
rect 16531 28676 16543 28679
rect 20530 28676 20536 28688
rect 16531 28648 20536 28676
rect 16531 28645 16543 28648
rect 16485 28639 16543 28645
rect 20530 28636 20536 28648
rect 20588 28636 20594 28688
rect 20806 28636 20812 28688
rect 20864 28676 20870 28688
rect 20864 28648 21588 28676
rect 20864 28636 20870 28648
rect 13541 28611 13599 28617
rect 13541 28608 13553 28611
rect 13504 28580 13553 28608
rect 13504 28568 13510 28580
rect 13541 28577 13553 28580
rect 13587 28577 13599 28611
rect 13541 28571 13599 28577
rect 14185 28611 14243 28617
rect 14185 28577 14197 28611
rect 14231 28577 14243 28611
rect 15378 28608 15384 28620
rect 15339 28580 15384 28608
rect 14185 28571 14243 28577
rect 13188 28512 13400 28540
rect 13556 28540 13584 28571
rect 15378 28568 15384 28580
rect 15436 28568 15442 28620
rect 15746 28608 15752 28620
rect 15707 28580 15752 28608
rect 15746 28568 15752 28580
rect 15804 28568 15810 28620
rect 16206 28608 16212 28620
rect 16167 28580 16212 28608
rect 16206 28568 16212 28580
rect 16264 28568 16270 28620
rect 16942 28608 16948 28620
rect 16903 28580 16948 28608
rect 16942 28568 16948 28580
rect 17000 28568 17006 28620
rect 17678 28608 17684 28620
rect 17639 28580 17684 28608
rect 17678 28568 17684 28580
rect 17736 28568 17742 28620
rect 18233 28611 18291 28617
rect 18233 28577 18245 28611
rect 18279 28577 18291 28611
rect 18233 28571 18291 28577
rect 16114 28540 16120 28552
rect 13556 28512 16120 28540
rect 12952 28500 12958 28512
rect 16114 28500 16120 28512
rect 16172 28500 16178 28552
rect 18248 28540 18276 28571
rect 18322 28568 18328 28620
rect 18380 28608 18386 28620
rect 18509 28611 18567 28617
rect 18509 28608 18521 28611
rect 18380 28580 18521 28608
rect 18380 28568 18386 28580
rect 18509 28577 18521 28580
rect 18555 28577 18567 28611
rect 18509 28571 18567 28577
rect 19521 28611 19579 28617
rect 19521 28577 19533 28611
rect 19567 28608 19579 28611
rect 19886 28608 19892 28620
rect 19567 28580 19892 28608
rect 19567 28577 19579 28580
rect 19521 28571 19579 28577
rect 19886 28568 19892 28580
rect 19944 28568 19950 28620
rect 20073 28611 20131 28617
rect 20073 28577 20085 28611
rect 20119 28608 20131 28611
rect 20714 28608 20720 28620
rect 20119 28580 20720 28608
rect 20119 28577 20131 28580
rect 20073 28571 20131 28577
rect 20714 28568 20720 28580
rect 20772 28568 20778 28620
rect 20901 28611 20959 28617
rect 20901 28577 20913 28611
rect 20947 28608 20959 28611
rect 21082 28608 21088 28620
rect 20947 28580 21088 28608
rect 20947 28577 20959 28580
rect 20901 28571 20959 28577
rect 21082 28568 21088 28580
rect 21140 28568 21146 28620
rect 21560 28617 21588 28648
rect 21726 28636 21732 28688
rect 21784 28676 21790 28688
rect 25792 28676 25820 28716
rect 32306 28704 32312 28716
rect 32364 28704 32370 28756
rect 33502 28744 33508 28756
rect 32508 28716 33508 28744
rect 21784 28648 25820 28676
rect 21784 28636 21790 28648
rect 26050 28636 26056 28688
rect 26108 28676 26114 28688
rect 26108 28648 28212 28676
rect 26108 28636 26114 28648
rect 21545 28611 21603 28617
rect 21545 28577 21557 28611
rect 21591 28577 21603 28611
rect 22186 28608 22192 28620
rect 22147 28580 22192 28608
rect 21545 28571 21603 28577
rect 22186 28568 22192 28580
rect 22244 28568 22250 28620
rect 23014 28608 23020 28620
rect 22975 28580 23020 28608
rect 23014 28568 23020 28580
rect 23072 28568 23078 28620
rect 23569 28611 23627 28617
rect 23569 28577 23581 28611
rect 23615 28577 23627 28611
rect 23569 28571 23627 28577
rect 18414 28540 18420 28552
rect 18248 28512 18420 28540
rect 18414 28500 18420 28512
rect 18472 28500 18478 28552
rect 18785 28543 18843 28549
rect 18785 28509 18797 28543
rect 18831 28540 18843 28543
rect 19426 28540 19432 28552
rect 18831 28512 19432 28540
rect 18831 28509 18843 28512
rect 18785 28503 18843 28509
rect 19426 28500 19432 28512
rect 19484 28500 19490 28552
rect 20165 28543 20223 28549
rect 20165 28509 20177 28543
rect 20211 28540 20223 28543
rect 20254 28540 20260 28552
rect 20211 28512 20260 28540
rect 20211 28509 20223 28512
rect 20165 28503 20223 28509
rect 20254 28500 20260 28512
rect 20312 28500 20318 28552
rect 23477 28543 23535 28549
rect 23477 28509 23489 28543
rect 23523 28509 23535 28543
rect 23584 28540 23612 28571
rect 23658 28568 23664 28620
rect 23716 28608 23722 28620
rect 24854 28608 24860 28620
rect 23716 28580 23761 28608
rect 24815 28580 24860 28608
rect 23716 28568 23722 28580
rect 24854 28568 24860 28580
rect 24912 28568 24918 28620
rect 24946 28568 24952 28620
rect 25004 28608 25010 28620
rect 25314 28608 25320 28620
rect 25004 28580 25049 28608
rect 25275 28580 25320 28608
rect 25004 28568 25010 28580
rect 25314 28568 25320 28580
rect 25372 28568 25378 28620
rect 26510 28608 26516 28620
rect 26471 28580 26516 28608
rect 26510 28568 26516 28580
rect 26568 28568 26574 28620
rect 28184 28617 28212 28648
rect 29362 28636 29368 28688
rect 29420 28676 29426 28688
rect 32508 28685 32536 28716
rect 33502 28704 33508 28716
rect 33560 28704 33566 28756
rect 33597 28747 33655 28753
rect 33597 28713 33609 28747
rect 33643 28744 33655 28747
rect 34146 28744 34152 28756
rect 33643 28716 34152 28744
rect 33643 28713 33655 28716
rect 33597 28707 33655 28713
rect 34146 28704 34152 28716
rect 34204 28704 34210 28756
rect 37642 28744 37648 28756
rect 36464 28716 37648 28744
rect 32493 28679 32551 28685
rect 32493 28676 32505 28679
rect 29420 28648 32505 28676
rect 29420 28636 29426 28648
rect 32493 28645 32505 28648
rect 32539 28645 32551 28679
rect 32493 28639 32551 28645
rect 33045 28679 33103 28685
rect 33045 28645 33057 28679
rect 33091 28676 33103 28679
rect 33134 28676 33140 28688
rect 33091 28648 33140 28676
rect 33091 28645 33103 28648
rect 33045 28639 33103 28645
rect 33134 28636 33140 28648
rect 33192 28636 33198 28688
rect 33520 28676 33548 28704
rect 35161 28679 35219 28685
rect 35161 28676 35173 28679
rect 33520 28648 35173 28676
rect 35161 28645 35173 28648
rect 35207 28645 35219 28679
rect 35161 28639 35219 28645
rect 36464 28620 36492 28716
rect 37642 28704 37648 28716
rect 37700 28744 37706 28756
rect 37921 28747 37979 28753
rect 37921 28744 37933 28747
rect 37700 28716 37933 28744
rect 37700 28704 37706 28716
rect 37921 28713 37933 28716
rect 37967 28713 37979 28747
rect 37921 28707 37979 28713
rect 27065 28611 27123 28617
rect 27065 28608 27077 28611
rect 26620 28580 27077 28608
rect 24872 28540 24900 28568
rect 23584 28512 24900 28540
rect 25777 28543 25835 28549
rect 23477 28503 23535 28509
rect 25777 28509 25789 28543
rect 25823 28540 25835 28543
rect 26620 28540 26648 28580
rect 27065 28577 27077 28580
rect 27111 28577 27123 28611
rect 27065 28571 27123 28577
rect 27709 28611 27767 28617
rect 27709 28577 27721 28611
rect 27755 28577 27767 28611
rect 27709 28571 27767 28577
rect 28169 28611 28227 28617
rect 28169 28577 28181 28611
rect 28215 28577 28227 28611
rect 28169 28571 28227 28577
rect 29181 28611 29239 28617
rect 29181 28577 29193 28611
rect 29227 28608 29239 28611
rect 29270 28608 29276 28620
rect 29227 28580 29276 28608
rect 29227 28577 29239 28580
rect 29181 28571 29239 28577
rect 26878 28540 26884 28552
rect 25823 28512 26648 28540
rect 26839 28512 26884 28540
rect 25823 28509 25835 28512
rect 25777 28503 25835 28509
rect 2406 28432 2412 28484
rect 2464 28472 2470 28484
rect 4893 28475 4951 28481
rect 4893 28472 4905 28475
rect 2464 28444 4905 28472
rect 2464 28432 2470 28444
rect 4893 28441 4905 28444
rect 4939 28441 4951 28475
rect 5718 28472 5724 28484
rect 5679 28444 5724 28472
rect 4893 28435 4951 28441
rect 5718 28432 5724 28444
rect 5776 28432 5782 28484
rect 12158 28432 12164 28484
rect 12216 28472 12222 28484
rect 13449 28475 13507 28481
rect 13449 28472 13461 28475
rect 12216 28444 13461 28472
rect 12216 28432 12222 28444
rect 13449 28441 13461 28444
rect 13495 28441 13507 28475
rect 23492 28472 23520 28503
rect 26878 28500 26884 28512
rect 26936 28500 26942 28552
rect 26970 28500 26976 28552
rect 27028 28540 27034 28552
rect 27724 28540 27752 28571
rect 29270 28568 29276 28580
rect 29328 28568 29334 28620
rect 29638 28608 29644 28620
rect 29599 28580 29644 28608
rect 29638 28568 29644 28580
rect 29696 28568 29702 28620
rect 30650 28608 30656 28620
rect 30611 28580 30656 28608
rect 30650 28568 30656 28580
rect 30708 28568 30714 28620
rect 31205 28611 31263 28617
rect 31205 28577 31217 28611
rect 31251 28608 31263 28611
rect 32398 28608 32404 28620
rect 31251 28580 32404 28608
rect 31251 28577 31263 28580
rect 31205 28571 31263 28577
rect 32398 28568 32404 28580
rect 32456 28568 32462 28620
rect 32677 28611 32735 28617
rect 32677 28577 32689 28611
rect 32723 28577 32735 28611
rect 32677 28571 32735 28577
rect 27028 28512 27752 28540
rect 27028 28500 27034 28512
rect 27890 28500 27896 28552
rect 27948 28540 27954 28552
rect 28261 28543 28319 28549
rect 28261 28540 28273 28543
rect 27948 28512 28273 28540
rect 27948 28500 27954 28512
rect 28261 28509 28273 28512
rect 28307 28509 28319 28543
rect 31478 28540 31484 28552
rect 31439 28512 31484 28540
rect 28261 28503 28319 28509
rect 31478 28500 31484 28512
rect 31536 28500 31542 28552
rect 32692 28540 32720 28571
rect 32766 28568 32772 28620
rect 32824 28608 32830 28620
rect 33505 28611 33563 28617
rect 33505 28608 33517 28611
rect 32824 28580 33517 28608
rect 32824 28568 32830 28580
rect 33505 28577 33517 28580
rect 33551 28577 33563 28611
rect 34238 28608 34244 28620
rect 34199 28580 34244 28608
rect 33505 28571 33563 28577
rect 34238 28568 34244 28580
rect 34296 28568 34302 28620
rect 35069 28611 35127 28617
rect 35069 28577 35081 28611
rect 35115 28577 35127 28611
rect 35069 28571 35127 28577
rect 33778 28540 33784 28552
rect 32692 28512 33784 28540
rect 33778 28500 33784 28512
rect 33836 28500 33842 28552
rect 34333 28543 34391 28549
rect 34333 28509 34345 28543
rect 34379 28509 34391 28543
rect 35084 28540 35112 28571
rect 35526 28568 35532 28620
rect 35584 28608 35590 28620
rect 35713 28611 35771 28617
rect 35713 28608 35725 28611
rect 35584 28580 35725 28608
rect 35584 28568 35590 28580
rect 35713 28577 35725 28580
rect 35759 28577 35771 28611
rect 36354 28608 36360 28620
rect 36315 28580 36360 28608
rect 35713 28571 35771 28577
rect 36354 28568 36360 28580
rect 36412 28568 36418 28620
rect 36446 28568 36452 28620
rect 36504 28608 36510 28620
rect 37185 28611 37243 28617
rect 36504 28580 36549 28608
rect 36504 28568 36510 28580
rect 37185 28577 37197 28611
rect 37231 28608 37243 28611
rect 37642 28608 37648 28620
rect 37231 28580 37648 28608
rect 37231 28577 37243 28580
rect 37185 28571 37243 28577
rect 37642 28568 37648 28580
rect 37700 28568 37706 28620
rect 37737 28611 37795 28617
rect 37737 28577 37749 28611
rect 37783 28577 37795 28611
rect 37737 28571 37795 28577
rect 36538 28540 36544 28552
rect 35084 28512 36544 28540
rect 34333 28503 34391 28509
rect 28534 28472 28540 28484
rect 23492 28444 28540 28472
rect 13449 28435 13507 28441
rect 28534 28432 28540 28444
rect 28592 28432 28598 28484
rect 28994 28472 29000 28484
rect 28955 28444 29000 28472
rect 28994 28432 29000 28444
rect 29052 28432 29058 28484
rect 30558 28472 30564 28484
rect 30519 28444 30564 28472
rect 30558 28432 30564 28444
rect 30616 28432 30622 28484
rect 32030 28432 32036 28484
rect 32088 28472 32094 28484
rect 34348 28472 34376 28503
rect 36538 28500 36544 28512
rect 36596 28540 36602 28552
rect 37752 28540 37780 28571
rect 36596 28512 37780 28540
rect 36596 28500 36602 28512
rect 32088 28444 34376 28472
rect 32088 28432 32094 28444
rect 2958 28404 2964 28416
rect 2919 28376 2964 28404
rect 2958 28364 2964 28376
rect 3016 28364 3022 28416
rect 8202 28364 8208 28416
rect 8260 28404 8266 28416
rect 8573 28407 8631 28413
rect 8573 28404 8585 28407
rect 8260 28376 8585 28404
rect 8260 28364 8266 28376
rect 8573 28373 8585 28376
rect 8619 28373 8631 28407
rect 8573 28367 8631 28373
rect 37093 28407 37151 28413
rect 37093 28373 37105 28407
rect 37139 28404 37151 28407
rect 37182 28404 37188 28416
rect 37139 28376 37188 28404
rect 37139 28373 37151 28376
rect 37093 28367 37151 28373
rect 37182 28364 37188 28376
rect 37240 28364 37246 28416
rect 1104 28314 38824 28336
rect 1104 28262 4246 28314
rect 4298 28262 4310 28314
rect 4362 28262 4374 28314
rect 4426 28262 4438 28314
rect 4490 28262 34966 28314
rect 35018 28262 35030 28314
rect 35082 28262 35094 28314
rect 35146 28262 35158 28314
rect 35210 28262 38824 28314
rect 1104 28240 38824 28262
rect 1854 28200 1860 28212
rect 1815 28172 1860 28200
rect 1854 28160 1860 28172
rect 1912 28160 1918 28212
rect 4341 28203 4399 28209
rect 4341 28169 4353 28203
rect 4387 28200 4399 28203
rect 4706 28200 4712 28212
rect 4387 28172 4712 28200
rect 4387 28169 4399 28172
rect 4341 28163 4399 28169
rect 4706 28160 4712 28172
rect 4764 28160 4770 28212
rect 8202 28160 8208 28212
rect 8260 28200 8266 28212
rect 8260 28172 14320 28200
rect 8260 28160 8266 28172
rect 3326 28132 3332 28144
rect 3287 28104 3332 28132
rect 3326 28092 3332 28104
rect 3384 28092 3390 28144
rect 5810 28132 5816 28144
rect 5771 28104 5816 28132
rect 5810 28092 5816 28104
rect 5868 28092 5874 28144
rect 7926 28132 7932 28144
rect 7024 28104 7932 28132
rect 2958 28024 2964 28076
rect 3016 28064 3022 28076
rect 5169 28067 5227 28073
rect 3016 28036 4200 28064
rect 3016 28024 3022 28036
rect 1765 27999 1823 28005
rect 1765 27965 1777 27999
rect 1811 27996 1823 27999
rect 2406 27996 2412 28008
rect 1811 27968 2412 27996
rect 1811 27965 1823 27968
rect 1765 27959 1823 27965
rect 2406 27956 2412 27968
rect 2464 27956 2470 28008
rect 2774 27956 2780 28008
rect 2832 27996 2838 28008
rect 3234 27996 3240 28008
rect 2832 27968 2877 27996
rect 3195 27968 3240 27996
rect 2832 27956 2838 27968
rect 3234 27956 3240 27968
rect 3292 27956 3298 28008
rect 3421 27999 3479 28005
rect 3421 27965 3433 27999
rect 3467 27996 3479 27999
rect 4062 27996 4068 28008
rect 3467 27968 4068 27996
rect 3467 27965 3479 27968
rect 3421 27959 3479 27965
rect 4062 27956 4068 27968
rect 4120 27956 4126 28008
rect 4172 28005 4200 28036
rect 5169 28033 5181 28067
rect 5215 28064 5227 28067
rect 5442 28064 5448 28076
rect 5215 28036 5448 28064
rect 5215 28033 5227 28036
rect 5169 28027 5227 28033
rect 5442 28024 5448 28036
rect 5500 28024 5506 28076
rect 4157 27999 4215 28005
rect 4157 27965 4169 27999
rect 4203 27965 4215 27999
rect 5350 27996 5356 28008
rect 5311 27968 5356 27996
rect 4157 27959 4215 27965
rect 5350 27956 5356 27968
rect 5408 27956 5414 28008
rect 5905 27999 5963 28005
rect 5905 27965 5917 27999
rect 5951 27996 5963 27999
rect 6362 27996 6368 28008
rect 5951 27968 6368 27996
rect 5951 27965 5963 27968
rect 5905 27959 5963 27965
rect 6362 27956 6368 27968
rect 6420 27956 6426 28008
rect 6914 27956 6920 28008
rect 6972 27996 6978 28008
rect 7024 28005 7052 28104
rect 7926 28092 7932 28104
rect 7984 28092 7990 28144
rect 8662 28132 8668 28144
rect 8623 28104 8668 28132
rect 8662 28092 8668 28104
rect 8720 28092 8726 28144
rect 9582 28132 9588 28144
rect 9324 28104 9588 28132
rect 7009 27999 7067 28005
rect 7009 27996 7021 27999
rect 6972 27968 7021 27996
rect 6972 27956 6978 27968
rect 7009 27965 7021 27968
rect 7055 27965 7067 27999
rect 7009 27959 7067 27965
rect 7745 27999 7803 28005
rect 7745 27965 7757 27999
rect 7791 27996 7803 27999
rect 8478 27996 8484 28008
rect 7791 27968 8484 27996
rect 7791 27965 7803 27968
rect 7745 27959 7803 27965
rect 8478 27956 8484 27968
rect 8536 27956 8542 28008
rect 8846 27996 8852 28008
rect 8807 27968 8852 27996
rect 8846 27956 8852 27968
rect 8904 27956 8910 28008
rect 9324 28005 9352 28104
rect 9582 28092 9588 28104
rect 9640 28092 9646 28144
rect 9674 28092 9680 28144
rect 9732 28132 9738 28144
rect 9732 28104 11652 28132
rect 9732 28092 9738 28104
rect 9950 28064 9956 28076
rect 9911 28036 9956 28064
rect 9950 28024 9956 28036
rect 10008 28024 10014 28076
rect 10594 28064 10600 28076
rect 10555 28036 10600 28064
rect 10594 28024 10600 28036
rect 10652 28024 10658 28076
rect 11149 28067 11207 28073
rect 11149 28033 11161 28067
rect 11195 28064 11207 28067
rect 11330 28064 11336 28076
rect 11195 28036 11336 28064
rect 11195 28033 11207 28036
rect 11149 28027 11207 28033
rect 11330 28024 11336 28036
rect 11388 28064 11394 28076
rect 11624 28073 11652 28104
rect 12434 28092 12440 28144
rect 12492 28132 12498 28144
rect 12529 28135 12587 28141
rect 12529 28132 12541 28135
rect 12492 28104 12541 28132
rect 12492 28092 12498 28104
rect 12529 28101 12541 28104
rect 12575 28101 12587 28135
rect 14292 28132 14320 28172
rect 14366 28160 14372 28212
rect 14424 28200 14430 28212
rect 17037 28203 17095 28209
rect 17037 28200 17049 28203
rect 14424 28172 17049 28200
rect 14424 28160 14430 28172
rect 15286 28132 15292 28144
rect 14292 28104 15292 28132
rect 12529 28095 12587 28101
rect 15286 28092 15292 28104
rect 15344 28092 15350 28144
rect 11609 28067 11667 28073
rect 11388 28036 11560 28064
rect 11388 28024 11394 28036
rect 9217 27999 9275 28005
rect 9217 27965 9229 27999
rect 9263 27965 9275 27999
rect 9217 27959 9275 27965
rect 9309 27999 9367 28005
rect 9309 27965 9321 27999
rect 9355 27965 9367 27999
rect 9766 27996 9772 28008
rect 9727 27968 9772 27996
rect 9309 27959 9367 27965
rect 9232 27928 9260 27959
rect 9766 27956 9772 27968
rect 9824 27956 9830 28008
rect 11422 27996 11428 28008
rect 11383 27968 11428 27996
rect 11422 27956 11428 27968
rect 11480 27956 11486 28008
rect 11532 27996 11560 28036
rect 11609 28033 11621 28067
rect 11655 28064 11667 28067
rect 14553 28067 14611 28073
rect 14553 28064 14565 28067
rect 11655 28036 14565 28064
rect 11655 28033 11667 28036
rect 11609 28027 11667 28033
rect 12066 27996 12072 28008
rect 11532 27968 12072 27996
rect 12066 27956 12072 27968
rect 12124 27956 12130 28008
rect 13188 28005 13216 28036
rect 14553 28033 14565 28036
rect 14599 28033 14611 28067
rect 14553 28027 14611 28033
rect 12529 27999 12587 28005
rect 12529 27965 12541 27999
rect 12575 27965 12587 27999
rect 12529 27959 12587 27965
rect 13173 27999 13231 28005
rect 13173 27965 13185 27999
rect 13219 27965 13231 27999
rect 13173 27959 13231 27965
rect 13725 27999 13783 28005
rect 13725 27965 13737 27999
rect 13771 27965 13783 27999
rect 13725 27959 13783 27965
rect 9232 27900 9352 27928
rect 7193 27863 7251 27869
rect 7193 27829 7205 27863
rect 7239 27860 7251 27863
rect 7558 27860 7564 27872
rect 7239 27832 7564 27860
rect 7239 27829 7251 27832
rect 7193 27823 7251 27829
rect 7558 27820 7564 27832
rect 7616 27820 7622 27872
rect 9324 27860 9352 27900
rect 11054 27860 11060 27872
rect 9324 27832 11060 27860
rect 11054 27820 11060 27832
rect 11112 27860 11118 27872
rect 12544 27860 12572 27959
rect 13740 27928 13768 27959
rect 13814 27956 13820 28008
rect 13872 27996 13878 28008
rect 15488 28005 15516 28172
rect 17037 28169 17049 28172
rect 17083 28200 17095 28203
rect 17126 28200 17132 28212
rect 17083 28172 17132 28200
rect 17083 28169 17095 28172
rect 17037 28163 17095 28169
rect 17126 28160 17132 28172
rect 17184 28160 17190 28212
rect 23014 28200 23020 28212
rect 22975 28172 23020 28200
rect 23014 28160 23020 28172
rect 23072 28160 23078 28212
rect 31849 28203 31907 28209
rect 31849 28169 31861 28203
rect 31895 28200 31907 28203
rect 31938 28200 31944 28212
rect 31895 28172 31944 28200
rect 31895 28169 31907 28172
rect 31849 28163 31907 28169
rect 31938 28160 31944 28172
rect 31996 28160 32002 28212
rect 32306 28160 32312 28212
rect 32364 28200 32370 28212
rect 32364 28172 33364 28200
rect 32364 28160 32370 28172
rect 15565 28135 15623 28141
rect 15565 28101 15577 28135
rect 15611 28132 15623 28135
rect 16206 28132 16212 28144
rect 15611 28104 16212 28132
rect 15611 28101 15623 28104
rect 15565 28095 15623 28101
rect 16206 28092 16212 28104
rect 16264 28092 16270 28144
rect 18322 28132 18328 28144
rect 18283 28104 18328 28132
rect 18322 28092 18328 28104
rect 18380 28092 18386 28144
rect 22649 28135 22707 28141
rect 22649 28101 22661 28135
rect 22695 28132 22707 28135
rect 23566 28132 23572 28144
rect 22695 28104 23572 28132
rect 22695 28101 22707 28104
rect 22649 28095 22707 28101
rect 23566 28092 23572 28104
rect 23624 28092 23630 28144
rect 24854 28092 24860 28144
rect 24912 28132 24918 28144
rect 25501 28135 25559 28141
rect 25501 28132 25513 28135
rect 24912 28104 25513 28132
rect 24912 28092 24918 28104
rect 25501 28101 25513 28104
rect 25547 28101 25559 28135
rect 25501 28095 25559 28101
rect 16114 28064 16120 28076
rect 16075 28036 16120 28064
rect 16114 28024 16120 28036
rect 16172 28024 16178 28076
rect 17678 28024 17684 28076
rect 17736 28064 17742 28076
rect 18877 28067 18935 28073
rect 18877 28064 18889 28067
rect 17736 28036 18889 28064
rect 17736 28024 17742 28036
rect 18877 28033 18889 28036
rect 18923 28033 18935 28067
rect 20622 28064 20628 28076
rect 18877 28027 18935 28033
rect 20272 28036 20628 28064
rect 14461 27999 14519 28005
rect 14461 27996 14473 27999
rect 13872 27968 14473 27996
rect 13872 27956 13878 27968
rect 14461 27965 14473 27968
rect 14507 27965 14519 27999
rect 14461 27959 14519 27965
rect 15473 27999 15531 28005
rect 15473 27965 15485 27999
rect 15519 27965 15531 27999
rect 15930 27996 15936 28008
rect 15891 27968 15936 27996
rect 15473 27959 15531 27965
rect 14366 27928 14372 27940
rect 13740 27900 14372 27928
rect 14366 27888 14372 27900
rect 14424 27888 14430 27940
rect 14476 27928 14504 27959
rect 15930 27956 15936 27968
rect 15988 27956 15994 28008
rect 16853 27999 16911 28005
rect 16853 27965 16865 27999
rect 16899 27996 16911 27999
rect 17494 27996 17500 28008
rect 16899 27968 17500 27996
rect 16899 27965 16911 27968
rect 16853 27959 16911 27965
rect 17494 27956 17500 27968
rect 17552 27956 17558 28008
rect 18046 27996 18052 28008
rect 18007 27968 18052 27996
rect 18046 27956 18052 27968
rect 18104 27956 18110 28008
rect 18414 27956 18420 28008
rect 18472 27996 18478 28008
rect 20272 28005 20300 28036
rect 20622 28024 20628 28036
rect 20680 28024 20686 28076
rect 22002 28024 22008 28076
rect 22060 28064 22066 28076
rect 22741 28067 22799 28073
rect 22741 28064 22753 28067
rect 22060 28036 22753 28064
rect 22060 28024 22066 28036
rect 22741 28033 22753 28036
rect 22787 28033 22799 28067
rect 26878 28064 26884 28076
rect 26839 28036 26884 28064
rect 22741 28027 22799 28033
rect 26878 28024 26884 28036
rect 26936 28024 26942 28076
rect 31956 28064 31984 28160
rect 32398 28092 32404 28144
rect 32456 28132 32462 28144
rect 33229 28135 33287 28141
rect 33229 28132 33241 28135
rect 32456 28104 33241 28132
rect 32456 28092 32462 28104
rect 33229 28101 33241 28104
rect 33275 28101 33287 28135
rect 33336 28132 33364 28172
rect 33410 28160 33416 28212
rect 33468 28200 33474 28212
rect 34149 28203 34207 28209
rect 34149 28200 34161 28203
rect 33468 28172 34161 28200
rect 33468 28160 33474 28172
rect 34149 28169 34161 28172
rect 34195 28169 34207 28203
rect 34149 28163 34207 28169
rect 34514 28160 34520 28212
rect 34572 28200 34578 28212
rect 35161 28203 35219 28209
rect 35161 28200 35173 28203
rect 34572 28172 35173 28200
rect 34572 28160 34578 28172
rect 35161 28169 35173 28172
rect 35207 28169 35219 28203
rect 37918 28200 37924 28212
rect 37879 28172 37924 28200
rect 35161 28163 35219 28169
rect 37918 28160 37924 28172
rect 37976 28160 37982 28212
rect 33336 28104 37780 28132
rect 33229 28095 33287 28101
rect 32493 28067 32551 28073
rect 32493 28064 32505 28067
rect 31956 28036 32505 28064
rect 32493 28033 32505 28036
rect 32539 28033 32551 28067
rect 36446 28064 36452 28076
rect 32493 28027 32551 28033
rect 32876 28036 36452 28064
rect 32876 28008 32904 28036
rect 18601 27999 18659 28005
rect 18601 27996 18613 27999
rect 18472 27968 18613 27996
rect 18472 27956 18478 27968
rect 18601 27965 18613 27968
rect 18647 27965 18659 27999
rect 18601 27959 18659 27965
rect 20257 27999 20315 28005
rect 20257 27965 20269 27999
rect 20303 27965 20315 27999
rect 20257 27959 20315 27965
rect 20533 27999 20591 28005
rect 20533 27965 20545 27999
rect 20579 27965 20591 27999
rect 21174 27996 21180 28008
rect 21135 27968 21180 27996
rect 20533 27959 20591 27965
rect 14918 27928 14924 27940
rect 14476 27900 14924 27928
rect 14918 27888 14924 27900
rect 14976 27928 14982 27940
rect 15948 27928 15976 27956
rect 14976 27900 15976 27928
rect 20548 27928 20576 27959
rect 21174 27956 21180 27968
rect 21232 27956 21238 28008
rect 22520 27999 22578 28005
rect 22520 27965 22532 27999
rect 22566 27996 22578 27999
rect 23290 27996 23296 28008
rect 22566 27968 23296 27996
rect 22566 27965 22578 27968
rect 22520 27959 22578 27965
rect 23290 27956 23296 27968
rect 23348 27956 23354 28008
rect 24397 27999 24455 28005
rect 24397 27965 24409 27999
rect 24443 27965 24455 27999
rect 24670 27996 24676 28008
rect 24631 27968 24676 27996
rect 24397 27959 24455 27965
rect 20990 27928 20996 27940
rect 20548 27900 20996 27928
rect 14976 27888 14982 27900
rect 20990 27888 20996 27900
rect 21048 27928 21054 27940
rect 21450 27928 21456 27940
rect 21048 27900 21456 27928
rect 21048 27888 21054 27900
rect 21450 27888 21456 27900
rect 21508 27888 21514 27940
rect 22373 27931 22431 27937
rect 22373 27897 22385 27931
rect 22419 27928 22431 27931
rect 22738 27928 22744 27940
rect 22419 27900 22744 27928
rect 22419 27897 22431 27900
rect 22373 27891 22431 27897
rect 22738 27888 22744 27900
rect 22796 27888 22802 27940
rect 24412 27928 24440 27959
rect 24670 27956 24676 27968
rect 24728 27956 24734 28008
rect 25130 27996 25136 28008
rect 25091 27968 25136 27996
rect 25130 27956 25136 27968
rect 25188 27956 25194 28008
rect 25501 27999 25559 28005
rect 25501 27965 25513 27999
rect 25547 27996 25559 27999
rect 26050 27996 26056 28008
rect 25547 27968 26056 27996
rect 25547 27965 25559 27968
rect 25501 27959 25559 27965
rect 26050 27956 26056 27968
rect 26108 27956 26114 28008
rect 26418 27956 26424 28008
rect 26476 27996 26482 28008
rect 26513 27999 26571 28005
rect 26513 27996 26525 27999
rect 26476 27968 26525 27996
rect 26476 27956 26482 27968
rect 26513 27965 26525 27968
rect 26559 27965 26571 27999
rect 26513 27959 26571 27965
rect 26605 27999 26663 28005
rect 26605 27965 26617 27999
rect 26651 27965 26663 27999
rect 26605 27959 26663 27965
rect 29273 27999 29331 28005
rect 29273 27965 29285 27999
rect 29319 27996 29331 27999
rect 29362 27996 29368 28008
rect 29319 27968 29368 27996
rect 29319 27965 29331 27968
rect 29273 27959 29331 27965
rect 26234 27928 26240 27940
rect 24412 27900 26240 27928
rect 26234 27888 26240 27900
rect 26292 27888 26298 27940
rect 11112 27832 12572 27860
rect 13817 27863 13875 27869
rect 11112 27820 11118 27832
rect 13817 27829 13829 27863
rect 13863 27860 13875 27863
rect 14458 27860 14464 27872
rect 13863 27832 14464 27860
rect 13863 27829 13875 27832
rect 13817 27823 13875 27829
rect 14458 27820 14464 27832
rect 14516 27820 14522 27872
rect 15286 27820 15292 27872
rect 15344 27860 15350 27872
rect 17402 27860 17408 27872
rect 15344 27832 17408 27860
rect 15344 27820 15350 27832
rect 17402 27820 17408 27832
rect 17460 27820 17466 27872
rect 20254 27860 20260 27872
rect 20215 27832 20260 27860
rect 20254 27820 20260 27832
rect 20312 27820 20318 27872
rect 21269 27863 21327 27869
rect 21269 27829 21281 27863
rect 21315 27860 21327 27863
rect 21542 27860 21548 27872
rect 21315 27832 21548 27860
rect 21315 27829 21327 27832
rect 21269 27823 21327 27829
rect 21542 27820 21548 27832
rect 21600 27820 21606 27872
rect 26329 27863 26387 27869
rect 26329 27829 26341 27863
rect 26375 27860 26387 27863
rect 26620 27860 26648 27959
rect 29362 27956 29368 27968
rect 29420 27956 29426 28008
rect 29457 27999 29515 28005
rect 29457 27965 29469 27999
rect 29503 27996 29515 27999
rect 30190 27996 30196 28008
rect 29503 27968 30196 27996
rect 29503 27965 29515 27968
rect 29457 27959 29515 27965
rect 30190 27956 30196 27968
rect 30248 27956 30254 28008
rect 30282 27956 30288 28008
rect 30340 27996 30346 28008
rect 30340 27968 30385 27996
rect 30340 27956 30346 27968
rect 30558 27956 30564 28008
rect 30616 27996 30622 28008
rect 32858 27996 32864 28008
rect 30616 27968 30661 27996
rect 32819 27968 32864 27996
rect 30616 27956 30622 27968
rect 32858 27956 32864 27968
rect 32916 27956 32922 28008
rect 33229 27999 33287 28005
rect 33229 27965 33241 27999
rect 33275 27965 33287 27999
rect 33229 27959 33287 27965
rect 28258 27928 28264 27940
rect 28219 27900 28264 27928
rect 28258 27888 28264 27900
rect 28316 27888 28322 27940
rect 29825 27931 29883 27937
rect 29825 27897 29837 27931
rect 29871 27897 29883 27931
rect 29825 27891 29883 27897
rect 27338 27860 27344 27872
rect 26375 27832 27344 27860
rect 26375 27829 26387 27832
rect 26329 27823 26387 27829
rect 27338 27820 27344 27832
rect 27396 27820 27402 27872
rect 29840 27860 29868 27891
rect 33244 27860 33272 27959
rect 33502 27956 33508 28008
rect 33560 27996 33566 28008
rect 34900 28005 34928 28036
rect 36446 28024 36452 28036
rect 36504 28024 36510 28076
rect 37090 28064 37096 28076
rect 37051 28036 37096 28064
rect 37090 28024 37096 28036
rect 37148 28024 37154 28076
rect 33965 27999 34023 28005
rect 33965 27996 33977 27999
rect 33560 27968 33977 27996
rect 33560 27956 33566 27968
rect 33965 27965 33977 27968
rect 34011 27965 34023 27999
rect 33965 27959 34023 27965
rect 34885 27999 34943 28005
rect 34885 27965 34897 27999
rect 34931 27965 34943 27999
rect 34885 27959 34943 27965
rect 35069 27999 35127 28005
rect 35069 27965 35081 27999
rect 35115 27996 35127 27999
rect 35250 27996 35256 28008
rect 35115 27968 35256 27996
rect 35115 27965 35127 27968
rect 35069 27959 35127 27965
rect 35250 27956 35256 27968
rect 35308 27956 35314 28008
rect 35526 27956 35532 28008
rect 35584 27996 35590 28008
rect 35989 27999 36047 28005
rect 35989 27996 36001 27999
rect 35584 27968 36001 27996
rect 35584 27956 35590 27968
rect 35989 27965 36001 27968
rect 36035 27965 36047 27999
rect 35989 27959 36047 27965
rect 36354 27956 36360 28008
rect 36412 27996 36418 28008
rect 36633 27999 36691 28005
rect 36633 27996 36645 27999
rect 36412 27968 36645 27996
rect 36412 27956 36418 27968
rect 36633 27965 36645 27968
rect 36679 27965 36691 27999
rect 36633 27959 36691 27965
rect 36648 27928 36676 27959
rect 36722 27956 36728 28008
rect 36780 27996 36786 28008
rect 37752 28005 37780 28104
rect 37737 27999 37795 28005
rect 36780 27968 36825 27996
rect 36780 27956 36786 27968
rect 37737 27965 37749 27999
rect 37783 27965 37795 27999
rect 37737 27959 37795 27965
rect 36998 27928 37004 27940
rect 36648 27900 37004 27928
rect 36998 27888 37004 27900
rect 37056 27888 37062 27940
rect 29840 27832 33272 27860
rect 1104 27770 38824 27792
rect 1104 27718 19606 27770
rect 19658 27718 19670 27770
rect 19722 27718 19734 27770
rect 19786 27718 19798 27770
rect 19850 27718 38824 27770
rect 1104 27696 38824 27718
rect 4249 27659 4307 27665
rect 4249 27625 4261 27659
rect 4295 27656 4307 27659
rect 4890 27656 4896 27668
rect 4295 27628 4896 27656
rect 4295 27625 4307 27628
rect 4249 27619 4307 27625
rect 4890 27616 4896 27628
rect 4948 27656 4954 27668
rect 5258 27656 5264 27668
rect 4948 27628 5264 27656
rect 4948 27616 4954 27628
rect 5258 27616 5264 27628
rect 5316 27616 5322 27668
rect 11146 27616 11152 27668
rect 11204 27656 11210 27668
rect 11425 27659 11483 27665
rect 11425 27656 11437 27659
rect 11204 27628 11437 27656
rect 11204 27616 11210 27628
rect 11425 27625 11437 27628
rect 11471 27625 11483 27659
rect 11425 27619 11483 27625
rect 14274 27616 14280 27668
rect 14332 27656 14338 27668
rect 15102 27656 15108 27668
rect 14332 27628 15108 27656
rect 14332 27616 14338 27628
rect 15102 27616 15108 27628
rect 15160 27616 15166 27668
rect 30098 27616 30104 27668
rect 30156 27656 30162 27668
rect 36630 27656 36636 27668
rect 30156 27628 36636 27656
rect 30156 27616 30162 27628
rect 36630 27616 36636 27628
rect 36688 27616 36694 27668
rect 6822 27588 6828 27600
rect 6783 27560 6828 27588
rect 6822 27548 6828 27560
rect 6880 27548 6886 27600
rect 8938 27588 8944 27600
rect 8899 27560 8944 27588
rect 8938 27548 8944 27560
rect 8996 27548 9002 27600
rect 12618 27588 12624 27600
rect 11624 27560 12624 27588
rect 2682 27520 2688 27532
rect 2643 27492 2688 27520
rect 2682 27480 2688 27492
rect 2740 27480 2746 27532
rect 3053 27523 3111 27529
rect 3053 27489 3065 27523
rect 3099 27520 3111 27523
rect 3234 27520 3240 27532
rect 3099 27492 3240 27520
rect 3099 27489 3111 27492
rect 3053 27483 3111 27489
rect 3234 27480 3240 27492
rect 3292 27480 3298 27532
rect 4062 27520 4068 27532
rect 4023 27492 4068 27520
rect 4062 27480 4068 27492
rect 4120 27480 4126 27532
rect 4982 27520 4988 27532
rect 4943 27492 4988 27520
rect 4982 27480 4988 27492
rect 5040 27480 5046 27532
rect 5445 27523 5503 27529
rect 5445 27489 5457 27523
rect 5491 27520 5503 27523
rect 5718 27520 5724 27532
rect 5491 27492 5724 27520
rect 5491 27489 5503 27492
rect 5445 27483 5503 27489
rect 5718 27480 5724 27492
rect 5776 27480 5782 27532
rect 7469 27523 7527 27529
rect 7469 27489 7481 27523
rect 7515 27520 7527 27523
rect 7650 27520 7656 27532
rect 7515 27492 7656 27520
rect 7515 27489 7527 27492
rect 7469 27483 7527 27489
rect 7650 27480 7656 27492
rect 7708 27480 7714 27532
rect 7745 27523 7803 27529
rect 7745 27489 7757 27523
rect 7791 27489 7803 27523
rect 8110 27520 8116 27532
rect 8071 27492 8116 27520
rect 7745 27483 7803 27489
rect 1486 27412 1492 27464
rect 1544 27452 1550 27464
rect 2225 27455 2283 27461
rect 2225 27452 2237 27455
rect 1544 27424 2237 27452
rect 1544 27412 1550 27424
rect 2225 27421 2237 27424
rect 2271 27421 2283 27455
rect 3142 27452 3148 27464
rect 3103 27424 3148 27452
rect 2225 27415 2283 27421
rect 3142 27412 3148 27424
rect 3200 27412 3206 27464
rect 5169 27455 5227 27461
rect 5169 27452 5181 27455
rect 4816 27424 5181 27452
rect 4614 27276 4620 27328
rect 4672 27316 4678 27328
rect 4816 27325 4844 27424
rect 5169 27421 5181 27424
rect 5215 27421 5227 27455
rect 5169 27415 5227 27421
rect 6362 27412 6368 27464
rect 6420 27452 6426 27464
rect 7760 27452 7788 27483
rect 8110 27480 8116 27492
rect 8168 27480 8174 27532
rect 8386 27480 8392 27532
rect 8444 27520 8450 27532
rect 8481 27523 8539 27529
rect 8481 27520 8493 27523
rect 8444 27492 8493 27520
rect 8444 27480 8450 27492
rect 8481 27489 8493 27492
rect 8527 27489 8539 27523
rect 8481 27483 8539 27489
rect 9677 27523 9735 27529
rect 9677 27489 9689 27523
rect 9723 27520 9735 27523
rect 10318 27520 10324 27532
rect 9723 27492 10324 27520
rect 9723 27489 9735 27492
rect 9677 27483 9735 27489
rect 10318 27480 10324 27492
rect 10376 27480 10382 27532
rect 11624 27529 11652 27560
rect 12618 27548 12624 27560
rect 12676 27548 12682 27600
rect 20070 27588 20076 27600
rect 20031 27560 20076 27588
rect 20070 27548 20076 27560
rect 20128 27548 20134 27600
rect 20714 27548 20720 27600
rect 20772 27588 20778 27600
rect 21269 27591 21327 27597
rect 21269 27588 21281 27591
rect 20772 27560 21281 27588
rect 20772 27548 20778 27560
rect 21269 27557 21281 27560
rect 21315 27557 21327 27591
rect 33410 27588 33416 27600
rect 21269 27551 21327 27557
rect 27264 27560 28304 27588
rect 10413 27523 10471 27529
rect 10413 27489 10425 27523
rect 10459 27489 10471 27523
rect 10413 27483 10471 27489
rect 11609 27523 11667 27529
rect 11609 27489 11621 27523
rect 11655 27489 11667 27523
rect 11790 27520 11796 27532
rect 11751 27492 11796 27520
rect 11609 27483 11667 27489
rect 6420 27424 7788 27452
rect 6420 27412 6426 27424
rect 7282 27384 7288 27396
rect 7243 27356 7288 27384
rect 7282 27344 7288 27356
rect 7340 27344 7346 27396
rect 7760 27384 7788 27424
rect 7926 27412 7932 27464
rect 7984 27452 7990 27464
rect 10428 27452 10456 27483
rect 11790 27480 11796 27492
rect 11848 27480 11854 27532
rect 12345 27523 12403 27529
rect 12345 27489 12357 27523
rect 12391 27520 12403 27523
rect 12434 27520 12440 27532
rect 12391 27492 12440 27520
rect 12391 27489 12403 27492
rect 12345 27483 12403 27489
rect 12434 27480 12440 27492
rect 12492 27480 12498 27532
rect 12713 27523 12771 27529
rect 12713 27489 12725 27523
rect 12759 27520 12771 27523
rect 13078 27520 13084 27532
rect 12759 27492 13084 27520
rect 12759 27489 12771 27492
rect 12713 27483 12771 27489
rect 7984 27424 10456 27452
rect 7984 27412 7990 27424
rect 10597 27387 10655 27393
rect 10597 27384 10609 27387
rect 7760 27356 10609 27384
rect 10597 27353 10609 27356
rect 10643 27353 10655 27387
rect 10597 27347 10655 27353
rect 11698 27344 11704 27396
rect 11756 27384 11762 27396
rect 12728 27384 12756 27483
rect 13078 27480 13084 27492
rect 13136 27480 13142 27532
rect 13814 27520 13820 27532
rect 13775 27492 13820 27520
rect 13814 27480 13820 27492
rect 13872 27480 13878 27532
rect 13998 27520 14004 27532
rect 13959 27492 14004 27520
rect 13998 27480 14004 27492
rect 14056 27480 14062 27532
rect 14458 27520 14464 27532
rect 14419 27492 14464 27520
rect 14458 27480 14464 27492
rect 14516 27480 14522 27532
rect 14550 27480 14556 27532
rect 14608 27520 14614 27532
rect 15657 27523 15715 27529
rect 15657 27520 15669 27523
rect 14608 27492 15669 27520
rect 14608 27480 14614 27492
rect 15657 27489 15669 27492
rect 15703 27489 15715 27523
rect 15657 27483 15715 27489
rect 15838 27480 15844 27532
rect 15896 27520 15902 27532
rect 16117 27523 16175 27529
rect 16117 27520 16129 27523
rect 15896 27492 16129 27520
rect 15896 27480 15902 27492
rect 16117 27489 16129 27492
rect 16163 27489 16175 27523
rect 16850 27520 16856 27532
rect 16811 27492 16856 27520
rect 16117 27483 16175 27489
rect 16850 27480 16856 27492
rect 16908 27480 16914 27532
rect 17865 27523 17923 27529
rect 17865 27489 17877 27523
rect 17911 27520 17923 27523
rect 18230 27520 18236 27532
rect 17911 27492 18236 27520
rect 17911 27489 17923 27492
rect 17865 27483 17923 27489
rect 18230 27480 18236 27492
rect 18288 27520 18294 27532
rect 19334 27520 19340 27532
rect 18288 27492 19340 27520
rect 18288 27480 18294 27492
rect 19334 27480 19340 27492
rect 19392 27480 19398 27532
rect 19518 27520 19524 27532
rect 19479 27492 19524 27520
rect 19518 27480 19524 27492
rect 19576 27480 19582 27532
rect 19978 27520 19984 27532
rect 19939 27492 19984 27520
rect 19978 27480 19984 27492
rect 20036 27480 20042 27532
rect 20438 27480 20444 27532
rect 20496 27520 20502 27532
rect 21361 27523 21419 27529
rect 21361 27520 21373 27523
rect 20496 27492 21373 27520
rect 20496 27480 20502 27492
rect 21361 27489 21373 27492
rect 21407 27489 21419 27523
rect 22002 27520 22008 27532
rect 21963 27492 22008 27520
rect 21361 27483 21419 27489
rect 22002 27480 22008 27492
rect 22060 27480 22066 27532
rect 22370 27520 22376 27532
rect 22331 27492 22376 27520
rect 22370 27480 22376 27492
rect 22428 27480 22434 27532
rect 22830 27520 22836 27532
rect 22791 27492 22836 27520
rect 22830 27480 22836 27492
rect 22888 27480 22894 27532
rect 23382 27520 23388 27532
rect 23343 27492 23388 27520
rect 23382 27480 23388 27492
rect 23440 27480 23446 27532
rect 23842 27520 23848 27532
rect 23803 27492 23848 27520
rect 23842 27480 23848 27492
rect 23900 27480 23906 27532
rect 24118 27520 24124 27532
rect 24079 27492 24124 27520
rect 24118 27480 24124 27492
rect 24176 27480 24182 27532
rect 24210 27480 24216 27532
rect 24268 27520 24274 27532
rect 24581 27523 24639 27529
rect 24581 27520 24593 27523
rect 24268 27492 24593 27520
rect 24268 27480 24274 27492
rect 24581 27489 24593 27492
rect 24627 27489 24639 27523
rect 24581 27483 24639 27489
rect 24949 27523 25007 27529
rect 24949 27489 24961 27523
rect 24995 27489 25007 27523
rect 24949 27483 25007 27489
rect 25685 27523 25743 27529
rect 25685 27489 25697 27523
rect 25731 27520 25743 27523
rect 26234 27520 26240 27532
rect 25731 27492 26240 27520
rect 25731 27489 25743 27492
rect 25685 27483 25743 27489
rect 14734 27452 14740 27464
rect 14695 27424 14740 27452
rect 14734 27412 14740 27424
rect 14792 27412 14798 27464
rect 15473 27455 15531 27461
rect 15473 27421 15485 27455
rect 15519 27452 15531 27455
rect 18141 27455 18199 27461
rect 15519 27424 15608 27452
rect 15519 27421 15531 27424
rect 15473 27415 15531 27421
rect 11756 27356 12756 27384
rect 11756 27344 11762 27356
rect 4801 27319 4859 27325
rect 4801 27316 4813 27319
rect 4672 27288 4813 27316
rect 4672 27276 4678 27288
rect 4801 27285 4813 27288
rect 4847 27285 4859 27319
rect 4801 27279 4859 27285
rect 8846 27276 8852 27328
rect 8904 27316 8910 27328
rect 9766 27316 9772 27328
rect 8904 27288 9772 27316
rect 8904 27276 8910 27288
rect 9766 27276 9772 27288
rect 9824 27316 9830 27328
rect 9861 27319 9919 27325
rect 9861 27316 9873 27319
rect 9824 27288 9873 27316
rect 9824 27276 9830 27288
rect 9861 27285 9873 27288
rect 9907 27285 9919 27319
rect 15580 27316 15608 27424
rect 18141 27421 18153 27455
rect 18187 27452 18199 27455
rect 22922 27452 22928 27464
rect 18187 27424 22928 27452
rect 18187 27421 18199 27424
rect 18141 27415 18199 27421
rect 22922 27412 22928 27424
rect 22980 27412 22986 27464
rect 23474 27452 23480 27464
rect 23435 27424 23480 27452
rect 23474 27412 23480 27424
rect 23532 27412 23538 27464
rect 16209 27387 16267 27393
rect 16209 27353 16221 27387
rect 16255 27384 16267 27387
rect 16255 27356 17908 27384
rect 16255 27353 16267 27356
rect 16209 27347 16267 27353
rect 15930 27316 15936 27328
rect 15580 27288 15936 27316
rect 9861 27279 9919 27285
rect 15930 27276 15936 27288
rect 15988 27316 15994 27328
rect 17037 27319 17095 27325
rect 17037 27316 17049 27319
rect 15988 27288 17049 27316
rect 15988 27276 15994 27288
rect 17037 27285 17049 27288
rect 17083 27285 17095 27319
rect 17880 27316 17908 27356
rect 19426 27344 19432 27396
rect 19484 27384 19490 27396
rect 20806 27384 20812 27396
rect 19484 27356 20812 27384
rect 19484 27344 19490 27356
rect 20806 27344 20812 27356
rect 20864 27344 20870 27396
rect 20901 27387 20959 27393
rect 20901 27353 20913 27387
rect 20947 27384 20959 27387
rect 21082 27384 21088 27396
rect 20947 27356 21088 27384
rect 20947 27353 20959 27356
rect 20901 27347 20959 27353
rect 21082 27344 21088 27356
rect 21140 27384 21146 27396
rect 24964 27384 24992 27483
rect 26234 27480 26240 27492
rect 26292 27520 26298 27532
rect 26786 27520 26792 27532
rect 26292 27492 26792 27520
rect 26292 27480 26298 27492
rect 26786 27480 26792 27492
rect 26844 27480 26850 27532
rect 27264 27529 27292 27560
rect 28276 27532 28304 27560
rect 32968 27560 33416 27588
rect 27249 27523 27307 27529
rect 27249 27489 27261 27523
rect 27295 27489 27307 27523
rect 27249 27483 27307 27489
rect 27617 27523 27675 27529
rect 27617 27489 27629 27523
rect 27663 27489 27675 27523
rect 27617 27483 27675 27489
rect 27154 27452 27160 27464
rect 25884 27424 27160 27452
rect 25884 27393 25912 27424
rect 27154 27412 27160 27424
rect 27212 27452 27218 27464
rect 27522 27452 27528 27464
rect 27212 27424 27528 27452
rect 27212 27412 27218 27424
rect 27522 27412 27528 27424
rect 27580 27452 27586 27464
rect 27632 27452 27660 27483
rect 28258 27480 28264 27532
rect 28316 27520 28322 27532
rect 30285 27523 30343 27529
rect 30285 27520 30297 27523
rect 28316 27492 30297 27520
rect 28316 27480 28322 27492
rect 30285 27489 30297 27492
rect 30331 27489 30343 27523
rect 30285 27483 30343 27489
rect 30374 27480 30380 27532
rect 30432 27520 30438 27532
rect 30653 27523 30711 27529
rect 30653 27520 30665 27523
rect 30432 27492 30665 27520
rect 30432 27480 30438 27492
rect 30653 27489 30665 27492
rect 30699 27489 30711 27523
rect 31202 27520 31208 27532
rect 31163 27492 31208 27520
rect 30653 27483 30711 27489
rect 31202 27480 31208 27492
rect 31260 27480 31266 27532
rect 32968 27529 32996 27560
rect 33410 27548 33416 27560
rect 33468 27548 33474 27600
rect 37093 27591 37151 27597
rect 37093 27588 37105 27591
rect 35360 27560 37105 27588
rect 32953 27523 33011 27529
rect 32953 27489 32965 27523
rect 32999 27489 33011 27523
rect 32953 27483 33011 27489
rect 33321 27523 33379 27529
rect 33321 27489 33333 27523
rect 33367 27520 33379 27523
rect 34698 27520 34704 27532
rect 33367 27492 34560 27520
rect 34659 27492 34704 27520
rect 33367 27489 33379 27492
rect 33321 27483 33379 27489
rect 27580 27424 27660 27452
rect 28169 27455 28227 27461
rect 27580 27412 27586 27424
rect 28169 27421 28181 27455
rect 28215 27421 28227 27455
rect 28442 27452 28448 27464
rect 28403 27424 28448 27452
rect 28169 27415 28227 27421
rect 21140 27356 24992 27384
rect 25869 27387 25927 27393
rect 21140 27344 21146 27356
rect 25869 27353 25881 27387
rect 25915 27353 25927 27387
rect 25869 27347 25927 27353
rect 26510 27344 26516 27396
rect 26568 27384 26574 27396
rect 27065 27387 27123 27393
rect 27065 27384 27077 27387
rect 26568 27356 27077 27384
rect 26568 27344 26574 27356
rect 27065 27353 27077 27356
rect 27111 27353 27123 27387
rect 27065 27347 27123 27353
rect 27430 27344 27436 27396
rect 27488 27384 27494 27396
rect 28184 27384 28212 27415
rect 28442 27412 28448 27424
rect 28500 27412 28506 27464
rect 32490 27452 32496 27464
rect 32451 27424 32496 27452
rect 32490 27412 32496 27424
rect 32548 27412 32554 27464
rect 34330 27412 34336 27464
rect 34388 27452 34394 27464
rect 34425 27455 34483 27461
rect 34425 27452 34437 27455
rect 34388 27424 34437 27452
rect 34388 27412 34394 27424
rect 34425 27421 34437 27424
rect 34471 27421 34483 27455
rect 34532 27452 34560 27492
rect 34698 27480 34704 27492
rect 34756 27480 34762 27532
rect 35360 27452 35388 27560
rect 37093 27557 37105 27560
rect 37139 27557 37151 27591
rect 37093 27551 37151 27557
rect 36538 27520 36544 27532
rect 36499 27492 36544 27520
rect 36538 27480 36544 27492
rect 36596 27480 36602 27532
rect 36725 27523 36783 27529
rect 36725 27489 36737 27523
rect 36771 27489 36783 27523
rect 37734 27520 37740 27532
rect 37695 27492 37740 27520
rect 36725 27483 36783 27489
rect 34532 27424 35388 27452
rect 34425 27415 34483 27421
rect 27488 27356 28212 27384
rect 27488 27344 27494 27356
rect 30650 27344 30656 27396
rect 30708 27384 30714 27396
rect 31113 27387 31171 27393
rect 31113 27384 31125 27387
rect 30708 27356 31125 27384
rect 30708 27344 30714 27356
rect 31113 27353 31125 27356
rect 31159 27353 31171 27387
rect 31113 27347 31171 27353
rect 32950 27344 32956 27396
rect 33008 27384 33014 27396
rect 33229 27387 33287 27393
rect 33229 27384 33241 27387
rect 33008 27356 33241 27384
rect 33008 27344 33014 27356
rect 33229 27353 33241 27356
rect 33275 27353 33287 27387
rect 36740 27384 36768 27483
rect 37734 27480 37740 27492
rect 37792 27480 37798 27532
rect 33229 27347 33287 27353
rect 35452 27356 36768 27384
rect 19150 27316 19156 27328
rect 17880 27288 19156 27316
rect 17037 27279 17095 27285
rect 19150 27276 19156 27288
rect 19208 27276 19214 27328
rect 19334 27276 19340 27328
rect 19392 27316 19398 27328
rect 20622 27316 20628 27328
rect 19392 27288 20628 27316
rect 19392 27276 19398 27288
rect 20622 27276 20628 27288
rect 20680 27276 20686 27328
rect 22278 27276 22284 27328
rect 22336 27316 22342 27328
rect 23382 27316 23388 27328
rect 22336 27288 23388 27316
rect 22336 27276 22342 27288
rect 23382 27276 23388 27288
rect 23440 27276 23446 27328
rect 29733 27319 29791 27325
rect 29733 27285 29745 27319
rect 29779 27316 29791 27319
rect 29914 27316 29920 27328
rect 29779 27288 29920 27316
rect 29779 27285 29791 27288
rect 29733 27279 29791 27285
rect 29914 27276 29920 27288
rect 29972 27276 29978 27328
rect 33778 27276 33784 27328
rect 33836 27316 33842 27328
rect 35452 27316 35480 27356
rect 33836 27288 35480 27316
rect 33836 27276 33842 27288
rect 35526 27276 35532 27328
rect 35584 27316 35590 27328
rect 35989 27319 36047 27325
rect 35989 27316 36001 27319
rect 35584 27288 36001 27316
rect 35584 27276 35590 27288
rect 35989 27285 36001 27288
rect 36035 27285 36047 27319
rect 37826 27316 37832 27328
rect 37787 27288 37832 27316
rect 35989 27279 36047 27285
rect 37826 27276 37832 27288
rect 37884 27276 37890 27328
rect 1104 27226 38824 27248
rect 1104 27174 4246 27226
rect 4298 27174 4310 27226
rect 4362 27174 4374 27226
rect 4426 27174 4438 27226
rect 4490 27174 34966 27226
rect 35018 27174 35030 27226
rect 35082 27174 35094 27226
rect 35146 27174 35158 27226
rect 35210 27174 38824 27226
rect 1104 27152 38824 27174
rect 1486 27112 1492 27124
rect 1447 27084 1492 27112
rect 1486 27072 1492 27084
rect 1544 27072 1550 27124
rect 1670 27072 1676 27124
rect 1728 27112 1734 27124
rect 1949 27115 2007 27121
rect 1949 27112 1961 27115
rect 1728 27084 1961 27112
rect 1728 27072 1734 27084
rect 1949 27081 1961 27084
rect 1995 27081 2007 27115
rect 4062 27112 4068 27124
rect 4023 27084 4068 27112
rect 1949 27075 2007 27081
rect 4062 27072 4068 27084
rect 4120 27072 4126 27124
rect 4798 27072 4804 27124
rect 4856 27112 4862 27124
rect 5077 27115 5135 27121
rect 5077 27112 5089 27115
rect 4856 27084 5089 27112
rect 4856 27072 4862 27084
rect 5077 27081 5089 27084
rect 5123 27081 5135 27115
rect 5077 27075 5135 27081
rect 6181 27115 6239 27121
rect 6181 27081 6193 27115
rect 6227 27112 6239 27115
rect 8110 27112 8116 27124
rect 6227 27084 8116 27112
rect 6227 27081 6239 27084
rect 6181 27075 6239 27081
rect 8110 27072 8116 27084
rect 8168 27072 8174 27124
rect 14734 27072 14740 27124
rect 14792 27112 14798 27124
rect 22922 27112 22928 27124
rect 14792 27084 22324 27112
rect 22883 27084 22928 27112
rect 14792 27072 14798 27084
rect 11790 27044 11796 27056
rect 11440 27016 11796 27044
rect 2608 26948 5028 26976
rect 1762 26908 1768 26920
rect 1723 26880 1768 26908
rect 1762 26868 1768 26880
rect 1820 26868 1826 26920
rect 1673 26843 1731 26849
rect 1673 26809 1685 26843
rect 1719 26840 1731 26843
rect 2608 26840 2636 26948
rect 2685 26911 2743 26917
rect 2685 26877 2697 26911
rect 2731 26877 2743 26911
rect 2685 26871 2743 26877
rect 1719 26812 2636 26840
rect 2700 26840 2728 26871
rect 2774 26868 2780 26920
rect 2832 26908 2838 26920
rect 3053 26911 3111 26917
rect 3053 26908 3065 26911
rect 2832 26880 3065 26908
rect 2832 26868 2838 26880
rect 3053 26877 3065 26880
rect 3099 26877 3111 26911
rect 3053 26871 3111 26877
rect 3142 26868 3148 26920
rect 3200 26908 3206 26920
rect 3421 26911 3479 26917
rect 3421 26908 3433 26911
rect 3200 26880 3433 26908
rect 3200 26868 3206 26880
rect 3421 26877 3433 26880
rect 3467 26877 3479 26911
rect 4062 26908 4068 26920
rect 4023 26880 4068 26908
rect 3421 26871 3479 26877
rect 4062 26868 4068 26880
rect 4120 26868 4126 26920
rect 4614 26908 4620 26920
rect 4575 26880 4620 26908
rect 4614 26868 4620 26880
rect 4672 26868 4678 26920
rect 4890 26908 4896 26920
rect 4851 26880 4896 26908
rect 4890 26868 4896 26880
rect 4948 26868 4954 26920
rect 4706 26840 4712 26852
rect 2700 26812 4712 26840
rect 1719 26809 1731 26812
rect 1673 26803 1731 26809
rect 4706 26800 4712 26812
rect 4764 26800 4770 26852
rect 4801 26843 4859 26849
rect 4801 26809 4813 26843
rect 4847 26840 4859 26843
rect 5000 26840 5028 26948
rect 7374 26936 7380 26988
rect 7432 26976 7438 26988
rect 8018 26976 8024 26988
rect 7432 26948 8024 26976
rect 7432 26936 7438 26948
rect 8018 26936 8024 26948
rect 8076 26936 8082 26988
rect 8662 26936 8668 26988
rect 8720 26976 8726 26988
rect 8941 26979 8999 26985
rect 8941 26976 8953 26979
rect 8720 26948 8953 26976
rect 8720 26936 8726 26948
rect 8941 26945 8953 26948
rect 8987 26945 8999 26979
rect 9214 26976 9220 26988
rect 9175 26948 9220 26976
rect 8941 26939 8999 26945
rect 6089 26911 6147 26917
rect 6089 26877 6101 26911
rect 6135 26908 6147 26911
rect 6914 26908 6920 26920
rect 6135 26880 6920 26908
rect 6135 26877 6147 26880
rect 6089 26871 6147 26877
rect 6914 26868 6920 26880
rect 6972 26868 6978 26920
rect 7190 26908 7196 26920
rect 7151 26880 7196 26908
rect 7190 26868 7196 26880
rect 7248 26868 7254 26920
rect 7926 26908 7932 26920
rect 7887 26880 7932 26908
rect 7926 26868 7932 26880
rect 7984 26868 7990 26920
rect 8956 26908 8984 26939
rect 9214 26936 9220 26948
rect 9272 26936 9278 26988
rect 9306 26936 9312 26988
rect 9364 26976 9370 26988
rect 9364 26948 11376 26976
rect 9364 26936 9370 26948
rect 9674 26908 9680 26920
rect 8956 26880 9680 26908
rect 9674 26868 9680 26880
rect 9732 26868 9738 26920
rect 10597 26911 10655 26917
rect 10597 26877 10609 26911
rect 10643 26908 10655 26911
rect 11238 26908 11244 26920
rect 10643 26880 11244 26908
rect 10643 26877 10655 26880
rect 10597 26871 10655 26877
rect 11238 26868 11244 26880
rect 11296 26868 11302 26920
rect 5994 26840 6000 26852
rect 4847 26812 6000 26840
rect 4847 26809 4859 26812
rect 4801 26803 4859 26809
rect 5994 26800 6000 26812
rect 6052 26800 6058 26852
rect 6932 26840 6960 26868
rect 6932 26812 9076 26840
rect 7374 26772 7380 26784
rect 7335 26744 7380 26772
rect 7374 26732 7380 26744
rect 7432 26732 7438 26784
rect 7466 26732 7472 26784
rect 7524 26772 7530 26784
rect 8113 26775 8171 26781
rect 8113 26772 8125 26775
rect 7524 26744 8125 26772
rect 7524 26732 7530 26744
rect 8113 26741 8125 26744
rect 8159 26741 8171 26775
rect 9048 26772 9076 26812
rect 10318 26800 10324 26852
rect 10376 26840 10382 26852
rect 10376 26812 11284 26840
rect 10376 26800 10382 26812
rect 11146 26772 11152 26784
rect 9048 26744 11152 26772
rect 8113 26735 8171 26741
rect 11146 26732 11152 26744
rect 11204 26732 11210 26784
rect 11256 26781 11284 26812
rect 11241 26775 11299 26781
rect 11241 26741 11253 26775
rect 11287 26741 11299 26775
rect 11348 26772 11376 26948
rect 11440 26917 11468 27016
rect 11790 27004 11796 27016
rect 11848 27044 11854 27056
rect 12710 27044 12716 27056
rect 11848 27016 12716 27044
rect 11848 27004 11854 27016
rect 11425 26911 11483 26917
rect 11425 26877 11437 26911
rect 11471 26877 11483 26911
rect 11698 26908 11704 26920
rect 11659 26880 11704 26908
rect 11425 26871 11483 26877
rect 11698 26868 11704 26880
rect 11756 26868 11762 26920
rect 12452 26917 12480 27016
rect 12710 27004 12716 27016
rect 12768 27004 12774 27056
rect 13814 27004 13820 27056
rect 13872 27044 13878 27056
rect 17218 27044 17224 27056
rect 13872 27016 17224 27044
rect 13872 27004 13878 27016
rect 17218 27004 17224 27016
rect 17276 27004 17282 27056
rect 17405 27047 17463 27053
rect 17405 27013 17417 27047
rect 17451 27044 17463 27047
rect 17678 27044 17684 27056
rect 17451 27016 17684 27044
rect 17451 27013 17463 27016
rect 17405 27007 17463 27013
rect 17678 27004 17684 27016
rect 17736 27004 17742 27056
rect 20714 27044 20720 27056
rect 17788 27016 20720 27044
rect 15838 26976 15844 26988
rect 14752 26948 15844 26976
rect 12437 26911 12495 26917
rect 12437 26877 12449 26911
rect 12483 26877 12495 26911
rect 12437 26871 12495 26877
rect 12526 26868 12532 26920
rect 12584 26908 12590 26920
rect 12897 26911 12955 26917
rect 12897 26908 12909 26911
rect 12584 26880 12909 26908
rect 12584 26868 12590 26880
rect 12897 26877 12909 26880
rect 12943 26908 12955 26911
rect 12986 26908 12992 26920
rect 12943 26880 12992 26908
rect 12943 26877 12955 26880
rect 12897 26871 12955 26877
rect 12986 26868 12992 26880
rect 13044 26868 13050 26920
rect 13078 26868 13084 26920
rect 13136 26908 13142 26920
rect 14752 26917 14780 26948
rect 15838 26936 15844 26948
rect 15896 26936 15902 26988
rect 17586 26936 17592 26988
rect 17644 26976 17650 26988
rect 17788 26976 17816 27016
rect 20714 27004 20720 27016
rect 20772 27004 20778 27056
rect 22296 27044 22324 27084
rect 22922 27072 22928 27084
rect 22980 27072 22986 27124
rect 24489 27115 24547 27121
rect 23032 27084 24256 27112
rect 23032 27044 23060 27084
rect 22296 27016 23060 27044
rect 23382 27004 23388 27056
rect 23440 27044 23446 27056
rect 23983 27047 24041 27053
rect 23983 27044 23995 27047
rect 23440 27016 23995 27044
rect 23440 27004 23446 27016
rect 23983 27013 23995 27016
rect 24029 27044 24041 27047
rect 24118 27044 24124 27056
rect 24029 27016 24124 27044
rect 24029 27013 24041 27016
rect 23983 27007 24041 27013
rect 24118 27004 24124 27016
rect 24176 27004 24182 27056
rect 24228 27044 24256 27084
rect 24489 27081 24501 27115
rect 24535 27112 24547 27115
rect 24946 27112 24952 27124
rect 24535 27084 24952 27112
rect 24535 27081 24547 27084
rect 24489 27075 24547 27081
rect 24946 27072 24952 27084
rect 25004 27072 25010 27124
rect 31849 27115 31907 27121
rect 31849 27081 31861 27115
rect 31895 27112 31907 27115
rect 32030 27112 32036 27124
rect 31895 27084 32036 27112
rect 31895 27081 31907 27084
rect 31849 27075 31907 27081
rect 32030 27072 32036 27084
rect 32088 27072 32094 27124
rect 33778 27112 33784 27124
rect 33739 27084 33784 27112
rect 33778 27072 33784 27084
rect 33836 27072 33842 27124
rect 25314 27044 25320 27056
rect 24228 27016 25320 27044
rect 25314 27004 25320 27016
rect 25372 27004 25378 27056
rect 28442 27044 28448 27056
rect 28403 27016 28448 27044
rect 28442 27004 28448 27016
rect 28500 27004 28506 27056
rect 30282 27004 30288 27056
rect 30340 27044 30346 27056
rect 34517 27047 34575 27053
rect 30340 27016 32444 27044
rect 30340 27004 30346 27016
rect 19334 26976 19340 26988
rect 17644 26948 17816 26976
rect 18064 26948 19340 26976
rect 17644 26936 17650 26948
rect 13265 26911 13323 26917
rect 13265 26908 13277 26911
rect 13136 26880 13277 26908
rect 13136 26868 13142 26880
rect 13265 26877 13277 26880
rect 13311 26877 13323 26911
rect 13265 26871 13323 26877
rect 14185 26911 14243 26917
rect 14185 26877 14197 26911
rect 14231 26877 14243 26911
rect 14185 26871 14243 26877
rect 14737 26911 14795 26917
rect 14737 26877 14749 26911
rect 14783 26877 14795 26911
rect 14737 26871 14795 26877
rect 15013 26911 15071 26917
rect 15013 26877 15025 26911
rect 15059 26908 15071 26911
rect 15102 26908 15108 26920
rect 15059 26880 15108 26908
rect 15059 26877 15071 26880
rect 15013 26871 15071 26877
rect 14200 26840 14228 26871
rect 15102 26868 15108 26880
rect 15160 26868 15166 26920
rect 15933 26911 15991 26917
rect 15933 26877 15945 26911
rect 15979 26877 15991 26911
rect 16390 26908 16396 26920
rect 16351 26880 16396 26908
rect 15933 26871 15991 26877
rect 15562 26840 15568 26852
rect 14200 26812 15568 26840
rect 15562 26800 15568 26812
rect 15620 26800 15626 26852
rect 15948 26840 15976 26871
rect 16390 26868 16396 26880
rect 16448 26868 16454 26920
rect 16574 26908 16580 26920
rect 16535 26880 16580 26908
rect 16574 26868 16580 26880
rect 16632 26868 16638 26920
rect 18064 26917 18092 26948
rect 17313 26911 17371 26917
rect 17313 26877 17325 26911
rect 17359 26908 17371 26911
rect 18049 26911 18107 26917
rect 17359 26880 18000 26908
rect 17359 26877 17371 26880
rect 17313 26871 17371 26877
rect 16942 26840 16948 26852
rect 15948 26812 16948 26840
rect 16942 26800 16948 26812
rect 17000 26800 17006 26852
rect 12529 26775 12587 26781
rect 12529 26772 12541 26775
rect 11348 26744 12541 26772
rect 11241 26735 11299 26741
rect 12529 26741 12541 26744
rect 12575 26741 12587 26775
rect 12529 26735 12587 26741
rect 14093 26775 14151 26781
rect 14093 26741 14105 26775
rect 14139 26772 14151 26775
rect 14366 26772 14372 26784
rect 14139 26744 14372 26772
rect 14139 26741 14151 26744
rect 14093 26735 14151 26741
rect 14366 26732 14372 26744
rect 14424 26732 14430 26784
rect 15841 26775 15899 26781
rect 15841 26741 15853 26775
rect 15887 26772 15899 26775
rect 17770 26772 17776 26784
rect 15887 26744 17776 26772
rect 15887 26741 15899 26744
rect 15841 26735 15899 26741
rect 17770 26732 17776 26744
rect 17828 26732 17834 26784
rect 17972 26772 18000 26880
rect 18049 26877 18061 26911
rect 18095 26877 18107 26911
rect 18049 26871 18107 26877
rect 18233 26911 18291 26917
rect 18233 26877 18245 26911
rect 18279 26908 18291 26911
rect 18966 26908 18972 26920
rect 18279 26880 18972 26908
rect 18279 26877 18291 26880
rect 18233 26871 18291 26877
rect 18966 26868 18972 26880
rect 19024 26868 19030 26920
rect 19260 26917 19288 26948
rect 19334 26936 19340 26948
rect 19392 26936 19398 26988
rect 20257 26979 20315 26985
rect 20257 26945 20269 26979
rect 20303 26976 20315 26979
rect 21174 26976 21180 26988
rect 20303 26948 21180 26976
rect 20303 26945 20315 26948
rect 20257 26939 20315 26945
rect 21174 26936 21180 26948
rect 21232 26936 21238 26988
rect 22094 26936 22100 26988
rect 22152 26976 22158 26988
rect 32416 26985 32444 27016
rect 34517 27013 34529 27047
rect 34563 27013 34575 27047
rect 34517 27007 34575 27013
rect 24213 26979 24271 26985
rect 24213 26976 24225 26979
rect 22152 26948 24225 26976
rect 22152 26936 22158 26948
rect 24213 26945 24225 26948
rect 24259 26945 24271 26979
rect 24213 26939 24271 26945
rect 25501 26979 25559 26985
rect 25501 26945 25513 26979
rect 25547 26976 25559 26979
rect 32401 26979 32459 26985
rect 25547 26948 27936 26976
rect 25547 26945 25559 26948
rect 25501 26939 25559 26945
rect 19245 26911 19303 26917
rect 19245 26877 19257 26911
rect 19291 26877 19303 26911
rect 19245 26871 19303 26877
rect 19518 26868 19524 26920
rect 19576 26908 19582 26920
rect 19705 26911 19763 26917
rect 19705 26908 19717 26911
rect 19576 26880 19717 26908
rect 19576 26868 19582 26880
rect 19705 26877 19717 26880
rect 19751 26877 19763 26911
rect 19705 26871 19763 26877
rect 19720 26840 19748 26871
rect 19886 26868 19892 26920
rect 19944 26908 19950 26920
rect 20073 26911 20131 26917
rect 20073 26908 20085 26911
rect 19944 26880 20085 26908
rect 19944 26868 19950 26880
rect 20073 26877 20085 26880
rect 20119 26908 20131 26911
rect 20438 26908 20444 26920
rect 20119 26880 20444 26908
rect 20119 26877 20131 26880
rect 20073 26871 20131 26877
rect 20438 26868 20444 26880
rect 20496 26868 20502 26920
rect 20622 26868 20628 26920
rect 20680 26908 20686 26920
rect 20717 26911 20775 26917
rect 20717 26908 20729 26911
rect 20680 26880 20729 26908
rect 20680 26868 20686 26880
rect 20717 26877 20729 26880
rect 20763 26877 20775 26911
rect 20990 26908 20996 26920
rect 20951 26880 20996 26908
rect 20717 26871 20775 26877
rect 20990 26868 20996 26880
rect 21048 26868 21054 26920
rect 21082 26868 21088 26920
rect 21140 26908 21146 26920
rect 22833 26911 22891 26917
rect 22833 26908 22845 26911
rect 21140 26880 22845 26908
rect 21140 26868 21146 26880
rect 22833 26877 22845 26880
rect 22879 26877 22891 26911
rect 22833 26871 22891 26877
rect 23566 26868 23572 26920
rect 23624 26908 23630 26920
rect 24075 26911 24133 26917
rect 24075 26908 24087 26911
rect 23624 26880 24087 26908
rect 23624 26868 23630 26880
rect 24075 26877 24087 26880
rect 24121 26877 24133 26911
rect 24075 26871 24133 26877
rect 24762 26868 24768 26920
rect 24820 26908 24826 26920
rect 25041 26911 25099 26917
rect 25041 26908 25053 26911
rect 24820 26880 25053 26908
rect 24820 26868 24826 26880
rect 25041 26877 25053 26880
rect 25087 26877 25099 26911
rect 25590 26908 25596 26920
rect 25551 26880 25596 26908
rect 25041 26871 25099 26877
rect 25590 26868 25596 26880
rect 25648 26868 25654 26920
rect 25866 26908 25872 26920
rect 25827 26880 25872 26908
rect 25866 26868 25872 26880
rect 25924 26868 25930 26920
rect 26050 26868 26056 26920
rect 26108 26908 26114 26920
rect 26237 26911 26295 26917
rect 26237 26908 26249 26911
rect 26108 26880 26249 26908
rect 26108 26868 26114 26880
rect 26237 26877 26249 26880
rect 26283 26877 26295 26911
rect 26237 26871 26295 26877
rect 27522 26868 27528 26920
rect 27580 26908 27586 26920
rect 27908 26917 27936 26948
rect 30392 26948 31708 26976
rect 30392 26920 30420 26948
rect 27617 26911 27675 26917
rect 27617 26908 27629 26911
rect 27580 26880 27629 26908
rect 27580 26868 27586 26880
rect 27617 26877 27629 26880
rect 27663 26877 27675 26911
rect 27617 26871 27675 26877
rect 27893 26911 27951 26917
rect 27893 26877 27905 26911
rect 27939 26877 27951 26911
rect 28442 26908 28448 26920
rect 28403 26880 28448 26908
rect 27893 26871 27951 26877
rect 28442 26868 28448 26880
rect 28500 26868 28506 26920
rect 29086 26868 29092 26920
rect 29144 26908 29150 26920
rect 29273 26911 29331 26917
rect 29273 26908 29285 26911
rect 29144 26880 29285 26908
rect 29144 26868 29150 26880
rect 29273 26877 29285 26880
rect 29319 26877 29331 26911
rect 29914 26908 29920 26920
rect 29875 26880 29920 26908
rect 29273 26871 29331 26877
rect 29914 26868 29920 26880
rect 29972 26868 29978 26920
rect 30374 26908 30380 26920
rect 30335 26880 30380 26908
rect 30374 26868 30380 26880
rect 30432 26868 30438 26920
rect 31680 26917 31708 26948
rect 32401 26945 32413 26979
rect 32447 26976 32459 26979
rect 32766 26976 32772 26988
rect 32447 26948 32772 26976
rect 32447 26945 32459 26948
rect 32401 26939 32459 26945
rect 32766 26936 32772 26948
rect 32824 26976 32830 26988
rect 34330 26976 34336 26988
rect 32824 26948 34336 26976
rect 32824 26936 32830 26948
rect 34330 26936 34336 26948
rect 34388 26976 34394 26988
rect 34532 26976 34560 27007
rect 34388 26948 34560 26976
rect 35069 26979 35127 26985
rect 34388 26936 34394 26948
rect 35069 26945 35081 26979
rect 35115 26976 35127 26979
rect 36725 26979 36783 26985
rect 35115 26948 36584 26976
rect 35115 26945 35127 26948
rect 35069 26939 35127 26945
rect 30837 26911 30895 26917
rect 30837 26877 30849 26911
rect 30883 26877 30895 26911
rect 30837 26871 30895 26877
rect 31665 26911 31723 26917
rect 31665 26877 31677 26911
rect 31711 26908 31723 26911
rect 32306 26908 32312 26920
rect 31711 26880 32312 26908
rect 31711 26877 31723 26880
rect 31665 26871 31723 26877
rect 19978 26840 19984 26852
rect 18156 26812 19984 26840
rect 18156 26772 18184 26812
rect 19978 26800 19984 26812
rect 20036 26800 20042 26852
rect 23658 26840 23664 26852
rect 21652 26812 23664 26840
rect 18322 26772 18328 26784
rect 17972 26744 18184 26772
rect 18283 26744 18328 26772
rect 18322 26732 18328 26744
rect 18380 26732 18386 26784
rect 19150 26732 19156 26784
rect 19208 26772 19214 26784
rect 21652 26772 21680 26812
rect 23658 26800 23664 26812
rect 23716 26800 23722 26852
rect 23842 26840 23848 26852
rect 23755 26812 23848 26840
rect 23842 26800 23848 26812
rect 23900 26840 23906 26852
rect 24486 26840 24492 26852
rect 23900 26812 24492 26840
rect 23900 26800 23906 26812
rect 24486 26800 24492 26812
rect 24544 26800 24550 26852
rect 19208 26744 21680 26772
rect 19208 26732 19214 26744
rect 22002 26732 22008 26784
rect 22060 26772 22066 26784
rect 22097 26775 22155 26781
rect 22097 26772 22109 26775
rect 22060 26744 22109 26772
rect 22060 26732 22066 26744
rect 22097 26741 22109 26744
rect 22143 26741 22155 26775
rect 22097 26735 22155 26741
rect 22738 26732 22744 26784
rect 22796 26772 22802 26784
rect 23860 26772 23888 26800
rect 22796 26744 23888 26772
rect 22796 26732 22802 26744
rect 27982 26732 27988 26784
rect 28040 26772 28046 26784
rect 29365 26775 29423 26781
rect 29365 26772 29377 26775
rect 28040 26744 29377 26772
rect 28040 26732 28046 26744
rect 29365 26741 29377 26744
rect 29411 26741 29423 26775
rect 30852 26772 30880 26871
rect 32306 26868 32312 26880
rect 32364 26868 32370 26920
rect 32674 26908 32680 26920
rect 32635 26880 32680 26908
rect 32674 26868 32680 26880
rect 32732 26868 32738 26920
rect 34606 26868 34612 26920
rect 34664 26908 34670 26920
rect 34701 26911 34759 26917
rect 34701 26908 34713 26911
rect 34664 26880 34713 26908
rect 34664 26868 34670 26880
rect 34701 26877 34713 26880
rect 34747 26877 34759 26911
rect 34701 26871 34759 26877
rect 35437 26911 35495 26917
rect 35437 26877 35449 26911
rect 35483 26877 35495 26911
rect 35710 26908 35716 26920
rect 35671 26880 35716 26908
rect 35437 26871 35495 26877
rect 31021 26843 31079 26849
rect 31021 26809 31033 26843
rect 31067 26840 31079 26843
rect 32214 26840 32220 26852
rect 31067 26812 32220 26840
rect 31067 26809 31079 26812
rect 31021 26803 31079 26809
rect 32214 26800 32220 26812
rect 32272 26800 32278 26852
rect 31110 26772 31116 26784
rect 30852 26744 31116 26772
rect 29365 26735 29423 26741
rect 31110 26732 31116 26744
rect 31168 26732 31174 26784
rect 35452 26772 35480 26871
rect 35710 26868 35716 26880
rect 35768 26868 35774 26920
rect 36354 26868 36360 26920
rect 36412 26908 36418 26920
rect 36449 26911 36507 26917
rect 36449 26908 36461 26911
rect 36412 26880 36461 26908
rect 36412 26868 36418 26880
rect 36449 26877 36461 26880
rect 36495 26877 36507 26911
rect 36556 26908 36584 26948
rect 36725 26945 36737 26979
rect 36771 26976 36783 26979
rect 37826 26976 37832 26988
rect 36771 26948 37832 26976
rect 36771 26945 36783 26948
rect 36725 26939 36783 26945
rect 37826 26936 37832 26948
rect 37884 26936 37890 26988
rect 36998 26908 37004 26920
rect 36556 26880 37004 26908
rect 36449 26871 36507 26877
rect 36998 26868 37004 26880
rect 37056 26868 37062 26920
rect 35986 26840 35992 26852
rect 35947 26812 35992 26840
rect 35986 26800 35992 26812
rect 36044 26800 36050 26852
rect 36814 26772 36820 26784
rect 35452 26744 36820 26772
rect 36814 26732 36820 26744
rect 36872 26732 36878 26784
rect 36998 26732 37004 26784
rect 37056 26772 37062 26784
rect 37829 26775 37887 26781
rect 37829 26772 37841 26775
rect 37056 26744 37841 26772
rect 37056 26732 37062 26744
rect 37829 26741 37841 26744
rect 37875 26741 37887 26775
rect 37829 26735 37887 26741
rect 1104 26682 38824 26704
rect 1104 26630 19606 26682
rect 19658 26630 19670 26682
rect 19722 26630 19734 26682
rect 19786 26630 19798 26682
rect 19850 26630 38824 26682
rect 1104 26608 38824 26630
rect 12434 26568 12440 26580
rect 10612 26540 12440 26568
rect 1394 26432 1400 26444
rect 1355 26404 1400 26432
rect 1394 26392 1400 26404
rect 1452 26392 1458 26444
rect 1670 26432 1676 26444
rect 1631 26404 1676 26432
rect 1670 26392 1676 26404
rect 1728 26392 1734 26444
rect 4798 26432 4804 26444
rect 4759 26404 4804 26432
rect 4798 26392 4804 26404
rect 4856 26392 4862 26444
rect 7190 26432 7196 26444
rect 7151 26404 7196 26432
rect 7190 26392 7196 26404
rect 7248 26392 7254 26444
rect 8570 26432 8576 26444
rect 8531 26404 8576 26432
rect 8570 26392 8576 26404
rect 8628 26392 8634 26444
rect 8754 26432 8760 26444
rect 8715 26404 8760 26432
rect 8754 26392 8760 26404
rect 8812 26392 8818 26444
rect 8846 26392 8852 26444
rect 8904 26432 8910 26444
rect 10612 26441 10640 26540
rect 12434 26528 12440 26540
rect 12492 26528 12498 26580
rect 12618 26528 12624 26580
rect 12676 26568 12682 26580
rect 15657 26571 15715 26577
rect 12676 26540 14872 26568
rect 12676 26528 12682 26540
rect 11146 26460 11152 26512
rect 11204 26500 11210 26512
rect 11204 26472 11836 26500
rect 11204 26460 11210 26472
rect 8941 26435 8999 26441
rect 8941 26432 8953 26435
rect 8904 26404 8953 26432
rect 8904 26392 8910 26404
rect 8941 26401 8953 26404
rect 8987 26401 8999 26435
rect 8941 26395 8999 26401
rect 10137 26435 10195 26441
rect 10137 26401 10149 26435
rect 10183 26432 10195 26435
rect 10597 26435 10655 26441
rect 10183 26404 10364 26432
rect 10183 26401 10195 26404
rect 10137 26395 10195 26401
rect 1412 26364 1440 26392
rect 4522 26364 4528 26376
rect 1412 26336 4528 26364
rect 2682 26256 2688 26308
rect 2740 26296 2746 26308
rect 2777 26299 2835 26305
rect 2777 26296 2789 26299
rect 2740 26268 2789 26296
rect 2740 26256 2746 26268
rect 2777 26265 2789 26268
rect 2823 26265 2835 26299
rect 2777 26259 2835 26265
rect 4448 26228 4476 26336
rect 4522 26324 4528 26336
rect 4580 26324 4586 26376
rect 4706 26324 4712 26376
rect 4764 26364 4770 26376
rect 5905 26367 5963 26373
rect 5905 26364 5917 26367
rect 4764 26336 5917 26364
rect 4764 26324 4770 26336
rect 5905 26333 5917 26336
rect 5951 26333 5963 26367
rect 5905 26327 5963 26333
rect 10229 26367 10287 26373
rect 10229 26333 10241 26367
rect 10275 26333 10287 26367
rect 10336 26364 10364 26404
rect 10597 26401 10609 26435
rect 10643 26401 10655 26435
rect 10597 26395 10655 26401
rect 10778 26392 10784 26444
rect 10836 26432 10842 26444
rect 11057 26435 11115 26441
rect 11057 26432 11069 26435
rect 10836 26404 11069 26432
rect 10836 26392 10842 26404
rect 11057 26401 11069 26404
rect 11103 26401 11115 26435
rect 11698 26432 11704 26444
rect 11659 26404 11704 26432
rect 11057 26395 11115 26401
rect 11698 26392 11704 26404
rect 11756 26392 11762 26444
rect 11808 26441 11836 26472
rect 11882 26460 11888 26512
rect 11940 26500 11946 26512
rect 14844 26500 14872 26540
rect 15657 26537 15669 26571
rect 15703 26568 15715 26571
rect 16574 26568 16580 26580
rect 15703 26540 16580 26568
rect 15703 26537 15715 26540
rect 15657 26531 15715 26537
rect 16574 26528 16580 26540
rect 16632 26528 16638 26580
rect 19978 26528 19984 26580
rect 20036 26568 20042 26580
rect 20254 26568 20260 26580
rect 20036 26540 20260 26568
rect 20036 26528 20042 26540
rect 20254 26528 20260 26540
rect 20312 26568 20318 26580
rect 22370 26568 22376 26580
rect 20312 26540 22376 26568
rect 20312 26528 20318 26540
rect 22370 26528 22376 26540
rect 22428 26568 22434 26580
rect 23106 26568 23112 26580
rect 22428 26540 23112 26568
rect 22428 26528 22434 26540
rect 23106 26528 23112 26540
rect 23164 26528 23170 26580
rect 25869 26571 25927 26577
rect 25869 26537 25881 26571
rect 25915 26568 25927 26571
rect 26050 26568 26056 26580
rect 25915 26540 26056 26568
rect 25915 26537 25927 26540
rect 25869 26531 25927 26537
rect 26050 26528 26056 26540
rect 26108 26528 26114 26580
rect 26973 26571 27031 26577
rect 26973 26537 26985 26571
rect 27019 26568 27031 26571
rect 29638 26568 29644 26580
rect 27019 26540 29644 26568
rect 27019 26537 27031 26540
rect 26973 26531 27031 26537
rect 29638 26528 29644 26540
rect 29696 26528 29702 26580
rect 32309 26571 32367 26577
rect 32309 26537 32321 26571
rect 32355 26568 32367 26571
rect 32674 26568 32680 26580
rect 32355 26540 32680 26568
rect 32355 26537 32367 26540
rect 32309 26531 32367 26537
rect 32674 26528 32680 26540
rect 32732 26528 32738 26580
rect 11940 26472 14780 26500
rect 14844 26472 16436 26500
rect 11940 26460 11946 26472
rect 11793 26435 11851 26441
rect 11793 26401 11805 26435
rect 11839 26401 11851 26435
rect 12526 26432 12532 26444
rect 12487 26404 12532 26432
rect 11793 26395 11851 26401
rect 12526 26392 12532 26404
rect 12584 26392 12590 26444
rect 12986 26432 12992 26444
rect 12947 26404 12992 26432
rect 12986 26392 12992 26404
rect 13044 26392 13050 26444
rect 13725 26435 13783 26441
rect 13725 26401 13737 26435
rect 13771 26432 13783 26435
rect 13814 26432 13820 26444
rect 13771 26404 13820 26432
rect 13771 26401 13783 26404
rect 13725 26395 13783 26401
rect 13814 26392 13820 26404
rect 13872 26392 13878 26444
rect 14752 26441 14780 26472
rect 14553 26435 14611 26441
rect 14553 26401 14565 26435
rect 14599 26401 14611 26435
rect 14553 26395 14611 26401
rect 14737 26435 14795 26441
rect 14737 26401 14749 26435
rect 14783 26401 14795 26435
rect 14737 26395 14795 26401
rect 15749 26435 15807 26441
rect 15749 26401 15761 26435
rect 15795 26432 15807 26435
rect 15838 26432 15844 26444
rect 15795 26404 15844 26432
rect 15795 26401 15807 26404
rect 15749 26395 15807 26401
rect 11149 26367 11207 26373
rect 11149 26364 11161 26367
rect 10336 26336 11161 26364
rect 10229 26327 10287 26333
rect 11149 26333 11161 26336
rect 11195 26333 11207 26367
rect 13078 26364 13084 26376
rect 13039 26336 13084 26364
rect 11149 26327 11207 26333
rect 8386 26296 8392 26308
rect 8347 26268 8392 26296
rect 8386 26256 8392 26268
rect 8444 26256 8450 26308
rect 10244 26296 10272 26327
rect 13078 26324 13084 26336
rect 13136 26324 13142 26376
rect 14274 26364 14280 26376
rect 14235 26336 14280 26364
rect 14274 26324 14280 26336
rect 14332 26324 14338 26376
rect 14568 26364 14596 26395
rect 15838 26392 15844 26404
rect 15896 26392 15902 26444
rect 16114 26432 16120 26444
rect 16075 26404 16120 26432
rect 16114 26392 16120 26404
rect 16172 26392 16178 26444
rect 16408 26441 16436 26472
rect 16758 26460 16764 26512
rect 16816 26500 16822 26512
rect 19334 26500 19340 26512
rect 16816 26472 17816 26500
rect 16816 26460 16822 26472
rect 16393 26435 16451 26441
rect 16393 26401 16405 26435
rect 16439 26401 16451 26435
rect 17586 26432 17592 26444
rect 17547 26404 17592 26432
rect 16393 26395 16451 26401
rect 17586 26392 17592 26404
rect 17644 26392 17650 26444
rect 17788 26441 17816 26472
rect 18892 26472 19340 26500
rect 17773 26435 17831 26441
rect 17773 26401 17785 26435
rect 17819 26401 17831 26435
rect 17773 26395 17831 26401
rect 17957 26435 18015 26441
rect 17957 26401 17969 26435
rect 18003 26432 18015 26435
rect 18046 26432 18052 26444
rect 18003 26404 18052 26432
rect 18003 26401 18015 26404
rect 17957 26395 18015 26401
rect 18046 26392 18052 26404
rect 18104 26392 18110 26444
rect 18892 26441 18920 26472
rect 19334 26460 19340 26472
rect 19392 26500 19398 26512
rect 19702 26500 19708 26512
rect 19392 26472 19708 26500
rect 19392 26460 19398 26472
rect 19702 26460 19708 26472
rect 19760 26460 19766 26512
rect 19797 26503 19855 26509
rect 19797 26469 19809 26503
rect 19843 26500 19855 26503
rect 21542 26500 21548 26512
rect 19843 26472 21548 26500
rect 19843 26469 19855 26472
rect 19797 26463 19855 26469
rect 21542 26460 21548 26472
rect 21600 26460 21606 26512
rect 22830 26460 22836 26512
rect 22888 26500 22894 26512
rect 25130 26500 25136 26512
rect 22888 26472 23796 26500
rect 22888 26460 22894 26472
rect 18877 26435 18935 26441
rect 18877 26401 18889 26435
rect 18923 26401 18935 26435
rect 18877 26395 18935 26401
rect 18966 26392 18972 26444
rect 19024 26432 19030 26444
rect 19245 26435 19303 26441
rect 19245 26432 19257 26435
rect 19024 26404 19257 26432
rect 19024 26392 19030 26404
rect 19245 26401 19257 26404
rect 19291 26432 19303 26435
rect 19886 26432 19892 26444
rect 19291 26404 19892 26432
rect 19291 26401 19303 26404
rect 19245 26395 19303 26401
rect 19886 26392 19892 26404
rect 19944 26392 19950 26444
rect 19978 26392 19984 26444
rect 20036 26432 20042 26444
rect 20036 26404 20081 26432
rect 20036 26392 20042 26404
rect 20622 26392 20628 26444
rect 20680 26432 20686 26444
rect 20680 26404 21036 26432
rect 20680 26392 20686 26404
rect 15102 26364 15108 26376
rect 14568 26336 15108 26364
rect 15102 26324 15108 26336
rect 15160 26324 15166 26376
rect 16482 26324 16488 26376
rect 16540 26364 16546 26376
rect 17129 26367 17187 26373
rect 17129 26364 17141 26367
rect 16540 26336 17141 26364
rect 16540 26324 16546 26336
rect 17129 26333 17141 26336
rect 17175 26333 17187 26367
rect 17129 26327 17187 26333
rect 17402 26324 17408 26376
rect 17460 26364 17466 26376
rect 20349 26367 20407 26373
rect 17460 26336 18828 26364
rect 17460 26324 17466 26336
rect 17310 26296 17316 26308
rect 10244 26268 17316 26296
rect 17310 26256 17316 26268
rect 17368 26256 17374 26308
rect 18414 26256 18420 26308
rect 18472 26296 18478 26308
rect 18693 26299 18751 26305
rect 18693 26296 18705 26299
rect 18472 26268 18705 26296
rect 18472 26256 18478 26268
rect 18693 26265 18705 26268
rect 18739 26265 18751 26299
rect 18800 26296 18828 26336
rect 20349 26333 20361 26367
rect 20395 26364 20407 26367
rect 20901 26367 20959 26373
rect 20901 26364 20913 26367
rect 20395 26336 20913 26364
rect 20395 26333 20407 26336
rect 20349 26327 20407 26333
rect 20901 26333 20913 26336
rect 20947 26333 20959 26367
rect 21008 26364 21036 26404
rect 21082 26392 21088 26444
rect 21140 26432 21146 26444
rect 21218 26435 21276 26441
rect 21140 26404 21185 26432
rect 21140 26392 21146 26404
rect 21218 26401 21230 26435
rect 21264 26432 21276 26435
rect 21450 26432 21456 26444
rect 21264 26404 21456 26432
rect 21264 26401 21276 26404
rect 21218 26395 21276 26401
rect 21450 26392 21456 26404
rect 21508 26392 21514 26444
rect 22278 26432 22284 26444
rect 22239 26404 22284 26432
rect 22278 26392 22284 26404
rect 22336 26392 22342 26444
rect 22738 26432 22744 26444
rect 22699 26404 22744 26432
rect 22738 26392 22744 26404
rect 22796 26392 22802 26444
rect 23201 26435 23259 26441
rect 23201 26401 23213 26435
rect 23247 26432 23259 26435
rect 23382 26432 23388 26444
rect 23247 26404 23388 26432
rect 23247 26401 23259 26404
rect 23201 26395 23259 26401
rect 23382 26392 23388 26404
rect 23440 26392 23446 26444
rect 23566 26432 23572 26444
rect 23527 26404 23572 26432
rect 23566 26392 23572 26404
rect 23624 26392 23630 26444
rect 23768 26441 23796 26472
rect 24504 26472 25136 26500
rect 24504 26441 24532 26472
rect 25130 26460 25136 26472
rect 25188 26500 25194 26512
rect 25314 26500 25320 26512
rect 25188 26472 25320 26500
rect 25188 26460 25194 26472
rect 25314 26460 25320 26472
rect 25372 26460 25378 26512
rect 28994 26500 29000 26512
rect 27540 26472 29000 26500
rect 23753 26435 23811 26441
rect 23753 26401 23765 26435
rect 23799 26401 23811 26435
rect 23753 26395 23811 26401
rect 24489 26435 24547 26441
rect 24489 26401 24501 26435
rect 24535 26401 24547 26435
rect 24489 26395 24547 26401
rect 24578 26392 24584 26444
rect 24636 26432 24642 26444
rect 25041 26435 25099 26441
rect 25041 26432 25053 26435
rect 24636 26404 25053 26432
rect 24636 26392 24642 26404
rect 25041 26401 25053 26404
rect 25087 26432 25099 26435
rect 25685 26435 25743 26441
rect 25685 26432 25697 26435
rect 25087 26404 25697 26432
rect 25087 26401 25099 26404
rect 25041 26395 25099 26401
rect 25685 26401 25697 26404
rect 25731 26401 25743 26435
rect 26786 26432 26792 26444
rect 26747 26404 26792 26432
rect 25685 26395 25743 26401
rect 26786 26392 26792 26404
rect 26844 26392 26850 26444
rect 27540 26441 27568 26472
rect 28994 26460 29000 26472
rect 29052 26460 29058 26512
rect 29914 26500 29920 26512
rect 29380 26472 29920 26500
rect 27525 26435 27583 26441
rect 27525 26401 27537 26435
rect 27571 26401 27583 26435
rect 27525 26395 27583 26401
rect 27614 26392 27620 26444
rect 27672 26432 27678 26444
rect 29380 26441 29408 26472
rect 29914 26460 29920 26472
rect 29972 26460 29978 26512
rect 33042 26460 33048 26512
rect 33100 26500 33106 26512
rect 33100 26472 33824 26500
rect 33100 26460 33106 26472
rect 28077 26435 28135 26441
rect 28077 26432 28089 26435
rect 27672 26404 28089 26432
rect 27672 26392 27678 26404
rect 28077 26401 28089 26404
rect 28123 26401 28135 26435
rect 28077 26395 28135 26401
rect 29365 26435 29423 26441
rect 29365 26401 29377 26435
rect 29411 26401 29423 26435
rect 29638 26432 29644 26444
rect 29599 26404 29644 26432
rect 29365 26395 29423 26401
rect 29638 26392 29644 26404
rect 29696 26392 29702 26444
rect 30561 26435 30619 26441
rect 30561 26401 30573 26435
rect 30607 26432 30619 26435
rect 31018 26432 31024 26444
rect 30607 26404 31024 26432
rect 30607 26401 30619 26404
rect 30561 26395 30619 26401
rect 31018 26392 31024 26404
rect 31076 26392 31082 26444
rect 31113 26435 31171 26441
rect 31113 26401 31125 26435
rect 31159 26432 31171 26435
rect 32030 26432 32036 26444
rect 31159 26404 32036 26432
rect 31159 26401 31171 26404
rect 31113 26395 31171 26401
rect 32030 26392 32036 26404
rect 32088 26392 32094 26444
rect 32214 26432 32220 26444
rect 32175 26404 32220 26432
rect 32214 26392 32220 26404
rect 32272 26392 32278 26444
rect 32950 26432 32956 26444
rect 32911 26404 32956 26432
rect 32950 26392 32956 26404
rect 33008 26392 33014 26444
rect 33796 26441 33824 26472
rect 35544 26472 37780 26500
rect 33781 26435 33839 26441
rect 33781 26401 33793 26435
rect 33827 26401 33839 26435
rect 33781 26395 33839 26401
rect 34609 26435 34667 26441
rect 34609 26401 34621 26435
rect 34655 26401 34667 26435
rect 34609 26395 34667 26401
rect 21008 26336 22968 26364
rect 20901 26327 20959 26333
rect 22940 26308 22968 26336
rect 23658 26324 23664 26376
rect 23716 26364 23722 26376
rect 24762 26364 24768 26376
rect 23716 26336 24768 26364
rect 23716 26324 23722 26336
rect 24762 26324 24768 26336
rect 24820 26364 24826 26376
rect 24949 26367 25007 26373
rect 24949 26364 24961 26367
rect 24820 26336 24961 26364
rect 24820 26324 24826 26336
rect 24949 26333 24961 26336
rect 24995 26333 25007 26367
rect 24949 26327 25007 26333
rect 28537 26367 28595 26373
rect 28537 26333 28549 26367
rect 28583 26364 28595 26367
rect 29270 26364 29276 26376
rect 28583 26336 29276 26364
rect 28583 26333 28595 26336
rect 28537 26327 28595 26333
rect 29270 26324 29276 26336
rect 29328 26324 29334 26376
rect 30742 26324 30748 26376
rect 30800 26364 30806 26376
rect 31205 26367 31263 26373
rect 31205 26364 31217 26367
rect 30800 26336 31217 26364
rect 30800 26324 30806 26336
rect 31205 26333 31217 26336
rect 31251 26333 31263 26367
rect 31205 26327 31263 26333
rect 31478 26324 31484 26376
rect 31536 26364 31542 26376
rect 33045 26367 33103 26373
rect 33045 26364 33057 26367
rect 31536 26336 33057 26364
rect 31536 26324 31542 26336
rect 33045 26333 33057 26336
rect 33091 26333 33103 26367
rect 34624 26364 34652 26395
rect 34698 26392 34704 26444
rect 34756 26432 34762 26444
rect 34885 26435 34943 26441
rect 34885 26432 34897 26435
rect 34756 26404 34897 26432
rect 34756 26392 34762 26404
rect 34885 26401 34897 26404
rect 34931 26401 34943 26435
rect 34885 26395 34943 26401
rect 35342 26392 35348 26444
rect 35400 26432 35406 26444
rect 35544 26441 35572 26472
rect 35529 26435 35587 26441
rect 35529 26432 35541 26435
rect 35400 26404 35541 26432
rect 35400 26392 35406 26404
rect 35529 26401 35541 26404
rect 35575 26401 35587 26435
rect 35529 26395 35587 26401
rect 35986 26392 35992 26444
rect 36044 26432 36050 26444
rect 36633 26435 36691 26441
rect 36633 26432 36645 26435
rect 36044 26404 36645 26432
rect 36044 26392 36050 26404
rect 36633 26401 36645 26404
rect 36679 26401 36691 26435
rect 36814 26432 36820 26444
rect 36775 26404 36820 26432
rect 36633 26395 36691 26401
rect 36814 26392 36820 26404
rect 36872 26392 36878 26444
rect 36998 26432 37004 26444
rect 36959 26404 37004 26432
rect 36998 26392 37004 26404
rect 37056 26392 37062 26444
rect 37752 26441 37780 26472
rect 37737 26435 37795 26441
rect 37737 26401 37749 26435
rect 37783 26401 37795 26435
rect 37737 26395 37795 26401
rect 34790 26364 34796 26376
rect 34624 26336 34796 26364
rect 33045 26327 33103 26333
rect 34790 26324 34796 26336
rect 34848 26324 34854 26376
rect 36832 26364 36860 26392
rect 37829 26367 37887 26373
rect 37829 26364 37841 26367
rect 36832 26336 37841 26364
rect 37829 26333 37841 26336
rect 37875 26333 37887 26367
rect 37829 26327 37887 26333
rect 21082 26296 21088 26308
rect 18800 26268 21088 26296
rect 18693 26259 18751 26265
rect 21082 26256 21088 26268
rect 21140 26256 21146 26308
rect 21266 26256 21272 26308
rect 21324 26296 21330 26308
rect 22002 26296 22008 26308
rect 21324 26268 22008 26296
rect 21324 26256 21330 26268
rect 22002 26256 22008 26268
rect 22060 26296 22066 26308
rect 22646 26296 22652 26308
rect 22060 26268 22652 26296
rect 22060 26256 22066 26268
rect 22646 26256 22652 26268
rect 22704 26256 22710 26308
rect 22922 26256 22928 26308
rect 22980 26256 22986 26308
rect 27801 26299 27859 26305
rect 27801 26265 27813 26299
rect 27847 26296 27859 26299
rect 28166 26296 28172 26308
rect 27847 26268 28172 26296
rect 27847 26265 27859 26268
rect 27801 26259 27859 26265
rect 28166 26256 28172 26268
rect 28224 26256 28230 26308
rect 28442 26256 28448 26308
rect 28500 26296 28506 26308
rect 29181 26299 29239 26305
rect 29181 26296 29193 26299
rect 28500 26268 29193 26296
rect 28500 26256 28506 26268
rect 29181 26265 29193 26268
rect 29227 26265 29239 26299
rect 30650 26296 30656 26308
rect 30611 26268 30656 26296
rect 29181 26259 29239 26265
rect 30650 26256 30656 26268
rect 30708 26256 30714 26308
rect 36449 26299 36507 26305
rect 36449 26265 36461 26299
rect 36495 26296 36507 26299
rect 37734 26296 37740 26308
rect 36495 26268 37740 26296
rect 36495 26265 36507 26268
rect 36449 26259 36507 26265
rect 37734 26256 37740 26268
rect 37792 26256 37798 26308
rect 4798 26228 4804 26240
rect 4448 26200 4804 26228
rect 4798 26188 4804 26200
rect 4856 26188 4862 26240
rect 4890 26188 4896 26240
rect 4948 26228 4954 26240
rect 6454 26228 6460 26240
rect 4948 26200 6460 26228
rect 4948 26188 4954 26200
rect 6454 26188 6460 26200
rect 6512 26228 6518 26240
rect 7377 26231 7435 26237
rect 7377 26228 7389 26231
rect 6512 26200 7389 26228
rect 6512 26188 6518 26200
rect 7377 26197 7389 26200
rect 7423 26197 7435 26231
rect 7377 26191 7435 26197
rect 9858 26188 9864 26240
rect 9916 26228 9922 26240
rect 13078 26228 13084 26240
rect 9916 26200 13084 26228
rect 9916 26188 9922 26200
rect 13078 26188 13084 26200
rect 13136 26188 13142 26240
rect 17586 26188 17592 26240
rect 17644 26228 17650 26240
rect 18230 26228 18236 26240
rect 17644 26200 18236 26228
rect 17644 26188 17650 26200
rect 18230 26188 18236 26200
rect 18288 26188 18294 26240
rect 20990 26188 20996 26240
rect 21048 26228 21054 26240
rect 21361 26231 21419 26237
rect 21361 26228 21373 26231
rect 21048 26200 21373 26228
rect 21048 26188 21054 26200
rect 21361 26197 21373 26200
rect 21407 26197 21419 26231
rect 22186 26228 22192 26240
rect 22147 26200 22192 26228
rect 21361 26191 21419 26197
rect 22186 26188 22192 26200
rect 22244 26188 22250 26240
rect 33962 26228 33968 26240
rect 33923 26200 33968 26228
rect 33962 26188 33968 26200
rect 34020 26188 34026 26240
rect 34606 26228 34612 26240
rect 34567 26200 34612 26228
rect 34606 26188 34612 26200
rect 34664 26188 34670 26240
rect 1104 26138 38824 26160
rect 1104 26086 4246 26138
rect 4298 26086 4310 26138
rect 4362 26086 4374 26138
rect 4426 26086 4438 26138
rect 4490 26086 34966 26138
rect 35018 26086 35030 26138
rect 35082 26086 35094 26138
rect 35146 26086 35158 26138
rect 35210 26086 38824 26138
rect 1104 26064 38824 26086
rect 1949 26027 2007 26033
rect 1949 25993 1961 26027
rect 1995 26024 2007 26027
rect 3970 26024 3976 26036
rect 1995 25996 3976 26024
rect 1995 25993 2007 25996
rect 1949 25987 2007 25993
rect 3970 25984 3976 25996
rect 4028 25984 4034 26036
rect 12529 26027 12587 26033
rect 12529 25993 12541 26027
rect 12575 26024 12587 26027
rect 12618 26024 12624 26036
rect 12575 25996 12624 26024
rect 12575 25993 12587 25996
rect 12529 25987 12587 25993
rect 12618 25984 12624 25996
rect 12676 25984 12682 26036
rect 16761 26027 16819 26033
rect 16761 25993 16773 26027
rect 16807 26024 16819 26027
rect 18322 26024 18328 26036
rect 16807 25996 18328 26024
rect 16807 25993 16819 25996
rect 16761 25987 16819 25993
rect 18322 25984 18328 25996
rect 18380 25984 18386 26036
rect 20993 26027 21051 26033
rect 20993 25993 21005 26027
rect 21039 26024 21051 26027
rect 21450 26024 21456 26036
rect 21039 25996 21456 26024
rect 21039 25993 21051 25996
rect 20993 25987 21051 25993
rect 21450 25984 21456 25996
rect 21508 25984 21514 26036
rect 23750 26024 23756 26036
rect 22848 25996 23756 26024
rect 1854 25916 1860 25968
rect 1912 25956 1918 25968
rect 5353 25959 5411 25965
rect 5353 25956 5365 25959
rect 1912 25928 5365 25956
rect 1912 25916 1918 25928
rect 5353 25925 5365 25928
rect 5399 25925 5411 25959
rect 7742 25956 7748 25968
rect 7703 25928 7748 25956
rect 5353 25919 5411 25925
rect 7742 25916 7748 25928
rect 7800 25916 7806 25968
rect 15378 25956 15384 25968
rect 15339 25928 15384 25956
rect 15378 25916 15384 25928
rect 15436 25916 15442 25968
rect 17770 25916 17776 25968
rect 17828 25956 17834 25968
rect 17828 25928 22416 25956
rect 17828 25916 17834 25928
rect 1762 25848 1768 25900
rect 1820 25888 1826 25900
rect 2593 25891 2651 25897
rect 2593 25888 2605 25891
rect 1820 25860 2605 25888
rect 1820 25848 1826 25860
rect 1872 25829 1900 25860
rect 2593 25857 2605 25860
rect 2639 25857 2651 25891
rect 4614 25888 4620 25900
rect 4575 25860 4620 25888
rect 2593 25851 2651 25857
rect 4614 25848 4620 25860
rect 4672 25848 4678 25900
rect 8570 25848 8576 25900
rect 8628 25888 8634 25900
rect 10873 25891 10931 25897
rect 8628 25860 8984 25888
rect 8628 25848 8634 25860
rect 1857 25823 1915 25829
rect 1857 25789 1869 25823
rect 1903 25789 1915 25823
rect 2682 25820 2688 25832
rect 2643 25792 2688 25820
rect 1857 25783 1915 25789
rect 2682 25780 2688 25792
rect 2740 25780 2746 25832
rect 3142 25820 3148 25832
rect 3103 25792 3148 25820
rect 3142 25780 3148 25792
rect 3200 25780 3206 25832
rect 3234 25780 3240 25832
rect 3292 25820 3298 25832
rect 3292 25792 3337 25820
rect 3292 25780 3298 25792
rect 3970 25780 3976 25832
rect 4028 25820 4034 25832
rect 4157 25823 4215 25829
rect 4157 25820 4169 25823
rect 4028 25792 4169 25820
rect 4028 25780 4034 25792
rect 4157 25789 4169 25792
rect 4203 25789 4215 25823
rect 4157 25783 4215 25789
rect 4341 25823 4399 25829
rect 4341 25789 4353 25823
rect 4387 25820 4399 25823
rect 4706 25820 4712 25832
rect 4387 25792 4712 25820
rect 4387 25789 4399 25792
rect 4341 25783 4399 25789
rect 4706 25780 4712 25792
rect 4764 25780 4770 25832
rect 5166 25820 5172 25832
rect 5127 25792 5172 25820
rect 5166 25780 5172 25792
rect 5224 25780 5230 25832
rect 5626 25780 5632 25832
rect 5684 25820 5690 25832
rect 5905 25823 5963 25829
rect 5905 25820 5917 25823
rect 5684 25792 5917 25820
rect 5684 25780 5690 25792
rect 5905 25789 5917 25792
rect 5951 25789 5963 25823
rect 5905 25783 5963 25789
rect 6917 25823 6975 25829
rect 6917 25789 6929 25823
rect 6963 25820 6975 25823
rect 7006 25820 7012 25832
rect 6963 25792 7012 25820
rect 6963 25789 6975 25792
rect 6917 25783 6975 25789
rect 7006 25780 7012 25792
rect 7064 25780 7070 25832
rect 7926 25820 7932 25832
rect 7887 25792 7932 25820
rect 7926 25780 7932 25792
rect 7984 25780 7990 25832
rect 8386 25820 8392 25832
rect 8347 25792 8392 25820
rect 8386 25780 8392 25792
rect 8444 25780 8450 25832
rect 8846 25820 8852 25832
rect 8807 25792 8852 25820
rect 8846 25780 8852 25792
rect 8904 25780 8910 25832
rect 8956 25829 8984 25860
rect 10873 25857 10885 25891
rect 10919 25888 10931 25891
rect 12526 25888 12532 25900
rect 10919 25860 12532 25888
rect 10919 25857 10931 25860
rect 10873 25851 10931 25857
rect 12526 25848 12532 25860
rect 12584 25888 12590 25900
rect 13538 25888 13544 25900
rect 12584 25860 13544 25888
rect 12584 25848 12590 25860
rect 13538 25848 13544 25860
rect 13596 25848 13602 25900
rect 14642 25888 14648 25900
rect 14603 25860 14648 25888
rect 14642 25848 14648 25860
rect 14700 25848 14706 25900
rect 16942 25848 16948 25900
rect 17000 25888 17006 25900
rect 18049 25891 18107 25897
rect 18049 25888 18061 25891
rect 17000 25860 18061 25888
rect 17000 25848 17006 25860
rect 18049 25857 18061 25860
rect 18095 25857 18107 25891
rect 18049 25851 18107 25857
rect 18230 25848 18236 25900
rect 18288 25888 18294 25900
rect 18288 25860 18552 25888
rect 18288 25848 18294 25860
rect 8941 25823 8999 25829
rect 8941 25789 8953 25823
rect 8987 25789 8999 25823
rect 8941 25783 8999 25789
rect 9309 25823 9367 25829
rect 9309 25789 9321 25823
rect 9355 25789 9367 25823
rect 9309 25783 9367 25789
rect 8754 25712 8760 25764
rect 8812 25752 8818 25764
rect 9324 25752 9352 25783
rect 9858 25780 9864 25832
rect 9916 25820 9922 25832
rect 10045 25823 10103 25829
rect 10045 25820 10057 25823
rect 9916 25792 10057 25820
rect 9916 25780 9922 25792
rect 10045 25789 10057 25792
rect 10091 25789 10103 25823
rect 12437 25823 12495 25829
rect 12437 25820 12449 25823
rect 10045 25783 10103 25789
rect 11256 25792 12449 25820
rect 11256 25764 11284 25792
rect 12437 25789 12449 25792
rect 12483 25789 12495 25823
rect 12437 25783 12495 25789
rect 13725 25823 13783 25829
rect 13725 25789 13737 25823
rect 13771 25820 13783 25823
rect 13814 25820 13820 25832
rect 13771 25792 13820 25820
rect 13771 25789 13783 25792
rect 13725 25783 13783 25789
rect 13814 25780 13820 25792
rect 13872 25780 13878 25832
rect 13909 25823 13967 25829
rect 13909 25789 13921 25823
rect 13955 25789 13967 25823
rect 14366 25820 14372 25832
rect 14327 25792 14372 25820
rect 13909 25783 13967 25789
rect 11238 25752 11244 25764
rect 8812 25724 10272 25752
rect 11199 25724 11244 25752
rect 8812 25712 8818 25724
rect 5994 25684 6000 25696
rect 5955 25656 6000 25684
rect 5994 25644 6000 25656
rect 6052 25644 6058 25696
rect 7101 25687 7159 25693
rect 7101 25653 7113 25687
rect 7147 25684 7159 25687
rect 8386 25684 8392 25696
rect 7147 25656 8392 25684
rect 7147 25653 7159 25656
rect 7101 25647 7159 25653
rect 8386 25644 8392 25656
rect 8444 25644 8450 25696
rect 10244 25693 10272 25724
rect 11238 25712 11244 25724
rect 11296 25712 11302 25764
rect 11606 25752 11612 25764
rect 11567 25724 11612 25752
rect 11606 25712 11612 25724
rect 11664 25712 11670 25764
rect 13446 25712 13452 25764
rect 13504 25752 13510 25764
rect 13924 25752 13952 25783
rect 14366 25780 14372 25792
rect 14424 25780 14430 25832
rect 15565 25823 15623 25829
rect 15565 25789 15577 25823
rect 15611 25789 15623 25823
rect 15565 25783 15623 25789
rect 13504 25724 13952 25752
rect 13504 25712 13510 25724
rect 10229 25687 10287 25693
rect 10229 25653 10241 25687
rect 10275 25653 10287 25687
rect 11054 25684 11060 25696
rect 11015 25656 11060 25684
rect 10229 25647 10287 25653
rect 11054 25644 11060 25656
rect 11112 25644 11118 25696
rect 11146 25644 11152 25696
rect 11204 25684 11210 25696
rect 11882 25684 11888 25696
rect 11204 25656 11888 25684
rect 11204 25644 11210 25656
rect 11882 25644 11888 25656
rect 11940 25644 11946 25696
rect 15580 25684 15608 25783
rect 15654 25780 15660 25832
rect 15712 25820 15718 25832
rect 15749 25823 15807 25829
rect 15749 25820 15761 25823
rect 15712 25792 15761 25820
rect 15712 25780 15718 25792
rect 15749 25789 15761 25792
rect 15795 25789 15807 25823
rect 15749 25783 15807 25789
rect 15933 25823 15991 25829
rect 15933 25789 15945 25823
rect 15979 25820 15991 25823
rect 16114 25820 16120 25832
rect 15979 25792 16120 25820
rect 15979 25789 15991 25792
rect 15933 25783 15991 25789
rect 16114 25780 16120 25792
rect 16172 25780 16178 25832
rect 17037 25823 17095 25829
rect 17037 25789 17049 25823
rect 17083 25820 17095 25823
rect 18414 25820 18420 25832
rect 17083 25792 18420 25820
rect 17083 25789 17095 25792
rect 17037 25783 17095 25789
rect 18414 25780 18420 25792
rect 18472 25780 18478 25832
rect 18524 25829 18552 25860
rect 18598 25848 18604 25900
rect 18656 25888 18662 25900
rect 18656 25860 18736 25888
rect 18656 25848 18662 25860
rect 18708 25829 18736 25860
rect 19978 25848 19984 25900
rect 20036 25888 20042 25900
rect 21266 25888 21272 25900
rect 20036 25860 21272 25888
rect 20036 25848 20042 25860
rect 18509 25823 18567 25829
rect 18509 25789 18521 25823
rect 18555 25789 18567 25823
rect 18509 25783 18567 25789
rect 18693 25823 18751 25829
rect 18693 25789 18705 25823
rect 18739 25789 18751 25823
rect 18693 25783 18751 25789
rect 18877 25823 18935 25829
rect 18877 25789 18889 25823
rect 18923 25789 18935 25823
rect 19886 25820 19892 25832
rect 19847 25792 19892 25820
rect 18877 25783 18935 25789
rect 16945 25755 17003 25761
rect 16945 25721 16957 25755
rect 16991 25752 17003 25755
rect 17402 25752 17408 25764
rect 16991 25724 17408 25752
rect 16991 25721 17003 25724
rect 16945 25715 17003 25721
rect 17402 25712 17408 25724
rect 17460 25712 17466 25764
rect 17497 25755 17555 25761
rect 17497 25721 17509 25755
rect 17543 25752 17555 25755
rect 17954 25752 17960 25764
rect 17543 25724 17960 25752
rect 17543 25721 17555 25724
rect 17497 25715 17555 25721
rect 17954 25712 17960 25724
rect 18012 25712 18018 25764
rect 15838 25684 15844 25696
rect 15580 25656 15844 25684
rect 15838 25644 15844 25656
rect 15896 25684 15902 25696
rect 16850 25684 16856 25696
rect 15896 25656 16856 25684
rect 15896 25644 15902 25656
rect 16850 25644 16856 25656
rect 16908 25684 16914 25696
rect 18892 25684 18920 25783
rect 19886 25780 19892 25792
rect 19944 25780 19950 25832
rect 20254 25820 20260 25832
rect 20215 25792 20260 25820
rect 20254 25780 20260 25792
rect 20312 25780 20318 25832
rect 20640 25829 20668 25860
rect 21266 25848 21272 25860
rect 21324 25848 21330 25900
rect 22186 25888 22192 25900
rect 22147 25860 22192 25888
rect 22186 25848 22192 25860
rect 22244 25848 22250 25900
rect 20625 25823 20683 25829
rect 20625 25789 20637 25823
rect 20671 25789 20683 25823
rect 20898 25820 20904 25832
rect 20859 25792 20904 25820
rect 20625 25783 20683 25789
rect 20898 25780 20904 25792
rect 20956 25780 20962 25832
rect 20990 25780 20996 25832
rect 21048 25820 21054 25832
rect 22388 25829 22416 25928
rect 21913 25823 21971 25829
rect 21913 25820 21925 25823
rect 21048 25792 21925 25820
rect 21048 25780 21054 25792
rect 21913 25789 21925 25792
rect 21959 25789 21971 25823
rect 21913 25783 21971 25789
rect 22373 25823 22431 25829
rect 22373 25789 22385 25823
rect 22419 25789 22431 25823
rect 22373 25783 22431 25789
rect 16908 25656 18920 25684
rect 21729 25687 21787 25693
rect 16908 25644 16914 25656
rect 21729 25653 21741 25687
rect 21775 25684 21787 25687
rect 22848 25684 22876 25996
rect 23750 25984 23756 25996
rect 23808 26024 23814 26036
rect 25038 26024 25044 26036
rect 23808 25996 25044 26024
rect 23808 25984 23814 25996
rect 25038 25984 25044 25996
rect 25096 25984 25102 26036
rect 25682 25984 25688 26036
rect 25740 26024 25746 26036
rect 28629 26027 28687 26033
rect 28629 26024 28641 26027
rect 25740 25996 28641 26024
rect 25740 25984 25746 25996
rect 28629 25993 28641 25996
rect 28675 25993 28687 26027
rect 28629 25987 28687 25993
rect 32030 25984 32036 26036
rect 32088 26024 32094 26036
rect 32585 26027 32643 26033
rect 32585 26024 32597 26027
rect 32088 25996 32597 26024
rect 32088 25984 32094 25996
rect 32585 25993 32597 25996
rect 32631 25993 32643 26027
rect 32585 25987 32643 25993
rect 34241 26027 34299 26033
rect 34241 25993 34253 26027
rect 34287 26024 34299 26027
rect 34422 26024 34428 26036
rect 34287 25996 34428 26024
rect 34287 25993 34299 25996
rect 34241 25987 34299 25993
rect 34422 25984 34428 25996
rect 34480 25984 34486 26036
rect 35342 26024 35348 26036
rect 35303 25996 35348 26024
rect 35342 25984 35348 25996
rect 35400 25984 35406 26036
rect 23937 25959 23995 25965
rect 23937 25956 23949 25959
rect 22940 25928 23949 25956
rect 22940 25829 22968 25928
rect 23937 25925 23949 25928
rect 23983 25925 23995 25959
rect 26418 25956 26424 25968
rect 23937 25919 23995 25925
rect 24136 25928 26424 25956
rect 23109 25891 23167 25897
rect 23109 25857 23121 25891
rect 23155 25888 23167 25891
rect 24136 25888 24164 25928
rect 26418 25916 26424 25928
rect 26476 25916 26482 25968
rect 26697 25891 26755 25897
rect 23155 25860 24164 25888
rect 24228 25860 26648 25888
rect 23155 25857 23167 25860
rect 23109 25851 23167 25857
rect 22925 25823 22983 25829
rect 22925 25789 22937 25823
rect 22971 25789 22983 25823
rect 23658 25820 23664 25832
rect 23619 25792 23664 25820
rect 22925 25783 22983 25789
rect 23658 25780 23664 25792
rect 23716 25780 23722 25832
rect 21775 25656 22876 25684
rect 21775 25653 21787 25656
rect 21729 25647 21787 25653
rect 23014 25644 23020 25696
rect 23072 25684 23078 25696
rect 24228 25684 24256 25860
rect 24394 25820 24400 25832
rect 24355 25792 24400 25820
rect 24394 25780 24400 25792
rect 24452 25780 24458 25832
rect 24670 25820 24676 25832
rect 24631 25792 24676 25820
rect 24670 25780 24676 25792
rect 24728 25780 24734 25832
rect 24762 25780 24768 25832
rect 24820 25820 24826 25832
rect 25409 25823 25467 25829
rect 25409 25820 25421 25823
rect 24820 25792 25421 25820
rect 24820 25780 24826 25792
rect 25409 25789 25421 25792
rect 25455 25789 25467 25823
rect 25409 25783 25467 25789
rect 26421 25823 26479 25829
rect 26421 25789 26433 25823
rect 26467 25820 26479 25823
rect 26510 25820 26516 25832
rect 26467 25792 26516 25820
rect 26467 25789 26479 25792
rect 26421 25783 26479 25789
rect 26510 25780 26516 25792
rect 26568 25780 26574 25832
rect 26620 25820 26648 25860
rect 26697 25857 26709 25891
rect 26743 25888 26755 25891
rect 27982 25888 27988 25900
rect 26743 25860 27988 25888
rect 26743 25857 26755 25860
rect 26697 25851 26755 25857
rect 27982 25848 27988 25860
rect 28040 25848 28046 25900
rect 30282 25848 30288 25900
rect 30340 25888 30346 25900
rect 30377 25891 30435 25897
rect 30377 25888 30389 25891
rect 30340 25860 30389 25888
rect 30340 25848 30346 25860
rect 30377 25857 30389 25860
rect 30423 25857 30435 25891
rect 30650 25888 30656 25900
rect 30611 25860 30656 25888
rect 30377 25851 30435 25857
rect 30650 25848 30656 25860
rect 30708 25848 30714 25900
rect 31754 25848 31760 25900
rect 31812 25888 31818 25900
rect 33962 25888 33968 25900
rect 31812 25860 33968 25888
rect 31812 25848 31818 25860
rect 28077 25823 28135 25829
rect 26620 25792 27384 25820
rect 27356 25752 27384 25792
rect 28077 25789 28089 25823
rect 28123 25820 28135 25823
rect 28537 25823 28595 25829
rect 28537 25820 28549 25823
rect 28123 25792 28549 25820
rect 28123 25789 28135 25792
rect 28077 25783 28135 25789
rect 28537 25789 28549 25792
rect 28583 25820 28595 25823
rect 29270 25820 29276 25832
rect 28583 25792 29276 25820
rect 28583 25789 28595 25792
rect 28537 25783 28595 25789
rect 29270 25780 29276 25792
rect 29328 25780 29334 25832
rect 29641 25823 29699 25829
rect 29641 25789 29653 25823
rect 29687 25789 29699 25823
rect 29641 25783 29699 25789
rect 32033 25823 32091 25829
rect 32033 25789 32045 25823
rect 32079 25820 32091 25823
rect 32490 25820 32496 25832
rect 32079 25792 32496 25820
rect 32079 25789 32091 25792
rect 32033 25783 32091 25789
rect 29656 25752 29684 25783
rect 32490 25780 32496 25792
rect 32548 25780 32554 25832
rect 32876 25829 32904 25860
rect 33962 25848 33968 25860
rect 34020 25848 34026 25900
rect 34514 25848 34520 25900
rect 34572 25888 34578 25900
rect 34572 25860 36124 25888
rect 34572 25848 34578 25860
rect 32861 25823 32919 25829
rect 32861 25789 32873 25823
rect 32907 25789 32919 25823
rect 33410 25820 33416 25832
rect 33371 25792 33416 25820
rect 32861 25783 32919 25789
rect 33410 25780 33416 25792
rect 33468 25780 33474 25832
rect 34149 25823 34207 25829
rect 34149 25789 34161 25823
rect 34195 25820 34207 25823
rect 34606 25820 34612 25832
rect 34195 25792 34612 25820
rect 34195 25789 34207 25792
rect 34149 25783 34207 25789
rect 34606 25780 34612 25792
rect 34664 25780 34670 25832
rect 35526 25820 35532 25832
rect 35487 25792 35532 25820
rect 35526 25780 35532 25792
rect 35584 25780 35590 25832
rect 35989 25823 36047 25829
rect 35989 25789 36001 25823
rect 36035 25789 36047 25823
rect 35989 25783 36047 25789
rect 27356 25724 29684 25752
rect 23072 25656 24256 25684
rect 23072 25644 23078 25656
rect 24486 25644 24492 25696
rect 24544 25684 24550 25696
rect 25593 25687 25651 25693
rect 25593 25684 25605 25687
rect 24544 25656 25605 25684
rect 24544 25644 24550 25656
rect 25593 25653 25605 25656
rect 25639 25653 25651 25687
rect 25593 25647 25651 25653
rect 29825 25687 29883 25693
rect 29825 25653 29837 25687
rect 29871 25684 29883 25687
rect 31110 25684 31116 25696
rect 29871 25656 31116 25684
rect 29871 25653 29883 25656
rect 29825 25647 29883 25653
rect 31110 25644 31116 25656
rect 31168 25644 31174 25696
rect 36004 25684 36032 25783
rect 36096 25752 36124 25860
rect 36354 25780 36360 25832
rect 36412 25820 36418 25832
rect 36449 25823 36507 25829
rect 36449 25820 36461 25823
rect 36412 25792 36461 25820
rect 36412 25780 36418 25792
rect 36449 25789 36461 25792
rect 36495 25789 36507 25823
rect 36725 25823 36783 25829
rect 36725 25820 36737 25823
rect 36449 25783 36507 25789
rect 36556 25792 36737 25820
rect 36556 25752 36584 25792
rect 36725 25789 36737 25792
rect 36771 25789 36783 25823
rect 36725 25783 36783 25789
rect 36096 25724 36584 25752
rect 36538 25684 36544 25696
rect 36004 25656 36544 25684
rect 36538 25644 36544 25656
rect 36596 25684 36602 25696
rect 37829 25687 37887 25693
rect 37829 25684 37841 25687
rect 36596 25656 37841 25684
rect 36596 25644 36602 25656
rect 37829 25653 37841 25656
rect 37875 25653 37887 25687
rect 37829 25647 37887 25653
rect 1104 25594 38824 25616
rect 1104 25542 19606 25594
rect 19658 25542 19670 25594
rect 19722 25542 19734 25594
rect 19786 25542 19798 25594
rect 19850 25542 38824 25594
rect 1104 25520 38824 25542
rect 3234 25440 3240 25492
rect 3292 25480 3298 25492
rect 4249 25483 4307 25489
rect 4249 25480 4261 25483
rect 3292 25452 4261 25480
rect 3292 25440 3298 25452
rect 4249 25449 4261 25452
rect 4295 25449 4307 25483
rect 4249 25443 4307 25449
rect 7006 25440 7012 25492
rect 7064 25480 7070 25492
rect 8021 25483 8079 25489
rect 8021 25480 8033 25483
rect 7064 25452 8033 25480
rect 7064 25440 7070 25452
rect 8021 25449 8033 25452
rect 8067 25480 8079 25483
rect 11146 25480 11152 25492
rect 8067 25452 11152 25480
rect 8067 25449 8079 25452
rect 8021 25443 8079 25449
rect 11146 25440 11152 25452
rect 11204 25440 11210 25492
rect 15654 25480 15660 25492
rect 11900 25452 15660 25480
rect 11238 25372 11244 25424
rect 11296 25412 11302 25424
rect 11296 25384 11836 25412
rect 11296 25372 11302 25384
rect 1394 25344 1400 25356
rect 1307 25316 1400 25344
rect 1394 25304 1400 25316
rect 1452 25344 1458 25356
rect 2682 25344 2688 25356
rect 1452 25316 2688 25344
rect 1452 25304 1458 25316
rect 2682 25304 2688 25316
rect 2740 25304 2746 25356
rect 4062 25344 4068 25356
rect 4023 25316 4068 25344
rect 4062 25304 4068 25316
rect 4120 25304 4126 25356
rect 5445 25347 5503 25353
rect 5445 25313 5457 25347
rect 5491 25313 5503 25347
rect 5626 25344 5632 25356
rect 5587 25316 5632 25344
rect 5445 25307 5503 25313
rect 1670 25276 1676 25288
rect 1631 25248 1676 25276
rect 1670 25236 1676 25248
rect 1728 25236 1734 25288
rect 5460 25276 5488 25307
rect 5626 25304 5632 25316
rect 5684 25304 5690 25356
rect 5997 25347 6055 25353
rect 5997 25313 6009 25347
rect 6043 25344 6055 25347
rect 7006 25344 7012 25356
rect 6043 25316 7012 25344
rect 6043 25313 6055 25316
rect 5997 25307 6055 25313
rect 7006 25304 7012 25316
rect 7064 25304 7070 25356
rect 8573 25347 8631 25353
rect 8573 25313 8585 25347
rect 8619 25344 8631 25347
rect 11606 25344 11612 25356
rect 8619 25316 11612 25344
rect 8619 25313 8631 25316
rect 8573 25307 8631 25313
rect 11606 25304 11612 25316
rect 11664 25304 11670 25356
rect 11808 25353 11836 25384
rect 11793 25347 11851 25353
rect 11793 25313 11805 25347
rect 11839 25313 11851 25347
rect 11793 25307 11851 25313
rect 5534 25276 5540 25288
rect 5460 25248 5540 25276
rect 5534 25236 5540 25248
rect 5592 25236 5598 25288
rect 6457 25279 6515 25285
rect 6457 25245 6469 25279
rect 6503 25245 6515 25279
rect 6457 25239 6515 25245
rect 6733 25279 6791 25285
rect 6733 25245 6745 25279
rect 6779 25276 6791 25279
rect 7190 25276 7196 25288
rect 6779 25248 7196 25276
rect 6779 25245 6791 25248
rect 6733 25239 6791 25245
rect 4706 25168 4712 25220
rect 4764 25208 4770 25220
rect 6472 25208 6500 25239
rect 7190 25236 7196 25248
rect 7248 25236 7254 25288
rect 9674 25236 9680 25288
rect 9732 25276 9738 25288
rect 9950 25276 9956 25288
rect 9732 25248 9777 25276
rect 9911 25248 9956 25276
rect 9732 25236 9738 25248
rect 9950 25236 9956 25248
rect 10008 25236 10014 25288
rect 11900 25276 11928 25452
rect 15654 25440 15660 25452
rect 15712 25440 15718 25492
rect 15838 25480 15844 25492
rect 15799 25452 15844 25480
rect 15838 25440 15844 25452
rect 15896 25440 15902 25492
rect 18046 25480 18052 25492
rect 15948 25452 18052 25480
rect 12618 25344 12624 25356
rect 12579 25316 12624 25344
rect 12618 25304 12624 25316
rect 12676 25304 12682 25356
rect 15194 25304 15200 25356
rect 15252 25344 15258 25356
rect 15657 25347 15715 25353
rect 15657 25344 15669 25347
rect 15252 25316 15669 25344
rect 15252 25304 15258 25316
rect 15657 25313 15669 25316
rect 15703 25344 15715 25347
rect 15948 25344 15976 25452
rect 16022 25372 16028 25424
rect 16080 25412 16086 25424
rect 16080 25384 17080 25412
rect 16080 25372 16086 25384
rect 16850 25344 16856 25356
rect 15703 25316 15976 25344
rect 16811 25316 16856 25344
rect 15703 25313 15715 25316
rect 15657 25307 15715 25313
rect 16850 25304 16856 25316
rect 16908 25304 16914 25356
rect 17052 25353 17080 25384
rect 17236 25353 17264 25452
rect 18046 25440 18052 25452
rect 18104 25440 18110 25492
rect 22278 25480 22284 25492
rect 21744 25452 22284 25480
rect 17037 25347 17095 25353
rect 17037 25313 17049 25347
rect 17083 25313 17095 25347
rect 17037 25307 17095 25313
rect 17221 25347 17279 25353
rect 17221 25313 17233 25347
rect 17267 25313 17279 25347
rect 17221 25307 17279 25313
rect 17310 25304 17316 25356
rect 17368 25344 17374 25356
rect 17865 25347 17923 25353
rect 17865 25344 17877 25347
rect 17368 25316 17877 25344
rect 17368 25304 17374 25316
rect 17865 25313 17877 25316
rect 17911 25313 17923 25347
rect 17865 25307 17923 25313
rect 17954 25304 17960 25356
rect 18012 25344 18018 25356
rect 18785 25347 18843 25353
rect 18785 25344 18797 25347
rect 18012 25316 18797 25344
rect 18012 25304 18018 25316
rect 18785 25313 18797 25316
rect 18831 25313 18843 25347
rect 18785 25307 18843 25313
rect 21266 25304 21272 25356
rect 21324 25344 21330 25356
rect 21744 25353 21772 25452
rect 22278 25440 22284 25452
rect 22336 25440 22342 25492
rect 35434 25480 35440 25492
rect 25700 25452 35440 25480
rect 22738 25412 22744 25424
rect 22204 25384 22744 25412
rect 21729 25347 21787 25353
rect 21729 25344 21741 25347
rect 21324 25316 21741 25344
rect 21324 25304 21330 25316
rect 21729 25313 21741 25316
rect 21775 25313 21787 25347
rect 22002 25344 22008 25356
rect 21963 25316 22008 25344
rect 21729 25307 21787 25313
rect 22002 25304 22008 25316
rect 22060 25304 22066 25356
rect 10612 25248 11928 25276
rect 12897 25279 12955 25285
rect 4764 25180 6500 25208
rect 7392 25180 8892 25208
rect 4764 25168 4770 25180
rect 2961 25143 3019 25149
rect 2961 25109 2973 25143
rect 3007 25140 3019 25143
rect 3142 25140 3148 25152
rect 3007 25112 3148 25140
rect 3007 25109 3019 25112
rect 2961 25103 3019 25109
rect 3142 25100 3148 25112
rect 3200 25100 3206 25152
rect 6822 25100 6828 25152
rect 6880 25140 6886 25152
rect 7392 25140 7420 25180
rect 6880 25112 7420 25140
rect 6880 25100 6886 25112
rect 8570 25100 8576 25152
rect 8628 25140 8634 25152
rect 8757 25143 8815 25149
rect 8757 25140 8769 25143
rect 8628 25112 8769 25140
rect 8628 25100 8634 25112
rect 8757 25109 8769 25112
rect 8803 25109 8815 25143
rect 8864 25140 8892 25180
rect 10612 25140 10640 25248
rect 12897 25245 12909 25279
rect 12943 25276 12955 25279
rect 18509 25279 18567 25285
rect 12943 25248 16804 25276
rect 12943 25245 12955 25248
rect 12897 25239 12955 25245
rect 16666 25208 16672 25220
rect 16627 25180 16672 25208
rect 16666 25168 16672 25180
rect 16724 25168 16730 25220
rect 16776 25208 16804 25248
rect 18509 25245 18521 25279
rect 18555 25276 18567 25279
rect 19426 25276 19432 25288
rect 18555 25248 19432 25276
rect 18555 25245 18567 25248
rect 18509 25239 18567 25245
rect 19426 25236 19432 25248
rect 19484 25236 19490 25288
rect 19886 25276 19892 25288
rect 19847 25248 19892 25276
rect 19886 25236 19892 25248
rect 19944 25236 19950 25288
rect 22097 25279 22155 25285
rect 22097 25245 22109 25279
rect 22143 25276 22155 25279
rect 22204 25276 22232 25384
rect 22738 25372 22744 25384
rect 22796 25372 22802 25424
rect 24762 25412 24768 25424
rect 23860 25384 24768 25412
rect 22281 25347 22339 25353
rect 22281 25313 22293 25347
rect 22327 25313 22339 25347
rect 22281 25307 22339 25313
rect 22925 25347 22983 25353
rect 22925 25313 22937 25347
rect 22971 25313 22983 25347
rect 23106 25344 23112 25356
rect 23067 25316 23112 25344
rect 22925 25307 22983 25313
rect 22143 25248 22232 25276
rect 22143 25245 22155 25248
rect 22097 25239 22155 25245
rect 17957 25211 18015 25217
rect 17957 25208 17969 25211
rect 16776 25180 17969 25208
rect 17957 25177 17969 25180
rect 18003 25177 18015 25211
rect 17957 25171 18015 25177
rect 21818 25168 21824 25220
rect 21876 25208 21882 25220
rect 22296 25208 22324 25307
rect 22940 25276 22968 25307
rect 23106 25304 23112 25316
rect 23164 25304 23170 25356
rect 23658 25276 23664 25288
rect 22940 25248 23664 25276
rect 23658 25236 23664 25248
rect 23716 25236 23722 25288
rect 21876 25180 22324 25208
rect 21876 25168 21882 25180
rect 8864 25112 10640 25140
rect 8757 25103 8815 25109
rect 11054 25100 11060 25152
rect 11112 25140 11118 25152
rect 11241 25143 11299 25149
rect 11241 25140 11253 25143
rect 11112 25112 11253 25140
rect 11112 25100 11118 25112
rect 11241 25109 11253 25112
rect 11287 25140 11299 25143
rect 11606 25140 11612 25152
rect 11287 25112 11612 25140
rect 11287 25109 11299 25112
rect 11241 25103 11299 25109
rect 11606 25100 11612 25112
rect 11664 25100 11670 25152
rect 11974 25140 11980 25152
rect 11935 25112 11980 25140
rect 11974 25100 11980 25112
rect 12032 25100 12038 25152
rect 13538 25100 13544 25152
rect 13596 25140 13602 25152
rect 14185 25143 14243 25149
rect 14185 25140 14197 25143
rect 13596 25112 14197 25140
rect 13596 25100 13602 25112
rect 14185 25109 14197 25112
rect 14231 25140 14243 25143
rect 14918 25140 14924 25152
rect 14231 25112 14924 25140
rect 14231 25109 14243 25112
rect 14185 25103 14243 25109
rect 14918 25100 14924 25112
rect 14976 25100 14982 25152
rect 15562 25100 15568 25152
rect 15620 25140 15626 25152
rect 16850 25140 16856 25152
rect 15620 25112 16856 25140
rect 15620 25100 15626 25112
rect 16850 25100 16856 25112
rect 16908 25140 16914 25152
rect 17586 25140 17592 25152
rect 16908 25112 17592 25140
rect 16908 25100 16914 25112
rect 17586 25100 17592 25112
rect 17644 25100 17650 25152
rect 21634 25100 21640 25152
rect 21692 25140 21698 25152
rect 22002 25140 22008 25152
rect 21692 25112 22008 25140
rect 21692 25100 21698 25112
rect 22002 25100 22008 25112
rect 22060 25140 22066 25152
rect 23860 25140 23888 25384
rect 24762 25372 24768 25384
rect 24820 25372 24826 25424
rect 24026 25344 24032 25356
rect 23987 25316 24032 25344
rect 24026 25304 24032 25316
rect 24084 25304 24090 25356
rect 24176 25347 24234 25353
rect 24176 25313 24188 25347
rect 24222 25344 24234 25347
rect 24486 25344 24492 25356
rect 24222 25316 24492 25344
rect 24222 25313 24234 25316
rect 24176 25307 24234 25313
rect 24486 25304 24492 25316
rect 24544 25304 24550 25356
rect 25501 25347 25559 25353
rect 25501 25313 25513 25347
rect 25547 25344 25559 25347
rect 25700 25344 25728 25452
rect 35434 25440 35440 25452
rect 35492 25440 35498 25492
rect 35618 25440 35624 25492
rect 35676 25480 35682 25492
rect 35676 25452 37780 25480
rect 35676 25440 35682 25452
rect 26418 25372 26424 25424
rect 26476 25412 26482 25424
rect 26476 25384 27108 25412
rect 26476 25372 26482 25384
rect 25547 25316 25728 25344
rect 25961 25347 26019 25353
rect 25547 25313 25559 25316
rect 25501 25307 25559 25313
rect 25961 25313 25973 25347
rect 26007 25344 26019 25347
rect 26142 25344 26148 25356
rect 26007 25316 26148 25344
rect 26007 25313 26019 25316
rect 25961 25307 26019 25313
rect 26142 25304 26148 25316
rect 26200 25304 26206 25356
rect 27080 25353 27108 25384
rect 29914 25372 29920 25424
rect 29972 25412 29978 25424
rect 29972 25384 32168 25412
rect 29972 25372 29978 25384
rect 26513 25347 26571 25353
rect 26513 25313 26525 25347
rect 26559 25313 26571 25347
rect 26513 25307 26571 25313
rect 27065 25347 27123 25353
rect 27065 25313 27077 25347
rect 27111 25313 27123 25347
rect 28166 25344 28172 25356
rect 28127 25316 28172 25344
rect 27065 25307 27123 25313
rect 24397 25279 24455 25285
rect 24397 25245 24409 25279
rect 24443 25245 24455 25279
rect 24397 25239 24455 25245
rect 24765 25279 24823 25285
rect 24765 25245 24777 25279
rect 24811 25276 24823 25279
rect 26528 25276 26556 25307
rect 28166 25304 28172 25316
rect 28224 25304 28230 25356
rect 30558 25344 30564 25356
rect 30519 25316 30564 25344
rect 30558 25304 30564 25316
rect 30616 25304 30622 25356
rect 30742 25344 30748 25356
rect 30703 25316 30748 25344
rect 30742 25304 30748 25316
rect 30800 25304 30806 25356
rect 32140 25353 32168 25384
rect 30929 25347 30987 25353
rect 30929 25313 30941 25347
rect 30975 25313 30987 25347
rect 30929 25307 30987 25313
rect 32125 25347 32183 25353
rect 32125 25313 32137 25347
rect 32171 25313 32183 25347
rect 32766 25344 32772 25356
rect 32727 25316 32772 25344
rect 32125 25307 32183 25313
rect 24811 25248 26556 25276
rect 26881 25279 26939 25285
rect 24811 25245 24823 25248
rect 24765 25239 24823 25245
rect 26881 25245 26893 25279
rect 26927 25276 26939 25279
rect 27614 25276 27620 25288
rect 26927 25248 27620 25276
rect 26927 25245 26939 25248
rect 26881 25239 26939 25245
rect 24302 25208 24308 25220
rect 24263 25180 24308 25208
rect 24302 25168 24308 25180
rect 24360 25168 24366 25220
rect 24412 25208 24440 25239
rect 27614 25236 27620 25248
rect 27672 25236 27678 25288
rect 27893 25279 27951 25285
rect 27893 25245 27905 25279
rect 27939 25245 27951 25279
rect 27893 25239 27951 25245
rect 29549 25279 29607 25285
rect 29549 25245 29561 25279
rect 29595 25276 29607 25279
rect 29822 25276 29828 25288
rect 29595 25248 29828 25276
rect 29595 25245 29607 25248
rect 29549 25239 29607 25245
rect 24486 25208 24492 25220
rect 24412 25180 24492 25208
rect 24486 25168 24492 25180
rect 24544 25168 24550 25220
rect 26510 25168 26516 25220
rect 26568 25208 26574 25220
rect 27430 25208 27436 25220
rect 26568 25180 27436 25208
rect 26568 25168 26574 25180
rect 27430 25168 27436 25180
rect 27488 25208 27494 25220
rect 27908 25208 27936 25239
rect 29822 25236 29828 25248
rect 29880 25276 29886 25288
rect 30944 25276 30972 25307
rect 32766 25304 32772 25316
rect 32824 25304 32830 25356
rect 33962 25304 33968 25356
rect 34020 25344 34026 25356
rect 37366 25344 37372 25356
rect 34020 25316 37372 25344
rect 34020 25304 34026 25316
rect 37366 25304 37372 25316
rect 37424 25304 37430 25356
rect 37752 25353 37780 25452
rect 37737 25347 37795 25353
rect 37737 25313 37749 25347
rect 37783 25313 37795 25347
rect 37737 25307 37795 25313
rect 29880 25248 30972 25276
rect 29880 25236 29886 25248
rect 31202 25236 31208 25288
rect 31260 25276 31266 25288
rect 32784 25276 32812 25304
rect 31260 25248 32812 25276
rect 31260 25236 31266 25248
rect 32950 25236 32956 25288
rect 33008 25276 33014 25288
rect 33045 25279 33103 25285
rect 33045 25276 33057 25279
rect 33008 25248 33057 25276
rect 33008 25236 33014 25248
rect 33045 25245 33057 25248
rect 33091 25245 33103 25279
rect 33045 25239 33103 25245
rect 34330 25236 34336 25288
rect 34388 25276 34394 25288
rect 35345 25279 35403 25285
rect 35345 25276 35357 25279
rect 34388 25248 35357 25276
rect 34388 25236 34394 25248
rect 35345 25245 35357 25248
rect 35391 25245 35403 25279
rect 35345 25239 35403 25245
rect 35621 25279 35679 25285
rect 35621 25245 35633 25279
rect 35667 25276 35679 25279
rect 35710 25276 35716 25288
rect 35667 25248 35716 25276
rect 35667 25245 35679 25248
rect 35621 25239 35679 25245
rect 35710 25236 35716 25248
rect 35768 25236 35774 25288
rect 37921 25211 37979 25217
rect 37921 25208 37933 25211
rect 27488 25180 27936 25208
rect 36280 25180 37933 25208
rect 27488 25168 27494 25180
rect 22060 25112 23888 25140
rect 25317 25143 25375 25149
rect 22060 25100 22066 25112
rect 25317 25109 25329 25143
rect 25363 25140 25375 25143
rect 25406 25140 25412 25152
rect 25363 25112 25412 25140
rect 25363 25109 25375 25112
rect 25317 25103 25375 25109
rect 25406 25100 25412 25112
rect 25464 25100 25470 25152
rect 31938 25100 31944 25152
rect 31996 25140 32002 25152
rect 32217 25143 32275 25149
rect 32217 25140 32229 25143
rect 31996 25112 32229 25140
rect 31996 25100 32002 25112
rect 32217 25109 32229 25112
rect 32263 25109 32275 25143
rect 32217 25103 32275 25109
rect 33778 25100 33784 25152
rect 33836 25140 33842 25152
rect 34149 25143 34207 25149
rect 34149 25140 34161 25143
rect 33836 25112 34161 25140
rect 33836 25100 33842 25112
rect 34149 25109 34161 25112
rect 34195 25109 34207 25143
rect 34149 25103 34207 25109
rect 35526 25100 35532 25152
rect 35584 25140 35590 25152
rect 36280 25140 36308 25180
rect 37921 25177 37933 25180
rect 37967 25177 37979 25211
rect 37921 25171 37979 25177
rect 35584 25112 36308 25140
rect 35584 25100 35590 25112
rect 36538 25100 36544 25152
rect 36596 25140 36602 25152
rect 36725 25143 36783 25149
rect 36725 25140 36737 25143
rect 36596 25112 36737 25140
rect 36596 25100 36602 25112
rect 36725 25109 36737 25112
rect 36771 25109 36783 25143
rect 36725 25103 36783 25109
rect 1104 25050 38824 25072
rect 1104 24998 4246 25050
rect 4298 24998 4310 25050
rect 4362 24998 4374 25050
rect 4426 24998 4438 25050
rect 4490 24998 34966 25050
rect 35018 24998 35030 25050
rect 35082 24998 35094 25050
rect 35146 24998 35158 25050
rect 35210 24998 38824 25050
rect 1104 24976 38824 24998
rect 9766 24896 9772 24948
rect 9824 24936 9830 24948
rect 12618 24936 12624 24948
rect 9824 24908 12624 24936
rect 9824 24896 9830 24908
rect 12618 24896 12624 24908
rect 12676 24896 12682 24948
rect 16316 24908 16528 24936
rect 8662 24828 8668 24880
rect 8720 24868 8726 24880
rect 11974 24868 11980 24880
rect 8720 24840 11980 24868
rect 8720 24828 8726 24840
rect 2317 24803 2375 24809
rect 2317 24769 2329 24803
rect 2363 24800 2375 24803
rect 3053 24803 3111 24809
rect 3053 24800 3065 24803
rect 2363 24772 3065 24800
rect 2363 24769 2375 24772
rect 2317 24763 2375 24769
rect 3053 24769 3065 24772
rect 3099 24769 3111 24803
rect 3053 24763 3111 24769
rect 3234 24760 3240 24812
rect 3292 24760 3298 24812
rect 4062 24760 4068 24812
rect 4120 24800 4126 24812
rect 4157 24803 4215 24809
rect 4157 24800 4169 24803
rect 4120 24772 4169 24800
rect 4120 24760 4126 24772
rect 4157 24769 4169 24772
rect 4203 24769 4215 24803
rect 5534 24800 5540 24812
rect 5495 24772 5540 24800
rect 4157 24763 4215 24769
rect 5534 24760 5540 24772
rect 5592 24760 5598 24812
rect 7190 24800 7196 24812
rect 7151 24772 7196 24800
rect 7190 24760 7196 24772
rect 7248 24760 7254 24812
rect 7742 24800 7748 24812
rect 7703 24772 7748 24800
rect 7742 24760 7748 24772
rect 7800 24760 7806 24812
rect 8205 24803 8263 24809
rect 8205 24769 8217 24803
rect 8251 24800 8263 24803
rect 8386 24800 8392 24812
rect 8251 24772 8392 24800
rect 8251 24769 8263 24772
rect 8205 24763 8263 24769
rect 8386 24760 8392 24772
rect 8444 24800 8450 24812
rect 10796 24800 10824 24840
rect 11974 24828 11980 24840
rect 12032 24828 12038 24880
rect 8444 24772 10640 24800
rect 10796 24772 10916 24800
rect 8444 24760 8450 24772
rect 1854 24732 1860 24744
rect 1815 24704 1860 24732
rect 1854 24692 1860 24704
rect 1912 24692 1918 24744
rect 2133 24735 2191 24741
rect 2133 24701 2145 24735
rect 2179 24701 2191 24735
rect 2133 24695 2191 24701
rect 2148 24664 2176 24695
rect 2682 24692 2688 24744
rect 2740 24732 2746 24744
rect 2777 24735 2835 24741
rect 2777 24732 2789 24735
rect 2740 24704 2789 24732
rect 2740 24692 2746 24704
rect 2777 24701 2789 24704
rect 2823 24701 2835 24735
rect 3252 24732 3280 24760
rect 2777 24695 2835 24701
rect 2884 24704 3280 24732
rect 5261 24735 5319 24741
rect 2884 24664 2912 24704
rect 5261 24701 5273 24735
rect 5307 24701 5319 24735
rect 5261 24695 5319 24701
rect 5353 24735 5411 24741
rect 5353 24701 5365 24735
rect 5399 24701 5411 24735
rect 5353 24695 5411 24701
rect 2148 24636 2912 24664
rect 5276 24596 5304 24695
rect 5368 24664 5396 24695
rect 5442 24692 5448 24744
rect 5500 24732 5506 24744
rect 5721 24735 5779 24741
rect 5721 24732 5733 24735
rect 5500 24704 5733 24732
rect 5500 24692 5506 24704
rect 5721 24701 5733 24704
rect 5767 24701 5779 24735
rect 5721 24695 5779 24701
rect 6914 24692 6920 24744
rect 6972 24732 6978 24744
rect 8021 24735 8079 24741
rect 8021 24732 8033 24735
rect 6972 24704 8033 24732
rect 6972 24692 6978 24704
rect 8021 24701 8033 24704
rect 8067 24701 8079 24735
rect 9214 24732 9220 24744
rect 9175 24704 9220 24732
rect 8021 24695 8079 24701
rect 9214 24692 9220 24704
rect 9272 24692 9278 24744
rect 9861 24735 9919 24741
rect 9861 24701 9873 24735
rect 9907 24701 9919 24735
rect 9861 24695 9919 24701
rect 7098 24664 7104 24676
rect 5368 24636 7104 24664
rect 7098 24624 7104 24636
rect 7156 24624 7162 24676
rect 9490 24624 9496 24676
rect 9548 24664 9554 24676
rect 9585 24667 9643 24673
rect 9585 24664 9597 24667
rect 9548 24636 9597 24664
rect 9548 24624 9554 24636
rect 9585 24633 9597 24636
rect 9631 24633 9643 24667
rect 9585 24627 9643 24633
rect 6822 24596 6828 24608
rect 5276 24568 6828 24596
rect 6822 24556 6828 24568
rect 6880 24556 6886 24608
rect 9876 24596 9904 24695
rect 10042 24692 10048 24744
rect 10100 24732 10106 24744
rect 10612 24741 10640 24772
rect 10137 24735 10195 24741
rect 10137 24732 10149 24735
rect 10100 24704 10149 24732
rect 10100 24692 10106 24704
rect 10137 24701 10149 24704
rect 10183 24701 10195 24735
rect 10137 24695 10195 24701
rect 10597 24735 10655 24741
rect 10597 24701 10609 24735
rect 10643 24732 10655 24735
rect 10778 24732 10784 24744
rect 10643 24704 10784 24732
rect 10643 24701 10655 24704
rect 10597 24695 10655 24701
rect 10778 24692 10784 24704
rect 10836 24692 10842 24744
rect 10888 24741 10916 24772
rect 12434 24760 12440 24812
rect 12492 24800 12498 24812
rect 13449 24803 13507 24809
rect 12492 24772 12537 24800
rect 12492 24760 12498 24772
rect 13449 24769 13461 24803
rect 13495 24800 13507 24803
rect 13538 24800 13544 24812
rect 13495 24772 13544 24800
rect 13495 24769 13507 24772
rect 13449 24763 13507 24769
rect 13538 24760 13544 24772
rect 13596 24760 13602 24812
rect 13909 24803 13967 24809
rect 13909 24769 13921 24803
rect 13955 24800 13967 24803
rect 16316 24800 16344 24908
rect 13955 24772 16344 24800
rect 16500 24800 16528 24908
rect 19426 24896 19432 24948
rect 19484 24936 19490 24948
rect 22278 24936 22284 24948
rect 19484 24908 22284 24936
rect 19484 24896 19490 24908
rect 22278 24896 22284 24908
rect 22336 24896 22342 24948
rect 25038 24896 25044 24948
rect 25096 24936 25102 24948
rect 27798 24936 27804 24948
rect 25096 24908 27804 24936
rect 25096 24896 25102 24908
rect 27798 24896 27804 24908
rect 27856 24896 27862 24948
rect 36262 24896 36268 24948
rect 36320 24936 36326 24948
rect 36449 24939 36507 24945
rect 36449 24936 36461 24939
rect 36320 24908 36461 24936
rect 36320 24896 36326 24908
rect 36449 24905 36461 24908
rect 36495 24936 36507 24939
rect 38010 24936 38016 24948
rect 36495 24908 38016 24936
rect 36495 24905 36507 24908
rect 36449 24899 36507 24905
rect 38010 24896 38016 24908
rect 38068 24896 38074 24948
rect 18046 24828 18052 24880
rect 18104 24868 18110 24880
rect 18966 24868 18972 24880
rect 18104 24840 18972 24868
rect 18104 24828 18110 24840
rect 18966 24828 18972 24840
rect 19024 24828 19030 24880
rect 20070 24868 20076 24880
rect 20031 24840 20076 24868
rect 20070 24828 20076 24840
rect 20128 24828 20134 24880
rect 23658 24868 23664 24880
rect 22480 24840 23664 24868
rect 17221 24803 17279 24809
rect 17221 24800 17233 24803
rect 16500 24772 17233 24800
rect 13955 24769 13967 24772
rect 13909 24763 13967 24769
rect 17221 24769 17233 24772
rect 17267 24769 17279 24803
rect 21082 24800 21088 24812
rect 17221 24763 17279 24769
rect 17420 24772 20024 24800
rect 21043 24772 21088 24800
rect 10873 24735 10931 24741
rect 10873 24701 10885 24735
rect 10919 24701 10931 24735
rect 11606 24732 11612 24744
rect 11567 24704 11612 24732
rect 10873 24695 10931 24701
rect 11606 24692 11612 24704
rect 11664 24692 11670 24744
rect 12066 24692 12072 24744
rect 12124 24732 12130 24744
rect 12989 24735 13047 24741
rect 12989 24732 13001 24735
rect 12124 24704 13001 24732
rect 12124 24692 12130 24704
rect 12989 24701 13001 24704
rect 13035 24701 13047 24735
rect 12989 24695 13047 24701
rect 13265 24735 13323 24741
rect 13265 24701 13277 24735
rect 13311 24701 13323 24735
rect 13265 24695 13323 24701
rect 10686 24624 10692 24676
rect 10744 24664 10750 24676
rect 13280 24664 13308 24695
rect 14274 24692 14280 24744
rect 14332 24732 14338 24744
rect 14461 24735 14519 24741
rect 14461 24732 14473 24735
rect 14332 24704 14473 24732
rect 14332 24692 14338 24704
rect 14461 24701 14473 24704
rect 14507 24732 14519 24735
rect 14642 24732 14648 24744
rect 14507 24704 14648 24732
rect 14507 24701 14519 24704
rect 14461 24695 14519 24701
rect 14642 24692 14648 24704
rect 14700 24692 14706 24744
rect 14737 24735 14795 24741
rect 14737 24701 14749 24735
rect 14783 24701 14795 24735
rect 14918 24732 14924 24744
rect 14879 24704 14924 24732
rect 14737 24695 14795 24701
rect 10744 24636 13308 24664
rect 14752 24664 14780 24695
rect 14918 24692 14924 24704
rect 14976 24692 14982 24744
rect 15654 24732 15660 24744
rect 15615 24704 15660 24732
rect 15654 24692 15660 24704
rect 15712 24692 15718 24744
rect 16485 24735 16543 24741
rect 16485 24701 16497 24735
rect 16531 24732 16543 24735
rect 16666 24732 16672 24744
rect 16531 24704 16672 24732
rect 16531 24701 16543 24704
rect 16485 24695 16543 24701
rect 16666 24692 16672 24704
rect 16724 24692 16730 24744
rect 17126 24732 17132 24744
rect 17087 24704 17132 24732
rect 17126 24692 17132 24704
rect 17184 24692 17190 24744
rect 14752 24636 14964 24664
rect 10744 24624 10750 24636
rect 14936 24608 14964 24636
rect 16206 24624 16212 24676
rect 16264 24664 16270 24676
rect 17420 24664 17448 24772
rect 18601 24735 18659 24741
rect 18601 24701 18613 24735
rect 18647 24701 18659 24735
rect 18782 24732 18788 24744
rect 18743 24704 18788 24732
rect 18601 24695 18659 24701
rect 18138 24664 18144 24676
rect 16264 24636 17448 24664
rect 18099 24636 18144 24664
rect 16264 24624 16270 24636
rect 18138 24624 18144 24636
rect 18196 24624 18202 24676
rect 18616 24664 18644 24695
rect 18782 24692 18788 24704
rect 18840 24692 18846 24744
rect 18966 24732 18972 24744
rect 18927 24704 18972 24732
rect 18966 24692 18972 24704
rect 19024 24692 19030 24744
rect 19886 24732 19892 24744
rect 19847 24704 19892 24732
rect 19886 24692 19892 24704
rect 19944 24692 19950 24744
rect 19996 24732 20024 24772
rect 21082 24760 21088 24772
rect 21140 24760 21146 24812
rect 21192 24772 22416 24800
rect 21192 24732 21220 24772
rect 19996 24704 21220 24732
rect 21266 24692 21272 24744
rect 21324 24732 21330 24744
rect 21634 24732 21640 24744
rect 21324 24704 21369 24732
rect 21595 24704 21640 24732
rect 21324 24692 21330 24704
rect 21634 24692 21640 24704
rect 21692 24692 21698 24744
rect 21818 24732 21824 24744
rect 21779 24704 21824 24732
rect 21818 24692 21824 24704
rect 21876 24692 21882 24744
rect 19334 24664 19340 24676
rect 18616 24636 19340 24664
rect 19334 24624 19340 24636
rect 19392 24624 19398 24676
rect 22388 24664 22416 24772
rect 22480 24741 22508 24840
rect 23658 24828 23664 24840
rect 23716 24828 23722 24880
rect 25501 24871 25559 24877
rect 25501 24837 25513 24871
rect 25547 24868 25559 24871
rect 25590 24868 25596 24880
rect 25547 24840 25596 24868
rect 25547 24837 25559 24840
rect 25501 24831 25559 24837
rect 25590 24828 25596 24840
rect 25648 24828 25654 24880
rect 28169 24871 28227 24877
rect 28169 24837 28181 24871
rect 28215 24868 28227 24871
rect 29086 24868 29092 24880
rect 28215 24840 29092 24868
rect 28215 24837 28227 24840
rect 28169 24831 28227 24837
rect 29086 24828 29092 24840
rect 29144 24828 29150 24880
rect 22738 24760 22744 24812
rect 22796 24800 22802 24812
rect 24673 24803 24731 24809
rect 24673 24800 24685 24803
rect 22796 24772 24685 24800
rect 22796 24760 22802 24772
rect 24673 24769 24685 24772
rect 24719 24769 24731 24803
rect 24673 24763 24731 24769
rect 27433 24803 27491 24809
rect 27433 24769 27445 24803
rect 27479 24800 27491 24803
rect 28258 24800 28264 24812
rect 27479 24772 28264 24800
rect 27479 24769 27491 24772
rect 27433 24763 27491 24769
rect 28258 24760 28264 24772
rect 28316 24760 28322 24812
rect 31938 24760 31944 24812
rect 31996 24800 32002 24812
rect 32125 24803 32183 24809
rect 32125 24800 32137 24803
rect 31996 24772 32137 24800
rect 31996 24760 32002 24772
rect 32125 24769 32137 24772
rect 32171 24769 32183 24803
rect 33962 24800 33968 24812
rect 32125 24763 32183 24769
rect 33888 24772 33968 24800
rect 22465 24735 22523 24741
rect 22465 24701 22477 24735
rect 22511 24701 22523 24735
rect 22646 24732 22652 24744
rect 22607 24704 22652 24732
rect 22465 24695 22523 24701
rect 22646 24692 22652 24704
rect 22704 24692 22710 24744
rect 23658 24732 23664 24744
rect 23571 24704 23664 24732
rect 23658 24692 23664 24704
rect 23716 24732 23722 24744
rect 24210 24732 24216 24744
rect 23716 24704 24216 24732
rect 23716 24692 23722 24704
rect 24210 24692 24216 24704
rect 24268 24692 24274 24744
rect 24946 24732 24952 24744
rect 24907 24704 24952 24732
rect 24946 24692 24952 24704
rect 25004 24692 25010 24744
rect 25406 24732 25412 24744
rect 25367 24704 25412 24732
rect 25406 24692 25412 24704
rect 25464 24692 25470 24744
rect 26142 24732 26148 24744
rect 26103 24704 26148 24732
rect 26142 24692 26148 24704
rect 26200 24692 26206 24744
rect 27706 24732 27712 24744
rect 27667 24704 27712 24732
rect 27706 24692 27712 24704
rect 27764 24692 27770 24744
rect 28074 24732 28080 24744
rect 28035 24704 28080 24732
rect 28074 24692 28080 24704
rect 28132 24692 28138 24744
rect 29270 24732 29276 24744
rect 29231 24704 29276 24732
rect 29270 24692 29276 24704
rect 29328 24692 29334 24744
rect 29822 24732 29828 24744
rect 29783 24704 29828 24732
rect 29822 24692 29828 24704
rect 29880 24692 29886 24744
rect 30466 24732 30472 24744
rect 30427 24704 30472 24732
rect 30466 24692 30472 24704
rect 30524 24692 30530 24744
rect 31386 24732 31392 24744
rect 31347 24704 31392 24732
rect 31386 24692 31392 24704
rect 31444 24692 31450 24744
rect 32030 24732 32036 24744
rect 31991 24704 32036 24732
rect 32030 24692 32036 24704
rect 32088 24692 32094 24744
rect 32861 24735 32919 24741
rect 32861 24701 32873 24735
rect 32907 24732 32919 24735
rect 33042 24732 33048 24744
rect 32907 24704 33048 24732
rect 32907 24701 32919 24704
rect 32861 24695 32919 24701
rect 33042 24692 33048 24704
rect 33100 24692 33106 24744
rect 33888 24741 33916 24772
rect 33962 24760 33968 24772
rect 34020 24760 34026 24812
rect 34333 24803 34391 24809
rect 34333 24769 34345 24803
rect 34379 24800 34391 24803
rect 34514 24800 34520 24812
rect 34379 24772 34520 24800
rect 34379 24769 34391 24772
rect 34333 24763 34391 24769
rect 34514 24760 34520 24772
rect 34572 24760 34578 24812
rect 34606 24760 34612 24812
rect 34664 24800 34670 24812
rect 35161 24803 35219 24809
rect 35161 24800 35173 24803
rect 34664 24772 35173 24800
rect 34664 24760 34670 24772
rect 35161 24769 35173 24772
rect 35207 24769 35219 24803
rect 35161 24763 35219 24769
rect 33873 24735 33931 24741
rect 33873 24701 33885 24735
rect 33919 24701 33931 24735
rect 33873 24695 33931 24701
rect 34885 24735 34943 24741
rect 34885 24701 34897 24735
rect 34931 24732 34943 24735
rect 36078 24732 36084 24744
rect 34931 24704 36084 24732
rect 34931 24701 34943 24704
rect 34885 24695 34943 24701
rect 32582 24664 32588 24676
rect 19996 24636 20300 24664
rect 22388 24636 32588 24664
rect 11698 24596 11704 24608
rect 9876 24568 11704 24596
rect 11698 24556 11704 24568
rect 11756 24596 11762 24608
rect 11793 24599 11851 24605
rect 11793 24596 11805 24599
rect 11756 24568 11805 24596
rect 11756 24556 11762 24568
rect 11793 24565 11805 24568
rect 11839 24565 11851 24599
rect 11793 24559 11851 24565
rect 14918 24556 14924 24608
rect 14976 24556 14982 24608
rect 15562 24556 15568 24608
rect 15620 24596 15626 24608
rect 15841 24599 15899 24605
rect 15841 24596 15853 24599
rect 15620 24568 15853 24596
rect 15620 24556 15626 24568
rect 15841 24565 15853 24568
rect 15887 24565 15899 24599
rect 15841 24559 15899 24565
rect 16485 24599 16543 24605
rect 16485 24565 16497 24599
rect 16531 24596 16543 24599
rect 19996 24596 20024 24636
rect 16531 24568 20024 24596
rect 20272 24596 20300 24636
rect 32582 24624 32588 24636
rect 32640 24624 32646 24676
rect 33594 24664 33600 24676
rect 33555 24636 33600 24664
rect 33594 24624 33600 24636
rect 33652 24624 33658 24676
rect 33962 24624 33968 24676
rect 34020 24664 34026 24676
rect 34020 24636 34065 24664
rect 34020 24624 34026 24636
rect 34330 24624 34336 24676
rect 34388 24664 34394 24676
rect 34900 24664 34928 24695
rect 36078 24692 36084 24704
rect 36136 24732 36142 24744
rect 36354 24732 36360 24744
rect 36136 24704 36360 24732
rect 36136 24692 36142 24704
rect 36354 24692 36360 24704
rect 36412 24692 36418 24744
rect 37182 24732 37188 24744
rect 37143 24704 37188 24732
rect 37182 24692 37188 24704
rect 37240 24692 37246 24744
rect 37553 24735 37611 24741
rect 37553 24701 37565 24735
rect 37599 24732 37611 24735
rect 37826 24732 37832 24744
rect 37599 24704 37832 24732
rect 37599 24701 37611 24704
rect 37553 24695 37611 24701
rect 37826 24692 37832 24704
rect 37884 24692 37890 24744
rect 34388 24636 34928 24664
rect 37737 24667 37795 24673
rect 34388 24624 34394 24636
rect 37737 24633 37749 24667
rect 37783 24664 37795 24667
rect 38010 24664 38016 24676
rect 37783 24636 38016 24664
rect 37783 24633 37795 24636
rect 37737 24627 37795 24633
rect 38010 24624 38016 24636
rect 38068 24624 38074 24676
rect 22462 24596 22468 24608
rect 20272 24568 22468 24596
rect 16531 24565 16543 24568
rect 16485 24559 16543 24565
rect 22462 24556 22468 24568
rect 22520 24556 22526 24608
rect 23566 24556 23572 24608
rect 23624 24596 23630 24608
rect 23845 24599 23903 24605
rect 23845 24596 23857 24599
rect 23624 24568 23857 24596
rect 23624 24556 23630 24568
rect 23845 24565 23857 24568
rect 23891 24596 23903 24599
rect 24394 24596 24400 24608
rect 23891 24568 24400 24596
rect 23891 24565 23903 24568
rect 23845 24559 23903 24565
rect 24394 24556 24400 24568
rect 24452 24556 24458 24608
rect 24670 24556 24676 24608
rect 24728 24596 24734 24608
rect 26329 24599 26387 24605
rect 26329 24596 26341 24599
rect 24728 24568 26341 24596
rect 24728 24556 24734 24568
rect 26329 24565 26341 24568
rect 26375 24565 26387 24599
rect 26329 24559 26387 24565
rect 28994 24556 29000 24608
rect 29052 24596 29058 24608
rect 29365 24599 29423 24605
rect 29365 24596 29377 24599
rect 29052 24568 29377 24596
rect 29052 24556 29058 24568
rect 29365 24565 29377 24568
rect 29411 24565 29423 24599
rect 29365 24559 29423 24565
rect 30561 24599 30619 24605
rect 30561 24565 30573 24599
rect 30607 24596 30619 24599
rect 30650 24596 30656 24608
rect 30607 24568 30656 24596
rect 30607 24565 30619 24568
rect 30561 24559 30619 24565
rect 30650 24556 30656 24568
rect 30708 24556 30714 24608
rect 31389 24599 31447 24605
rect 31389 24565 31401 24599
rect 31435 24596 31447 24599
rect 31478 24596 31484 24608
rect 31435 24568 31484 24596
rect 31435 24565 31447 24568
rect 31389 24559 31447 24565
rect 31478 24556 31484 24568
rect 31536 24556 31542 24608
rect 32306 24556 32312 24608
rect 32364 24596 32370 24608
rect 32858 24596 32864 24608
rect 32364 24568 32864 24596
rect 32364 24556 32370 24568
rect 32858 24556 32864 24568
rect 32916 24596 32922 24608
rect 33045 24599 33103 24605
rect 33045 24596 33057 24599
rect 32916 24568 33057 24596
rect 32916 24556 32922 24568
rect 33045 24565 33057 24568
rect 33091 24565 33103 24599
rect 33045 24559 33103 24565
rect 33781 24599 33839 24605
rect 33781 24565 33793 24599
rect 33827 24596 33839 24599
rect 36814 24596 36820 24608
rect 33827 24568 36820 24596
rect 33827 24565 33839 24568
rect 33781 24559 33839 24565
rect 36814 24556 36820 24568
rect 36872 24556 36878 24608
rect 1104 24506 38824 24528
rect 1104 24454 19606 24506
rect 19658 24454 19670 24506
rect 19722 24454 19734 24506
rect 19786 24454 19798 24506
rect 19850 24454 38824 24506
rect 1104 24432 38824 24454
rect 1765 24395 1823 24401
rect 1765 24361 1777 24395
rect 1811 24392 1823 24395
rect 16206 24392 16212 24404
rect 1811 24364 16212 24392
rect 1811 24361 1823 24364
rect 1765 24355 1823 24361
rect 16206 24352 16212 24364
rect 16264 24352 16270 24404
rect 16301 24395 16359 24401
rect 16301 24361 16313 24395
rect 16347 24392 16359 24395
rect 24946 24392 24952 24404
rect 16347 24364 21312 24392
rect 16347 24361 16359 24364
rect 16301 24355 16359 24361
rect 4890 24324 4896 24336
rect 2332 24296 4896 24324
rect 1673 24259 1731 24265
rect 1673 24225 1685 24259
rect 1719 24256 1731 24259
rect 1719 24228 2176 24256
rect 1719 24225 1731 24228
rect 1673 24219 1731 24225
rect 2148 24188 2176 24228
rect 2222 24216 2228 24268
rect 2280 24256 2286 24268
rect 2332 24265 2360 24296
rect 4890 24284 4896 24296
rect 4948 24284 4954 24336
rect 6917 24327 6975 24333
rect 6917 24293 6929 24327
rect 6963 24324 6975 24327
rect 7006 24324 7012 24336
rect 6963 24296 7012 24324
rect 6963 24293 6975 24296
rect 6917 24287 6975 24293
rect 7006 24284 7012 24296
rect 7064 24284 7070 24336
rect 8386 24284 8392 24336
rect 8444 24324 8450 24336
rect 8573 24327 8631 24333
rect 8573 24324 8585 24327
rect 8444 24296 8585 24324
rect 8444 24284 8450 24296
rect 8573 24293 8585 24296
rect 8619 24293 8631 24327
rect 8754 24324 8760 24336
rect 8715 24296 8760 24324
rect 8573 24287 8631 24293
rect 8754 24284 8760 24296
rect 8812 24284 8818 24336
rect 9677 24327 9735 24333
rect 9677 24293 9689 24327
rect 9723 24324 9735 24327
rect 11054 24324 11060 24336
rect 9723 24296 9812 24324
rect 9723 24293 9735 24296
rect 9677 24287 9735 24293
rect 2317 24259 2375 24265
rect 2317 24256 2329 24259
rect 2280 24228 2329 24256
rect 2280 24216 2286 24228
rect 2317 24225 2329 24228
rect 2363 24225 2375 24259
rect 2317 24219 2375 24225
rect 2866 24216 2872 24268
rect 2924 24256 2930 24268
rect 3053 24259 3111 24265
rect 3053 24256 3065 24259
rect 2924 24228 3065 24256
rect 2924 24216 2930 24228
rect 3053 24225 3065 24228
rect 3099 24256 3111 24259
rect 3234 24256 3240 24268
rect 3099 24228 3240 24256
rect 3099 24225 3111 24228
rect 3053 24219 3111 24225
rect 3234 24216 3240 24228
rect 3292 24216 3298 24268
rect 5077 24259 5135 24265
rect 5077 24225 5089 24259
rect 5123 24256 5135 24259
rect 5994 24256 6000 24268
rect 5123 24228 6000 24256
rect 5123 24225 5135 24228
rect 5077 24219 5135 24225
rect 5994 24216 6000 24228
rect 6052 24216 6058 24268
rect 6457 24259 6515 24265
rect 6457 24225 6469 24259
rect 6503 24256 6515 24259
rect 7098 24256 7104 24268
rect 6503 24228 7104 24256
rect 6503 24225 6515 24228
rect 6457 24219 6515 24225
rect 7098 24216 7104 24228
rect 7156 24256 7162 24268
rect 7742 24256 7748 24268
rect 7156 24228 7604 24256
rect 7703 24228 7748 24256
rect 7156 24216 7162 24228
rect 2774 24188 2780 24200
rect 2148 24160 2780 24188
rect 2774 24148 2780 24160
rect 2832 24148 2838 24200
rect 3142 24188 3148 24200
rect 3103 24160 3148 24188
rect 3142 24148 3148 24160
rect 3200 24148 3206 24200
rect 4706 24148 4712 24200
rect 4764 24188 4770 24200
rect 4801 24191 4859 24197
rect 4801 24188 4813 24191
rect 4764 24160 4813 24188
rect 4764 24148 4770 24160
rect 4801 24157 4813 24160
rect 4847 24157 4859 24191
rect 7466 24188 7472 24200
rect 7427 24160 7472 24188
rect 4801 24151 4859 24157
rect 7466 24148 7472 24160
rect 7524 24148 7530 24200
rect 7576 24188 7604 24228
rect 7742 24216 7748 24228
rect 7800 24216 7806 24268
rect 8662 24256 8668 24268
rect 8623 24228 8668 24256
rect 8662 24216 8668 24228
rect 8720 24216 8726 24268
rect 9122 24256 9128 24268
rect 9083 24228 9128 24256
rect 9122 24216 9128 24228
rect 9180 24216 9186 24268
rect 9490 24216 9496 24268
rect 9548 24256 9554 24268
rect 9784 24256 9812 24296
rect 10704 24296 11060 24324
rect 9950 24256 9956 24268
rect 9548 24228 9720 24256
rect 9784 24228 9956 24256
rect 9548 24216 9554 24228
rect 7929 24191 7987 24197
rect 7929 24188 7941 24191
rect 7576 24160 7941 24188
rect 7929 24157 7941 24160
rect 7975 24188 7987 24191
rect 8018 24188 8024 24200
rect 7975 24160 8024 24188
rect 7975 24157 7987 24160
rect 7929 24151 7987 24157
rect 8018 24148 8024 24160
rect 8076 24148 8082 24200
rect 8389 24191 8447 24197
rect 8389 24157 8401 24191
rect 8435 24188 8447 24191
rect 8846 24188 8852 24200
rect 8435 24160 8852 24188
rect 8435 24157 8447 24160
rect 8389 24151 8447 24157
rect 8846 24148 8852 24160
rect 8904 24188 8910 24200
rect 9582 24188 9588 24200
rect 8904 24160 9588 24188
rect 8904 24148 8910 24160
rect 9582 24148 9588 24160
rect 9640 24148 9646 24200
rect 9692 24188 9720 24228
rect 9950 24216 9956 24228
rect 10008 24216 10014 24268
rect 10229 24259 10287 24265
rect 10229 24256 10241 24259
rect 10060 24228 10241 24256
rect 10060 24188 10088 24228
rect 10229 24225 10241 24228
rect 10275 24225 10287 24259
rect 10502 24256 10508 24268
rect 10463 24228 10508 24256
rect 10229 24219 10287 24225
rect 10502 24216 10508 24228
rect 10560 24216 10566 24268
rect 10704 24265 10732 24296
rect 11054 24284 11060 24296
rect 11112 24324 11118 24336
rect 11698 24324 11704 24336
rect 11112 24296 11704 24324
rect 11112 24284 11118 24296
rect 11698 24284 11704 24296
rect 11756 24284 11762 24336
rect 14918 24324 14924 24336
rect 13832 24296 14924 24324
rect 10689 24259 10747 24265
rect 10689 24225 10701 24259
rect 10735 24225 10747 24259
rect 10689 24219 10747 24225
rect 12345 24259 12403 24265
rect 12345 24225 12357 24259
rect 12391 24256 12403 24259
rect 13170 24256 13176 24268
rect 12391 24228 13176 24256
rect 12391 24225 12403 24228
rect 12345 24219 12403 24225
rect 13170 24216 13176 24228
rect 13228 24216 13234 24268
rect 13262 24216 13268 24268
rect 13320 24256 13326 24268
rect 13832 24265 13860 24296
rect 14918 24284 14924 24296
rect 14976 24284 14982 24336
rect 16758 24284 16764 24336
rect 16816 24324 16822 24336
rect 16816 24296 18644 24324
rect 16816 24284 16822 24296
rect 13817 24259 13875 24265
rect 13320 24228 13365 24256
rect 13320 24216 13326 24228
rect 13817 24225 13829 24259
rect 13863 24225 13875 24259
rect 13817 24219 13875 24225
rect 14185 24259 14243 24265
rect 14185 24225 14197 24259
rect 14231 24256 14243 24259
rect 14642 24256 14648 24268
rect 14231 24228 14648 24256
rect 14231 24225 14243 24228
rect 14185 24219 14243 24225
rect 14642 24216 14648 24228
rect 14700 24216 14706 24268
rect 15102 24216 15108 24268
rect 15160 24256 15166 24268
rect 15289 24259 15347 24265
rect 15289 24256 15301 24259
rect 15160 24228 15301 24256
rect 15160 24216 15166 24228
rect 15289 24225 15301 24228
rect 15335 24225 15347 24259
rect 15289 24219 15347 24225
rect 16393 24259 16451 24265
rect 16393 24225 16405 24259
rect 16439 24256 16451 24259
rect 16482 24256 16488 24268
rect 16439 24228 16488 24256
rect 16439 24225 16451 24228
rect 16393 24219 16451 24225
rect 16482 24216 16488 24228
rect 16540 24216 16546 24268
rect 16942 24256 16948 24268
rect 16903 24228 16948 24256
rect 16942 24216 16948 24228
rect 17000 24216 17006 24268
rect 18138 24256 18144 24268
rect 18099 24228 18144 24256
rect 18138 24216 18144 24228
rect 18196 24216 18202 24268
rect 18616 24265 18644 24296
rect 19334 24284 19340 24336
rect 19392 24324 19398 24336
rect 19978 24324 19984 24336
rect 19392 24296 19984 24324
rect 19392 24284 19398 24296
rect 19978 24284 19984 24296
rect 20036 24284 20042 24336
rect 18601 24259 18659 24265
rect 18601 24225 18613 24259
rect 18647 24225 18659 24259
rect 18601 24219 18659 24225
rect 19426 24216 19432 24268
rect 19484 24256 19490 24268
rect 20073 24259 20131 24265
rect 20073 24256 20085 24259
rect 19484 24228 20085 24256
rect 19484 24216 19490 24228
rect 20073 24225 20085 24228
rect 20119 24256 20131 24259
rect 20898 24256 20904 24268
rect 20119 24228 20904 24256
rect 20119 24225 20131 24228
rect 20073 24219 20131 24225
rect 20898 24216 20904 24228
rect 20956 24216 20962 24268
rect 21082 24256 21088 24268
rect 21043 24228 21088 24256
rect 21082 24216 21088 24228
rect 21140 24216 21146 24268
rect 21284 24265 21312 24364
rect 21376 24364 24952 24392
rect 21269 24259 21327 24265
rect 21269 24225 21281 24259
rect 21315 24225 21327 24259
rect 21269 24219 21327 24225
rect 9692 24160 10088 24188
rect 11517 24191 11575 24197
rect 11517 24157 11529 24191
rect 11563 24188 11575 24191
rect 11698 24188 11704 24200
rect 11563 24160 11704 24188
rect 11563 24157 11575 24160
rect 11517 24151 11575 24157
rect 11698 24148 11704 24160
rect 11756 24148 11762 24200
rect 12066 24188 12072 24200
rect 11979 24160 12072 24188
rect 12066 24148 12072 24160
rect 12124 24148 12130 24200
rect 12158 24148 12164 24200
rect 12216 24197 12222 24200
rect 12216 24191 12265 24197
rect 12216 24157 12219 24191
rect 12253 24157 12265 24191
rect 17037 24191 17095 24197
rect 17037 24188 17049 24191
rect 12216 24151 12265 24157
rect 13464 24160 17049 24188
rect 12216 24148 12222 24151
rect 2406 24120 2412 24132
rect 2367 24092 2412 24120
rect 2406 24080 2412 24092
rect 2464 24080 2470 24132
rect 7484 24120 7512 24148
rect 12084 24120 12112 24148
rect 7484 24092 12112 24120
rect 12526 24080 12532 24132
rect 12584 24120 12590 24132
rect 13464 24120 13492 24160
rect 17037 24157 17049 24160
rect 17083 24157 17095 24191
rect 17037 24151 17095 24157
rect 17218 24148 17224 24200
rect 17276 24188 17282 24200
rect 18877 24191 18935 24197
rect 18877 24188 18889 24191
rect 17276 24160 18889 24188
rect 17276 24148 17282 24160
rect 18877 24157 18889 24160
rect 18923 24157 18935 24191
rect 18877 24151 18935 24157
rect 12584 24092 13492 24120
rect 12584 24080 12590 24092
rect 13814 24080 13820 24132
rect 13872 24120 13878 24132
rect 14093 24123 14151 24129
rect 14093 24120 14105 24123
rect 13872 24092 14105 24120
rect 13872 24080 13878 24092
rect 14093 24089 14105 24092
rect 14139 24089 14151 24123
rect 14093 24083 14151 24089
rect 18325 24123 18383 24129
rect 18325 24089 18337 24123
rect 18371 24120 18383 24123
rect 21376 24120 21404 24364
rect 24946 24352 24952 24364
rect 25004 24352 25010 24404
rect 27617 24395 27675 24401
rect 27617 24361 27629 24395
rect 27663 24392 27675 24395
rect 28074 24392 28080 24404
rect 27663 24364 28080 24392
rect 27663 24361 27675 24364
rect 27617 24355 27675 24361
rect 28074 24352 28080 24364
rect 28132 24352 28138 24404
rect 28718 24392 28724 24404
rect 28184 24364 28724 24392
rect 22005 24327 22063 24333
rect 22005 24293 22017 24327
rect 22051 24324 22063 24327
rect 25222 24324 25228 24336
rect 22051 24296 25228 24324
rect 22051 24293 22063 24296
rect 22005 24287 22063 24293
rect 25222 24284 25228 24296
rect 25280 24284 25286 24336
rect 28184 24324 28212 24364
rect 28718 24352 28724 24364
rect 28776 24392 28782 24404
rect 34698 24392 34704 24404
rect 28776 24364 34704 24392
rect 28776 24352 28782 24364
rect 34698 24352 34704 24364
rect 34756 24352 34762 24404
rect 37826 24392 37832 24404
rect 37787 24364 37832 24392
rect 37826 24352 37832 24364
rect 37884 24352 37890 24404
rect 34790 24324 34796 24336
rect 26528 24296 28212 24324
rect 34532 24296 34796 24324
rect 21726 24256 21732 24268
rect 21687 24228 21732 24256
rect 21726 24216 21732 24228
rect 21784 24216 21790 24268
rect 22646 24216 22652 24268
rect 22704 24256 22710 24268
rect 22741 24259 22799 24265
rect 22741 24256 22753 24259
rect 22704 24228 22753 24256
rect 22704 24216 22710 24228
rect 22741 24225 22753 24228
rect 22787 24225 22799 24259
rect 23658 24256 23664 24268
rect 23619 24228 23664 24256
rect 22741 24219 22799 24225
rect 23658 24216 23664 24228
rect 23716 24216 23722 24268
rect 24026 24216 24032 24268
rect 24084 24256 24090 24268
rect 24305 24259 24363 24265
rect 24305 24256 24317 24259
rect 24084 24228 24317 24256
rect 24084 24216 24090 24228
rect 24305 24225 24317 24228
rect 24351 24225 24363 24259
rect 24305 24219 24363 24225
rect 24489 24259 24547 24265
rect 24489 24225 24501 24259
rect 24535 24256 24547 24259
rect 24762 24256 24768 24268
rect 24535 24228 24768 24256
rect 24535 24225 24547 24228
rect 24489 24219 24547 24225
rect 18371 24092 21404 24120
rect 22925 24123 22983 24129
rect 18371 24089 18383 24092
rect 18325 24083 18383 24089
rect 22925 24089 22937 24123
rect 22971 24120 22983 24123
rect 23676 24120 23704 24216
rect 24320 24188 24348 24219
rect 24762 24216 24768 24228
rect 24820 24216 24826 24268
rect 25038 24256 25044 24268
rect 24999 24228 25044 24256
rect 25038 24216 25044 24228
rect 25096 24216 25102 24268
rect 25682 24256 25688 24268
rect 25643 24228 25688 24256
rect 25682 24216 25688 24228
rect 25740 24216 25746 24268
rect 26528 24265 26556 24296
rect 34532 24268 34560 24296
rect 34790 24284 34796 24296
rect 34848 24284 34854 24336
rect 35894 24284 35900 24336
rect 35952 24324 35958 24336
rect 35952 24296 37780 24324
rect 35952 24284 35958 24296
rect 26513 24259 26571 24265
rect 26513 24225 26525 24259
rect 26559 24225 26571 24259
rect 26513 24219 26571 24225
rect 27430 24216 27436 24268
rect 27488 24256 27494 24268
rect 27525 24259 27583 24265
rect 27525 24256 27537 24259
rect 27488 24228 27537 24256
rect 27488 24216 27494 24228
rect 27525 24225 27537 24228
rect 27571 24225 27583 24259
rect 28258 24256 28264 24268
rect 28219 24228 28264 24256
rect 27525 24219 27583 24225
rect 28258 24216 28264 24228
rect 28316 24216 28322 24268
rect 28994 24216 29000 24268
rect 29052 24256 29058 24268
rect 29089 24259 29147 24265
rect 29089 24256 29101 24259
rect 29052 24228 29101 24256
rect 29052 24216 29058 24228
rect 29089 24225 29101 24228
rect 29135 24256 29147 24259
rect 31202 24256 31208 24268
rect 29135 24228 31208 24256
rect 29135 24225 29147 24228
rect 29089 24219 29147 24225
rect 31202 24216 31208 24228
rect 31260 24216 31266 24268
rect 31297 24259 31355 24265
rect 31297 24225 31309 24259
rect 31343 24225 31355 24259
rect 32122 24256 32128 24268
rect 32083 24228 32128 24256
rect 31297 24219 31355 24225
rect 24578 24188 24584 24200
rect 24320 24160 24584 24188
rect 24578 24148 24584 24160
rect 24636 24148 24642 24200
rect 24670 24148 24676 24200
rect 24728 24148 24734 24200
rect 26786 24188 26792 24200
rect 25884 24160 26792 24188
rect 24688 24120 24716 24148
rect 25884 24129 25912 24160
rect 26786 24148 26792 24160
rect 26844 24188 26850 24200
rect 28353 24191 28411 24197
rect 28353 24188 28365 24191
rect 26844 24160 28365 24188
rect 26844 24148 26850 24160
rect 28353 24157 28365 24160
rect 28399 24157 28411 24191
rect 29362 24188 29368 24200
rect 29323 24160 29368 24188
rect 28353 24151 28411 24157
rect 29362 24148 29368 24160
rect 29420 24148 29426 24200
rect 22971 24092 23704 24120
rect 24596 24092 24716 24120
rect 25869 24123 25927 24129
rect 22971 24089 22983 24092
rect 22925 24083 22983 24089
rect 9122 24012 9128 24064
rect 9180 24052 9186 24064
rect 10502 24052 10508 24064
rect 9180 24024 10508 24052
rect 9180 24012 9186 24024
rect 10502 24012 10508 24024
rect 10560 24012 10566 24064
rect 14918 24012 14924 24064
rect 14976 24052 14982 24064
rect 15473 24055 15531 24061
rect 15473 24052 15485 24055
rect 14976 24024 15485 24052
rect 14976 24012 14982 24024
rect 15473 24021 15485 24024
rect 15519 24021 15531 24055
rect 15473 24015 15531 24021
rect 15654 24012 15660 24064
rect 15712 24052 15718 24064
rect 19334 24052 19340 24064
rect 15712 24024 19340 24052
rect 15712 24012 15718 24024
rect 19334 24012 19340 24024
rect 19392 24012 19398 24064
rect 20254 24052 20260 24064
rect 20215 24024 20260 24052
rect 20254 24012 20260 24024
rect 20312 24012 20318 24064
rect 24596 24061 24624 24092
rect 25869 24089 25881 24123
rect 25915 24089 25927 24123
rect 25869 24083 25927 24089
rect 24581 24055 24639 24061
rect 24581 24021 24593 24055
rect 24627 24021 24639 24055
rect 24581 24015 24639 24021
rect 24670 24012 24676 24064
rect 24728 24052 24734 24064
rect 25133 24055 25191 24061
rect 25133 24052 25145 24055
rect 24728 24024 25145 24052
rect 24728 24012 24734 24024
rect 25133 24021 25145 24024
rect 25179 24021 25191 24055
rect 26694 24052 26700 24064
rect 26655 24024 26700 24052
rect 25133 24015 25191 24021
rect 26694 24012 26700 24024
rect 26752 24012 26758 24064
rect 27890 24012 27896 24064
rect 27948 24052 27954 24064
rect 30466 24052 30472 24064
rect 27948 24024 30472 24052
rect 27948 24012 27954 24024
rect 30466 24012 30472 24024
rect 30524 24012 30530 24064
rect 31312 24052 31340 24219
rect 32122 24216 32128 24228
rect 32180 24216 32186 24268
rect 32677 24259 32735 24265
rect 32677 24225 32689 24259
rect 32723 24225 32735 24259
rect 32677 24219 32735 24225
rect 32692 24188 32720 24219
rect 33410 24216 33416 24268
rect 33468 24256 33474 24268
rect 34149 24259 34207 24265
rect 34149 24256 34161 24259
rect 33468 24228 34161 24256
rect 33468 24216 33474 24228
rect 34149 24225 34161 24228
rect 34195 24225 34207 24259
rect 34514 24256 34520 24268
rect 34475 24228 34520 24256
rect 34149 24219 34207 24225
rect 34514 24216 34520 24228
rect 34572 24216 34578 24268
rect 34698 24256 34704 24268
rect 34659 24228 34704 24256
rect 34698 24216 34704 24228
rect 34756 24216 34762 24268
rect 35529 24259 35587 24265
rect 35529 24225 35541 24259
rect 35575 24225 35587 24259
rect 36262 24256 36268 24268
rect 36223 24228 36268 24256
rect 35529 24219 35587 24225
rect 33318 24188 33324 24200
rect 31588 24160 33324 24188
rect 31588 24132 31616 24160
rect 33318 24148 33324 24160
rect 33376 24148 33382 24200
rect 34238 24188 34244 24200
rect 34151 24160 34244 24188
rect 34238 24148 34244 24160
rect 34296 24188 34302 24200
rect 35544 24188 35572 24219
rect 36262 24216 36268 24228
rect 36320 24216 36326 24268
rect 36538 24256 36544 24268
rect 36499 24228 36544 24256
rect 36538 24216 36544 24228
rect 36596 24216 36602 24268
rect 36814 24256 36820 24268
rect 36775 24228 36820 24256
rect 36814 24216 36820 24228
rect 36872 24216 36878 24268
rect 37752 24265 37780 24296
rect 37737 24259 37795 24265
rect 37737 24225 37749 24259
rect 37783 24225 37795 24259
rect 37737 24219 37795 24225
rect 34296 24160 35572 24188
rect 34296 24148 34302 24160
rect 31481 24123 31539 24129
rect 31481 24089 31493 24123
rect 31527 24120 31539 24123
rect 31570 24120 31576 24132
rect 31527 24092 31576 24120
rect 31527 24089 31539 24092
rect 31481 24083 31539 24089
rect 31570 24080 31576 24092
rect 31628 24080 31634 24132
rect 32030 24080 32036 24132
rect 32088 24120 32094 24132
rect 32217 24123 32275 24129
rect 32217 24120 32229 24123
rect 32088 24092 32229 24120
rect 32088 24080 32094 24092
rect 32217 24089 32229 24092
rect 32263 24089 32275 24123
rect 32217 24083 32275 24089
rect 36354 24080 36360 24132
rect 36412 24120 36418 24132
rect 36909 24123 36967 24129
rect 36909 24120 36921 24123
rect 36412 24092 36921 24120
rect 36412 24080 36418 24092
rect 36909 24089 36921 24092
rect 36955 24089 36967 24123
rect 36909 24083 36967 24089
rect 32582 24052 32588 24064
rect 31312 24024 32588 24052
rect 32582 24012 32588 24024
rect 32640 24052 32646 24064
rect 33042 24052 33048 24064
rect 32640 24024 33048 24052
rect 32640 24012 32646 24024
rect 33042 24012 33048 24024
rect 33100 24012 33106 24064
rect 33597 24055 33655 24061
rect 33597 24021 33609 24055
rect 33643 24052 33655 24055
rect 33686 24052 33692 24064
rect 33643 24024 33692 24052
rect 33643 24021 33655 24024
rect 33597 24015 33655 24021
rect 33686 24012 33692 24024
rect 33744 24012 33750 24064
rect 1104 23962 38824 23984
rect 1104 23910 4246 23962
rect 4298 23910 4310 23962
rect 4362 23910 4374 23962
rect 4426 23910 4438 23962
rect 4490 23910 34966 23962
rect 35018 23910 35030 23962
rect 35082 23910 35094 23962
rect 35146 23910 35158 23962
rect 35210 23910 38824 23962
rect 1104 23888 38824 23910
rect 7377 23851 7435 23857
rect 7377 23817 7389 23851
rect 7423 23848 7435 23851
rect 7926 23848 7932 23860
rect 7423 23820 7932 23848
rect 7423 23817 7435 23820
rect 7377 23811 7435 23817
rect 7926 23808 7932 23820
rect 7984 23848 7990 23860
rect 9214 23848 9220 23860
rect 7984 23820 9220 23848
rect 7984 23808 7990 23820
rect 9214 23808 9220 23820
rect 9272 23808 9278 23860
rect 23014 23848 23020 23860
rect 22975 23820 23020 23848
rect 23014 23808 23020 23820
rect 23072 23808 23078 23860
rect 23198 23808 23204 23860
rect 23256 23848 23262 23860
rect 23937 23851 23995 23857
rect 23937 23848 23949 23851
rect 23256 23820 23949 23848
rect 23256 23808 23262 23820
rect 23937 23817 23949 23820
rect 23983 23817 23995 23851
rect 23937 23811 23995 23817
rect 24026 23808 24032 23860
rect 24084 23848 24090 23860
rect 25038 23848 25044 23860
rect 24084 23820 25044 23848
rect 24084 23808 24090 23820
rect 25038 23808 25044 23820
rect 25096 23808 25102 23860
rect 29362 23808 29368 23860
rect 29420 23848 29426 23860
rect 29641 23851 29699 23857
rect 29641 23848 29653 23851
rect 29420 23820 29653 23848
rect 29420 23808 29426 23820
rect 29641 23817 29653 23820
rect 29687 23817 29699 23851
rect 32122 23848 32128 23860
rect 29641 23811 29699 23817
rect 30668 23820 32128 23848
rect 14277 23783 14335 23789
rect 11072 23752 13584 23780
rect 11072 23724 11100 23752
rect 1670 23672 1676 23724
rect 1728 23712 1734 23724
rect 1857 23715 1915 23721
rect 1857 23712 1869 23715
rect 1728 23684 1869 23712
rect 1728 23672 1734 23684
rect 1857 23681 1869 23684
rect 1903 23681 1915 23715
rect 2406 23712 2412 23724
rect 2367 23684 2412 23712
rect 1857 23675 1915 23681
rect 2406 23672 2412 23684
rect 2464 23672 2470 23724
rect 3142 23712 3148 23724
rect 2700 23684 3148 23712
rect 2700 23653 2728 23684
rect 3142 23672 3148 23684
rect 3200 23672 3206 23724
rect 5813 23715 5871 23721
rect 5813 23712 5825 23715
rect 4356 23684 5825 23712
rect 2685 23647 2743 23653
rect 2685 23613 2697 23647
rect 2731 23613 2743 23647
rect 2866 23644 2872 23656
rect 2827 23616 2872 23644
rect 2685 23607 2743 23613
rect 2866 23604 2872 23616
rect 2924 23604 2930 23656
rect 3326 23644 3332 23656
rect 3287 23616 3332 23644
rect 3326 23604 3332 23616
rect 3384 23604 3390 23656
rect 4356 23653 4384 23684
rect 5813 23681 5825 23684
rect 5859 23681 5871 23715
rect 5813 23675 5871 23681
rect 6178 23672 6184 23724
rect 6236 23712 6242 23724
rect 8021 23715 8079 23721
rect 8021 23712 8033 23715
rect 6236 23684 8033 23712
rect 6236 23672 6242 23684
rect 8021 23681 8033 23684
rect 8067 23681 8079 23715
rect 9858 23712 9864 23724
rect 8021 23675 8079 23681
rect 8956 23684 9864 23712
rect 4341 23647 4399 23653
rect 4341 23613 4353 23647
rect 4387 23613 4399 23647
rect 4341 23607 4399 23613
rect 5169 23647 5227 23653
rect 5169 23613 5181 23647
rect 5215 23613 5227 23647
rect 5442 23644 5448 23656
rect 5403 23616 5448 23644
rect 5169 23607 5227 23613
rect 3421 23579 3479 23585
rect 3421 23545 3433 23579
rect 3467 23576 3479 23579
rect 4614 23576 4620 23588
rect 3467 23548 4620 23576
rect 3467 23545 3479 23548
rect 3421 23539 3479 23545
rect 4614 23536 4620 23548
rect 4672 23536 4678 23588
rect 5184 23576 5212 23607
rect 5442 23604 5448 23616
rect 5500 23604 5506 23656
rect 5905 23647 5963 23653
rect 5905 23613 5917 23647
rect 5951 23644 5963 23647
rect 6546 23644 6552 23656
rect 5951 23616 6552 23644
rect 5951 23613 5963 23616
rect 5905 23607 5963 23613
rect 6546 23604 6552 23616
rect 6604 23604 6610 23656
rect 7193 23647 7251 23653
rect 7193 23613 7205 23647
rect 7239 23644 7251 23647
rect 7282 23644 7288 23656
rect 7239 23616 7288 23644
rect 7239 23613 7251 23616
rect 7193 23607 7251 23613
rect 7282 23604 7288 23616
rect 7340 23604 7346 23656
rect 8110 23644 8116 23656
rect 8071 23616 8116 23644
rect 8110 23604 8116 23616
rect 8168 23604 8174 23656
rect 8570 23644 8576 23656
rect 8531 23616 8576 23644
rect 8570 23604 8576 23616
rect 8628 23604 8634 23656
rect 8956 23653 8984 23684
rect 9858 23672 9864 23684
rect 9916 23672 9922 23724
rect 10318 23712 10324 23724
rect 10060 23684 10324 23712
rect 8941 23647 8999 23653
rect 8941 23613 8953 23647
rect 8987 23613 8999 23647
rect 8941 23607 8999 23613
rect 9401 23647 9459 23653
rect 9401 23613 9413 23647
rect 9447 23644 9459 23647
rect 10060 23644 10088 23684
rect 10318 23672 10324 23684
rect 10376 23672 10382 23724
rect 10686 23712 10692 23724
rect 10647 23684 10692 23712
rect 10686 23672 10692 23684
rect 10744 23672 10750 23724
rect 11054 23712 11060 23724
rect 10980 23684 11060 23712
rect 9447 23616 10088 23644
rect 10137 23647 10195 23653
rect 9447 23613 9459 23616
rect 9401 23607 9459 23613
rect 10137 23613 10149 23647
rect 10183 23644 10195 23647
rect 10980 23644 11008 23684
rect 11054 23672 11060 23684
rect 11112 23672 11118 23724
rect 11517 23715 11575 23721
rect 11517 23681 11529 23715
rect 11563 23712 11575 23715
rect 12618 23712 12624 23724
rect 11563 23684 12624 23712
rect 11563 23681 11575 23684
rect 11517 23675 11575 23681
rect 12618 23672 12624 23684
rect 12676 23672 12682 23724
rect 13556 23721 13584 23752
rect 14277 23749 14289 23783
rect 14323 23780 14335 23783
rect 14550 23780 14556 23792
rect 14323 23752 14556 23780
rect 14323 23749 14335 23752
rect 14277 23743 14335 23749
rect 14550 23740 14556 23752
rect 14608 23740 14614 23792
rect 17126 23780 17132 23792
rect 17087 23752 17132 23780
rect 17126 23740 17132 23752
rect 17184 23740 17190 23792
rect 21358 23780 21364 23792
rect 19076 23752 21364 23780
rect 13081 23715 13139 23721
rect 13081 23681 13093 23715
rect 13127 23712 13139 23715
rect 13541 23715 13599 23721
rect 13127 23684 13492 23712
rect 13127 23681 13139 23684
rect 13081 23675 13139 23681
rect 11146 23644 11152 23656
rect 10183 23616 11008 23644
rect 11107 23616 11152 23644
rect 10183 23613 10195 23616
rect 10137 23607 10195 23613
rect 11146 23604 11152 23616
rect 11204 23604 11210 23656
rect 11698 23644 11704 23656
rect 11659 23616 11704 23644
rect 11698 23604 11704 23616
rect 11756 23604 11762 23656
rect 12526 23644 12532 23656
rect 12487 23616 12532 23644
rect 12526 23604 12532 23616
rect 12584 23604 12590 23656
rect 13357 23647 13415 23653
rect 13357 23613 13369 23647
rect 13403 23613 13415 23647
rect 13464 23644 13492 23684
rect 13541 23681 13553 23715
rect 13587 23681 13599 23715
rect 14642 23712 14648 23724
rect 13541 23675 13599 23681
rect 14108 23684 14648 23712
rect 14108 23644 14136 23684
rect 14642 23672 14648 23684
rect 14700 23672 14706 23724
rect 15930 23712 15936 23724
rect 14752 23684 15936 23712
rect 14752 23653 14780 23684
rect 15930 23672 15936 23684
rect 15988 23672 15994 23724
rect 13464 23616 14136 23644
rect 14185 23647 14243 23653
rect 13357 23607 13415 23613
rect 14185 23613 14197 23647
rect 14231 23613 14243 23647
rect 14185 23607 14243 23613
rect 14737 23647 14795 23653
rect 14737 23613 14749 23647
rect 14783 23613 14795 23647
rect 14918 23644 14924 23656
rect 14879 23616 14924 23644
rect 14737 23607 14795 23613
rect 6822 23576 6828 23588
rect 5184 23548 6828 23576
rect 6822 23536 6828 23548
rect 6880 23536 6886 23588
rect 9950 23576 9956 23588
rect 9911 23548 9956 23576
rect 9950 23536 9956 23548
rect 10008 23536 10014 23588
rect 10321 23579 10379 23585
rect 10321 23576 10333 23579
rect 10060 23548 10333 23576
rect 4433 23511 4491 23517
rect 4433 23477 4445 23511
rect 4479 23508 4491 23511
rect 4522 23508 4528 23520
rect 4479 23480 4528 23508
rect 4479 23477 4491 23480
rect 4433 23471 4491 23477
rect 4522 23468 4528 23480
rect 4580 23468 4586 23520
rect 8662 23468 8668 23520
rect 8720 23508 8726 23520
rect 10060 23508 10088 23548
rect 10321 23545 10333 23548
rect 10367 23545 10379 23579
rect 10321 23539 10379 23545
rect 8720 23480 10088 23508
rect 10229 23511 10287 23517
rect 8720 23468 8726 23480
rect 10229 23477 10241 23511
rect 10275 23508 10287 23511
rect 10962 23508 10968 23520
rect 10275 23480 10968 23508
rect 10275 23477 10287 23480
rect 10229 23471 10287 23477
rect 10962 23468 10968 23480
rect 11020 23468 11026 23520
rect 13372 23508 13400 23607
rect 14200 23576 14228 23607
rect 14918 23604 14924 23616
rect 14976 23604 14982 23656
rect 15470 23604 15476 23656
rect 15528 23644 15534 23656
rect 15565 23647 15623 23653
rect 15565 23644 15577 23647
rect 15528 23616 15577 23644
rect 15528 23604 15534 23616
rect 15565 23613 15577 23616
rect 15611 23644 15623 23647
rect 16206 23644 16212 23656
rect 15611 23616 16212 23644
rect 15611 23613 15623 23616
rect 15565 23607 15623 23613
rect 16206 23604 16212 23616
rect 16264 23604 16270 23656
rect 16393 23647 16451 23653
rect 16393 23613 16405 23647
rect 16439 23644 16451 23647
rect 16574 23644 16580 23656
rect 16439 23616 16580 23644
rect 16439 23613 16451 23616
rect 16393 23607 16451 23613
rect 16574 23604 16580 23616
rect 16632 23604 16638 23656
rect 16761 23647 16819 23653
rect 16761 23613 16773 23647
rect 16807 23613 16819 23647
rect 17126 23644 17132 23656
rect 17087 23616 17132 23644
rect 16761 23607 16819 23613
rect 15378 23576 15384 23588
rect 14200 23548 15384 23576
rect 15378 23536 15384 23548
rect 15436 23536 15442 23588
rect 16776 23576 16804 23607
rect 17126 23604 17132 23616
rect 17184 23604 17190 23656
rect 18506 23644 18512 23656
rect 18467 23616 18512 23644
rect 18506 23604 18512 23616
rect 18564 23604 18570 23656
rect 18969 23647 19027 23653
rect 18969 23613 18981 23647
rect 19015 23644 19027 23647
rect 19076 23644 19104 23752
rect 21358 23740 21364 23752
rect 21416 23740 21422 23792
rect 22370 23740 22376 23792
rect 22428 23780 22434 23792
rect 22428 23752 24992 23780
rect 22428 23740 22434 23752
rect 19334 23712 19340 23724
rect 19295 23684 19340 23712
rect 19334 23672 19340 23684
rect 19392 23672 19398 23724
rect 20441 23715 20499 23721
rect 20441 23681 20453 23715
rect 20487 23712 20499 23715
rect 21726 23712 21732 23724
rect 20487 23684 21732 23712
rect 20487 23681 20499 23684
rect 20441 23675 20499 23681
rect 21726 23672 21732 23684
rect 21784 23672 21790 23724
rect 22002 23672 22008 23724
rect 22060 23712 22066 23724
rect 22189 23715 22247 23721
rect 22189 23712 22201 23715
rect 22060 23684 22201 23712
rect 22060 23672 22066 23684
rect 22189 23681 22201 23684
rect 22235 23681 22247 23715
rect 23934 23712 23940 23724
rect 22189 23675 22247 23681
rect 22848 23684 23940 23712
rect 19242 23644 19248 23656
rect 19015 23616 19104 23644
rect 19203 23616 19248 23644
rect 19015 23613 19027 23616
rect 18969 23607 19027 23613
rect 19242 23604 19248 23616
rect 19300 23604 19306 23656
rect 20349 23647 20407 23653
rect 20349 23613 20361 23647
rect 20395 23644 20407 23647
rect 20622 23644 20628 23656
rect 20395 23616 20628 23644
rect 20395 23613 20407 23616
rect 20349 23607 20407 23613
rect 20622 23604 20628 23616
rect 20680 23604 20686 23656
rect 20809 23647 20867 23653
rect 20809 23613 20821 23647
rect 20855 23613 20867 23647
rect 20809 23607 20867 23613
rect 17402 23576 17408 23588
rect 16776 23548 17408 23576
rect 17402 23536 17408 23548
rect 17460 23536 17466 23588
rect 20824 23576 20852 23607
rect 21174 23604 21180 23656
rect 21232 23644 21238 23656
rect 21545 23647 21603 23653
rect 21545 23644 21557 23647
rect 21232 23616 21557 23644
rect 21232 23604 21238 23616
rect 21545 23613 21557 23616
rect 21591 23644 21603 23647
rect 21591 23616 21680 23644
rect 21591 23613 21603 23616
rect 21545 23607 21603 23613
rect 21652 23576 21680 23616
rect 22094 23604 22100 23656
rect 22152 23644 22158 23656
rect 22738 23644 22744 23656
rect 22152 23616 22744 23644
rect 22152 23604 22158 23616
rect 22738 23604 22744 23616
rect 22796 23604 22802 23656
rect 22848 23653 22876 23684
rect 23934 23672 23940 23684
rect 23992 23712 23998 23724
rect 24670 23712 24676 23724
rect 23992 23684 24676 23712
rect 23992 23672 23998 23684
rect 24670 23672 24676 23684
rect 24728 23672 24734 23724
rect 24964 23721 24992 23752
rect 24949 23715 25007 23721
rect 24949 23681 24961 23715
rect 24995 23681 25007 23715
rect 24949 23675 25007 23681
rect 26513 23715 26571 23721
rect 26513 23681 26525 23715
rect 26559 23712 26571 23715
rect 26694 23712 26700 23724
rect 26559 23684 26700 23712
rect 26559 23681 26571 23684
rect 26513 23675 26571 23681
rect 26694 23672 26700 23684
rect 26752 23672 26758 23724
rect 30668 23721 30696 23820
rect 32122 23808 32128 23820
rect 32180 23848 32186 23860
rect 32585 23851 32643 23857
rect 32585 23848 32597 23851
rect 32180 23820 32597 23848
rect 32180 23808 32186 23820
rect 32585 23817 32597 23820
rect 32631 23817 32643 23851
rect 32585 23811 32643 23817
rect 30101 23715 30159 23721
rect 30101 23681 30113 23715
rect 30147 23681 30159 23715
rect 30101 23675 30159 23681
rect 30653 23715 30711 23721
rect 30653 23681 30665 23715
rect 30699 23681 30711 23715
rect 30653 23675 30711 23681
rect 22833 23647 22891 23653
rect 22833 23613 22845 23647
rect 22879 23613 22891 23647
rect 24486 23644 24492 23656
rect 24447 23616 24492 23644
rect 22833 23607 22891 23613
rect 24486 23604 24492 23616
rect 24544 23604 24550 23656
rect 24581 23647 24639 23653
rect 24581 23613 24593 23647
rect 24627 23613 24639 23647
rect 24854 23644 24860 23656
rect 24815 23616 24860 23644
rect 24581 23607 24639 23613
rect 22646 23576 22652 23588
rect 20824 23548 21588 23576
rect 21652 23548 22652 23576
rect 15102 23508 15108 23520
rect 13372 23480 15108 23508
rect 15102 23468 15108 23480
rect 15160 23508 15166 23520
rect 21560 23517 21588 23548
rect 22646 23536 22652 23548
rect 22704 23536 22710 23588
rect 24596 23576 24624 23607
rect 24854 23604 24860 23616
rect 24912 23604 24918 23656
rect 26786 23644 26792 23656
rect 26747 23616 26792 23644
rect 26786 23604 26792 23616
rect 26844 23604 26850 23656
rect 26970 23644 26976 23656
rect 26931 23616 26976 23644
rect 26970 23604 26976 23616
rect 27028 23604 27034 23656
rect 27709 23647 27767 23653
rect 27709 23613 27721 23647
rect 27755 23613 27767 23647
rect 27709 23607 27767 23613
rect 25682 23576 25688 23588
rect 22940 23548 24532 23576
rect 24596 23548 25688 23576
rect 15657 23511 15715 23517
rect 15657 23508 15669 23511
rect 15160 23480 15669 23508
rect 15160 23468 15166 23480
rect 15657 23477 15669 23480
rect 15703 23477 15715 23511
rect 15657 23471 15715 23477
rect 21545 23511 21603 23517
rect 21545 23477 21557 23511
rect 21591 23508 21603 23511
rect 22940 23508 22968 23548
rect 21591 23480 22968 23508
rect 24504 23508 24532 23548
rect 25682 23536 25688 23548
rect 25740 23536 25746 23588
rect 25961 23579 26019 23585
rect 25961 23545 25973 23579
rect 26007 23576 26019 23579
rect 26602 23576 26608 23588
rect 26007 23548 26608 23576
rect 26007 23545 26019 23548
rect 25961 23539 26019 23545
rect 26602 23536 26608 23548
rect 26660 23536 26666 23588
rect 27724 23576 27752 23607
rect 27890 23604 27896 23656
rect 27948 23644 27954 23656
rect 28261 23647 28319 23653
rect 28261 23644 28273 23647
rect 27948 23616 28273 23644
rect 27948 23604 27954 23616
rect 28261 23613 28273 23616
rect 28307 23613 28319 23647
rect 28261 23607 28319 23613
rect 28445 23647 28503 23653
rect 28445 23613 28457 23647
rect 28491 23644 28503 23647
rect 28626 23644 28632 23656
rect 28491 23616 28632 23644
rect 28491 23613 28503 23616
rect 28445 23607 28503 23613
rect 28626 23604 28632 23616
rect 28684 23604 28690 23656
rect 29546 23576 29552 23588
rect 27724 23548 29552 23576
rect 29546 23536 29552 23548
rect 29604 23576 29610 23588
rect 29914 23576 29920 23588
rect 29604 23548 29920 23576
rect 29604 23536 29610 23548
rect 29914 23536 29920 23548
rect 29972 23536 29978 23588
rect 26142 23508 26148 23520
rect 24504 23480 26148 23508
rect 21591 23477 21603 23480
rect 21545 23471 21603 23477
rect 26142 23468 26148 23480
rect 26200 23468 26206 23520
rect 27706 23508 27712 23520
rect 27667 23480 27712 23508
rect 27706 23468 27712 23480
rect 27764 23468 27770 23520
rect 29638 23468 29644 23520
rect 29696 23508 29702 23520
rect 30116 23508 30144 23675
rect 31018 23672 31024 23724
rect 31076 23712 31082 23724
rect 31478 23712 31484 23724
rect 31076 23684 31340 23712
rect 31439 23684 31484 23712
rect 31076 23672 31082 23684
rect 30193 23647 30251 23653
rect 30193 23613 30205 23647
rect 30239 23613 30251 23647
rect 30558 23644 30564 23656
rect 30519 23616 30564 23644
rect 30193 23607 30251 23613
rect 30208 23576 30236 23607
rect 30558 23604 30564 23616
rect 30616 23604 30622 23656
rect 31202 23644 31208 23656
rect 31163 23616 31208 23644
rect 31202 23604 31208 23616
rect 31260 23604 31266 23656
rect 31312 23644 31340 23684
rect 31478 23672 31484 23684
rect 31536 23672 31542 23724
rect 35710 23712 35716 23724
rect 33888 23684 35480 23712
rect 35671 23684 35716 23712
rect 33888 23653 33916 23684
rect 33873 23647 33931 23653
rect 33873 23644 33885 23647
rect 31312 23616 33885 23644
rect 33873 23613 33885 23616
rect 33919 23613 33931 23647
rect 33873 23607 33931 23613
rect 34149 23647 34207 23653
rect 34149 23613 34161 23647
rect 34195 23644 34207 23647
rect 34790 23644 34796 23656
rect 34195 23616 34796 23644
rect 34195 23613 34207 23616
rect 34149 23607 34207 23613
rect 34790 23604 34796 23616
rect 34848 23604 34854 23656
rect 35452 23653 35480 23684
rect 35710 23672 35716 23684
rect 35768 23672 35774 23724
rect 36078 23672 36084 23724
rect 36136 23712 36142 23724
rect 36449 23715 36507 23721
rect 36449 23712 36461 23715
rect 36136 23684 36461 23712
rect 36136 23672 36142 23684
rect 36449 23681 36461 23684
rect 36495 23681 36507 23715
rect 36814 23712 36820 23724
rect 36449 23675 36507 23681
rect 36556 23684 36820 23712
rect 35437 23647 35495 23653
rect 35437 23613 35449 23647
rect 35483 23644 35495 23647
rect 35526 23644 35532 23656
rect 35483 23616 35532 23644
rect 35483 23613 35495 23616
rect 35437 23607 35495 23613
rect 35526 23604 35532 23616
rect 35584 23604 35590 23656
rect 35621 23647 35679 23653
rect 35621 23613 35633 23647
rect 35667 23644 35679 23647
rect 36556 23644 36584 23684
rect 36814 23672 36820 23684
rect 36872 23672 36878 23724
rect 36722 23644 36728 23656
rect 35667 23616 36584 23644
rect 36683 23616 36728 23644
rect 35667 23613 35679 23616
rect 35621 23607 35679 23613
rect 36722 23604 36728 23616
rect 36780 23604 36786 23656
rect 30374 23576 30380 23588
rect 30208 23548 30380 23576
rect 30374 23536 30380 23548
rect 30432 23536 30438 23588
rect 34330 23576 34336 23588
rect 34291 23548 34336 23576
rect 34330 23536 34336 23548
rect 34388 23536 34394 23588
rect 34238 23508 34244 23520
rect 29696 23480 34244 23508
rect 29696 23468 29702 23480
rect 34238 23468 34244 23480
rect 34296 23468 34302 23520
rect 37826 23508 37832 23520
rect 37787 23480 37832 23508
rect 37826 23468 37832 23480
rect 37884 23468 37890 23520
rect 1104 23418 38824 23440
rect 1104 23366 19606 23418
rect 19658 23366 19670 23418
rect 19722 23366 19734 23418
rect 19786 23366 19798 23418
rect 19850 23366 38824 23418
rect 1104 23344 38824 23366
rect 7558 23304 7564 23316
rect 2976 23276 7564 23304
rect 2976 23177 3004 23276
rect 7558 23264 7564 23276
rect 7616 23264 7622 23316
rect 8478 23264 8484 23316
rect 8536 23304 8542 23316
rect 8662 23304 8668 23316
rect 8536 23276 8668 23304
rect 8536 23264 8542 23276
rect 8662 23264 8668 23276
rect 8720 23264 8726 23316
rect 14366 23264 14372 23316
rect 14424 23304 14430 23316
rect 15010 23304 15016 23316
rect 14424 23276 15016 23304
rect 14424 23264 14430 23276
rect 15010 23264 15016 23276
rect 15068 23304 15074 23316
rect 17126 23304 17132 23316
rect 15068 23276 16804 23304
rect 17087 23276 17132 23304
rect 15068 23264 15074 23276
rect 7282 23236 7288 23248
rect 6748 23208 7288 23236
rect 1673 23171 1731 23177
rect 1673 23137 1685 23171
rect 1719 23137 1731 23171
rect 1673 23131 1731 23137
rect 2593 23171 2651 23177
rect 2593 23137 2605 23171
rect 2639 23137 2651 23171
rect 2593 23131 2651 23137
rect 2961 23171 3019 23177
rect 2961 23137 2973 23171
rect 3007 23137 3019 23171
rect 2961 23131 3019 23137
rect 3329 23171 3387 23177
rect 3329 23137 3341 23171
rect 3375 23168 3387 23171
rect 3602 23168 3608 23180
rect 3375 23140 3608 23168
rect 3375 23137 3387 23140
rect 3329 23131 3387 23137
rect 1688 23100 1716 23131
rect 2409 23103 2467 23109
rect 2409 23100 2421 23103
rect 1688 23072 2421 23100
rect 2409 23069 2421 23072
rect 2455 23069 2467 23103
rect 2608 23100 2636 23131
rect 3602 23128 3608 23140
rect 3660 23128 3666 23180
rect 4522 23168 4528 23180
rect 4483 23140 4528 23168
rect 4522 23128 4528 23140
rect 4580 23128 4586 23180
rect 6748 23177 6776 23208
rect 7282 23196 7288 23208
rect 7340 23196 7346 23248
rect 9398 23196 9404 23248
rect 9456 23236 9462 23248
rect 12526 23236 12532 23248
rect 9456 23208 12532 23236
rect 9456 23196 9462 23208
rect 6733 23171 6791 23177
rect 6733 23137 6745 23171
rect 6779 23137 6791 23171
rect 6733 23131 6791 23137
rect 6822 23128 6828 23180
rect 6880 23168 6886 23180
rect 6917 23171 6975 23177
rect 6917 23168 6929 23171
rect 6880 23140 6929 23168
rect 6880 23128 6886 23140
rect 6917 23137 6929 23140
rect 6963 23137 6975 23171
rect 7374 23168 7380 23180
rect 7335 23140 7380 23168
rect 6917 23131 6975 23137
rect 7374 23128 7380 23140
rect 7432 23128 7438 23180
rect 7929 23171 7987 23177
rect 7929 23137 7941 23171
rect 7975 23137 7987 23171
rect 8110 23168 8116 23180
rect 8071 23140 8116 23168
rect 7929 23131 7987 23137
rect 4062 23100 4068 23112
rect 2608 23072 4068 23100
rect 2409 23063 2467 23069
rect 4062 23060 4068 23072
rect 4120 23060 4126 23112
rect 4249 23103 4307 23109
rect 4249 23069 4261 23103
rect 4295 23100 4307 23103
rect 4706 23100 4712 23112
rect 4295 23072 4712 23100
rect 4295 23069 4307 23072
rect 4249 23063 4307 23069
rect 1394 22992 1400 23044
rect 1452 23032 1458 23044
rect 4264 23032 4292 23063
rect 4706 23060 4712 23072
rect 4764 23060 4770 23112
rect 7944 23100 7972 23131
rect 8110 23128 8116 23140
rect 8168 23128 8174 23180
rect 8846 23168 8852 23180
rect 8759 23140 8852 23168
rect 8846 23128 8852 23140
rect 8904 23168 8910 23180
rect 9306 23168 9312 23180
rect 8904 23140 9312 23168
rect 8904 23128 8910 23140
rect 9306 23128 9312 23140
rect 9364 23128 9370 23180
rect 11348 23177 11376 23208
rect 12526 23196 12532 23208
rect 12584 23236 12590 23248
rect 13262 23236 13268 23248
rect 12584 23208 13268 23236
rect 12584 23196 12590 23208
rect 13262 23196 13268 23208
rect 13320 23196 13326 23248
rect 16666 23236 16672 23248
rect 15488 23208 16672 23236
rect 10689 23171 10747 23177
rect 10689 23137 10701 23171
rect 10735 23137 10747 23171
rect 10689 23131 10747 23137
rect 11333 23171 11391 23177
rect 11333 23137 11345 23171
rect 11379 23137 11391 23171
rect 11333 23131 11391 23137
rect 11425 23171 11483 23177
rect 11425 23137 11437 23171
rect 11471 23137 11483 23171
rect 12158 23168 12164 23180
rect 12119 23140 12164 23168
rect 11425 23131 11483 23137
rect 10318 23100 10324 23112
rect 7944 23072 10324 23100
rect 10318 23060 10324 23072
rect 10376 23100 10382 23112
rect 10704 23100 10732 23131
rect 11146 23100 11152 23112
rect 10376 23072 10732 23100
rect 11107 23072 11152 23100
rect 10376 23060 10382 23072
rect 11146 23060 11152 23072
rect 11204 23060 11210 23112
rect 11440 23100 11468 23131
rect 12158 23128 12164 23140
rect 12216 23128 12222 23180
rect 12618 23168 12624 23180
rect 12579 23140 12624 23168
rect 12618 23128 12624 23140
rect 12676 23128 12682 23180
rect 13817 23171 13875 23177
rect 13817 23137 13829 23171
rect 13863 23168 13875 23171
rect 13906 23168 13912 23180
rect 13863 23140 13912 23168
rect 13863 23137 13875 23140
rect 13817 23131 13875 23137
rect 13906 23128 13912 23140
rect 13964 23128 13970 23180
rect 14369 23171 14427 23177
rect 14369 23137 14381 23171
rect 14415 23168 14427 23171
rect 15286 23168 15292 23180
rect 14415 23140 15292 23168
rect 14415 23137 14427 23140
rect 14369 23131 14427 23137
rect 15286 23128 15292 23140
rect 15344 23128 15350 23180
rect 15488 23177 15516 23208
rect 16666 23196 16672 23208
rect 16724 23196 16730 23248
rect 16776 23177 16804 23276
rect 17126 23264 17132 23276
rect 17184 23264 17190 23316
rect 17328 23276 19932 23304
rect 15473 23171 15531 23177
rect 15473 23137 15485 23171
rect 15519 23137 15531 23171
rect 15473 23131 15531 23137
rect 16209 23171 16267 23177
rect 16209 23137 16221 23171
rect 16255 23137 16267 23171
rect 16209 23131 16267 23137
rect 16761 23171 16819 23177
rect 16761 23137 16773 23171
rect 16807 23168 16819 23171
rect 17328 23168 17356 23276
rect 18874 23236 18880 23248
rect 17880 23208 18880 23236
rect 17880 23177 17908 23208
rect 18874 23196 18880 23208
rect 18932 23236 18938 23248
rect 19242 23236 19248 23248
rect 18932 23208 19248 23236
rect 18932 23196 18938 23208
rect 19242 23196 19248 23208
rect 19300 23236 19306 23248
rect 19904 23236 19932 23276
rect 19978 23264 19984 23316
rect 20036 23304 20042 23316
rect 20993 23307 21051 23313
rect 20993 23304 21005 23307
rect 20036 23276 21005 23304
rect 20036 23264 20042 23276
rect 20993 23273 21005 23276
rect 21039 23273 21051 23307
rect 20993 23267 21051 23273
rect 21542 23264 21548 23316
rect 21600 23304 21606 23316
rect 27706 23304 27712 23316
rect 21600 23276 27712 23304
rect 21600 23264 21606 23276
rect 20806 23236 20812 23248
rect 19300 23208 19380 23236
rect 19904 23208 20812 23236
rect 19300 23196 19306 23208
rect 16807 23140 17356 23168
rect 17405 23171 17463 23177
rect 16807 23137 16819 23140
rect 16761 23131 16819 23137
rect 17405 23137 17417 23171
rect 17451 23137 17463 23171
rect 17405 23131 17463 23137
rect 17865 23171 17923 23177
rect 17865 23137 17877 23171
rect 17911 23137 17923 23171
rect 18506 23168 18512 23180
rect 18467 23140 18512 23168
rect 17865 23131 17923 23137
rect 14458 23100 14464 23112
rect 11348 23072 11468 23100
rect 14419 23072 14464 23100
rect 1452 23004 4292 23032
rect 1452 22992 1458 23004
rect 6546 22992 6552 23044
rect 6604 23032 6610 23044
rect 6604 23004 6649 23032
rect 6604 22992 6610 23004
rect 7374 22992 7380 23044
rect 7432 23032 7438 23044
rect 9033 23035 9091 23041
rect 9033 23032 9045 23035
rect 7432 23004 9045 23032
rect 7432 22992 7438 23004
rect 9033 23001 9045 23004
rect 9079 23032 9091 23035
rect 9950 23032 9956 23044
rect 9079 23004 9956 23032
rect 9079 23001 9091 23004
rect 9033 22995 9091 23001
rect 9950 22992 9956 23004
rect 10008 23032 10014 23044
rect 11348 23032 11376 23072
rect 14458 23060 14464 23072
rect 14516 23100 14522 23112
rect 14918 23100 14924 23112
rect 14516 23072 14924 23100
rect 14516 23060 14522 23072
rect 14918 23060 14924 23072
rect 14976 23060 14982 23112
rect 10008 23004 11376 23032
rect 13909 23035 13967 23041
rect 10008 22992 10014 23004
rect 13909 23001 13921 23035
rect 13955 23032 13967 23035
rect 13998 23032 14004 23044
rect 13955 23004 14004 23032
rect 13955 23001 13967 23004
rect 13909 22995 13967 23001
rect 13998 22992 14004 23004
rect 14056 22992 14062 23044
rect 15102 22992 15108 23044
rect 15160 23032 15166 23044
rect 15657 23035 15715 23041
rect 15657 23032 15669 23035
rect 15160 23004 15669 23032
rect 15160 22992 15166 23004
rect 15657 23001 15669 23004
rect 15703 23032 15715 23035
rect 16224 23032 16252 23131
rect 17420 23100 17448 23131
rect 18506 23128 18512 23140
rect 18564 23128 18570 23180
rect 19058 23168 19064 23180
rect 19019 23140 19064 23168
rect 19058 23128 19064 23140
rect 19116 23128 19122 23180
rect 19352 23177 19380 23208
rect 20806 23196 20812 23208
rect 20864 23236 20870 23248
rect 22370 23236 22376 23248
rect 20864 23208 22376 23236
rect 20864 23196 20870 23208
rect 22370 23196 22376 23208
rect 22428 23196 22434 23248
rect 24026 23236 24032 23248
rect 22480 23208 24032 23236
rect 19337 23171 19395 23177
rect 19337 23137 19349 23171
rect 19383 23137 19395 23171
rect 20070 23168 20076 23180
rect 20031 23140 20076 23168
rect 19337 23131 19395 23137
rect 20070 23128 20076 23140
rect 20128 23128 20134 23180
rect 21174 23168 21180 23180
rect 21135 23140 21180 23168
rect 21174 23128 21180 23140
rect 21232 23128 21238 23180
rect 21729 23171 21787 23177
rect 21729 23137 21741 23171
rect 21775 23168 21787 23171
rect 21910 23168 21916 23180
rect 21775 23140 21916 23168
rect 21775 23137 21787 23140
rect 21729 23131 21787 23137
rect 21910 23128 21916 23140
rect 21968 23128 21974 23180
rect 22480 23177 22508 23208
rect 24026 23196 24032 23208
rect 24084 23196 24090 23248
rect 24320 23245 24348 23276
rect 27706 23264 27712 23276
rect 27764 23264 27770 23316
rect 28077 23307 28135 23313
rect 28077 23273 28089 23307
rect 28123 23304 28135 23307
rect 28994 23304 29000 23316
rect 28123 23276 29000 23304
rect 28123 23273 28135 23276
rect 28077 23267 28135 23273
rect 28994 23264 29000 23276
rect 29052 23304 29058 23316
rect 29052 23276 30328 23304
rect 29052 23264 29058 23276
rect 24305 23239 24363 23245
rect 24305 23205 24317 23239
rect 24351 23205 24363 23239
rect 24305 23199 24363 23205
rect 28258 23196 28264 23248
rect 28316 23236 28322 23248
rect 29273 23239 29331 23245
rect 29273 23236 29285 23239
rect 28316 23208 29285 23236
rect 28316 23196 28322 23208
rect 29273 23205 29285 23208
rect 29319 23205 29331 23239
rect 29273 23199 29331 23205
rect 30300 23180 30328 23276
rect 30466 23264 30472 23316
rect 30524 23264 30530 23316
rect 31386 23264 31392 23316
rect 31444 23304 31450 23316
rect 31481 23307 31539 23313
rect 31481 23304 31493 23307
rect 31444 23276 31493 23304
rect 31444 23264 31450 23276
rect 31481 23273 31493 23276
rect 31527 23273 31539 23307
rect 31481 23267 31539 23273
rect 31680 23276 33272 23304
rect 22465 23171 22523 23177
rect 22465 23137 22477 23171
rect 22511 23137 22523 23171
rect 22465 23131 22523 23137
rect 23201 23171 23259 23177
rect 23201 23137 23213 23171
rect 23247 23137 23259 23171
rect 23201 23131 23259 23137
rect 21634 23100 21640 23112
rect 15703 23004 16252 23032
rect 16316 23072 17448 23100
rect 21595 23072 21640 23100
rect 15703 23001 15715 23004
rect 15657 22995 15715 23001
rect 1670 22924 1676 22976
rect 1728 22964 1734 22976
rect 1765 22967 1823 22973
rect 1765 22964 1777 22967
rect 1728 22936 1777 22964
rect 1728 22924 1734 22936
rect 1765 22933 1777 22936
rect 1811 22933 1823 22967
rect 5626 22964 5632 22976
rect 5587 22936 5632 22964
rect 1765 22927 1823 22933
rect 5626 22924 5632 22936
rect 5684 22924 5690 22976
rect 12710 22964 12716 22976
rect 12671 22936 12716 22964
rect 12710 22924 12716 22936
rect 12768 22924 12774 22976
rect 12894 22924 12900 22976
rect 12952 22964 12958 22976
rect 16316 22964 16344 23072
rect 21634 23060 21640 23072
rect 21692 23100 21698 23112
rect 21818 23100 21824 23112
rect 21692 23072 21824 23100
rect 21692 23060 21698 23072
rect 21818 23060 21824 23072
rect 21876 23100 21882 23112
rect 23216 23100 23244 23131
rect 23842 23128 23848 23180
rect 23900 23168 23906 23180
rect 24121 23171 24179 23177
rect 24121 23168 24133 23171
rect 23900 23140 24133 23168
rect 23900 23128 23906 23140
rect 24121 23137 24133 23140
rect 24167 23137 24179 23171
rect 24121 23131 24179 23137
rect 24210 23128 24216 23180
rect 24268 23168 24274 23180
rect 24673 23171 24731 23177
rect 24268 23140 24313 23168
rect 24268 23128 24274 23140
rect 24673 23137 24685 23171
rect 24719 23168 24731 23171
rect 25133 23171 25191 23177
rect 25133 23168 25145 23171
rect 24719 23140 25145 23168
rect 24719 23137 24731 23140
rect 24673 23131 24731 23137
rect 25133 23137 25145 23140
rect 25179 23137 25191 23171
rect 25133 23131 25191 23137
rect 26602 23128 26608 23180
rect 26660 23168 26666 23180
rect 26789 23171 26847 23177
rect 26789 23168 26801 23171
rect 26660 23140 26801 23168
rect 26660 23128 26666 23140
rect 26789 23137 26801 23140
rect 26835 23137 26847 23171
rect 26789 23131 26847 23137
rect 27614 23128 27620 23180
rect 27672 23168 27678 23180
rect 28629 23171 28687 23177
rect 28629 23168 28641 23171
rect 27672 23140 28641 23168
rect 27672 23128 27678 23140
rect 28629 23137 28641 23140
rect 28675 23137 28687 23171
rect 28629 23131 28687 23137
rect 29917 23171 29975 23177
rect 29917 23137 29929 23171
rect 29963 23168 29975 23171
rect 29963 23140 30236 23168
rect 29963 23137 29975 23140
rect 29917 23131 29975 23137
rect 21876 23072 23244 23100
rect 23937 23103 23995 23109
rect 21876 23060 21882 23072
rect 23937 23069 23949 23103
rect 23983 23100 23995 23103
rect 24394 23100 24400 23112
rect 23983 23072 24400 23100
rect 23983 23069 23995 23072
rect 23937 23063 23995 23069
rect 24394 23060 24400 23072
rect 24452 23100 24458 23112
rect 24854 23100 24860 23112
rect 24452 23072 24860 23100
rect 24452 23060 24458 23072
rect 24854 23060 24860 23072
rect 24912 23060 24918 23112
rect 26510 23100 26516 23112
rect 26471 23072 26516 23100
rect 26510 23060 26516 23072
rect 26568 23060 26574 23112
rect 26694 23060 26700 23112
rect 26752 23100 26758 23112
rect 29822 23100 29828 23112
rect 26752 23072 29828 23100
rect 26752 23060 26758 23072
rect 29822 23060 29828 23072
rect 29880 23060 29886 23112
rect 30006 23100 30012 23112
rect 29967 23072 30012 23100
rect 30006 23060 30012 23072
rect 30064 23060 30070 23112
rect 30208 23100 30236 23140
rect 30282 23128 30288 23180
rect 30340 23168 30346 23180
rect 30484 23177 30512 23264
rect 31202 23196 31208 23248
rect 31260 23236 31266 23248
rect 31680 23236 31708 23276
rect 32398 23236 32404 23248
rect 31260 23208 31708 23236
rect 32359 23208 32404 23236
rect 31260 23196 31266 23208
rect 32398 23196 32404 23208
rect 32456 23196 32462 23248
rect 32950 23236 32956 23248
rect 32911 23208 32956 23236
rect 32950 23196 32956 23208
rect 33008 23196 33014 23248
rect 30469 23171 30527 23177
rect 30340 23140 30433 23168
rect 30340 23128 30346 23140
rect 30469 23137 30481 23171
rect 30515 23137 30527 23171
rect 31294 23168 31300 23180
rect 31255 23140 31300 23168
rect 30469 23131 30527 23137
rect 31294 23128 31300 23140
rect 31352 23128 31358 23180
rect 32585 23171 32643 23177
rect 32585 23137 32597 23171
rect 32631 23168 32643 23171
rect 32674 23168 32680 23180
rect 32631 23140 32680 23168
rect 32631 23137 32643 23140
rect 32585 23131 32643 23137
rect 32674 23128 32680 23140
rect 32732 23128 32738 23180
rect 33244 23168 33272 23276
rect 34514 23264 34520 23316
rect 34572 23304 34578 23316
rect 37829 23307 37887 23313
rect 37829 23304 37841 23307
rect 34572 23276 37841 23304
rect 34572 23264 34578 23276
rect 37829 23273 37841 23276
rect 37875 23273 37887 23307
rect 37829 23267 37887 23273
rect 33413 23171 33471 23177
rect 33413 23168 33425 23171
rect 33244 23140 33425 23168
rect 33413 23137 33425 23140
rect 33459 23137 33471 23171
rect 33686 23168 33692 23180
rect 33647 23140 33692 23168
rect 33413 23131 33471 23137
rect 33686 23128 33692 23140
rect 33744 23128 33750 23180
rect 35986 23168 35992 23180
rect 35947 23140 35992 23168
rect 35986 23128 35992 23140
rect 36044 23128 36050 23180
rect 36446 23168 36452 23180
rect 36407 23140 36452 23168
rect 36446 23128 36452 23140
rect 36504 23168 36510 23180
rect 37737 23171 37795 23177
rect 37737 23168 37749 23171
rect 36504 23140 37749 23168
rect 36504 23128 36510 23140
rect 37737 23137 37749 23140
rect 37783 23168 37795 23171
rect 37826 23168 37832 23180
rect 37783 23140 37832 23168
rect 37783 23137 37795 23140
rect 37737 23131 37795 23137
rect 37826 23128 37832 23140
rect 37884 23128 37890 23180
rect 30374 23100 30380 23112
rect 30208 23072 30380 23100
rect 30374 23060 30380 23072
rect 30432 23060 30438 23112
rect 31110 23060 31116 23112
rect 31168 23100 31174 23112
rect 31386 23100 31392 23112
rect 31168 23072 31392 23100
rect 31168 23060 31174 23072
rect 31386 23060 31392 23072
rect 31444 23060 31450 23112
rect 35894 23060 35900 23112
rect 35952 23100 35958 23112
rect 36541 23103 36599 23109
rect 36541 23100 36553 23103
rect 35952 23072 36553 23100
rect 35952 23060 35958 23072
rect 36541 23069 36553 23072
rect 36587 23069 36599 23103
rect 36541 23063 36599 23069
rect 16574 22992 16580 23044
rect 16632 23032 16638 23044
rect 19337 23035 19395 23041
rect 19337 23032 19349 23035
rect 16632 23004 19349 23032
rect 16632 22992 16638 23004
rect 19337 23001 19349 23004
rect 19383 23001 19395 23035
rect 25314 23032 25320 23044
rect 25275 23004 25320 23032
rect 19337 22995 19395 23001
rect 25314 22992 25320 23004
rect 25372 22992 25378 23044
rect 12952 22936 16344 22964
rect 12952 22924 12958 22936
rect 18966 22924 18972 22976
rect 19024 22964 19030 22976
rect 20257 22967 20315 22973
rect 20257 22964 20269 22967
rect 19024 22936 20269 22964
rect 19024 22924 19030 22936
rect 20257 22933 20269 22936
rect 20303 22933 20315 22967
rect 20257 22927 20315 22933
rect 22370 22924 22376 22976
rect 22428 22964 22434 22976
rect 22649 22967 22707 22973
rect 22649 22964 22661 22967
rect 22428 22936 22661 22964
rect 22428 22924 22434 22936
rect 22649 22933 22661 22936
rect 22695 22933 22707 22967
rect 23382 22964 23388 22976
rect 23343 22936 23388 22964
rect 22649 22927 22707 22933
rect 23382 22924 23388 22936
rect 23440 22924 23446 22976
rect 24578 22924 24584 22976
rect 24636 22964 24642 22976
rect 28721 22967 28779 22973
rect 28721 22964 28733 22967
rect 24636 22936 28733 22964
rect 24636 22924 24642 22936
rect 28721 22933 28733 22936
rect 28767 22933 28779 22967
rect 28721 22927 28779 22933
rect 34698 22924 34704 22976
rect 34756 22964 34762 22976
rect 34977 22967 35035 22973
rect 34977 22964 34989 22967
rect 34756 22936 34989 22964
rect 34756 22924 34762 22936
rect 34977 22933 34989 22936
rect 35023 22964 35035 22967
rect 35802 22964 35808 22976
rect 35023 22936 35808 22964
rect 35023 22933 35035 22936
rect 34977 22927 35035 22933
rect 35802 22924 35808 22936
rect 35860 22924 35866 22976
rect 1104 22874 38824 22896
rect 1104 22822 4246 22874
rect 4298 22822 4310 22874
rect 4362 22822 4374 22874
rect 4426 22822 4438 22874
rect 4490 22822 34966 22874
rect 35018 22822 35030 22874
rect 35082 22822 35094 22874
rect 35146 22822 35158 22874
rect 35210 22822 38824 22874
rect 1104 22800 38824 22822
rect 3142 22720 3148 22772
rect 3200 22760 3206 22772
rect 3602 22760 3608 22772
rect 3200 22732 3608 22760
rect 3200 22720 3206 22732
rect 3602 22720 3608 22732
rect 3660 22720 3666 22772
rect 4614 22720 4620 22772
rect 4672 22760 4678 22772
rect 4672 22732 15056 22760
rect 4672 22720 4678 22732
rect 7282 22652 7288 22704
rect 7340 22692 7346 22704
rect 8665 22695 8723 22701
rect 8665 22692 8677 22695
rect 7340 22664 8677 22692
rect 7340 22652 7346 22664
rect 8665 22661 8677 22664
rect 8711 22661 8723 22695
rect 8665 22655 8723 22661
rect 9674 22652 9680 22704
rect 9732 22692 9738 22704
rect 11241 22695 11299 22701
rect 11241 22692 11253 22695
rect 9732 22664 11253 22692
rect 9732 22652 9738 22664
rect 11241 22661 11253 22664
rect 11287 22661 11299 22695
rect 11241 22655 11299 22661
rect 1394 22624 1400 22636
rect 1355 22596 1400 22624
rect 1394 22584 1400 22596
rect 1452 22584 1458 22636
rect 1670 22624 1676 22636
rect 1631 22596 1676 22624
rect 1670 22584 1676 22596
rect 1728 22584 1734 22636
rect 5626 22624 5632 22636
rect 5460 22596 5632 22624
rect 3694 22556 3700 22568
rect 3655 22528 3700 22556
rect 3694 22516 3700 22528
rect 3752 22516 3758 22568
rect 3881 22559 3939 22565
rect 3881 22525 3893 22559
rect 3927 22525 3939 22559
rect 3881 22519 3939 22525
rect 4525 22559 4583 22565
rect 4525 22525 4537 22559
rect 4571 22556 4583 22559
rect 4706 22556 4712 22568
rect 4571 22528 4712 22556
rect 4571 22525 4583 22528
rect 4525 22519 4583 22525
rect 3326 22488 3332 22500
rect 2976 22460 3332 22488
rect 2976 22432 3004 22460
rect 3326 22448 3332 22460
rect 3384 22488 3390 22500
rect 3896 22488 3924 22519
rect 4706 22516 4712 22528
rect 4764 22556 4770 22568
rect 5350 22556 5356 22568
rect 4764 22528 5356 22556
rect 4764 22516 4770 22528
rect 5350 22516 5356 22528
rect 5408 22516 5414 22568
rect 5460 22565 5488 22596
rect 5626 22584 5632 22596
rect 5684 22584 5690 22636
rect 7374 22624 7380 22636
rect 7335 22596 7380 22624
rect 7374 22584 7380 22596
rect 7432 22584 7438 22636
rect 7742 22584 7748 22636
rect 7800 22624 7806 22636
rect 8113 22627 8171 22633
rect 8113 22624 8125 22627
rect 7800 22596 8125 22624
rect 7800 22584 7806 22596
rect 8113 22593 8125 22596
rect 8159 22593 8171 22627
rect 8113 22587 8171 22593
rect 8754 22584 8760 22636
rect 8812 22624 8818 22636
rect 13170 22624 13176 22636
rect 8812 22596 10088 22624
rect 8812 22584 8818 22596
rect 10060 22568 10088 22596
rect 10336 22596 12848 22624
rect 13131 22596 13176 22624
rect 10336 22568 10364 22596
rect 5445 22559 5503 22565
rect 5445 22525 5457 22559
rect 5491 22525 5503 22559
rect 5445 22519 5503 22525
rect 5534 22516 5540 22568
rect 5592 22556 5598 22568
rect 5721 22559 5779 22565
rect 5721 22556 5733 22559
rect 5592 22528 5733 22556
rect 5592 22516 5598 22528
rect 5721 22525 5733 22528
rect 5767 22525 5779 22559
rect 5721 22519 5779 22525
rect 6089 22559 6147 22565
rect 6089 22525 6101 22559
rect 6135 22556 6147 22559
rect 6135 22528 6776 22556
rect 6135 22525 6147 22528
rect 6089 22519 6147 22525
rect 3384 22460 3924 22488
rect 3384 22448 3390 22460
rect 2958 22420 2964 22432
rect 2919 22392 2964 22420
rect 2958 22380 2964 22392
rect 3016 22380 3022 22432
rect 6748 22420 6776 22528
rect 6822 22516 6828 22568
rect 6880 22556 6886 22568
rect 7561 22559 7619 22565
rect 7561 22556 7573 22559
rect 6880 22528 7573 22556
rect 6880 22516 6886 22528
rect 7561 22525 7573 22528
rect 7607 22525 7619 22559
rect 7561 22519 7619 22525
rect 7653 22559 7711 22565
rect 7653 22525 7665 22559
rect 7699 22556 7711 22559
rect 8570 22556 8576 22568
rect 7699 22528 8576 22556
rect 7699 22525 7711 22528
rect 7653 22519 7711 22525
rect 8570 22516 8576 22528
rect 8628 22516 8634 22568
rect 9398 22556 9404 22568
rect 9359 22528 9404 22556
rect 9398 22516 9404 22528
rect 9456 22516 9462 22568
rect 9582 22556 9588 22568
rect 9543 22528 9588 22556
rect 9582 22516 9588 22528
rect 9640 22516 9646 22568
rect 10042 22556 10048 22568
rect 10003 22528 10048 22556
rect 10042 22516 10048 22528
rect 10100 22516 10106 22568
rect 10318 22556 10324 22568
rect 10279 22528 10324 22556
rect 10318 22516 10324 22528
rect 10376 22516 10382 22568
rect 11330 22556 11336 22568
rect 11291 22528 11336 22556
rect 11330 22516 11336 22528
rect 11388 22516 11394 22568
rect 11885 22559 11943 22565
rect 11885 22525 11897 22559
rect 11931 22556 11943 22559
rect 12158 22556 12164 22568
rect 11931 22528 12164 22556
rect 11931 22525 11943 22528
rect 11885 22519 11943 22525
rect 12158 22516 12164 22528
rect 12216 22516 12222 22568
rect 12526 22516 12532 22568
rect 12584 22556 12590 22568
rect 12621 22559 12679 22565
rect 12621 22556 12633 22559
rect 12584 22528 12633 22556
rect 12584 22516 12590 22528
rect 12621 22525 12633 22528
rect 12667 22525 12679 22559
rect 12621 22519 12679 22525
rect 7742 22488 7748 22500
rect 7655 22460 7748 22488
rect 7742 22448 7748 22460
rect 7800 22488 7806 22500
rect 8110 22488 8116 22500
rect 7800 22460 8116 22488
rect 7800 22448 7806 22460
rect 8110 22448 8116 22460
rect 8168 22448 8174 22500
rect 9033 22491 9091 22497
rect 9033 22457 9045 22491
rect 9079 22488 9091 22491
rect 9858 22488 9864 22500
rect 9079 22460 9864 22488
rect 9079 22457 9091 22460
rect 9033 22451 9091 22457
rect 9858 22448 9864 22460
rect 9916 22448 9922 22500
rect 10410 22448 10416 22500
rect 10468 22488 10474 22500
rect 12820 22497 12848 22596
rect 13170 22584 13176 22596
rect 13228 22584 13234 22636
rect 14366 22556 14372 22568
rect 14327 22528 14372 22556
rect 14366 22516 14372 22528
rect 14424 22516 14430 22568
rect 15028 22565 15056 22732
rect 16666 22720 16672 22772
rect 16724 22760 16730 22772
rect 17218 22760 17224 22772
rect 16724 22732 17224 22760
rect 16724 22720 16730 22732
rect 17218 22720 17224 22732
rect 17276 22720 17282 22772
rect 19334 22760 19340 22772
rect 17972 22732 19340 22760
rect 16942 22652 16948 22704
rect 17000 22692 17006 22704
rect 17129 22695 17187 22701
rect 17129 22692 17141 22695
rect 17000 22664 17141 22692
rect 17000 22652 17006 22664
rect 17129 22661 17141 22664
rect 17175 22661 17187 22695
rect 17129 22655 17187 22661
rect 16485 22627 16543 22633
rect 16485 22593 16497 22627
rect 16531 22624 16543 22627
rect 17972 22624 18000 22732
rect 19334 22720 19340 22732
rect 19392 22720 19398 22772
rect 22738 22760 22744 22772
rect 22699 22732 22744 22760
rect 22738 22720 22744 22732
rect 22796 22720 22802 22772
rect 26878 22720 26884 22772
rect 26936 22760 26942 22772
rect 37458 22760 37464 22772
rect 26936 22732 28396 22760
rect 37419 22732 37464 22760
rect 26936 22720 26942 22732
rect 20257 22695 20315 22701
rect 20257 22692 20269 22695
rect 16531 22596 18000 22624
rect 19260 22664 20269 22692
rect 16531 22593 16543 22596
rect 16485 22587 16543 22593
rect 14461 22559 14519 22565
rect 14461 22525 14473 22559
rect 14507 22525 14519 22559
rect 14461 22519 14519 22525
rect 15013 22559 15071 22565
rect 15013 22525 15025 22559
rect 15059 22525 15071 22559
rect 15013 22519 15071 22525
rect 15473 22559 15531 22565
rect 15473 22525 15485 22559
rect 15519 22556 15531 22559
rect 15562 22556 15568 22568
rect 15519 22528 15568 22556
rect 15519 22525 15531 22528
rect 15473 22519 15531 22525
rect 12437 22491 12495 22497
rect 12437 22488 12449 22491
rect 10468 22460 12449 22488
rect 10468 22448 10474 22460
rect 12437 22457 12449 22460
rect 12483 22457 12495 22491
rect 12437 22451 12495 22457
rect 12805 22491 12863 22497
rect 12805 22457 12817 22491
rect 12851 22457 12863 22491
rect 14476 22488 14504 22519
rect 15562 22516 15568 22528
rect 15620 22516 15626 22568
rect 16666 22556 16672 22568
rect 16627 22528 16672 22556
rect 16666 22516 16672 22528
rect 16724 22516 16730 22568
rect 17221 22559 17279 22565
rect 17221 22525 17233 22559
rect 17267 22556 17279 22559
rect 17494 22556 17500 22568
rect 17267 22528 17500 22556
rect 17267 22525 17279 22528
rect 17221 22519 17279 22525
rect 17494 22516 17500 22528
rect 17552 22516 17558 22568
rect 19260 22565 19288 22664
rect 20257 22661 20269 22664
rect 20303 22692 20315 22695
rect 21910 22692 21916 22704
rect 20303 22664 21916 22692
rect 20303 22661 20315 22664
rect 20257 22655 20315 22661
rect 21910 22652 21916 22664
rect 21968 22692 21974 22704
rect 21968 22664 22600 22692
rect 21968 22652 21974 22664
rect 21542 22624 21548 22636
rect 20364 22596 21548 22624
rect 18049 22559 18107 22565
rect 18049 22525 18061 22559
rect 18095 22525 18107 22559
rect 18049 22519 18107 22525
rect 19245 22559 19303 22565
rect 19245 22525 19257 22559
rect 19291 22525 19303 22559
rect 19426 22556 19432 22568
rect 19387 22528 19432 22556
rect 19245 22519 19303 22525
rect 15102 22488 15108 22500
rect 14476 22460 15108 22488
rect 12805 22451 12863 22457
rect 15102 22448 15108 22460
rect 15160 22448 15166 22500
rect 18064 22488 18092 22519
rect 19426 22516 19432 22528
rect 19484 22516 19490 22568
rect 19978 22516 19984 22568
rect 20036 22556 20042 22568
rect 20364 22565 20392 22596
rect 21542 22584 21548 22596
rect 21600 22584 21606 22636
rect 20349 22559 20407 22565
rect 20349 22556 20361 22559
rect 20036 22528 20361 22556
rect 20036 22516 20042 22528
rect 20349 22525 20361 22528
rect 20395 22525 20407 22559
rect 20349 22519 20407 22525
rect 20901 22559 20959 22565
rect 20901 22525 20913 22559
rect 20947 22525 20959 22559
rect 20901 22519 20959 22525
rect 21821 22559 21879 22565
rect 21821 22525 21833 22559
rect 21867 22556 21879 22559
rect 21910 22556 21916 22568
rect 21867 22528 21916 22556
rect 21867 22525 21879 22528
rect 21821 22519 21879 22525
rect 19705 22491 19763 22497
rect 18064 22460 19656 22488
rect 8018 22420 8024 22432
rect 6748 22392 8024 22420
rect 8018 22380 8024 22392
rect 8076 22420 8082 22432
rect 12526 22420 12532 22432
rect 8076 22392 12532 22420
rect 8076 22380 8082 22392
rect 12526 22380 12532 22392
rect 12584 22380 12590 22432
rect 12713 22423 12771 22429
rect 12713 22389 12725 22423
rect 12759 22420 12771 22423
rect 13078 22420 13084 22432
rect 12759 22392 13084 22420
rect 12759 22389 12771 22392
rect 12713 22383 12771 22389
rect 13078 22380 13084 22392
rect 13136 22380 13142 22432
rect 14737 22423 14795 22429
rect 14737 22389 14749 22423
rect 14783 22420 14795 22423
rect 16114 22420 16120 22432
rect 14783 22392 16120 22420
rect 14783 22389 14795 22392
rect 14737 22383 14795 22389
rect 16114 22380 16120 22392
rect 16172 22380 16178 22432
rect 16206 22380 16212 22432
rect 16264 22420 16270 22432
rect 18233 22423 18291 22429
rect 18233 22420 18245 22423
rect 16264 22392 18245 22420
rect 16264 22380 16270 22392
rect 18233 22389 18245 22392
rect 18279 22389 18291 22423
rect 19628 22420 19656 22460
rect 19705 22457 19717 22491
rect 19751 22488 19763 22491
rect 20438 22488 20444 22500
rect 19751 22460 20444 22488
rect 19751 22457 19763 22460
rect 19705 22451 19763 22457
rect 20438 22448 20444 22460
rect 20496 22448 20502 22500
rect 20714 22448 20720 22500
rect 20772 22488 20778 22500
rect 20916 22488 20944 22519
rect 21910 22516 21916 22528
rect 21968 22556 21974 22568
rect 22370 22556 22376 22568
rect 21968 22528 22376 22556
rect 21968 22516 21974 22528
rect 22370 22516 22376 22528
rect 22428 22516 22434 22568
rect 22572 22565 22600 22664
rect 23382 22652 23388 22704
rect 23440 22652 23446 22704
rect 27724 22664 28212 22692
rect 23400 22624 23428 22652
rect 24394 22624 24400 22636
rect 23400 22596 24256 22624
rect 24307 22596 24400 22624
rect 22557 22559 22615 22565
rect 22557 22525 22569 22559
rect 22603 22525 22615 22559
rect 22557 22519 22615 22525
rect 22646 22516 22652 22568
rect 22704 22556 22710 22568
rect 23382 22556 23388 22568
rect 22704 22528 23388 22556
rect 22704 22516 22710 22528
rect 23382 22516 23388 22528
rect 23440 22556 23446 22568
rect 23661 22559 23719 22565
rect 23661 22556 23673 22559
rect 23440 22528 23673 22556
rect 23440 22516 23446 22528
rect 23661 22525 23673 22528
rect 23707 22525 23719 22559
rect 24118 22556 24124 22568
rect 24079 22528 24124 22556
rect 23661 22519 23719 22525
rect 24118 22516 24124 22528
rect 24176 22516 24182 22568
rect 24228 22556 24256 22596
rect 24394 22584 24400 22596
rect 24452 22624 24458 22636
rect 26694 22624 26700 22636
rect 24452 22596 26700 22624
rect 24452 22584 24458 22596
rect 26694 22584 26700 22596
rect 26752 22584 26758 22636
rect 26970 22584 26976 22636
rect 27028 22624 27034 22636
rect 27341 22627 27399 22633
rect 27341 22624 27353 22627
rect 27028 22596 27353 22624
rect 27028 22584 27034 22596
rect 27341 22593 27353 22596
rect 27387 22593 27399 22627
rect 27341 22587 27399 22593
rect 25869 22559 25927 22565
rect 25869 22556 25881 22559
rect 24228 22528 25881 22556
rect 25869 22525 25881 22528
rect 25915 22525 25927 22559
rect 25869 22519 25927 22525
rect 26145 22559 26203 22565
rect 26145 22525 26157 22559
rect 26191 22525 26203 22559
rect 26145 22519 26203 22525
rect 26329 22559 26387 22565
rect 26329 22525 26341 22559
rect 26375 22556 26387 22559
rect 26878 22556 26884 22568
rect 26375 22528 26884 22556
rect 26375 22525 26387 22528
rect 26329 22519 26387 22525
rect 24210 22488 24216 22500
rect 20772 22460 24216 22488
rect 20772 22448 20778 22460
rect 24210 22448 24216 22460
rect 24268 22448 24274 22500
rect 24946 22448 24952 22500
rect 25004 22488 25010 22500
rect 25317 22491 25375 22497
rect 25317 22488 25329 22491
rect 25004 22460 25329 22488
rect 25004 22448 25010 22460
rect 25317 22457 25329 22460
rect 25363 22457 25375 22491
rect 26160 22488 26188 22519
rect 26878 22516 26884 22528
rect 26936 22516 26942 22568
rect 27338 22488 27344 22500
rect 26160 22460 27344 22488
rect 25317 22451 25375 22457
rect 27338 22448 27344 22460
rect 27396 22488 27402 22500
rect 27724 22488 27752 22664
rect 27890 22624 27896 22636
rect 27851 22596 27896 22624
rect 27890 22584 27896 22596
rect 27948 22584 27954 22636
rect 27396 22460 27752 22488
rect 27908 22488 27936 22584
rect 28184 22565 28212 22664
rect 28368 22633 28396 22732
rect 37458 22720 37464 22732
rect 37516 22720 37522 22772
rect 30006 22692 30012 22704
rect 29967 22664 30012 22692
rect 30006 22652 30012 22664
rect 30064 22652 30070 22704
rect 31021 22695 31079 22701
rect 31021 22661 31033 22695
rect 31067 22661 31079 22695
rect 31021 22655 31079 22661
rect 28353 22627 28411 22633
rect 28353 22593 28365 22627
rect 28399 22624 28411 22627
rect 28626 22624 28632 22636
rect 28399 22596 28632 22624
rect 28399 22593 28411 22596
rect 28353 22587 28411 22593
rect 28626 22584 28632 22596
rect 28684 22584 28690 22636
rect 31036 22624 31064 22655
rect 28920 22596 31064 22624
rect 28169 22559 28227 22565
rect 28169 22525 28181 22559
rect 28215 22556 28227 22559
rect 28920 22556 28948 22596
rect 29546 22556 29552 22568
rect 28215 22528 28948 22556
rect 29507 22528 29552 22556
rect 28215 22525 28227 22528
rect 28169 22519 28227 22525
rect 29546 22516 29552 22528
rect 29604 22516 29610 22568
rect 29733 22559 29791 22565
rect 29733 22525 29745 22559
rect 29779 22525 29791 22559
rect 29733 22519 29791 22525
rect 30101 22559 30159 22565
rect 30101 22525 30113 22559
rect 30147 22556 30159 22559
rect 30282 22556 30288 22568
rect 30147 22528 30288 22556
rect 30147 22525 30159 22528
rect 30101 22519 30159 22525
rect 29748 22488 29776 22519
rect 30282 22516 30288 22528
rect 30340 22516 30346 22568
rect 30834 22556 30840 22568
rect 30795 22528 30840 22556
rect 30834 22516 30840 22528
rect 30892 22516 30898 22568
rect 27908 22460 29776 22488
rect 27396 22448 27402 22460
rect 20346 22420 20352 22432
rect 19628 22392 20352 22420
rect 18233 22383 18291 22389
rect 20346 22380 20352 22392
rect 20404 22380 20410 22432
rect 22005 22423 22063 22429
rect 22005 22389 22017 22423
rect 22051 22420 22063 22423
rect 22094 22420 22100 22432
rect 22051 22392 22100 22420
rect 22051 22389 22063 22392
rect 22005 22383 22063 22389
rect 22094 22380 22100 22392
rect 22152 22380 22158 22432
rect 31036 22420 31064 22596
rect 31202 22584 31208 22636
rect 31260 22624 31266 22636
rect 31573 22627 31631 22633
rect 31573 22624 31585 22627
rect 31260 22596 31585 22624
rect 31260 22584 31266 22596
rect 31573 22593 31585 22596
rect 31619 22593 31631 22627
rect 31573 22587 31631 22593
rect 31754 22584 31760 22636
rect 31812 22624 31818 22636
rect 32674 22624 32680 22636
rect 31812 22596 32680 22624
rect 31812 22584 31818 22596
rect 32674 22584 32680 22596
rect 32732 22624 32738 22636
rect 34333 22627 34391 22633
rect 32732 22596 34008 22624
rect 32732 22584 32738 22596
rect 31846 22556 31852 22568
rect 31807 22528 31852 22556
rect 31846 22516 31852 22528
rect 31904 22516 31910 22568
rect 33778 22556 33784 22568
rect 33739 22528 33784 22556
rect 33778 22516 33784 22528
rect 33836 22516 33842 22568
rect 33980 22565 34008 22596
rect 34333 22593 34345 22627
rect 34379 22624 34391 22627
rect 34606 22624 34612 22636
rect 34379 22596 34612 22624
rect 34379 22593 34391 22596
rect 34333 22587 34391 22593
rect 34606 22584 34612 22596
rect 34664 22584 34670 22636
rect 35253 22627 35311 22633
rect 35253 22593 35265 22627
rect 35299 22624 35311 22627
rect 36357 22627 36415 22633
rect 36357 22624 36369 22627
rect 35299 22596 36369 22624
rect 35299 22593 35311 22596
rect 35253 22587 35311 22593
rect 36357 22593 36369 22596
rect 36403 22593 36415 22627
rect 36357 22587 36415 22593
rect 33965 22559 34023 22565
rect 33965 22525 33977 22559
rect 34011 22525 34023 22559
rect 33965 22519 34023 22525
rect 33594 22488 33600 22500
rect 32692 22460 33600 22488
rect 32692 22420 32720 22460
rect 33594 22448 33600 22460
rect 33652 22448 33658 22500
rect 33980 22488 34008 22519
rect 34054 22516 34060 22568
rect 34112 22556 34118 22568
rect 34885 22559 34943 22565
rect 34885 22556 34897 22559
rect 34112 22528 34897 22556
rect 34112 22516 34118 22528
rect 34885 22525 34897 22528
rect 34931 22525 34943 22559
rect 34885 22519 34943 22525
rect 35342 22516 35348 22568
rect 35400 22556 35406 22568
rect 35437 22559 35495 22565
rect 35437 22556 35449 22559
rect 35400 22528 35449 22556
rect 35400 22516 35406 22528
rect 35437 22525 35449 22528
rect 35483 22525 35495 22559
rect 36078 22556 36084 22568
rect 36039 22528 36084 22556
rect 35437 22519 35495 22525
rect 36078 22516 36084 22528
rect 36136 22516 36142 22568
rect 35618 22488 35624 22500
rect 33980 22460 35624 22488
rect 35618 22448 35624 22460
rect 35676 22448 35682 22500
rect 33134 22420 33140 22432
rect 31036 22392 32720 22420
rect 33095 22392 33140 22420
rect 33134 22380 33140 22392
rect 33192 22380 33198 22432
rect 1104 22330 38824 22352
rect 1104 22278 19606 22330
rect 19658 22278 19670 22330
rect 19722 22278 19734 22330
rect 19786 22278 19798 22330
rect 19850 22278 38824 22330
rect 1104 22256 38824 22278
rect 5721 22219 5779 22225
rect 5721 22185 5733 22219
rect 5767 22216 5779 22219
rect 6822 22216 6828 22228
rect 5767 22188 6828 22216
rect 5767 22185 5779 22188
rect 5721 22179 5779 22185
rect 6822 22176 6828 22188
rect 6880 22176 6886 22228
rect 7466 22216 7472 22228
rect 7116 22188 7472 22216
rect 7116 22148 7144 22188
rect 7466 22176 7472 22188
rect 7524 22216 7530 22228
rect 8754 22216 8760 22228
rect 7524 22188 8760 22216
rect 7524 22176 7530 22188
rect 8754 22176 8760 22188
rect 8812 22176 8818 22228
rect 12250 22176 12256 22228
rect 12308 22216 12314 22228
rect 13265 22219 13323 22225
rect 13265 22216 13277 22219
rect 12308 22188 13277 22216
rect 12308 22176 12314 22188
rect 13265 22185 13277 22188
rect 13311 22216 13323 22219
rect 17494 22216 17500 22228
rect 13311 22188 15516 22216
rect 17455 22188 17500 22216
rect 13311 22185 13323 22188
rect 13265 22179 13323 22185
rect 7742 22148 7748 22160
rect 2608 22120 7144 22148
rect 7208 22120 7748 22148
rect 1762 22080 1768 22092
rect 1723 22052 1768 22080
rect 1762 22040 1768 22052
rect 1820 22040 1826 22092
rect 2608 22089 2636 22120
rect 2593 22083 2651 22089
rect 2593 22049 2605 22083
rect 2639 22049 2651 22083
rect 3142 22080 3148 22092
rect 3103 22052 3148 22080
rect 2593 22043 2651 22049
rect 3142 22040 3148 22052
rect 3200 22040 3206 22092
rect 4341 22083 4399 22089
rect 4341 22049 4353 22083
rect 4387 22080 4399 22083
rect 4614 22080 4620 22092
rect 4387 22052 4620 22080
rect 4387 22049 4399 22052
rect 4341 22043 4399 22049
rect 4614 22040 4620 22052
rect 4672 22040 4678 22092
rect 4801 22083 4859 22089
rect 4801 22049 4813 22083
rect 4847 22080 4859 22083
rect 4890 22080 4896 22092
rect 4847 22052 4896 22080
rect 4847 22049 4859 22052
rect 4801 22043 4859 22049
rect 4890 22040 4896 22052
rect 4948 22040 4954 22092
rect 5537 22083 5595 22089
rect 5537 22049 5549 22083
rect 5583 22080 5595 22083
rect 5626 22080 5632 22092
rect 5583 22052 5632 22080
rect 5583 22049 5595 22052
rect 5537 22043 5595 22049
rect 5626 22040 5632 22052
rect 5684 22040 5690 22092
rect 7208 22089 7236 22120
rect 7742 22108 7748 22120
rect 7800 22108 7806 22160
rect 8846 22148 8852 22160
rect 8496 22120 8852 22148
rect 6641 22083 6699 22089
rect 6641 22049 6653 22083
rect 6687 22049 6699 22083
rect 6641 22043 6699 22049
rect 7193 22083 7251 22089
rect 7193 22049 7205 22083
rect 7239 22080 7251 22083
rect 7653 22083 7711 22089
rect 7239 22052 7273 22080
rect 7239 22049 7251 22052
rect 7193 22043 7251 22049
rect 7653 22049 7665 22083
rect 7699 22049 7711 22083
rect 7653 22043 7711 22049
rect 8113 22083 8171 22089
rect 8113 22049 8125 22083
rect 8159 22080 8171 22083
rect 8496 22080 8524 22120
rect 8846 22108 8852 22120
rect 8904 22108 8910 22160
rect 10318 22148 10324 22160
rect 9876 22120 10324 22148
rect 8159 22052 8524 22080
rect 8159 22049 8171 22052
rect 8113 22043 8171 22049
rect 3418 22012 3424 22024
rect 3379 21984 3424 22012
rect 3418 21972 3424 21984
rect 3476 21972 3482 22024
rect 3694 21972 3700 22024
rect 3752 22012 3758 22024
rect 4062 22012 4068 22024
rect 3752 21984 4068 22012
rect 3752 21972 3758 21984
rect 4062 21972 4068 21984
rect 4120 22012 4126 22024
rect 6656 22012 6684 22043
rect 7282 22012 7288 22024
rect 4120 21984 6684 22012
rect 7243 21984 7288 22012
rect 4120 21972 4126 21984
rect 7282 21972 7288 21984
rect 7340 21972 7346 22024
rect 7668 22012 7696 22043
rect 8570 22040 8576 22092
rect 8628 22080 8634 22092
rect 9490 22080 9496 22092
rect 8628 22052 8721 22080
rect 9451 22052 9496 22080
rect 8628 22040 8634 22052
rect 9490 22040 9496 22052
rect 9548 22040 9554 22092
rect 9677 22083 9735 22089
rect 9677 22049 9689 22083
rect 9723 22080 9735 22083
rect 9876 22080 9904 22120
rect 10318 22108 10324 22120
rect 10376 22108 10382 22160
rect 14001 22151 14059 22157
rect 14001 22148 14013 22151
rect 12820 22120 14013 22148
rect 10042 22080 10048 22092
rect 9723 22052 9904 22080
rect 10003 22052 10048 22080
rect 9723 22049 9735 22052
rect 9677 22043 9735 22049
rect 8588 22012 8616 22040
rect 9692 22012 9720 22043
rect 10042 22040 10048 22052
rect 10100 22040 10106 22092
rect 10410 22080 10416 22092
rect 10371 22052 10416 22080
rect 10410 22040 10416 22052
rect 10468 22040 10474 22092
rect 12618 22040 12624 22092
rect 12676 22080 12682 22092
rect 12820 22080 12848 22120
rect 14001 22117 14013 22120
rect 14047 22117 14059 22151
rect 15102 22148 15108 22160
rect 14001 22111 14059 22117
rect 14108 22120 15108 22148
rect 14108 22089 14136 22120
rect 15102 22108 15108 22120
rect 15160 22148 15166 22160
rect 15488 22157 15516 22188
rect 17494 22176 17500 22188
rect 17552 22176 17558 22228
rect 19613 22219 19671 22225
rect 19613 22185 19625 22219
rect 19659 22216 19671 22219
rect 23106 22216 23112 22228
rect 19659 22188 23112 22216
rect 19659 22185 19671 22188
rect 19613 22179 19671 22185
rect 23106 22176 23112 22188
rect 23164 22176 23170 22228
rect 23382 22176 23388 22228
rect 23440 22216 23446 22228
rect 24121 22219 24179 22225
rect 24121 22216 24133 22219
rect 23440 22188 24133 22216
rect 23440 22176 23446 22188
rect 24121 22185 24133 22188
rect 24167 22185 24179 22219
rect 26786 22216 26792 22228
rect 26747 22188 26792 22216
rect 24121 22179 24179 22185
rect 26786 22176 26792 22188
rect 26844 22176 26850 22228
rect 28166 22176 28172 22228
rect 28224 22216 28230 22228
rect 28353 22219 28411 22225
rect 28353 22216 28365 22219
rect 28224 22188 28365 22216
rect 28224 22176 28230 22188
rect 28353 22185 28365 22188
rect 28399 22185 28411 22219
rect 28353 22179 28411 22185
rect 30101 22219 30159 22225
rect 30101 22185 30113 22219
rect 30147 22216 30159 22219
rect 30374 22216 30380 22228
rect 30147 22188 30380 22216
rect 30147 22185 30159 22188
rect 30101 22179 30159 22185
rect 30374 22176 30380 22188
rect 30432 22176 30438 22228
rect 33502 22176 33508 22228
rect 33560 22216 33566 22228
rect 33560 22188 34560 22216
rect 33560 22176 33566 22188
rect 15473 22151 15531 22157
rect 15160 22120 15424 22148
rect 15160 22108 15166 22120
rect 12676 22052 12848 22080
rect 14093 22083 14151 22089
rect 12676 22040 12682 22052
rect 14093 22049 14105 22083
rect 14139 22080 14151 22083
rect 15396 22080 15424 22120
rect 15473 22117 15485 22151
rect 15519 22117 15531 22151
rect 15473 22111 15531 22117
rect 19797 22151 19855 22157
rect 19797 22117 19809 22151
rect 19843 22148 19855 22151
rect 19978 22148 19984 22160
rect 19843 22120 19984 22148
rect 19843 22117 19855 22120
rect 19797 22111 19855 22117
rect 19978 22108 19984 22120
rect 20036 22108 20042 22160
rect 20070 22108 20076 22160
rect 20128 22148 20134 22160
rect 20165 22151 20223 22157
rect 20165 22148 20177 22151
rect 20128 22120 20177 22148
rect 20128 22108 20134 22120
rect 20165 22117 20177 22120
rect 20211 22117 20223 22151
rect 20165 22111 20223 22117
rect 24486 22108 24492 22160
rect 24544 22148 24550 22160
rect 29546 22148 29552 22160
rect 24544 22120 25728 22148
rect 24544 22108 24550 22120
rect 15565 22083 15623 22089
rect 15565 22080 15577 22083
rect 14139 22052 14173 22080
rect 15396 22052 15577 22080
rect 14139 22049 14151 22052
rect 14093 22043 14151 22049
rect 15565 22049 15577 22052
rect 15611 22080 15623 22083
rect 16577 22083 16635 22089
rect 16577 22080 16589 22083
rect 15611 22052 16589 22080
rect 15611 22049 15623 22052
rect 15565 22043 15623 22049
rect 16577 22049 16589 22052
rect 16623 22049 16635 22083
rect 16577 22043 16635 22049
rect 16945 22083 17003 22089
rect 16945 22049 16957 22083
rect 16991 22049 17003 22083
rect 16945 22043 17003 22049
rect 10594 22012 10600 22024
rect 7668 21984 8616 22012
rect 8772 21984 9720 22012
rect 10555 21984 10600 22012
rect 2314 21904 2320 21956
rect 2372 21944 2378 21956
rect 2501 21947 2559 21953
rect 2501 21944 2513 21947
rect 2372 21916 2513 21944
rect 2372 21904 2378 21916
rect 2501 21913 2513 21916
rect 2547 21913 2559 21947
rect 4154 21944 4160 21956
rect 4115 21916 4160 21944
rect 2501 21907 2559 21913
rect 4154 21904 4160 21916
rect 4212 21904 4218 21956
rect 8772 21953 8800 21984
rect 10594 21972 10600 21984
rect 10652 21972 10658 22024
rect 11701 22015 11759 22021
rect 11701 21981 11713 22015
rect 11747 21981 11759 22015
rect 11701 21975 11759 21981
rect 11977 22015 12035 22021
rect 11977 21981 11989 22015
rect 12023 22012 12035 22015
rect 12710 22012 12716 22024
rect 12023 21984 12716 22012
rect 12023 21981 12035 21984
rect 11977 21975 12035 21981
rect 8757 21947 8815 21953
rect 8757 21913 8769 21947
rect 8803 21913 8815 21947
rect 8757 21907 8815 21913
rect 9766 21904 9772 21956
rect 9824 21944 9830 21956
rect 11716 21944 11744 21975
rect 12710 21972 12716 21984
rect 12768 21972 12774 22024
rect 16960 22012 16988 22043
rect 17034 22040 17040 22092
rect 17092 22080 17098 22092
rect 17773 22083 17831 22089
rect 17773 22080 17785 22083
rect 17092 22052 17785 22080
rect 17092 22040 17098 22052
rect 17773 22049 17785 22052
rect 17819 22049 17831 22083
rect 17773 22043 17831 22049
rect 18233 22083 18291 22089
rect 18233 22049 18245 22083
rect 18279 22080 18291 22083
rect 18874 22080 18880 22092
rect 18279 22052 18880 22080
rect 18279 22049 18291 22052
rect 18233 22043 18291 22049
rect 18874 22040 18880 22052
rect 18932 22040 18938 22092
rect 19058 22080 19064 22092
rect 19019 22052 19064 22080
rect 19058 22040 19064 22052
rect 19116 22040 19122 22092
rect 19702 22080 19708 22092
rect 19663 22052 19708 22080
rect 19702 22040 19708 22052
rect 19760 22040 19766 22092
rect 20901 22083 20959 22089
rect 20901 22049 20913 22083
rect 20947 22080 20959 22083
rect 21726 22080 21732 22092
rect 20947 22052 21732 22080
rect 20947 22049 20959 22052
rect 20901 22043 20959 22049
rect 21726 22040 21732 22052
rect 21784 22040 21790 22092
rect 21818 22040 21824 22092
rect 21876 22080 21882 22092
rect 22005 22083 22063 22089
rect 22005 22080 22017 22083
rect 21876 22052 22017 22080
rect 21876 22040 21882 22052
rect 22005 22049 22017 22052
rect 22051 22049 22063 22083
rect 22005 22043 22063 22049
rect 22186 22040 22192 22092
rect 22244 22080 22250 22092
rect 22373 22083 22431 22089
rect 22373 22080 22385 22083
rect 22244 22052 22385 22080
rect 22244 22040 22250 22052
rect 22373 22049 22385 22052
rect 22419 22049 22431 22083
rect 22738 22080 22744 22092
rect 22699 22052 22744 22080
rect 22373 22043 22431 22049
rect 22738 22040 22744 22052
rect 22796 22040 22802 22092
rect 23382 22080 23388 22092
rect 23343 22052 23388 22080
rect 23382 22040 23388 22052
rect 23440 22040 23446 22092
rect 23937 22083 23995 22089
rect 23937 22049 23949 22083
rect 23983 22049 23995 22083
rect 25406 22080 25412 22092
rect 25367 22052 25412 22080
rect 23937 22043 23995 22049
rect 16960 21984 17080 22012
rect 9824 21916 11744 21944
rect 13817 21947 13875 21953
rect 9824 21904 9830 21916
rect 13817 21913 13829 21947
rect 13863 21944 13875 21947
rect 15010 21944 15016 21956
rect 13863 21916 15016 21944
rect 13863 21913 13875 21916
rect 13817 21907 13875 21913
rect 15010 21904 15016 21916
rect 15068 21944 15074 21956
rect 15289 21947 15347 21953
rect 15289 21944 15301 21947
rect 15068 21916 15301 21944
rect 15068 21904 15074 21916
rect 15289 21913 15301 21916
rect 15335 21913 15347 21947
rect 17052 21944 17080 21984
rect 17218 21972 17224 22024
rect 17276 22012 17282 22024
rect 19429 22015 19487 22021
rect 19429 22012 19441 22015
rect 17276 21984 19441 22012
rect 17276 21972 17282 21984
rect 19429 21981 19441 21984
rect 19475 21981 19487 22015
rect 23952 22012 23980 22043
rect 25406 22040 25412 22052
rect 25464 22040 25470 22092
rect 25700 22089 25728 22120
rect 29012 22120 29552 22148
rect 25685 22083 25743 22089
rect 25685 22049 25697 22083
rect 25731 22049 25743 22083
rect 26878 22080 26884 22092
rect 26839 22052 26884 22080
rect 25685 22043 25743 22049
rect 26878 22040 26884 22052
rect 26936 22040 26942 22092
rect 27338 22080 27344 22092
rect 27299 22052 27344 22080
rect 27338 22040 27344 22052
rect 27396 22040 27402 22092
rect 27522 22080 27528 22092
rect 27483 22052 27528 22080
rect 27522 22040 27528 22052
rect 27580 22040 27586 22092
rect 28537 22083 28595 22089
rect 28537 22049 28549 22083
rect 28583 22080 28595 22083
rect 29012 22080 29040 22120
rect 29546 22108 29552 22120
rect 29604 22108 29610 22160
rect 34238 22148 34244 22160
rect 30024 22120 30604 22148
rect 28583 22052 29040 22080
rect 29089 22083 29147 22089
rect 28583 22049 28595 22052
rect 28537 22043 28595 22049
rect 29089 22049 29101 22083
rect 29135 22049 29147 22083
rect 29089 22043 29147 22049
rect 24394 22012 24400 22024
rect 23952 21984 24400 22012
rect 19429 21975 19487 21981
rect 17770 21944 17776 21956
rect 17052 21916 17776 21944
rect 15289 21907 15347 21913
rect 17770 21904 17776 21916
rect 17828 21904 17834 21956
rect 18782 21904 18788 21956
rect 18840 21944 18846 21956
rect 18877 21947 18935 21953
rect 18877 21944 18889 21947
rect 18840 21916 18889 21944
rect 18840 21904 18846 21916
rect 18877 21913 18889 21916
rect 18923 21913 18935 21947
rect 19444 21944 19472 21975
rect 24394 21972 24400 21984
rect 24452 21972 24458 22024
rect 24946 22012 24952 22024
rect 24907 21984 24952 22012
rect 24946 21972 24952 21984
rect 25004 21972 25010 22024
rect 25961 22015 26019 22021
rect 25961 21981 25973 22015
rect 26007 22012 26019 22015
rect 26970 22012 26976 22024
rect 26007 21984 26976 22012
rect 26007 21981 26019 21984
rect 25961 21975 26019 21981
rect 26970 21972 26976 21984
rect 27028 21972 27034 22024
rect 27982 22012 27988 22024
rect 27080 21984 27988 22012
rect 21085 21947 21143 21953
rect 21085 21944 21097 21947
rect 19444 21916 21097 21944
rect 18877 21907 18935 21913
rect 21085 21913 21097 21916
rect 21131 21913 21143 21947
rect 21085 21907 21143 21913
rect 23385 21947 23443 21953
rect 23385 21913 23397 21947
rect 23431 21944 23443 21947
rect 27080 21944 27108 21984
rect 27982 21972 27988 21984
rect 28040 21972 28046 22024
rect 28994 22012 29000 22024
rect 28955 21984 29000 22012
rect 28994 21972 29000 21984
rect 29052 21972 29058 22024
rect 29104 22012 29132 22043
rect 29362 22040 29368 22092
rect 29420 22080 29426 22092
rect 29825 22083 29883 22089
rect 29825 22080 29837 22083
rect 29420 22052 29837 22080
rect 29420 22040 29426 22052
rect 29825 22049 29837 22052
rect 29871 22049 29883 22083
rect 29825 22043 29883 22049
rect 30024 22012 30052 22120
rect 30576 22080 30604 22120
rect 33796 22120 34244 22148
rect 30650 22080 30656 22092
rect 30576 22052 30656 22080
rect 30650 22040 30656 22052
rect 30708 22040 30714 22092
rect 30834 22080 30840 22092
rect 30795 22052 30840 22080
rect 30834 22040 30840 22052
rect 30892 22040 30898 22092
rect 31202 22040 31208 22092
rect 31260 22080 31266 22092
rect 31389 22083 31447 22089
rect 31389 22080 31401 22083
rect 31260 22052 31401 22080
rect 31260 22040 31266 22052
rect 31389 22049 31401 22052
rect 31435 22049 31447 22083
rect 32122 22080 32128 22092
rect 32083 22052 32128 22080
rect 31389 22043 31447 22049
rect 29104 21984 30052 22012
rect 23431 21916 27108 21944
rect 31404 21944 31432 22043
rect 32122 22040 32128 22052
rect 32180 22040 32186 22092
rect 32674 22080 32680 22092
rect 32635 22052 32680 22080
rect 32674 22040 32680 22052
rect 32732 22040 32738 22092
rect 33137 22083 33195 22089
rect 33137 22049 33149 22083
rect 33183 22049 33195 22083
rect 33318 22080 33324 22092
rect 33279 22052 33324 22080
rect 33137 22043 33195 22049
rect 31846 21972 31852 22024
rect 31904 22012 31910 22024
rect 32217 22015 32275 22021
rect 32217 22012 32229 22015
rect 31904 21984 32229 22012
rect 31904 21972 31910 21984
rect 32217 21981 32229 21984
rect 32263 21981 32275 22015
rect 33152 22012 33180 22043
rect 33318 22040 33324 22052
rect 33376 22040 33382 22092
rect 33796 22089 33824 22120
rect 34238 22108 34244 22120
rect 34296 22108 34302 22160
rect 34532 22089 34560 22188
rect 36633 22151 36691 22157
rect 36633 22117 36645 22151
rect 36679 22148 36691 22151
rect 37274 22148 37280 22160
rect 36679 22120 37280 22148
rect 36679 22117 36691 22120
rect 36633 22111 36691 22117
rect 37274 22108 37280 22120
rect 37332 22108 37338 22160
rect 33781 22083 33839 22089
rect 33781 22049 33793 22083
rect 33827 22049 33839 22083
rect 33781 22043 33839 22049
rect 34517 22083 34575 22089
rect 34517 22049 34529 22083
rect 34563 22049 34575 22083
rect 35069 22083 35127 22089
rect 35069 22080 35081 22083
rect 34517 22043 34575 22049
rect 34624 22052 35081 22080
rect 33336 22012 33364 22040
rect 34624 22012 34652 22052
rect 35069 22049 35081 22052
rect 35115 22049 35127 22083
rect 35069 22043 35127 22049
rect 35529 22083 35587 22089
rect 35529 22049 35541 22083
rect 35575 22049 35587 22083
rect 35802 22080 35808 22092
rect 35763 22052 35808 22080
rect 35529 22043 35587 22049
rect 34790 22012 34796 22024
rect 33152 21984 33272 22012
rect 33336 21984 34652 22012
rect 34751 21984 34796 22012
rect 32217 21975 32275 21981
rect 33244 21956 33272 21984
rect 34790 21972 34796 21984
rect 34848 21972 34854 22024
rect 35544 22012 35572 22043
rect 35802 22040 35808 22052
rect 35860 22040 35866 22092
rect 36725 22083 36783 22089
rect 36725 22049 36737 22083
rect 36771 22080 36783 22083
rect 37642 22080 37648 22092
rect 36771 22052 37648 22080
rect 36771 22049 36783 22052
rect 36725 22043 36783 22049
rect 37642 22040 37648 22052
rect 37700 22040 37706 22092
rect 37737 22083 37795 22089
rect 37737 22049 37749 22083
rect 37783 22049 37795 22083
rect 37737 22043 37795 22049
rect 36446 22012 36452 22024
rect 35544 21984 36452 22012
rect 36446 21972 36452 21984
rect 36504 21972 36510 22024
rect 33134 21944 33140 21956
rect 31404 21916 33140 21944
rect 23431 21913 23443 21916
rect 23385 21907 23443 21913
rect 33134 21904 33140 21916
rect 33192 21904 33198 21956
rect 33226 21904 33232 21956
rect 33284 21944 33290 21956
rect 34422 21944 34428 21956
rect 33284 21916 34428 21944
rect 33284 21904 33290 21916
rect 34422 21904 34428 21916
rect 34480 21904 34486 21956
rect 35526 21904 35532 21956
rect 35584 21944 35590 21956
rect 37752 21944 37780 22043
rect 35584 21916 37780 21944
rect 35584 21904 35590 21916
rect 1857 21879 1915 21885
rect 1857 21845 1869 21879
rect 1903 21876 1915 21879
rect 3142 21876 3148 21888
rect 1903 21848 3148 21876
rect 1903 21845 1915 21848
rect 1857 21839 1915 21845
rect 3142 21836 3148 21848
rect 3200 21876 3206 21888
rect 4706 21876 4712 21888
rect 3200 21848 4712 21876
rect 3200 21836 3206 21848
rect 4706 21836 4712 21848
rect 4764 21836 4770 21888
rect 7650 21836 7656 21888
rect 7708 21876 7714 21888
rect 9309 21879 9367 21885
rect 9309 21876 9321 21879
rect 7708 21848 9321 21876
rect 7708 21836 7714 21848
rect 9309 21845 9321 21848
rect 9355 21845 9367 21879
rect 9309 21839 9367 21845
rect 13906 21836 13912 21888
rect 13964 21876 13970 21888
rect 14277 21879 14335 21885
rect 14277 21876 14289 21879
rect 13964 21848 14289 21876
rect 13964 21836 13970 21848
rect 14277 21845 14289 21848
rect 14323 21845 14335 21879
rect 14277 21839 14335 21845
rect 15378 21836 15384 21888
rect 15436 21876 15442 21888
rect 15749 21879 15807 21885
rect 15749 21876 15761 21879
rect 15436 21848 15761 21876
rect 15436 21836 15442 21848
rect 15749 21845 15761 21848
rect 15795 21845 15807 21879
rect 15749 21839 15807 21845
rect 31481 21879 31539 21885
rect 31481 21845 31493 21879
rect 31527 21876 31539 21879
rect 32674 21876 32680 21888
rect 31527 21848 32680 21876
rect 31527 21845 31539 21848
rect 31481 21839 31539 21845
rect 32674 21836 32680 21848
rect 32732 21836 32738 21888
rect 33686 21836 33692 21888
rect 33744 21876 33750 21888
rect 34238 21876 34244 21888
rect 33744 21848 34244 21876
rect 33744 21836 33750 21848
rect 34238 21836 34244 21848
rect 34296 21876 34302 21888
rect 36449 21879 36507 21885
rect 36449 21876 36461 21879
rect 34296 21848 36461 21876
rect 34296 21836 34302 21848
rect 36449 21845 36461 21848
rect 36495 21845 36507 21879
rect 36449 21839 36507 21845
rect 36722 21836 36728 21888
rect 36780 21876 36786 21888
rect 36909 21879 36967 21885
rect 36909 21876 36921 21879
rect 36780 21848 36921 21876
rect 36780 21836 36786 21848
rect 36909 21845 36921 21848
rect 36955 21845 36967 21879
rect 36909 21839 36967 21845
rect 36998 21836 37004 21888
rect 37056 21876 37062 21888
rect 37829 21879 37887 21885
rect 37829 21876 37841 21879
rect 37056 21848 37841 21876
rect 37056 21836 37062 21848
rect 37829 21845 37841 21848
rect 37875 21845 37887 21879
rect 37829 21839 37887 21845
rect 1104 21786 38824 21808
rect 1104 21734 4246 21786
rect 4298 21734 4310 21786
rect 4362 21734 4374 21786
rect 4426 21734 4438 21786
rect 4490 21734 34966 21786
rect 35018 21734 35030 21786
rect 35082 21734 35094 21786
rect 35146 21734 35158 21786
rect 35210 21734 38824 21786
rect 1104 21712 38824 21734
rect 7742 21632 7748 21684
rect 7800 21672 7806 21684
rect 8481 21675 8539 21681
rect 8481 21672 8493 21675
rect 7800 21644 8493 21672
rect 7800 21632 7806 21644
rect 8481 21641 8493 21644
rect 8527 21641 8539 21675
rect 8481 21635 8539 21641
rect 8570 21632 8576 21684
rect 8628 21672 8634 21684
rect 17034 21672 17040 21684
rect 8628 21644 17040 21672
rect 8628 21632 8634 21644
rect 17034 21632 17040 21644
rect 17092 21632 17098 21684
rect 17586 21672 17592 21684
rect 17547 21644 17592 21672
rect 17586 21632 17592 21644
rect 17644 21632 17650 21684
rect 20162 21632 20168 21684
rect 20220 21632 20226 21684
rect 21634 21672 21640 21684
rect 21595 21644 21640 21672
rect 21634 21632 21640 21644
rect 21692 21632 21698 21684
rect 21726 21632 21732 21684
rect 21784 21672 21790 21684
rect 23937 21675 23995 21681
rect 23937 21672 23949 21675
rect 21784 21644 23949 21672
rect 21784 21632 21790 21644
rect 23937 21641 23949 21644
rect 23983 21641 23995 21675
rect 28626 21672 28632 21684
rect 28587 21644 28632 21672
rect 23937 21635 23995 21641
rect 28626 21632 28632 21644
rect 28684 21632 28690 21684
rect 30558 21632 30564 21684
rect 30616 21672 30622 21684
rect 32490 21672 32496 21684
rect 30616 21644 32496 21672
rect 30616 21632 30622 21644
rect 32490 21632 32496 21644
rect 32548 21632 32554 21684
rect 32582 21632 32588 21684
rect 32640 21672 32646 21684
rect 33965 21675 34023 21681
rect 33965 21672 33977 21675
rect 32640 21644 33977 21672
rect 32640 21632 32646 21644
rect 33965 21641 33977 21644
rect 34011 21641 34023 21675
rect 33965 21635 34023 21641
rect 34422 21632 34428 21684
rect 34480 21672 34486 21684
rect 36998 21672 37004 21684
rect 34480 21644 37004 21672
rect 34480 21632 34486 21644
rect 36998 21632 37004 21644
rect 37056 21632 37062 21684
rect 1762 21564 1768 21616
rect 1820 21604 1826 21616
rect 1820 21576 5120 21604
rect 1820 21564 1826 21576
rect 1854 21496 1860 21548
rect 1912 21536 1918 21548
rect 2225 21539 2283 21545
rect 2225 21536 2237 21539
rect 1912 21508 2237 21536
rect 1912 21496 1918 21508
rect 2225 21505 2237 21508
rect 2271 21505 2283 21539
rect 2958 21536 2964 21548
rect 2225 21499 2283 21505
rect 2792 21508 2964 21536
rect 1486 21468 1492 21480
rect 1447 21440 1492 21468
rect 1486 21428 1492 21440
rect 1544 21428 1550 21480
rect 2792 21477 2820 21508
rect 2958 21496 2964 21508
rect 3016 21496 3022 21548
rect 5092 21536 5120 21576
rect 9398 21564 9404 21616
rect 9456 21564 9462 21616
rect 11517 21607 11575 21613
rect 11517 21573 11529 21607
rect 11563 21604 11575 21607
rect 12526 21604 12532 21616
rect 11563 21576 12532 21604
rect 11563 21573 11575 21576
rect 11517 21567 11575 21573
rect 12526 21564 12532 21576
rect 12584 21564 12590 21616
rect 15562 21564 15568 21616
rect 15620 21604 15626 21616
rect 16022 21604 16028 21616
rect 15620 21576 16028 21604
rect 15620 21564 15626 21576
rect 16022 21564 16028 21576
rect 16080 21604 16086 21616
rect 16482 21604 16488 21616
rect 16080 21576 16488 21604
rect 16080 21564 16086 21576
rect 16482 21564 16488 21576
rect 16540 21564 16546 21616
rect 19150 21604 19156 21616
rect 17328 21576 19156 21604
rect 6178 21536 6184 21548
rect 5092 21508 6184 21536
rect 2409 21471 2467 21477
rect 2409 21437 2421 21471
rect 2455 21437 2467 21471
rect 2409 21431 2467 21437
rect 2777 21471 2835 21477
rect 2777 21437 2789 21471
rect 2823 21437 2835 21471
rect 3142 21468 3148 21480
rect 3103 21440 3148 21468
rect 2777 21431 2835 21437
rect 2424 21400 2452 21431
rect 3142 21428 3148 21440
rect 3200 21428 3206 21480
rect 3418 21468 3424 21480
rect 3379 21440 3424 21468
rect 3418 21428 3424 21440
rect 3476 21428 3482 21480
rect 4798 21428 4804 21480
rect 4856 21468 4862 21480
rect 5092 21477 5120 21508
rect 6178 21496 6184 21508
rect 6236 21496 6242 21548
rect 9217 21539 9275 21545
rect 9217 21505 9229 21539
rect 9263 21536 9275 21539
rect 9416 21536 9444 21564
rect 9674 21536 9680 21548
rect 9263 21508 9444 21536
rect 9508 21508 9680 21536
rect 9263 21505 9275 21508
rect 9217 21499 9275 21505
rect 4893 21471 4951 21477
rect 4893 21468 4905 21471
rect 4856 21440 4905 21468
rect 4856 21428 4862 21440
rect 4893 21437 4905 21440
rect 4939 21437 4951 21471
rect 4893 21431 4951 21437
rect 5077 21471 5135 21477
rect 5077 21437 5089 21471
rect 5123 21437 5135 21471
rect 5077 21431 5135 21437
rect 5169 21471 5227 21477
rect 5169 21437 5181 21471
rect 5215 21437 5227 21471
rect 5169 21431 5227 21437
rect 5445 21471 5503 21477
rect 5445 21437 5457 21471
rect 5491 21468 5503 21471
rect 5534 21468 5540 21480
rect 5491 21440 5540 21468
rect 5491 21437 5503 21440
rect 5445 21431 5503 21437
rect 4062 21400 4068 21412
rect 2424 21372 4068 21400
rect 4062 21360 4068 21372
rect 4120 21360 4126 21412
rect 4706 21360 4712 21412
rect 4764 21400 4770 21412
rect 5184 21400 5212 21431
rect 5534 21428 5540 21440
rect 5592 21428 5598 21480
rect 5813 21471 5871 21477
rect 5813 21437 5825 21471
rect 5859 21437 5871 21471
rect 5813 21431 5871 21437
rect 7377 21471 7435 21477
rect 7377 21437 7389 21471
rect 7423 21437 7435 21471
rect 7377 21431 7435 21437
rect 8389 21471 8447 21477
rect 8389 21437 8401 21471
rect 8435 21468 8447 21471
rect 9508 21468 9536 21508
rect 9674 21496 9680 21508
rect 9732 21496 9738 21548
rect 10137 21539 10195 21545
rect 10137 21505 10149 21539
rect 10183 21536 10195 21539
rect 16390 21536 16396 21548
rect 10183 21508 12480 21536
rect 16351 21508 16396 21536
rect 10183 21505 10195 21508
rect 10137 21499 10195 21505
rect 8435 21440 9536 21468
rect 9585 21471 9643 21477
rect 8435 21437 8447 21440
rect 8389 21431 8447 21437
rect 9585 21437 9597 21471
rect 9631 21437 9643 21471
rect 9858 21468 9864 21480
rect 9819 21440 9864 21468
rect 9585 21431 9643 21437
rect 4764 21372 5212 21400
rect 4764 21360 4770 21372
rect 1578 21332 1584 21344
rect 1539 21304 1584 21332
rect 1578 21292 1584 21304
rect 1636 21292 1642 21344
rect 4433 21335 4491 21341
rect 4433 21301 4445 21335
rect 4479 21332 4491 21335
rect 4614 21332 4620 21344
rect 4479 21304 4620 21332
rect 4479 21301 4491 21304
rect 4433 21295 4491 21301
rect 4614 21292 4620 21304
rect 4672 21292 4678 21344
rect 5258 21292 5264 21344
rect 5316 21332 5322 21344
rect 5828 21332 5856 21431
rect 7392 21400 7420 21431
rect 8570 21400 8576 21412
rect 7392 21372 8576 21400
rect 8570 21360 8576 21372
rect 8628 21360 8634 21412
rect 9600 21400 9628 21431
rect 9858 21428 9864 21440
rect 9916 21428 9922 21480
rect 10594 21468 10600 21480
rect 10555 21440 10600 21468
rect 10594 21428 10600 21440
rect 10652 21428 10658 21480
rect 11330 21468 11336 21480
rect 11291 21440 11336 21468
rect 11330 21428 11336 21440
rect 11388 21428 11394 21480
rect 12452 21477 12480 21508
rect 16390 21496 16396 21508
rect 16448 21496 16454 21548
rect 17328 21545 17356 21576
rect 19150 21564 19156 21576
rect 19208 21604 19214 21616
rect 20180 21604 20208 21632
rect 19208 21576 20208 21604
rect 19208 21564 19214 21576
rect 22278 21564 22284 21616
rect 22336 21604 22342 21616
rect 23201 21607 23259 21613
rect 23201 21604 23213 21607
rect 22336 21576 23213 21604
rect 22336 21564 22342 21576
rect 23201 21573 23213 21576
rect 23247 21573 23259 21607
rect 23201 21567 23259 21573
rect 26881 21607 26939 21613
rect 26881 21573 26893 21607
rect 26927 21573 26939 21607
rect 26881 21567 26939 21573
rect 17313 21539 17371 21545
rect 17313 21505 17325 21539
rect 17359 21505 17371 21539
rect 19334 21536 19340 21548
rect 17313 21499 17371 21505
rect 18616 21508 19340 21536
rect 12437 21471 12495 21477
rect 12437 21437 12449 21471
rect 12483 21437 12495 21471
rect 12437 21431 12495 21437
rect 13725 21471 13783 21477
rect 13725 21437 13737 21471
rect 13771 21468 13783 21471
rect 13814 21468 13820 21480
rect 13771 21440 13820 21468
rect 13771 21437 13783 21440
rect 13725 21431 13783 21437
rect 13814 21428 13820 21440
rect 13872 21428 13878 21480
rect 13998 21468 14004 21480
rect 13959 21440 14004 21468
rect 13998 21428 14004 21440
rect 14056 21428 14062 21480
rect 14185 21471 14243 21477
rect 14185 21437 14197 21471
rect 14231 21437 14243 21471
rect 14185 21431 14243 21437
rect 14645 21471 14703 21477
rect 14645 21437 14657 21471
rect 14691 21468 14703 21471
rect 15378 21468 15384 21480
rect 14691 21440 15384 21468
rect 14691 21437 14703 21440
rect 14645 21431 14703 21437
rect 10689 21403 10747 21409
rect 10689 21400 10701 21403
rect 9600 21372 10701 21400
rect 10689 21369 10701 21372
rect 10735 21369 10747 21403
rect 10689 21363 10747 21369
rect 13173 21403 13231 21409
rect 13173 21369 13185 21403
rect 13219 21400 13231 21403
rect 14090 21400 14096 21412
rect 13219 21372 14096 21400
rect 13219 21369 13231 21372
rect 13173 21363 13231 21369
rect 14090 21360 14096 21372
rect 14148 21360 14154 21412
rect 7561 21335 7619 21341
rect 7561 21332 7573 21335
rect 5316 21304 7573 21332
rect 5316 21292 5322 21304
rect 7561 21301 7573 21304
rect 7607 21332 7619 21335
rect 8110 21332 8116 21344
rect 7607 21304 8116 21332
rect 7607 21301 7619 21304
rect 7561 21295 7619 21301
rect 8110 21292 8116 21304
rect 8168 21292 8174 21344
rect 12526 21332 12532 21344
rect 12487 21304 12532 21332
rect 12526 21292 12532 21304
rect 12584 21292 12590 21344
rect 13722 21292 13728 21344
rect 13780 21332 13786 21344
rect 14200 21332 14228 21431
rect 15378 21428 15384 21440
rect 15436 21428 15442 21480
rect 15473 21471 15531 21477
rect 15473 21437 15485 21471
rect 15519 21468 15531 21471
rect 15562 21468 15568 21480
rect 15519 21440 15568 21468
rect 15519 21437 15531 21440
rect 15473 21431 15531 21437
rect 15562 21428 15568 21440
rect 15620 21428 15626 21480
rect 15749 21471 15807 21477
rect 15749 21437 15761 21471
rect 15795 21437 15807 21471
rect 16114 21468 16120 21480
rect 16075 21440 16120 21468
rect 15749 21431 15807 21437
rect 13780 21304 14228 21332
rect 13780 21292 13786 21304
rect 14366 21292 14372 21344
rect 14424 21332 14430 21344
rect 14737 21335 14795 21341
rect 14737 21332 14749 21335
rect 14424 21304 14749 21332
rect 14424 21292 14430 21304
rect 14737 21301 14749 21304
rect 14783 21301 14795 21335
rect 15764 21332 15792 21431
rect 16114 21428 16120 21440
rect 16172 21428 16178 21480
rect 16853 21471 16911 21477
rect 16853 21437 16865 21471
rect 16899 21468 16911 21471
rect 17034 21468 17040 21480
rect 16899 21440 17040 21468
rect 16899 21437 16911 21440
rect 16853 21431 16911 21437
rect 17034 21428 17040 21440
rect 17092 21428 17098 21480
rect 17405 21471 17463 21477
rect 17405 21437 17417 21471
rect 17451 21468 17463 21471
rect 17954 21468 17960 21480
rect 17451 21440 17960 21468
rect 17451 21437 17463 21440
rect 17405 21431 17463 21437
rect 17954 21428 17960 21440
rect 18012 21428 18018 21480
rect 18233 21471 18291 21477
rect 18233 21437 18245 21471
rect 18279 21468 18291 21471
rect 18506 21468 18512 21480
rect 18279 21440 18512 21468
rect 18279 21437 18291 21440
rect 18233 21431 18291 21437
rect 18506 21428 18512 21440
rect 18564 21428 18570 21480
rect 18616 21477 18644 21508
rect 19334 21496 19340 21508
rect 19392 21496 19398 21548
rect 19886 21536 19892 21548
rect 19536 21508 19892 21536
rect 18601 21471 18659 21477
rect 18601 21437 18613 21471
rect 18647 21437 18659 21471
rect 18966 21468 18972 21480
rect 18927 21440 18972 21468
rect 18601 21431 18659 21437
rect 18966 21428 18972 21440
rect 19024 21428 19030 21480
rect 19536 21477 19564 21508
rect 19886 21496 19892 21508
rect 19944 21496 19950 21548
rect 23661 21539 23719 21545
rect 23661 21505 23673 21539
rect 23707 21536 23719 21539
rect 24118 21536 24124 21548
rect 23707 21508 24124 21536
rect 23707 21505 23719 21508
rect 23661 21499 23719 21505
rect 24118 21496 24124 21508
rect 24176 21496 24182 21548
rect 24949 21539 25007 21545
rect 24949 21505 24961 21539
rect 24995 21536 25007 21539
rect 26896 21536 26924 21567
rect 30374 21564 30380 21616
rect 30432 21604 30438 21616
rect 31294 21604 31300 21616
rect 30432 21576 31300 21604
rect 30432 21564 30438 21576
rect 31294 21564 31300 21576
rect 31352 21604 31358 21616
rect 32398 21604 32404 21616
rect 31352 21576 32404 21604
rect 31352 21564 31358 21576
rect 32398 21564 32404 21576
rect 32456 21564 32462 21616
rect 33226 21604 33232 21616
rect 32600 21576 33232 21604
rect 24995 21508 26924 21536
rect 24995 21505 25007 21508
rect 24949 21499 25007 21505
rect 26970 21496 26976 21548
rect 27028 21536 27034 21548
rect 27617 21539 27675 21545
rect 27617 21536 27629 21539
rect 27028 21508 27629 21536
rect 27028 21496 27034 21508
rect 27617 21505 27629 21508
rect 27663 21505 27675 21539
rect 31202 21536 31208 21548
rect 27617 21499 27675 21505
rect 29380 21508 31208 21536
rect 29380 21480 29408 21508
rect 19521 21471 19579 21477
rect 19521 21437 19533 21471
rect 19567 21437 19579 21471
rect 19794 21468 19800 21480
rect 19755 21440 19800 21468
rect 19521 21431 19579 21437
rect 19794 21428 19800 21440
rect 19852 21428 19858 21480
rect 19981 21471 20039 21477
rect 19981 21437 19993 21471
rect 20027 21437 20039 21471
rect 19981 21431 20039 21437
rect 15838 21360 15844 21412
rect 15896 21400 15902 21412
rect 19153 21403 19211 21409
rect 19153 21400 19165 21403
rect 15896 21372 19165 21400
rect 15896 21360 15902 21372
rect 19153 21369 19165 21372
rect 19199 21369 19211 21403
rect 19153 21363 19211 21369
rect 19426 21360 19432 21412
rect 19484 21400 19490 21412
rect 19996 21400 20024 21431
rect 20254 21428 20260 21480
rect 20312 21468 20318 21480
rect 20533 21471 20591 21477
rect 20533 21468 20545 21471
rect 20312 21440 20545 21468
rect 20312 21428 20318 21440
rect 20533 21437 20545 21440
rect 20579 21437 20591 21471
rect 20533 21431 20591 21437
rect 21174 21428 21180 21480
rect 21232 21468 21238 21480
rect 21818 21468 21824 21480
rect 21232 21440 21824 21468
rect 21232 21428 21238 21440
rect 21818 21428 21824 21440
rect 21876 21428 21882 21480
rect 22189 21471 22247 21477
rect 22189 21437 22201 21471
rect 22235 21468 22247 21471
rect 22278 21468 22284 21480
rect 22235 21440 22284 21468
rect 22235 21437 22247 21440
rect 22189 21431 22247 21437
rect 22278 21428 22284 21440
rect 22336 21428 22342 21480
rect 22557 21471 22615 21477
rect 22557 21437 22569 21471
rect 22603 21468 22615 21471
rect 22738 21468 22744 21480
rect 22603 21440 22744 21468
rect 22603 21437 22615 21440
rect 22557 21431 22615 21437
rect 22738 21428 22744 21440
rect 22796 21428 22802 21480
rect 23385 21471 23443 21477
rect 23385 21437 23397 21471
rect 23431 21468 23443 21471
rect 23566 21468 23572 21480
rect 23431 21440 23572 21468
rect 23431 21437 23443 21440
rect 23385 21431 23443 21437
rect 23566 21428 23572 21440
rect 23624 21428 23630 21480
rect 23753 21471 23811 21477
rect 23753 21437 23765 21471
rect 23799 21437 23811 21471
rect 23753 21431 23811 21437
rect 19484 21372 20024 21400
rect 20441 21403 20499 21409
rect 19484 21360 19490 21372
rect 20441 21369 20453 21403
rect 20487 21369 20499 21403
rect 20441 21363 20499 21369
rect 16206 21332 16212 21344
rect 15764 21304 16212 21332
rect 14737 21295 14795 21301
rect 16206 21292 16212 21304
rect 16264 21292 16270 21344
rect 16482 21292 16488 21344
rect 16540 21332 16546 21344
rect 17037 21335 17095 21341
rect 17037 21332 17049 21335
rect 16540 21304 17049 21332
rect 16540 21292 16546 21304
rect 17037 21301 17049 21304
rect 17083 21301 17095 21335
rect 20456 21332 20484 21363
rect 20530 21332 20536 21344
rect 20456 21304 20536 21332
rect 17037 21295 17095 21301
rect 20530 21292 20536 21304
rect 20588 21292 20594 21344
rect 22756 21332 22784 21428
rect 23658 21332 23664 21344
rect 22756 21304 23664 21332
rect 23658 21292 23664 21304
rect 23716 21292 23722 21344
rect 23768 21332 23796 21431
rect 24026 21428 24032 21480
rect 24084 21468 24090 21480
rect 24673 21471 24731 21477
rect 24673 21468 24685 21471
rect 24084 21440 24685 21468
rect 24084 21428 24090 21440
rect 24673 21437 24685 21440
rect 24719 21468 24731 21471
rect 26510 21468 26516 21480
rect 24719 21440 26516 21468
rect 24719 21437 24731 21440
rect 24673 21431 24731 21437
rect 26510 21428 26516 21440
rect 26568 21428 26574 21480
rect 26881 21471 26939 21477
rect 26881 21437 26893 21471
rect 26927 21437 26939 21471
rect 26881 21431 26939 21437
rect 26896 21400 26924 21431
rect 27062 21428 27068 21480
rect 27120 21468 27126 21480
rect 27341 21471 27399 21477
rect 27341 21468 27353 21471
rect 27120 21440 27353 21468
rect 27120 21428 27126 21440
rect 27341 21437 27353 21440
rect 27387 21437 27399 21471
rect 27341 21431 27399 21437
rect 28445 21471 28503 21477
rect 28445 21437 28457 21471
rect 28491 21468 28503 21471
rect 29362 21468 29368 21480
rect 28491 21440 29368 21468
rect 28491 21437 28503 21440
rect 28445 21431 28503 21437
rect 29362 21428 29368 21440
rect 29420 21428 29426 21480
rect 29549 21471 29607 21477
rect 29549 21437 29561 21471
rect 29595 21468 29607 21471
rect 29638 21468 29644 21480
rect 29595 21440 29644 21468
rect 29595 21437 29607 21440
rect 29549 21431 29607 21437
rect 29638 21428 29644 21440
rect 29696 21428 29702 21480
rect 29733 21471 29791 21477
rect 29733 21437 29745 21471
rect 29779 21437 29791 21471
rect 29733 21431 29791 21437
rect 27246 21400 27252 21412
rect 26896 21372 27252 21400
rect 27246 21360 27252 21372
rect 27304 21360 27310 21412
rect 27522 21360 27528 21412
rect 27580 21400 27586 21412
rect 29748 21400 29776 21431
rect 29914 21428 29920 21480
rect 29972 21468 29978 21480
rect 30852 21477 30880 21508
rect 31202 21496 31208 21508
rect 31260 21496 31266 21548
rect 32600 21536 32628 21576
rect 33226 21564 33232 21576
rect 33284 21564 33290 21616
rect 32766 21536 32772 21548
rect 32508 21508 32628 21536
rect 32727 21508 32772 21536
rect 30101 21471 30159 21477
rect 30101 21468 30113 21471
rect 29972 21440 30113 21468
rect 29972 21428 29978 21440
rect 30101 21437 30113 21440
rect 30147 21437 30159 21471
rect 30101 21431 30159 21437
rect 30837 21471 30895 21477
rect 30837 21437 30849 21471
rect 30883 21437 30895 21471
rect 30837 21431 30895 21437
rect 30926 21428 30932 21480
rect 30984 21468 30990 21480
rect 32508 21477 32536 21508
rect 32766 21496 32772 21508
rect 32824 21496 32830 21548
rect 33042 21536 33048 21548
rect 32876 21508 33048 21536
rect 32876 21477 32904 21508
rect 33042 21496 33048 21508
rect 33100 21496 33106 21548
rect 34330 21496 34336 21548
rect 34388 21536 34394 21548
rect 35161 21539 35219 21545
rect 35161 21536 35173 21539
rect 34388 21508 35173 21536
rect 34388 21496 34394 21508
rect 35161 21505 35173 21508
rect 35207 21505 35219 21539
rect 35161 21499 35219 21505
rect 37274 21496 37280 21548
rect 37332 21536 37338 21548
rect 37332 21508 37872 21536
rect 37332 21496 37338 21508
rect 37844 21480 37872 21508
rect 31297 21471 31355 21477
rect 31297 21468 31309 21471
rect 30984 21440 31309 21468
rect 30984 21428 30990 21440
rect 31297 21437 31309 21440
rect 31343 21437 31355 21471
rect 31297 21431 31355 21437
rect 32493 21471 32551 21477
rect 32493 21437 32505 21471
rect 32539 21437 32551 21471
rect 32493 21431 32551 21437
rect 32861 21471 32919 21477
rect 32861 21437 32873 21471
rect 32907 21437 32919 21471
rect 32861 21431 32919 21437
rect 32953 21471 33011 21477
rect 32953 21437 32965 21471
rect 32999 21437 33011 21471
rect 32953 21431 33011 21437
rect 33873 21471 33931 21477
rect 33873 21437 33885 21471
rect 33919 21468 33931 21471
rect 33962 21468 33968 21480
rect 33919 21440 33968 21468
rect 33919 21437 33931 21440
rect 33873 21431 33931 21437
rect 27580 21372 29776 21400
rect 27580 21360 27586 21372
rect 30466 21360 30472 21412
rect 30524 21400 30530 21412
rect 31570 21400 31576 21412
rect 30524 21372 31576 21400
rect 30524 21360 30530 21372
rect 31570 21360 31576 21372
rect 31628 21360 31634 21412
rect 31754 21360 31760 21412
rect 31812 21400 31818 21412
rect 32030 21400 32036 21412
rect 31812 21372 32036 21400
rect 31812 21360 31818 21372
rect 32030 21360 32036 21372
rect 32088 21360 32094 21412
rect 32214 21360 32220 21412
rect 32272 21400 32278 21412
rect 32674 21400 32680 21412
rect 32272 21372 32680 21400
rect 32272 21360 32278 21372
rect 32674 21360 32680 21372
rect 32732 21400 32738 21412
rect 32968 21400 32996 21431
rect 33962 21428 33968 21440
rect 34020 21428 34026 21480
rect 34885 21471 34943 21477
rect 34885 21437 34897 21471
rect 34931 21468 34943 21471
rect 35250 21468 35256 21480
rect 34931 21440 35256 21468
rect 34931 21437 34943 21440
rect 34885 21431 34943 21437
rect 35250 21428 35256 21440
rect 35308 21428 35314 21480
rect 36078 21468 36084 21480
rect 35820 21440 36084 21468
rect 32732 21372 32996 21400
rect 32732 21360 32738 21372
rect 24394 21332 24400 21344
rect 23768 21304 24400 21332
rect 24394 21292 24400 21304
rect 24452 21332 24458 21344
rect 26053 21335 26111 21341
rect 26053 21332 26065 21335
rect 24452 21304 26065 21332
rect 24452 21292 24458 21304
rect 26053 21301 26065 21304
rect 26099 21301 26111 21335
rect 26053 21295 26111 21301
rect 29178 21292 29184 21344
rect 29236 21332 29242 21344
rect 29365 21335 29423 21341
rect 29365 21332 29377 21335
rect 29236 21304 29377 21332
rect 29236 21292 29242 21304
rect 29365 21301 29377 21304
rect 29411 21301 29423 21335
rect 29365 21295 29423 21301
rect 31478 21292 31484 21344
rect 31536 21332 31542 21344
rect 35820 21332 35848 21440
rect 36078 21428 36084 21440
rect 36136 21468 36142 21480
rect 37001 21471 37059 21477
rect 37001 21468 37013 21471
rect 36136 21440 37013 21468
rect 36136 21428 36142 21440
rect 37001 21437 37013 21440
rect 37047 21437 37059 21471
rect 37642 21468 37648 21480
rect 37603 21440 37648 21468
rect 37001 21431 37059 21437
rect 37642 21428 37648 21440
rect 37700 21428 37706 21480
rect 37826 21468 37832 21480
rect 37787 21440 37832 21468
rect 37826 21428 37832 21440
rect 37884 21428 37890 21480
rect 31536 21304 35848 21332
rect 31536 21292 31542 21304
rect 35894 21292 35900 21344
rect 35952 21332 35958 21344
rect 36265 21335 36323 21341
rect 36265 21332 36277 21335
rect 35952 21304 36277 21332
rect 35952 21292 35958 21304
rect 36265 21301 36277 21304
rect 36311 21301 36323 21335
rect 36265 21295 36323 21301
rect 37277 21335 37335 21341
rect 37277 21301 37289 21335
rect 37323 21332 37335 21335
rect 37366 21332 37372 21344
rect 37323 21304 37372 21332
rect 37323 21301 37335 21304
rect 37277 21295 37335 21301
rect 37366 21292 37372 21304
rect 37424 21292 37430 21344
rect 1104 21242 38824 21264
rect 1104 21190 19606 21242
rect 19658 21190 19670 21242
rect 19722 21190 19734 21242
rect 19786 21190 19798 21242
rect 19850 21190 38824 21242
rect 1104 21168 38824 21190
rect 4062 21088 4068 21140
rect 4120 21128 4126 21140
rect 4249 21131 4307 21137
rect 4249 21128 4261 21131
rect 4120 21100 4261 21128
rect 4120 21088 4126 21100
rect 4249 21097 4261 21100
rect 4295 21097 4307 21131
rect 4249 21091 4307 21097
rect 8389 21131 8447 21137
rect 8389 21097 8401 21131
rect 8435 21128 8447 21131
rect 8570 21128 8576 21140
rect 8435 21100 8576 21128
rect 8435 21097 8447 21100
rect 8389 21091 8447 21097
rect 8570 21088 8576 21100
rect 8628 21088 8634 21140
rect 11330 21128 11336 21140
rect 11291 21100 11336 21128
rect 11330 21088 11336 21100
rect 11388 21088 11394 21140
rect 14642 21128 14648 21140
rect 14603 21100 14648 21128
rect 14642 21088 14648 21100
rect 14700 21088 14706 21140
rect 15378 21088 15384 21140
rect 15436 21128 15442 21140
rect 19797 21131 19855 21137
rect 19797 21128 19809 21131
rect 15436 21100 19809 21128
rect 15436 21088 15442 21100
rect 19797 21097 19809 21100
rect 19843 21128 19855 21131
rect 21450 21128 21456 21140
rect 19843 21100 21456 21128
rect 19843 21097 19855 21100
rect 19797 21091 19855 21097
rect 21450 21088 21456 21100
rect 21508 21088 21514 21140
rect 27246 21088 27252 21140
rect 27304 21128 27310 21140
rect 29270 21128 29276 21140
rect 27304 21100 29276 21128
rect 27304 21088 27310 21100
rect 29270 21088 29276 21100
rect 29328 21088 29334 21140
rect 29546 21088 29552 21140
rect 29604 21128 29610 21140
rect 30285 21131 30343 21137
rect 30285 21128 30297 21131
rect 29604 21100 30297 21128
rect 29604 21088 29610 21100
rect 30285 21097 30297 21100
rect 30331 21097 30343 21131
rect 30285 21091 30343 21097
rect 32306 21088 32312 21140
rect 32364 21128 32370 21140
rect 33042 21128 33048 21140
rect 32364 21100 33048 21128
rect 32364 21088 32370 21100
rect 33042 21088 33048 21100
rect 33100 21128 33106 21140
rect 37829 21131 37887 21137
rect 37829 21128 37841 21131
rect 33100 21100 37841 21128
rect 33100 21088 33106 21100
rect 37829 21097 37841 21100
rect 37875 21097 37887 21131
rect 37829 21091 37887 21097
rect 8202 21060 8208 21072
rect 4172 21032 5488 21060
rect 1854 20992 1860 21004
rect 1815 20964 1860 20992
rect 1854 20952 1860 20964
rect 1912 20952 1918 21004
rect 2314 20992 2320 21004
rect 2275 20964 2320 20992
rect 2314 20952 2320 20964
rect 2372 20952 2378 21004
rect 2958 20992 2964 21004
rect 2919 20964 2964 20992
rect 2958 20952 2964 20964
rect 3016 20952 3022 21004
rect 3418 20992 3424 21004
rect 3379 20964 3424 20992
rect 3418 20952 3424 20964
rect 3476 20952 3482 21004
rect 4172 21001 4200 21032
rect 4157 20995 4215 21001
rect 4157 20961 4169 20995
rect 4203 20961 4215 20995
rect 4157 20955 4215 20961
rect 5077 20995 5135 21001
rect 5077 20961 5089 20995
rect 5123 20992 5135 20995
rect 5258 20992 5264 21004
rect 5123 20964 5264 20992
rect 5123 20961 5135 20964
rect 5077 20955 5135 20961
rect 5258 20952 5264 20964
rect 5316 20952 5322 21004
rect 5460 21001 5488 21032
rect 7300 21032 8208 21060
rect 5445 20995 5503 21001
rect 5445 20961 5457 20995
rect 5491 20992 5503 20995
rect 5534 20992 5540 21004
rect 5491 20964 5540 20992
rect 5491 20961 5503 20964
rect 5445 20955 5503 20961
rect 5534 20952 5540 20964
rect 5592 20952 5598 21004
rect 5629 20995 5687 21001
rect 5629 20961 5641 20995
rect 5675 20961 5687 20995
rect 6178 20992 6184 21004
rect 6139 20964 6184 20992
rect 5629 20955 5687 20961
rect 3145 20927 3203 20933
rect 3145 20893 3157 20927
rect 3191 20924 3203 20927
rect 5644 20924 5672 20955
rect 6178 20952 6184 20964
rect 6236 20952 6242 21004
rect 6454 20952 6460 21004
rect 6512 20992 6518 21004
rect 7300 21001 7328 21032
rect 8202 21020 8208 21032
rect 8260 21020 8266 21072
rect 16758 21060 16764 21072
rect 16719 21032 16764 21060
rect 16758 21020 16764 21032
rect 16816 21020 16822 21072
rect 17034 21020 17040 21072
rect 17092 21060 17098 21072
rect 19978 21060 19984 21072
rect 17092 21032 18920 21060
rect 19939 21032 19984 21060
rect 17092 21020 17098 21032
rect 7285 20995 7343 21001
rect 7285 20992 7297 20995
rect 6512 20964 7297 20992
rect 6512 20952 6518 20964
rect 7285 20961 7297 20964
rect 7331 20961 7343 20995
rect 7285 20955 7343 20961
rect 7374 20952 7380 21004
rect 7432 20992 7438 21004
rect 8297 20995 8355 21001
rect 8297 20992 8309 20995
rect 7432 20964 7477 20992
rect 7576 20964 8309 20992
rect 7432 20952 7438 20964
rect 5902 20924 5908 20936
rect 3191 20896 5908 20924
rect 3191 20893 3203 20896
rect 3145 20887 3203 20893
rect 5902 20884 5908 20896
rect 5960 20884 5966 20936
rect 6270 20924 6276 20936
rect 6231 20896 6276 20924
rect 6270 20884 6276 20896
rect 6328 20884 6334 20936
rect 7006 20884 7012 20936
rect 7064 20924 7070 20936
rect 7576 20924 7604 20964
rect 8297 20961 8309 20964
rect 8343 20961 8355 20995
rect 8938 20992 8944 21004
rect 8899 20964 8944 20992
rect 8297 20955 8355 20961
rect 8938 20952 8944 20964
rect 8996 20952 9002 21004
rect 9766 20992 9772 21004
rect 9727 20964 9772 20992
rect 9766 20952 9772 20964
rect 9824 20952 9830 21004
rect 10045 20995 10103 21001
rect 10045 20961 10057 20995
rect 10091 20992 10103 20995
rect 12526 20992 12532 21004
rect 10091 20964 12532 20992
rect 10091 20961 10103 20964
rect 10045 20955 10103 20961
rect 12526 20952 12532 20964
rect 12584 20952 12590 21004
rect 13357 20995 13415 21001
rect 13357 20961 13369 20995
rect 13403 20961 13415 20995
rect 13357 20955 13415 20961
rect 13725 20995 13783 21001
rect 13725 20961 13737 20995
rect 13771 20992 13783 20995
rect 14458 20992 14464 21004
rect 13771 20964 14464 20992
rect 13771 20961 13783 20964
rect 13725 20955 13783 20961
rect 7064 20896 7604 20924
rect 7837 20927 7895 20933
rect 7064 20884 7070 20896
rect 7837 20893 7849 20927
rect 7883 20924 7895 20927
rect 9490 20924 9496 20936
rect 7883 20896 9496 20924
rect 7883 20893 7895 20896
rect 7837 20887 7895 20893
rect 9490 20884 9496 20896
rect 9548 20884 9554 20936
rect 12897 20927 12955 20933
rect 12897 20924 12909 20927
rect 9600 20896 12909 20924
rect 1486 20816 1492 20868
rect 1544 20856 1550 20868
rect 1673 20859 1731 20865
rect 1673 20856 1685 20859
rect 1544 20828 1685 20856
rect 1544 20816 1550 20828
rect 1673 20825 1685 20828
rect 1719 20825 1731 20859
rect 9030 20856 9036 20868
rect 8943 20828 9036 20856
rect 1673 20819 1731 20825
rect 9030 20816 9036 20828
rect 9088 20856 9094 20868
rect 9600 20856 9628 20896
rect 12897 20893 12909 20896
rect 12943 20893 12955 20927
rect 13372 20924 13400 20955
rect 14458 20952 14464 20964
rect 14516 20952 14522 21004
rect 14553 20995 14611 21001
rect 14553 20961 14565 20995
rect 14599 20992 14611 20995
rect 15194 20992 15200 21004
rect 14599 20964 15200 20992
rect 14599 20961 14611 20964
rect 14553 20955 14611 20961
rect 15194 20952 15200 20964
rect 15252 20952 15258 21004
rect 15838 20992 15844 21004
rect 15799 20964 15844 20992
rect 15838 20952 15844 20964
rect 15896 20952 15902 21004
rect 16025 20995 16083 21001
rect 16025 20961 16037 20995
rect 16071 20961 16083 20995
rect 16025 20955 16083 20961
rect 16485 20995 16543 21001
rect 16485 20961 16497 20995
rect 16531 20961 16543 20995
rect 17218 20992 17224 21004
rect 17179 20964 17224 20992
rect 16485 20955 16543 20961
rect 13814 20924 13820 20936
rect 13372 20896 13820 20924
rect 12897 20887 12955 20893
rect 13814 20884 13820 20896
rect 13872 20924 13878 20936
rect 14182 20924 14188 20936
rect 13872 20896 14188 20924
rect 13872 20884 13878 20896
rect 14182 20884 14188 20896
rect 14240 20884 14246 20936
rect 15654 20884 15660 20936
rect 15712 20924 15718 20936
rect 16040 20924 16068 20955
rect 15712 20896 16068 20924
rect 15712 20884 15718 20896
rect 9088 20828 9628 20856
rect 9088 20816 9094 20828
rect 13538 20816 13544 20868
rect 13596 20856 13602 20868
rect 13633 20859 13691 20865
rect 13633 20856 13645 20859
rect 13596 20828 13645 20856
rect 13596 20816 13602 20828
rect 13633 20825 13645 20828
rect 13679 20825 13691 20859
rect 16500 20856 16528 20955
rect 17218 20952 17224 20964
rect 17276 20952 17282 21004
rect 17770 20992 17776 21004
rect 17683 20964 17776 20992
rect 17770 20952 17776 20964
rect 17828 20992 17834 21004
rect 18414 20992 18420 21004
rect 17828 20964 18276 20992
rect 18375 20964 18420 20992
rect 17828 20952 17834 20964
rect 18141 20859 18199 20865
rect 18141 20856 18153 20859
rect 16500 20828 18153 20856
rect 13633 20819 13691 20825
rect 18141 20825 18153 20828
rect 18187 20825 18199 20859
rect 18248 20856 18276 20964
rect 18414 20952 18420 20964
rect 18472 20952 18478 21004
rect 18892 21001 18920 21032
rect 19978 21020 19984 21032
rect 20036 21020 20042 21072
rect 20346 21060 20352 21072
rect 20307 21032 20352 21060
rect 20346 21020 20352 21032
rect 20404 21020 20410 21072
rect 21358 21020 21364 21072
rect 21416 21060 21422 21072
rect 21416 21032 22140 21060
rect 21416 21020 21422 21032
rect 18877 20995 18935 21001
rect 18877 20961 18889 20995
rect 18923 20992 18935 20995
rect 19886 20992 19892 21004
rect 18923 20964 19748 20992
rect 19799 20964 19892 20992
rect 18923 20961 18935 20964
rect 18877 20955 18935 20961
rect 19426 20884 19432 20936
rect 19484 20924 19490 20936
rect 19521 20927 19579 20933
rect 19521 20924 19533 20927
rect 19484 20896 19533 20924
rect 19484 20884 19490 20896
rect 19521 20893 19533 20896
rect 19567 20924 19579 20927
rect 19613 20927 19671 20933
rect 19613 20924 19625 20927
rect 19567 20896 19625 20924
rect 19567 20893 19579 20896
rect 19521 20887 19579 20893
rect 19613 20893 19625 20896
rect 19659 20893 19671 20927
rect 19720 20924 19748 20964
rect 19886 20952 19892 20964
rect 19944 20992 19950 21004
rect 20714 20992 20720 21004
rect 19944 20964 20720 20992
rect 19944 20952 19950 20964
rect 20714 20952 20720 20964
rect 20772 20952 20778 21004
rect 21637 20995 21695 21001
rect 21637 20961 21649 20995
rect 21683 20961 21695 20995
rect 21637 20955 21695 20961
rect 20530 20924 20536 20936
rect 19720 20896 20536 20924
rect 19613 20887 19671 20893
rect 20530 20884 20536 20896
rect 20588 20884 20594 20936
rect 21652 20924 21680 20955
rect 21726 20952 21732 21004
rect 21784 20992 21790 21004
rect 22112 21001 22140 21032
rect 24302 21020 24308 21072
rect 24360 21060 24366 21072
rect 32122 21060 32128 21072
rect 24360 21032 28304 21060
rect 32083 21032 32128 21060
rect 24360 21020 24366 21032
rect 22097 20995 22155 21001
rect 21784 20964 21829 20992
rect 21784 20952 21790 20964
rect 22097 20961 22109 20995
rect 22143 20961 22155 20995
rect 22097 20955 22155 20961
rect 23017 20995 23075 21001
rect 23017 20961 23029 20995
rect 23063 20992 23075 20995
rect 24026 20992 24032 21004
rect 23063 20964 24032 20992
rect 23063 20961 23075 20964
rect 23017 20955 23075 20961
rect 24026 20952 24032 20964
rect 24084 20952 24090 21004
rect 24118 20952 24124 21004
rect 24176 20992 24182 21004
rect 25133 20995 25191 21001
rect 25133 20992 25145 20995
rect 24176 20964 25145 20992
rect 24176 20952 24182 20964
rect 25133 20961 25145 20964
rect 25179 20961 25191 20995
rect 25133 20955 25191 20961
rect 27249 20995 27307 21001
rect 27249 20961 27261 20995
rect 27295 20992 27307 20995
rect 27522 20992 27528 21004
rect 27295 20964 27528 20992
rect 27295 20961 27307 20964
rect 27249 20955 27307 20961
rect 27522 20952 27528 20964
rect 27580 20952 27586 21004
rect 28276 21001 28304 21032
rect 32122 21020 32128 21032
rect 32180 21020 32186 21072
rect 32398 21020 32404 21072
rect 32456 21060 32462 21072
rect 37550 21060 37556 21072
rect 32456 21032 32628 21060
rect 32456 21020 32462 21032
rect 27617 20995 27675 21001
rect 27617 20961 27629 20995
rect 27663 20961 27675 20995
rect 27617 20955 27675 20961
rect 27985 20995 28043 21001
rect 27985 20961 27997 20995
rect 28031 20961 28043 20995
rect 27985 20955 28043 20961
rect 28261 20995 28319 21001
rect 28261 20961 28273 20995
rect 28307 20961 28319 20995
rect 28902 20992 28908 21004
rect 28863 20964 28908 20992
rect 28261 20955 28319 20961
rect 22278 20924 22284 20936
rect 21652 20896 22284 20924
rect 22278 20884 22284 20896
rect 22336 20884 22342 20936
rect 23293 20927 23351 20933
rect 23293 20893 23305 20927
rect 23339 20924 23351 20927
rect 23474 20924 23480 20936
rect 23339 20896 23480 20924
rect 23339 20893 23351 20896
rect 23293 20887 23351 20893
rect 23474 20884 23480 20896
rect 23532 20884 23538 20936
rect 23658 20884 23664 20936
rect 23716 20924 23722 20936
rect 24397 20927 24455 20933
rect 24397 20924 24409 20927
rect 23716 20896 24409 20924
rect 23716 20884 23722 20896
rect 24397 20893 24409 20896
rect 24443 20893 24455 20927
rect 24397 20887 24455 20893
rect 20438 20856 20444 20868
rect 18248 20828 20444 20856
rect 18141 20819 18199 20825
rect 20438 20816 20444 20828
rect 20496 20816 20502 20868
rect 27632 20856 27660 20955
rect 28000 20924 28028 20955
rect 28902 20952 28908 20964
rect 28960 20952 28966 21004
rect 29178 20992 29184 21004
rect 29139 20964 29184 20992
rect 29178 20952 29184 20964
rect 29236 20952 29242 21004
rect 29270 20952 29276 21004
rect 29328 20992 29334 21004
rect 30190 20992 30196 21004
rect 29328 20964 30196 20992
rect 29328 20952 29334 20964
rect 30190 20952 30196 20964
rect 30248 20952 30254 21004
rect 31297 20995 31355 21001
rect 31297 20961 31309 20995
rect 31343 20992 31355 20995
rect 32030 20992 32036 21004
rect 31343 20964 32036 20992
rect 31343 20961 31355 20964
rect 31297 20955 31355 20961
rect 32030 20952 32036 20964
rect 32088 20952 32094 21004
rect 32600 21001 32628 21032
rect 33060 21032 34744 21060
rect 32585 20995 32643 21001
rect 32585 20961 32597 20995
rect 32631 20961 32643 20995
rect 32585 20955 32643 20961
rect 32858 20952 32864 21004
rect 32916 20992 32922 21004
rect 33060 21001 33088 21032
rect 34716 21004 34744 21032
rect 36648 21032 37556 21060
rect 36648 21004 36676 21032
rect 37550 21020 37556 21032
rect 37608 21020 37614 21072
rect 32953 20995 33011 21001
rect 32953 20992 32965 20995
rect 32916 20964 32965 20992
rect 32916 20952 32922 20964
rect 32953 20961 32965 20964
rect 32999 20961 33011 20995
rect 32953 20955 33011 20961
rect 33045 20995 33103 21001
rect 33045 20961 33057 20995
rect 33091 20961 33103 20995
rect 33870 20992 33876 21004
rect 33831 20964 33876 20992
rect 33045 20955 33103 20961
rect 33870 20952 33876 20964
rect 33928 20952 33934 21004
rect 34333 20995 34391 21001
rect 33980 20964 34284 20992
rect 31754 20924 31760 20936
rect 28000 20896 31760 20924
rect 31754 20884 31760 20896
rect 31812 20884 31818 20936
rect 32490 20884 32496 20936
rect 32548 20924 32554 20936
rect 33980 20924 34008 20964
rect 34146 20924 34152 20936
rect 32548 20896 34008 20924
rect 34107 20896 34152 20924
rect 32548 20884 32554 20896
rect 34146 20884 34152 20896
rect 34204 20884 34210 20936
rect 34256 20924 34284 20964
rect 34333 20961 34345 20995
rect 34379 20992 34391 20995
rect 34422 20992 34428 21004
rect 34379 20964 34428 20992
rect 34379 20961 34391 20964
rect 34333 20955 34391 20961
rect 34422 20952 34428 20964
rect 34480 20952 34486 21004
rect 34698 20992 34704 21004
rect 34659 20964 34704 20992
rect 34698 20952 34704 20964
rect 34756 20952 34762 21004
rect 34885 20995 34943 21001
rect 34885 20961 34897 20995
rect 34931 20961 34943 20995
rect 34885 20955 34943 20961
rect 35529 20995 35587 21001
rect 35529 20961 35541 20995
rect 35575 20992 35587 20995
rect 35710 20992 35716 21004
rect 35575 20964 35716 20992
rect 35575 20961 35587 20964
rect 35529 20955 35587 20961
rect 34900 20924 34928 20955
rect 35710 20952 35716 20964
rect 35768 20952 35774 21004
rect 36630 20992 36636 21004
rect 36591 20964 36636 20992
rect 36630 20952 36636 20964
rect 36688 20952 36694 21004
rect 36998 20992 37004 21004
rect 36959 20964 37004 20992
rect 36998 20952 37004 20964
rect 37056 20952 37062 21004
rect 37737 20995 37795 21001
rect 37737 20961 37749 20995
rect 37783 20961 37795 20995
rect 37737 20955 37795 20961
rect 36814 20924 36820 20936
rect 34256 20896 34928 20924
rect 36775 20896 36820 20924
rect 36814 20884 36820 20896
rect 36872 20884 36878 20936
rect 27632 20828 28948 20856
rect 7098 20788 7104 20800
rect 7059 20760 7104 20788
rect 7098 20748 7104 20760
rect 7156 20748 7162 20800
rect 17218 20748 17224 20800
rect 17276 20788 17282 20800
rect 19521 20791 19579 20797
rect 19521 20788 19533 20791
rect 17276 20760 19533 20788
rect 17276 20748 17282 20760
rect 19521 20757 19533 20760
rect 19567 20757 19579 20791
rect 19521 20751 19579 20757
rect 21453 20791 21511 20797
rect 21453 20757 21465 20791
rect 21499 20788 21511 20791
rect 22002 20788 22008 20800
rect 21499 20760 22008 20788
rect 21499 20757 21511 20760
rect 21453 20751 21511 20757
rect 22002 20748 22008 20760
rect 22060 20748 22066 20800
rect 23014 20748 23020 20800
rect 23072 20788 23078 20800
rect 25317 20791 25375 20797
rect 25317 20788 25329 20791
rect 23072 20760 25329 20788
rect 23072 20748 23078 20760
rect 25317 20757 25329 20760
rect 25363 20757 25375 20791
rect 25317 20751 25375 20757
rect 28074 20748 28080 20800
rect 28132 20788 28138 20800
rect 28169 20791 28227 20797
rect 28169 20788 28181 20791
rect 28132 20760 28181 20788
rect 28132 20748 28138 20760
rect 28169 20757 28181 20760
rect 28215 20757 28227 20791
rect 28920 20788 28948 20828
rect 30190 20816 30196 20868
rect 30248 20856 30254 20868
rect 31481 20859 31539 20865
rect 31481 20856 31493 20859
rect 30248 20828 31493 20856
rect 30248 20816 30254 20828
rect 31481 20825 31493 20828
rect 31527 20825 31539 20859
rect 31481 20819 31539 20825
rect 30650 20788 30656 20800
rect 28920 20760 30656 20788
rect 28169 20751 28227 20757
rect 30650 20748 30656 20760
rect 30708 20748 30714 20800
rect 31662 20748 31668 20800
rect 31720 20788 31726 20800
rect 37752 20788 37780 20955
rect 31720 20760 37780 20788
rect 31720 20748 31726 20760
rect 1104 20698 38824 20720
rect 1104 20646 4246 20698
rect 4298 20646 4310 20698
rect 4362 20646 4374 20698
rect 4426 20646 4438 20698
rect 4490 20646 34966 20698
rect 35018 20646 35030 20698
rect 35082 20646 35094 20698
rect 35146 20646 35158 20698
rect 35210 20646 38824 20698
rect 1104 20624 38824 20646
rect 3510 20544 3516 20596
rect 3568 20584 3574 20596
rect 3605 20587 3663 20593
rect 3605 20584 3617 20587
rect 3568 20556 3617 20584
rect 3568 20544 3574 20556
rect 3605 20553 3617 20556
rect 3651 20553 3663 20587
rect 3605 20547 3663 20553
rect 8938 20544 8944 20596
rect 8996 20584 9002 20596
rect 10597 20587 10655 20593
rect 10597 20584 10609 20587
rect 8996 20556 10609 20584
rect 8996 20544 9002 20556
rect 10597 20553 10609 20556
rect 10643 20553 10655 20587
rect 13998 20584 14004 20596
rect 13959 20556 14004 20584
rect 10597 20547 10655 20553
rect 13998 20544 14004 20556
rect 14056 20544 14062 20596
rect 14550 20584 14556 20596
rect 14463 20556 14556 20584
rect 14550 20544 14556 20556
rect 14608 20584 14614 20596
rect 14826 20584 14832 20596
rect 14608 20556 14832 20584
rect 14608 20544 14614 20556
rect 14826 20544 14832 20556
rect 14884 20544 14890 20596
rect 19334 20544 19340 20596
rect 19392 20584 19398 20596
rect 20073 20587 20131 20593
rect 20073 20584 20085 20587
rect 19392 20556 20085 20584
rect 19392 20544 19398 20556
rect 20073 20553 20085 20556
rect 20119 20553 20131 20587
rect 20073 20547 20131 20553
rect 20625 20587 20683 20593
rect 20625 20553 20637 20587
rect 20671 20584 20683 20587
rect 20806 20584 20812 20596
rect 20671 20556 20812 20584
rect 20671 20553 20683 20556
rect 20625 20547 20683 20553
rect 20806 20544 20812 20556
rect 20864 20544 20870 20596
rect 22922 20544 22928 20596
rect 22980 20584 22986 20596
rect 23293 20587 23351 20593
rect 23293 20584 23305 20587
rect 22980 20556 23305 20584
rect 22980 20544 22986 20556
rect 23293 20553 23305 20556
rect 23339 20553 23351 20587
rect 23293 20547 23351 20553
rect 24118 20544 24124 20596
rect 24176 20584 24182 20596
rect 24489 20587 24547 20593
rect 24489 20584 24501 20587
rect 24176 20556 24501 20584
rect 24176 20544 24182 20556
rect 24489 20553 24501 20556
rect 24535 20553 24547 20587
rect 27430 20584 27436 20596
rect 24489 20547 24547 20553
rect 25424 20556 27436 20584
rect 4982 20476 4988 20528
rect 5040 20516 5046 20528
rect 5169 20519 5227 20525
rect 5169 20516 5181 20519
rect 5040 20488 5181 20516
rect 5040 20476 5046 20488
rect 5169 20485 5181 20488
rect 5215 20485 5227 20519
rect 5169 20479 5227 20485
rect 7742 20476 7748 20528
rect 7800 20516 7806 20528
rect 12434 20516 12440 20528
rect 7800 20488 9260 20516
rect 7800 20476 7806 20488
rect 1578 20408 1584 20460
rect 1636 20448 1642 20460
rect 1673 20451 1731 20457
rect 1673 20448 1685 20451
rect 1636 20420 1685 20448
rect 1636 20408 1642 20420
rect 1673 20417 1685 20420
rect 1719 20417 1731 20451
rect 7098 20448 7104 20460
rect 7059 20420 7104 20448
rect 1673 20411 1731 20417
rect 7098 20408 7104 20420
rect 7156 20408 7162 20460
rect 9030 20448 9036 20460
rect 7208 20420 9036 20448
rect 1394 20380 1400 20392
rect 1355 20352 1400 20380
rect 1394 20340 1400 20352
rect 1452 20340 1458 20392
rect 3053 20383 3111 20389
rect 3053 20349 3065 20383
rect 3099 20380 3111 20383
rect 3418 20380 3424 20392
rect 3099 20352 3424 20380
rect 3099 20349 3111 20352
rect 3053 20343 3111 20349
rect 3418 20340 3424 20352
rect 3476 20380 3482 20392
rect 3513 20383 3571 20389
rect 3513 20380 3525 20383
rect 3476 20352 3525 20380
rect 3476 20340 3482 20352
rect 3513 20349 3525 20352
rect 3559 20349 3571 20383
rect 3513 20343 3571 20349
rect 4525 20383 4583 20389
rect 4525 20349 4537 20383
rect 4571 20380 4583 20383
rect 4706 20380 4712 20392
rect 4571 20352 4712 20380
rect 4571 20349 4583 20352
rect 4525 20343 4583 20349
rect 4706 20340 4712 20352
rect 4764 20340 4770 20392
rect 4890 20380 4896 20392
rect 4851 20352 4896 20380
rect 4890 20340 4896 20352
rect 4948 20340 4954 20392
rect 5258 20380 5264 20392
rect 5219 20352 5264 20380
rect 5258 20340 5264 20352
rect 5316 20340 5322 20392
rect 5902 20380 5908 20392
rect 5863 20352 5908 20380
rect 5902 20340 5908 20352
rect 5960 20340 5966 20392
rect 7009 20383 7067 20389
rect 7009 20349 7021 20383
rect 7055 20380 7067 20383
rect 7208 20380 7236 20420
rect 9030 20408 9036 20420
rect 9088 20408 9094 20460
rect 9232 20457 9260 20488
rect 10152 20488 12440 20516
rect 9217 20451 9275 20457
rect 9217 20417 9229 20451
rect 9263 20417 9275 20451
rect 9490 20448 9496 20460
rect 9451 20420 9496 20448
rect 9217 20411 9275 20417
rect 9490 20408 9496 20420
rect 9548 20408 9554 20460
rect 7055 20352 7236 20380
rect 7055 20349 7067 20352
rect 7009 20343 7067 20349
rect 7282 20340 7288 20392
rect 7340 20380 7346 20392
rect 7653 20383 7711 20389
rect 7340 20352 7385 20380
rect 7340 20340 7346 20352
rect 7653 20349 7665 20383
rect 7699 20349 7711 20383
rect 8110 20380 8116 20392
rect 8071 20352 8116 20380
rect 7653 20343 7711 20349
rect 6089 20247 6147 20253
rect 6089 20213 6101 20247
rect 6135 20244 6147 20247
rect 6362 20244 6368 20256
rect 6135 20216 6368 20244
rect 6135 20213 6147 20216
rect 6089 20207 6147 20213
rect 6362 20204 6368 20216
rect 6420 20244 6426 20256
rect 7668 20244 7696 20343
rect 8110 20340 8116 20352
rect 8168 20340 8174 20392
rect 8202 20340 8208 20392
rect 8260 20380 8266 20392
rect 8757 20383 8815 20389
rect 8757 20380 8769 20383
rect 8260 20352 8769 20380
rect 8260 20340 8266 20352
rect 8757 20349 8769 20352
rect 8803 20380 8815 20383
rect 10152 20380 10180 20488
rect 12434 20476 12440 20488
rect 12492 20476 12498 20528
rect 15746 20516 15752 20528
rect 15707 20488 15752 20516
rect 15746 20476 15752 20488
rect 15804 20476 15810 20528
rect 21266 20516 21272 20528
rect 20272 20488 21272 20516
rect 11885 20451 11943 20457
rect 11885 20417 11897 20451
rect 11931 20448 11943 20451
rect 12713 20451 12771 20457
rect 12713 20448 12725 20451
rect 11931 20420 12725 20448
rect 11931 20417 11943 20420
rect 11885 20411 11943 20417
rect 12713 20417 12725 20420
rect 12759 20417 12771 20451
rect 12713 20411 12771 20417
rect 14921 20451 14979 20457
rect 14921 20417 14933 20451
rect 14967 20448 14979 20451
rect 20272 20448 20300 20488
rect 21266 20476 21272 20488
rect 21324 20476 21330 20528
rect 21542 20476 21548 20528
rect 21600 20516 21606 20528
rect 21726 20516 21732 20528
rect 21600 20488 21732 20516
rect 21600 20476 21606 20488
rect 21726 20476 21732 20488
rect 21784 20516 21790 20528
rect 23845 20519 23903 20525
rect 23845 20516 23857 20519
rect 21784 20488 23857 20516
rect 21784 20476 21790 20488
rect 23845 20485 23857 20488
rect 23891 20485 23903 20519
rect 23845 20479 23903 20485
rect 14967 20420 20300 20448
rect 14967 20417 14979 20420
rect 14921 20411 14979 20417
rect 20898 20408 20904 20460
rect 20956 20448 20962 20460
rect 21358 20448 21364 20460
rect 20956 20420 21364 20448
rect 20956 20408 20962 20420
rect 21358 20408 21364 20420
rect 21416 20448 21422 20460
rect 21416 20420 21864 20448
rect 21416 20408 21422 20420
rect 8803 20352 10180 20380
rect 11333 20383 11391 20389
rect 8803 20349 8815 20352
rect 8757 20343 8815 20349
rect 11333 20349 11345 20383
rect 11379 20349 11391 20383
rect 11333 20343 11391 20349
rect 6420 20216 7696 20244
rect 11348 20244 11376 20343
rect 11422 20340 11428 20392
rect 11480 20380 11486 20392
rect 12437 20383 12495 20389
rect 11480 20352 11525 20380
rect 11480 20340 11486 20352
rect 12437 20349 12449 20383
rect 12483 20380 12495 20383
rect 12526 20380 12532 20392
rect 12483 20352 12532 20380
rect 12483 20349 12495 20352
rect 12437 20343 12495 20349
rect 12526 20340 12532 20352
rect 12584 20380 12590 20392
rect 14550 20380 14556 20392
rect 12584 20352 14556 20380
rect 12584 20340 12590 20352
rect 14550 20340 14556 20352
rect 14608 20340 14614 20392
rect 14734 20380 14740 20392
rect 14695 20352 14740 20380
rect 14734 20340 14740 20352
rect 14792 20340 14798 20392
rect 14826 20340 14832 20392
rect 14884 20380 14890 20392
rect 15470 20380 15476 20392
rect 14884 20352 14929 20380
rect 15431 20352 15476 20380
rect 14884 20340 14890 20352
rect 15470 20340 15476 20352
rect 15528 20340 15534 20392
rect 16117 20383 16175 20389
rect 16117 20349 16129 20383
rect 16163 20349 16175 20383
rect 16298 20380 16304 20392
rect 16259 20352 16304 20380
rect 16117 20343 16175 20349
rect 16132 20312 16160 20343
rect 16298 20340 16304 20352
rect 16356 20340 16362 20392
rect 17034 20380 17040 20392
rect 16995 20352 17040 20380
rect 17034 20340 17040 20352
rect 17092 20340 17098 20392
rect 18414 20340 18420 20392
rect 18472 20380 18478 20392
rect 18601 20383 18659 20389
rect 18601 20380 18613 20383
rect 18472 20352 18613 20380
rect 18472 20340 18478 20352
rect 18601 20349 18613 20352
rect 18647 20349 18659 20383
rect 18601 20343 18659 20349
rect 18693 20383 18751 20389
rect 18693 20349 18705 20383
rect 18739 20380 18751 20383
rect 18782 20380 18788 20392
rect 18739 20352 18788 20380
rect 18739 20349 18751 20352
rect 18693 20343 18751 20349
rect 18782 20340 18788 20352
rect 18840 20340 18846 20392
rect 18969 20383 19027 20389
rect 18969 20349 18981 20383
rect 19015 20380 19027 20383
rect 19886 20380 19892 20392
rect 19015 20352 19892 20380
rect 19015 20349 19027 20352
rect 18969 20343 19027 20349
rect 19886 20340 19892 20352
rect 19944 20340 19950 20392
rect 20438 20380 20444 20392
rect 20399 20352 20444 20380
rect 20438 20340 20444 20352
rect 20496 20340 20502 20392
rect 20530 20340 20536 20392
rect 20588 20380 20594 20392
rect 21836 20389 21864 20420
rect 22738 20408 22744 20460
rect 22796 20448 22802 20460
rect 25424 20448 25452 20556
rect 27430 20544 27436 20556
rect 27488 20544 27494 20596
rect 29457 20587 29515 20593
rect 29457 20553 29469 20587
rect 29503 20584 29515 20587
rect 29638 20584 29644 20596
rect 29503 20556 29644 20584
rect 29503 20553 29515 20556
rect 29457 20547 29515 20553
rect 29638 20544 29644 20556
rect 29696 20544 29702 20596
rect 30926 20544 30932 20596
rect 30984 20584 30990 20596
rect 31389 20587 31447 20593
rect 31389 20584 31401 20587
rect 30984 20556 31401 20584
rect 30984 20544 30990 20556
rect 31389 20553 31401 20556
rect 31435 20584 31447 20587
rect 31570 20584 31576 20596
rect 31435 20556 31576 20584
rect 31435 20553 31447 20556
rect 31389 20547 31447 20553
rect 31570 20544 31576 20556
rect 31628 20544 31634 20596
rect 37642 20584 37648 20596
rect 37603 20556 37648 20584
rect 37642 20544 37648 20556
rect 37700 20544 37706 20596
rect 27798 20476 27804 20528
rect 27856 20516 27862 20528
rect 28445 20519 28503 20525
rect 28445 20516 28457 20519
rect 27856 20488 28457 20516
rect 27856 20476 27862 20488
rect 28445 20485 28457 20488
rect 28491 20485 28503 20519
rect 28445 20479 28503 20485
rect 35250 20476 35256 20528
rect 35308 20516 35314 20528
rect 36262 20516 36268 20528
rect 35308 20488 36268 20516
rect 35308 20476 35314 20488
rect 36262 20476 36268 20488
rect 36320 20476 36326 20528
rect 22796 20420 25452 20448
rect 25501 20451 25559 20457
rect 22796 20408 22802 20420
rect 25501 20417 25513 20451
rect 25547 20448 25559 20451
rect 27154 20448 27160 20460
rect 25547 20420 27160 20448
rect 25547 20417 25559 20420
rect 25501 20411 25559 20417
rect 27154 20408 27160 20420
rect 27212 20408 27218 20460
rect 30285 20451 30343 20457
rect 30285 20417 30297 20451
rect 30331 20448 30343 20451
rect 33045 20451 33103 20457
rect 33045 20448 33057 20451
rect 30331 20420 33057 20448
rect 30331 20417 30343 20420
rect 30285 20411 30343 20417
rect 33045 20417 33057 20420
rect 33091 20417 33103 20451
rect 33045 20411 33103 20417
rect 35437 20451 35495 20457
rect 35437 20417 35449 20451
rect 35483 20448 35495 20451
rect 36541 20451 36599 20457
rect 36541 20448 36553 20451
rect 35483 20420 36553 20448
rect 35483 20417 35495 20420
rect 35437 20411 35495 20417
rect 36541 20417 36553 20420
rect 36587 20417 36599 20451
rect 36541 20411 36599 20417
rect 20809 20383 20867 20389
rect 20809 20380 20821 20383
rect 20588 20352 20821 20380
rect 20588 20340 20594 20352
rect 20809 20349 20821 20352
rect 20855 20349 20867 20383
rect 20809 20343 20867 20349
rect 21637 20383 21695 20389
rect 21637 20349 21649 20383
rect 21683 20349 21695 20383
rect 21637 20343 21695 20349
rect 21821 20383 21879 20389
rect 21821 20349 21833 20383
rect 21867 20349 21879 20383
rect 21821 20343 21879 20349
rect 22557 20383 22615 20389
rect 22557 20349 22569 20383
rect 22603 20349 22615 20383
rect 22557 20343 22615 20349
rect 23477 20383 23535 20389
rect 23477 20349 23489 20383
rect 23523 20380 23535 20383
rect 23566 20380 23572 20392
rect 23523 20352 23572 20380
rect 23523 20349 23535 20352
rect 23477 20343 23535 20349
rect 17678 20312 17684 20324
rect 16132 20284 17684 20312
rect 17678 20272 17684 20284
rect 17736 20272 17742 20324
rect 21652 20312 21680 20343
rect 22186 20312 22192 20324
rect 21652 20284 22192 20312
rect 22186 20272 22192 20284
rect 22244 20312 22250 20324
rect 22572 20312 22600 20343
rect 23566 20340 23572 20352
rect 23624 20340 23630 20392
rect 23658 20340 23664 20392
rect 23716 20380 23722 20392
rect 24397 20383 24455 20389
rect 24397 20380 24409 20383
rect 23716 20352 24409 20380
rect 23716 20340 23722 20352
rect 24397 20349 24409 20352
rect 24443 20349 24455 20383
rect 24397 20343 24455 20349
rect 25777 20383 25835 20389
rect 25777 20349 25789 20383
rect 25823 20380 25835 20383
rect 26050 20380 26056 20392
rect 25823 20352 26056 20380
rect 25823 20349 25835 20352
rect 25777 20343 25835 20349
rect 26050 20340 26056 20352
rect 26108 20340 26114 20392
rect 26786 20340 26792 20392
rect 26844 20380 26850 20392
rect 27617 20383 27675 20389
rect 27617 20380 27629 20383
rect 26844 20352 27629 20380
rect 26844 20340 26850 20352
rect 27617 20349 27629 20352
rect 27663 20349 27675 20383
rect 28166 20380 28172 20392
rect 28127 20352 28172 20380
rect 27617 20343 27675 20349
rect 28166 20340 28172 20352
rect 28224 20340 28230 20392
rect 28442 20380 28448 20392
rect 28403 20352 28448 20380
rect 28442 20340 28448 20352
rect 28500 20340 28506 20392
rect 29270 20380 29276 20392
rect 29231 20352 29276 20380
rect 29270 20340 29276 20352
rect 29328 20340 29334 20392
rect 30006 20380 30012 20392
rect 29967 20352 30012 20380
rect 30006 20340 30012 20352
rect 30064 20340 30070 20392
rect 32306 20380 32312 20392
rect 32267 20352 32312 20380
rect 32306 20340 32312 20352
rect 32364 20340 32370 20392
rect 32493 20383 32551 20389
rect 32493 20349 32505 20383
rect 32539 20349 32551 20383
rect 32493 20343 32551 20349
rect 32953 20383 33011 20389
rect 32953 20349 32965 20383
rect 32999 20380 33011 20383
rect 33226 20380 33232 20392
rect 32999 20352 33232 20380
rect 32999 20349 33011 20352
rect 32953 20343 33011 20349
rect 22244 20284 22600 20312
rect 29288 20312 29316 20340
rect 30098 20312 30104 20324
rect 29288 20284 30104 20312
rect 22244 20272 22250 20284
rect 30098 20272 30104 20284
rect 30156 20272 30162 20324
rect 32122 20272 32128 20324
rect 32180 20312 32186 20324
rect 32508 20312 32536 20343
rect 33226 20340 33232 20352
rect 33284 20340 33290 20392
rect 33962 20380 33968 20392
rect 33923 20352 33968 20380
rect 33962 20340 33968 20352
rect 34020 20340 34026 20392
rect 35345 20383 35403 20389
rect 35345 20349 35357 20383
rect 35391 20349 35403 20383
rect 35710 20380 35716 20392
rect 35671 20352 35716 20380
rect 35345 20343 35403 20349
rect 32180 20284 32536 20312
rect 33781 20315 33839 20321
rect 32180 20272 32186 20284
rect 33781 20281 33793 20315
rect 33827 20281 33839 20315
rect 33781 20275 33839 20281
rect 34333 20315 34391 20321
rect 34333 20281 34345 20315
rect 34379 20312 34391 20315
rect 34422 20312 34428 20324
rect 34379 20284 34428 20312
rect 34379 20281 34391 20284
rect 34333 20275 34391 20281
rect 12434 20244 12440 20256
rect 11348 20216 12440 20244
rect 6420 20204 6426 20216
rect 12434 20204 12440 20216
rect 12492 20204 12498 20256
rect 17221 20247 17279 20253
rect 17221 20213 17233 20247
rect 17267 20244 17279 20247
rect 17310 20244 17316 20256
rect 17267 20216 17316 20244
rect 17267 20213 17279 20216
rect 17221 20207 17279 20213
rect 17310 20204 17316 20216
rect 17368 20204 17374 20256
rect 17862 20204 17868 20256
rect 17920 20244 17926 20256
rect 18417 20247 18475 20253
rect 18417 20244 18429 20247
rect 17920 20216 18429 20244
rect 17920 20204 17926 20216
rect 18417 20213 18429 20216
rect 18463 20213 18475 20247
rect 18417 20207 18475 20213
rect 18966 20204 18972 20256
rect 19024 20244 19030 20256
rect 20993 20247 21051 20253
rect 20993 20244 21005 20247
rect 19024 20216 21005 20244
rect 19024 20204 19030 20216
rect 20993 20213 21005 20216
rect 21039 20213 21051 20247
rect 21450 20244 21456 20256
rect 21411 20216 21456 20244
rect 20993 20207 21051 20213
rect 21450 20204 21456 20216
rect 21508 20204 21514 20256
rect 22370 20204 22376 20256
rect 22428 20244 22434 20256
rect 22741 20247 22799 20253
rect 22741 20244 22753 20247
rect 22428 20216 22753 20244
rect 22428 20204 22434 20216
rect 22741 20213 22753 20216
rect 22787 20213 22799 20247
rect 22741 20207 22799 20213
rect 22922 20204 22928 20256
rect 22980 20244 22986 20256
rect 23842 20244 23848 20256
rect 22980 20216 23848 20244
rect 22980 20204 22986 20216
rect 23842 20204 23848 20216
rect 23900 20204 23906 20256
rect 25866 20204 25872 20256
rect 25924 20244 25930 20256
rect 26881 20247 26939 20253
rect 26881 20244 26893 20247
rect 25924 20216 26893 20244
rect 25924 20204 25930 20216
rect 26881 20213 26893 20216
rect 26927 20213 26939 20247
rect 26881 20207 26939 20213
rect 27430 20204 27436 20256
rect 27488 20244 27494 20256
rect 30374 20244 30380 20256
rect 27488 20216 30380 20244
rect 27488 20204 27494 20216
rect 30374 20204 30380 20216
rect 30432 20204 30438 20256
rect 32950 20204 32956 20256
rect 33008 20244 33014 20256
rect 33796 20244 33824 20275
rect 34422 20272 34428 20284
rect 34480 20272 34486 20324
rect 35360 20312 35388 20343
rect 35710 20340 35716 20352
rect 35768 20340 35774 20392
rect 36262 20380 36268 20392
rect 36223 20352 36268 20380
rect 36262 20340 36268 20352
rect 36320 20340 36326 20392
rect 37826 20380 37832 20392
rect 36372 20352 37832 20380
rect 36372 20312 36400 20352
rect 37826 20340 37832 20352
rect 37884 20340 37890 20392
rect 35360 20284 36400 20312
rect 34698 20244 34704 20256
rect 33008 20216 34704 20244
rect 33008 20204 33014 20216
rect 34698 20204 34704 20216
rect 34756 20204 34762 20256
rect 35342 20204 35348 20256
rect 35400 20244 35406 20256
rect 35710 20244 35716 20256
rect 35400 20216 35716 20244
rect 35400 20204 35406 20216
rect 35710 20204 35716 20216
rect 35768 20204 35774 20256
rect 1104 20154 38824 20176
rect 1104 20102 19606 20154
rect 19658 20102 19670 20154
rect 19722 20102 19734 20154
rect 19786 20102 19798 20154
rect 19850 20102 38824 20154
rect 1104 20080 38824 20102
rect 2866 20040 2872 20052
rect 2424 20012 2872 20040
rect 1946 19864 1952 19916
rect 2004 19904 2010 19916
rect 2424 19913 2452 20012
rect 2866 20000 2872 20012
rect 2924 20000 2930 20052
rect 4065 20043 4123 20049
rect 4065 20009 4077 20043
rect 4111 20040 4123 20043
rect 4249 20043 4307 20049
rect 4249 20040 4261 20043
rect 4111 20012 4261 20040
rect 4111 20009 4123 20012
rect 4065 20003 4123 20009
rect 4249 20009 4261 20012
rect 4295 20009 4307 20043
rect 4249 20003 4307 20009
rect 4614 20000 4620 20052
rect 4672 20000 4678 20052
rect 11422 20000 11428 20052
rect 11480 20040 11486 20052
rect 11517 20043 11575 20049
rect 11517 20040 11529 20043
rect 11480 20012 11529 20040
rect 11480 20000 11486 20012
rect 11517 20009 11529 20012
rect 11563 20009 11575 20043
rect 11517 20003 11575 20009
rect 11882 20000 11888 20052
rect 11940 20040 11946 20052
rect 12526 20040 12532 20052
rect 11940 20012 12532 20040
rect 11940 20000 11946 20012
rect 12526 20000 12532 20012
rect 12584 20000 12590 20052
rect 13446 20040 13452 20052
rect 13407 20012 13452 20040
rect 13446 20000 13452 20012
rect 13504 20000 13510 20052
rect 17862 20040 17868 20052
rect 15120 20012 17868 20040
rect 4632 19972 4660 20000
rect 3252 19944 4660 19972
rect 3252 19913 3280 19944
rect 4890 19932 4896 19984
rect 4948 19972 4954 19984
rect 8386 19972 8392 19984
rect 4948 19944 6960 19972
rect 4948 19932 4954 19944
rect 2409 19907 2467 19913
rect 2409 19904 2421 19907
rect 2004 19876 2421 19904
rect 2004 19864 2010 19876
rect 2409 19873 2421 19876
rect 2455 19873 2467 19907
rect 2409 19867 2467 19873
rect 3237 19907 3295 19913
rect 3237 19873 3249 19907
rect 3283 19873 3295 19907
rect 3237 19867 3295 19873
rect 3421 19907 3479 19913
rect 3421 19873 3433 19907
rect 3467 19904 3479 19907
rect 4065 19907 4123 19913
rect 4065 19904 4077 19907
rect 3467 19876 4077 19904
rect 3467 19873 3479 19876
rect 3421 19867 3479 19873
rect 4065 19873 4077 19876
rect 4111 19873 4123 19907
rect 4065 19867 4123 19873
rect 4433 19907 4491 19913
rect 4433 19873 4445 19907
rect 4479 19904 4491 19907
rect 4522 19904 4528 19916
rect 4479 19876 4528 19904
rect 4479 19873 4491 19876
rect 4433 19867 4491 19873
rect 3142 19796 3148 19848
rect 3200 19836 3206 19848
rect 3436 19836 3464 19867
rect 4522 19864 4528 19876
rect 4580 19864 4586 19916
rect 4617 19907 4675 19913
rect 4617 19873 4629 19907
rect 4663 19873 4675 19907
rect 4617 19867 4675 19873
rect 3200 19808 3464 19836
rect 4632 19836 4660 19867
rect 4706 19864 4712 19916
rect 4764 19904 4770 19916
rect 5460 19913 5488 19944
rect 5169 19907 5227 19913
rect 5169 19904 5181 19907
rect 4764 19876 5181 19904
rect 4764 19864 4770 19876
rect 5169 19873 5181 19876
rect 5215 19873 5227 19907
rect 5169 19867 5227 19873
rect 5445 19907 5503 19913
rect 5445 19873 5457 19907
rect 5491 19873 5503 19907
rect 6362 19904 6368 19916
rect 6323 19876 6368 19904
rect 5445 19867 5503 19873
rect 5184 19836 5212 19867
rect 6362 19864 6368 19876
rect 6420 19864 6426 19916
rect 6932 19913 6960 19944
rect 8220 19944 8392 19972
rect 6917 19907 6975 19913
rect 6917 19873 6929 19907
rect 6963 19904 6975 19907
rect 7282 19904 7288 19916
rect 6963 19876 7288 19904
rect 6963 19873 6975 19876
rect 6917 19867 6975 19873
rect 7282 19864 7288 19876
rect 7340 19864 7346 19916
rect 8220 19913 8248 19944
rect 8386 19932 8392 19944
rect 8444 19972 8450 19984
rect 8938 19972 8944 19984
rect 8444 19944 8944 19972
rect 8444 19932 8450 19944
rect 8938 19932 8944 19944
rect 8996 19932 9002 19984
rect 7561 19907 7619 19913
rect 7561 19873 7573 19907
rect 7607 19873 7619 19907
rect 7561 19867 7619 19873
rect 8205 19907 8263 19913
rect 8205 19873 8217 19907
rect 8251 19873 8263 19907
rect 8205 19867 8263 19873
rect 8297 19907 8355 19913
rect 8297 19873 8309 19907
rect 8343 19873 8355 19907
rect 9030 19904 9036 19916
rect 8991 19876 9036 19904
rect 8297 19867 8355 19873
rect 6380 19836 6408 19864
rect 4632 19808 4752 19836
rect 5184 19808 6408 19836
rect 7101 19839 7159 19845
rect 3200 19796 3206 19808
rect 2958 19728 2964 19780
rect 3016 19768 3022 19780
rect 3237 19771 3295 19777
rect 3237 19768 3249 19771
rect 3016 19740 3249 19768
rect 3016 19728 3022 19740
rect 3237 19737 3249 19740
rect 3283 19737 3295 19771
rect 4724 19768 4752 19808
rect 7101 19805 7113 19839
rect 7147 19836 7159 19839
rect 7466 19836 7472 19848
rect 7147 19808 7472 19836
rect 7147 19805 7159 19808
rect 7101 19799 7159 19805
rect 7466 19796 7472 19808
rect 7524 19796 7530 19848
rect 5258 19768 5264 19780
rect 4724 19740 5264 19768
rect 3237 19731 3295 19737
rect 5258 19728 5264 19740
rect 5316 19728 5322 19780
rect 7282 19728 7288 19780
rect 7340 19768 7346 19780
rect 7576 19768 7604 19867
rect 8312 19836 8340 19867
rect 9030 19864 9036 19876
rect 9088 19864 9094 19916
rect 10137 19907 10195 19913
rect 10137 19873 10149 19907
rect 10183 19904 10195 19907
rect 11882 19904 11888 19916
rect 10183 19876 11888 19904
rect 10183 19873 10195 19876
rect 10137 19867 10195 19873
rect 11882 19864 11888 19876
rect 11940 19864 11946 19916
rect 12342 19904 12348 19916
rect 12303 19876 12348 19904
rect 12342 19864 12348 19876
rect 12400 19864 12406 19916
rect 13538 19904 13544 19916
rect 13499 19876 13544 19904
rect 13538 19864 13544 19876
rect 13596 19864 13602 19916
rect 13998 19904 14004 19916
rect 13959 19876 14004 19904
rect 13998 19864 14004 19876
rect 14056 19864 14062 19916
rect 14090 19864 14096 19916
rect 14148 19904 14154 19916
rect 15120 19913 15148 20012
rect 17862 20000 17868 20012
rect 17920 20000 17926 20052
rect 20254 20000 20260 20052
rect 20312 20040 20318 20052
rect 21453 20043 21511 20049
rect 21453 20040 21465 20043
rect 20312 20012 21465 20040
rect 20312 20000 20318 20012
rect 21453 20009 21465 20012
rect 21499 20040 21511 20043
rect 21499 20012 23152 20040
rect 21499 20009 21511 20012
rect 21453 20003 21511 20009
rect 15289 19975 15347 19981
rect 15289 19941 15301 19975
rect 15335 19972 15347 19975
rect 15841 19975 15899 19981
rect 15335 19944 15608 19972
rect 15335 19941 15347 19944
rect 15289 19935 15347 19941
rect 14185 19907 14243 19913
rect 14185 19904 14197 19907
rect 14148 19876 14197 19904
rect 14148 19864 14154 19876
rect 14185 19873 14197 19876
rect 14231 19873 14243 19907
rect 14185 19867 14243 19873
rect 15105 19907 15163 19913
rect 15105 19873 15117 19907
rect 15151 19873 15163 19907
rect 15470 19904 15476 19916
rect 15431 19876 15476 19904
rect 15105 19867 15163 19873
rect 15470 19864 15476 19876
rect 15528 19864 15534 19916
rect 15580 19904 15608 19944
rect 15841 19941 15853 19975
rect 15887 19972 15899 19975
rect 16298 19972 16304 19984
rect 15887 19944 16304 19972
rect 15887 19941 15899 19944
rect 15841 19935 15899 19941
rect 16298 19932 16304 19944
rect 16356 19932 16362 19984
rect 20714 19932 20720 19984
rect 20772 19972 20778 19984
rect 21174 19972 21180 19984
rect 20772 19944 21180 19972
rect 20772 19932 20778 19944
rect 21174 19932 21180 19944
rect 21232 19972 21238 19984
rect 23124 19972 23152 20012
rect 23566 20000 23572 20052
rect 23624 20040 23630 20052
rect 23753 20043 23811 20049
rect 23753 20040 23765 20043
rect 23624 20012 23765 20040
rect 23624 20000 23630 20012
rect 23753 20009 23765 20012
rect 23799 20009 23811 20043
rect 23753 20003 23811 20009
rect 23842 20000 23848 20052
rect 23900 20040 23906 20052
rect 25869 20043 25927 20049
rect 23900 20012 24440 20040
rect 23900 20000 23906 20012
rect 21232 19944 23060 19972
rect 23124 19944 24164 19972
rect 21232 19932 21238 19944
rect 16022 19904 16028 19916
rect 15580 19876 16028 19904
rect 16022 19864 16028 19876
rect 16080 19864 16086 19916
rect 16577 19907 16635 19913
rect 16577 19873 16589 19907
rect 16623 19904 16635 19907
rect 17586 19904 17592 19916
rect 16623 19876 17592 19904
rect 16623 19873 16635 19876
rect 16577 19867 16635 19873
rect 17586 19864 17592 19876
rect 17644 19864 17650 19916
rect 18966 19904 18972 19916
rect 18927 19876 18972 19904
rect 18966 19864 18972 19876
rect 19024 19864 19030 19916
rect 21376 19913 21404 19944
rect 21361 19907 21419 19913
rect 21361 19873 21373 19907
rect 21407 19904 21419 19907
rect 21910 19904 21916 19916
rect 21407 19876 21441 19904
rect 21871 19876 21916 19904
rect 21407 19873 21419 19876
rect 21361 19867 21419 19873
rect 21910 19864 21916 19876
rect 21968 19864 21974 19916
rect 22186 19864 22192 19916
rect 22244 19904 22250 19916
rect 23032 19913 23060 19944
rect 22557 19907 22615 19913
rect 22557 19904 22569 19907
rect 22244 19876 22569 19904
rect 22244 19864 22250 19876
rect 22557 19873 22569 19876
rect 22603 19873 22615 19907
rect 22557 19867 22615 19873
rect 23017 19907 23075 19913
rect 23017 19873 23029 19907
rect 23063 19873 23075 19907
rect 23017 19867 23075 19873
rect 23934 19864 23940 19916
rect 23992 19904 23998 19916
rect 24136 19913 24164 19944
rect 24412 19913 24440 20012
rect 25869 20009 25881 20043
rect 25915 20040 25927 20043
rect 25915 20012 26004 20040
rect 25915 20009 25927 20012
rect 25869 20003 25927 20009
rect 25130 19972 25136 19984
rect 25091 19944 25136 19972
rect 25130 19932 25136 19944
rect 25188 19932 25194 19984
rect 25976 19972 26004 20012
rect 26050 20000 26056 20052
rect 26108 20040 26114 20052
rect 27157 20043 27215 20049
rect 27157 20040 27169 20043
rect 26108 20012 27169 20040
rect 26108 20000 26114 20012
rect 27157 20009 27169 20012
rect 27203 20009 27215 20043
rect 27157 20003 27215 20009
rect 28629 20043 28687 20049
rect 28629 20009 28641 20043
rect 28675 20040 28687 20043
rect 29178 20040 29184 20052
rect 28675 20012 29184 20040
rect 28675 20009 28687 20012
rect 28629 20003 28687 20009
rect 29178 20000 29184 20012
rect 29236 20040 29242 20052
rect 29454 20040 29460 20052
rect 29236 20012 29460 20040
rect 29236 20000 29242 20012
rect 29454 20000 29460 20012
rect 29512 20000 29518 20052
rect 29917 20043 29975 20049
rect 29917 20009 29929 20043
rect 29963 20040 29975 20043
rect 30374 20040 30380 20052
rect 29963 20012 30380 20040
rect 29963 20009 29975 20012
rect 29917 20003 29975 20009
rect 30374 20000 30380 20012
rect 30432 20000 30438 20052
rect 30653 20043 30711 20049
rect 30653 20009 30665 20043
rect 30699 20040 30711 20043
rect 32030 20040 32036 20052
rect 30699 20012 32036 20040
rect 30699 20009 30711 20012
rect 30653 20003 30711 20009
rect 32030 20000 32036 20012
rect 32088 20000 32094 20052
rect 35986 20040 35992 20052
rect 32140 20012 35992 20040
rect 27522 19972 27528 19984
rect 25700 19944 25912 19972
rect 25976 19944 27528 19972
rect 24121 19907 24179 19913
rect 23992 19876 24037 19904
rect 23992 19864 23998 19876
rect 24121 19873 24133 19907
rect 24167 19873 24179 19907
rect 24121 19867 24179 19873
rect 24397 19907 24455 19913
rect 24397 19873 24409 19907
rect 24443 19873 24455 19907
rect 24397 19867 24455 19873
rect 24949 19907 25007 19913
rect 24949 19873 24961 19907
rect 24995 19904 25007 19907
rect 25700 19904 25728 19944
rect 24995 19876 25728 19904
rect 25777 19907 25835 19913
rect 24995 19873 25007 19876
rect 24949 19867 25007 19873
rect 25777 19873 25789 19907
rect 25823 19873 25835 19907
rect 25884 19904 25912 19944
rect 27522 19932 27528 19944
rect 27580 19932 27586 19984
rect 28994 19972 29000 19984
rect 28644 19944 29000 19972
rect 26970 19904 26976 19916
rect 25884 19876 26976 19904
rect 25777 19867 25835 19873
rect 7340 19740 7604 19768
rect 8220 19808 8340 19836
rect 10413 19839 10471 19845
rect 7340 19728 7346 19740
rect 6270 19660 6276 19712
rect 6328 19700 6334 19712
rect 8220 19700 8248 19808
rect 10413 19805 10425 19839
rect 10459 19836 10471 19839
rect 11054 19836 11060 19848
rect 10459 19808 11060 19836
rect 10459 19805 10471 19808
rect 10413 19799 10471 19805
rect 11054 19796 11060 19808
rect 11112 19796 11118 19848
rect 12253 19839 12311 19845
rect 12253 19805 12265 19839
rect 12299 19836 12311 19839
rect 12434 19836 12440 19848
rect 12299 19808 12440 19836
rect 12299 19805 12311 19808
rect 12253 19799 12311 19805
rect 12434 19796 12440 19808
rect 12492 19796 12498 19848
rect 16301 19839 16359 19845
rect 16301 19805 16313 19839
rect 16347 19836 16359 19839
rect 18782 19836 18788 19848
rect 16347 19808 18788 19836
rect 16347 19805 16359 19808
rect 16301 19799 16359 19805
rect 18782 19796 18788 19808
rect 18840 19796 18846 19848
rect 23106 19836 23112 19848
rect 23067 19808 23112 19836
rect 23106 19796 23112 19808
rect 23164 19796 23170 19848
rect 25792 19836 25820 19867
rect 26970 19864 26976 19876
rect 27028 19864 27034 19916
rect 27246 19904 27252 19916
rect 27207 19876 27252 19904
rect 27246 19864 27252 19876
rect 27304 19864 27310 19916
rect 27798 19904 27804 19916
rect 27759 19876 27804 19904
rect 27798 19864 27804 19876
rect 27856 19864 27862 19916
rect 28074 19904 28080 19916
rect 28035 19876 28080 19904
rect 28074 19864 28080 19876
rect 28132 19864 28138 19916
rect 28644 19836 28672 19944
rect 28994 19932 29000 19944
rect 29052 19932 29058 19984
rect 32140 19972 32168 20012
rect 35986 20000 35992 20012
rect 36044 20000 36050 20052
rect 29748 19944 32168 19972
rect 28813 19907 28871 19913
rect 28813 19873 28825 19907
rect 28859 19873 28871 19907
rect 28813 19867 28871 19873
rect 29089 19907 29147 19913
rect 29089 19873 29101 19907
rect 29135 19904 29147 19907
rect 29638 19904 29644 19916
rect 29135 19876 29644 19904
rect 29135 19873 29147 19876
rect 29089 19867 29147 19873
rect 25792 19808 28672 19836
rect 20070 19728 20076 19780
rect 20128 19768 20134 19780
rect 20257 19771 20315 19777
rect 20257 19768 20269 19771
rect 20128 19740 20269 19768
rect 20128 19728 20134 19740
rect 20257 19737 20269 19740
rect 20303 19737 20315 19771
rect 20257 19731 20315 19737
rect 21450 19728 21456 19780
rect 21508 19768 21514 19780
rect 22922 19768 22928 19780
rect 21508 19740 22928 19768
rect 21508 19728 21514 19740
rect 22922 19728 22928 19740
rect 22980 19728 22986 19780
rect 28828 19768 28856 19867
rect 29638 19864 29644 19876
rect 29696 19864 29702 19916
rect 29748 19913 29776 19944
rect 32582 19932 32588 19984
rect 32640 19972 32646 19984
rect 32861 19975 32919 19981
rect 32861 19972 32873 19975
rect 32640 19944 32873 19972
rect 32640 19932 32646 19944
rect 32861 19941 32873 19944
rect 32907 19941 32919 19975
rect 33410 19972 33416 19984
rect 33371 19944 33416 19972
rect 32861 19935 32919 19941
rect 33410 19932 33416 19944
rect 33468 19932 33474 19984
rect 35526 19972 35532 19984
rect 35487 19944 35532 19972
rect 35526 19932 35532 19944
rect 35584 19932 35590 19984
rect 29733 19907 29791 19913
rect 29733 19873 29745 19907
rect 29779 19873 29791 19907
rect 29733 19867 29791 19873
rect 29748 19768 29776 19867
rect 30098 19864 30104 19916
rect 30156 19904 30162 19916
rect 30469 19907 30527 19913
rect 30469 19904 30481 19907
rect 30156 19876 30481 19904
rect 30156 19864 30162 19876
rect 30469 19873 30481 19876
rect 30515 19873 30527 19907
rect 30469 19867 30527 19873
rect 31018 19864 31024 19916
rect 31076 19904 31082 19916
rect 31205 19907 31263 19913
rect 31205 19904 31217 19907
rect 31076 19876 31217 19904
rect 31076 19864 31082 19876
rect 31205 19873 31217 19876
rect 31251 19873 31263 19907
rect 32766 19904 32772 19916
rect 32727 19876 32772 19904
rect 31205 19867 31263 19873
rect 32766 19864 32772 19876
rect 32824 19864 32830 19916
rect 32950 19904 32956 19916
rect 32911 19876 32956 19904
rect 32950 19864 32956 19876
rect 33008 19864 33014 19916
rect 34146 19904 34152 19916
rect 34107 19876 34152 19904
rect 34146 19864 34152 19876
rect 34204 19864 34210 19916
rect 36078 19904 36084 19916
rect 36039 19876 36084 19904
rect 36078 19864 36084 19876
rect 36136 19864 36142 19916
rect 36725 19907 36783 19913
rect 36725 19873 36737 19907
rect 36771 19873 36783 19907
rect 36725 19867 36783 19873
rect 33873 19839 33931 19845
rect 33873 19805 33885 19839
rect 33919 19836 33931 19839
rect 35250 19836 35256 19848
rect 33919 19808 35256 19836
rect 33919 19805 33931 19808
rect 33873 19799 33931 19805
rect 35250 19796 35256 19808
rect 35308 19796 35314 19848
rect 36740 19836 36768 19867
rect 36814 19864 36820 19916
rect 36872 19904 36878 19916
rect 36909 19907 36967 19913
rect 36909 19904 36921 19907
rect 36872 19876 36921 19904
rect 36872 19864 36878 19876
rect 36909 19873 36921 19876
rect 36955 19873 36967 19907
rect 36909 19867 36967 19873
rect 37274 19864 37280 19916
rect 37332 19904 37338 19916
rect 37737 19907 37795 19913
rect 37737 19904 37749 19907
rect 37332 19876 37749 19904
rect 37332 19864 37338 19876
rect 37737 19873 37749 19876
rect 37783 19873 37795 19907
rect 37737 19867 37795 19873
rect 36740 19808 36952 19836
rect 36924 19780 36952 19808
rect 30466 19768 30472 19780
rect 23032 19740 28856 19768
rect 29104 19740 29776 19768
rect 29840 19740 30472 19768
rect 6328 19672 8248 19700
rect 8941 19703 8999 19709
rect 6328 19660 6334 19672
rect 8941 19669 8953 19703
rect 8987 19700 8999 19703
rect 9674 19700 9680 19712
rect 8987 19672 9680 19700
rect 8987 19669 8999 19672
rect 8941 19663 8999 19669
rect 9674 19660 9680 19672
rect 9732 19660 9738 19712
rect 12526 19700 12532 19712
rect 12487 19672 12532 19700
rect 12526 19660 12532 19672
rect 12584 19660 12590 19712
rect 13814 19660 13820 19712
rect 13872 19700 13878 19712
rect 14734 19700 14740 19712
rect 13872 19672 14740 19700
rect 13872 19660 13878 19672
rect 14734 19660 14740 19672
rect 14792 19700 14798 19712
rect 14921 19703 14979 19709
rect 14921 19700 14933 19703
rect 14792 19672 14933 19700
rect 14792 19660 14798 19672
rect 14921 19669 14933 19672
rect 14967 19669 14979 19703
rect 14921 19663 14979 19669
rect 16758 19660 16764 19712
rect 16816 19700 16822 19712
rect 17681 19703 17739 19709
rect 17681 19700 17693 19703
rect 16816 19672 17693 19700
rect 16816 19660 16822 19672
rect 17681 19669 17693 19672
rect 17727 19669 17739 19703
rect 17681 19663 17739 19669
rect 21174 19660 21180 19712
rect 21232 19700 21238 19712
rect 23032 19700 23060 19740
rect 21232 19672 23060 19700
rect 21232 19660 21238 19672
rect 25222 19660 25228 19712
rect 25280 19700 25286 19712
rect 29104 19700 29132 19740
rect 25280 19672 29132 19700
rect 29181 19703 29239 19709
rect 25280 19660 25286 19672
rect 29181 19669 29193 19703
rect 29227 19700 29239 19703
rect 29840 19700 29868 19740
rect 30466 19728 30472 19740
rect 30524 19728 30530 19780
rect 36357 19771 36415 19777
rect 36357 19737 36369 19771
rect 36403 19768 36415 19771
rect 36722 19768 36728 19780
rect 36403 19740 36728 19768
rect 36403 19737 36415 19740
rect 36357 19731 36415 19737
rect 36722 19728 36728 19740
rect 36780 19728 36786 19780
rect 36906 19728 36912 19780
rect 36964 19728 36970 19780
rect 29227 19672 29868 19700
rect 29227 19669 29239 19672
rect 29181 19663 29239 19669
rect 30650 19660 30656 19712
rect 30708 19700 30714 19712
rect 31389 19703 31447 19709
rect 31389 19700 31401 19703
rect 30708 19672 31401 19700
rect 30708 19660 30714 19672
rect 31389 19669 31401 19672
rect 31435 19669 31447 19703
rect 31389 19663 31447 19669
rect 36998 19660 37004 19712
rect 37056 19700 37062 19712
rect 37829 19703 37887 19709
rect 37829 19700 37841 19703
rect 37056 19672 37841 19700
rect 37056 19660 37062 19672
rect 37829 19669 37841 19672
rect 37875 19669 37887 19703
rect 37829 19663 37887 19669
rect 1104 19610 38824 19632
rect 1104 19558 4246 19610
rect 4298 19558 4310 19610
rect 4362 19558 4374 19610
rect 4426 19558 4438 19610
rect 4490 19558 34966 19610
rect 35018 19558 35030 19610
rect 35082 19558 35094 19610
rect 35146 19558 35158 19610
rect 35210 19558 38824 19610
rect 1104 19536 38824 19558
rect 4614 19496 4620 19508
rect 4527 19468 4620 19496
rect 4614 19456 4620 19468
rect 4672 19496 4678 19508
rect 8202 19496 8208 19508
rect 4672 19468 8208 19496
rect 4672 19456 4678 19468
rect 8202 19456 8208 19468
rect 8260 19456 8266 19508
rect 10873 19499 10931 19505
rect 10873 19465 10885 19499
rect 10919 19496 10931 19499
rect 11054 19496 11060 19508
rect 10919 19468 11060 19496
rect 10919 19465 10931 19468
rect 10873 19459 10931 19465
rect 11054 19456 11060 19468
rect 11112 19456 11118 19508
rect 14826 19456 14832 19508
rect 14884 19496 14890 19508
rect 25866 19496 25872 19508
rect 14884 19468 25872 19496
rect 14884 19456 14890 19468
rect 25866 19456 25872 19468
rect 25924 19456 25930 19508
rect 27154 19456 27160 19508
rect 27212 19496 27218 19508
rect 27985 19499 28043 19505
rect 27212 19468 27936 19496
rect 27212 19456 27218 19468
rect 3973 19431 4031 19437
rect 3973 19397 3985 19431
rect 4019 19428 4031 19431
rect 4522 19428 4528 19440
rect 4019 19400 4528 19428
rect 4019 19397 4031 19400
rect 3973 19391 4031 19397
rect 4522 19388 4528 19400
rect 4580 19428 4586 19440
rect 4706 19428 4712 19440
rect 4580 19400 4712 19428
rect 4580 19388 4586 19400
rect 4706 19388 4712 19400
rect 4764 19428 4770 19440
rect 5994 19428 6000 19440
rect 4764 19400 6000 19428
rect 4764 19388 4770 19400
rect 5994 19388 6000 19400
rect 6052 19388 6058 19440
rect 8018 19388 8024 19440
rect 8076 19428 8082 19440
rect 18966 19428 18972 19440
rect 8076 19400 18972 19428
rect 8076 19388 8082 19400
rect 18966 19388 18972 19400
rect 19024 19388 19030 19440
rect 22186 19388 22192 19440
rect 22244 19428 22250 19440
rect 22373 19431 22431 19437
rect 22373 19428 22385 19431
rect 22244 19400 22385 19428
rect 22244 19388 22250 19400
rect 22373 19397 22385 19400
rect 22419 19397 22431 19431
rect 23753 19431 23811 19437
rect 23753 19428 23765 19431
rect 22373 19391 22431 19397
rect 23032 19400 23765 19428
rect 7374 19360 7380 19372
rect 7335 19332 7380 19360
rect 7374 19320 7380 19332
rect 7432 19360 7438 19372
rect 13449 19363 13507 19369
rect 7432 19332 9168 19360
rect 7432 19320 7438 19332
rect 1394 19252 1400 19304
rect 1452 19292 1458 19304
rect 2409 19295 2467 19301
rect 2409 19292 2421 19295
rect 1452 19264 2421 19292
rect 1452 19252 1458 19264
rect 2409 19261 2421 19264
rect 2455 19261 2467 19295
rect 2409 19255 2467 19261
rect 2685 19295 2743 19301
rect 2685 19261 2697 19295
rect 2731 19292 2743 19295
rect 2958 19292 2964 19304
rect 2731 19264 2964 19292
rect 2731 19261 2743 19264
rect 2685 19255 2743 19261
rect 2958 19252 2964 19264
rect 3016 19252 3022 19304
rect 4522 19292 4528 19304
rect 4483 19264 4528 19292
rect 4522 19252 4528 19264
rect 4580 19252 4586 19304
rect 5258 19292 5264 19304
rect 5219 19264 5264 19292
rect 5258 19252 5264 19264
rect 5316 19252 5322 19304
rect 5442 19292 5448 19304
rect 5403 19264 5448 19292
rect 5442 19252 5448 19264
rect 5500 19252 5506 19304
rect 6454 19292 6460 19304
rect 5736 19264 6460 19292
rect 4062 19184 4068 19236
rect 4120 19224 4126 19236
rect 5353 19227 5411 19233
rect 4120 19196 4752 19224
rect 4120 19184 4126 19196
rect 4724 19156 4752 19196
rect 5353 19193 5365 19227
rect 5399 19224 5411 19227
rect 5736 19224 5764 19264
rect 6454 19252 6460 19264
rect 6512 19252 6518 19304
rect 7006 19292 7012 19304
rect 6967 19264 7012 19292
rect 7006 19252 7012 19264
rect 7064 19252 7070 19304
rect 7282 19292 7288 19304
rect 7243 19264 7288 19292
rect 7282 19252 7288 19264
rect 7340 19252 7346 19304
rect 7466 19252 7472 19304
rect 7524 19292 7530 19304
rect 7561 19295 7619 19301
rect 7561 19292 7573 19295
rect 7524 19264 7573 19292
rect 7524 19252 7530 19264
rect 7561 19261 7573 19264
rect 7607 19261 7619 19295
rect 7561 19255 7619 19261
rect 8297 19295 8355 19301
rect 8297 19261 8309 19295
rect 8343 19292 8355 19295
rect 8386 19292 8392 19304
rect 8343 19264 8392 19292
rect 8343 19261 8355 19264
rect 8297 19255 8355 19261
rect 8386 19252 8392 19264
rect 8444 19252 8450 19304
rect 8754 19252 8760 19304
rect 8812 19292 8818 19304
rect 9033 19295 9091 19301
rect 9033 19292 9045 19295
rect 8812 19264 9045 19292
rect 8812 19252 8818 19264
rect 9033 19261 9045 19264
rect 9079 19261 9091 19295
rect 9140 19292 9168 19332
rect 9968 19332 10732 19360
rect 9677 19295 9735 19301
rect 9677 19292 9689 19295
rect 9140 19264 9689 19292
rect 9033 19255 9091 19261
rect 9677 19261 9689 19264
rect 9723 19261 9735 19295
rect 9677 19255 9735 19261
rect 5902 19224 5908 19236
rect 5399 19196 5764 19224
rect 5863 19196 5908 19224
rect 5399 19193 5411 19196
rect 5353 19187 5411 19193
rect 5902 19184 5908 19196
rect 5960 19184 5966 19236
rect 5994 19184 6000 19236
rect 6052 19224 6058 19236
rect 7300 19224 7328 19252
rect 9968 19224 9996 19332
rect 10045 19295 10103 19301
rect 10045 19261 10057 19295
rect 10091 19261 10103 19295
rect 10594 19292 10600 19304
rect 10555 19264 10600 19292
rect 10045 19255 10103 19261
rect 6052 19196 7328 19224
rect 8128 19196 9996 19224
rect 10060 19224 10088 19255
rect 10594 19252 10600 19264
rect 10652 19252 10658 19304
rect 10704 19301 10732 19332
rect 13449 19329 13461 19363
rect 13495 19360 13507 19363
rect 13722 19360 13728 19372
rect 13495 19332 13728 19360
rect 13495 19329 13507 19332
rect 13449 19323 13507 19329
rect 13722 19320 13728 19332
rect 13780 19320 13786 19372
rect 15930 19360 15936 19372
rect 14200 19332 15792 19360
rect 15891 19332 15936 19360
rect 14200 19304 14228 19332
rect 10689 19295 10747 19301
rect 10689 19261 10701 19295
rect 10735 19261 10747 19295
rect 11606 19292 11612 19304
rect 11567 19264 11612 19292
rect 10689 19255 10747 19261
rect 11606 19252 11612 19264
rect 11664 19252 11670 19304
rect 13538 19252 13544 19304
rect 13596 19292 13602 19304
rect 13633 19295 13691 19301
rect 13633 19292 13645 19295
rect 13596 19264 13645 19292
rect 13596 19252 13602 19264
rect 13633 19261 13645 19264
rect 13679 19261 13691 19295
rect 14182 19292 14188 19304
rect 14095 19264 14188 19292
rect 13633 19255 13691 19261
rect 14182 19252 14188 19264
rect 14240 19252 14246 19304
rect 14369 19295 14427 19301
rect 14369 19261 14381 19295
rect 14415 19292 14427 19295
rect 14829 19295 14887 19301
rect 14829 19292 14841 19295
rect 14415 19264 14841 19292
rect 14415 19261 14427 19264
rect 14369 19255 14427 19261
rect 14829 19261 14841 19264
rect 14875 19261 14887 19295
rect 15194 19292 15200 19304
rect 15155 19264 15200 19292
rect 14829 19255 14887 19261
rect 15194 19252 15200 19264
rect 15252 19252 15258 19304
rect 15286 19252 15292 19304
rect 15344 19292 15350 19304
rect 15657 19295 15715 19301
rect 15657 19292 15669 19295
rect 15344 19264 15669 19292
rect 15344 19252 15350 19264
rect 15657 19261 15669 19264
rect 15703 19261 15715 19295
rect 15764 19292 15792 19332
rect 15930 19320 15936 19332
rect 15988 19320 15994 19372
rect 17310 19360 17316 19372
rect 16040 19332 17316 19360
rect 16040 19292 16068 19332
rect 17310 19320 17316 19332
rect 17368 19320 17374 19372
rect 20070 19320 20076 19372
rect 20128 19360 20134 19372
rect 20901 19363 20959 19369
rect 20901 19360 20913 19363
rect 20128 19332 20913 19360
rect 20128 19320 20134 19332
rect 20901 19329 20913 19332
rect 20947 19360 20959 19363
rect 21174 19360 21180 19372
rect 20947 19332 21180 19360
rect 20947 19329 20959 19332
rect 20901 19323 20959 19329
rect 21174 19320 21180 19332
rect 21232 19320 21238 19372
rect 21726 19320 21732 19372
rect 21784 19360 21790 19372
rect 21784 19332 22232 19360
rect 21784 19320 21790 19332
rect 16390 19292 16396 19304
rect 15764 19264 16068 19292
rect 16351 19264 16396 19292
rect 15657 19255 15715 19261
rect 16390 19252 16396 19264
rect 16448 19252 16454 19304
rect 16482 19252 16488 19304
rect 16540 19292 16546 19304
rect 17862 19292 17868 19304
rect 16540 19264 16585 19292
rect 17823 19264 17868 19292
rect 16540 19252 16546 19264
rect 17862 19252 17868 19264
rect 17920 19252 17926 19304
rect 18046 19292 18052 19304
rect 18007 19264 18052 19292
rect 18046 19252 18052 19264
rect 18104 19252 18110 19304
rect 18141 19295 18199 19301
rect 18141 19261 18153 19295
rect 18187 19292 18199 19295
rect 18230 19292 18236 19304
rect 18187 19264 18236 19292
rect 18187 19261 18199 19264
rect 18141 19255 18199 19261
rect 18230 19252 18236 19264
rect 18288 19252 18294 19304
rect 20530 19252 20536 19304
rect 20588 19292 20594 19304
rect 20993 19295 21051 19301
rect 20993 19292 21005 19295
rect 20588 19264 21005 19292
rect 20588 19252 20594 19264
rect 20993 19261 21005 19264
rect 21039 19261 21051 19295
rect 20993 19255 21051 19261
rect 21269 19295 21327 19301
rect 21269 19261 21281 19295
rect 21315 19292 21327 19295
rect 22002 19292 22008 19304
rect 21315 19264 22008 19292
rect 21315 19261 21327 19264
rect 21269 19255 21327 19261
rect 22002 19252 22008 19264
rect 22060 19252 22066 19304
rect 22204 19292 22232 19332
rect 22741 19295 22799 19301
rect 22741 19292 22753 19295
rect 22204 19264 22753 19292
rect 22741 19261 22753 19264
rect 22787 19261 22799 19295
rect 22741 19255 22799 19261
rect 16942 19224 16948 19236
rect 10060 19196 11744 19224
rect 16903 19196 16948 19224
rect 6052 19184 6058 19196
rect 8128 19156 8156 19196
rect 4724 19128 8156 19156
rect 9125 19159 9183 19165
rect 9125 19125 9137 19159
rect 9171 19156 9183 19159
rect 10226 19156 10232 19168
rect 9171 19128 10232 19156
rect 9171 19125 9183 19128
rect 9125 19119 9183 19125
rect 10226 19116 10232 19128
rect 10284 19116 10290 19168
rect 11716 19165 11744 19196
rect 16942 19184 16948 19196
rect 17000 19184 17006 19236
rect 17126 19184 17132 19236
rect 17184 19224 17190 19236
rect 18601 19227 18659 19233
rect 18601 19224 18613 19227
rect 17184 19196 18613 19224
rect 17184 19184 17190 19196
rect 18601 19193 18613 19196
rect 18647 19193 18659 19227
rect 18601 19187 18659 19193
rect 19153 19227 19211 19233
rect 19153 19193 19165 19227
rect 19199 19224 19211 19227
rect 19199 19196 20668 19224
rect 19199 19193 19211 19196
rect 19153 19187 19211 19193
rect 11701 19159 11759 19165
rect 11701 19125 11713 19159
rect 11747 19156 11759 19159
rect 14274 19156 14280 19168
rect 11747 19128 14280 19156
rect 11747 19125 11759 19128
rect 11701 19119 11759 19125
rect 14274 19116 14280 19128
rect 14332 19116 14338 19168
rect 17681 19159 17739 19165
rect 17681 19125 17693 19159
rect 17727 19156 17739 19159
rect 18966 19156 18972 19168
rect 17727 19128 18972 19156
rect 17727 19125 17739 19128
rect 17681 19119 17739 19125
rect 18966 19116 18972 19128
rect 19024 19116 19030 19168
rect 20640 19156 20668 19196
rect 22094 19184 22100 19236
rect 22152 19224 22158 19236
rect 23032 19224 23060 19400
rect 23753 19397 23765 19400
rect 23799 19397 23811 19431
rect 27908 19428 27936 19468
rect 27985 19465 27997 19499
rect 28031 19496 28043 19499
rect 28442 19496 28448 19508
rect 28031 19468 28448 19496
rect 28031 19465 28043 19468
rect 27985 19459 28043 19465
rect 28442 19456 28448 19468
rect 28500 19456 28506 19508
rect 29178 19456 29184 19508
rect 29236 19496 29242 19508
rect 32122 19496 32128 19508
rect 29236 19468 32128 19496
rect 29236 19456 29242 19468
rect 32122 19456 32128 19468
rect 32180 19456 32186 19508
rect 28994 19428 29000 19440
rect 27908 19400 29000 19428
rect 23753 19391 23811 19397
rect 28994 19388 29000 19400
rect 29052 19428 29058 19440
rect 30006 19428 30012 19440
rect 29052 19400 30012 19428
rect 29052 19388 29058 19400
rect 30006 19388 30012 19400
rect 30064 19388 30070 19440
rect 30837 19431 30895 19437
rect 30837 19397 30849 19431
rect 30883 19428 30895 19431
rect 31018 19428 31024 19440
rect 30883 19400 31024 19428
rect 30883 19397 30895 19400
rect 30837 19391 30895 19397
rect 31018 19388 31024 19400
rect 31076 19388 31082 19440
rect 26510 19320 26516 19372
rect 26568 19360 26574 19372
rect 26789 19363 26847 19369
rect 26789 19360 26801 19363
rect 26568 19332 26801 19360
rect 26568 19320 26574 19332
rect 26789 19329 26801 19332
rect 26835 19329 26847 19363
rect 26789 19323 26847 19329
rect 29086 19320 29092 19372
rect 29144 19360 29150 19372
rect 29454 19360 29460 19372
rect 29144 19332 29460 19360
rect 29144 19320 29150 19332
rect 29454 19320 29460 19332
rect 29512 19320 29518 19372
rect 29638 19320 29644 19372
rect 29696 19360 29702 19372
rect 30374 19360 30380 19372
rect 29696 19332 30380 19360
rect 29696 19320 29702 19332
rect 30374 19320 30380 19332
rect 30432 19320 30438 19372
rect 33318 19360 33324 19372
rect 33279 19332 33324 19360
rect 33318 19320 33324 19332
rect 33376 19320 33382 19372
rect 36262 19320 36268 19372
rect 36320 19360 36326 19372
rect 36449 19363 36507 19369
rect 36449 19360 36461 19363
rect 36320 19332 36461 19360
rect 36320 19320 36326 19332
rect 36449 19329 36461 19332
rect 36495 19360 36507 19363
rect 36495 19332 36584 19360
rect 36495 19329 36507 19332
rect 36449 19323 36507 19329
rect 36556 19304 36584 19332
rect 23290 19252 23296 19304
rect 23348 19292 23354 19304
rect 23661 19295 23719 19301
rect 23661 19292 23673 19295
rect 23348 19264 23673 19292
rect 23348 19252 23354 19264
rect 23661 19261 23673 19264
rect 23707 19261 23719 19295
rect 24394 19292 24400 19304
rect 24355 19264 24400 19292
rect 23661 19255 23719 19261
rect 24394 19252 24400 19264
rect 24452 19252 24458 19304
rect 24854 19292 24860 19304
rect 24815 19264 24860 19292
rect 24854 19252 24860 19264
rect 24912 19252 24918 19304
rect 25038 19292 25044 19304
rect 24999 19264 25044 19292
rect 25038 19252 25044 19264
rect 25096 19252 25102 19304
rect 25130 19252 25136 19304
rect 25188 19292 25194 19304
rect 25317 19295 25375 19301
rect 25317 19292 25329 19295
rect 25188 19264 25329 19292
rect 25188 19252 25194 19264
rect 25317 19261 25329 19264
rect 25363 19261 25375 19295
rect 26142 19292 26148 19304
rect 26103 19264 26148 19292
rect 25317 19255 25375 19261
rect 26142 19252 26148 19264
rect 26200 19252 26206 19304
rect 26878 19252 26884 19304
rect 26936 19292 26942 19304
rect 26973 19295 27031 19301
rect 26973 19292 26985 19295
rect 26936 19264 26985 19292
rect 26936 19252 26942 19264
rect 26973 19261 26985 19264
rect 27019 19261 27031 19295
rect 26973 19255 27031 19261
rect 27522 19252 27528 19304
rect 27580 19292 27586 19304
rect 27709 19295 27767 19301
rect 27580 19264 27625 19292
rect 27580 19252 27586 19264
rect 27709 19261 27721 19295
rect 27755 19292 27767 19295
rect 27890 19292 27896 19304
rect 27755 19264 27896 19292
rect 27755 19261 27767 19264
rect 27709 19255 27767 19261
rect 27890 19252 27896 19264
rect 27948 19252 27954 19304
rect 28902 19252 28908 19304
rect 28960 19292 28966 19304
rect 29273 19295 29331 19301
rect 29273 19292 29285 19295
rect 28960 19264 29285 19292
rect 28960 19252 28966 19264
rect 29273 19261 29285 19264
rect 29319 19261 29331 19295
rect 29273 19255 29331 19261
rect 29362 19252 29368 19304
rect 29420 19292 29426 19304
rect 29733 19295 29791 19301
rect 29733 19292 29745 19295
rect 29420 19264 29745 19292
rect 29420 19252 29426 19264
rect 29733 19261 29745 19264
rect 29779 19261 29791 19295
rect 29733 19255 29791 19261
rect 31021 19295 31079 19301
rect 31021 19261 31033 19295
rect 31067 19261 31079 19295
rect 31021 19255 31079 19261
rect 31389 19295 31447 19301
rect 31389 19261 31401 19295
rect 31435 19261 31447 19295
rect 31389 19255 31447 19261
rect 22152 19196 23060 19224
rect 22152 19184 22158 19196
rect 24762 19184 24768 19236
rect 24820 19224 24826 19236
rect 25056 19224 25084 19252
rect 24820 19196 25084 19224
rect 24820 19184 24826 19196
rect 27246 19184 27252 19236
rect 27304 19224 27310 19236
rect 30282 19224 30288 19236
rect 27304 19196 30288 19224
rect 27304 19184 27310 19196
rect 30282 19184 30288 19196
rect 30340 19184 30346 19236
rect 22278 19156 22284 19168
rect 20640 19128 22284 19156
rect 22278 19116 22284 19128
rect 22336 19116 22342 19168
rect 22830 19116 22836 19168
rect 22888 19156 22894 19168
rect 22925 19159 22983 19165
rect 22925 19156 22937 19159
rect 22888 19128 22937 19156
rect 22888 19116 22894 19128
rect 22925 19125 22937 19128
rect 22971 19156 22983 19159
rect 25958 19156 25964 19168
rect 22971 19128 25964 19156
rect 22971 19125 22983 19128
rect 22925 19119 22983 19125
rect 25958 19116 25964 19128
rect 26016 19116 26022 19168
rect 26234 19156 26240 19168
rect 26195 19128 26240 19156
rect 26234 19116 26240 19128
rect 26292 19116 26298 19168
rect 26970 19116 26976 19168
rect 27028 19156 27034 19168
rect 27430 19156 27436 19168
rect 27028 19128 27436 19156
rect 27028 19116 27034 19128
rect 27430 19116 27436 19128
rect 27488 19116 27494 19168
rect 27706 19116 27712 19168
rect 27764 19156 27770 19168
rect 29365 19159 29423 19165
rect 29365 19156 29377 19159
rect 27764 19128 29377 19156
rect 27764 19116 27770 19128
rect 29365 19125 29377 19128
rect 29411 19125 29423 19159
rect 29365 19119 29423 19125
rect 29730 19116 29736 19168
rect 29788 19156 29794 19168
rect 30190 19156 30196 19168
rect 29788 19128 30196 19156
rect 29788 19116 29794 19128
rect 30190 19116 30196 19128
rect 30248 19116 30254 19168
rect 31036 19156 31064 19255
rect 31404 19224 31432 19255
rect 31478 19252 31484 19304
rect 31536 19292 31542 19304
rect 31536 19264 31581 19292
rect 31536 19252 31542 19264
rect 31754 19252 31760 19304
rect 31812 19292 31818 19304
rect 32033 19295 32091 19301
rect 32033 19292 32045 19295
rect 31812 19264 32045 19292
rect 31812 19252 31818 19264
rect 32033 19261 32045 19264
rect 32079 19261 32091 19295
rect 32950 19292 32956 19304
rect 32911 19264 32956 19292
rect 32033 19255 32091 19261
rect 32950 19252 32956 19264
rect 33008 19252 33014 19304
rect 33134 19292 33140 19304
rect 33095 19264 33140 19292
rect 33134 19252 33140 19264
rect 33192 19252 33198 19304
rect 33413 19295 33471 19301
rect 33413 19261 33425 19295
rect 33459 19261 33471 19295
rect 33413 19255 33471 19261
rect 32968 19224 32996 19252
rect 31404 19196 32996 19224
rect 33042 19184 33048 19236
rect 33100 19224 33106 19236
rect 33428 19224 33456 19255
rect 33594 19252 33600 19304
rect 33652 19292 33658 19304
rect 34238 19292 34244 19304
rect 33652 19264 34244 19292
rect 33652 19252 33658 19264
rect 34238 19252 34244 19264
rect 34296 19292 34302 19304
rect 34885 19295 34943 19301
rect 34885 19292 34897 19295
rect 34296 19264 34897 19292
rect 34296 19252 34302 19264
rect 34885 19261 34897 19264
rect 34931 19261 34943 19295
rect 34885 19255 34943 19261
rect 34974 19252 34980 19304
rect 35032 19292 35038 19304
rect 35437 19295 35495 19301
rect 35437 19292 35449 19295
rect 35032 19264 35449 19292
rect 35032 19252 35038 19264
rect 35437 19261 35449 19264
rect 35483 19292 35495 19295
rect 35526 19292 35532 19304
rect 35483 19264 35532 19292
rect 35483 19261 35495 19264
rect 35437 19255 35495 19261
rect 35526 19252 35532 19264
rect 35584 19252 35590 19304
rect 36538 19252 36544 19304
rect 36596 19252 36602 19304
rect 36725 19295 36783 19301
rect 36725 19261 36737 19295
rect 36771 19292 36783 19295
rect 37366 19292 37372 19304
rect 36771 19264 37372 19292
rect 36771 19261 36783 19264
rect 36725 19255 36783 19261
rect 37366 19252 37372 19264
rect 37424 19252 37430 19304
rect 33100 19196 33456 19224
rect 33100 19184 33106 19196
rect 34698 19184 34704 19236
rect 34756 19224 34762 19236
rect 34756 19196 35112 19224
rect 34756 19184 34762 19196
rect 32766 19156 32772 19168
rect 31036 19128 32772 19156
rect 32766 19116 32772 19128
rect 32824 19116 32830 19168
rect 34790 19116 34796 19168
rect 34848 19156 34854 19168
rect 34977 19159 35035 19165
rect 34977 19156 34989 19159
rect 34848 19128 34989 19156
rect 34848 19116 34854 19128
rect 34977 19125 34989 19128
rect 35023 19125 35035 19159
rect 35084 19156 35112 19196
rect 37829 19159 37887 19165
rect 37829 19156 37841 19159
rect 35084 19128 37841 19156
rect 34977 19119 35035 19125
rect 37829 19125 37841 19128
rect 37875 19125 37887 19159
rect 37829 19119 37887 19125
rect 1104 19066 38824 19088
rect 1104 19014 19606 19066
rect 19658 19014 19670 19066
rect 19722 19014 19734 19066
rect 19786 19014 19798 19066
rect 19850 19014 38824 19066
rect 1104 18992 38824 19014
rect 3970 18912 3976 18964
rect 4028 18952 4034 18964
rect 5902 18952 5908 18964
rect 4028 18924 5908 18952
rect 4028 18912 4034 18924
rect 5902 18912 5908 18924
rect 5960 18912 5966 18964
rect 6086 18912 6092 18964
rect 6144 18952 6150 18964
rect 15470 18952 15476 18964
rect 6144 18924 15476 18952
rect 6144 18912 6150 18924
rect 15470 18912 15476 18924
rect 15528 18912 15534 18964
rect 15764 18924 17816 18952
rect 6104 18884 6132 18912
rect 7466 18884 7472 18896
rect 5092 18856 6132 18884
rect 7116 18856 7472 18884
rect 2314 18816 2320 18828
rect 2275 18788 2320 18816
rect 2314 18776 2320 18788
rect 2372 18776 2378 18828
rect 2682 18816 2688 18828
rect 2643 18788 2688 18816
rect 2682 18776 2688 18788
rect 2740 18776 2746 18828
rect 3053 18819 3111 18825
rect 3053 18785 3065 18819
rect 3099 18816 3111 18819
rect 3142 18816 3148 18828
rect 3099 18788 3148 18816
rect 3099 18785 3111 18788
rect 3053 18779 3111 18785
rect 3142 18776 3148 18788
rect 3200 18776 3206 18828
rect 3418 18816 3424 18828
rect 3379 18788 3424 18816
rect 3418 18776 3424 18788
rect 3476 18816 3482 18828
rect 5092 18825 5120 18856
rect 4065 18819 4123 18825
rect 4065 18816 4077 18819
rect 3476 18788 4077 18816
rect 3476 18776 3482 18788
rect 4065 18785 4077 18788
rect 4111 18785 4123 18819
rect 4065 18779 4123 18785
rect 5077 18819 5135 18825
rect 5077 18785 5089 18819
rect 5123 18785 5135 18819
rect 5258 18816 5264 18828
rect 5219 18788 5264 18816
rect 5077 18779 5135 18785
rect 5258 18776 5264 18788
rect 5316 18776 5322 18828
rect 5626 18776 5632 18828
rect 5684 18816 5690 18828
rect 5684 18788 5729 18816
rect 5684 18776 5690 18788
rect 5902 18776 5908 18828
rect 5960 18816 5966 18828
rect 6089 18819 6147 18825
rect 6089 18816 6101 18819
rect 5960 18788 6101 18816
rect 5960 18776 5966 18788
rect 6089 18785 6101 18788
rect 6135 18816 6147 18819
rect 6178 18816 6184 18828
rect 6135 18788 6184 18816
rect 6135 18785 6147 18788
rect 6089 18779 6147 18785
rect 6178 18776 6184 18788
rect 6236 18776 6242 18828
rect 6733 18819 6791 18825
rect 6733 18785 6745 18819
rect 6779 18816 6791 18819
rect 7006 18816 7012 18828
rect 6779 18788 7012 18816
rect 6779 18785 6791 18788
rect 6733 18779 6791 18785
rect 7006 18776 7012 18788
rect 7064 18776 7070 18828
rect 7116 18825 7144 18856
rect 7466 18844 7472 18856
rect 7524 18844 7530 18896
rect 13538 18884 13544 18896
rect 13499 18856 13544 18884
rect 13538 18844 13544 18856
rect 13596 18844 13602 18896
rect 13722 18844 13728 18896
rect 13780 18884 13786 18896
rect 14645 18887 14703 18893
rect 13780 18856 14412 18884
rect 13780 18844 13786 18856
rect 7101 18819 7159 18825
rect 7101 18785 7113 18819
rect 7147 18785 7159 18819
rect 7101 18779 7159 18785
rect 7282 18776 7288 18828
rect 7340 18816 7346 18828
rect 7377 18819 7435 18825
rect 7377 18816 7389 18819
rect 7340 18788 7389 18816
rect 7340 18776 7346 18788
rect 7377 18785 7389 18788
rect 7423 18785 7435 18819
rect 8386 18816 8392 18828
rect 8347 18788 8392 18816
rect 7377 18779 7435 18785
rect 8386 18776 8392 18788
rect 8444 18776 8450 18828
rect 8941 18819 8999 18825
rect 8941 18785 8953 18819
rect 8987 18816 8999 18819
rect 9030 18816 9036 18828
rect 8987 18788 9036 18816
rect 8987 18785 8999 18788
rect 8941 18779 8999 18785
rect 9030 18776 9036 18788
rect 9088 18776 9094 18828
rect 9674 18816 9680 18828
rect 9635 18788 9680 18816
rect 9674 18776 9680 18788
rect 9732 18776 9738 18828
rect 10226 18816 10232 18828
rect 10187 18788 10232 18816
rect 10226 18776 10232 18788
rect 10284 18776 10290 18828
rect 10781 18819 10839 18825
rect 10781 18785 10793 18819
rect 10827 18816 10839 18819
rect 10965 18819 11023 18825
rect 10965 18816 10977 18819
rect 10827 18788 10977 18816
rect 10827 18785 10839 18788
rect 10781 18779 10839 18785
rect 10965 18785 10977 18788
rect 11011 18816 11023 18819
rect 11698 18816 11704 18828
rect 11011 18788 11704 18816
rect 11011 18785 11023 18788
rect 10965 18779 11023 18785
rect 11698 18776 11704 18788
rect 11756 18776 11762 18828
rect 11882 18816 11888 18828
rect 11843 18788 11888 18816
rect 11882 18776 11888 18788
rect 11940 18776 11946 18828
rect 12161 18819 12219 18825
rect 12161 18785 12173 18819
rect 12207 18816 12219 18819
rect 12526 18816 12532 18828
rect 12207 18788 12532 18816
rect 12207 18785 12219 18788
rect 12161 18779 12219 18785
rect 12526 18776 12532 18788
rect 12584 18776 12590 18828
rect 14001 18819 14059 18825
rect 14001 18785 14013 18819
rect 14047 18816 14059 18819
rect 14093 18819 14151 18825
rect 14093 18816 14105 18819
rect 14047 18788 14105 18816
rect 14047 18785 14059 18788
rect 14001 18779 14059 18785
rect 14093 18785 14105 18788
rect 14139 18785 14151 18819
rect 14274 18816 14280 18828
rect 14235 18788 14280 18816
rect 14093 18779 14151 18785
rect 14274 18776 14280 18788
rect 14332 18776 14338 18828
rect 14384 18816 14412 18856
rect 14645 18853 14657 18887
rect 14691 18884 14703 18887
rect 15286 18884 15292 18896
rect 14691 18856 15292 18884
rect 14691 18853 14703 18856
rect 14645 18847 14703 18853
rect 15286 18844 15292 18856
rect 15344 18844 15350 18896
rect 15473 18819 15531 18825
rect 15473 18816 15485 18819
rect 14384 18788 15485 18816
rect 15473 18785 15485 18788
rect 15519 18816 15531 18819
rect 15764 18816 15792 18924
rect 16758 18884 16764 18896
rect 15856 18856 16764 18884
rect 15856 18825 15884 18856
rect 16758 18844 16764 18856
rect 16816 18844 16822 18896
rect 17788 18884 17816 18924
rect 17954 18912 17960 18964
rect 18012 18952 18018 18964
rect 18233 18955 18291 18961
rect 18233 18952 18245 18955
rect 18012 18924 18245 18952
rect 18012 18912 18018 18924
rect 18233 18921 18245 18924
rect 18279 18921 18291 18955
rect 22186 18952 22192 18964
rect 18233 18915 18291 18921
rect 20916 18924 22192 18952
rect 19978 18884 19984 18896
rect 17788 18856 19984 18884
rect 19978 18844 19984 18856
rect 20036 18844 20042 18896
rect 15519 18788 15792 18816
rect 15841 18819 15899 18825
rect 15519 18785 15531 18788
rect 15473 18779 15531 18785
rect 15841 18785 15853 18819
rect 15887 18785 15899 18819
rect 15841 18779 15899 18785
rect 16022 18776 16028 18828
rect 16080 18816 16086 18828
rect 16117 18819 16175 18825
rect 16117 18816 16129 18819
rect 16080 18788 16129 18816
rect 16080 18776 16086 18788
rect 16117 18785 16129 18788
rect 16163 18785 16175 18819
rect 17126 18816 17132 18828
rect 17087 18788 17132 18816
rect 16117 18779 16175 18785
rect 17126 18776 17132 18788
rect 17184 18776 17190 18828
rect 18874 18776 18880 18828
rect 18932 18816 18938 18828
rect 19061 18819 19119 18825
rect 19061 18816 19073 18819
rect 18932 18788 19073 18816
rect 18932 18776 18938 18788
rect 19061 18785 19073 18788
rect 19107 18785 19119 18819
rect 19702 18816 19708 18828
rect 19663 18788 19708 18816
rect 19061 18779 19119 18785
rect 19702 18776 19708 18788
rect 19760 18776 19766 18828
rect 20257 18819 20315 18825
rect 20257 18785 20269 18819
rect 20303 18816 20315 18819
rect 20714 18816 20720 18828
rect 20303 18788 20720 18816
rect 20303 18785 20315 18788
rect 20257 18779 20315 18785
rect 20714 18776 20720 18788
rect 20772 18776 20778 18828
rect 20916 18825 20944 18924
rect 22186 18912 22192 18924
rect 22244 18912 22250 18964
rect 22278 18912 22284 18964
rect 22336 18952 22342 18964
rect 22336 18924 32904 18952
rect 22336 18912 22342 18924
rect 20990 18844 20996 18896
rect 21048 18884 21054 18896
rect 24578 18884 24584 18896
rect 21048 18856 21956 18884
rect 24491 18856 24584 18884
rect 21048 18844 21054 18856
rect 21928 18828 21956 18856
rect 20901 18819 20959 18825
rect 20901 18785 20913 18819
rect 20947 18785 20959 18819
rect 20901 18779 20959 18785
rect 21082 18776 21088 18828
rect 21140 18816 21146 18828
rect 21542 18816 21548 18828
rect 21140 18788 21548 18816
rect 21140 18776 21146 18788
rect 21542 18776 21548 18788
rect 21600 18776 21606 18828
rect 21910 18776 21916 18828
rect 21968 18816 21974 18828
rect 22373 18819 22431 18825
rect 22373 18816 22385 18819
rect 21968 18788 22385 18816
rect 21968 18776 21974 18788
rect 22373 18785 22385 18788
rect 22419 18816 22431 18819
rect 23658 18816 23664 18828
rect 22419 18788 23664 18816
rect 22419 18785 22431 18788
rect 22373 18779 22431 18785
rect 23658 18776 23664 18788
rect 23716 18776 23722 18828
rect 24029 18819 24087 18825
rect 24029 18785 24041 18819
rect 24075 18816 24087 18819
rect 24394 18816 24400 18828
rect 24075 18788 24400 18816
rect 24075 18785 24087 18788
rect 24029 18779 24087 18785
rect 24394 18776 24400 18788
rect 24452 18776 24458 18828
rect 24504 18825 24532 18856
rect 24578 18844 24584 18856
rect 24636 18884 24642 18896
rect 24854 18884 24860 18896
rect 24636 18856 24860 18884
rect 24636 18844 24642 18856
rect 24854 18844 24860 18856
rect 24912 18884 24918 18896
rect 26050 18884 26056 18896
rect 24912 18856 26056 18884
rect 24912 18844 24918 18856
rect 26050 18844 26056 18856
rect 26108 18844 26114 18896
rect 28813 18887 28871 18893
rect 28813 18853 28825 18887
rect 28859 18884 28871 18887
rect 29362 18884 29368 18896
rect 28859 18856 29368 18884
rect 28859 18853 28871 18856
rect 28813 18847 28871 18853
rect 24489 18819 24547 18825
rect 24489 18785 24501 18819
rect 24535 18785 24547 18819
rect 24762 18816 24768 18828
rect 24723 18788 24768 18816
rect 24489 18779 24547 18785
rect 24762 18776 24768 18788
rect 24820 18776 24826 18828
rect 25130 18816 25136 18828
rect 25091 18788 25136 18816
rect 25130 18776 25136 18788
rect 25188 18776 25194 18828
rect 25685 18819 25743 18825
rect 25685 18785 25697 18819
rect 25731 18816 25743 18819
rect 25866 18816 25872 18828
rect 25731 18788 25872 18816
rect 25731 18785 25743 18788
rect 25685 18779 25743 18785
rect 25866 18776 25872 18788
rect 25924 18776 25930 18828
rect 26513 18819 26571 18825
rect 26513 18785 26525 18819
rect 26559 18816 26571 18819
rect 28828 18816 28856 18847
rect 29362 18844 29368 18856
rect 29420 18844 29426 18896
rect 32876 18884 32904 18924
rect 32950 18912 32956 18964
rect 33008 18952 33014 18964
rect 37829 18955 37887 18961
rect 37829 18952 37841 18955
rect 33008 18924 37841 18952
rect 33008 18912 33014 18924
rect 37829 18921 37841 18924
rect 37875 18921 37887 18955
rect 37829 18915 37887 18921
rect 30208 18856 32352 18884
rect 32876 18856 32996 18884
rect 30208 18828 30236 18856
rect 26559 18788 28856 18816
rect 26559 18785 26571 18788
rect 26513 18779 26571 18785
rect 28994 18776 29000 18828
rect 29052 18816 29058 18828
rect 29273 18819 29331 18825
rect 29273 18816 29285 18819
rect 29052 18788 29285 18816
rect 29052 18776 29058 18788
rect 29273 18785 29285 18788
rect 29319 18785 29331 18819
rect 29273 18779 29331 18785
rect 30190 18776 30196 18828
rect 30248 18776 30254 18828
rect 31294 18776 31300 18828
rect 31352 18816 31358 18828
rect 31389 18819 31447 18825
rect 31389 18816 31401 18819
rect 31352 18788 31401 18816
rect 31352 18776 31358 18788
rect 31389 18785 31401 18788
rect 31435 18816 31447 18819
rect 31478 18816 31484 18828
rect 31435 18788 31484 18816
rect 31435 18785 31447 18788
rect 31389 18779 31447 18785
rect 31478 18776 31484 18788
rect 31536 18776 31542 18828
rect 32324 18816 32352 18856
rect 32861 18819 32919 18825
rect 32861 18816 32873 18819
rect 32324 18788 32873 18816
rect 32861 18785 32873 18788
rect 32907 18785 32919 18819
rect 32861 18779 32919 18785
rect 2866 18748 2872 18760
rect 2827 18720 2872 18748
rect 2866 18708 2872 18720
rect 2924 18708 2930 18760
rect 10594 18708 10600 18760
rect 10652 18748 10658 18760
rect 10873 18751 10931 18757
rect 10873 18748 10885 18751
rect 10652 18720 10885 18748
rect 10652 18708 10658 18720
rect 10873 18717 10885 18720
rect 10919 18748 10931 18751
rect 11238 18748 11244 18760
rect 10919 18720 11244 18748
rect 10919 18717 10931 18720
rect 10873 18711 10931 18717
rect 11238 18708 11244 18720
rect 11296 18708 11302 18760
rect 16040 18748 16068 18776
rect 15488 18720 16068 18748
rect 16853 18751 16911 18757
rect 4157 18683 4215 18689
rect 4157 18649 4169 18683
rect 4203 18680 4215 18683
rect 4614 18680 4620 18692
rect 4203 18652 4620 18680
rect 4203 18649 4215 18652
rect 4157 18643 4215 18649
rect 4614 18640 4620 18652
rect 4672 18680 4678 18692
rect 11330 18680 11336 18692
rect 4672 18652 11336 18680
rect 4672 18640 4678 18652
rect 11330 18640 11336 18652
rect 11388 18640 11394 18692
rect 13906 18640 13912 18692
rect 13964 18680 13970 18692
rect 14001 18683 14059 18689
rect 14001 18680 14013 18683
rect 13964 18652 14013 18680
rect 13964 18640 13970 18652
rect 14001 18649 14013 18652
rect 14047 18680 14059 18683
rect 15488 18680 15516 18720
rect 16853 18717 16865 18751
rect 16899 18748 16911 18751
rect 18782 18748 18788 18760
rect 16899 18720 18788 18748
rect 16899 18717 16911 18720
rect 16853 18711 16911 18717
rect 18782 18708 18788 18720
rect 18840 18708 18846 18760
rect 18969 18751 19027 18757
rect 18969 18717 18981 18751
rect 19015 18717 19027 18751
rect 18969 18711 19027 18717
rect 14047 18652 15516 18680
rect 14047 18649 14059 18652
rect 14001 18643 14059 18649
rect 15562 18640 15568 18692
rect 15620 18680 15626 18692
rect 16117 18683 16175 18689
rect 16117 18680 16129 18683
rect 15620 18652 16129 18680
rect 15620 18640 15626 18652
rect 16117 18649 16129 18652
rect 16163 18649 16175 18683
rect 16117 18643 16175 18649
rect 17862 18640 17868 18692
rect 17920 18680 17926 18692
rect 18984 18680 19012 18711
rect 19242 18708 19248 18760
rect 19300 18748 19306 18760
rect 19613 18751 19671 18757
rect 19613 18748 19625 18751
rect 19300 18720 19625 18748
rect 19300 18708 19306 18720
rect 19613 18717 19625 18720
rect 19659 18717 19671 18751
rect 22094 18748 22100 18760
rect 19613 18711 19671 18717
rect 20456 18720 22100 18748
rect 17920 18652 19012 18680
rect 17920 18640 17926 18652
rect 19058 18640 19064 18692
rect 19116 18680 19122 18692
rect 20346 18680 20352 18692
rect 19116 18652 20352 18680
rect 19116 18640 19122 18652
rect 20346 18640 20352 18652
rect 20404 18640 20410 18692
rect 20456 18689 20484 18720
rect 22094 18708 22100 18720
rect 22152 18748 22158 18760
rect 22281 18751 22339 18757
rect 22281 18748 22293 18751
rect 22152 18720 22293 18748
rect 22152 18708 22158 18720
rect 22281 18717 22293 18720
rect 22327 18717 22339 18751
rect 22281 18711 22339 18717
rect 22649 18751 22707 18757
rect 22649 18717 22661 18751
rect 22695 18748 22707 18751
rect 26970 18748 26976 18760
rect 22695 18720 26976 18748
rect 22695 18717 22707 18720
rect 22649 18711 22707 18717
rect 26970 18708 26976 18720
rect 27028 18708 27034 18760
rect 27154 18748 27160 18760
rect 27115 18720 27160 18748
rect 27154 18708 27160 18720
rect 27212 18708 27218 18760
rect 27433 18751 27491 18757
rect 27433 18717 27445 18751
rect 27479 18748 27491 18751
rect 28350 18748 28356 18760
rect 27479 18720 28356 18748
rect 27479 18717 27491 18720
rect 27433 18711 27491 18717
rect 28350 18708 28356 18720
rect 28408 18708 28414 18760
rect 29546 18748 29552 18760
rect 29507 18720 29552 18748
rect 29546 18708 29552 18720
rect 29604 18708 29610 18760
rect 29638 18708 29644 18760
rect 29696 18748 29702 18760
rect 32968 18748 32996 18856
rect 33244 18856 33824 18884
rect 33244 18825 33272 18856
rect 33796 18828 33824 18856
rect 34238 18844 34244 18896
rect 34296 18884 34302 18896
rect 34296 18856 35572 18884
rect 34296 18844 34302 18856
rect 33229 18819 33287 18825
rect 33229 18785 33241 18819
rect 33275 18785 33287 18819
rect 33229 18779 33287 18785
rect 33318 18776 33324 18828
rect 33376 18816 33382 18828
rect 33376 18788 33421 18816
rect 33376 18776 33382 18788
rect 33778 18776 33784 18828
rect 33836 18816 33842 18828
rect 33873 18819 33931 18825
rect 33873 18816 33885 18819
rect 33836 18788 33885 18816
rect 33836 18776 33842 18788
rect 33873 18785 33885 18788
rect 33919 18785 33931 18819
rect 33873 18779 33931 18785
rect 34425 18819 34483 18825
rect 34425 18785 34437 18819
rect 34471 18816 34483 18819
rect 34974 18816 34980 18828
rect 34471 18788 34836 18816
rect 34935 18788 34980 18816
rect 34471 18785 34483 18788
rect 34425 18779 34483 18785
rect 34146 18748 34152 18760
rect 29696 18720 31524 18748
rect 32968 18720 34152 18748
rect 29696 18708 29702 18720
rect 20441 18683 20499 18689
rect 20441 18649 20453 18683
rect 20487 18649 20499 18683
rect 23290 18680 23296 18692
rect 23251 18652 23296 18680
rect 20441 18643 20499 18649
rect 23290 18640 23296 18652
rect 23348 18640 23354 18692
rect 23385 18683 23443 18689
rect 23385 18649 23397 18683
rect 23431 18680 23443 18683
rect 23566 18680 23572 18692
rect 23431 18652 23572 18680
rect 23431 18649 23443 18652
rect 23385 18643 23443 18649
rect 23566 18640 23572 18652
rect 23624 18640 23630 18692
rect 30282 18640 30288 18692
rect 30340 18680 30346 18692
rect 31496 18689 31524 18720
rect 34146 18708 34152 18720
rect 34204 18708 34210 18760
rect 34514 18748 34520 18760
rect 34475 18720 34520 18748
rect 34514 18708 34520 18720
rect 34572 18708 34578 18760
rect 31481 18683 31539 18689
rect 30340 18652 30788 18680
rect 30340 18640 30346 18652
rect 5626 18572 5632 18624
rect 5684 18612 5690 18624
rect 6181 18615 6239 18621
rect 6181 18612 6193 18615
rect 5684 18584 6193 18612
rect 5684 18572 5690 18584
rect 6181 18581 6193 18584
rect 6227 18581 6239 18615
rect 6181 18575 6239 18581
rect 7466 18572 7472 18624
rect 7524 18612 7530 18624
rect 8297 18615 8355 18621
rect 8297 18612 8309 18615
rect 7524 18584 8309 18612
rect 7524 18572 7530 18584
rect 8297 18581 8309 18584
rect 8343 18581 8355 18615
rect 9766 18612 9772 18624
rect 9727 18584 9772 18612
rect 8297 18575 8355 18581
rect 9766 18572 9772 18584
rect 9824 18572 9830 18624
rect 11146 18612 11152 18624
rect 11107 18584 11152 18612
rect 11146 18572 11152 18584
rect 11204 18572 11210 18624
rect 18598 18572 18604 18624
rect 18656 18612 18662 18624
rect 19245 18615 19303 18621
rect 19245 18612 19257 18615
rect 18656 18584 19257 18612
rect 18656 18572 18662 18584
rect 19245 18581 19257 18584
rect 19291 18581 19303 18615
rect 19886 18612 19892 18624
rect 19847 18584 19892 18612
rect 19245 18575 19303 18581
rect 19886 18572 19892 18584
rect 19944 18572 19950 18624
rect 23198 18572 23204 18624
rect 23256 18612 23262 18624
rect 25869 18615 25927 18621
rect 25869 18612 25881 18615
rect 23256 18584 25881 18612
rect 23256 18572 23262 18584
rect 25869 18581 25881 18584
rect 25915 18581 25927 18615
rect 25869 18575 25927 18581
rect 26605 18615 26663 18621
rect 26605 18581 26617 18615
rect 26651 18612 26663 18615
rect 27522 18612 27528 18624
rect 26651 18584 27528 18612
rect 26651 18581 26663 18584
rect 26605 18575 26663 18581
rect 27522 18572 27528 18584
rect 27580 18572 27586 18624
rect 28534 18572 28540 18624
rect 28592 18612 28598 18624
rect 28902 18612 28908 18624
rect 28592 18584 28908 18612
rect 28592 18572 28598 18584
rect 28902 18572 28908 18584
rect 28960 18612 28966 18624
rect 30653 18615 30711 18621
rect 30653 18612 30665 18615
rect 28960 18584 30665 18612
rect 28960 18572 28966 18584
rect 30653 18581 30665 18584
rect 30699 18581 30711 18615
rect 30760 18612 30788 18652
rect 31481 18649 31493 18683
rect 31527 18649 31539 18683
rect 31481 18643 31539 18649
rect 32677 18683 32735 18689
rect 32677 18649 32689 18683
rect 32723 18680 32735 18683
rect 34698 18680 34704 18692
rect 32723 18652 34704 18680
rect 32723 18649 32735 18652
rect 32677 18643 32735 18649
rect 34698 18640 34704 18652
rect 34756 18640 34762 18692
rect 34808 18680 34836 18788
rect 34974 18776 34980 18788
rect 35032 18776 35038 18828
rect 35345 18819 35403 18825
rect 35345 18785 35357 18819
rect 35391 18816 35403 18819
rect 35434 18816 35440 18828
rect 35391 18788 35440 18816
rect 35391 18785 35403 18788
rect 35345 18779 35403 18785
rect 35434 18776 35440 18788
rect 35492 18776 35498 18828
rect 35544 18825 35572 18856
rect 35529 18819 35587 18825
rect 35529 18785 35541 18819
rect 35575 18785 35587 18819
rect 36446 18816 36452 18828
rect 36407 18788 36452 18816
rect 35529 18779 35587 18785
rect 36446 18776 36452 18788
rect 36504 18776 36510 18828
rect 36998 18816 37004 18828
rect 36911 18788 37004 18816
rect 36998 18776 37004 18788
rect 37056 18776 37062 18828
rect 37737 18819 37795 18825
rect 37737 18785 37749 18819
rect 37783 18785 37795 18819
rect 37737 18779 37795 18785
rect 36262 18708 36268 18760
rect 36320 18748 36326 18760
rect 37016 18748 37044 18776
rect 36320 18720 37044 18748
rect 36320 18708 36326 18720
rect 35802 18680 35808 18692
rect 34808 18652 35808 18680
rect 35802 18640 35808 18652
rect 35860 18680 35866 18692
rect 37752 18680 37780 18779
rect 35860 18652 37780 18680
rect 35860 18640 35866 18652
rect 35526 18612 35532 18624
rect 30760 18584 35532 18612
rect 30653 18575 30711 18581
rect 35526 18572 35532 18584
rect 35584 18572 35590 18624
rect 35986 18572 35992 18624
rect 36044 18612 36050 18624
rect 36541 18615 36599 18621
rect 36541 18612 36553 18615
rect 36044 18584 36553 18612
rect 36044 18572 36050 18584
rect 36541 18581 36553 18584
rect 36587 18581 36599 18615
rect 36541 18575 36599 18581
rect 1104 18522 38824 18544
rect 1104 18470 4246 18522
rect 4298 18470 4310 18522
rect 4362 18470 4374 18522
rect 4426 18470 4438 18522
rect 4490 18470 34966 18522
rect 35018 18470 35030 18522
rect 35082 18470 35094 18522
rect 35146 18470 35158 18522
rect 35210 18470 38824 18522
rect 1104 18448 38824 18470
rect 2682 18368 2688 18420
rect 2740 18408 2746 18420
rect 2777 18411 2835 18417
rect 2777 18408 2789 18411
rect 2740 18380 2789 18408
rect 2740 18368 2746 18380
rect 2777 18377 2789 18380
rect 2823 18377 2835 18411
rect 5442 18408 5448 18420
rect 5403 18380 5448 18408
rect 2777 18371 2835 18377
rect 2792 18340 2820 18371
rect 5442 18368 5448 18380
rect 5500 18368 5506 18420
rect 6086 18408 6092 18420
rect 6047 18380 6092 18408
rect 6086 18368 6092 18380
rect 6144 18368 6150 18420
rect 6178 18368 6184 18420
rect 6236 18408 6242 18420
rect 7561 18411 7619 18417
rect 7561 18408 7573 18411
rect 6236 18380 7573 18408
rect 6236 18368 6242 18380
rect 7561 18377 7573 18380
rect 7607 18377 7619 18411
rect 7561 18371 7619 18377
rect 9030 18368 9036 18420
rect 9088 18408 9094 18420
rect 9677 18411 9735 18417
rect 9677 18408 9689 18411
rect 9088 18380 9689 18408
rect 9088 18368 9094 18380
rect 9677 18377 9689 18380
rect 9723 18408 9735 18411
rect 11606 18408 11612 18420
rect 9723 18380 11612 18408
rect 9723 18377 9735 18380
rect 9677 18371 9735 18377
rect 11606 18368 11612 18380
rect 11664 18368 11670 18420
rect 11793 18411 11851 18417
rect 11793 18377 11805 18411
rect 11839 18408 11851 18411
rect 12342 18408 12348 18420
rect 11839 18380 12348 18408
rect 11839 18377 11851 18380
rect 11793 18371 11851 18377
rect 12342 18368 12348 18380
rect 12400 18368 12406 18420
rect 12526 18368 12532 18420
rect 12584 18408 12590 18420
rect 12713 18411 12771 18417
rect 12713 18408 12725 18411
rect 12584 18380 12725 18408
rect 12584 18368 12590 18380
rect 12713 18377 12725 18380
rect 12759 18377 12771 18411
rect 12713 18371 12771 18377
rect 16390 18368 16396 18420
rect 16448 18408 16454 18420
rect 19058 18408 19064 18420
rect 16448 18380 19064 18408
rect 16448 18368 16454 18380
rect 19058 18368 19064 18380
rect 19116 18368 19122 18420
rect 19702 18408 19708 18420
rect 19663 18380 19708 18408
rect 19702 18368 19708 18380
rect 19760 18368 19766 18420
rect 22462 18368 22468 18420
rect 22520 18408 22526 18420
rect 23198 18408 23204 18420
rect 22520 18380 23204 18408
rect 22520 18368 22526 18380
rect 23198 18368 23204 18380
rect 23256 18368 23262 18420
rect 26973 18411 27031 18417
rect 26973 18377 26985 18411
rect 27019 18408 27031 18411
rect 27246 18408 27252 18420
rect 27019 18380 27252 18408
rect 27019 18377 27031 18380
rect 26973 18371 27031 18377
rect 27246 18368 27252 18380
rect 27304 18368 27310 18420
rect 27338 18368 27344 18420
rect 27396 18408 27402 18420
rect 36446 18408 36452 18420
rect 27396 18380 36452 18408
rect 27396 18368 27402 18380
rect 36446 18368 36452 18380
rect 36504 18408 36510 18420
rect 37734 18408 37740 18420
rect 36504 18380 37740 18408
rect 36504 18368 36510 18380
rect 37734 18368 37740 18380
rect 37792 18368 37798 18420
rect 2792 18312 5396 18340
rect 2314 18232 2320 18284
rect 2372 18272 2378 18284
rect 2372 18244 5304 18272
rect 2372 18232 2378 18244
rect 1394 18204 1400 18216
rect 1355 18176 1400 18204
rect 1394 18164 1400 18176
rect 1452 18164 1458 18216
rect 1673 18207 1731 18213
rect 1673 18173 1685 18207
rect 1719 18204 1731 18207
rect 3970 18204 3976 18216
rect 1719 18176 3976 18204
rect 1719 18173 1731 18176
rect 1673 18167 1731 18173
rect 3970 18164 3976 18176
rect 4028 18164 4034 18216
rect 4080 18213 4108 18244
rect 4065 18207 4123 18213
rect 4065 18173 4077 18207
rect 4111 18173 4123 18207
rect 4706 18204 4712 18216
rect 4667 18176 4712 18204
rect 4065 18167 4123 18173
rect 4706 18164 4712 18176
rect 4764 18164 4770 18216
rect 5077 18207 5135 18213
rect 5077 18173 5089 18207
rect 5123 18173 5135 18207
rect 5077 18167 5135 18173
rect 5092 18068 5120 18167
rect 5276 18136 5304 18244
rect 5368 18213 5396 18312
rect 19978 18300 19984 18352
rect 20036 18340 20042 18352
rect 20036 18312 25728 18340
rect 20036 18300 20042 18312
rect 10505 18275 10563 18281
rect 10505 18241 10517 18275
rect 10551 18272 10563 18275
rect 11146 18272 11152 18284
rect 10551 18244 11152 18272
rect 10551 18241 10563 18244
rect 10505 18235 10563 18241
rect 11146 18232 11152 18244
rect 11204 18232 11210 18284
rect 11330 18232 11336 18284
rect 11388 18272 11394 18284
rect 14461 18275 14519 18281
rect 11388 18244 14136 18272
rect 11388 18232 11394 18244
rect 5353 18207 5411 18213
rect 5353 18173 5365 18207
rect 5399 18204 5411 18207
rect 5997 18207 6055 18213
rect 5997 18204 6009 18207
rect 5399 18176 6009 18204
rect 5399 18173 5411 18176
rect 5353 18167 5411 18173
rect 5997 18173 6009 18176
rect 6043 18173 6055 18207
rect 5997 18167 6055 18173
rect 6270 18164 6276 18216
rect 6328 18204 6334 18216
rect 6825 18207 6883 18213
rect 6825 18204 6837 18207
rect 6328 18176 6837 18204
rect 6328 18164 6334 18176
rect 6825 18173 6837 18176
rect 6871 18173 6883 18207
rect 7466 18204 7472 18216
rect 7427 18176 7472 18204
rect 6825 18167 6883 18173
rect 7466 18164 7472 18176
rect 7524 18164 7530 18216
rect 7742 18164 7748 18216
rect 7800 18204 7806 18216
rect 8113 18207 8171 18213
rect 8113 18204 8125 18207
rect 7800 18176 8125 18204
rect 7800 18164 7806 18176
rect 8113 18173 8125 18176
rect 8159 18173 8171 18207
rect 8386 18204 8392 18216
rect 8347 18176 8392 18204
rect 8113 18167 8171 18173
rect 8386 18164 8392 18176
rect 8444 18164 8450 18216
rect 10134 18164 10140 18216
rect 10192 18204 10198 18216
rect 10229 18207 10287 18213
rect 10229 18204 10241 18207
rect 10192 18176 10241 18204
rect 10192 18164 10198 18176
rect 10229 18173 10241 18176
rect 10275 18173 10287 18207
rect 12434 18204 12440 18216
rect 12395 18176 12440 18204
rect 10229 18167 10287 18173
rect 12434 18164 12440 18176
rect 12492 18164 12498 18216
rect 12618 18213 12624 18216
rect 12570 18207 12624 18213
rect 12570 18173 12582 18207
rect 12616 18173 12624 18207
rect 12570 18167 12624 18173
rect 12618 18164 12624 18167
rect 12676 18164 12682 18216
rect 13814 18204 13820 18216
rect 13775 18176 13820 18204
rect 13814 18164 13820 18176
rect 13872 18164 13878 18216
rect 13906 18164 13912 18216
rect 13964 18204 13970 18216
rect 14108 18213 14136 18244
rect 14461 18241 14473 18275
rect 14507 18272 14519 18275
rect 16114 18272 16120 18284
rect 14507 18244 16120 18272
rect 14507 18241 14519 18244
rect 14461 18235 14519 18241
rect 16114 18232 16120 18244
rect 16172 18232 16178 18284
rect 18598 18272 18604 18284
rect 18559 18244 18604 18272
rect 18598 18232 18604 18244
rect 18656 18232 18662 18284
rect 18782 18232 18788 18284
rect 18840 18232 18846 18284
rect 20901 18275 20959 18281
rect 20901 18241 20913 18275
rect 20947 18272 20959 18275
rect 20990 18272 20996 18284
rect 20947 18244 20996 18272
rect 20947 18241 20959 18244
rect 20901 18235 20959 18241
rect 20990 18232 20996 18244
rect 21048 18232 21054 18284
rect 22097 18275 22155 18281
rect 22097 18241 22109 18275
rect 22143 18272 22155 18275
rect 23198 18272 23204 18284
rect 22143 18244 23204 18272
rect 22143 18241 22155 18244
rect 22097 18235 22155 18241
rect 23198 18232 23204 18244
rect 23256 18232 23262 18284
rect 14093 18207 14151 18213
rect 13964 18176 14009 18204
rect 13964 18164 13970 18176
rect 14093 18173 14105 18207
rect 14139 18173 14151 18207
rect 14093 18167 14151 18173
rect 14550 18164 14556 18216
rect 14608 18204 14614 18216
rect 14921 18207 14979 18213
rect 14921 18204 14933 18207
rect 14608 18176 14933 18204
rect 14608 18164 14614 18176
rect 14921 18173 14933 18176
rect 14967 18173 14979 18207
rect 14921 18167 14979 18173
rect 15197 18207 15255 18213
rect 15197 18173 15209 18207
rect 15243 18204 15255 18207
rect 16942 18204 16948 18216
rect 15243 18176 16948 18204
rect 15243 18173 15255 18176
rect 15197 18167 15255 18173
rect 16942 18164 16948 18176
rect 17000 18164 17006 18216
rect 17126 18164 17132 18216
rect 17184 18204 17190 18216
rect 17221 18207 17279 18213
rect 17221 18204 17233 18207
rect 17184 18176 17233 18204
rect 17184 18164 17190 18176
rect 17221 18173 17233 18176
rect 17267 18173 17279 18207
rect 17221 18167 17279 18173
rect 18325 18207 18383 18213
rect 18325 18173 18337 18207
rect 18371 18204 18383 18207
rect 18800 18204 18828 18232
rect 18371 18176 18828 18204
rect 18371 18173 18383 18176
rect 18325 18167 18383 18173
rect 18966 18164 18972 18216
rect 19024 18204 19030 18216
rect 20625 18207 20683 18213
rect 20625 18204 20637 18207
rect 19024 18176 20637 18204
rect 19024 18164 19030 18176
rect 20625 18173 20637 18176
rect 20671 18173 20683 18207
rect 20625 18167 20683 18173
rect 20806 18164 20812 18216
rect 20864 18204 20870 18216
rect 21637 18207 21695 18213
rect 21637 18204 21649 18207
rect 20864 18176 21649 18204
rect 20864 18164 20870 18176
rect 21637 18173 21649 18176
rect 21683 18173 21695 18207
rect 21637 18167 21695 18173
rect 22278 18164 22284 18216
rect 22336 18204 22342 18216
rect 22557 18207 22615 18213
rect 22557 18204 22569 18207
rect 22336 18176 22569 18204
rect 22336 18164 22342 18176
rect 22557 18173 22569 18176
rect 22603 18204 22615 18207
rect 22738 18204 22744 18216
rect 22603 18176 22744 18204
rect 22603 18173 22615 18176
rect 22557 18167 22615 18173
rect 22738 18164 22744 18176
rect 22796 18164 22802 18216
rect 22922 18204 22928 18216
rect 22883 18176 22928 18204
rect 22922 18164 22928 18176
rect 22980 18164 22986 18216
rect 23014 18164 23020 18216
rect 23072 18204 23078 18216
rect 23658 18204 23664 18216
rect 23072 18176 23117 18204
rect 23619 18176 23664 18204
rect 23072 18164 23078 18176
rect 23658 18164 23664 18176
rect 23716 18164 23722 18216
rect 24397 18207 24455 18213
rect 24397 18173 24409 18207
rect 24443 18173 24455 18207
rect 25498 18204 25504 18216
rect 25459 18176 25504 18204
rect 24397 18167 24455 18173
rect 5902 18136 5908 18148
rect 5276 18108 5908 18136
rect 5902 18096 5908 18108
rect 5960 18096 5966 18148
rect 6288 18068 6316 18164
rect 11238 18096 11244 18148
rect 11296 18136 11302 18148
rect 16577 18139 16635 18145
rect 11296 18108 15056 18136
rect 11296 18096 11302 18108
rect 6914 18068 6920 18080
rect 5092 18040 6316 18068
rect 6875 18040 6920 18068
rect 6914 18028 6920 18040
rect 6972 18028 6978 18080
rect 12710 18028 12716 18080
rect 12768 18068 12774 18080
rect 13633 18071 13691 18077
rect 13633 18068 13645 18071
rect 12768 18040 13645 18068
rect 12768 18028 12774 18040
rect 13633 18037 13645 18040
rect 13679 18037 13691 18071
rect 15028 18068 15056 18108
rect 16577 18105 16589 18139
rect 16623 18136 16635 18139
rect 17770 18136 17776 18148
rect 16623 18108 17776 18136
rect 16623 18105 16635 18108
rect 16577 18099 16635 18105
rect 17770 18096 17776 18108
rect 17828 18096 17834 18148
rect 21269 18139 21327 18145
rect 21269 18105 21281 18139
rect 21315 18136 21327 18139
rect 22462 18136 22468 18148
rect 21315 18108 22468 18136
rect 21315 18105 21327 18108
rect 21269 18099 21327 18105
rect 22462 18096 22468 18108
rect 22520 18096 22526 18148
rect 22646 18096 22652 18148
rect 22704 18136 22710 18148
rect 24412 18136 24440 18167
rect 25498 18164 25504 18176
rect 25556 18164 25562 18216
rect 25700 18213 25728 18312
rect 26234 18300 26240 18352
rect 26292 18340 26298 18352
rect 29178 18340 29184 18352
rect 26292 18312 29184 18340
rect 26292 18300 26298 18312
rect 29178 18300 29184 18312
rect 29236 18300 29242 18352
rect 29546 18340 29552 18352
rect 29507 18312 29552 18340
rect 29546 18300 29552 18312
rect 29604 18300 29610 18352
rect 30374 18300 30380 18352
rect 30432 18340 30438 18352
rect 30432 18312 34008 18340
rect 30432 18300 30438 18312
rect 25884 18244 27292 18272
rect 25884 18216 25912 18244
rect 25685 18207 25743 18213
rect 25685 18173 25697 18207
rect 25731 18173 25743 18207
rect 25866 18204 25872 18216
rect 25827 18176 25872 18204
rect 25685 18167 25743 18173
rect 25866 18164 25872 18176
rect 25924 18164 25930 18216
rect 27154 18204 27160 18216
rect 27115 18176 27160 18204
rect 27154 18164 27160 18176
rect 27212 18164 27218 18216
rect 27264 18204 27292 18244
rect 27338 18232 27344 18284
rect 27396 18272 27402 18284
rect 28166 18272 28172 18284
rect 27396 18244 28172 18272
rect 27396 18232 27402 18244
rect 28166 18232 28172 18244
rect 28224 18232 28230 18284
rect 33980 18281 34008 18312
rect 34146 18300 34152 18352
rect 34204 18340 34210 18352
rect 36170 18340 36176 18352
rect 34204 18312 36176 18340
rect 34204 18300 34210 18312
rect 36170 18300 36176 18312
rect 36228 18300 36234 18352
rect 37550 18300 37556 18352
rect 37608 18340 37614 18352
rect 37829 18343 37887 18349
rect 37829 18340 37841 18343
rect 37608 18312 37841 18340
rect 37608 18300 37614 18312
rect 37829 18309 37841 18312
rect 37875 18309 37887 18343
rect 37829 18303 37887 18309
rect 31481 18275 31539 18281
rect 31481 18272 31493 18275
rect 28276 18244 31493 18272
rect 27433 18207 27491 18213
rect 27433 18204 27445 18207
rect 27264 18176 27445 18204
rect 27433 18173 27445 18176
rect 27479 18173 27491 18207
rect 27433 18167 27491 18173
rect 27522 18164 27528 18216
rect 27580 18204 27586 18216
rect 28077 18207 28135 18213
rect 28077 18204 28089 18207
rect 27580 18176 28089 18204
rect 27580 18164 27586 18176
rect 28077 18173 28089 18176
rect 28123 18173 28135 18207
rect 28077 18167 28135 18173
rect 25038 18136 25044 18148
rect 22704 18108 24440 18136
rect 24999 18108 25044 18136
rect 22704 18096 22710 18108
rect 25038 18096 25044 18108
rect 25096 18096 25102 18148
rect 25406 18096 25412 18148
rect 25464 18136 25470 18148
rect 25884 18136 25912 18164
rect 25464 18108 25912 18136
rect 25464 18096 25470 18108
rect 26050 18096 26056 18148
rect 26108 18136 26114 18148
rect 28276 18136 28304 18244
rect 31481 18241 31493 18244
rect 31527 18241 31539 18275
rect 31481 18235 31539 18241
rect 33965 18275 34023 18281
rect 33965 18241 33977 18275
rect 34011 18241 34023 18275
rect 33965 18235 34023 18241
rect 34514 18232 34520 18284
rect 34572 18272 34578 18284
rect 35713 18275 35771 18281
rect 35713 18272 35725 18275
rect 34572 18244 35725 18272
rect 34572 18232 34578 18244
rect 35713 18241 35725 18244
rect 35759 18241 35771 18275
rect 36722 18272 36728 18284
rect 36683 18244 36728 18272
rect 35713 18235 35771 18241
rect 36722 18232 36728 18244
rect 36780 18232 36786 18284
rect 29457 18207 29515 18213
rect 29457 18173 29469 18207
rect 29503 18173 29515 18207
rect 29822 18204 29828 18216
rect 29783 18176 29828 18204
rect 29457 18167 29515 18173
rect 26108 18108 28304 18136
rect 29472 18136 29500 18167
rect 29822 18164 29828 18176
rect 29880 18164 29886 18216
rect 30190 18204 30196 18216
rect 30151 18176 30196 18204
rect 30190 18164 30196 18176
rect 30248 18164 30254 18216
rect 30837 18207 30895 18213
rect 30837 18173 30849 18207
rect 30883 18173 30895 18207
rect 32030 18204 32036 18216
rect 31991 18176 32036 18204
rect 30837 18167 30895 18173
rect 29730 18136 29736 18148
rect 29472 18108 29736 18136
rect 26108 18096 26114 18108
rect 29730 18096 29736 18108
rect 29788 18096 29794 18148
rect 17405 18071 17463 18077
rect 17405 18068 17417 18071
rect 15028 18040 17417 18068
rect 13633 18031 13691 18037
rect 17405 18037 17417 18040
rect 17451 18068 17463 18071
rect 17862 18068 17868 18080
rect 17451 18040 17868 18068
rect 17451 18037 17463 18040
rect 17405 18031 17463 18037
rect 17862 18028 17868 18040
rect 17920 18028 17926 18080
rect 20441 18071 20499 18077
rect 20441 18037 20453 18071
rect 20487 18068 20499 18071
rect 20530 18068 20536 18080
rect 20487 18040 20536 18068
rect 20487 18037 20499 18040
rect 20441 18031 20499 18037
rect 20530 18028 20536 18040
rect 20588 18028 20594 18080
rect 21082 18068 21088 18080
rect 21043 18040 21088 18068
rect 21082 18028 21088 18040
rect 21140 18028 21146 18080
rect 21177 18071 21235 18077
rect 21177 18037 21189 18071
rect 21223 18068 21235 18071
rect 22094 18068 22100 18080
rect 21223 18040 22100 18068
rect 21223 18037 21235 18040
rect 21177 18031 21235 18037
rect 22094 18028 22100 18040
rect 22152 18028 22158 18080
rect 22186 18028 22192 18080
rect 22244 18068 22250 18080
rect 23014 18068 23020 18080
rect 22244 18040 23020 18068
rect 22244 18028 22250 18040
rect 23014 18028 23020 18040
rect 23072 18028 23078 18080
rect 23842 18068 23848 18080
rect 23803 18040 23848 18068
rect 23842 18028 23848 18040
rect 23900 18028 23906 18080
rect 24486 18068 24492 18080
rect 24447 18040 24492 18068
rect 24486 18028 24492 18040
rect 24544 18028 24550 18080
rect 27154 18028 27160 18080
rect 27212 18068 27218 18080
rect 27798 18068 27804 18080
rect 27212 18040 27804 18068
rect 27212 18028 27218 18040
rect 27798 18028 27804 18040
rect 27856 18068 27862 18080
rect 28261 18071 28319 18077
rect 28261 18068 28273 18071
rect 27856 18040 28273 18068
rect 27856 18028 27862 18040
rect 28261 18037 28273 18040
rect 28307 18037 28319 18071
rect 30852 18068 30880 18167
rect 32030 18164 32036 18176
rect 32088 18164 32094 18216
rect 32214 18204 32220 18216
rect 32175 18176 32220 18204
rect 32214 18164 32220 18176
rect 32272 18164 32278 18216
rect 32306 18164 32312 18216
rect 32364 18204 32370 18216
rect 32493 18207 32551 18213
rect 32364 18176 32409 18204
rect 32364 18164 32370 18176
rect 32493 18173 32505 18207
rect 32539 18173 32551 18207
rect 32766 18204 32772 18216
rect 32727 18176 32772 18204
rect 32493 18167 32551 18173
rect 30929 18139 30987 18145
rect 30929 18105 30941 18139
rect 30975 18136 30987 18139
rect 31754 18136 31760 18148
rect 30975 18108 31760 18136
rect 30975 18105 30987 18108
rect 30929 18099 30987 18105
rect 31754 18096 31760 18108
rect 31812 18136 31818 18148
rect 32508 18136 32536 18167
rect 32766 18164 32772 18176
rect 32824 18164 32830 18216
rect 33134 18164 33140 18216
rect 33192 18204 33198 18216
rect 33413 18207 33471 18213
rect 33413 18204 33425 18207
rect 33192 18176 33425 18204
rect 33192 18164 33198 18176
rect 33413 18173 33425 18176
rect 33459 18173 33471 18207
rect 33413 18167 33471 18173
rect 33873 18207 33931 18213
rect 33873 18173 33885 18207
rect 33919 18173 33931 18207
rect 33873 18167 33931 18173
rect 33888 18136 33916 18167
rect 34698 18164 34704 18216
rect 34756 18204 34762 18216
rect 34885 18207 34943 18213
rect 34885 18204 34897 18207
rect 34756 18176 34897 18204
rect 34756 18164 34762 18176
rect 34885 18173 34897 18176
rect 34931 18173 34943 18207
rect 34885 18167 34943 18173
rect 35621 18207 35679 18213
rect 35621 18173 35633 18207
rect 35667 18204 35679 18207
rect 36262 18204 36268 18216
rect 35667 18176 36268 18204
rect 35667 18173 35679 18176
rect 35621 18167 35679 18173
rect 36262 18164 36268 18176
rect 36320 18164 36326 18216
rect 36449 18207 36507 18213
rect 36449 18173 36461 18207
rect 36495 18204 36507 18207
rect 36538 18204 36544 18216
rect 36495 18176 36544 18204
rect 36495 18173 36507 18176
rect 36449 18167 36507 18173
rect 31812 18108 33916 18136
rect 31812 18096 31818 18108
rect 32582 18068 32588 18080
rect 30852 18040 32588 18068
rect 28261 18031 28319 18037
rect 32582 18028 32588 18040
rect 32640 18028 32646 18080
rect 34974 18068 34980 18080
rect 34935 18040 34980 18068
rect 34974 18028 34980 18040
rect 35032 18028 35038 18080
rect 36262 18028 36268 18080
rect 36320 18068 36326 18080
rect 36464 18068 36492 18167
rect 36538 18164 36544 18176
rect 36596 18164 36602 18216
rect 36320 18040 36492 18068
rect 36320 18028 36326 18040
rect 1104 17978 38824 18000
rect 1104 17926 19606 17978
rect 19658 17926 19670 17978
rect 19722 17926 19734 17978
rect 19786 17926 19798 17978
rect 19850 17926 38824 17978
rect 1104 17904 38824 17926
rect 3418 17864 3424 17876
rect 3379 17836 3424 17864
rect 3418 17824 3424 17836
rect 3476 17824 3482 17876
rect 8386 17824 8392 17876
rect 8444 17864 8450 17876
rect 8757 17867 8815 17873
rect 8757 17864 8769 17867
rect 8444 17836 8769 17864
rect 8444 17824 8450 17836
rect 8757 17833 8769 17836
rect 8803 17833 8815 17867
rect 8757 17827 8815 17833
rect 11701 17867 11759 17873
rect 11701 17833 11713 17867
rect 11747 17864 11759 17867
rect 12618 17864 12624 17876
rect 11747 17836 12624 17864
rect 11747 17833 11759 17836
rect 11701 17827 11759 17833
rect 12618 17824 12624 17836
rect 12676 17824 12682 17876
rect 19613 17867 19671 17873
rect 19613 17833 19625 17867
rect 19659 17864 19671 17867
rect 19978 17864 19984 17876
rect 19659 17836 19984 17864
rect 19659 17833 19671 17836
rect 19613 17827 19671 17833
rect 19978 17824 19984 17836
rect 20036 17824 20042 17876
rect 20714 17824 20720 17876
rect 20772 17864 20778 17876
rect 21177 17867 21235 17873
rect 21177 17864 21189 17867
rect 20772 17836 21189 17864
rect 20772 17824 20778 17836
rect 21177 17833 21189 17836
rect 21223 17833 21235 17867
rect 21177 17827 21235 17833
rect 24394 17824 24400 17876
rect 24452 17824 24458 17876
rect 25958 17824 25964 17876
rect 26016 17864 26022 17876
rect 28810 17864 28816 17876
rect 26016 17836 28816 17864
rect 26016 17824 26022 17836
rect 28810 17824 28816 17836
rect 28868 17824 28874 17876
rect 29270 17824 29276 17876
rect 29328 17864 29334 17876
rect 29825 17867 29883 17873
rect 29825 17864 29837 17867
rect 29328 17836 29837 17864
rect 29328 17824 29334 17836
rect 29825 17833 29837 17836
rect 29871 17864 29883 17867
rect 30098 17864 30104 17876
rect 29871 17836 30104 17864
rect 29871 17833 29883 17836
rect 29825 17827 29883 17833
rect 30098 17824 30104 17836
rect 30156 17824 30162 17876
rect 32030 17824 32036 17876
rect 32088 17864 32094 17876
rect 33962 17864 33968 17876
rect 32088 17836 33968 17864
rect 32088 17824 32094 17836
rect 33962 17824 33968 17836
rect 34020 17824 34026 17876
rect 7006 17796 7012 17808
rect 6967 17768 7012 17796
rect 7006 17756 7012 17768
rect 7064 17756 7070 17808
rect 14645 17799 14703 17805
rect 14645 17765 14657 17799
rect 14691 17796 14703 17799
rect 14691 17768 16896 17796
rect 14691 17765 14703 17768
rect 14645 17759 14703 17765
rect 4341 17731 4399 17737
rect 4341 17697 4353 17731
rect 4387 17728 4399 17731
rect 4614 17728 4620 17740
rect 4387 17700 4620 17728
rect 4387 17697 4399 17700
rect 4341 17691 4399 17697
rect 4614 17688 4620 17700
rect 4672 17688 4678 17740
rect 4801 17731 4859 17737
rect 4801 17697 4813 17731
rect 4847 17728 4859 17731
rect 5442 17728 5448 17740
rect 4847 17700 5448 17728
rect 4847 17697 4859 17700
rect 4801 17691 4859 17697
rect 5442 17688 5448 17700
rect 5500 17688 5506 17740
rect 5902 17688 5908 17740
rect 5960 17728 5966 17740
rect 7653 17731 7711 17737
rect 5960 17700 7604 17728
rect 5960 17688 5966 17700
rect 1394 17620 1400 17672
rect 1452 17660 1458 17672
rect 1857 17663 1915 17669
rect 1857 17660 1869 17663
rect 1452 17632 1869 17660
rect 1452 17620 1458 17632
rect 1857 17629 1869 17632
rect 1903 17629 1915 17663
rect 2130 17660 2136 17672
rect 2091 17632 2136 17660
rect 1857 17623 1915 17629
rect 2130 17620 2136 17632
rect 2188 17620 2194 17672
rect 5350 17660 5356 17672
rect 5311 17632 5356 17660
rect 5350 17620 5356 17632
rect 5408 17620 5414 17672
rect 7576 17669 7604 17700
rect 7653 17697 7665 17731
rect 7699 17728 7711 17731
rect 8386 17728 8392 17740
rect 7699 17700 8392 17728
rect 7699 17697 7711 17700
rect 7653 17691 7711 17697
rect 8386 17688 8392 17700
rect 8444 17688 8450 17740
rect 8665 17731 8723 17737
rect 8665 17697 8677 17731
rect 8711 17728 8723 17731
rect 9766 17728 9772 17740
rect 8711 17700 9772 17728
rect 8711 17697 8723 17700
rect 8665 17691 8723 17697
rect 9766 17688 9772 17700
rect 9824 17688 9830 17740
rect 10413 17731 10471 17737
rect 10413 17697 10425 17731
rect 10459 17728 10471 17731
rect 12526 17728 12532 17740
rect 10459 17700 12388 17728
rect 12487 17700 12532 17728
rect 10459 17697 10471 17700
rect 10413 17691 10471 17697
rect 5629 17663 5687 17669
rect 5629 17629 5641 17663
rect 5675 17660 5687 17663
rect 7561 17663 7619 17669
rect 5675 17632 7512 17660
rect 5675 17629 5687 17632
rect 5629 17623 5687 17629
rect 7484 17592 7512 17632
rect 7561 17629 7573 17663
rect 7607 17660 7619 17663
rect 9674 17660 9680 17672
rect 7607 17632 9680 17660
rect 7607 17629 7619 17632
rect 7561 17623 7619 17629
rect 9674 17620 9680 17632
rect 9732 17620 9738 17672
rect 10134 17660 10140 17672
rect 10047 17632 10140 17660
rect 10134 17620 10140 17632
rect 10192 17620 10198 17672
rect 11882 17620 11888 17672
rect 11940 17660 11946 17672
rect 12253 17663 12311 17669
rect 12253 17660 12265 17663
rect 11940 17632 12265 17660
rect 11940 17620 11946 17632
rect 12253 17629 12265 17632
rect 12299 17629 12311 17663
rect 12360 17660 12388 17700
rect 12526 17688 12532 17700
rect 12584 17688 12590 17740
rect 14553 17731 14611 17737
rect 14553 17697 14565 17731
rect 14599 17728 14611 17731
rect 15286 17728 15292 17740
rect 14599 17700 15292 17728
rect 14599 17697 14611 17700
rect 14553 17691 14611 17697
rect 15286 17688 15292 17700
rect 15344 17688 15350 17740
rect 15654 17728 15660 17740
rect 15615 17700 15660 17728
rect 15654 17688 15660 17700
rect 15712 17688 15718 17740
rect 16114 17728 16120 17740
rect 16075 17700 16120 17728
rect 16114 17688 16120 17700
rect 16172 17688 16178 17740
rect 16868 17737 16896 17768
rect 18598 17756 18604 17808
rect 18656 17796 18662 17808
rect 18656 17768 19472 17796
rect 18656 17756 18662 17768
rect 16853 17731 16911 17737
rect 16853 17697 16865 17731
rect 16899 17697 16911 17731
rect 17218 17728 17224 17740
rect 17179 17700 17224 17728
rect 16853 17691 16911 17697
rect 17218 17688 17224 17700
rect 17276 17688 17282 17740
rect 17310 17688 17316 17740
rect 17368 17728 17374 17740
rect 17681 17731 17739 17737
rect 17681 17728 17693 17731
rect 17368 17700 17693 17728
rect 17368 17688 17374 17700
rect 17681 17697 17693 17700
rect 17727 17697 17739 17731
rect 17681 17691 17739 17697
rect 18509 17731 18567 17737
rect 18509 17697 18521 17731
rect 18555 17728 18567 17731
rect 18690 17728 18696 17740
rect 18555 17700 18696 17728
rect 18555 17697 18567 17700
rect 18509 17691 18567 17697
rect 18690 17688 18696 17700
rect 18748 17688 18754 17740
rect 19444 17737 19472 17768
rect 23474 17756 23480 17808
rect 23532 17796 23538 17808
rect 23569 17799 23627 17805
rect 23569 17796 23581 17799
rect 23532 17768 23581 17796
rect 23532 17756 23538 17768
rect 23569 17765 23581 17768
rect 23615 17765 23627 17799
rect 24412 17796 24440 17824
rect 27062 17796 27068 17808
rect 23569 17759 23627 17765
rect 23952 17768 24440 17796
rect 25700 17768 26740 17796
rect 27023 17768 27068 17796
rect 19429 17731 19487 17737
rect 19429 17697 19441 17731
rect 19475 17697 19487 17731
rect 19429 17691 19487 17697
rect 20165 17731 20223 17737
rect 20165 17697 20177 17731
rect 20211 17728 20223 17731
rect 20438 17728 20444 17740
rect 20211 17700 20444 17728
rect 20211 17697 20223 17700
rect 20165 17691 20223 17697
rect 20438 17688 20444 17700
rect 20496 17728 20502 17740
rect 20993 17731 21051 17737
rect 20993 17728 21005 17731
rect 20496 17700 21005 17728
rect 20496 17688 20502 17700
rect 20993 17697 21005 17700
rect 21039 17697 21051 17731
rect 20993 17691 21051 17697
rect 22189 17731 22247 17737
rect 22189 17697 22201 17731
rect 22235 17728 22247 17731
rect 22278 17728 22284 17740
rect 22235 17700 22284 17728
rect 22235 17697 22247 17700
rect 22189 17691 22247 17697
rect 22278 17688 22284 17700
rect 22336 17688 22342 17740
rect 22557 17731 22615 17737
rect 22557 17697 22569 17731
rect 22603 17728 22615 17731
rect 22922 17728 22928 17740
rect 22603 17700 22928 17728
rect 22603 17697 22615 17700
rect 22557 17691 22615 17697
rect 22922 17688 22928 17700
rect 22980 17688 22986 17740
rect 23198 17728 23204 17740
rect 23159 17700 23204 17728
rect 23198 17688 23204 17700
rect 23256 17688 23262 17740
rect 23658 17688 23664 17740
rect 23716 17728 23722 17740
rect 23952 17737 23980 17768
rect 25700 17740 25728 17768
rect 23937 17731 23995 17737
rect 23937 17728 23949 17731
rect 23716 17700 23949 17728
rect 23716 17688 23722 17700
rect 23937 17697 23949 17700
rect 23983 17697 23995 17731
rect 23937 17691 23995 17697
rect 24118 17688 24124 17740
rect 24176 17728 24182 17740
rect 24397 17731 24455 17737
rect 24397 17728 24409 17731
rect 24176 17700 24409 17728
rect 24176 17688 24182 17700
rect 24397 17697 24409 17700
rect 24443 17728 24455 17731
rect 24578 17728 24584 17740
rect 24443 17700 24584 17728
rect 24443 17697 24455 17700
rect 24397 17691 24455 17697
rect 24578 17688 24584 17700
rect 24636 17688 24642 17740
rect 24673 17731 24731 17737
rect 24673 17697 24685 17731
rect 24719 17697 24731 17731
rect 24854 17728 24860 17740
rect 24815 17700 24860 17728
rect 24673 17691 24731 17697
rect 12360 17632 14596 17660
rect 12253 17623 12311 17629
rect 8938 17592 8944 17604
rect 7484 17564 8944 17592
rect 8938 17552 8944 17564
rect 8996 17552 9002 17604
rect 3694 17484 3700 17536
rect 3752 17524 3758 17536
rect 4157 17527 4215 17533
rect 4157 17524 4169 17527
rect 3752 17496 4169 17524
rect 3752 17484 3758 17496
rect 4157 17493 4169 17496
rect 4203 17493 4215 17527
rect 7834 17524 7840 17536
rect 7795 17496 7840 17524
rect 4157 17487 4215 17493
rect 7834 17484 7840 17496
rect 7892 17484 7898 17536
rect 10152 17524 10180 17620
rect 12710 17524 12716 17536
rect 10152 17496 12716 17524
rect 12710 17484 12716 17496
rect 12768 17484 12774 17536
rect 13814 17524 13820 17536
rect 13775 17496 13820 17524
rect 13814 17484 13820 17496
rect 13872 17484 13878 17536
rect 14568 17524 14596 17632
rect 14642 17620 14648 17672
rect 14700 17660 14706 17672
rect 15381 17663 15439 17669
rect 15381 17660 15393 17663
rect 14700 17632 15393 17660
rect 14700 17620 14706 17632
rect 15381 17629 15393 17632
rect 15427 17629 15439 17663
rect 15381 17623 15439 17629
rect 18417 17663 18475 17669
rect 18417 17629 18429 17663
rect 18463 17660 18475 17663
rect 19058 17660 19064 17672
rect 18463 17632 19064 17660
rect 18463 17629 18475 17632
rect 18417 17623 18475 17629
rect 19058 17620 19064 17632
rect 19116 17620 19122 17672
rect 22649 17663 22707 17669
rect 22649 17629 22661 17663
rect 22695 17660 22707 17663
rect 23382 17660 23388 17672
rect 22695 17632 23388 17660
rect 22695 17629 22707 17632
rect 22649 17623 22707 17629
rect 23382 17620 23388 17632
rect 23440 17660 23446 17672
rect 23842 17660 23848 17672
rect 23440 17632 23848 17660
rect 23440 17620 23446 17632
rect 23842 17620 23848 17632
rect 23900 17620 23906 17672
rect 24688 17604 24716 17691
rect 24854 17688 24860 17700
rect 24912 17688 24918 17740
rect 25682 17728 25688 17740
rect 25643 17700 25688 17728
rect 25682 17688 25688 17700
rect 25740 17688 25746 17740
rect 26510 17728 26516 17740
rect 26471 17700 26516 17728
rect 26510 17688 26516 17700
rect 26568 17688 26574 17740
rect 26712 17737 26740 17768
rect 27062 17756 27068 17768
rect 27120 17756 27126 17808
rect 33042 17796 33048 17808
rect 27540 17768 30604 17796
rect 26697 17731 26755 17737
rect 26697 17697 26709 17731
rect 26743 17728 26755 17731
rect 27540 17728 27568 17768
rect 26743 17700 27568 17728
rect 26743 17697 26755 17700
rect 26697 17691 26755 17697
rect 27614 17688 27620 17740
rect 27672 17728 27678 17740
rect 28368 17737 28396 17768
rect 28261 17731 28319 17737
rect 28261 17728 28273 17731
rect 27672 17700 28273 17728
rect 27672 17688 27678 17700
rect 28261 17697 28273 17700
rect 28307 17697 28319 17731
rect 28261 17691 28319 17697
rect 28353 17731 28411 17737
rect 28353 17697 28365 17731
rect 28399 17697 28411 17731
rect 28626 17728 28632 17740
rect 28587 17700 28632 17728
rect 28353 17691 28411 17697
rect 28626 17688 28632 17700
rect 28684 17688 28690 17740
rect 28810 17688 28816 17740
rect 28868 17728 28874 17740
rect 29362 17728 29368 17740
rect 28868 17700 29368 17728
rect 28868 17688 28874 17700
rect 29362 17688 29368 17700
rect 29420 17728 29426 17740
rect 29641 17731 29699 17737
rect 29641 17728 29653 17731
rect 29420 17700 29653 17728
rect 29420 17688 29426 17700
rect 29641 17697 29653 17700
rect 29687 17697 29699 17731
rect 30466 17728 30472 17740
rect 30427 17700 30472 17728
rect 29641 17691 29699 17697
rect 30466 17688 30472 17700
rect 30524 17688 30530 17740
rect 25774 17620 25780 17672
rect 25832 17660 25838 17672
rect 26234 17660 26240 17672
rect 25832 17632 26240 17660
rect 25832 17620 25838 17632
rect 26234 17620 26240 17632
rect 26292 17660 26298 17672
rect 28721 17663 28779 17669
rect 28721 17660 28733 17663
rect 26292 17632 28733 17660
rect 26292 17620 26298 17632
rect 28721 17629 28733 17632
rect 28767 17660 28779 17663
rect 28994 17660 29000 17672
rect 28767 17632 29000 17660
rect 28767 17629 28779 17632
rect 28721 17623 28779 17629
rect 28994 17620 29000 17632
rect 29052 17620 29058 17672
rect 30576 17669 30604 17768
rect 32600 17768 33048 17796
rect 31018 17728 31024 17740
rect 30979 17700 31024 17728
rect 31018 17688 31024 17700
rect 31076 17688 31082 17740
rect 31202 17728 31208 17740
rect 31163 17700 31208 17728
rect 31202 17688 31208 17700
rect 31260 17728 31266 17740
rect 32600 17737 32628 17768
rect 33042 17756 33048 17768
rect 33100 17756 33106 17808
rect 33778 17796 33784 17808
rect 33739 17768 33784 17796
rect 33778 17756 33784 17768
rect 33836 17756 33842 17808
rect 37185 17799 37243 17805
rect 37185 17765 37197 17799
rect 37231 17796 37243 17799
rect 37274 17796 37280 17808
rect 37231 17768 37280 17796
rect 37231 17765 37243 17768
rect 37185 17759 37243 17765
rect 37274 17756 37280 17768
rect 37332 17756 37338 17808
rect 32125 17731 32183 17737
rect 32125 17728 32137 17731
rect 31260 17700 32137 17728
rect 31260 17688 31266 17700
rect 32125 17697 32137 17700
rect 32171 17697 32183 17731
rect 32125 17691 32183 17697
rect 32585 17731 32643 17737
rect 32585 17697 32597 17731
rect 32631 17697 32643 17731
rect 32766 17728 32772 17740
rect 32727 17700 32772 17728
rect 32585 17691 32643 17697
rect 32766 17688 32772 17700
rect 32824 17688 32830 17740
rect 32953 17731 33011 17737
rect 32953 17697 32965 17731
rect 32999 17697 33011 17731
rect 32953 17691 33011 17697
rect 30561 17663 30619 17669
rect 30561 17629 30573 17663
rect 30607 17629 30619 17663
rect 30561 17623 30619 17629
rect 30742 17620 30748 17672
rect 30800 17660 30806 17672
rect 31294 17660 31300 17672
rect 30800 17632 31300 17660
rect 30800 17620 30806 17632
rect 31294 17620 31300 17632
rect 31352 17660 31358 17672
rect 32968 17660 32996 17691
rect 34422 17688 34428 17740
rect 34480 17728 34486 17740
rect 34609 17731 34667 17737
rect 34609 17728 34621 17731
rect 34480 17700 34621 17728
rect 34480 17688 34486 17700
rect 34609 17697 34621 17700
rect 34655 17697 34667 17731
rect 34790 17728 34796 17740
rect 34751 17700 34796 17728
rect 34609 17691 34667 17697
rect 34790 17688 34796 17700
rect 34848 17688 34854 17740
rect 34974 17688 34980 17740
rect 35032 17728 35038 17740
rect 35805 17731 35863 17737
rect 35805 17728 35817 17731
rect 35032 17700 35817 17728
rect 35032 17688 35038 17700
rect 35805 17697 35817 17700
rect 35851 17697 35863 17731
rect 35805 17691 35863 17697
rect 37737 17731 37795 17737
rect 37737 17697 37749 17731
rect 37783 17697 37795 17731
rect 37737 17691 37795 17697
rect 34330 17660 34336 17672
rect 31352 17632 32996 17660
rect 34291 17632 34336 17660
rect 31352 17620 31358 17632
rect 34330 17620 34336 17632
rect 34388 17620 34394 17672
rect 35529 17663 35587 17669
rect 35529 17629 35541 17663
rect 35575 17629 35587 17663
rect 35529 17623 35587 17629
rect 15470 17552 15476 17604
rect 15528 17592 15534 17604
rect 16117 17595 16175 17601
rect 16117 17592 16129 17595
rect 15528 17564 16129 17592
rect 15528 17552 15534 17564
rect 16117 17561 16129 17564
rect 16163 17561 16175 17595
rect 17678 17592 17684 17604
rect 17639 17564 17684 17592
rect 16117 17555 16175 17561
rect 17678 17552 17684 17564
rect 17736 17552 17742 17604
rect 17770 17552 17776 17604
rect 17828 17592 17834 17604
rect 18138 17592 18144 17604
rect 17828 17564 18144 17592
rect 17828 17552 17834 17564
rect 18138 17552 18144 17564
rect 18196 17552 18202 17604
rect 21174 17552 21180 17604
rect 21232 17592 21238 17604
rect 21726 17592 21732 17604
rect 21232 17564 21732 17592
rect 21232 17552 21238 17564
rect 21726 17552 21732 17564
rect 21784 17552 21790 17604
rect 22005 17595 22063 17601
rect 22005 17561 22017 17595
rect 22051 17592 22063 17595
rect 23290 17592 23296 17604
rect 22051 17564 23296 17592
rect 22051 17561 22063 17564
rect 22005 17555 22063 17561
rect 23290 17552 23296 17564
rect 23348 17552 23354 17604
rect 24670 17592 24676 17604
rect 24583 17564 24676 17592
rect 24670 17552 24676 17564
rect 24728 17592 24734 17604
rect 34606 17592 34612 17604
rect 24728 17564 34612 17592
rect 24728 17552 24734 17564
rect 34606 17552 34612 17564
rect 34664 17552 34670 17604
rect 18693 17527 18751 17533
rect 18693 17524 18705 17527
rect 14568 17496 18705 17524
rect 18693 17493 18705 17496
rect 18739 17493 18751 17527
rect 18693 17487 18751 17493
rect 19886 17484 19892 17536
rect 19944 17524 19950 17536
rect 20162 17524 20168 17536
rect 19944 17496 20168 17524
rect 19944 17484 19950 17496
rect 20162 17484 20168 17496
rect 20220 17484 20226 17536
rect 20257 17527 20315 17533
rect 20257 17493 20269 17527
rect 20303 17524 20315 17527
rect 20346 17524 20352 17536
rect 20303 17496 20352 17524
rect 20303 17493 20315 17496
rect 20257 17487 20315 17493
rect 20346 17484 20352 17496
rect 20404 17524 20410 17536
rect 20898 17524 20904 17536
rect 20404 17496 20904 17524
rect 20404 17484 20410 17496
rect 20898 17484 20904 17496
rect 20956 17484 20962 17536
rect 21266 17484 21272 17536
rect 21324 17524 21330 17536
rect 23566 17524 23572 17536
rect 21324 17496 23572 17524
rect 21324 17484 21330 17496
rect 23566 17484 23572 17496
rect 23624 17484 23630 17536
rect 25866 17524 25872 17536
rect 25827 17496 25872 17524
rect 25866 17484 25872 17496
rect 25924 17484 25930 17536
rect 27709 17527 27767 17533
rect 27709 17493 27721 17527
rect 27755 17524 27767 17527
rect 27890 17524 27896 17536
rect 27755 17496 27896 17524
rect 27755 17493 27767 17496
rect 27709 17487 27767 17493
rect 27890 17484 27896 17496
rect 27948 17484 27954 17536
rect 30374 17484 30380 17536
rect 30432 17524 30438 17536
rect 30558 17524 30564 17536
rect 30432 17496 30564 17524
rect 30432 17484 30438 17496
rect 30558 17484 30564 17496
rect 30616 17484 30622 17536
rect 34514 17484 34520 17536
rect 34572 17524 34578 17536
rect 35544 17524 35572 17623
rect 35710 17620 35716 17672
rect 35768 17660 35774 17672
rect 37752 17660 37780 17691
rect 35768 17632 37780 17660
rect 35768 17620 35774 17632
rect 36262 17524 36268 17536
rect 34572 17496 36268 17524
rect 34572 17484 34578 17496
rect 36262 17484 36268 17496
rect 36320 17484 36326 17536
rect 37826 17524 37832 17536
rect 37787 17496 37832 17524
rect 37826 17484 37832 17496
rect 37884 17484 37890 17536
rect 1104 17434 38824 17456
rect 1104 17382 4246 17434
rect 4298 17382 4310 17434
rect 4362 17382 4374 17434
rect 4426 17382 4438 17434
rect 4490 17382 34966 17434
rect 35018 17382 35030 17434
rect 35082 17382 35094 17434
rect 35146 17382 35158 17434
rect 35210 17382 38824 17434
rect 1104 17360 38824 17382
rect 2130 17320 2136 17332
rect 2091 17292 2136 17320
rect 2130 17280 2136 17292
rect 2188 17280 2194 17332
rect 5994 17280 6000 17332
rect 6052 17320 6058 17332
rect 23566 17320 23572 17332
rect 6052 17292 23572 17320
rect 6052 17280 6058 17292
rect 23566 17280 23572 17292
rect 23624 17280 23630 17332
rect 24394 17280 24400 17332
rect 24452 17320 24458 17332
rect 27890 17320 27896 17332
rect 24452 17292 26648 17320
rect 27851 17292 27896 17320
rect 24452 17280 24458 17292
rect 12342 17252 12348 17264
rect 10428 17224 12348 17252
rect 2777 17187 2835 17193
rect 2777 17184 2789 17187
rect 2056 17156 2789 17184
rect 2056 17125 2084 17156
rect 2777 17153 2789 17156
rect 2823 17153 2835 17187
rect 5626 17184 5632 17196
rect 2777 17147 2835 17153
rect 3344 17156 5632 17184
rect 2041 17119 2099 17125
rect 2041 17085 2053 17119
rect 2087 17085 2099 17119
rect 2866 17116 2872 17128
rect 2827 17088 2872 17116
rect 2041 17079 2099 17085
rect 2866 17076 2872 17088
rect 2924 17076 2930 17128
rect 3344 17125 3372 17156
rect 3329 17119 3387 17125
rect 3329 17085 3341 17119
rect 3375 17085 3387 17119
rect 3694 17116 3700 17128
rect 3655 17088 3700 17116
rect 3329 17079 3387 17085
rect 3694 17076 3700 17088
rect 3752 17076 3758 17128
rect 4982 17116 4988 17128
rect 4943 17088 4988 17116
rect 4982 17076 4988 17088
rect 5040 17076 5046 17128
rect 5368 17125 5396 17156
rect 5626 17144 5632 17156
rect 5684 17184 5690 17196
rect 5902 17184 5908 17196
rect 5684 17156 5908 17184
rect 5684 17144 5690 17156
rect 5902 17144 5908 17156
rect 5960 17144 5966 17196
rect 8662 17184 8668 17196
rect 7024 17156 8668 17184
rect 5353 17119 5411 17125
rect 5353 17085 5365 17119
rect 5399 17085 5411 17119
rect 5353 17079 5411 17085
rect 5721 17119 5779 17125
rect 5721 17085 5733 17119
rect 5767 17116 5779 17119
rect 6914 17116 6920 17128
rect 5767 17088 6920 17116
rect 5767 17085 5779 17088
rect 5721 17079 5779 17085
rect 6914 17076 6920 17088
rect 6972 17076 6978 17128
rect 7024 17125 7052 17156
rect 8662 17144 8668 17156
rect 8720 17144 8726 17196
rect 7009 17119 7067 17125
rect 7009 17085 7021 17119
rect 7055 17085 7067 17119
rect 7742 17116 7748 17128
rect 7703 17088 7748 17116
rect 7009 17079 7067 17085
rect 7742 17076 7748 17088
rect 7800 17076 7806 17128
rect 8018 17116 8024 17128
rect 7979 17088 8024 17116
rect 8018 17076 8024 17088
rect 8076 17076 8082 17128
rect 9858 17116 9864 17128
rect 9819 17088 9864 17116
rect 9858 17076 9864 17088
rect 9916 17076 9922 17128
rect 10428 17125 10456 17224
rect 12342 17212 12348 17224
rect 12400 17212 12406 17264
rect 12710 17212 12716 17264
rect 12768 17252 12774 17264
rect 12768 17224 15148 17252
rect 12768 17212 12774 17224
rect 15120 17196 15148 17224
rect 16114 17212 16120 17264
rect 16172 17252 16178 17264
rect 20438 17252 20444 17264
rect 16172 17224 18736 17252
rect 20399 17224 20444 17252
rect 16172 17212 16178 17224
rect 10686 17184 10692 17196
rect 10647 17156 10692 17184
rect 10686 17144 10692 17156
rect 10744 17144 10750 17196
rect 14553 17187 14611 17193
rect 14553 17153 14565 17187
rect 14599 17184 14611 17187
rect 14642 17184 14648 17196
rect 14599 17156 14648 17184
rect 14599 17153 14611 17156
rect 14553 17147 14611 17153
rect 14642 17144 14648 17156
rect 14700 17144 14706 17196
rect 15102 17184 15108 17196
rect 15015 17156 15108 17184
rect 15102 17144 15108 17156
rect 15160 17144 15166 17196
rect 15381 17187 15439 17193
rect 15381 17153 15393 17187
rect 15427 17184 15439 17187
rect 18601 17187 18659 17193
rect 18601 17184 18613 17187
rect 15427 17156 18613 17184
rect 15427 17153 15439 17156
rect 15381 17147 15439 17153
rect 18601 17153 18613 17156
rect 18647 17153 18659 17187
rect 18708 17184 18736 17224
rect 20438 17212 20444 17224
rect 20496 17212 20502 17264
rect 21082 17212 21088 17264
rect 21140 17252 21146 17264
rect 21140 17224 21404 17252
rect 21140 17212 21146 17224
rect 18708 17156 21312 17184
rect 18601 17147 18659 17153
rect 10413 17119 10471 17125
rect 10413 17085 10425 17119
rect 10459 17085 10471 17119
rect 10413 17079 10471 17085
rect 10781 17119 10839 17125
rect 10781 17085 10793 17119
rect 10827 17116 10839 17119
rect 11054 17116 11060 17128
rect 10827 17088 11060 17116
rect 10827 17085 10839 17088
rect 10781 17079 10839 17085
rect 11054 17076 11060 17088
rect 11112 17076 11118 17128
rect 12805 17119 12863 17125
rect 12805 17085 12817 17119
rect 12851 17085 12863 17119
rect 13630 17116 13636 17128
rect 13591 17088 13636 17116
rect 12805 17079 12863 17085
rect 5902 17048 5908 17060
rect 5863 17020 5908 17048
rect 5902 17008 5908 17020
rect 5960 17008 5966 17060
rect 12618 17048 12624 17060
rect 9232 17020 12624 17048
rect 7190 16980 7196 16992
rect 7151 16952 7196 16980
rect 7190 16940 7196 16952
rect 7248 16940 7254 16992
rect 7558 16940 7564 16992
rect 7616 16980 7622 16992
rect 9232 16980 9260 17020
rect 12618 17008 12624 17020
rect 12676 17008 12682 17060
rect 12820 17048 12848 17079
rect 13630 17076 13636 17088
rect 13688 17076 13694 17128
rect 13814 17116 13820 17128
rect 13775 17088 13820 17116
rect 13814 17076 13820 17088
rect 13872 17076 13878 17128
rect 14182 17076 14188 17128
rect 14240 17116 14246 17128
rect 14277 17119 14335 17125
rect 14277 17116 14289 17119
rect 14240 17088 14289 17116
rect 14240 17076 14246 17088
rect 14277 17085 14289 17088
rect 14323 17085 14335 17119
rect 16114 17116 16120 17128
rect 14277 17079 14335 17085
rect 15212 17088 16120 17116
rect 15212 17048 15240 17088
rect 16114 17076 16120 17088
rect 16172 17076 16178 17128
rect 17126 17076 17132 17128
rect 17184 17116 17190 17128
rect 17221 17119 17279 17125
rect 17221 17116 17233 17119
rect 17184 17088 17233 17116
rect 17184 17076 17190 17088
rect 17221 17085 17233 17088
rect 17267 17116 17279 17119
rect 17310 17116 17316 17128
rect 17267 17088 17316 17116
rect 17267 17085 17279 17088
rect 17221 17079 17279 17085
rect 17310 17076 17316 17088
rect 17368 17076 17374 17128
rect 18046 17116 18052 17128
rect 18007 17088 18052 17116
rect 18046 17076 18052 17088
rect 18104 17076 18110 17128
rect 18138 17076 18144 17128
rect 18196 17116 18202 17128
rect 19061 17119 19119 17125
rect 18196 17088 18241 17116
rect 18196 17076 18202 17088
rect 19061 17085 19073 17119
rect 19107 17085 19119 17119
rect 19334 17116 19340 17128
rect 19295 17088 19340 17116
rect 19061 17079 19119 17085
rect 12820 17020 15240 17048
rect 7616 16952 9260 16980
rect 9309 16983 9367 16989
rect 7616 16940 7622 16952
rect 9309 16949 9321 16983
rect 9355 16980 9367 16983
rect 9766 16980 9772 16992
rect 9355 16952 9772 16980
rect 9355 16949 9367 16952
rect 9309 16943 9367 16949
rect 9766 16940 9772 16952
rect 9824 16940 9830 16992
rect 12434 16940 12440 16992
rect 12492 16980 12498 16992
rect 12897 16983 12955 16989
rect 12897 16980 12909 16983
rect 12492 16952 12909 16980
rect 12492 16940 12498 16952
rect 12897 16949 12909 16952
rect 12943 16949 12955 16983
rect 12897 16943 12955 16949
rect 16114 16940 16120 16992
rect 16172 16980 16178 16992
rect 16485 16983 16543 16989
rect 16485 16980 16497 16983
rect 16172 16952 16497 16980
rect 16172 16940 16178 16952
rect 16485 16949 16497 16952
rect 16531 16949 16543 16983
rect 16485 16943 16543 16949
rect 17405 16983 17463 16989
rect 17405 16949 17417 16983
rect 17451 16980 17463 16983
rect 18064 16980 18092 17076
rect 18506 17008 18512 17060
rect 18564 17048 18570 17060
rect 18966 17048 18972 17060
rect 18564 17020 18972 17048
rect 18564 17008 18570 17020
rect 18966 17008 18972 17020
rect 19024 17008 19030 17060
rect 17451 16952 18092 16980
rect 17451 16949 17463 16952
rect 17405 16943 17463 16949
rect 18138 16940 18144 16992
rect 18196 16980 18202 16992
rect 19076 16980 19104 17079
rect 19334 17076 19340 17088
rect 19392 17076 19398 17128
rect 21174 17116 21180 17128
rect 21135 17088 21180 17116
rect 21174 17076 21180 17088
rect 21232 17076 21238 17128
rect 20162 16980 20168 16992
rect 18196 16952 20168 16980
rect 18196 16940 18202 16952
rect 20162 16940 20168 16952
rect 20220 16980 20226 16992
rect 20530 16980 20536 16992
rect 20220 16952 20536 16980
rect 20220 16940 20226 16952
rect 20530 16940 20536 16952
rect 20588 16940 20594 16992
rect 21284 16989 21312 17156
rect 21376 17116 21404 17224
rect 21818 17212 21824 17264
rect 21876 17252 21882 17264
rect 22186 17252 22192 17264
rect 21876 17224 22192 17252
rect 21876 17212 21882 17224
rect 22186 17212 22192 17224
rect 22244 17212 22250 17264
rect 24854 17252 24860 17264
rect 24815 17224 24860 17252
rect 24854 17212 24860 17224
rect 24912 17212 24918 17264
rect 25869 17255 25927 17261
rect 25869 17221 25881 17255
rect 25915 17252 25927 17255
rect 26510 17252 26516 17264
rect 25915 17224 26516 17252
rect 25915 17221 25927 17224
rect 25869 17215 25927 17221
rect 26510 17212 26516 17224
rect 26568 17212 26574 17264
rect 26620 17252 26648 17292
rect 27890 17280 27896 17292
rect 27948 17280 27954 17332
rect 28350 17320 28356 17332
rect 28311 17292 28356 17320
rect 28350 17280 28356 17292
rect 28408 17280 28414 17332
rect 28994 17280 29000 17332
rect 29052 17320 29058 17332
rect 37826 17320 37832 17332
rect 29052 17292 37832 17320
rect 29052 17280 29058 17292
rect 37826 17280 37832 17292
rect 37884 17280 37890 17332
rect 30650 17252 30656 17264
rect 26620 17224 30656 17252
rect 30650 17212 30656 17224
rect 30708 17212 30714 17264
rect 31110 17212 31116 17264
rect 31168 17252 31174 17264
rect 33318 17252 33324 17264
rect 31168 17224 33324 17252
rect 31168 17212 31174 17224
rect 33318 17212 33324 17224
rect 33376 17212 33382 17264
rect 35161 17255 35219 17261
rect 33428 17224 35112 17252
rect 26418 17184 26424 17196
rect 26160 17156 26424 17184
rect 21913 17119 21971 17125
rect 21913 17116 21925 17119
rect 21376 17088 21925 17116
rect 21913 17085 21925 17088
rect 21959 17085 21971 17119
rect 21913 17079 21971 17085
rect 21928 17048 21956 17079
rect 22002 17076 22008 17128
rect 22060 17116 22066 17128
rect 22557 17119 22615 17125
rect 22060 17088 22105 17116
rect 22060 17076 22066 17088
rect 22557 17085 22569 17119
rect 22603 17116 22615 17119
rect 22646 17116 22652 17128
rect 22603 17088 22652 17116
rect 22603 17085 22615 17088
rect 22557 17079 22615 17085
rect 22646 17076 22652 17088
rect 22704 17076 22710 17128
rect 23477 17119 23535 17125
rect 23477 17085 23489 17119
rect 23523 17116 23535 17119
rect 23750 17116 23756 17128
rect 23523 17088 23756 17116
rect 23523 17085 23535 17088
rect 23477 17079 23535 17085
rect 23750 17076 23756 17088
rect 23808 17076 23814 17128
rect 23842 17076 23848 17128
rect 23900 17116 23906 17128
rect 23937 17119 23995 17125
rect 23937 17116 23949 17119
rect 23900 17088 23949 17116
rect 23900 17076 23906 17088
rect 23937 17085 23949 17088
rect 23983 17085 23995 17119
rect 24486 17116 24492 17128
rect 24399 17088 24492 17116
rect 23937 17079 23995 17085
rect 24486 17076 24492 17088
rect 24544 17076 24550 17128
rect 24857 17119 24915 17125
rect 24857 17085 24869 17119
rect 24903 17116 24915 17119
rect 24946 17116 24952 17128
rect 24903 17088 24952 17116
rect 24903 17085 24915 17088
rect 24857 17079 24915 17085
rect 24946 17076 24952 17088
rect 25004 17076 25010 17128
rect 25774 17116 25780 17128
rect 25735 17088 25780 17116
rect 25774 17076 25780 17088
rect 25832 17076 25838 17128
rect 26160 17125 26188 17156
rect 26418 17144 26424 17156
rect 26476 17144 26482 17196
rect 29457 17187 29515 17193
rect 29457 17153 29469 17187
rect 29503 17184 29515 17187
rect 29822 17184 29828 17196
rect 29503 17156 29828 17184
rect 29503 17153 29515 17156
rect 29457 17147 29515 17153
rect 29822 17144 29828 17156
rect 29880 17144 29886 17196
rect 31202 17184 31208 17196
rect 30392 17156 31208 17184
rect 26145 17119 26203 17125
rect 26145 17085 26157 17119
rect 26191 17085 26203 17119
rect 26510 17116 26516 17128
rect 26471 17088 26516 17116
rect 26145 17079 26203 17085
rect 26510 17076 26516 17088
rect 26568 17076 26574 17128
rect 26694 17116 26700 17128
rect 26655 17088 26700 17116
rect 26694 17076 26700 17088
rect 26752 17076 26758 17128
rect 27157 17119 27215 17125
rect 27157 17085 27169 17119
rect 27203 17085 27215 17119
rect 28166 17116 28172 17128
rect 28127 17088 28172 17116
rect 27157 17079 27215 17085
rect 24394 17048 24400 17060
rect 21928 17020 24400 17048
rect 24394 17008 24400 17020
rect 24452 17008 24458 17060
rect 24504 17048 24532 17076
rect 27172 17048 27200 17079
rect 28166 17076 28172 17088
rect 28224 17076 28230 17128
rect 28258 17076 28264 17128
rect 28316 17116 28322 17128
rect 29638 17116 29644 17128
rect 28316 17088 29644 17116
rect 28316 17076 28322 17088
rect 29638 17076 29644 17088
rect 29696 17076 29702 17128
rect 29917 17119 29975 17125
rect 29917 17085 29929 17119
rect 29963 17085 29975 17119
rect 30098 17116 30104 17128
rect 30059 17088 30104 17116
rect 29917 17079 29975 17085
rect 24504 17020 27200 17048
rect 28077 17051 28135 17057
rect 28077 17017 28089 17051
rect 28123 17048 28135 17051
rect 28350 17048 28356 17060
rect 28123 17020 28356 17048
rect 28123 17017 28135 17020
rect 28077 17011 28135 17017
rect 28350 17008 28356 17020
rect 28408 17008 28414 17060
rect 21269 16983 21327 16989
rect 21269 16949 21281 16983
rect 21315 16949 21327 16983
rect 21269 16943 21327 16949
rect 23293 16983 23351 16989
rect 23293 16949 23305 16983
rect 23339 16980 23351 16983
rect 23934 16980 23940 16992
rect 23339 16952 23940 16980
rect 23339 16949 23351 16952
rect 23293 16943 23351 16949
rect 23934 16940 23940 16952
rect 23992 16980 23998 16992
rect 24578 16980 24584 16992
rect 23992 16952 24584 16980
rect 23992 16940 23998 16952
rect 24578 16940 24584 16952
rect 24636 16940 24642 16992
rect 27430 16940 27436 16992
rect 27488 16980 27494 16992
rect 29932 16980 29960 17079
rect 30098 17076 30104 17088
rect 30156 17076 30162 17128
rect 30392 17125 30420 17156
rect 31202 17144 31208 17156
rect 31260 17184 31266 17196
rect 31260 17156 32168 17184
rect 31260 17144 31266 17156
rect 30377 17119 30435 17125
rect 30377 17085 30389 17119
rect 30423 17085 30435 17119
rect 30377 17079 30435 17085
rect 30469 17119 30527 17125
rect 30469 17085 30481 17119
rect 30515 17085 30527 17119
rect 30469 17079 30527 17085
rect 30484 17048 30512 17079
rect 30558 17076 30564 17128
rect 30616 17116 30622 17128
rect 30745 17119 30803 17125
rect 30745 17116 30757 17119
rect 30616 17088 30757 17116
rect 30616 17076 30622 17088
rect 30745 17085 30757 17088
rect 30791 17085 30803 17119
rect 30745 17079 30803 17085
rect 30650 17048 30656 17060
rect 30484 17020 30656 17048
rect 30650 17008 30656 17020
rect 30708 17008 30714 17060
rect 27488 16952 29960 16980
rect 30760 16980 30788 17079
rect 31018 17076 31024 17128
rect 31076 17116 31082 17128
rect 31389 17119 31447 17125
rect 31389 17116 31401 17119
rect 31076 17088 31401 17116
rect 31076 17076 31082 17088
rect 31389 17085 31401 17088
rect 31435 17085 31447 17119
rect 31389 17079 31447 17085
rect 31754 17076 31760 17128
rect 31812 17116 31818 17128
rect 32140 17125 32168 17156
rect 33428 17125 33456 17224
rect 33502 17144 33508 17196
rect 33560 17184 33566 17196
rect 34057 17187 34115 17193
rect 34057 17184 34069 17187
rect 33560 17156 34069 17184
rect 33560 17144 33566 17156
rect 34057 17153 34069 17156
rect 34103 17153 34115 17187
rect 34057 17147 34115 17153
rect 32125 17119 32183 17125
rect 31812 17088 31857 17116
rect 31812 17076 31818 17088
rect 32125 17085 32137 17119
rect 32171 17085 32183 17119
rect 32125 17079 32183 17085
rect 33413 17119 33471 17125
rect 33413 17085 33425 17119
rect 33459 17085 33471 17119
rect 33413 17079 33471 17085
rect 33781 17119 33839 17125
rect 33781 17085 33793 17119
rect 33827 17116 33839 17119
rect 34330 17116 34336 17128
rect 33827 17088 34336 17116
rect 33827 17085 33839 17088
rect 33781 17079 33839 17085
rect 32585 17051 32643 17057
rect 32585 17017 32597 17051
rect 32631 17048 32643 17051
rect 32950 17048 32956 17060
rect 32631 17020 32956 17048
rect 32631 17017 32643 17020
rect 32585 17011 32643 17017
rect 32950 17008 32956 17020
rect 33008 17008 33014 17060
rect 33796 17048 33824 17079
rect 34330 17076 34336 17088
rect 34388 17076 34394 17128
rect 35084 17125 35112 17224
rect 35161 17221 35173 17255
rect 35207 17221 35219 17255
rect 35161 17215 35219 17221
rect 35176 17184 35204 17215
rect 36725 17187 36783 17193
rect 36725 17184 36737 17187
rect 35176 17156 36737 17184
rect 36725 17153 36737 17156
rect 36771 17153 36783 17187
rect 36725 17147 36783 17153
rect 37734 17144 37740 17196
rect 37792 17184 37798 17196
rect 37829 17187 37887 17193
rect 37829 17184 37841 17187
rect 37792 17156 37841 17184
rect 37792 17144 37798 17156
rect 37829 17153 37841 17156
rect 37875 17153 37887 17187
rect 37829 17147 37887 17153
rect 35069 17119 35127 17125
rect 35069 17085 35081 17119
rect 35115 17116 35127 17119
rect 35621 17119 35679 17125
rect 35115 17088 35204 17116
rect 35115 17085 35127 17088
rect 35069 17079 35127 17085
rect 33244 17020 33824 17048
rect 33244 16980 33272 17020
rect 30760 16952 33272 16980
rect 33321 16983 33379 16989
rect 27488 16940 27494 16952
rect 33321 16949 33333 16983
rect 33367 16980 33379 16983
rect 34790 16980 34796 16992
rect 33367 16952 34796 16980
rect 33367 16949 33379 16952
rect 33321 16943 33379 16949
rect 34790 16940 34796 16952
rect 34848 16940 34854 16992
rect 35176 16980 35204 17088
rect 35621 17085 35633 17119
rect 35667 17085 35679 17119
rect 35621 17079 35679 17085
rect 35805 17119 35863 17125
rect 35805 17085 35817 17119
rect 35851 17116 35863 17119
rect 35986 17116 35992 17128
rect 35851 17088 35992 17116
rect 35851 17085 35863 17088
rect 35805 17079 35863 17085
rect 35636 17048 35664 17079
rect 35986 17076 35992 17088
rect 36044 17076 36050 17128
rect 36262 17076 36268 17128
rect 36320 17116 36326 17128
rect 36449 17119 36507 17125
rect 36449 17116 36461 17119
rect 36320 17088 36461 17116
rect 36320 17076 36326 17088
rect 36449 17085 36461 17088
rect 36495 17085 36507 17119
rect 36449 17079 36507 17085
rect 36538 17048 36544 17060
rect 35636 17020 36544 17048
rect 36538 17008 36544 17020
rect 36596 17008 36602 17060
rect 36078 16980 36084 16992
rect 35176 16952 36084 16980
rect 36078 16940 36084 16952
rect 36136 16940 36142 16992
rect 1104 16890 38824 16912
rect 1104 16838 19606 16890
rect 19658 16838 19670 16890
rect 19722 16838 19734 16890
rect 19786 16838 19798 16890
rect 19850 16838 38824 16890
rect 1104 16816 38824 16838
rect 2961 16779 3019 16785
rect 2961 16745 2973 16779
rect 3007 16776 3019 16779
rect 3050 16776 3056 16788
rect 3007 16748 3056 16776
rect 3007 16745 3019 16748
rect 2961 16739 3019 16745
rect 3050 16736 3056 16748
rect 3108 16736 3114 16788
rect 3142 16736 3148 16788
rect 3200 16776 3206 16788
rect 7929 16779 7987 16785
rect 3200 16748 5856 16776
rect 3200 16736 3206 16748
rect 5626 16708 5632 16720
rect 5368 16680 5632 16708
rect 1670 16640 1676 16652
rect 1631 16612 1676 16640
rect 1670 16600 1676 16612
rect 1728 16600 1734 16652
rect 4154 16640 4160 16652
rect 4115 16612 4160 16640
rect 4154 16600 4160 16612
rect 4212 16600 4218 16652
rect 5368 16640 5396 16680
rect 5626 16668 5632 16680
rect 5684 16668 5690 16720
rect 5534 16640 5540 16652
rect 4264 16612 5396 16640
rect 5495 16612 5540 16640
rect 1394 16572 1400 16584
rect 1355 16544 1400 16572
rect 1394 16532 1400 16544
rect 1452 16532 1458 16584
rect 4065 16575 4123 16581
rect 4065 16541 4077 16575
rect 4111 16572 4123 16575
rect 4264 16572 4292 16612
rect 5534 16600 5540 16612
rect 5592 16600 5598 16652
rect 5442 16572 5448 16584
rect 4111 16544 4292 16572
rect 5403 16544 5448 16572
rect 4111 16541 4123 16544
rect 4065 16535 4123 16541
rect 5442 16532 5448 16544
rect 5500 16532 5506 16584
rect 5828 16572 5856 16748
rect 7929 16745 7941 16779
rect 7975 16776 7987 16779
rect 8018 16776 8024 16788
rect 7975 16748 8024 16776
rect 7975 16745 7987 16748
rect 7929 16739 7987 16745
rect 8018 16736 8024 16748
rect 8076 16736 8082 16788
rect 8938 16776 8944 16788
rect 8899 16748 8944 16776
rect 8938 16736 8944 16748
rect 8996 16736 9002 16788
rect 12802 16776 12808 16788
rect 10244 16748 12808 16776
rect 5902 16668 5908 16720
rect 5960 16708 5966 16720
rect 10244 16717 10272 16748
rect 12802 16736 12808 16748
rect 12860 16736 12866 16788
rect 21266 16776 21272 16788
rect 14200 16748 21272 16776
rect 10229 16711 10287 16717
rect 5960 16680 8892 16708
rect 5960 16668 5966 16680
rect 5994 16640 6000 16652
rect 5955 16612 6000 16640
rect 5994 16600 6000 16612
rect 6052 16600 6058 16652
rect 6457 16643 6515 16649
rect 6457 16640 6469 16643
rect 6104 16612 6469 16640
rect 6104 16572 6132 16612
rect 6457 16609 6469 16612
rect 6503 16640 6515 16643
rect 7009 16643 7067 16649
rect 6503 16612 6960 16640
rect 6503 16609 6515 16612
rect 6457 16603 6515 16609
rect 5828 16544 6132 16572
rect 6932 16504 6960 16612
rect 7009 16609 7021 16643
rect 7055 16640 7067 16643
rect 7558 16640 7564 16652
rect 7055 16612 7564 16640
rect 7055 16609 7067 16612
rect 7009 16603 7067 16609
rect 7558 16600 7564 16612
rect 7616 16600 7622 16652
rect 8864 16649 8892 16680
rect 8956 16680 10180 16708
rect 7653 16643 7711 16649
rect 7653 16609 7665 16643
rect 7699 16609 7711 16643
rect 7653 16603 7711 16609
rect 8205 16643 8263 16649
rect 8205 16609 8217 16643
rect 8251 16640 8263 16643
rect 8849 16643 8907 16649
rect 8251 16612 8800 16640
rect 8251 16609 8263 16612
rect 8205 16603 8263 16609
rect 7098 16572 7104 16584
rect 7059 16544 7104 16572
rect 7098 16532 7104 16544
rect 7156 16532 7162 16584
rect 7668 16572 7696 16603
rect 7576 16544 7696 16572
rect 8772 16572 8800 16612
rect 8849 16609 8861 16643
rect 8895 16609 8907 16643
rect 8849 16603 8907 16609
rect 8956 16572 8984 16680
rect 9766 16640 9772 16652
rect 9727 16612 9772 16640
rect 9766 16600 9772 16612
rect 9824 16600 9830 16652
rect 10152 16640 10180 16680
rect 10229 16677 10241 16711
rect 10275 16677 10287 16711
rect 11238 16708 11244 16720
rect 10229 16671 10287 16677
rect 10980 16680 11244 16708
rect 10980 16649 11008 16680
rect 11238 16668 11244 16680
rect 11296 16668 11302 16720
rect 10965 16643 11023 16649
rect 10152 16612 10916 16640
rect 9674 16572 9680 16584
rect 8772 16544 8984 16572
rect 9635 16544 9680 16572
rect 7576 16504 7604 16544
rect 9674 16532 9680 16544
rect 9732 16532 9738 16584
rect 6932 16476 7604 16504
rect 10888 16504 10916 16612
rect 10965 16609 10977 16643
rect 11011 16609 11023 16643
rect 11422 16640 11428 16652
rect 11383 16612 11428 16640
rect 10965 16603 11023 16609
rect 11422 16600 11428 16612
rect 11480 16600 11486 16652
rect 11793 16643 11851 16649
rect 11793 16609 11805 16643
rect 11839 16640 11851 16643
rect 12434 16640 12440 16652
rect 11839 16612 12440 16640
rect 11839 16609 11851 16612
rect 11793 16603 11851 16609
rect 12434 16600 12440 16612
rect 12492 16600 12498 16652
rect 12710 16640 12716 16652
rect 12671 16612 12716 16640
rect 12710 16600 12716 16612
rect 12768 16600 12774 16652
rect 12989 16643 13047 16649
rect 12989 16609 13001 16643
rect 13035 16640 13047 16643
rect 14200 16640 14228 16748
rect 21266 16736 21272 16748
rect 21324 16736 21330 16788
rect 25774 16776 25780 16788
rect 25687 16748 25780 16776
rect 25774 16736 25780 16748
rect 25832 16776 25838 16788
rect 26142 16776 26148 16788
rect 25832 16748 26148 16776
rect 25832 16736 25838 16748
rect 26142 16736 26148 16748
rect 26200 16736 26206 16788
rect 30834 16776 30840 16788
rect 27264 16748 30840 16776
rect 22002 16708 22008 16720
rect 19812 16680 22008 16708
rect 14366 16640 14372 16652
rect 13035 16612 14228 16640
rect 14327 16612 14372 16640
rect 13035 16609 13047 16612
rect 12989 16603 13047 16609
rect 14366 16600 14372 16612
rect 14424 16600 14430 16652
rect 16114 16640 16120 16652
rect 16075 16612 16120 16640
rect 16114 16600 16120 16612
rect 16172 16600 16178 16652
rect 16390 16640 16396 16652
rect 16351 16612 16396 16640
rect 16390 16600 16396 16612
rect 16448 16600 16454 16652
rect 16482 16600 16488 16652
rect 16540 16640 16546 16652
rect 17313 16643 17371 16649
rect 16540 16612 17172 16640
rect 16540 16600 16546 16612
rect 11054 16572 11060 16584
rect 11015 16544 11060 16572
rect 11054 16532 11060 16544
rect 11112 16532 11118 16584
rect 17037 16575 17095 16581
rect 17037 16541 17049 16575
rect 17083 16541 17095 16575
rect 17144 16572 17172 16612
rect 17313 16609 17325 16643
rect 17359 16640 17371 16643
rect 18506 16640 18512 16652
rect 17359 16612 18512 16640
rect 17359 16609 17371 16612
rect 17313 16603 17371 16609
rect 18506 16600 18512 16612
rect 18564 16600 18570 16652
rect 19812 16649 19840 16680
rect 22002 16668 22008 16680
rect 22060 16668 22066 16720
rect 23566 16668 23572 16720
rect 23624 16708 23630 16720
rect 27264 16708 27292 16748
rect 30834 16736 30840 16748
rect 30892 16736 30898 16788
rect 32582 16736 32588 16788
rect 32640 16776 32646 16788
rect 35897 16779 35955 16785
rect 35897 16776 35909 16779
rect 32640 16748 35909 16776
rect 32640 16736 32646 16748
rect 29825 16711 29883 16717
rect 29825 16708 29837 16711
rect 23624 16680 27292 16708
rect 27356 16680 29837 16708
rect 23624 16668 23630 16680
rect 19153 16643 19211 16649
rect 19153 16640 19165 16643
rect 18616 16612 19165 16640
rect 18616 16572 18644 16612
rect 19153 16609 19165 16612
rect 19199 16609 19211 16643
rect 19153 16603 19211 16609
rect 19797 16643 19855 16649
rect 19797 16609 19809 16643
rect 19843 16609 19855 16643
rect 19797 16603 19855 16609
rect 20165 16643 20223 16649
rect 20165 16609 20177 16643
rect 20211 16640 20223 16643
rect 20714 16640 20720 16652
rect 20211 16612 20720 16640
rect 20211 16609 20223 16612
rect 20165 16603 20223 16609
rect 20714 16600 20720 16612
rect 20772 16600 20778 16652
rect 21082 16640 21088 16652
rect 21043 16612 21088 16640
rect 21082 16600 21088 16612
rect 21140 16600 21146 16652
rect 21174 16600 21180 16652
rect 21232 16640 21238 16652
rect 21545 16643 21603 16649
rect 21545 16640 21557 16643
rect 21232 16612 21557 16640
rect 21232 16600 21238 16612
rect 21545 16609 21557 16612
rect 21591 16609 21603 16643
rect 21818 16640 21824 16652
rect 21779 16612 21824 16640
rect 21545 16603 21603 16609
rect 21818 16600 21824 16612
rect 21876 16600 21882 16652
rect 21913 16643 21971 16649
rect 21913 16609 21925 16643
rect 21959 16609 21971 16643
rect 22186 16640 22192 16652
rect 22147 16612 22192 16640
rect 21913 16603 21971 16609
rect 19426 16572 19432 16584
rect 17144 16544 18644 16572
rect 18984 16544 19432 16572
rect 17037 16535 17095 16541
rect 11790 16504 11796 16516
rect 10888 16476 11796 16504
rect 11790 16464 11796 16476
rect 11848 16464 11854 16516
rect 15286 16464 15292 16516
rect 15344 16504 15350 16516
rect 15933 16507 15991 16513
rect 15933 16504 15945 16507
rect 15344 16476 15945 16504
rect 15344 16464 15350 16476
rect 15933 16473 15945 16476
rect 15979 16473 15991 16507
rect 15933 16467 15991 16473
rect 1854 16396 1860 16448
rect 1912 16436 1918 16448
rect 4341 16439 4399 16445
rect 4341 16436 4353 16439
rect 1912 16408 4353 16436
rect 1912 16396 1918 16408
rect 4341 16405 4353 16408
rect 4387 16405 4399 16439
rect 4341 16399 4399 16405
rect 12618 16396 12624 16448
rect 12676 16436 12682 16448
rect 16942 16436 16948 16448
rect 12676 16408 16948 16436
rect 12676 16396 12682 16408
rect 16942 16396 16948 16408
rect 17000 16396 17006 16448
rect 17052 16436 17080 16535
rect 18046 16464 18052 16516
rect 18104 16504 18110 16516
rect 18984 16504 19012 16544
rect 19426 16532 19432 16544
rect 19484 16532 19490 16584
rect 21928 16572 21956 16603
rect 22186 16600 22192 16612
rect 22244 16600 22250 16652
rect 22462 16640 22468 16652
rect 22423 16612 22468 16640
rect 22462 16600 22468 16612
rect 22520 16600 22526 16652
rect 23198 16640 23204 16652
rect 23159 16612 23204 16640
rect 23198 16600 23204 16612
rect 23256 16600 23262 16652
rect 23658 16640 23664 16652
rect 23619 16612 23664 16640
rect 23658 16600 23664 16612
rect 23716 16600 23722 16652
rect 24118 16640 24124 16652
rect 24079 16612 24124 16640
rect 24118 16600 24124 16612
rect 24176 16600 24182 16652
rect 24670 16640 24676 16652
rect 24631 16612 24676 16640
rect 24670 16600 24676 16612
rect 24728 16600 24734 16652
rect 24854 16640 24860 16652
rect 24815 16612 24860 16640
rect 24854 16600 24860 16612
rect 24912 16600 24918 16652
rect 24946 16600 24952 16652
rect 25004 16640 25010 16652
rect 25593 16643 25651 16649
rect 25593 16640 25605 16643
rect 25004 16612 25605 16640
rect 25004 16600 25010 16612
rect 25593 16609 25605 16612
rect 25639 16640 25651 16643
rect 25682 16640 25688 16652
rect 25639 16612 25688 16640
rect 25639 16609 25651 16612
rect 25593 16603 25651 16609
rect 25682 16600 25688 16612
rect 25740 16600 25746 16652
rect 26510 16640 26516 16652
rect 26471 16612 26516 16640
rect 26510 16600 26516 16612
rect 26568 16600 26574 16652
rect 27356 16649 27384 16680
rect 29825 16677 29837 16680
rect 29871 16708 29883 16711
rect 30098 16708 30104 16720
rect 29871 16680 30104 16708
rect 29871 16677 29883 16680
rect 29825 16671 29883 16677
rect 30098 16668 30104 16680
rect 30156 16668 30162 16720
rect 32030 16668 32036 16720
rect 32088 16708 32094 16720
rect 32088 16680 32904 16708
rect 32088 16668 32094 16680
rect 27341 16643 27399 16649
rect 27341 16609 27353 16643
rect 27387 16609 27399 16643
rect 27614 16640 27620 16652
rect 27341 16603 27399 16609
rect 27448 16612 27620 16640
rect 21928 16544 23244 16572
rect 23216 16516 23244 16544
rect 18104 16476 19012 16504
rect 18104 16464 18110 16476
rect 19058 16464 19064 16516
rect 19116 16504 19122 16516
rect 19116 16476 21312 16504
rect 19116 16464 19122 16476
rect 18138 16436 18144 16448
rect 17052 16408 18144 16436
rect 18138 16396 18144 16408
rect 18196 16396 18202 16448
rect 18601 16439 18659 16445
rect 18601 16405 18613 16439
rect 18647 16436 18659 16439
rect 18782 16436 18788 16448
rect 18647 16408 18788 16436
rect 18647 16405 18659 16408
rect 18601 16399 18659 16405
rect 18782 16396 18788 16408
rect 18840 16396 18846 16448
rect 18966 16396 18972 16448
rect 19024 16436 19030 16448
rect 19245 16439 19303 16445
rect 19245 16436 19257 16439
rect 19024 16408 19257 16436
rect 19024 16396 19030 16408
rect 19245 16405 19257 16408
rect 19291 16405 19303 16439
rect 21284 16436 21312 16476
rect 23198 16464 23204 16516
rect 23256 16464 23262 16516
rect 23293 16507 23351 16513
rect 23293 16473 23305 16507
rect 23339 16473 23351 16507
rect 23293 16467 23351 16473
rect 23308 16436 23336 16467
rect 25498 16464 25504 16516
rect 25556 16504 25562 16516
rect 27448 16513 27476 16612
rect 27614 16600 27620 16612
rect 27672 16600 27678 16652
rect 27798 16640 27804 16652
rect 27759 16612 27804 16640
rect 27798 16600 27804 16612
rect 27856 16600 27862 16652
rect 29273 16643 29331 16649
rect 29273 16640 29285 16643
rect 28736 16612 29285 16640
rect 28166 16572 28172 16584
rect 28079 16544 28172 16572
rect 28166 16532 28172 16544
rect 28224 16572 28230 16584
rect 28736 16572 28764 16612
rect 29273 16609 29285 16612
rect 29319 16640 29331 16643
rect 29454 16640 29460 16652
rect 29319 16612 29460 16640
rect 29319 16609 29331 16612
rect 29273 16603 29331 16609
rect 29454 16600 29460 16612
rect 29512 16600 29518 16652
rect 29638 16640 29644 16652
rect 29599 16612 29644 16640
rect 29638 16600 29644 16612
rect 29696 16600 29702 16652
rect 31110 16640 31116 16652
rect 31071 16612 31116 16640
rect 31110 16600 31116 16612
rect 31168 16600 31174 16652
rect 31573 16643 31631 16649
rect 31573 16609 31585 16643
rect 31619 16609 31631 16643
rect 31573 16603 31631 16609
rect 28224 16544 28764 16572
rect 28905 16575 28963 16581
rect 28224 16532 28230 16544
rect 28905 16541 28917 16575
rect 28951 16572 28963 16575
rect 28994 16572 29000 16584
rect 28951 16544 29000 16572
rect 28951 16541 28963 16544
rect 28905 16535 28963 16541
rect 28994 16532 29000 16544
rect 29052 16532 29058 16584
rect 31205 16575 31263 16581
rect 31205 16541 31217 16575
rect 31251 16541 31263 16575
rect 31588 16572 31616 16603
rect 31662 16600 31668 16652
rect 31720 16640 31726 16652
rect 32876 16649 32904 16680
rect 32309 16643 32367 16649
rect 32309 16640 32321 16643
rect 31720 16612 32321 16640
rect 31720 16600 31726 16612
rect 32309 16609 32321 16612
rect 32355 16609 32367 16643
rect 32309 16603 32367 16609
rect 32861 16643 32919 16649
rect 32861 16609 32873 16643
rect 32907 16609 32919 16643
rect 32968 16640 32996 16748
rect 35897 16745 35909 16748
rect 35943 16776 35955 16779
rect 35986 16776 35992 16788
rect 35943 16748 35992 16776
rect 35943 16745 35955 16748
rect 35897 16739 35955 16745
rect 35986 16736 35992 16748
rect 36044 16776 36050 16788
rect 36817 16779 36875 16785
rect 36817 16776 36829 16779
rect 36044 16748 36676 16776
rect 36044 16736 36050 16748
rect 33042 16668 33048 16720
rect 33100 16708 33106 16720
rect 33100 16680 33824 16708
rect 33100 16668 33106 16680
rect 33137 16643 33195 16649
rect 32968 16612 33088 16640
rect 32861 16603 32919 16609
rect 32490 16572 32496 16584
rect 31588 16544 32496 16572
rect 31205 16535 31263 16541
rect 27433 16507 27491 16513
rect 25556 16476 26740 16504
rect 25556 16464 25562 16476
rect 26602 16436 26608 16448
rect 21284 16408 23336 16436
rect 26563 16408 26608 16436
rect 19245 16399 19303 16405
rect 26602 16396 26608 16408
rect 26660 16396 26666 16448
rect 26712 16436 26740 16476
rect 27433 16473 27445 16507
rect 27479 16473 27491 16507
rect 31220 16504 31248 16535
rect 32490 16532 32496 16544
rect 32548 16532 32554 16584
rect 33060 16572 33088 16612
rect 33137 16609 33149 16643
rect 33183 16640 33195 16643
rect 33410 16640 33416 16652
rect 33183 16612 33416 16640
rect 33183 16609 33195 16612
rect 33137 16603 33195 16609
rect 33410 16600 33416 16612
rect 33468 16600 33474 16652
rect 33796 16649 33824 16680
rect 33781 16643 33839 16649
rect 33781 16609 33793 16643
rect 33827 16609 33839 16643
rect 34514 16640 34520 16652
rect 34475 16612 34520 16640
rect 33781 16603 33839 16609
rect 34514 16600 34520 16612
rect 34572 16600 34578 16652
rect 34790 16640 34796 16652
rect 34751 16612 34796 16640
rect 34790 16600 34796 16612
rect 34848 16600 34854 16652
rect 35434 16600 35440 16652
rect 35492 16640 35498 16652
rect 36648 16649 36676 16748
rect 36740 16748 36829 16776
rect 36633 16643 36691 16649
rect 35492 16612 36584 16640
rect 35492 16600 35498 16612
rect 33318 16572 33324 16584
rect 33060 16544 33324 16572
rect 33318 16532 33324 16544
rect 33376 16532 33382 16584
rect 36556 16572 36584 16612
rect 36633 16609 36645 16643
rect 36679 16609 36691 16643
rect 36633 16603 36691 16609
rect 36740 16572 36768 16748
rect 36817 16745 36829 16748
rect 36863 16745 36875 16779
rect 36817 16739 36875 16745
rect 37737 16643 37795 16649
rect 37737 16609 37749 16643
rect 37783 16640 37795 16643
rect 38102 16640 38108 16652
rect 37783 16612 38108 16640
rect 37783 16609 37795 16612
rect 37737 16603 37795 16609
rect 38102 16600 38108 16612
rect 38160 16600 38166 16652
rect 36556 16544 36768 16572
rect 33502 16504 33508 16516
rect 31220 16476 33508 16504
rect 27433 16467 27491 16473
rect 33502 16464 33508 16476
rect 33560 16464 33566 16516
rect 33962 16504 33968 16516
rect 33923 16476 33968 16504
rect 33962 16464 33968 16476
rect 34020 16464 34026 16516
rect 29270 16436 29276 16448
rect 26712 16408 29276 16436
rect 29270 16396 29276 16408
rect 29328 16396 29334 16448
rect 37918 16436 37924 16448
rect 37879 16408 37924 16436
rect 37918 16396 37924 16408
rect 37976 16396 37982 16448
rect 1104 16346 38824 16368
rect 1104 16294 4246 16346
rect 4298 16294 4310 16346
rect 4362 16294 4374 16346
rect 4426 16294 4438 16346
rect 4490 16294 34966 16346
rect 35018 16294 35030 16346
rect 35082 16294 35094 16346
rect 35146 16294 35158 16346
rect 35210 16294 38824 16346
rect 1104 16272 38824 16294
rect 3513 16235 3571 16241
rect 3513 16201 3525 16235
rect 3559 16232 3571 16235
rect 4062 16232 4068 16244
rect 3559 16204 4068 16232
rect 3559 16201 3571 16204
rect 3513 16195 3571 16201
rect 4062 16192 4068 16204
rect 4120 16192 4126 16244
rect 5534 16192 5540 16244
rect 5592 16232 5598 16244
rect 5629 16235 5687 16241
rect 5629 16232 5641 16235
rect 5592 16204 5641 16232
rect 5592 16192 5598 16204
rect 5629 16201 5641 16204
rect 5675 16201 5687 16235
rect 8386 16232 8392 16244
rect 8347 16204 8392 16232
rect 5629 16195 5687 16201
rect 8386 16192 8392 16204
rect 8444 16192 8450 16244
rect 11149 16235 11207 16241
rect 11149 16201 11161 16235
rect 11195 16232 11207 16235
rect 11238 16232 11244 16244
rect 11195 16204 11244 16232
rect 11195 16201 11207 16204
rect 11149 16195 11207 16201
rect 11238 16192 11244 16204
rect 11296 16192 11302 16244
rect 11790 16232 11796 16244
rect 11751 16204 11796 16232
rect 11790 16192 11796 16204
rect 11848 16192 11854 16244
rect 15197 16235 15255 16241
rect 15197 16201 15209 16235
rect 15243 16232 15255 16235
rect 16114 16232 16120 16244
rect 15243 16204 16120 16232
rect 15243 16201 15255 16204
rect 15197 16195 15255 16201
rect 16114 16192 16120 16204
rect 16172 16232 16178 16244
rect 18046 16232 18052 16244
rect 16172 16204 18052 16232
rect 16172 16192 16178 16204
rect 18046 16192 18052 16204
rect 18104 16192 18110 16244
rect 18233 16235 18291 16241
rect 18233 16201 18245 16235
rect 18279 16232 18291 16235
rect 19242 16232 19248 16244
rect 18279 16204 19248 16232
rect 18279 16201 18291 16204
rect 18233 16195 18291 16201
rect 19242 16192 19248 16204
rect 19300 16192 19306 16244
rect 20714 16192 20720 16244
rect 20772 16232 20778 16244
rect 24121 16235 24179 16241
rect 24121 16232 24133 16235
rect 20772 16204 24133 16232
rect 20772 16192 20778 16204
rect 24121 16201 24133 16204
rect 24167 16201 24179 16235
rect 24121 16195 24179 16201
rect 25869 16235 25927 16241
rect 25869 16201 25881 16235
rect 25915 16232 25927 16235
rect 27430 16232 27436 16244
rect 25915 16204 27436 16232
rect 25915 16201 25927 16204
rect 25869 16195 25927 16201
rect 27430 16192 27436 16204
rect 27488 16192 27494 16244
rect 30742 16232 30748 16244
rect 28460 16204 30748 16232
rect 23106 16164 23112 16176
rect 21192 16136 23112 16164
rect 4249 16099 4307 16105
rect 4249 16096 4261 16099
rect 1964 16068 4261 16096
rect 1394 15988 1400 16040
rect 1452 16028 1458 16040
rect 1964 16037 1992 16068
rect 4249 16065 4261 16068
rect 4295 16096 4307 16099
rect 5350 16096 5356 16108
rect 4295 16068 5356 16096
rect 4295 16065 4307 16068
rect 4249 16059 4307 16065
rect 5350 16056 5356 16068
rect 5408 16056 5414 16108
rect 7098 16096 7104 16108
rect 7059 16068 7104 16096
rect 7098 16056 7104 16068
rect 7156 16056 7162 16108
rect 9861 16099 9919 16105
rect 9324 16068 9720 16096
rect 1949 16031 2007 16037
rect 1949 16028 1961 16031
rect 1452 16000 1961 16028
rect 1452 15988 1458 16000
rect 1949 15997 1961 16000
rect 1995 15997 2007 16031
rect 1949 15991 2007 15997
rect 2225 16031 2283 16037
rect 2225 15997 2237 16031
rect 2271 16028 2283 16031
rect 2682 16028 2688 16040
rect 2271 16000 2688 16028
rect 2271 15997 2283 16000
rect 2225 15991 2283 15997
rect 2682 15988 2688 16000
rect 2740 15988 2746 16040
rect 4522 16028 4528 16040
rect 4483 16000 4528 16028
rect 4522 15988 4528 16000
rect 4580 15988 4586 16040
rect 6825 16031 6883 16037
rect 6825 15997 6837 16031
rect 6871 16028 6883 16031
rect 7742 16028 7748 16040
rect 6871 16000 7748 16028
rect 6871 15997 6883 16000
rect 6825 15991 6883 15997
rect 7742 15988 7748 16000
rect 7800 16028 7806 16040
rect 9324 16028 9352 16068
rect 7800 16000 9352 16028
rect 7800 15988 7806 16000
rect 9490 15988 9496 16040
rect 9548 16028 9554 16040
rect 9585 16031 9643 16037
rect 9585 16028 9597 16031
rect 9548 16000 9597 16028
rect 9548 15988 9554 16000
rect 9585 15997 9597 16000
rect 9631 15997 9643 16031
rect 9692 16028 9720 16068
rect 9861 16065 9873 16099
rect 9907 16096 9919 16099
rect 10686 16096 10692 16108
rect 9907 16068 10692 16096
rect 9907 16065 9919 16068
rect 9861 16059 9919 16065
rect 10686 16056 10692 16068
rect 10744 16056 10750 16108
rect 18785 16099 18843 16105
rect 18785 16096 18797 16099
rect 10796 16068 18797 16096
rect 10502 16028 10508 16040
rect 9692 16000 10508 16028
rect 9585 15991 9643 15997
rect 10502 15988 10508 16000
rect 10560 16028 10566 16040
rect 10796 16028 10824 16068
rect 18785 16065 18797 16068
rect 18831 16065 18843 16099
rect 21192 16096 21220 16136
rect 23106 16124 23112 16136
rect 23164 16124 23170 16176
rect 27062 16164 27068 16176
rect 25148 16136 27068 16164
rect 18785 16059 18843 16065
rect 18892 16068 21220 16096
rect 22281 16099 22339 16105
rect 10560 16000 10824 16028
rect 10560 15988 10566 16000
rect 11238 15988 11244 16040
rect 11296 16028 11302 16040
rect 11701 16031 11759 16037
rect 11701 16028 11713 16031
rect 11296 16000 11713 16028
rect 11296 15988 11302 16000
rect 11701 15997 11713 16000
rect 11747 15997 11759 16031
rect 11701 15991 11759 15997
rect 12434 15988 12440 16040
rect 12492 16028 12498 16040
rect 12713 16031 12771 16037
rect 12713 16028 12725 16031
rect 12492 16000 12725 16028
rect 12492 15988 12498 16000
rect 12713 15997 12725 16000
rect 12759 15997 12771 16031
rect 12713 15991 12771 15997
rect 12802 15988 12808 16040
rect 12860 16028 12866 16040
rect 13633 16031 13691 16037
rect 13633 16028 13645 16031
rect 12860 16000 13645 16028
rect 12860 15988 12866 16000
rect 13633 15997 13645 16000
rect 13679 15997 13691 16031
rect 13906 16028 13912 16040
rect 13867 16000 13912 16028
rect 13633 15991 13691 15997
rect 13906 15988 13912 16000
rect 13964 15988 13970 16040
rect 15102 15988 15108 16040
rect 15160 16028 15166 16040
rect 15749 16031 15807 16037
rect 15749 16028 15761 16031
rect 15160 16000 15761 16028
rect 15160 15988 15166 16000
rect 15749 15997 15761 16000
rect 15795 15997 15807 16031
rect 16022 16028 16028 16040
rect 15983 16000 16028 16028
rect 15749 15991 15807 15997
rect 16022 15988 16028 16000
rect 16080 15988 16086 16040
rect 17310 15988 17316 16040
rect 17368 16028 17374 16040
rect 18049 16031 18107 16037
rect 18049 16028 18061 16031
rect 17368 16000 18061 16028
rect 17368 15988 17374 16000
rect 18049 15997 18061 16000
rect 18095 16028 18107 16031
rect 18892 16028 18920 16068
rect 22281 16065 22293 16099
rect 22327 16096 22339 16099
rect 22646 16096 22652 16108
rect 22327 16068 22652 16096
rect 22327 16065 22339 16068
rect 22281 16059 22339 16065
rect 22646 16056 22652 16068
rect 22704 16056 22710 16108
rect 24762 16096 24768 16108
rect 24723 16068 24768 16096
rect 24762 16056 24768 16068
rect 24820 16056 24826 16108
rect 25148 16105 25176 16136
rect 27062 16124 27068 16136
rect 27120 16164 27126 16176
rect 27338 16164 27344 16176
rect 27120 16136 27344 16164
rect 27120 16124 27126 16136
rect 27338 16124 27344 16136
rect 27396 16124 27402 16176
rect 25133 16099 25191 16105
rect 25133 16065 25145 16099
rect 25179 16065 25191 16099
rect 25133 16059 25191 16065
rect 26436 16068 27660 16096
rect 19058 16028 19064 16040
rect 18095 16000 18920 16028
rect 19019 16000 19064 16028
rect 18095 15997 18107 16000
rect 18049 15991 18107 15997
rect 19058 15988 19064 16000
rect 19116 15988 19122 16040
rect 20898 16028 20904 16040
rect 20859 16000 20904 16028
rect 20898 15988 20904 16000
rect 20956 15988 20962 16040
rect 20993 16031 21051 16037
rect 20993 15997 21005 16031
rect 21039 15997 21051 16031
rect 21450 16028 21456 16040
rect 21411 16000 21456 16028
rect 20993 15991 21051 15997
rect 18138 15960 18144 15972
rect 10520 15932 13768 15960
rect 9858 15852 9864 15904
rect 9916 15892 9922 15904
rect 10520 15892 10548 15932
rect 9916 15864 10548 15892
rect 9916 15852 9922 15864
rect 12342 15852 12348 15904
rect 12400 15892 12406 15904
rect 12897 15895 12955 15901
rect 12897 15892 12909 15895
rect 12400 15864 12909 15892
rect 12400 15852 12406 15864
rect 12897 15861 12909 15864
rect 12943 15861 12955 15895
rect 13740 15892 13768 15932
rect 14936 15932 15884 15960
rect 14936 15892 14964 15932
rect 13740 15864 14964 15892
rect 15856 15892 15884 15932
rect 16776 15932 18144 15960
rect 16776 15892 16804 15932
rect 18138 15920 18144 15932
rect 18196 15920 18202 15972
rect 20441 15963 20499 15969
rect 20441 15929 20453 15963
rect 20487 15960 20499 15963
rect 21008 15960 21036 15991
rect 21450 15988 21456 16000
rect 21508 15988 21514 16040
rect 22005 16031 22063 16037
rect 22005 15997 22017 16031
rect 22051 15997 22063 16031
rect 22005 15991 22063 15997
rect 20487 15932 21036 15960
rect 22020 15960 22048 15991
rect 22186 15988 22192 16040
rect 22244 16028 22250 16040
rect 22465 16031 22523 16037
rect 22465 16028 22477 16031
rect 22244 16000 22477 16028
rect 22244 15988 22250 16000
rect 22465 15997 22477 16000
rect 22511 15997 22523 16031
rect 22465 15991 22523 15997
rect 24673 16031 24731 16037
rect 24673 15997 24685 16031
rect 24719 16028 24731 16031
rect 24946 16028 24952 16040
rect 24719 16000 24952 16028
rect 24719 15997 24731 16000
rect 24673 15991 24731 15997
rect 24946 15988 24952 16000
rect 25004 15988 25010 16040
rect 26436 16037 26464 16068
rect 25041 16031 25099 16037
rect 25041 15997 25053 16031
rect 25087 15997 25099 16031
rect 25041 15991 25099 15997
rect 25777 16031 25835 16037
rect 25777 15997 25789 16031
rect 25823 15997 25835 16031
rect 25777 15991 25835 15997
rect 26421 16031 26479 16037
rect 26421 15997 26433 16031
rect 26467 15997 26479 16031
rect 26421 15991 26479 15997
rect 26528 16000 27292 16028
rect 22094 15960 22100 15972
rect 22020 15932 22100 15960
rect 20487 15929 20499 15932
rect 20441 15923 20499 15929
rect 22094 15920 22100 15932
rect 22152 15920 22158 15972
rect 23198 15920 23204 15972
rect 23256 15960 23262 15972
rect 25056 15960 25084 15991
rect 23256 15932 25084 15960
rect 23256 15920 23262 15932
rect 15856 15864 16804 15892
rect 12897 15855 12955 15861
rect 16850 15852 16856 15904
rect 16908 15892 16914 15904
rect 17129 15895 17187 15901
rect 17129 15892 17141 15895
rect 16908 15864 17141 15892
rect 16908 15852 16914 15864
rect 17129 15861 17141 15864
rect 17175 15861 17187 15895
rect 18156 15892 18184 15920
rect 19978 15892 19984 15904
rect 18156 15864 19984 15892
rect 17129 15855 17187 15861
rect 19978 15852 19984 15864
rect 20036 15852 20042 15904
rect 25792 15892 25820 15991
rect 26528 15892 26556 16000
rect 27264 15960 27292 16000
rect 27338 15988 27344 16040
rect 27396 16028 27402 16040
rect 27433 16031 27491 16037
rect 27433 16028 27445 16031
rect 27396 16000 27445 16028
rect 27396 15988 27402 16000
rect 27433 15997 27445 16000
rect 27479 16028 27491 16031
rect 27522 16028 27528 16040
rect 27479 16000 27528 16028
rect 27479 15997 27491 16000
rect 27433 15991 27491 15997
rect 27522 15988 27528 16000
rect 27580 15988 27586 16040
rect 27632 16037 27660 16068
rect 27617 16031 27675 16037
rect 27617 15997 27629 16031
rect 27663 16028 27675 16031
rect 27982 16028 27988 16040
rect 27663 16000 27988 16028
rect 27663 15997 27675 16000
rect 27617 15991 27675 15997
rect 27982 15988 27988 16000
rect 28040 15988 28046 16040
rect 28460 16037 28488 16204
rect 30742 16192 30748 16204
rect 30800 16192 30806 16244
rect 32677 16235 32735 16241
rect 32677 16201 32689 16235
rect 32723 16232 32735 16235
rect 33042 16232 33048 16244
rect 32723 16204 33048 16232
rect 32723 16201 32735 16204
rect 32677 16195 32735 16201
rect 33042 16192 33048 16204
rect 33100 16192 33106 16244
rect 36538 16232 36544 16244
rect 36499 16204 36544 16232
rect 36538 16192 36544 16204
rect 36596 16192 36602 16244
rect 30190 16164 30196 16176
rect 30151 16136 30196 16164
rect 30190 16124 30196 16136
rect 30248 16124 30254 16176
rect 35710 16164 35716 16176
rect 33980 16136 35716 16164
rect 29457 16099 29515 16105
rect 29457 16065 29469 16099
rect 29503 16096 29515 16099
rect 31570 16096 31576 16108
rect 29503 16068 31576 16096
rect 29503 16065 29515 16068
rect 29457 16059 29515 16065
rect 31570 16056 31576 16068
rect 31628 16056 31634 16108
rect 33980 16105 34008 16136
rect 35710 16124 35716 16136
rect 35768 16124 35774 16176
rect 33965 16099 34023 16105
rect 33965 16065 33977 16099
rect 34011 16065 34023 16099
rect 34974 16096 34980 16108
rect 34935 16068 34980 16096
rect 33965 16059 34023 16065
rect 34974 16056 34980 16068
rect 35032 16056 35038 16108
rect 35986 16096 35992 16108
rect 35084 16068 35848 16096
rect 35947 16068 35992 16096
rect 28445 16031 28503 16037
rect 28445 15997 28457 16031
rect 28491 15997 28503 16031
rect 29730 16028 29736 16040
rect 29691 16000 29736 16028
rect 28445 15991 28503 15997
rect 29730 15988 29736 16000
rect 29788 15988 29794 16040
rect 30101 16031 30159 16037
rect 30101 15997 30113 16031
rect 30147 15997 30159 16031
rect 30101 15991 30159 15997
rect 28534 15960 28540 15972
rect 27264 15932 28540 15960
rect 28534 15920 28540 15932
rect 28592 15920 28598 15972
rect 29178 15920 29184 15972
rect 29236 15960 29242 15972
rect 30116 15960 30144 15991
rect 30190 15988 30196 16040
rect 30248 16028 30254 16040
rect 31113 16031 31171 16037
rect 31113 16028 31125 16031
rect 30248 16000 31125 16028
rect 30248 15988 30254 16000
rect 31113 15997 31125 16000
rect 31159 15997 31171 16031
rect 31386 16028 31392 16040
rect 31347 16000 31392 16028
rect 31113 15991 31171 15997
rect 31386 15988 31392 16000
rect 31444 15988 31450 16040
rect 33318 16028 33324 16040
rect 33279 16000 33324 16028
rect 33318 15988 33324 16000
rect 33376 15988 33382 16040
rect 33410 15988 33416 16040
rect 33468 16028 33474 16040
rect 33781 16031 33839 16037
rect 33781 16028 33793 16031
rect 33468 16000 33793 16028
rect 33468 15988 33474 16000
rect 33781 15997 33793 16000
rect 33827 16028 33839 16031
rect 35084 16028 35112 16068
rect 35820 16037 35848 16068
rect 35986 16056 35992 16068
rect 36044 16056 36050 16108
rect 37274 16096 37280 16108
rect 37016 16068 37280 16096
rect 33827 16000 35112 16028
rect 35529 16031 35587 16037
rect 33827 15997 33839 16000
rect 33781 15991 33839 15997
rect 35529 15997 35541 16031
rect 35575 15997 35587 16031
rect 35529 15991 35587 15997
rect 35805 16031 35863 16037
rect 35805 15997 35817 16031
rect 35851 16028 35863 16031
rect 35894 16028 35900 16040
rect 35851 16000 35900 16028
rect 35851 15997 35863 16000
rect 35805 15991 35863 15997
rect 29236 15932 30144 15960
rect 29236 15920 29242 15932
rect 25792 15864 26556 15892
rect 26605 15895 26663 15901
rect 26605 15861 26617 15895
rect 26651 15892 26663 15895
rect 26786 15892 26792 15904
rect 26651 15864 26792 15892
rect 26651 15861 26663 15864
rect 26605 15855 26663 15861
rect 26786 15852 26792 15864
rect 26844 15852 26850 15904
rect 27246 15892 27252 15904
rect 27207 15864 27252 15892
rect 27246 15852 27252 15864
rect 27304 15852 27310 15904
rect 28629 15895 28687 15901
rect 28629 15861 28641 15895
rect 28675 15892 28687 15895
rect 29362 15892 29368 15904
rect 28675 15864 29368 15892
rect 28675 15861 28687 15864
rect 28629 15855 28687 15861
rect 29362 15852 29368 15864
rect 29420 15852 29426 15904
rect 35544 15892 35572 15991
rect 35894 15988 35900 16000
rect 35952 15988 35958 16040
rect 37016 16037 37044 16068
rect 37274 16056 37280 16068
rect 37332 16056 37338 16108
rect 36725 16031 36783 16037
rect 36725 15997 36737 16031
rect 36771 15997 36783 16031
rect 36725 15991 36783 15997
rect 37001 16031 37059 16037
rect 37001 15997 37013 16031
rect 37047 15997 37059 16031
rect 37182 16028 37188 16040
rect 37143 16000 37188 16028
rect 37001 15991 37059 15997
rect 36740 15960 36768 15991
rect 37182 15988 37188 16000
rect 37240 15988 37246 16040
rect 37366 15960 37372 15972
rect 36740 15932 37372 15960
rect 37366 15920 37372 15932
rect 37424 15920 37430 15972
rect 36998 15892 37004 15904
rect 35544 15864 37004 15892
rect 36998 15852 37004 15864
rect 37056 15852 37062 15904
rect 1104 15802 38824 15824
rect 1104 15750 19606 15802
rect 19658 15750 19670 15802
rect 19722 15750 19734 15802
rect 19786 15750 19798 15802
rect 19850 15750 38824 15802
rect 1104 15728 38824 15750
rect 2682 15688 2688 15700
rect 2643 15660 2688 15688
rect 2682 15648 2688 15660
rect 2740 15648 2746 15700
rect 4433 15691 4491 15697
rect 4433 15657 4445 15691
rect 4479 15688 4491 15691
rect 4522 15688 4528 15700
rect 4479 15660 4528 15688
rect 4479 15657 4491 15660
rect 4433 15651 4491 15657
rect 4522 15648 4528 15660
rect 4580 15648 4586 15700
rect 5537 15691 5595 15697
rect 5537 15657 5549 15691
rect 5583 15688 5595 15691
rect 5626 15688 5632 15700
rect 5583 15660 5632 15688
rect 5583 15657 5595 15660
rect 5537 15651 5595 15657
rect 5626 15648 5632 15660
rect 5684 15648 5690 15700
rect 7653 15691 7711 15697
rect 7653 15688 7665 15691
rect 6380 15660 7665 15688
rect 4062 15580 4068 15632
rect 4120 15620 4126 15632
rect 6380 15620 6408 15660
rect 7653 15657 7665 15660
rect 7699 15688 7711 15691
rect 9582 15688 9588 15700
rect 7699 15660 9588 15688
rect 7699 15657 7711 15660
rect 7653 15651 7711 15657
rect 9582 15648 9588 15660
rect 9640 15648 9646 15700
rect 10134 15648 10140 15700
rect 10192 15688 10198 15700
rect 11422 15688 11428 15700
rect 10192 15660 11428 15688
rect 10192 15648 10198 15660
rect 11422 15648 11428 15660
rect 11480 15688 11486 15700
rect 15933 15691 15991 15697
rect 11480 15660 13952 15688
rect 11480 15648 11486 15660
rect 4120 15592 6408 15620
rect 13924 15620 13952 15660
rect 15933 15657 15945 15691
rect 15979 15688 15991 15691
rect 16022 15688 16028 15700
rect 15979 15660 16028 15688
rect 15979 15657 15991 15660
rect 15933 15651 15991 15657
rect 16022 15648 16028 15660
rect 16080 15648 16086 15700
rect 16298 15648 16304 15700
rect 16356 15688 16362 15700
rect 19061 15691 19119 15697
rect 16356 15660 18368 15688
rect 16356 15648 16362 15660
rect 18340 15620 18368 15660
rect 19061 15657 19073 15691
rect 19107 15688 19119 15691
rect 19334 15688 19340 15700
rect 19107 15660 19340 15688
rect 19107 15657 19119 15660
rect 19061 15651 19119 15657
rect 19334 15648 19340 15660
rect 19392 15648 19398 15700
rect 22830 15688 22836 15700
rect 19904 15660 22836 15688
rect 19794 15620 19800 15632
rect 13924 15592 14320 15620
rect 4120 15580 4126 15592
rect 2869 15555 2927 15561
rect 2869 15521 2881 15555
rect 2915 15552 2927 15555
rect 2958 15552 2964 15564
rect 2915 15524 2964 15552
rect 2915 15521 2927 15524
rect 2869 15515 2927 15521
rect 2958 15512 2964 15524
rect 3016 15512 3022 15564
rect 3142 15552 3148 15564
rect 3103 15524 3148 15552
rect 3142 15512 3148 15524
rect 3200 15512 3206 15564
rect 4157 15555 4215 15561
rect 4157 15521 4169 15555
rect 4203 15521 4215 15555
rect 4706 15552 4712 15564
rect 4667 15524 4712 15552
rect 4157 15515 4215 15521
rect 1762 15444 1768 15496
rect 1820 15484 1826 15496
rect 4172 15484 4200 15515
rect 4706 15512 4712 15524
rect 4764 15512 4770 15564
rect 5353 15555 5411 15561
rect 5353 15521 5365 15555
rect 5399 15552 5411 15555
rect 5626 15552 5632 15564
rect 5399 15524 5632 15552
rect 5399 15521 5411 15524
rect 5353 15515 5411 15521
rect 5626 15512 5632 15524
rect 5684 15552 5690 15564
rect 7190 15552 7196 15564
rect 5684 15524 7196 15552
rect 5684 15512 5690 15524
rect 7190 15512 7196 15524
rect 7248 15512 7254 15564
rect 9490 15512 9496 15564
rect 9548 15552 9554 15564
rect 13924 15561 13952 15592
rect 11149 15555 11207 15561
rect 11149 15552 11161 15555
rect 9548 15524 11161 15552
rect 9548 15512 9554 15524
rect 11149 15521 11161 15524
rect 11195 15521 11207 15555
rect 11149 15515 11207 15521
rect 13633 15555 13691 15561
rect 13633 15521 13645 15555
rect 13679 15552 13691 15555
rect 13909 15555 13967 15561
rect 13679 15524 13860 15552
rect 13679 15521 13691 15524
rect 13633 15515 13691 15521
rect 5810 15484 5816 15496
rect 1820 15456 5816 15484
rect 1820 15444 1826 15456
rect 5810 15444 5816 15456
rect 5868 15444 5874 15496
rect 6270 15484 6276 15496
rect 6231 15456 6276 15484
rect 6270 15444 6276 15456
rect 6328 15444 6334 15496
rect 6549 15487 6607 15493
rect 6549 15453 6561 15487
rect 6595 15484 6607 15487
rect 9674 15484 9680 15496
rect 6595 15456 9680 15484
rect 6595 15453 6607 15456
rect 6549 15447 6607 15453
rect 9674 15444 9680 15456
rect 9732 15444 9738 15496
rect 11425 15487 11483 15493
rect 11425 15453 11437 15487
rect 11471 15484 11483 15487
rect 13262 15484 13268 15496
rect 11471 15456 13268 15484
rect 11471 15453 11483 15456
rect 11425 15447 11483 15453
rect 13262 15444 13268 15456
rect 13320 15444 13326 15496
rect 13832 15416 13860 15524
rect 13909 15521 13921 15555
rect 13955 15521 13967 15555
rect 14182 15552 14188 15564
rect 14143 15524 14188 15552
rect 13909 15515 13967 15521
rect 14182 15512 14188 15524
rect 14240 15512 14246 15564
rect 13998 15484 14004 15496
rect 13959 15456 14004 15484
rect 13998 15444 14004 15456
rect 14056 15444 14062 15496
rect 14292 15484 14320 15592
rect 15856 15592 18276 15620
rect 18340 15592 19800 15620
rect 15856 15561 15884 15592
rect 15841 15555 15899 15561
rect 15841 15521 15853 15555
rect 15887 15521 15899 15555
rect 15841 15515 15899 15521
rect 16669 15555 16727 15561
rect 16669 15521 16681 15555
rect 16715 15521 16727 15555
rect 16942 15552 16948 15564
rect 16903 15524 16948 15552
rect 16669 15515 16727 15521
rect 16482 15484 16488 15496
rect 14292 15456 16488 15484
rect 16482 15444 16488 15456
rect 16540 15444 16546 15496
rect 16684 15484 16712 15515
rect 16942 15512 16948 15524
rect 17000 15512 17006 15564
rect 17497 15555 17555 15561
rect 17497 15521 17509 15555
rect 17543 15521 17555 15555
rect 17862 15552 17868 15564
rect 17823 15524 17868 15552
rect 17497 15515 17555 15521
rect 17126 15484 17132 15496
rect 16684 15456 17132 15484
rect 17126 15444 17132 15456
rect 17184 15444 17190 15496
rect 17512 15484 17540 15515
rect 17862 15512 17868 15524
rect 17920 15512 17926 15564
rect 18138 15552 18144 15564
rect 18099 15524 18144 15552
rect 18138 15512 18144 15524
rect 18196 15512 18202 15564
rect 18248 15552 18276 15592
rect 19794 15580 19800 15592
rect 19852 15580 19858 15632
rect 18966 15552 18972 15564
rect 18248 15524 18972 15552
rect 18966 15512 18972 15524
rect 19024 15512 19030 15564
rect 19904 15561 19932 15660
rect 22830 15648 22836 15660
rect 22888 15648 22894 15700
rect 22922 15648 22928 15700
rect 22980 15688 22986 15700
rect 22980 15660 23612 15688
rect 22980 15648 22986 15660
rect 23584 15620 23612 15660
rect 27430 15648 27436 15700
rect 27488 15688 27494 15700
rect 29730 15688 29736 15700
rect 27488 15660 27660 15688
rect 29691 15660 29736 15688
rect 27488 15648 27494 15660
rect 20088 15592 21772 15620
rect 20088 15561 20116 15592
rect 19889 15555 19947 15561
rect 19889 15521 19901 15555
rect 19935 15521 19947 15555
rect 19889 15515 19947 15521
rect 20073 15555 20131 15561
rect 20073 15521 20085 15555
rect 20119 15521 20131 15555
rect 21174 15552 21180 15564
rect 21135 15524 21180 15552
rect 20073 15515 20131 15521
rect 21174 15512 21180 15524
rect 21232 15512 21238 15564
rect 21744 15561 21772 15592
rect 23584 15592 25820 15620
rect 21729 15555 21787 15561
rect 21729 15521 21741 15555
rect 21775 15552 21787 15555
rect 21910 15552 21916 15564
rect 21775 15524 21916 15552
rect 21775 15521 21787 15524
rect 21729 15515 21787 15521
rect 21910 15512 21916 15524
rect 21968 15512 21974 15564
rect 23198 15552 23204 15564
rect 23159 15524 23204 15552
rect 23198 15512 23204 15524
rect 23256 15512 23262 15564
rect 23584 15561 23612 15592
rect 25792 15564 25820 15592
rect 23569 15555 23627 15561
rect 23569 15521 23581 15555
rect 23615 15521 23627 15555
rect 23569 15515 23627 15521
rect 24121 15555 24179 15561
rect 24121 15521 24133 15555
rect 24167 15552 24179 15555
rect 24394 15552 24400 15564
rect 24167 15524 24400 15552
rect 24167 15521 24179 15524
rect 24121 15515 24179 15521
rect 24394 15512 24400 15524
rect 24452 15512 24458 15564
rect 25409 15555 25467 15561
rect 25409 15521 25421 15555
rect 25455 15552 25467 15555
rect 25498 15552 25504 15564
rect 25455 15524 25504 15552
rect 25455 15521 25467 15524
rect 25409 15515 25467 15521
rect 25498 15512 25504 15524
rect 25556 15512 25562 15564
rect 25774 15552 25780 15564
rect 25735 15524 25780 15552
rect 25774 15512 25780 15524
rect 25832 15512 25838 15564
rect 25869 15555 25927 15561
rect 25869 15521 25881 15555
rect 25915 15552 25927 15555
rect 26602 15552 26608 15564
rect 25915 15524 26608 15552
rect 25915 15521 25927 15524
rect 25869 15515 25927 15521
rect 26602 15512 26608 15524
rect 26660 15512 26666 15564
rect 27062 15552 27068 15564
rect 27023 15524 27068 15552
rect 27062 15512 27068 15524
rect 27120 15512 27126 15564
rect 27249 15555 27307 15561
rect 27249 15521 27261 15555
rect 27295 15521 27307 15555
rect 27249 15515 27307 15521
rect 27433 15555 27491 15561
rect 27433 15521 27445 15555
rect 27479 15552 27491 15555
rect 27522 15552 27528 15564
rect 27479 15524 27528 15552
rect 27479 15521 27491 15524
rect 27433 15515 27491 15521
rect 17954 15484 17960 15496
rect 17512 15456 17960 15484
rect 17954 15444 17960 15456
rect 18012 15444 18018 15496
rect 18322 15444 18328 15496
rect 18380 15484 18386 15496
rect 20165 15487 20223 15493
rect 20165 15484 20177 15487
rect 18380 15456 20177 15484
rect 18380 15444 18386 15456
rect 20165 15453 20177 15456
rect 20211 15453 20223 15487
rect 21818 15484 21824 15496
rect 20165 15447 20223 15453
rect 20456 15456 21680 15484
rect 21779 15456 21824 15484
rect 16298 15416 16304 15428
rect 13832 15388 16304 15416
rect 16298 15376 16304 15388
rect 16356 15376 16362 15428
rect 16574 15416 16580 15428
rect 16535 15388 16580 15416
rect 16574 15376 16580 15388
rect 16632 15376 16638 15428
rect 16758 15376 16764 15428
rect 16816 15416 16822 15428
rect 20456 15416 20484 15456
rect 21652 15425 21680 15456
rect 21818 15444 21824 15456
rect 21876 15444 21882 15496
rect 24946 15484 24952 15496
rect 24907 15456 24952 15484
rect 24946 15444 24952 15456
rect 25004 15444 25010 15496
rect 26786 15444 26792 15496
rect 26844 15484 26850 15496
rect 27264 15484 27292 15515
rect 27522 15512 27528 15524
rect 27580 15512 27586 15564
rect 27632 15561 27660 15660
rect 29730 15648 29736 15660
rect 29788 15648 29794 15700
rect 32217 15691 32275 15697
rect 32217 15657 32229 15691
rect 32263 15688 32275 15691
rect 32766 15688 32772 15700
rect 32263 15660 32772 15688
rect 32263 15657 32275 15660
rect 32217 15651 32275 15657
rect 32766 15648 32772 15660
rect 32824 15648 32830 15700
rect 35894 15648 35900 15700
rect 35952 15688 35958 15700
rect 35952 15660 37780 15688
rect 35952 15648 35958 15660
rect 28166 15620 28172 15632
rect 27724 15592 28172 15620
rect 27617 15555 27675 15561
rect 27617 15521 27629 15555
rect 27663 15521 27675 15555
rect 27617 15515 27675 15521
rect 27724 15484 27752 15592
rect 28166 15580 28172 15592
rect 28224 15580 28230 15632
rect 30926 15620 30932 15632
rect 30852 15592 30932 15620
rect 27801 15555 27859 15561
rect 27801 15521 27813 15555
rect 27847 15521 27859 15555
rect 28534 15552 28540 15564
rect 28495 15524 28540 15552
rect 27801 15515 27859 15521
rect 26844 15456 27752 15484
rect 26844 15444 26850 15456
rect 16816 15388 20484 15416
rect 21637 15419 21695 15425
rect 16816 15376 16822 15388
rect 21637 15385 21649 15419
rect 21683 15385 21695 15419
rect 21637 15379 21695 15385
rect 22002 15376 22008 15428
rect 22060 15416 22066 15428
rect 23017 15419 23075 15425
rect 23017 15416 23029 15419
rect 22060 15388 23029 15416
rect 22060 15376 22066 15388
rect 23017 15385 23029 15388
rect 23063 15385 23075 15419
rect 23017 15379 23075 15385
rect 26694 15376 26700 15428
rect 26752 15416 26758 15428
rect 27816 15416 27844 15515
rect 28534 15512 28540 15524
rect 28592 15512 28598 15564
rect 28994 15552 29000 15564
rect 28955 15524 29000 15552
rect 28994 15512 29000 15524
rect 29052 15512 29058 15564
rect 29362 15552 29368 15564
rect 29323 15524 29368 15552
rect 29362 15512 29368 15524
rect 29420 15512 29426 15564
rect 29454 15512 29460 15564
rect 29512 15552 29518 15564
rect 29733 15555 29791 15561
rect 29733 15552 29745 15555
rect 29512 15524 29745 15552
rect 29512 15512 29518 15524
rect 29733 15521 29745 15524
rect 29779 15521 29791 15555
rect 29733 15515 29791 15521
rect 30742 15512 30748 15564
rect 30800 15552 30806 15564
rect 30852 15561 30880 15592
rect 30926 15580 30932 15592
rect 30984 15580 30990 15632
rect 33410 15620 33416 15632
rect 32140 15592 33416 15620
rect 32140 15561 32168 15592
rect 33410 15580 33416 15592
rect 33468 15580 33474 15632
rect 33962 15580 33968 15632
rect 34020 15620 34026 15632
rect 36906 15620 36912 15632
rect 34020 15592 34744 15620
rect 36867 15592 36912 15620
rect 34020 15580 34026 15592
rect 30837 15555 30895 15561
rect 30837 15552 30849 15555
rect 30800 15524 30849 15552
rect 30800 15512 30806 15524
rect 30837 15521 30849 15524
rect 30883 15521 30895 15555
rect 31297 15555 31355 15561
rect 31297 15552 31309 15555
rect 30837 15515 30895 15521
rect 30944 15524 31309 15552
rect 30006 15444 30012 15496
rect 30064 15484 30070 15496
rect 30944 15484 30972 15524
rect 31297 15521 31309 15524
rect 31343 15521 31355 15555
rect 31297 15515 31355 15521
rect 32125 15555 32183 15561
rect 32125 15521 32137 15555
rect 32171 15521 32183 15555
rect 33042 15552 33048 15564
rect 33003 15524 33048 15552
rect 32125 15515 32183 15521
rect 33042 15512 33048 15524
rect 33100 15512 33106 15564
rect 33137 15555 33195 15561
rect 33137 15521 33149 15555
rect 33183 15521 33195 15555
rect 33137 15515 33195 15521
rect 33689 15555 33747 15561
rect 33689 15521 33701 15555
rect 33735 15521 33747 15555
rect 34054 15552 34060 15564
rect 34015 15524 34060 15552
rect 33689 15515 33747 15521
rect 31386 15484 31392 15496
rect 30064 15456 30972 15484
rect 31347 15456 31392 15484
rect 30064 15444 30070 15456
rect 31386 15444 31392 15456
rect 31444 15444 31450 15496
rect 32490 15444 32496 15496
rect 32548 15484 32554 15496
rect 33152 15484 33180 15515
rect 33318 15484 33324 15496
rect 32548 15456 33180 15484
rect 33279 15456 33324 15484
rect 32548 15444 32554 15456
rect 26752 15388 27844 15416
rect 33060 15416 33088 15456
rect 33318 15444 33324 15456
rect 33376 15444 33382 15496
rect 33704 15484 33732 15515
rect 34054 15512 34060 15524
rect 34112 15512 34118 15564
rect 34716 15561 34744 15592
rect 36906 15580 36912 15592
rect 36964 15580 36970 15632
rect 34701 15555 34759 15561
rect 34701 15521 34713 15555
rect 34747 15521 34759 15555
rect 35710 15552 35716 15564
rect 35671 15524 35716 15552
rect 34701 15515 34759 15521
rect 35710 15512 35716 15524
rect 35768 15512 35774 15564
rect 36357 15555 36415 15561
rect 36357 15521 36369 15555
rect 36403 15521 36415 15555
rect 36630 15552 36636 15564
rect 36591 15524 36636 15552
rect 36357 15515 36415 15521
rect 35342 15484 35348 15496
rect 33704 15456 35348 15484
rect 35342 15444 35348 15456
rect 35400 15444 35406 15496
rect 36372 15484 36400 15515
rect 36630 15512 36636 15524
rect 36688 15512 36694 15564
rect 37185 15555 37243 15561
rect 37185 15521 37197 15555
rect 37231 15552 37243 15555
rect 37274 15552 37280 15564
rect 37231 15524 37280 15552
rect 37231 15521 37243 15524
rect 37185 15515 37243 15521
rect 37274 15512 37280 15524
rect 37332 15512 37338 15564
rect 37752 15561 37780 15660
rect 37737 15555 37795 15561
rect 37737 15521 37749 15555
rect 37783 15521 37795 15555
rect 37737 15515 37795 15521
rect 37366 15484 37372 15496
rect 36372 15456 37372 15484
rect 37366 15444 37372 15456
rect 37424 15444 37430 15496
rect 34885 15419 34943 15425
rect 34885 15416 34897 15419
rect 33060 15388 34897 15416
rect 26752 15376 26758 15388
rect 34885 15385 34897 15388
rect 34931 15385 34943 15419
rect 34885 15379 34943 15385
rect 3786 15308 3792 15360
rect 3844 15348 3850 15360
rect 11330 15348 11336 15360
rect 3844 15320 11336 15348
rect 3844 15308 3850 15320
rect 11330 15308 11336 15320
rect 11388 15348 11394 15360
rect 12526 15348 12532 15360
rect 11388 15320 12532 15348
rect 11388 15308 11394 15320
rect 12526 15308 12532 15320
rect 12584 15308 12590 15360
rect 23750 15308 23756 15360
rect 23808 15348 23814 15360
rect 24305 15351 24363 15357
rect 24305 15348 24317 15351
rect 23808 15320 24317 15348
rect 23808 15308 23814 15320
rect 24305 15317 24317 15320
rect 24351 15317 24363 15351
rect 26602 15348 26608 15360
rect 26563 15320 26608 15348
rect 24305 15311 24363 15317
rect 26602 15308 26608 15320
rect 26660 15308 26666 15360
rect 35434 15308 35440 15360
rect 35492 15348 35498 15360
rect 37921 15351 37979 15357
rect 37921 15348 37933 15351
rect 35492 15320 37933 15348
rect 35492 15308 35498 15320
rect 37921 15317 37933 15320
rect 37967 15317 37979 15351
rect 37921 15311 37979 15317
rect 1104 15258 38824 15280
rect 1104 15206 4246 15258
rect 4298 15206 4310 15258
rect 4362 15206 4374 15258
rect 4426 15206 4438 15258
rect 4490 15206 34966 15258
rect 35018 15206 35030 15258
rect 35082 15206 35094 15258
rect 35146 15206 35158 15258
rect 35210 15206 38824 15258
rect 1104 15184 38824 15206
rect 1670 15104 1676 15156
rect 1728 15144 1734 15156
rect 2409 15147 2467 15153
rect 2409 15144 2421 15147
rect 1728 15116 2421 15144
rect 1728 15104 1734 15116
rect 2409 15113 2421 15116
rect 2455 15113 2467 15147
rect 2409 15107 2467 15113
rect 3896 15116 5304 15144
rect 1854 15036 1860 15088
rect 1912 15076 1918 15088
rect 3896 15076 3924 15116
rect 1912 15048 3924 15076
rect 5276 15076 5304 15116
rect 5350 15104 5356 15156
rect 5408 15144 5414 15156
rect 6181 15147 6239 15153
rect 6181 15144 6193 15147
rect 5408 15116 6193 15144
rect 5408 15104 5414 15116
rect 6181 15113 6193 15116
rect 6227 15144 6239 15147
rect 14458 15144 14464 15156
rect 6227 15116 14464 15144
rect 6227 15113 6239 15116
rect 6181 15107 6239 15113
rect 14458 15104 14464 15116
rect 14516 15104 14522 15156
rect 16758 15144 16764 15156
rect 15396 15116 16764 15144
rect 5994 15076 6000 15088
rect 5276 15048 6000 15076
rect 1912 15036 1918 15048
rect 3896 15017 3924 15048
rect 5994 15036 6000 15048
rect 6052 15076 6058 15088
rect 6270 15076 6276 15088
rect 6052 15048 6276 15076
rect 6052 15036 6058 15048
rect 6270 15036 6276 15048
rect 6328 15036 6334 15088
rect 10226 15036 10232 15088
rect 10284 15076 10290 15088
rect 11793 15079 11851 15085
rect 11793 15076 11805 15079
rect 10284 15048 11805 15076
rect 10284 15036 10290 15048
rect 11793 15045 11805 15048
rect 11839 15045 11851 15079
rect 11793 15039 11851 15045
rect 3881 15011 3939 15017
rect 3881 14977 3893 15011
rect 3927 14977 3939 15011
rect 4614 15008 4620 15020
rect 3881 14971 3939 14977
rect 3988 14980 4620 15008
rect 2130 14940 2136 14952
rect 2091 14912 2136 14940
rect 2130 14900 2136 14912
rect 2188 14900 2194 14952
rect 2225 14943 2283 14949
rect 2225 14909 2237 14943
rect 2271 14940 2283 14943
rect 2774 14940 2780 14952
rect 2271 14912 2780 14940
rect 2271 14909 2283 14912
rect 2225 14903 2283 14909
rect 2774 14900 2780 14912
rect 2832 14900 2838 14952
rect 3237 14943 3295 14949
rect 3237 14909 3249 14943
rect 3283 14909 3295 14943
rect 3237 14903 3295 14909
rect 3252 14804 3280 14903
rect 3329 14875 3387 14881
rect 3329 14841 3341 14875
rect 3375 14872 3387 14875
rect 3988 14872 4016 14980
rect 4614 14968 4620 14980
rect 4672 14968 4678 15020
rect 5445 15011 5503 15017
rect 5445 14977 5457 15011
rect 5491 15008 5503 15011
rect 7374 15008 7380 15020
rect 5491 14980 7380 15008
rect 5491 14977 5503 14980
rect 5445 14971 5503 14977
rect 4154 14940 4160 14952
rect 4115 14912 4160 14940
rect 4154 14900 4160 14912
rect 4212 14900 4218 14952
rect 3375 14844 4016 14872
rect 3375 14841 3387 14844
rect 3329 14835 3387 14841
rect 5460 14804 5488 14971
rect 7374 14968 7380 14980
rect 7432 14968 7438 15020
rect 7558 15008 7564 15020
rect 7471 14980 7564 15008
rect 5626 14900 5632 14952
rect 5684 14940 5690 14952
rect 5997 14943 6055 14949
rect 5997 14940 6009 14943
rect 5684 14912 6009 14940
rect 5684 14900 5690 14912
rect 5997 14909 6009 14912
rect 6043 14909 6055 14943
rect 5997 14903 6055 14909
rect 6178 14900 6184 14952
rect 6236 14940 6242 14952
rect 6822 14940 6828 14952
rect 6236 14912 6828 14940
rect 6236 14900 6242 14912
rect 6822 14900 6828 14912
rect 6880 14900 6886 14952
rect 7098 14900 7104 14952
rect 7156 14940 7162 14952
rect 7484 14940 7512 14980
rect 7558 14968 7564 14980
rect 7616 15008 7622 15020
rect 10502 15008 10508 15020
rect 7616 14980 10364 15008
rect 10463 14980 10508 15008
rect 7616 14968 7622 14980
rect 7156 14912 7512 14940
rect 7745 14943 7803 14949
rect 7156 14900 7162 14912
rect 7745 14909 7757 14943
rect 7791 14909 7803 14943
rect 8018 14940 8024 14952
rect 7979 14912 8024 14940
rect 7745 14903 7803 14909
rect 6270 14832 6276 14884
rect 6328 14872 6334 14884
rect 7760 14872 7788 14903
rect 8018 14900 8024 14912
rect 8076 14900 8082 14952
rect 9030 14900 9036 14952
rect 9088 14940 9094 14952
rect 9582 14940 9588 14952
rect 9088 14912 9588 14940
rect 9088 14900 9094 14912
rect 9582 14900 9588 14912
rect 9640 14940 9646 14952
rect 9861 14943 9919 14949
rect 9861 14940 9873 14943
rect 9640 14912 9873 14940
rect 9640 14900 9646 14912
rect 9861 14909 9873 14912
rect 9907 14909 9919 14943
rect 9861 14903 9919 14909
rect 10134 14900 10140 14952
rect 10192 14940 10198 14952
rect 10229 14943 10287 14949
rect 10229 14940 10241 14943
rect 10192 14912 10241 14940
rect 10192 14900 10198 14912
rect 10229 14909 10241 14912
rect 10275 14909 10287 14943
rect 10336 14940 10364 14980
rect 10502 14968 10508 14980
rect 10560 14968 10566 15020
rect 11808 15008 11836 15039
rect 12434 15036 12440 15088
rect 12492 15076 12498 15088
rect 13262 15076 13268 15088
rect 12492 15048 12940 15076
rect 13223 15048 13268 15076
rect 12492 15036 12498 15048
rect 12912 15008 12940 15048
rect 13262 15036 13268 15048
rect 13320 15036 13326 15088
rect 15286 15008 15292 15020
rect 10612 14980 11284 15008
rect 11808 14980 12848 15008
rect 12912 14980 14044 15008
rect 15247 14980 15292 15008
rect 10612 14940 10640 14980
rect 10870 14940 10876 14952
rect 10336 14912 10640 14940
rect 10831 14912 10876 14940
rect 10229 14903 10287 14909
rect 10870 14900 10876 14912
rect 10928 14900 10934 14952
rect 6328 14844 7788 14872
rect 6328 14832 6334 14844
rect 7006 14804 7012 14816
rect 3252 14776 5488 14804
rect 6967 14776 7012 14804
rect 7006 14764 7012 14776
rect 7064 14764 7070 14816
rect 7760 14804 7788 14844
rect 9401 14875 9459 14881
rect 9401 14841 9413 14875
rect 9447 14872 9459 14875
rect 9766 14872 9772 14884
rect 9447 14844 9772 14872
rect 9447 14841 9459 14844
rect 9401 14835 9459 14841
rect 9766 14832 9772 14844
rect 9824 14832 9830 14884
rect 9490 14804 9496 14816
rect 7760 14776 9496 14804
rect 9490 14764 9496 14776
rect 9548 14764 9554 14816
rect 9582 14764 9588 14816
rect 9640 14804 9646 14816
rect 10152 14804 10180 14900
rect 9640 14776 10180 14804
rect 11256 14804 11284 14980
rect 12820 14952 12848 14980
rect 11609 14943 11667 14949
rect 11609 14909 11621 14943
rect 11655 14940 11667 14943
rect 12434 14940 12440 14952
rect 11655 14912 12440 14940
rect 11655 14909 11667 14912
rect 11609 14903 11667 14909
rect 12434 14900 12440 14912
rect 12492 14900 12498 14952
rect 12529 14943 12587 14949
rect 12529 14909 12541 14943
rect 12575 14909 12587 14943
rect 12802 14940 12808 14952
rect 12763 14912 12808 14940
rect 12529 14903 12587 14909
rect 12250 14832 12256 14884
rect 12308 14872 12314 14884
rect 12544 14872 12572 14903
rect 12802 14900 12808 14912
rect 12860 14900 12866 14952
rect 13262 14940 13268 14952
rect 13223 14912 13268 14940
rect 13262 14900 13268 14912
rect 13320 14900 13326 14952
rect 14016 14949 14044 14980
rect 15286 14968 15292 14980
rect 15344 14968 15350 15020
rect 14001 14943 14059 14949
rect 14001 14909 14013 14943
rect 14047 14909 14059 14943
rect 14001 14903 14059 14909
rect 15197 14943 15255 14949
rect 15197 14909 15209 14943
rect 15243 14940 15255 14943
rect 15396 14940 15424 15116
rect 16758 15104 16764 15116
rect 16816 15104 16822 15156
rect 17034 15104 17040 15156
rect 17092 15144 17098 15156
rect 18141 15147 18199 15153
rect 18141 15144 18153 15147
rect 17092 15116 18153 15144
rect 17092 15104 17098 15116
rect 18141 15113 18153 15116
rect 18187 15113 18199 15147
rect 18141 15107 18199 15113
rect 20533 15147 20591 15153
rect 20533 15113 20545 15147
rect 20579 15144 20591 15147
rect 23198 15144 23204 15156
rect 20579 15116 23204 15144
rect 20579 15113 20591 15116
rect 20533 15107 20591 15113
rect 23198 15104 23204 15116
rect 23256 15104 23262 15156
rect 28350 15104 28356 15156
rect 28408 15144 28414 15156
rect 34238 15144 34244 15156
rect 28408 15116 34244 15144
rect 28408 15104 28414 15116
rect 34238 15104 34244 15116
rect 34296 15104 34302 15156
rect 37366 15104 37372 15156
rect 37424 15144 37430 15156
rect 37829 15147 37887 15153
rect 37829 15144 37841 15147
rect 37424 15116 37841 15144
rect 37424 15104 37430 15116
rect 37829 15113 37841 15116
rect 37875 15113 37887 15147
rect 37829 15107 37887 15113
rect 16942 15036 16948 15088
rect 17000 15076 17006 15088
rect 20898 15076 20904 15088
rect 17000 15048 20904 15076
rect 17000 15036 17006 15048
rect 20898 15036 20904 15048
rect 20956 15076 20962 15088
rect 21266 15076 21272 15088
rect 20956 15048 21272 15076
rect 20956 15036 20962 15048
rect 21266 15036 21272 15048
rect 21324 15036 21330 15088
rect 21818 15036 21824 15088
rect 21876 15076 21882 15088
rect 28626 15076 28632 15088
rect 21876 15048 23704 15076
rect 21876 15036 21882 15048
rect 16117 15011 16175 15017
rect 16117 14977 16129 15011
rect 16163 15008 16175 15011
rect 16574 15008 16580 15020
rect 16163 14980 16580 15008
rect 16163 14977 16175 14980
rect 16117 14971 16175 14977
rect 16574 14968 16580 14980
rect 16632 14968 16638 15020
rect 16758 14968 16764 15020
rect 16816 15008 16822 15020
rect 16816 14980 18736 15008
rect 16816 14968 16822 14980
rect 18708 14949 18736 14980
rect 19058 14968 19064 15020
rect 19116 15008 19122 15020
rect 19245 15011 19303 15017
rect 19245 15008 19257 15011
rect 19116 14980 19257 15008
rect 19116 14968 19122 14980
rect 19245 14977 19257 14980
rect 19291 14977 19303 15011
rect 21634 15008 21640 15020
rect 19245 14971 19303 14977
rect 21560 14980 21640 15008
rect 15243 14912 15424 14940
rect 15841 14943 15899 14949
rect 15243 14909 15255 14912
rect 15197 14903 15255 14909
rect 15841 14909 15853 14943
rect 15887 14909 15899 14943
rect 15841 14903 15899 14909
rect 18049 14943 18107 14949
rect 18049 14909 18061 14943
rect 18095 14909 18107 14943
rect 18049 14903 18107 14909
rect 18693 14943 18751 14949
rect 18693 14909 18705 14943
rect 18739 14909 18751 14943
rect 18693 14903 18751 14909
rect 19153 14943 19211 14949
rect 19153 14909 19165 14943
rect 19199 14909 19211 14943
rect 20346 14940 20352 14952
rect 20307 14912 20352 14940
rect 19153 14903 19211 14909
rect 14274 14872 14280 14884
rect 12308 14844 12572 14872
rect 14016 14844 14280 14872
rect 12308 14832 12314 14844
rect 14016 14804 14044 14844
rect 14274 14832 14280 14844
rect 14332 14832 14338 14884
rect 15102 14832 15108 14884
rect 15160 14872 15166 14884
rect 15856 14872 15884 14903
rect 15160 14844 15884 14872
rect 17497 14875 17555 14881
rect 15160 14832 15166 14844
rect 17497 14841 17509 14875
rect 17543 14872 17555 14875
rect 17586 14872 17592 14884
rect 17543 14844 17592 14872
rect 17543 14841 17555 14844
rect 17497 14835 17555 14841
rect 17586 14832 17592 14844
rect 17644 14872 17650 14884
rect 18064 14872 18092 14903
rect 17644 14844 18092 14872
rect 17644 14832 17650 14844
rect 14182 14804 14188 14816
rect 11256 14776 14044 14804
rect 14143 14776 14188 14804
rect 9640 14764 9646 14776
rect 14182 14764 14188 14776
rect 14240 14764 14246 14816
rect 14458 14764 14464 14816
rect 14516 14804 14522 14816
rect 18414 14804 18420 14816
rect 14516 14776 18420 14804
rect 14516 14764 14522 14776
rect 18414 14764 18420 14776
rect 18472 14764 18478 14816
rect 18708 14804 18736 14903
rect 19058 14832 19064 14884
rect 19116 14872 19122 14884
rect 19168 14872 19196 14903
rect 20346 14900 20352 14912
rect 20404 14900 20410 14952
rect 21560 14949 21588 14980
rect 21634 14968 21640 14980
rect 21692 15008 21698 15020
rect 21910 15008 21916 15020
rect 21692 14980 21916 15008
rect 21692 14968 21698 14980
rect 21910 14968 21916 14980
rect 21968 14968 21974 15020
rect 21545 14943 21603 14949
rect 21545 14909 21557 14943
rect 21591 14909 21603 14943
rect 21726 14940 21732 14952
rect 21687 14912 21732 14940
rect 21545 14903 21603 14909
rect 21726 14900 21732 14912
rect 21784 14900 21790 14952
rect 22005 14943 22063 14949
rect 22005 14909 22017 14943
rect 22051 14909 22063 14943
rect 22005 14903 22063 14909
rect 19116 14844 19196 14872
rect 19116 14832 19122 14844
rect 19242 14832 19248 14884
rect 19300 14872 19306 14884
rect 21085 14875 21143 14881
rect 21085 14872 21097 14875
rect 19300 14844 21097 14872
rect 19300 14832 19306 14844
rect 21085 14841 21097 14844
rect 21131 14841 21143 14875
rect 22020 14872 22048 14903
rect 22094 14900 22100 14952
rect 22152 14940 22158 14952
rect 22462 14940 22468 14952
rect 22152 14912 22197 14940
rect 22423 14912 22468 14940
rect 22152 14900 22158 14912
rect 22462 14900 22468 14912
rect 22520 14940 22526 14952
rect 23290 14940 23296 14952
rect 22520 14912 23296 14940
rect 22520 14900 22526 14912
rect 23290 14900 23296 14912
rect 23348 14900 23354 14952
rect 23676 14949 23704 15048
rect 24504 15048 28632 15076
rect 23661 14943 23719 14949
rect 23661 14909 23673 14943
rect 23707 14940 23719 14943
rect 23750 14940 23756 14952
rect 23707 14912 23756 14940
rect 23707 14909 23719 14912
rect 23661 14903 23719 14909
rect 23750 14900 23756 14912
rect 23808 14900 23814 14952
rect 24394 14900 24400 14952
rect 24452 14940 24458 14952
rect 24504 14949 24532 15048
rect 28626 15036 28632 15048
rect 28684 15036 28690 15088
rect 29178 15036 29184 15088
rect 29236 15076 29242 15088
rect 29733 15079 29791 15085
rect 29733 15076 29745 15079
rect 29236 15048 29745 15076
rect 29236 15036 29242 15048
rect 29733 15045 29745 15048
rect 29779 15076 29791 15079
rect 29914 15076 29920 15088
rect 29779 15048 29920 15076
rect 29779 15045 29791 15048
rect 29733 15039 29791 15045
rect 29914 15036 29920 15048
rect 29972 15036 29978 15088
rect 33962 15076 33968 15088
rect 33612 15048 33968 15076
rect 25958 15008 25964 15020
rect 25919 14980 25964 15008
rect 25958 14968 25964 14980
rect 26016 14968 26022 15020
rect 27338 14968 27344 15020
rect 27396 15008 27402 15020
rect 27396 14980 27844 15008
rect 27396 14968 27402 14980
rect 24489 14943 24547 14949
rect 24489 14940 24501 14943
rect 24452 14912 24501 14940
rect 24452 14900 24458 14912
rect 24489 14909 24501 14912
rect 24535 14909 24547 14943
rect 24489 14903 24547 14909
rect 25317 14943 25375 14949
rect 25317 14909 25329 14943
rect 25363 14909 25375 14943
rect 25682 14940 25688 14952
rect 25643 14912 25688 14940
rect 25317 14903 25375 14909
rect 22186 14872 22192 14884
rect 22020 14844 22192 14872
rect 21085 14835 21143 14841
rect 22186 14832 22192 14844
rect 22244 14832 22250 14884
rect 24581 14875 24639 14881
rect 24581 14872 24593 14875
rect 23676 14844 24593 14872
rect 19426 14804 19432 14816
rect 18708 14776 19432 14804
rect 19426 14764 19432 14776
rect 19484 14764 19490 14816
rect 22002 14764 22008 14816
rect 22060 14804 22066 14816
rect 23676 14804 23704 14844
rect 24581 14841 24593 14844
rect 24627 14841 24639 14875
rect 25332 14872 25360 14903
rect 25682 14900 25688 14912
rect 25740 14900 25746 14952
rect 26053 14943 26111 14949
rect 26053 14909 26065 14943
rect 26099 14940 26111 14943
rect 26602 14940 26608 14952
rect 26099 14912 26608 14940
rect 26099 14909 26111 14912
rect 26053 14903 26111 14909
rect 26602 14900 26608 14912
rect 26660 14900 26666 14952
rect 26694 14900 26700 14952
rect 26752 14940 26758 14952
rect 26973 14943 27031 14949
rect 26973 14940 26985 14943
rect 26752 14912 26985 14940
rect 26752 14900 26758 14912
rect 26973 14909 26985 14912
rect 27019 14909 27031 14943
rect 27430 14940 27436 14952
rect 27391 14912 27436 14940
rect 26973 14903 27031 14909
rect 27430 14900 27436 14912
rect 27488 14900 27494 14952
rect 27816 14949 27844 14980
rect 30098 14968 30104 15020
rect 30156 15008 30162 15020
rect 30285 15011 30343 15017
rect 30285 15008 30297 15011
rect 30156 14980 30297 15008
rect 30156 14968 30162 14980
rect 30285 14977 30297 14980
rect 30331 14977 30343 15011
rect 30285 14971 30343 14977
rect 27801 14943 27859 14949
rect 27801 14909 27813 14943
rect 27847 14909 27859 14943
rect 28166 14940 28172 14952
rect 28127 14912 28172 14940
rect 27801 14903 27859 14909
rect 28166 14900 28172 14912
rect 28224 14900 28230 14952
rect 29362 14900 29368 14952
rect 29420 14940 29426 14952
rect 29549 14943 29607 14949
rect 29549 14940 29561 14943
rect 29420 14912 29561 14940
rect 29420 14900 29426 14912
rect 29549 14909 29561 14912
rect 29595 14940 29607 14943
rect 30190 14940 30196 14952
rect 29595 14912 30196 14940
rect 29595 14909 29607 14912
rect 29549 14903 29607 14909
rect 30190 14900 30196 14912
rect 30248 14900 30254 14952
rect 30558 14940 30564 14952
rect 30519 14912 30564 14940
rect 30558 14900 30564 14912
rect 30616 14900 30622 14952
rect 33042 14900 33048 14952
rect 33100 14940 33106 14952
rect 33137 14943 33195 14949
rect 33137 14940 33149 14943
rect 33100 14912 33149 14940
rect 33100 14900 33106 14912
rect 33137 14909 33149 14912
rect 33183 14909 33195 14943
rect 33137 14903 33195 14909
rect 33505 14943 33563 14949
rect 33505 14909 33517 14943
rect 33551 14940 33563 14943
rect 33612 14940 33640 15048
rect 33962 15036 33968 15048
rect 34020 15036 34026 15088
rect 35526 15036 35532 15088
rect 35584 15076 35590 15088
rect 35713 15079 35771 15085
rect 35713 15076 35725 15079
rect 35584 15048 35725 15076
rect 35584 15036 35590 15048
rect 35713 15045 35725 15048
rect 35759 15045 35771 15079
rect 35713 15039 35771 15045
rect 33870 15008 33876 15020
rect 33831 14980 33876 15008
rect 33870 14968 33876 14980
rect 33928 14968 33934 15020
rect 34514 14968 34520 15020
rect 34572 15008 34578 15020
rect 35069 15011 35127 15017
rect 35069 15008 35081 15011
rect 34572 14980 35081 15008
rect 34572 14968 34578 14980
rect 35069 14977 35081 14980
rect 35115 15008 35127 15011
rect 35250 15008 35256 15020
rect 35115 14980 35256 15008
rect 35115 14977 35127 14980
rect 35069 14971 35127 14977
rect 35250 14968 35256 14980
rect 35308 14968 35314 15020
rect 35986 14968 35992 15020
rect 36044 15008 36050 15020
rect 36725 15011 36783 15017
rect 36725 15008 36737 15011
rect 36044 14980 36737 15008
rect 36044 14968 36050 14980
rect 36725 14977 36737 14980
rect 36771 14977 36783 15011
rect 36725 14971 36783 14977
rect 33551 14912 33640 14940
rect 33781 14943 33839 14949
rect 33551 14909 33563 14912
rect 33505 14903 33563 14909
rect 33781 14909 33793 14943
rect 33827 14940 33839 14943
rect 33962 14940 33968 14952
rect 33827 14912 33968 14940
rect 33827 14909 33839 14912
rect 33781 14903 33839 14909
rect 26510 14872 26516 14884
rect 25332 14844 26516 14872
rect 24581 14835 24639 14841
rect 23842 14804 23848 14816
rect 22060 14776 23704 14804
rect 23803 14776 23848 14804
rect 22060 14764 22066 14776
rect 23842 14764 23848 14776
rect 23900 14764 23906 14816
rect 24596 14804 24624 14835
rect 26510 14832 26516 14844
rect 26568 14872 26574 14884
rect 27890 14872 27896 14884
rect 26568 14844 27896 14872
rect 26568 14832 26574 14844
rect 27890 14832 27896 14844
rect 27948 14832 27954 14884
rect 33152 14872 33180 14903
rect 33962 14900 33968 14912
rect 34020 14900 34026 14952
rect 34146 14940 34152 14952
rect 34107 14912 34152 14940
rect 34146 14900 34152 14912
rect 34204 14900 34210 14952
rect 35434 14940 35440 14952
rect 35395 14912 35440 14940
rect 35434 14900 35440 14912
rect 35492 14900 35498 14952
rect 35526 14900 35532 14952
rect 35584 14940 35590 14952
rect 35713 14943 35771 14949
rect 35713 14940 35725 14943
rect 35584 14912 35725 14940
rect 35584 14900 35590 14912
rect 35713 14909 35725 14912
rect 35759 14909 35771 14943
rect 35713 14903 35771 14909
rect 36262 14900 36268 14952
rect 36320 14940 36326 14952
rect 36446 14940 36452 14952
rect 36320 14912 36452 14940
rect 36320 14900 36326 14912
rect 36446 14900 36452 14912
rect 36504 14900 36510 14952
rect 34514 14872 34520 14884
rect 33152 14844 34520 14872
rect 34514 14832 34520 14844
rect 34572 14832 34578 14884
rect 27522 14804 27528 14816
rect 24596 14776 27528 14804
rect 27522 14764 27528 14776
rect 27580 14764 27586 14816
rect 27614 14764 27620 14816
rect 27672 14804 27678 14816
rect 28169 14807 28227 14813
rect 28169 14804 28181 14807
rect 27672 14776 28181 14804
rect 27672 14764 27678 14776
rect 28169 14773 28181 14776
rect 28215 14773 28227 14807
rect 28169 14767 28227 14773
rect 30650 14764 30656 14816
rect 30708 14804 30714 14816
rect 31665 14807 31723 14813
rect 31665 14804 31677 14807
rect 30708 14776 31677 14804
rect 30708 14764 30714 14776
rect 31665 14773 31677 14776
rect 31711 14773 31723 14807
rect 31665 14767 31723 14773
rect 1104 14714 38824 14736
rect 1104 14662 19606 14714
rect 19658 14662 19670 14714
rect 19722 14662 19734 14714
rect 19786 14662 19798 14714
rect 19850 14662 38824 14714
rect 1104 14640 38824 14662
rect 2774 14560 2780 14612
rect 2832 14600 2838 14612
rect 19242 14600 19248 14612
rect 2832 14572 2877 14600
rect 4632 14572 19248 14600
rect 2832 14560 2838 14572
rect 3881 14467 3939 14473
rect 3881 14433 3893 14467
rect 3927 14433 3939 14467
rect 3881 14427 3939 14433
rect 1394 14396 1400 14408
rect 1355 14368 1400 14396
rect 1394 14356 1400 14368
rect 1452 14356 1458 14408
rect 1670 14396 1676 14408
rect 1631 14368 1676 14396
rect 1670 14356 1676 14368
rect 1728 14356 1734 14408
rect 3896 14328 3924 14427
rect 3970 14424 3976 14476
rect 4028 14464 4034 14476
rect 4525 14467 4583 14473
rect 4525 14464 4537 14467
rect 4028 14436 4537 14464
rect 4028 14424 4034 14436
rect 4525 14433 4537 14436
rect 4571 14464 4583 14467
rect 4632 14464 4660 14572
rect 19242 14560 19248 14572
rect 19300 14560 19306 14612
rect 22186 14600 22192 14612
rect 19352 14572 20944 14600
rect 19352 14544 19380 14572
rect 7006 14532 7012 14544
rect 5368 14504 7012 14532
rect 4571 14436 4660 14464
rect 4571 14433 4583 14436
rect 4525 14427 4583 14433
rect 4706 14424 4712 14476
rect 4764 14464 4770 14476
rect 4801 14467 4859 14473
rect 4801 14464 4813 14467
rect 4764 14436 4813 14464
rect 4764 14424 4770 14436
rect 4801 14433 4813 14436
rect 4847 14433 4859 14467
rect 4801 14427 4859 14433
rect 4982 14424 4988 14476
rect 5040 14464 5046 14476
rect 5368 14473 5396 14504
rect 7006 14492 7012 14504
rect 7064 14492 7070 14544
rect 8588 14504 10272 14532
rect 5353 14467 5411 14473
rect 5353 14464 5365 14467
rect 5040 14436 5365 14464
rect 5040 14424 5046 14436
rect 5353 14433 5365 14436
rect 5399 14433 5411 14467
rect 5353 14427 5411 14433
rect 5721 14467 5779 14473
rect 5721 14433 5733 14467
rect 5767 14433 5779 14467
rect 5721 14427 5779 14433
rect 6273 14467 6331 14473
rect 6273 14433 6285 14467
rect 6319 14464 6331 14467
rect 6914 14464 6920 14476
rect 6319 14436 6920 14464
rect 6319 14433 6331 14436
rect 6273 14427 6331 14433
rect 4154 14356 4160 14408
rect 4212 14396 4218 14408
rect 4433 14399 4491 14405
rect 4433 14396 4445 14399
rect 4212 14368 4445 14396
rect 4212 14356 4218 14368
rect 4433 14365 4445 14368
rect 4479 14365 4491 14399
rect 4433 14359 4491 14365
rect 5442 14356 5448 14408
rect 5500 14396 5506 14408
rect 5736 14396 5764 14427
rect 6914 14424 6920 14436
rect 6972 14424 6978 14476
rect 8588 14473 8616 14504
rect 10244 14476 10272 14504
rect 10870 14492 10876 14544
rect 10928 14532 10934 14544
rect 12437 14535 12495 14541
rect 10928 14504 12020 14532
rect 10928 14492 10934 14504
rect 7285 14467 7343 14473
rect 7285 14433 7297 14467
rect 7331 14433 7343 14467
rect 7285 14427 7343 14433
rect 8573 14467 8631 14473
rect 8573 14433 8585 14467
rect 8619 14433 8631 14467
rect 8938 14464 8944 14476
rect 8899 14436 8944 14464
rect 8573 14427 8631 14433
rect 7098 14396 7104 14408
rect 5500 14368 7104 14396
rect 5500 14356 5506 14368
rect 7098 14356 7104 14368
rect 7156 14356 7162 14408
rect 5074 14328 5080 14340
rect 3896 14300 5080 14328
rect 5074 14288 5080 14300
rect 5132 14288 5138 14340
rect 7300 14328 7328 14427
rect 8938 14424 8944 14436
rect 8996 14424 9002 14476
rect 9125 14467 9183 14473
rect 9125 14433 9137 14467
rect 9171 14464 9183 14467
rect 9950 14464 9956 14476
rect 9171 14436 9956 14464
rect 9171 14433 9183 14436
rect 9125 14427 9183 14433
rect 9950 14424 9956 14436
rect 10008 14424 10014 14476
rect 10226 14464 10232 14476
rect 10187 14436 10232 14464
rect 10226 14424 10232 14436
rect 10284 14424 10290 14476
rect 10502 14464 10508 14476
rect 10463 14436 10508 14464
rect 10502 14424 10508 14436
rect 10560 14424 10566 14476
rect 11330 14464 11336 14476
rect 11291 14436 11336 14464
rect 11330 14424 11336 14436
rect 11388 14424 11394 14476
rect 11882 14464 11888 14476
rect 11843 14436 11888 14464
rect 11882 14424 11888 14436
rect 11940 14424 11946 14476
rect 11992 14473 12020 14504
rect 12437 14501 12449 14535
rect 12483 14532 12495 14535
rect 13262 14532 13268 14544
rect 12483 14504 13268 14532
rect 12483 14501 12495 14504
rect 12437 14495 12495 14501
rect 13262 14492 13268 14504
rect 13320 14492 13326 14544
rect 14182 14532 14188 14544
rect 13372 14504 14188 14532
rect 11977 14467 12035 14473
rect 11977 14433 11989 14467
rect 12023 14464 12035 14467
rect 13372 14464 13400 14504
rect 14182 14492 14188 14504
rect 14240 14492 14246 14544
rect 18322 14532 18328 14544
rect 16868 14504 18328 14532
rect 12023 14436 13400 14464
rect 13449 14467 13507 14473
rect 12023 14433 12035 14436
rect 11977 14427 12035 14433
rect 13449 14433 13461 14467
rect 13495 14433 13507 14467
rect 13998 14464 14004 14476
rect 13959 14436 14004 14464
rect 13449 14427 13507 14433
rect 8205 14399 8263 14405
rect 8205 14365 8217 14399
rect 8251 14396 8263 14399
rect 8754 14396 8760 14408
rect 8251 14368 8760 14396
rect 8251 14365 8263 14368
rect 8205 14359 8263 14365
rect 8754 14356 8760 14368
rect 8812 14356 8818 14408
rect 9858 14396 9864 14408
rect 9819 14368 9864 14396
rect 9858 14356 9864 14368
rect 9916 14356 9922 14408
rect 13170 14396 13176 14408
rect 13131 14368 13176 14396
rect 13170 14356 13176 14368
rect 13228 14356 13234 14408
rect 8478 14328 8484 14340
rect 7300 14300 8484 14328
rect 8478 14288 8484 14300
rect 8536 14328 8542 14340
rect 9214 14328 9220 14340
rect 8536 14300 9220 14328
rect 8536 14288 8542 14300
rect 9214 14288 9220 14300
rect 9272 14288 9278 14340
rect 9674 14288 9680 14340
rect 9732 14328 9738 14340
rect 10505 14331 10563 14337
rect 10505 14328 10517 14331
rect 9732 14300 10517 14328
rect 9732 14288 9738 14300
rect 10505 14297 10517 14300
rect 10551 14297 10563 14331
rect 10505 14291 10563 14297
rect 11422 14288 11428 14340
rect 11480 14328 11486 14340
rect 12342 14328 12348 14340
rect 11480 14300 12348 14328
rect 11480 14288 11486 14300
rect 12342 14288 12348 14300
rect 12400 14328 12406 14340
rect 13464 14328 13492 14427
rect 13998 14424 14004 14436
rect 14056 14424 14062 14476
rect 15746 14464 15752 14476
rect 15707 14436 15752 14464
rect 15746 14424 15752 14436
rect 15804 14424 15810 14476
rect 16114 14464 16120 14476
rect 16075 14436 16120 14464
rect 16114 14424 16120 14436
rect 16172 14424 16178 14476
rect 16868 14473 16896 14504
rect 18322 14492 18328 14504
rect 18380 14492 18386 14544
rect 19334 14532 19340 14544
rect 18432 14504 19340 14532
rect 16853 14467 16911 14473
rect 16853 14433 16865 14467
rect 16899 14433 16911 14467
rect 16853 14427 16911 14433
rect 17505 14467 17563 14473
rect 17505 14433 17517 14467
rect 17551 14433 17563 14467
rect 17505 14427 17563 14433
rect 15473 14399 15531 14405
rect 15473 14365 15485 14399
rect 15519 14396 15531 14399
rect 15838 14396 15844 14408
rect 15519 14368 15844 14396
rect 15519 14365 15531 14368
rect 15473 14359 15531 14365
rect 15838 14356 15844 14368
rect 15896 14356 15902 14408
rect 17512 14396 17540 14427
rect 17770 14424 17776 14476
rect 17828 14464 17834 14476
rect 18432 14473 18460 14504
rect 19334 14492 19340 14504
rect 19392 14492 19398 14544
rect 20916 14541 20944 14572
rect 21652 14572 22192 14600
rect 20901 14535 20959 14541
rect 20901 14501 20913 14535
rect 20947 14501 20959 14535
rect 20901 14495 20959 14501
rect 18417 14467 18475 14473
rect 18417 14464 18429 14467
rect 17828 14436 18429 14464
rect 17828 14424 17834 14436
rect 18417 14433 18429 14436
rect 18463 14433 18475 14467
rect 19058 14464 19064 14476
rect 19019 14436 19064 14464
rect 18417 14427 18475 14433
rect 19058 14424 19064 14436
rect 19116 14424 19122 14476
rect 19150 14424 19156 14476
rect 19208 14464 19214 14476
rect 19794 14464 19800 14476
rect 19208 14436 19253 14464
rect 19755 14436 19800 14464
rect 19208 14424 19214 14436
rect 19794 14424 19800 14436
rect 19852 14424 19858 14476
rect 19886 14424 19892 14476
rect 19944 14464 19950 14476
rect 21652 14473 21680 14572
rect 22186 14560 22192 14572
rect 22244 14600 22250 14612
rect 23382 14600 23388 14612
rect 22244 14572 23388 14600
rect 22244 14560 22250 14572
rect 23382 14560 23388 14572
rect 23440 14560 23446 14612
rect 25682 14560 25688 14612
rect 25740 14600 25746 14612
rect 26142 14600 26148 14612
rect 25740 14572 26148 14600
rect 25740 14560 25746 14572
rect 26142 14560 26148 14572
rect 26200 14600 26206 14612
rect 26973 14603 27031 14609
rect 26973 14600 26985 14603
rect 26200 14572 26985 14600
rect 26200 14560 26206 14572
rect 26973 14569 26985 14572
rect 27019 14569 27031 14603
rect 26973 14563 27031 14569
rect 27062 14560 27068 14612
rect 27120 14600 27126 14612
rect 28626 14600 28632 14612
rect 27120 14572 28632 14600
rect 27120 14560 27126 14572
rect 28626 14560 28632 14572
rect 28684 14560 28690 14612
rect 28721 14603 28779 14609
rect 28721 14569 28733 14603
rect 28767 14600 28779 14603
rect 30098 14600 30104 14612
rect 28767 14572 30104 14600
rect 28767 14569 28779 14572
rect 28721 14563 28779 14569
rect 21910 14492 21916 14544
rect 21968 14532 21974 14544
rect 27430 14532 27436 14544
rect 21968 14504 23336 14532
rect 21968 14492 21974 14504
rect 20073 14467 20131 14473
rect 20073 14464 20085 14467
rect 19944 14436 20085 14464
rect 19944 14424 19950 14436
rect 20073 14433 20085 14436
rect 20119 14464 20131 14467
rect 21453 14467 21511 14473
rect 20119 14436 20576 14464
rect 20119 14433 20131 14436
rect 20073 14427 20131 14433
rect 18046 14396 18052 14408
rect 17512 14368 18052 14396
rect 18046 14356 18052 14368
rect 18104 14396 18110 14408
rect 19242 14396 19248 14408
rect 18104 14368 19248 14396
rect 18104 14356 18110 14368
rect 19242 14356 19248 14368
rect 19300 14356 19306 14408
rect 19429 14399 19487 14405
rect 19429 14365 19441 14399
rect 19475 14396 19487 14399
rect 20438 14396 20444 14408
rect 19475 14368 20444 14396
rect 19475 14365 19487 14368
rect 19429 14359 19487 14365
rect 20438 14356 20444 14368
rect 20496 14356 20502 14408
rect 13906 14328 13912 14340
rect 12400 14300 13492 14328
rect 13867 14300 13912 14328
rect 12400 14288 12406 14300
rect 13906 14288 13912 14300
rect 13964 14288 13970 14340
rect 14274 14288 14280 14340
rect 14332 14328 14338 14340
rect 16117 14331 16175 14337
rect 16117 14328 16129 14331
rect 14332 14300 16129 14328
rect 14332 14288 14338 14300
rect 16117 14297 16129 14300
rect 16163 14297 16175 14331
rect 16117 14291 16175 14297
rect 17494 14288 17500 14340
rect 17552 14328 17558 14340
rect 17589 14331 17647 14337
rect 17589 14328 17601 14331
rect 17552 14300 17601 14328
rect 17552 14288 17558 14300
rect 17589 14297 17601 14300
rect 17635 14297 17647 14331
rect 20548 14328 20576 14436
rect 21453 14433 21465 14467
rect 21499 14433 21511 14467
rect 21453 14427 21511 14433
rect 21637 14467 21695 14473
rect 21637 14433 21649 14467
rect 21683 14433 21695 14467
rect 21818 14464 21824 14476
rect 21779 14436 21824 14464
rect 21637 14427 21695 14433
rect 21468 14396 21496 14427
rect 21818 14424 21824 14436
rect 21876 14424 21882 14476
rect 22005 14467 22063 14473
rect 22005 14433 22017 14467
rect 22051 14464 22063 14467
rect 22094 14464 22100 14476
rect 22051 14436 22100 14464
rect 22051 14433 22063 14436
rect 22005 14427 22063 14433
rect 22094 14424 22100 14436
rect 22152 14424 22158 14476
rect 22278 14464 22284 14476
rect 22239 14436 22284 14464
rect 22278 14424 22284 14436
rect 22336 14424 22342 14476
rect 22738 14464 22744 14476
rect 22388 14436 22744 14464
rect 22388 14396 22416 14436
rect 22738 14424 22744 14436
rect 22796 14424 22802 14476
rect 23308 14473 23336 14504
rect 27172 14504 27436 14532
rect 23293 14467 23351 14473
rect 23293 14433 23305 14467
rect 23339 14433 23351 14467
rect 23293 14427 23351 14433
rect 23382 14424 23388 14476
rect 23440 14464 23446 14476
rect 23477 14467 23535 14473
rect 23477 14464 23489 14467
rect 23440 14436 23489 14464
rect 23440 14424 23446 14436
rect 23477 14433 23489 14436
rect 23523 14433 23535 14467
rect 23477 14427 23535 14433
rect 23661 14467 23719 14473
rect 23661 14433 23673 14467
rect 23707 14433 23719 14467
rect 23661 14427 23719 14433
rect 22830 14396 22836 14408
rect 21468 14368 22416 14396
rect 22791 14368 22836 14396
rect 22830 14356 22836 14368
rect 22888 14356 22894 14408
rect 23198 14356 23204 14408
rect 23256 14396 23262 14408
rect 23676 14396 23704 14427
rect 23750 14424 23756 14476
rect 23808 14464 23814 14476
rect 23845 14467 23903 14473
rect 23845 14464 23857 14467
rect 23808 14436 23857 14464
rect 23808 14424 23814 14436
rect 23845 14433 23857 14436
rect 23891 14433 23903 14467
rect 24118 14464 24124 14476
rect 24079 14436 24124 14464
rect 23845 14427 23903 14433
rect 24118 14424 24124 14436
rect 24176 14424 24182 14476
rect 24765 14467 24823 14473
rect 24765 14433 24777 14467
rect 24811 14464 24823 14467
rect 24946 14464 24952 14476
rect 24811 14436 24952 14464
rect 24811 14433 24823 14436
rect 24765 14427 24823 14433
rect 24946 14424 24952 14436
rect 25004 14424 25010 14476
rect 25501 14467 25559 14473
rect 25501 14433 25513 14467
rect 25547 14464 25559 14467
rect 25958 14464 25964 14476
rect 25547 14436 25964 14464
rect 25547 14433 25559 14436
rect 25501 14427 25559 14433
rect 25958 14424 25964 14436
rect 26016 14424 26022 14476
rect 27172 14473 27200 14504
rect 27430 14492 27436 14504
rect 27488 14492 27494 14544
rect 27157 14467 27215 14473
rect 27157 14433 27169 14467
rect 27203 14433 27215 14467
rect 27338 14464 27344 14476
rect 27299 14436 27344 14464
rect 27157 14427 27215 14433
rect 27338 14424 27344 14436
rect 27396 14424 27402 14476
rect 27709 14467 27767 14473
rect 27709 14433 27721 14467
rect 27755 14464 27767 14467
rect 27982 14464 27988 14476
rect 27755 14436 27988 14464
rect 27755 14433 27767 14436
rect 27709 14427 27767 14433
rect 27982 14424 27988 14436
rect 28040 14424 28046 14476
rect 23256 14368 23704 14396
rect 25777 14399 25835 14405
rect 23256 14356 23262 14368
rect 25777 14365 25789 14399
rect 25823 14396 25835 14399
rect 26786 14396 26792 14408
rect 25823 14368 26792 14396
rect 25823 14365 25835 14368
rect 25777 14359 25835 14365
rect 26786 14356 26792 14368
rect 26844 14356 26850 14408
rect 28736 14396 28764 14563
rect 30098 14560 30104 14572
rect 30156 14560 30162 14612
rect 30558 14600 30564 14612
rect 30519 14572 30564 14600
rect 30558 14560 30564 14572
rect 30616 14560 30622 14612
rect 32858 14600 32864 14612
rect 32819 14572 32864 14600
rect 32858 14560 32864 14572
rect 32916 14560 32922 14612
rect 33962 14560 33968 14612
rect 34020 14600 34026 14612
rect 37829 14603 37887 14609
rect 37829 14600 37841 14603
rect 34020 14572 37841 14600
rect 34020 14560 34026 14572
rect 37829 14569 37841 14572
rect 37875 14569 37887 14603
rect 37829 14563 37887 14569
rect 33502 14532 33508 14544
rect 29472 14504 33508 14532
rect 28905 14467 28963 14473
rect 28905 14433 28917 14467
rect 28951 14464 28963 14467
rect 28994 14464 29000 14476
rect 28951 14436 29000 14464
rect 28951 14433 28963 14436
rect 28905 14427 28963 14433
rect 28994 14424 29000 14436
rect 29052 14424 29058 14476
rect 29472 14473 29500 14504
rect 33502 14492 33508 14504
rect 33560 14492 33566 14544
rect 34514 14532 34520 14544
rect 34440 14504 34520 14532
rect 29457 14467 29515 14473
rect 29457 14433 29469 14467
rect 29503 14433 29515 14467
rect 29638 14464 29644 14476
rect 29599 14436 29644 14464
rect 29457 14427 29515 14433
rect 29638 14424 29644 14436
rect 29696 14424 29702 14476
rect 29825 14467 29883 14473
rect 29825 14433 29837 14467
rect 29871 14464 29883 14467
rect 30374 14464 30380 14476
rect 29871 14436 30380 14464
rect 29871 14433 29883 14436
rect 29825 14427 29883 14433
rect 30374 14424 30380 14436
rect 30432 14424 30438 14476
rect 30742 14464 30748 14476
rect 30703 14436 30748 14464
rect 30742 14424 30748 14436
rect 30800 14424 30806 14476
rect 30926 14464 30932 14476
rect 30887 14436 30932 14464
rect 30926 14424 30932 14436
rect 30984 14424 30990 14476
rect 32677 14467 32735 14473
rect 32677 14433 32689 14467
rect 32723 14464 32735 14467
rect 32766 14464 32772 14476
rect 32723 14436 32772 14464
rect 32723 14433 32735 14436
rect 32677 14427 32735 14433
rect 32766 14424 32772 14436
rect 32824 14424 32830 14476
rect 32950 14424 32956 14476
rect 33008 14464 33014 14476
rect 34440 14473 34468 14504
rect 34514 14492 34520 14504
rect 34572 14492 34578 14544
rect 34790 14532 34796 14544
rect 34624 14504 34796 14532
rect 34624 14473 34652 14504
rect 34790 14492 34796 14504
rect 34848 14532 34854 14544
rect 35434 14532 35440 14544
rect 34848 14504 35440 14532
rect 34848 14492 34854 14504
rect 35434 14492 35440 14504
rect 35492 14492 35498 14544
rect 36096 14504 37780 14532
rect 33413 14467 33471 14473
rect 33413 14464 33425 14467
rect 33008 14436 33425 14464
rect 33008 14424 33014 14436
rect 33413 14433 33425 14436
rect 33459 14433 33471 14467
rect 33413 14427 33471 14433
rect 34425 14467 34483 14473
rect 34425 14433 34437 14467
rect 34471 14433 34483 14467
rect 34425 14427 34483 14433
rect 34609 14467 34667 14473
rect 34609 14433 34621 14467
rect 34655 14433 34667 14467
rect 34609 14427 34667 14433
rect 34698 14424 34704 14476
rect 34756 14464 34762 14476
rect 35069 14467 35127 14473
rect 35069 14464 35081 14467
rect 34756 14436 35081 14464
rect 34756 14424 34762 14436
rect 35069 14433 35081 14436
rect 35115 14433 35127 14467
rect 35069 14427 35127 14433
rect 35342 14424 35348 14476
rect 35400 14464 35406 14476
rect 36096 14464 36124 14504
rect 36262 14464 36268 14476
rect 35400 14436 36124 14464
rect 36223 14436 36268 14464
rect 35400 14424 35406 14436
rect 36262 14424 36268 14436
rect 36320 14424 36326 14476
rect 36449 14467 36507 14473
rect 36449 14433 36461 14467
rect 36495 14433 36507 14467
rect 36630 14464 36636 14476
rect 36591 14436 36636 14464
rect 36449 14427 36507 14433
rect 27172 14368 28764 14396
rect 27172 14340 27200 14368
rect 32214 14356 32220 14408
rect 32272 14396 32278 14408
rect 32968 14396 32996 14424
rect 32272 14368 32996 14396
rect 32272 14356 32278 14368
rect 34514 14356 34520 14408
rect 34572 14396 34578 14408
rect 35710 14396 35716 14408
rect 34572 14368 35716 14396
rect 34572 14356 34578 14368
rect 35710 14356 35716 14368
rect 35768 14396 35774 14408
rect 36464 14396 36492 14427
rect 36630 14424 36636 14436
rect 36688 14424 36694 14476
rect 37752 14473 37780 14504
rect 37737 14467 37795 14473
rect 37737 14433 37749 14467
rect 37783 14433 37795 14467
rect 37737 14427 37795 14433
rect 35768 14368 36492 14396
rect 35768 14356 35774 14368
rect 23658 14328 23664 14340
rect 20548 14300 23664 14328
rect 17589 14291 17647 14297
rect 23658 14288 23664 14300
rect 23716 14288 23722 14340
rect 24026 14288 24032 14340
rect 24084 14328 24090 14340
rect 24857 14331 24915 14337
rect 24857 14328 24869 14331
rect 24084 14300 24869 14328
rect 24084 14288 24090 14300
rect 24857 14297 24869 14300
rect 24903 14297 24915 14331
rect 24857 14291 24915 14297
rect 27154 14288 27160 14340
rect 27212 14288 27218 14340
rect 29273 14331 29331 14337
rect 29273 14297 29285 14331
rect 29319 14328 29331 14331
rect 30466 14328 30472 14340
rect 29319 14300 30472 14328
rect 29319 14297 29331 14300
rect 29273 14291 29331 14297
rect 30466 14288 30472 14300
rect 30524 14288 30530 14340
rect 34606 14288 34612 14340
rect 34664 14328 34670 14340
rect 35069 14331 35127 14337
rect 35069 14328 35081 14331
rect 34664 14300 35081 14328
rect 34664 14288 34670 14300
rect 35069 14297 35081 14300
rect 35115 14297 35127 14331
rect 35069 14291 35127 14297
rect 36081 14331 36139 14337
rect 36081 14297 36093 14331
rect 36127 14328 36139 14331
rect 37182 14328 37188 14340
rect 36127 14300 37188 14328
rect 36127 14297 36139 14300
rect 36081 14291 36139 14297
rect 37182 14288 37188 14300
rect 37240 14288 37246 14340
rect 1394 14220 1400 14272
rect 1452 14260 1458 14272
rect 3697 14263 3755 14269
rect 3697 14260 3709 14263
rect 1452 14232 3709 14260
rect 1452 14220 1458 14232
rect 3697 14229 3709 14232
rect 3743 14229 3755 14263
rect 3697 14223 3755 14229
rect 5810 14220 5816 14272
rect 5868 14260 5874 14272
rect 7469 14263 7527 14269
rect 7469 14260 7481 14263
rect 5868 14232 7481 14260
rect 5868 14220 5874 14232
rect 7469 14229 7481 14232
rect 7515 14260 7527 14263
rect 16758 14260 16764 14272
rect 7515 14232 16764 14260
rect 7515 14229 7527 14232
rect 7469 14223 7527 14229
rect 16758 14220 16764 14232
rect 16816 14220 16822 14272
rect 16942 14260 16948 14272
rect 16903 14232 16948 14260
rect 16942 14220 16948 14232
rect 17000 14220 17006 14272
rect 17678 14220 17684 14272
rect 17736 14260 17742 14272
rect 22922 14260 22928 14272
rect 17736 14232 22928 14260
rect 17736 14220 17742 14232
rect 22922 14220 22928 14232
rect 22980 14220 22986 14272
rect 28718 14220 28724 14272
rect 28776 14260 28782 14272
rect 29546 14260 29552 14272
rect 28776 14232 29552 14260
rect 28776 14220 28782 14232
rect 29546 14220 29552 14232
rect 29604 14260 29610 14272
rect 32766 14260 32772 14272
rect 29604 14232 32772 14260
rect 29604 14220 29610 14232
rect 32766 14220 32772 14232
rect 32824 14220 32830 14272
rect 33502 14220 33508 14272
rect 33560 14260 33566 14272
rect 33597 14263 33655 14269
rect 33597 14260 33609 14263
rect 33560 14232 33609 14260
rect 33560 14220 33566 14232
rect 33597 14229 33609 14232
rect 33643 14229 33655 14263
rect 33597 14223 33655 14229
rect 1104 14170 38824 14192
rect 1104 14118 4246 14170
rect 4298 14118 4310 14170
rect 4362 14118 4374 14170
rect 4426 14118 4438 14170
rect 4490 14118 34966 14170
rect 35018 14118 35030 14170
rect 35082 14118 35094 14170
rect 35146 14118 35158 14170
rect 35210 14118 38824 14170
rect 1104 14096 38824 14118
rect 2130 14016 2136 14068
rect 2188 14056 2194 14068
rect 5350 14056 5356 14068
rect 2188 14028 5356 14056
rect 2188 14016 2194 14028
rect 5350 14016 5356 14028
rect 5408 14016 5414 14068
rect 7760 14028 8892 14056
rect 1854 13920 1860 13932
rect 1815 13892 1860 13920
rect 1854 13880 1860 13892
rect 1912 13880 1918 13932
rect 2133 13923 2191 13929
rect 2133 13889 2145 13923
rect 2179 13920 2191 13923
rect 4065 13923 4123 13929
rect 4065 13920 4077 13923
rect 2179 13892 4077 13920
rect 2179 13889 2191 13892
rect 2133 13883 2191 13889
rect 4065 13889 4077 13892
rect 4111 13889 4123 13923
rect 4065 13883 4123 13889
rect 3970 13852 3976 13864
rect 3931 13824 3976 13852
rect 3970 13812 3976 13824
rect 4028 13812 4034 13864
rect 4617 13855 4675 13861
rect 4617 13821 4629 13855
rect 4663 13821 4675 13855
rect 4982 13852 4988 13864
rect 4943 13824 4988 13852
rect 4617 13815 4675 13821
rect 4632 13784 4660 13815
rect 4982 13812 4988 13824
rect 5040 13812 5046 13864
rect 5353 13855 5411 13861
rect 5353 13821 5365 13855
rect 5399 13852 5411 13855
rect 5442 13852 5448 13864
rect 5399 13824 5448 13852
rect 5399 13821 5411 13824
rect 5353 13815 5411 13821
rect 5442 13812 5448 13824
rect 5500 13812 5506 13864
rect 5902 13852 5908 13864
rect 5863 13824 5908 13852
rect 5902 13812 5908 13824
rect 5960 13812 5966 13864
rect 6914 13812 6920 13864
rect 6972 13852 6978 13864
rect 7760 13861 7788 14028
rect 8018 13988 8024 14000
rect 7979 13960 8024 13988
rect 8018 13948 8024 13960
rect 8076 13948 8082 14000
rect 8864 13988 8892 14028
rect 8938 14016 8944 14068
rect 8996 14056 9002 14068
rect 10505 14059 10563 14065
rect 10505 14056 10517 14059
rect 8996 14028 10517 14056
rect 8996 14016 9002 14028
rect 10505 14025 10517 14028
rect 10551 14025 10563 14059
rect 10505 14019 10563 14025
rect 16301 14059 16359 14065
rect 16301 14025 16313 14059
rect 16347 14056 16359 14059
rect 16482 14056 16488 14068
rect 16347 14028 16488 14056
rect 16347 14025 16359 14028
rect 16301 14019 16359 14025
rect 16482 14016 16488 14028
rect 16540 14016 16546 14068
rect 17126 14016 17132 14068
rect 17184 14056 17190 14068
rect 17770 14056 17776 14068
rect 17184 14028 17776 14056
rect 17184 14016 17190 14028
rect 17770 14016 17776 14028
rect 17828 14016 17834 14068
rect 18966 14016 18972 14068
rect 19024 14056 19030 14068
rect 21545 14059 21603 14065
rect 21545 14056 21557 14059
rect 19024 14028 21557 14056
rect 19024 14016 19030 14028
rect 21545 14025 21557 14028
rect 21591 14025 21603 14059
rect 21545 14019 21603 14025
rect 21818 14016 21824 14068
rect 21876 14056 21882 14068
rect 21876 14028 24532 14056
rect 21876 14016 21882 14028
rect 11422 13988 11428 14000
rect 8864 13960 11428 13988
rect 11422 13948 11428 13960
rect 11480 13948 11486 14000
rect 13262 13988 13268 14000
rect 13223 13960 13268 13988
rect 13262 13948 13268 13960
rect 13320 13948 13326 14000
rect 15286 13948 15292 14000
rect 15344 13988 15350 14000
rect 17037 13991 17095 13997
rect 17037 13988 17049 13991
rect 15344 13960 17049 13988
rect 15344 13948 15350 13960
rect 17037 13957 17049 13960
rect 17083 13957 17095 13991
rect 17037 13951 17095 13957
rect 19242 13948 19248 14000
rect 19300 13988 19306 14000
rect 19429 13991 19487 13997
rect 19429 13988 19441 13991
rect 19300 13960 19441 13988
rect 19300 13948 19306 13960
rect 19429 13957 19441 13960
rect 19475 13957 19487 13991
rect 19429 13951 19487 13957
rect 8849 13923 8907 13929
rect 8849 13920 8861 13923
rect 8128 13892 8861 13920
rect 8128 13861 8156 13892
rect 8849 13889 8861 13892
rect 8895 13889 8907 13923
rect 9766 13920 9772 13932
rect 8849 13883 8907 13889
rect 9048 13892 9772 13920
rect 9048 13861 9076 13892
rect 9766 13880 9772 13892
rect 9824 13880 9830 13932
rect 10870 13920 10876 13932
rect 10520 13892 10876 13920
rect 7377 13855 7435 13861
rect 7377 13852 7389 13855
rect 6972 13824 7389 13852
rect 6972 13812 6978 13824
rect 7377 13821 7389 13824
rect 7423 13821 7435 13855
rect 7377 13815 7435 13821
rect 7745 13855 7803 13861
rect 7745 13821 7757 13855
rect 7791 13821 7803 13855
rect 7745 13815 7803 13821
rect 8113 13855 8171 13861
rect 8113 13821 8125 13855
rect 8159 13821 8171 13855
rect 8113 13815 8171 13821
rect 9033 13855 9091 13861
rect 9033 13821 9045 13855
rect 9079 13821 9091 13855
rect 9033 13815 9091 13821
rect 9401 13855 9459 13861
rect 9401 13821 9413 13855
rect 9447 13852 9459 13855
rect 9582 13852 9588 13864
rect 9447 13824 9588 13852
rect 9447 13821 9459 13824
rect 9401 13815 9459 13821
rect 4890 13784 4896 13796
rect 4632 13756 4896 13784
rect 4890 13744 4896 13756
rect 4948 13744 4954 13796
rect 7392 13784 7420 13815
rect 9582 13812 9588 13824
rect 9640 13812 9646 13864
rect 9677 13855 9735 13861
rect 9677 13821 9689 13855
rect 9723 13852 9735 13855
rect 10520 13852 10548 13892
rect 10870 13880 10876 13892
rect 10928 13920 10934 13932
rect 12621 13923 12679 13929
rect 10928 13892 11192 13920
rect 10928 13880 10934 13892
rect 10686 13852 10692 13864
rect 9723 13824 10548 13852
rect 10647 13824 10692 13852
rect 9723 13821 9735 13824
rect 9677 13815 9735 13821
rect 10686 13812 10692 13824
rect 10744 13812 10750 13864
rect 11054 13852 11060 13864
rect 11015 13824 11060 13852
rect 11054 13812 11060 13824
rect 11112 13812 11118 13864
rect 11164 13861 11192 13892
rect 12621 13889 12633 13923
rect 12667 13920 12679 13923
rect 12710 13920 12716 13932
rect 12667 13892 12716 13920
rect 12667 13889 12679 13892
rect 12621 13883 12679 13889
rect 12710 13880 12716 13892
rect 12768 13880 12774 13932
rect 14274 13920 14280 13932
rect 14235 13892 14280 13920
rect 14274 13880 14280 13892
rect 14332 13880 14338 13932
rect 15102 13880 15108 13932
rect 15160 13920 15166 13932
rect 15381 13923 15439 13929
rect 15381 13920 15393 13923
rect 15160 13892 15393 13920
rect 15160 13880 15166 13892
rect 15381 13889 15393 13892
rect 15427 13889 15439 13923
rect 15381 13883 15439 13889
rect 18049 13923 18107 13929
rect 18049 13889 18061 13923
rect 18095 13920 18107 13923
rect 18095 13892 18460 13920
rect 18095 13889 18107 13892
rect 18049 13883 18107 13889
rect 11149 13855 11207 13861
rect 11149 13821 11161 13855
rect 11195 13821 11207 13855
rect 12802 13852 12808 13864
rect 11149 13815 11207 13821
rect 12360 13824 12480 13852
rect 12763 13824 12808 13852
rect 12360 13784 12388 13824
rect 7392 13756 12388 13784
rect 3326 13676 3332 13728
rect 3384 13716 3390 13728
rect 3421 13719 3479 13725
rect 3421 13716 3433 13719
rect 3384 13688 3433 13716
rect 3384 13676 3390 13688
rect 3421 13685 3433 13688
rect 3467 13685 3479 13719
rect 12452 13716 12480 13824
rect 12802 13812 12808 13824
rect 12860 13812 12866 13864
rect 13357 13855 13415 13861
rect 13357 13821 13369 13855
rect 13403 13852 13415 13855
rect 13446 13852 13452 13864
rect 13403 13824 13452 13852
rect 13403 13821 13415 13824
rect 13357 13815 13415 13821
rect 13446 13812 13452 13824
rect 13504 13812 13510 13864
rect 14001 13855 14059 13861
rect 14001 13821 14013 13855
rect 14047 13852 14059 13855
rect 15010 13852 15016 13864
rect 14047 13824 15016 13852
rect 14047 13821 14059 13824
rect 14001 13815 14059 13821
rect 15010 13812 15016 13824
rect 15068 13812 15074 13864
rect 16117 13855 16175 13861
rect 16117 13821 16129 13855
rect 16163 13852 16175 13855
rect 16853 13855 16911 13861
rect 16853 13852 16865 13855
rect 16163 13824 16865 13852
rect 16163 13821 16175 13824
rect 16117 13815 16175 13821
rect 16853 13821 16865 13824
rect 16899 13852 16911 13855
rect 17678 13852 17684 13864
rect 16899 13824 17684 13852
rect 16899 13821 16911 13824
rect 16853 13815 16911 13821
rect 17678 13812 17684 13824
rect 17736 13812 17742 13864
rect 18322 13852 18328 13864
rect 18283 13824 18328 13852
rect 18322 13812 18328 13824
rect 18380 13812 18386 13864
rect 18432 13852 18460 13892
rect 18506 13880 18512 13932
rect 18564 13920 18570 13932
rect 20438 13920 20444 13932
rect 18564 13892 20300 13920
rect 20399 13892 20444 13920
rect 18564 13880 18570 13892
rect 20162 13852 20168 13864
rect 18432 13824 20168 13852
rect 20162 13812 20168 13824
rect 20220 13812 20226 13864
rect 20272 13852 20300 13892
rect 20438 13880 20444 13892
rect 20496 13880 20502 13932
rect 22370 13920 22376 13932
rect 22283 13892 22376 13920
rect 22370 13880 22376 13892
rect 22428 13920 22434 13932
rect 23014 13920 23020 13932
rect 22428 13892 23020 13920
rect 22428 13880 22434 13892
rect 23014 13880 23020 13892
rect 23072 13920 23078 13932
rect 23661 13923 23719 13929
rect 23661 13920 23673 13923
rect 23072 13892 23673 13920
rect 23072 13880 23078 13892
rect 23661 13889 23673 13892
rect 23707 13889 23719 13923
rect 23661 13883 23719 13889
rect 24397 13923 24455 13929
rect 24397 13889 24409 13923
rect 24443 13920 24455 13923
rect 24504 13920 24532 14028
rect 26234 14016 26240 14068
rect 26292 14056 26298 14068
rect 28626 14056 28632 14068
rect 26292 14028 27568 14056
rect 28539 14028 28632 14056
rect 26292 14016 26298 14028
rect 26786 13988 26792 14000
rect 26747 13960 26792 13988
rect 26786 13948 26792 13960
rect 26844 13948 26850 14000
rect 27540 13929 27568 14028
rect 28626 14016 28632 14028
rect 28684 14056 28690 14068
rect 29638 14056 29644 14068
rect 28684 14028 29644 14056
rect 28684 14016 28690 14028
rect 29638 14016 29644 14028
rect 29696 14016 29702 14068
rect 34330 14056 34336 14068
rect 34243 14028 34336 14056
rect 34330 14016 34336 14028
rect 34388 14056 34394 14068
rect 36078 14056 36084 14068
rect 34388 14028 36084 14056
rect 34388 14016 34394 14028
rect 36078 14016 36084 14028
rect 36136 14056 36142 14068
rect 36446 14056 36452 14068
rect 36136 14028 36452 14056
rect 36136 14016 36142 14028
rect 36446 14016 36452 14028
rect 36504 14016 36510 14068
rect 31386 13988 31392 14000
rect 29564 13960 31392 13988
rect 24443 13892 24532 13920
rect 27525 13923 27583 13929
rect 24443 13889 24455 13892
rect 24397 13883 24455 13889
rect 27525 13889 27537 13923
rect 27571 13889 27583 13923
rect 27525 13883 27583 13889
rect 23109 13855 23167 13861
rect 23109 13852 23121 13855
rect 20272 13824 23121 13852
rect 23109 13821 23121 13824
rect 23155 13821 23167 13855
rect 23109 13815 23167 13821
rect 23290 13812 23296 13864
rect 23348 13852 23354 13864
rect 23348 13824 23704 13852
rect 23348 13812 23354 13824
rect 18138 13784 18144 13796
rect 16868 13756 18144 13784
rect 16868 13716 16896 13756
rect 18138 13744 18144 13756
rect 18196 13744 18202 13796
rect 22649 13787 22707 13793
rect 22649 13784 22661 13787
rect 22480 13756 22661 13784
rect 12452 13688 16896 13716
rect 3421 13679 3479 13685
rect 17310 13676 17316 13728
rect 17368 13716 17374 13728
rect 20070 13716 20076 13728
rect 17368 13688 20076 13716
rect 17368 13676 17374 13688
rect 20070 13676 20076 13688
rect 20128 13676 20134 13728
rect 21726 13676 21732 13728
rect 21784 13716 21790 13728
rect 22480 13716 22508 13756
rect 22649 13753 22661 13756
rect 22695 13753 22707 13787
rect 22649 13747 22707 13753
rect 22741 13787 22799 13793
rect 22741 13753 22753 13787
rect 22787 13784 22799 13787
rect 23474 13784 23480 13796
rect 22787 13756 23480 13784
rect 22787 13753 22799 13756
rect 22741 13747 22799 13753
rect 23474 13744 23480 13756
rect 23532 13744 23538 13796
rect 23676 13784 23704 13824
rect 23750 13812 23756 13864
rect 23808 13852 23814 13864
rect 23937 13855 23995 13861
rect 23937 13852 23949 13855
rect 23808 13824 23949 13852
rect 23808 13812 23814 13824
rect 23937 13821 23949 13824
rect 23983 13821 23995 13855
rect 23937 13815 23995 13821
rect 24578 13812 24584 13864
rect 24636 13852 24642 13864
rect 25041 13855 25099 13861
rect 25041 13852 25053 13855
rect 24636 13824 25053 13852
rect 24636 13812 24642 13824
rect 25041 13821 25053 13824
rect 25087 13821 25099 13855
rect 25041 13815 25099 13821
rect 25225 13855 25283 13861
rect 25225 13821 25237 13855
rect 25271 13821 25283 13855
rect 25225 13815 25283 13821
rect 24029 13787 24087 13793
rect 24029 13784 24041 13787
rect 23676 13756 24041 13784
rect 24029 13753 24041 13756
rect 24075 13753 24087 13787
rect 25240 13784 25268 13815
rect 25314 13812 25320 13864
rect 25372 13852 25378 13864
rect 25685 13855 25743 13861
rect 25685 13852 25697 13855
rect 25372 13824 25697 13852
rect 25372 13812 25378 13824
rect 25685 13821 25697 13824
rect 25731 13821 25743 13855
rect 25685 13815 25743 13821
rect 26145 13855 26203 13861
rect 26145 13821 26157 13855
rect 26191 13852 26203 13855
rect 26234 13852 26240 13864
rect 26191 13824 26240 13852
rect 26191 13821 26203 13824
rect 26145 13815 26203 13821
rect 26234 13812 26240 13824
rect 26292 13812 26298 13864
rect 26697 13855 26755 13861
rect 26697 13821 26709 13855
rect 26743 13821 26755 13855
rect 26697 13815 26755 13821
rect 25866 13784 25872 13796
rect 25240 13756 25872 13784
rect 24029 13747 24087 13753
rect 25866 13744 25872 13756
rect 25924 13784 25930 13796
rect 26712 13784 26740 13815
rect 27062 13812 27068 13864
rect 27120 13852 27126 13864
rect 27249 13855 27307 13861
rect 27249 13852 27261 13855
rect 27120 13824 27261 13852
rect 27120 13812 27126 13824
rect 27249 13821 27261 13824
rect 27295 13821 27307 13855
rect 27249 13815 27307 13821
rect 28445 13855 28503 13861
rect 28445 13821 28457 13855
rect 28491 13852 28503 13855
rect 28626 13852 28632 13864
rect 28491 13824 28632 13852
rect 28491 13821 28503 13824
rect 28445 13815 28503 13821
rect 28626 13812 28632 13824
rect 28684 13812 28690 13864
rect 29564 13861 29592 13960
rect 31386 13948 31392 13960
rect 31444 13948 31450 14000
rect 33778 13988 33784 14000
rect 32600 13960 33784 13988
rect 29733 13923 29791 13929
rect 29733 13889 29745 13923
rect 29779 13920 29791 13923
rect 30926 13920 30932 13932
rect 29779 13892 30932 13920
rect 29779 13889 29791 13892
rect 29733 13883 29791 13889
rect 30926 13880 30932 13892
rect 30984 13880 30990 13932
rect 29549 13855 29607 13861
rect 29549 13821 29561 13855
rect 29595 13821 29607 13855
rect 29822 13852 29828 13864
rect 29783 13824 29828 13852
rect 29549 13815 29607 13821
rect 29822 13812 29828 13824
rect 29880 13812 29886 13864
rect 30193 13855 30251 13861
rect 30193 13821 30205 13855
rect 30239 13821 30251 13855
rect 30466 13852 30472 13864
rect 30427 13824 30472 13852
rect 30193 13815 30251 13821
rect 25924 13756 26740 13784
rect 25924 13744 25930 13756
rect 21784 13688 22508 13716
rect 22557 13719 22615 13725
rect 21784 13676 21790 13688
rect 22557 13685 22569 13719
rect 22603 13716 22615 13719
rect 23566 13716 23572 13728
rect 22603 13688 23572 13716
rect 22603 13685 22615 13688
rect 22557 13679 22615 13685
rect 23566 13676 23572 13688
rect 23624 13716 23630 13728
rect 23845 13719 23903 13725
rect 23845 13716 23857 13719
rect 23624 13688 23857 13716
rect 23624 13676 23630 13688
rect 23845 13685 23857 13688
rect 23891 13716 23903 13719
rect 23934 13716 23940 13728
rect 23891 13688 23940 13716
rect 23891 13685 23903 13688
rect 23845 13679 23903 13685
rect 23934 13676 23940 13688
rect 23992 13676 23998 13728
rect 24854 13716 24860 13728
rect 24815 13688 24860 13716
rect 24854 13676 24860 13688
rect 24912 13676 24918 13728
rect 25225 13719 25283 13725
rect 25225 13685 25237 13719
rect 25271 13716 25283 13719
rect 25682 13716 25688 13728
rect 25271 13688 25688 13716
rect 25271 13685 25283 13688
rect 25225 13679 25283 13685
rect 25682 13676 25688 13688
rect 25740 13676 25746 13728
rect 30208 13716 30236 13815
rect 30466 13812 30472 13824
rect 30524 13812 30530 13864
rect 31205 13855 31263 13861
rect 31205 13852 31217 13855
rect 30576 13824 31217 13852
rect 30282 13744 30288 13796
rect 30340 13784 30346 13796
rect 30576 13784 30604 13824
rect 31205 13821 31217 13824
rect 31251 13821 31263 13855
rect 32122 13852 32128 13864
rect 32083 13824 32128 13852
rect 31205 13815 31263 13821
rect 32122 13812 32128 13824
rect 32180 13812 32186 13864
rect 32600 13861 32628 13960
rect 33778 13948 33784 13960
rect 33836 13988 33842 14000
rect 36262 13988 36268 14000
rect 33836 13960 36268 13988
rect 33836 13948 33842 13960
rect 36262 13948 36268 13960
rect 36320 13948 36326 14000
rect 33226 13920 33232 13932
rect 33187 13892 33232 13920
rect 33226 13880 33232 13892
rect 33284 13880 33290 13932
rect 33962 13920 33968 13932
rect 33888 13892 33968 13920
rect 32585 13855 32643 13861
rect 32585 13821 32597 13855
rect 32631 13821 32643 13855
rect 32766 13852 32772 13864
rect 32727 13824 32772 13852
rect 32585 13815 32643 13821
rect 32766 13812 32772 13824
rect 32824 13812 32830 13864
rect 33318 13852 33324 13864
rect 33279 13824 33324 13852
rect 33318 13812 33324 13824
rect 33376 13812 33382 13864
rect 33888 13861 33916 13892
rect 33962 13880 33968 13892
rect 34020 13880 34026 13932
rect 34238 13880 34244 13932
rect 34296 13920 34302 13932
rect 35434 13920 35440 13932
rect 34296 13892 35440 13920
rect 34296 13880 34302 13892
rect 35434 13880 35440 13892
rect 35492 13880 35498 13932
rect 37829 13923 37887 13929
rect 37829 13920 37841 13923
rect 35544 13892 37841 13920
rect 35544 13861 35572 13892
rect 37829 13889 37841 13892
rect 37875 13889 37887 13923
rect 37829 13883 37887 13889
rect 33873 13855 33931 13861
rect 33873 13821 33885 13855
rect 33919 13821 33931 13855
rect 34517 13855 34575 13861
rect 34517 13852 34529 13855
rect 33873 13815 33931 13821
rect 33980 13824 34529 13852
rect 33980 13784 34008 13824
rect 34517 13821 34529 13824
rect 34563 13821 34575 13855
rect 34517 13815 34575 13821
rect 35529 13855 35587 13861
rect 35529 13821 35541 13855
rect 35575 13821 35587 13855
rect 35986 13852 35992 13864
rect 35947 13824 35992 13852
rect 35529 13815 35587 13821
rect 35986 13812 35992 13824
rect 36044 13812 36050 13864
rect 36446 13852 36452 13864
rect 36407 13824 36452 13852
rect 36446 13812 36452 13824
rect 36504 13812 36510 13864
rect 36538 13812 36544 13864
rect 36596 13852 36602 13864
rect 36725 13855 36783 13861
rect 36725 13852 36737 13855
rect 36596 13824 36737 13852
rect 36596 13812 36602 13824
rect 36725 13821 36737 13824
rect 36771 13821 36783 13855
rect 36725 13815 36783 13821
rect 30340 13756 30604 13784
rect 33704 13756 34008 13784
rect 30340 13744 30346 13756
rect 33704 13728 33732 13756
rect 30650 13716 30656 13728
rect 30208 13688 30656 13716
rect 30650 13676 30656 13688
rect 30708 13676 30714 13728
rect 31386 13716 31392 13728
rect 31347 13688 31392 13716
rect 31386 13676 31392 13688
rect 31444 13676 31450 13728
rect 31938 13716 31944 13728
rect 31899 13688 31944 13716
rect 31938 13676 31944 13688
rect 31996 13676 32002 13728
rect 33686 13676 33692 13728
rect 33744 13676 33750 13728
rect 1104 13626 38824 13648
rect 1104 13574 19606 13626
rect 19658 13574 19670 13626
rect 19722 13574 19734 13626
rect 19786 13574 19798 13626
rect 19850 13574 38824 13626
rect 1104 13552 38824 13574
rect 1670 13512 1676 13524
rect 1631 13484 1676 13512
rect 1670 13472 1676 13484
rect 1728 13472 1734 13524
rect 10686 13472 10692 13524
rect 10744 13512 10750 13524
rect 10962 13512 10968 13524
rect 10744 13484 10968 13512
rect 10744 13472 10750 13484
rect 10962 13472 10968 13484
rect 11020 13512 11026 13524
rect 11057 13515 11115 13521
rect 11057 13512 11069 13515
rect 11020 13484 11069 13512
rect 11020 13472 11026 13484
rect 11057 13481 11069 13484
rect 11103 13481 11115 13515
rect 14645 13515 14703 13521
rect 14645 13512 14657 13515
rect 11057 13475 11115 13481
rect 11164 13484 14657 13512
rect 3970 13404 3976 13456
rect 4028 13444 4034 13456
rect 4028 13416 5396 13444
rect 4028 13404 4034 13416
rect 1762 13376 1768 13388
rect 1723 13348 1768 13376
rect 1762 13336 1768 13348
rect 1820 13336 1826 13388
rect 2133 13379 2191 13385
rect 2133 13345 2145 13379
rect 2179 13345 2191 13379
rect 3326 13376 3332 13388
rect 3287 13348 3332 13376
rect 2133 13339 2191 13345
rect 2148 13308 2176 13339
rect 3326 13336 3332 13348
rect 3384 13336 3390 13388
rect 4065 13379 4123 13385
rect 4065 13345 4077 13379
rect 4111 13376 4123 13379
rect 4614 13376 4620 13388
rect 4111 13348 4620 13376
rect 4111 13345 4123 13348
rect 4065 13339 4123 13345
rect 4614 13336 4620 13348
rect 4672 13336 4678 13388
rect 5368 13385 5396 13416
rect 4709 13379 4767 13385
rect 4709 13345 4721 13379
rect 4755 13376 4767 13379
rect 5353 13379 5411 13385
rect 4755 13348 5304 13376
rect 4755 13345 4767 13348
rect 4709 13339 4767 13345
rect 3421 13311 3479 13317
rect 3421 13308 3433 13311
rect 2148 13280 3433 13308
rect 3421 13277 3433 13280
rect 3467 13308 3479 13311
rect 4890 13308 4896 13320
rect 3467 13280 4896 13308
rect 3467 13277 3479 13280
rect 3421 13271 3479 13277
rect 4890 13268 4896 13280
rect 4948 13268 4954 13320
rect 5276 13308 5304 13348
rect 5353 13345 5365 13379
rect 5399 13345 5411 13379
rect 5353 13339 5411 13345
rect 5994 13336 6000 13388
rect 6052 13376 6058 13388
rect 6089 13379 6147 13385
rect 6089 13376 6101 13379
rect 6052 13348 6101 13376
rect 6052 13336 6058 13348
rect 6089 13345 6101 13348
rect 6135 13345 6147 13379
rect 8662 13376 8668 13388
rect 6089 13339 6147 13345
rect 6196 13348 7512 13376
rect 8623 13348 8668 13376
rect 6196 13308 6224 13348
rect 6362 13308 6368 13320
rect 5276 13280 6224 13308
rect 6323 13280 6368 13308
rect 6362 13268 6368 13280
rect 6420 13268 6426 13320
rect 7484 13317 7512 13348
rect 8662 13336 8668 13348
rect 8720 13336 8726 13388
rect 9674 13376 9680 13388
rect 9635 13348 9680 13376
rect 9674 13336 9680 13348
rect 9732 13336 9738 13388
rect 9950 13376 9956 13388
rect 9911 13348 9956 13376
rect 9950 13336 9956 13348
rect 10008 13336 10014 13388
rect 10226 13336 10232 13388
rect 10284 13376 10290 13388
rect 11164 13376 11192 13484
rect 14645 13481 14657 13484
rect 14691 13481 14703 13515
rect 19058 13512 19064 13524
rect 19019 13484 19064 13512
rect 14645 13475 14703 13481
rect 19058 13472 19064 13484
rect 19116 13472 19122 13524
rect 23474 13512 23480 13524
rect 23387 13484 23480 13512
rect 23474 13472 23480 13484
rect 23532 13512 23538 13524
rect 24213 13515 24271 13521
rect 23532 13484 24072 13512
rect 23532 13472 23538 13484
rect 15470 13444 15476 13456
rect 13924 13416 15476 13444
rect 10284 13348 11192 13376
rect 12437 13379 12495 13385
rect 10284 13336 10290 13348
rect 12437 13345 12449 13379
rect 12483 13376 12495 13379
rect 13262 13376 13268 13388
rect 12483 13348 13268 13376
rect 12483 13345 12495 13348
rect 12437 13339 12495 13345
rect 13262 13336 13268 13348
rect 13320 13336 13326 13388
rect 7469 13311 7527 13317
rect 7469 13277 7481 13311
rect 7515 13277 7527 13311
rect 7469 13271 7527 13277
rect 12161 13311 12219 13317
rect 12161 13277 12173 13311
rect 12207 13308 12219 13311
rect 13924 13308 13952 13416
rect 15470 13404 15476 13416
rect 15528 13404 15534 13456
rect 17494 13444 17500 13456
rect 17236 13416 17500 13444
rect 14461 13379 14519 13385
rect 14461 13345 14473 13379
rect 14507 13345 14519 13379
rect 14461 13339 14519 13345
rect 12207 13280 13952 13308
rect 14476 13308 14504 13339
rect 14550 13336 14556 13388
rect 14608 13376 14614 13388
rect 14608 13348 14653 13376
rect 14608 13336 14614 13348
rect 14918 13336 14924 13388
rect 14976 13376 14982 13388
rect 15289 13379 15347 13385
rect 15289 13376 15301 13379
rect 14976 13348 15301 13376
rect 14976 13336 14982 13348
rect 15289 13345 15301 13348
rect 15335 13345 15347 13379
rect 16022 13376 16028 13388
rect 15983 13348 16028 13376
rect 15289 13339 15347 13345
rect 16022 13336 16028 13348
rect 16080 13336 16086 13388
rect 16761 13379 16819 13385
rect 16761 13345 16773 13379
rect 16807 13376 16819 13379
rect 17126 13376 17132 13388
rect 16807 13348 17132 13376
rect 16807 13345 16819 13348
rect 16761 13339 16819 13345
rect 17126 13336 17132 13348
rect 17184 13336 17190 13388
rect 17236 13385 17264 13416
rect 17494 13404 17500 13416
rect 17552 13404 17558 13456
rect 17954 13444 17960 13456
rect 17696 13416 17960 13444
rect 17221 13379 17279 13385
rect 17221 13345 17233 13379
rect 17267 13345 17279 13379
rect 17221 13339 17279 13345
rect 17405 13379 17463 13385
rect 17405 13345 17417 13379
rect 17451 13376 17463 13379
rect 17696 13376 17724 13416
rect 17954 13404 17960 13416
rect 18012 13444 18018 13456
rect 19242 13444 19248 13456
rect 18012 13416 19248 13444
rect 18012 13404 18018 13416
rect 19242 13404 19248 13416
rect 19300 13404 19306 13456
rect 21726 13404 21732 13456
rect 21784 13444 21790 13456
rect 23492 13444 23520 13472
rect 21784 13416 22140 13444
rect 21784 13404 21790 13416
rect 17862 13376 17868 13388
rect 17451 13348 17724 13376
rect 17823 13348 17868 13376
rect 17451 13345 17463 13348
rect 17405 13339 17463 13345
rect 17862 13336 17868 13348
rect 17920 13336 17926 13388
rect 18138 13336 18144 13388
rect 18196 13376 18202 13388
rect 18233 13379 18291 13385
rect 18233 13376 18245 13379
rect 18196 13348 18245 13376
rect 18196 13336 18202 13348
rect 18233 13345 18245 13348
rect 18279 13376 18291 13379
rect 18414 13376 18420 13388
rect 18279 13348 18420 13376
rect 18279 13345 18291 13348
rect 18233 13339 18291 13345
rect 18414 13336 18420 13348
rect 18472 13336 18478 13388
rect 18966 13376 18972 13388
rect 18927 13348 18972 13376
rect 18966 13336 18972 13348
rect 19024 13336 19030 13388
rect 19426 13336 19432 13388
rect 19484 13376 19490 13388
rect 19613 13379 19671 13385
rect 19613 13376 19625 13379
rect 19484 13348 19625 13376
rect 19484 13336 19490 13348
rect 19613 13345 19625 13348
rect 19659 13345 19671 13379
rect 19613 13339 19671 13345
rect 19978 13336 19984 13388
rect 20036 13376 20042 13388
rect 20073 13379 20131 13385
rect 20073 13376 20085 13379
rect 20036 13348 20085 13376
rect 20036 13336 20042 13348
rect 20073 13345 20085 13348
rect 20119 13345 20131 13379
rect 21910 13376 21916 13388
rect 21871 13348 21916 13376
rect 20073 13339 20131 13345
rect 21910 13336 21916 13348
rect 21968 13336 21974 13388
rect 22112 13385 22140 13416
rect 22756 13416 23520 13444
rect 22097 13379 22155 13385
rect 22097 13345 22109 13379
rect 22143 13345 22155 13379
rect 22097 13339 22155 13345
rect 22186 13336 22192 13388
rect 22244 13376 22250 13388
rect 22756 13385 22784 13416
rect 22465 13379 22523 13385
rect 22244 13348 22289 13376
rect 22244 13336 22250 13348
rect 22465 13345 22477 13379
rect 22511 13345 22523 13379
rect 22465 13339 22523 13345
rect 22741 13379 22799 13385
rect 22741 13345 22753 13379
rect 22787 13345 22799 13379
rect 23290 13376 23296 13388
rect 23251 13348 23296 13376
rect 22741 13339 22799 13345
rect 17310 13308 17316 13320
rect 14476 13280 17316 13308
rect 12207 13277 12219 13280
rect 12161 13271 12219 13277
rect 17310 13268 17316 13280
rect 17368 13268 17374 13320
rect 17589 13311 17647 13317
rect 17589 13277 17601 13311
rect 17635 13308 17647 13311
rect 18322 13308 18328 13320
rect 17635 13280 18328 13308
rect 17635 13277 17647 13280
rect 17589 13271 17647 13277
rect 18322 13268 18328 13280
rect 18380 13268 18386 13320
rect 20349 13311 20407 13317
rect 20349 13277 20361 13311
rect 20395 13308 20407 13311
rect 21174 13308 21180 13320
rect 20395 13280 21180 13308
rect 20395 13277 20407 13280
rect 20349 13271 20407 13277
rect 21174 13268 21180 13280
rect 21232 13268 21238 13320
rect 21358 13308 21364 13320
rect 21319 13280 21364 13308
rect 21358 13268 21364 13280
rect 21416 13268 21422 13320
rect 22480 13308 22508 13339
rect 23290 13336 23296 13348
rect 23348 13336 23354 13388
rect 24044 13385 24072 13484
rect 24213 13481 24225 13515
rect 24259 13512 24271 13515
rect 24302 13512 24308 13524
rect 24259 13484 24308 13512
rect 24259 13481 24271 13484
rect 24213 13475 24271 13481
rect 24302 13472 24308 13484
rect 24360 13472 24366 13524
rect 28350 13512 28356 13524
rect 28311 13484 28356 13512
rect 28350 13472 28356 13484
rect 28408 13472 28414 13524
rect 32858 13512 32864 13524
rect 29288 13484 32864 13512
rect 27614 13444 27620 13456
rect 27080 13416 27620 13444
rect 24029 13379 24087 13385
rect 24029 13345 24041 13379
rect 24075 13376 24087 13379
rect 24118 13376 24124 13388
rect 24075 13348 24124 13376
rect 24075 13345 24087 13348
rect 24029 13339 24087 13345
rect 24118 13336 24124 13348
rect 24176 13336 24182 13388
rect 25038 13376 25044 13388
rect 24999 13348 25044 13376
rect 25038 13336 25044 13348
rect 25096 13336 25102 13388
rect 25501 13379 25559 13385
rect 25501 13345 25513 13379
rect 25547 13345 25559 13379
rect 25682 13376 25688 13388
rect 25643 13348 25688 13376
rect 25501 13339 25559 13345
rect 23198 13308 23204 13320
rect 22480 13280 23204 13308
rect 23198 13268 23204 13280
rect 23256 13268 23262 13320
rect 4801 13243 4859 13249
rect 4801 13209 4813 13243
rect 4847 13240 4859 13243
rect 5994 13240 6000 13252
rect 4847 13212 6000 13240
rect 4847 13209 4859 13212
rect 4801 13203 4859 13209
rect 5994 13200 6000 13212
rect 6052 13200 6058 13252
rect 11422 13200 11428 13252
rect 11480 13240 11486 13252
rect 11480 13212 11744 13240
rect 11480 13200 11486 13212
rect 4157 13175 4215 13181
rect 4157 13141 4169 13175
rect 4203 13172 4215 13175
rect 4614 13172 4620 13184
rect 4203 13144 4620 13172
rect 4203 13141 4215 13144
rect 4157 13135 4215 13141
rect 4614 13132 4620 13144
rect 4672 13132 4678 13184
rect 5537 13175 5595 13181
rect 5537 13141 5549 13175
rect 5583 13172 5595 13175
rect 7006 13172 7012 13184
rect 5583 13144 7012 13172
rect 5583 13141 5595 13144
rect 5537 13135 5595 13141
rect 7006 13132 7012 13144
rect 7064 13132 7070 13184
rect 8849 13175 8907 13181
rect 8849 13141 8861 13175
rect 8895 13172 8907 13175
rect 9398 13172 9404 13184
rect 8895 13144 9404 13172
rect 8895 13141 8907 13144
rect 8849 13135 8907 13141
rect 9398 13132 9404 13144
rect 9456 13132 9462 13184
rect 11716 13172 11744 13212
rect 14182 13200 14188 13252
rect 14240 13240 14246 13252
rect 14277 13243 14335 13249
rect 14277 13240 14289 13243
rect 14240 13212 14289 13240
rect 14240 13200 14246 13212
rect 14277 13209 14289 13212
rect 14323 13240 14335 13243
rect 14458 13240 14464 13252
rect 14323 13212 14464 13240
rect 14323 13209 14335 13212
rect 14277 13203 14335 13209
rect 14458 13200 14464 13212
rect 14516 13200 14522 13252
rect 14550 13200 14556 13252
rect 14608 13240 14614 13252
rect 14608 13212 23888 13240
rect 14608 13200 14614 13212
rect 13354 13172 13360 13184
rect 11716 13144 13360 13172
rect 13354 13132 13360 13144
rect 13412 13132 13418 13184
rect 13725 13175 13783 13181
rect 13725 13141 13737 13175
rect 13771 13172 13783 13175
rect 13906 13172 13912 13184
rect 13771 13144 13912 13172
rect 13771 13141 13783 13144
rect 13725 13135 13783 13141
rect 13906 13132 13912 13144
rect 13964 13132 13970 13184
rect 15378 13172 15384 13184
rect 15339 13144 15384 13172
rect 15378 13132 15384 13144
rect 15436 13132 15442 13184
rect 16942 13132 16948 13184
rect 17000 13172 17006 13184
rect 17862 13172 17868 13184
rect 17000 13144 17868 13172
rect 17000 13132 17006 13144
rect 17862 13132 17868 13144
rect 17920 13172 17926 13184
rect 19886 13172 19892 13184
rect 17920 13144 19892 13172
rect 17920 13132 17926 13144
rect 19886 13132 19892 13144
rect 19944 13172 19950 13184
rect 20530 13172 20536 13184
rect 19944 13144 20536 13172
rect 19944 13132 19950 13144
rect 20530 13132 20536 13144
rect 20588 13132 20594 13184
rect 23860 13172 23888 13212
rect 23934 13200 23940 13252
rect 23992 13240 23998 13252
rect 24949 13243 25007 13249
rect 24949 13240 24961 13243
rect 23992 13212 24961 13240
rect 23992 13200 23998 13212
rect 24949 13209 24961 13212
rect 24995 13209 25007 13243
rect 25516 13240 25544 13339
rect 25682 13336 25688 13348
rect 25740 13336 25746 13388
rect 27080 13385 27108 13416
rect 27614 13404 27620 13416
rect 27672 13404 27678 13456
rect 27065 13379 27123 13385
rect 27065 13345 27077 13379
rect 27111 13345 27123 13379
rect 27338 13376 27344 13388
rect 27299 13348 27344 13376
rect 27065 13339 27123 13345
rect 27338 13336 27344 13348
rect 27396 13336 27402 13388
rect 27522 13336 27528 13388
rect 27580 13376 27586 13388
rect 28166 13376 28172 13388
rect 27580 13348 27844 13376
rect 28127 13348 28172 13376
rect 27580 13336 27586 13348
rect 26697 13311 26755 13317
rect 26697 13277 26709 13311
rect 26743 13308 26755 13311
rect 27706 13308 27712 13320
rect 26743 13280 27712 13308
rect 26743 13277 26755 13280
rect 26697 13271 26755 13277
rect 27706 13268 27712 13280
rect 27764 13268 27770 13320
rect 27816 13308 27844 13348
rect 28166 13336 28172 13348
rect 28224 13336 28230 13388
rect 28810 13336 28816 13388
rect 28868 13376 28874 13388
rect 29089 13379 29147 13385
rect 29089 13376 29101 13379
rect 28868 13348 29101 13376
rect 28868 13336 28874 13348
rect 29089 13345 29101 13348
rect 29135 13376 29147 13379
rect 29288 13376 29316 13484
rect 29135 13348 29316 13376
rect 29365 13379 29423 13385
rect 29135 13345 29147 13348
rect 29089 13339 29147 13345
rect 29365 13345 29377 13379
rect 29411 13345 29423 13379
rect 29365 13339 29423 13345
rect 29917 13379 29975 13385
rect 29917 13345 29929 13379
rect 29963 13345 29975 13379
rect 30190 13376 30196 13388
rect 30151 13348 30196 13376
rect 29917 13339 29975 13345
rect 29380 13308 29408 13339
rect 29822 13308 29828 13320
rect 27816 13280 29408 13308
rect 29783 13280 29828 13308
rect 29822 13268 29828 13280
rect 29880 13268 29886 13320
rect 29932 13308 29960 13339
rect 30190 13336 30196 13348
rect 30248 13336 30254 13388
rect 30650 13376 30656 13388
rect 30611 13348 30656 13376
rect 30650 13336 30656 13348
rect 30708 13336 30714 13388
rect 31297 13379 31355 13385
rect 31297 13345 31309 13379
rect 31343 13345 31355 13379
rect 31297 13339 31355 13345
rect 30374 13308 30380 13320
rect 29932 13280 30380 13308
rect 30374 13268 30380 13280
rect 30432 13268 30438 13320
rect 27341 13243 27399 13249
rect 27341 13240 27353 13243
rect 25516 13212 27353 13240
rect 24949 13203 25007 13209
rect 27341 13209 27353 13212
rect 27387 13209 27399 13243
rect 27341 13203 27399 13209
rect 27798 13200 27804 13252
rect 27856 13240 27862 13252
rect 31312 13240 31340 13339
rect 31846 13336 31852 13388
rect 31904 13376 31910 13388
rect 32600 13385 32628 13484
rect 32858 13472 32864 13484
rect 32916 13472 32922 13524
rect 34054 13472 34060 13524
rect 34112 13512 34118 13524
rect 34330 13512 34336 13524
rect 34112 13484 34336 13512
rect 34112 13472 34118 13484
rect 34330 13472 34336 13484
rect 34388 13472 34394 13524
rect 34606 13472 34612 13524
rect 34664 13512 34670 13524
rect 35342 13512 35348 13524
rect 34664 13484 35348 13512
rect 34664 13472 34670 13484
rect 35342 13472 35348 13484
rect 35400 13512 35406 13524
rect 35437 13515 35495 13521
rect 35437 13512 35449 13515
rect 35400 13484 35449 13512
rect 35400 13472 35406 13484
rect 35437 13481 35449 13484
rect 35483 13481 35495 13515
rect 35437 13475 35495 13481
rect 32217 13379 32275 13385
rect 32217 13376 32229 13379
rect 31904 13348 32229 13376
rect 31904 13336 31910 13348
rect 32217 13345 32229 13348
rect 32263 13345 32275 13379
rect 32217 13339 32275 13345
rect 32585 13379 32643 13385
rect 32585 13345 32597 13379
rect 32631 13345 32643 13379
rect 32585 13339 32643 13345
rect 33045 13379 33103 13385
rect 33045 13345 33057 13379
rect 33091 13376 33103 13379
rect 33226 13376 33232 13388
rect 33091 13348 33232 13376
rect 33091 13345 33103 13348
rect 33045 13339 33103 13345
rect 33226 13336 33232 13348
rect 33284 13336 33290 13388
rect 33965 13379 34023 13385
rect 33965 13376 33977 13379
rect 33336 13348 33977 13376
rect 31938 13268 31944 13320
rect 31996 13308 32002 13320
rect 33336 13308 33364 13348
rect 33965 13345 33977 13348
rect 34011 13345 34023 13379
rect 37001 13379 37059 13385
rect 37001 13376 37013 13379
rect 33965 13339 34023 13345
rect 34992 13348 37013 13376
rect 34054 13308 34060 13320
rect 31996 13280 33364 13308
rect 34015 13280 34060 13308
rect 31996 13268 32002 13280
rect 34054 13268 34060 13280
rect 34112 13268 34118 13320
rect 34330 13308 34336 13320
rect 34291 13280 34336 13308
rect 34330 13268 34336 13280
rect 34388 13268 34394 13320
rect 27856 13212 31340 13240
rect 27856 13200 27862 13212
rect 32766 13200 32772 13252
rect 32824 13240 32830 13252
rect 33045 13243 33103 13249
rect 33045 13240 33057 13243
rect 32824 13212 33057 13240
rect 32824 13200 32830 13212
rect 33045 13209 33057 13212
rect 33091 13209 33103 13243
rect 33045 13203 33103 13209
rect 33134 13200 33140 13252
rect 33192 13240 33198 13252
rect 33192 13212 33916 13240
rect 33192 13200 33198 13212
rect 27062 13172 27068 13184
rect 23860 13144 27068 13172
rect 27062 13132 27068 13144
rect 27120 13172 27126 13184
rect 28718 13172 28724 13184
rect 27120 13144 28724 13172
rect 27120 13132 27126 13144
rect 28718 13132 28724 13144
rect 28776 13132 28782 13184
rect 31481 13175 31539 13181
rect 31481 13141 31493 13175
rect 31527 13172 31539 13175
rect 31570 13172 31576 13184
rect 31527 13144 31576 13172
rect 31527 13141 31539 13144
rect 31481 13135 31539 13141
rect 31570 13132 31576 13144
rect 31628 13172 31634 13184
rect 33318 13172 33324 13184
rect 31628 13144 33324 13172
rect 31628 13132 31634 13144
rect 33318 13132 33324 13144
rect 33376 13132 33382 13184
rect 33686 13132 33692 13184
rect 33744 13172 33750 13184
rect 33781 13175 33839 13181
rect 33781 13172 33793 13175
rect 33744 13144 33793 13172
rect 33744 13132 33750 13144
rect 33781 13141 33793 13144
rect 33827 13141 33839 13175
rect 33888 13172 33916 13212
rect 34992 13172 35020 13348
rect 37001 13345 37013 13348
rect 37047 13345 37059 13379
rect 37734 13376 37740 13388
rect 37695 13348 37740 13376
rect 37001 13339 37059 13345
rect 37734 13336 37740 13348
rect 37792 13336 37798 13388
rect 36170 13308 36176 13320
rect 36131 13280 36176 13308
rect 36170 13268 36176 13280
rect 36228 13268 36234 13320
rect 36262 13268 36268 13320
rect 36320 13308 36326 13320
rect 36725 13311 36783 13317
rect 36725 13308 36737 13311
rect 36320 13280 36737 13308
rect 36320 13268 36326 13280
rect 36725 13277 36737 13280
rect 36771 13277 36783 13311
rect 37182 13308 37188 13320
rect 37143 13280 37188 13308
rect 36725 13271 36783 13277
rect 37182 13268 37188 13280
rect 37240 13268 37246 13320
rect 33888 13144 35020 13172
rect 33781 13135 33839 13141
rect 35526 13132 35532 13184
rect 35584 13172 35590 13184
rect 37921 13175 37979 13181
rect 37921 13172 37933 13175
rect 35584 13144 37933 13172
rect 35584 13132 35590 13144
rect 37921 13141 37933 13144
rect 37967 13141 37979 13175
rect 37921 13135 37979 13141
rect 1104 13082 38824 13104
rect 1104 13030 4246 13082
rect 4298 13030 4310 13082
rect 4362 13030 4374 13082
rect 4426 13030 4438 13082
rect 4490 13030 34966 13082
rect 35018 13030 35030 13082
rect 35082 13030 35094 13082
rect 35146 13030 35158 13082
rect 35210 13030 38824 13082
rect 1104 13008 38824 13030
rect 6638 12928 6644 12980
rect 6696 12968 6702 12980
rect 7650 12968 7656 12980
rect 6696 12940 7656 12968
rect 6696 12928 6702 12940
rect 7650 12928 7656 12940
rect 7708 12928 7714 12980
rect 9398 12928 9404 12980
rect 9456 12968 9462 12980
rect 11238 12968 11244 12980
rect 9456 12940 11244 12968
rect 9456 12928 9462 12940
rect 11238 12928 11244 12940
rect 11296 12928 11302 12980
rect 11330 12928 11336 12980
rect 11388 12968 11394 12980
rect 22002 12968 22008 12980
rect 11388 12940 22008 12968
rect 11388 12928 11394 12940
rect 22002 12928 22008 12940
rect 22060 12928 22066 12980
rect 22278 12968 22284 12980
rect 22239 12940 22284 12968
rect 22278 12928 22284 12940
rect 22336 12968 22342 12980
rect 22646 12968 22652 12980
rect 22336 12940 22652 12968
rect 22336 12928 22342 12940
rect 22646 12928 22652 12940
rect 22704 12928 22710 12980
rect 28166 12928 28172 12980
rect 28224 12968 28230 12980
rect 36814 12968 36820 12980
rect 28224 12940 36820 12968
rect 28224 12928 28230 12940
rect 36814 12928 36820 12940
rect 36872 12928 36878 12980
rect 4982 12860 4988 12912
rect 5040 12860 5046 12912
rect 6362 12860 6368 12912
rect 6420 12900 6426 12912
rect 6917 12903 6975 12909
rect 6917 12900 6929 12903
rect 6420 12872 6929 12900
rect 6420 12860 6426 12872
rect 6917 12869 6929 12872
rect 6963 12869 6975 12903
rect 13170 12900 13176 12912
rect 6917 12863 6975 12869
rect 7024 12872 13176 12900
rect 1673 12835 1731 12841
rect 1673 12801 1685 12835
rect 1719 12832 1731 12835
rect 1854 12832 1860 12844
rect 1719 12804 1860 12832
rect 1719 12801 1731 12804
rect 1673 12795 1731 12801
rect 1854 12792 1860 12804
rect 1912 12792 1918 12844
rect 1949 12835 2007 12841
rect 1949 12801 1961 12835
rect 1995 12832 2007 12835
rect 3881 12835 3939 12841
rect 3881 12832 3893 12835
rect 1995 12804 3893 12832
rect 1995 12801 2007 12804
rect 1949 12795 2007 12801
rect 3881 12801 3893 12804
rect 3927 12801 3939 12835
rect 4614 12832 4620 12844
rect 3881 12795 3939 12801
rect 4448 12804 4620 12832
rect 3970 12764 3976 12776
rect 3931 12736 3976 12764
rect 3970 12724 3976 12736
rect 4028 12724 4034 12776
rect 4154 12724 4160 12776
rect 4212 12764 4218 12776
rect 4448 12773 4476 12804
rect 4614 12792 4620 12804
rect 4672 12792 4678 12844
rect 5000 12832 5028 12860
rect 7024 12832 7052 12872
rect 13170 12860 13176 12872
rect 13228 12860 13234 12912
rect 16666 12900 16672 12912
rect 13280 12872 15240 12900
rect 16627 12872 16672 12900
rect 4816 12804 5028 12832
rect 5736 12804 7052 12832
rect 9585 12835 9643 12841
rect 4816 12773 4844 12804
rect 4433 12767 4491 12773
rect 4433 12764 4445 12767
rect 4212 12736 4445 12764
rect 4212 12724 4218 12736
rect 4433 12733 4445 12736
rect 4479 12733 4491 12767
rect 4433 12727 4491 12733
rect 4801 12767 4859 12773
rect 4801 12733 4813 12767
rect 4847 12733 4859 12767
rect 4801 12727 4859 12733
rect 5169 12767 5227 12773
rect 5169 12733 5181 12767
rect 5215 12764 5227 12767
rect 5442 12764 5448 12776
rect 5215 12736 5448 12764
rect 5215 12733 5227 12736
rect 5169 12727 5227 12733
rect 5442 12724 5448 12736
rect 5500 12724 5506 12776
rect 5736 12773 5764 12804
rect 9585 12801 9597 12835
rect 9631 12832 9643 12835
rect 10870 12832 10876 12844
rect 9631 12804 10876 12832
rect 9631 12801 9643 12804
rect 9585 12795 9643 12801
rect 10870 12792 10876 12804
rect 10928 12792 10934 12844
rect 11146 12832 11152 12844
rect 11107 12804 11152 12832
rect 11146 12792 11152 12804
rect 11204 12792 11210 12844
rect 11882 12832 11888 12844
rect 11256 12804 11888 12832
rect 5721 12767 5779 12773
rect 5721 12733 5733 12767
rect 5767 12733 5779 12767
rect 6638 12764 6644 12776
rect 6599 12736 6644 12764
rect 5721 12727 5779 12733
rect 6638 12724 6644 12736
rect 6696 12724 6702 12776
rect 7006 12764 7012 12776
rect 6967 12736 7012 12764
rect 7006 12724 7012 12736
rect 7064 12724 7070 12776
rect 7285 12767 7343 12773
rect 7285 12733 7297 12767
rect 7331 12733 7343 12767
rect 7285 12727 7343 12733
rect 7561 12767 7619 12773
rect 7561 12733 7573 12767
rect 7607 12733 7619 12767
rect 8018 12764 8024 12776
rect 7979 12736 8024 12764
rect 7561 12727 7619 12733
rect 3329 12699 3387 12705
rect 3329 12665 3341 12699
rect 3375 12696 3387 12699
rect 4706 12696 4712 12708
rect 3375 12668 4712 12696
rect 3375 12665 3387 12668
rect 3329 12659 3387 12665
rect 4706 12656 4712 12668
rect 4764 12656 4770 12708
rect 5994 12656 6000 12708
rect 6052 12696 6058 12708
rect 7300 12696 7328 12727
rect 6052 12668 7328 12696
rect 6052 12656 6058 12668
rect 6656 12640 6684 12668
rect 6454 12628 6460 12640
rect 6415 12600 6460 12628
rect 6454 12588 6460 12600
rect 6512 12588 6518 12640
rect 6638 12588 6644 12640
rect 6696 12588 6702 12640
rect 6822 12588 6828 12640
rect 6880 12628 6886 12640
rect 7576 12628 7604 12727
rect 8018 12724 8024 12736
rect 8076 12724 8082 12776
rect 8754 12764 8760 12776
rect 8715 12736 8760 12764
rect 8754 12724 8760 12736
rect 8812 12724 8818 12776
rect 9398 12764 9404 12776
rect 9359 12736 9404 12764
rect 9398 12724 9404 12736
rect 9456 12724 9462 12776
rect 9766 12764 9772 12776
rect 9727 12736 9772 12764
rect 9766 12724 9772 12736
rect 9824 12724 9830 12776
rect 10597 12767 10655 12773
rect 10597 12733 10609 12767
rect 10643 12733 10655 12767
rect 10597 12727 10655 12733
rect 10965 12767 11023 12773
rect 10965 12733 10977 12767
rect 11011 12733 11023 12767
rect 10965 12727 11023 12733
rect 8294 12656 8300 12708
rect 8352 12696 8358 12708
rect 9490 12696 9496 12708
rect 8352 12668 9496 12696
rect 8352 12656 8358 12668
rect 9490 12656 9496 12668
rect 9548 12696 9554 12708
rect 10612 12696 10640 12727
rect 9548 12668 10640 12696
rect 10980 12696 11008 12727
rect 11054 12724 11060 12776
rect 11112 12764 11118 12776
rect 11256 12773 11284 12804
rect 11882 12792 11888 12804
rect 11940 12832 11946 12844
rect 13280 12832 13308 12872
rect 13446 12832 13452 12844
rect 11940 12804 13308 12832
rect 13407 12804 13452 12832
rect 11940 12792 11946 12804
rect 11241 12767 11299 12773
rect 11241 12764 11253 12767
rect 11112 12736 11253 12764
rect 11112 12724 11118 12736
rect 11241 12733 11253 12736
rect 11287 12733 11299 12767
rect 11422 12764 11428 12776
rect 11383 12736 11428 12764
rect 11241 12727 11299 12733
rect 11422 12724 11428 12736
rect 11480 12724 11486 12776
rect 13188 12773 13216 12804
rect 13446 12792 13452 12804
rect 13504 12792 13510 12844
rect 15212 12832 15240 12872
rect 16666 12860 16672 12872
rect 16724 12860 16730 12912
rect 16758 12860 16764 12912
rect 16816 12900 16822 12912
rect 28184 12900 28212 12928
rect 16816 12872 20852 12900
rect 16816 12860 16822 12872
rect 15286 12832 15292 12844
rect 15212 12804 15292 12832
rect 12897 12767 12955 12773
rect 12897 12733 12909 12767
rect 12943 12733 12955 12767
rect 12897 12727 12955 12733
rect 13173 12767 13231 12773
rect 13173 12733 13185 12767
rect 13219 12733 13231 12767
rect 13354 12764 13360 12776
rect 13315 12736 13360 12764
rect 13173 12727 13231 12733
rect 11330 12696 11336 12708
rect 10980 12668 11336 12696
rect 9548 12656 9554 12668
rect 11330 12656 11336 12668
rect 11388 12656 11394 12708
rect 12912 12696 12940 12727
rect 13354 12724 13360 12736
rect 13412 12724 13418 12776
rect 14642 12724 14648 12776
rect 14700 12764 14706 12776
rect 14921 12767 14979 12773
rect 14921 12764 14933 12767
rect 14700 12736 14933 12764
rect 14700 12724 14706 12736
rect 14921 12733 14933 12736
rect 14967 12764 14979 12767
rect 15102 12764 15108 12776
rect 14967 12736 15108 12764
rect 14967 12733 14979 12736
rect 14921 12727 14979 12733
rect 15102 12724 15108 12736
rect 15160 12724 15166 12776
rect 15212 12773 15240 12804
rect 15286 12792 15292 12804
rect 15344 12792 15350 12844
rect 15841 12835 15899 12841
rect 15841 12801 15853 12835
rect 15887 12832 15899 12835
rect 16114 12832 16120 12844
rect 15887 12804 16120 12832
rect 15887 12801 15899 12804
rect 15841 12795 15899 12801
rect 16114 12792 16120 12804
rect 16172 12792 16178 12844
rect 18785 12835 18843 12841
rect 18785 12801 18797 12835
rect 18831 12832 18843 12835
rect 19886 12832 19892 12844
rect 18831 12804 19564 12832
rect 19847 12804 19892 12832
rect 18831 12801 18843 12804
rect 18785 12795 18843 12801
rect 15197 12767 15255 12773
rect 15197 12733 15209 12767
rect 15243 12733 15255 12767
rect 15197 12727 15255 12733
rect 15657 12767 15715 12773
rect 15657 12733 15669 12767
rect 15703 12764 15715 12767
rect 15746 12764 15752 12776
rect 15703 12736 15752 12764
rect 15703 12733 15715 12736
rect 15657 12727 15715 12733
rect 15746 12724 15752 12736
rect 15804 12724 15810 12776
rect 16390 12764 16396 12776
rect 16351 12736 16396 12764
rect 16390 12724 16396 12736
rect 16448 12724 16454 12776
rect 16945 12767 17003 12773
rect 16945 12733 16957 12767
rect 16991 12733 17003 12767
rect 16945 12727 17003 12733
rect 17405 12767 17463 12773
rect 17405 12733 17417 12767
rect 17451 12764 17463 12767
rect 17954 12764 17960 12776
rect 17451 12736 17960 12764
rect 17451 12733 17463 12736
rect 17405 12727 17463 12733
rect 13906 12696 13912 12708
rect 12912 12668 13912 12696
rect 13906 12656 13912 12668
rect 13964 12656 13970 12708
rect 15286 12656 15292 12708
rect 15344 12696 15350 12708
rect 16960 12696 16988 12727
rect 17954 12724 17960 12736
rect 18012 12724 18018 12776
rect 18049 12767 18107 12773
rect 18049 12733 18061 12767
rect 18095 12764 18107 12767
rect 18506 12764 18512 12776
rect 18095 12736 18512 12764
rect 18095 12733 18107 12736
rect 18049 12727 18107 12733
rect 18506 12724 18512 12736
rect 18564 12724 18570 12776
rect 18693 12767 18751 12773
rect 18693 12733 18705 12767
rect 18739 12733 18751 12767
rect 19334 12764 19340 12776
rect 19295 12736 19340 12764
rect 18693 12727 18751 12733
rect 15344 12668 16988 12696
rect 18708 12696 18736 12727
rect 19334 12724 19340 12736
rect 19392 12724 19398 12776
rect 19536 12764 19564 12804
rect 19886 12792 19892 12804
rect 19944 12792 19950 12844
rect 19978 12764 19984 12776
rect 19536 12736 19984 12764
rect 19978 12724 19984 12736
rect 20036 12724 20042 12776
rect 20346 12764 20352 12776
rect 20307 12736 20352 12764
rect 20346 12724 20352 12736
rect 20404 12724 20410 12776
rect 20530 12764 20536 12776
rect 20491 12736 20536 12764
rect 20530 12724 20536 12736
rect 20588 12724 20594 12776
rect 20824 12764 20852 12872
rect 26160 12872 28212 12900
rect 30929 12903 30987 12909
rect 23474 12832 23480 12844
rect 22112 12804 23480 12832
rect 20990 12764 20996 12776
rect 20824 12736 20996 12764
rect 20990 12724 20996 12736
rect 21048 12724 21054 12776
rect 22112 12773 22140 12804
rect 23474 12792 23480 12804
rect 23532 12792 23538 12844
rect 23934 12832 23940 12844
rect 23895 12804 23940 12832
rect 23934 12792 23940 12804
rect 23992 12792 23998 12844
rect 22097 12767 22155 12773
rect 22097 12733 22109 12767
rect 22143 12733 22155 12767
rect 22097 12727 22155 12733
rect 22833 12767 22891 12773
rect 22833 12733 22845 12767
rect 22879 12764 22891 12767
rect 23566 12764 23572 12776
rect 22879 12736 23572 12764
rect 22879 12733 22891 12736
rect 22833 12727 22891 12733
rect 23566 12724 23572 12736
rect 23624 12724 23630 12776
rect 23661 12767 23719 12773
rect 23661 12733 23673 12767
rect 23707 12764 23719 12767
rect 23750 12764 23756 12776
rect 23707 12736 23756 12764
rect 23707 12733 23719 12736
rect 23661 12727 23719 12733
rect 19426 12696 19432 12708
rect 18708 12668 19432 12696
rect 15344 12656 15350 12668
rect 19426 12656 19432 12668
rect 19484 12656 19490 12708
rect 20254 12656 20260 12708
rect 20312 12696 20318 12708
rect 23676 12696 23704 12727
rect 23750 12724 23756 12736
rect 23808 12724 23814 12776
rect 24210 12724 24216 12776
rect 24268 12764 24274 12776
rect 24670 12764 24676 12776
rect 24268 12736 24676 12764
rect 24268 12724 24274 12736
rect 24670 12724 24676 12736
rect 24728 12724 24734 12776
rect 24854 12724 24860 12776
rect 24912 12764 24918 12776
rect 26053 12767 26111 12773
rect 26053 12764 26065 12767
rect 24912 12736 26065 12764
rect 24912 12724 24918 12736
rect 26053 12733 26065 12736
rect 26099 12733 26111 12767
rect 26053 12727 26111 12733
rect 20312 12668 23704 12696
rect 25317 12699 25375 12705
rect 20312 12656 20318 12668
rect 25317 12665 25329 12699
rect 25363 12696 25375 12699
rect 25498 12696 25504 12708
rect 25363 12668 25504 12696
rect 25363 12665 25375 12668
rect 25317 12659 25375 12665
rect 25498 12656 25504 12668
rect 25556 12656 25562 12708
rect 26160 12696 26188 12872
rect 30929 12869 30941 12903
rect 30975 12869 30987 12903
rect 31386 12900 31392 12912
rect 30929 12863 30987 12869
rect 31128 12872 31392 12900
rect 26697 12835 26755 12841
rect 26697 12801 26709 12835
rect 26743 12832 26755 12835
rect 27338 12832 27344 12844
rect 26743 12804 27344 12832
rect 26743 12801 26755 12804
rect 26697 12795 26755 12801
rect 27338 12792 27344 12804
rect 27396 12792 27402 12844
rect 30944 12832 30972 12863
rect 29932 12804 30972 12832
rect 26418 12724 26424 12776
rect 26476 12764 26482 12776
rect 26605 12767 26663 12773
rect 26605 12764 26617 12767
rect 26476 12736 26617 12764
rect 26476 12724 26482 12736
rect 26605 12733 26617 12736
rect 26651 12764 26663 12767
rect 27065 12767 27123 12773
rect 26651 12736 27016 12764
rect 26651 12733 26663 12736
rect 26605 12727 26663 12733
rect 25608 12668 26188 12696
rect 10410 12628 10416 12640
rect 6880 12600 7604 12628
rect 10371 12600 10416 12628
rect 6880 12588 6886 12600
rect 10410 12588 10416 12600
rect 10468 12588 10474 12640
rect 15746 12588 15752 12640
rect 15804 12628 15810 12640
rect 18141 12631 18199 12637
rect 18141 12628 18153 12631
rect 15804 12600 18153 12628
rect 15804 12588 15810 12600
rect 18141 12597 18153 12600
rect 18187 12597 18199 12631
rect 18141 12591 18199 12597
rect 18598 12588 18604 12640
rect 18656 12628 18662 12640
rect 20714 12628 20720 12640
rect 18656 12600 20720 12628
rect 18656 12588 18662 12600
rect 20714 12588 20720 12600
rect 20772 12588 20778 12640
rect 22922 12588 22928 12640
rect 22980 12628 22986 12640
rect 23017 12631 23075 12637
rect 23017 12628 23029 12631
rect 22980 12600 23029 12628
rect 22980 12588 22986 12600
rect 23017 12597 23029 12600
rect 23063 12628 23075 12631
rect 25608 12628 25636 12668
rect 25866 12628 25872 12640
rect 23063 12600 25636 12628
rect 25827 12600 25872 12628
rect 23063 12597 23075 12600
rect 23017 12591 23075 12597
rect 25866 12588 25872 12600
rect 25924 12588 25930 12640
rect 26988 12628 27016 12736
rect 27065 12733 27077 12767
rect 27111 12733 27123 12767
rect 27246 12764 27252 12776
rect 27207 12736 27252 12764
rect 27065 12727 27123 12733
rect 27080 12696 27108 12727
rect 27246 12724 27252 12736
rect 27304 12724 27310 12776
rect 27801 12767 27859 12773
rect 27801 12733 27813 12767
rect 27847 12764 27859 12767
rect 27890 12764 27896 12776
rect 27847 12736 27896 12764
rect 27847 12733 27859 12736
rect 27801 12727 27859 12733
rect 27890 12724 27896 12736
rect 27948 12724 27954 12776
rect 28261 12767 28319 12773
rect 28261 12733 28273 12767
rect 28307 12764 28319 12767
rect 28534 12764 28540 12776
rect 28307 12736 28540 12764
rect 28307 12733 28319 12736
rect 28261 12727 28319 12733
rect 28534 12724 28540 12736
rect 28592 12724 28598 12776
rect 29365 12767 29423 12773
rect 29365 12733 29377 12767
rect 29411 12764 29423 12767
rect 29638 12764 29644 12776
rect 29411 12736 29644 12764
rect 29411 12733 29423 12736
rect 29365 12727 29423 12733
rect 29638 12724 29644 12736
rect 29696 12724 29702 12776
rect 29932 12773 29960 12804
rect 29917 12767 29975 12773
rect 29917 12733 29929 12767
rect 29963 12733 29975 12767
rect 30098 12764 30104 12776
rect 30059 12736 30104 12764
rect 29917 12727 29975 12733
rect 30098 12724 30104 12736
rect 30156 12724 30162 12776
rect 31128 12773 31156 12872
rect 31386 12860 31392 12872
rect 31444 12900 31450 12912
rect 33505 12903 33563 12909
rect 31444 12872 32260 12900
rect 31444 12860 31450 12872
rect 32232 12773 32260 12872
rect 33505 12869 33517 12903
rect 33551 12900 33563 12903
rect 34330 12900 34336 12912
rect 33551 12872 34336 12900
rect 33551 12869 33563 12872
rect 33505 12863 33563 12869
rect 34330 12860 34336 12872
rect 34388 12860 34394 12912
rect 32401 12835 32459 12841
rect 32401 12801 32413 12835
rect 32447 12832 32459 12835
rect 35161 12835 35219 12841
rect 32447 12804 33824 12832
rect 32447 12801 32459 12804
rect 32401 12795 32459 12801
rect 31113 12767 31171 12773
rect 31113 12733 31125 12767
rect 31159 12733 31171 12767
rect 31113 12727 31171 12733
rect 31389 12767 31447 12773
rect 31389 12733 31401 12767
rect 31435 12733 31447 12767
rect 31389 12727 31447 12733
rect 32217 12767 32275 12773
rect 32217 12733 32229 12767
rect 32263 12733 32275 12767
rect 32766 12764 32772 12776
rect 32727 12736 32772 12764
rect 32217 12727 32275 12733
rect 27706 12696 27712 12708
rect 27080 12668 27712 12696
rect 27706 12656 27712 12668
rect 27764 12656 27770 12708
rect 29454 12656 29460 12708
rect 29512 12696 29518 12708
rect 31404 12696 31432 12727
rect 29512 12668 31432 12696
rect 32232 12696 32260 12727
rect 32766 12724 32772 12736
rect 32824 12724 32830 12776
rect 33796 12773 33824 12804
rect 35161 12801 35173 12835
rect 35207 12832 35219 12835
rect 35434 12832 35440 12844
rect 35207 12804 35440 12832
rect 35207 12801 35219 12804
rect 35161 12795 35219 12801
rect 35434 12792 35440 12804
rect 35492 12792 35498 12844
rect 35713 12835 35771 12841
rect 35713 12801 35725 12835
rect 35759 12832 35771 12835
rect 36538 12832 36544 12844
rect 35759 12804 36544 12832
rect 35759 12801 35771 12804
rect 35713 12795 35771 12801
rect 36538 12792 36544 12804
rect 36596 12792 36602 12844
rect 33229 12767 33287 12773
rect 33229 12733 33241 12767
rect 33275 12733 33287 12767
rect 33229 12727 33287 12733
rect 33781 12767 33839 12773
rect 33781 12733 33793 12767
rect 33827 12733 33839 12767
rect 34238 12764 34244 12776
rect 34199 12736 34244 12764
rect 33781 12727 33839 12733
rect 32950 12696 32956 12708
rect 32232 12668 32956 12696
rect 29512 12656 29518 12668
rect 32950 12656 32956 12668
rect 33008 12656 33014 12708
rect 29178 12628 29184 12640
rect 26988 12600 29184 12628
rect 29178 12588 29184 12600
rect 29236 12588 29242 12640
rect 29362 12628 29368 12640
rect 29323 12600 29368 12628
rect 29362 12588 29368 12600
rect 29420 12588 29426 12640
rect 29638 12588 29644 12640
rect 29696 12628 29702 12640
rect 29914 12628 29920 12640
rect 29696 12600 29920 12628
rect 29696 12588 29702 12600
rect 29914 12588 29920 12600
rect 29972 12628 29978 12640
rect 33244 12628 33272 12727
rect 34238 12724 34244 12736
rect 34296 12724 34302 12776
rect 35250 12724 35256 12776
rect 35308 12764 35314 12776
rect 35308 12736 35353 12764
rect 35308 12724 35314 12736
rect 36078 12724 36084 12776
rect 36136 12764 36142 12776
rect 36173 12767 36231 12773
rect 36173 12764 36185 12767
rect 36136 12736 36185 12764
rect 36136 12724 36142 12736
rect 36173 12733 36185 12736
rect 36219 12733 36231 12767
rect 36173 12727 36231 12733
rect 36449 12767 36507 12773
rect 36449 12733 36461 12767
rect 36495 12764 36507 12767
rect 36722 12764 36728 12776
rect 36495 12736 36728 12764
rect 36495 12733 36507 12736
rect 36449 12727 36507 12733
rect 36722 12724 36728 12736
rect 36780 12724 36786 12776
rect 37550 12628 37556 12640
rect 29972 12600 33272 12628
rect 37511 12600 37556 12628
rect 29972 12588 29978 12600
rect 37550 12588 37556 12600
rect 37608 12588 37614 12640
rect 1104 12538 38824 12560
rect 1104 12486 19606 12538
rect 19658 12486 19670 12538
rect 19722 12486 19734 12538
rect 19786 12486 19798 12538
rect 19850 12486 38824 12538
rect 1104 12464 38824 12486
rect 9858 12424 9864 12436
rect 4540 12396 7236 12424
rect 1394 12288 1400 12300
rect 1355 12260 1400 12288
rect 1394 12248 1400 12260
rect 1452 12248 1458 12300
rect 4341 12291 4399 12297
rect 4341 12257 4353 12291
rect 4387 12288 4399 12291
rect 4540 12288 4568 12396
rect 7006 12356 7012 12368
rect 6104 12328 7012 12356
rect 4706 12288 4712 12300
rect 4387 12260 4568 12288
rect 4667 12260 4712 12288
rect 4387 12257 4399 12260
rect 4341 12251 4399 12257
rect 4706 12248 4712 12260
rect 4764 12248 4770 12300
rect 5258 12288 5264 12300
rect 5219 12260 5264 12288
rect 5258 12248 5264 12260
rect 5316 12248 5322 12300
rect 6104 12297 6132 12328
rect 7006 12316 7012 12328
rect 7064 12316 7070 12368
rect 6089 12291 6147 12297
rect 6089 12257 6101 12291
rect 6135 12257 6147 12291
rect 6546 12288 6552 12300
rect 6507 12260 6552 12288
rect 6089 12251 6147 12257
rect 6546 12248 6552 12260
rect 6604 12248 6610 12300
rect 6822 12288 6828 12300
rect 6783 12260 6828 12288
rect 6822 12248 6828 12260
rect 6880 12248 6886 12300
rect 1670 12220 1676 12232
rect 1631 12192 1676 12220
rect 1670 12180 1676 12192
rect 1728 12180 1734 12232
rect 4433 12223 4491 12229
rect 4433 12189 4445 12223
rect 4479 12220 4491 12223
rect 4798 12220 4804 12232
rect 4479 12192 4804 12220
rect 4479 12189 4491 12192
rect 4433 12183 4491 12189
rect 4798 12180 4804 12192
rect 4856 12180 4862 12232
rect 5353 12223 5411 12229
rect 5353 12189 5365 12223
rect 5399 12220 5411 12223
rect 6564 12220 6592 12248
rect 5399 12192 6592 12220
rect 5399 12189 5411 12192
rect 5353 12183 5411 12189
rect 2958 12112 2964 12164
rect 3016 12152 3022 12164
rect 5997 12155 6055 12161
rect 5997 12152 6009 12155
rect 3016 12124 6009 12152
rect 3016 12112 3022 12124
rect 5997 12121 6009 12124
rect 6043 12121 6055 12155
rect 5997 12115 6055 12121
rect 7098 12112 7104 12164
rect 7156 12152 7162 12164
rect 7208 12152 7236 12396
rect 7852 12396 9864 12424
rect 7852 12297 7880 12396
rect 9858 12384 9864 12396
rect 9916 12424 9922 12436
rect 10686 12424 10692 12436
rect 9916 12396 10692 12424
rect 9916 12384 9922 12396
rect 10686 12384 10692 12396
rect 10744 12384 10750 12436
rect 10870 12384 10876 12436
rect 10928 12424 10934 12436
rect 15562 12424 15568 12436
rect 10928 12396 12756 12424
rect 15523 12396 15568 12424
rect 10928 12384 10934 12396
rect 9398 12356 9404 12368
rect 8588 12328 9404 12356
rect 8588 12297 8616 12328
rect 9398 12316 9404 12328
rect 9456 12316 9462 12368
rect 7285 12291 7343 12297
rect 7285 12257 7297 12291
rect 7331 12257 7343 12291
rect 7285 12251 7343 12257
rect 7837 12291 7895 12297
rect 7837 12257 7849 12291
rect 7883 12257 7895 12291
rect 7837 12251 7895 12257
rect 8573 12291 8631 12297
rect 8573 12257 8585 12291
rect 8619 12257 8631 12291
rect 9030 12288 9036 12300
rect 8991 12260 9036 12288
rect 8573 12251 8631 12257
rect 7300 12220 7328 12251
rect 9030 12248 9036 12260
rect 9088 12248 9094 12300
rect 9674 12248 9680 12300
rect 9732 12288 9738 12300
rect 9953 12291 10011 12297
rect 9953 12288 9965 12291
rect 9732 12260 9965 12288
rect 9732 12248 9738 12260
rect 9953 12257 9965 12260
rect 9999 12257 10011 12291
rect 9953 12251 10011 12257
rect 11974 12248 11980 12300
rect 12032 12288 12038 12300
rect 12728 12297 12756 12396
rect 15562 12384 15568 12396
rect 15620 12384 15626 12436
rect 18966 12424 18972 12436
rect 18524 12396 18972 12424
rect 16390 12356 16396 12368
rect 15948 12328 16396 12356
rect 12069 12291 12127 12297
rect 12069 12288 12081 12291
rect 12032 12260 12081 12288
rect 12032 12248 12038 12260
rect 12069 12257 12081 12260
rect 12115 12257 12127 12291
rect 12069 12251 12127 12257
rect 12713 12291 12771 12297
rect 12713 12257 12725 12291
rect 12759 12257 12771 12291
rect 13170 12288 13176 12300
rect 13131 12260 13176 12288
rect 12713 12251 12771 12257
rect 13170 12248 13176 12260
rect 13228 12248 13234 12300
rect 13725 12291 13783 12297
rect 13725 12257 13737 12291
rect 13771 12257 13783 12291
rect 14366 12288 14372 12300
rect 14327 12260 14372 12288
rect 13725 12251 13783 12257
rect 8018 12220 8024 12232
rect 7300 12192 8024 12220
rect 8018 12180 8024 12192
rect 8076 12180 8082 12232
rect 10229 12223 10287 12229
rect 10229 12189 10241 12223
rect 10275 12220 10287 12223
rect 10870 12220 10876 12232
rect 10275 12192 10876 12220
rect 10275 12189 10287 12192
rect 10229 12183 10287 12189
rect 10870 12180 10876 12192
rect 10928 12180 10934 12232
rect 13354 12220 13360 12232
rect 13315 12192 13360 12220
rect 13354 12180 13360 12192
rect 13412 12180 13418 12232
rect 13740 12220 13768 12251
rect 14366 12248 14372 12260
rect 14424 12248 14430 12300
rect 15657 12291 15715 12297
rect 15657 12257 15669 12291
rect 15703 12288 15715 12291
rect 15948 12288 15976 12328
rect 16390 12316 16396 12328
rect 16448 12356 16454 12368
rect 16448 12328 17908 12356
rect 16448 12316 16454 12328
rect 15703 12260 15976 12288
rect 16209 12291 16267 12297
rect 15703 12257 15715 12260
rect 15657 12251 15715 12257
rect 16209 12257 16221 12291
rect 16255 12257 16267 12291
rect 16209 12251 16267 12257
rect 16114 12220 16120 12232
rect 13740 12192 16120 12220
rect 16114 12180 16120 12192
rect 16172 12180 16178 12232
rect 7156 12124 8524 12152
rect 7156 12112 7162 12124
rect 2406 12044 2412 12096
rect 2464 12084 2470 12096
rect 2777 12087 2835 12093
rect 2777 12084 2789 12087
rect 2464 12056 2789 12084
rect 2464 12044 2470 12056
rect 2777 12053 2789 12056
rect 2823 12053 2835 12087
rect 8386 12084 8392 12096
rect 8347 12056 8392 12084
rect 2777 12047 2835 12053
rect 8386 12044 8392 12056
rect 8444 12044 8450 12096
rect 8496 12084 8524 12124
rect 14734 12112 14740 12164
rect 14792 12152 14798 12164
rect 16224 12152 16252 12251
rect 17494 12248 17500 12300
rect 17552 12288 17558 12300
rect 17681 12291 17739 12297
rect 17681 12288 17693 12291
rect 17552 12260 17693 12288
rect 17552 12248 17558 12260
rect 17681 12257 17693 12260
rect 17727 12257 17739 12291
rect 17681 12251 17739 12257
rect 16485 12223 16543 12229
rect 16485 12189 16497 12223
rect 16531 12220 16543 12223
rect 17037 12223 17095 12229
rect 17037 12220 17049 12223
rect 16531 12192 17049 12220
rect 16531 12189 16543 12192
rect 16485 12183 16543 12189
rect 17037 12189 17049 12192
rect 17083 12189 17095 12223
rect 17037 12183 17095 12189
rect 17773 12223 17831 12229
rect 17773 12189 17785 12223
rect 17819 12189 17831 12223
rect 17880 12220 17908 12328
rect 18046 12288 18052 12300
rect 18007 12260 18052 12288
rect 18046 12248 18052 12260
rect 18104 12248 18110 12300
rect 18233 12291 18291 12297
rect 18233 12257 18245 12291
rect 18279 12288 18291 12291
rect 18524 12288 18552 12396
rect 18966 12384 18972 12396
rect 19024 12424 19030 12436
rect 20717 12427 20775 12433
rect 19024 12396 19840 12424
rect 19024 12384 19030 12396
rect 19426 12316 19432 12368
rect 19484 12316 19490 12368
rect 18279 12260 18552 12288
rect 18279 12257 18291 12260
rect 18233 12251 18291 12257
rect 18598 12248 18604 12300
rect 18656 12288 18662 12300
rect 18874 12288 18880 12300
rect 18656 12260 18880 12288
rect 18656 12248 18662 12260
rect 18874 12248 18880 12260
rect 18932 12248 18938 12300
rect 19334 12288 19340 12300
rect 19295 12260 19340 12288
rect 19334 12248 19340 12260
rect 19392 12248 19398 12300
rect 19444 12288 19472 12316
rect 19702 12288 19708 12300
rect 19444 12260 19708 12288
rect 19702 12248 19708 12260
rect 19760 12248 19766 12300
rect 19812 12297 19840 12396
rect 20717 12393 20729 12427
rect 20763 12424 20775 12427
rect 23201 12427 23259 12433
rect 23201 12424 23213 12427
rect 20763 12396 23213 12424
rect 20763 12393 20775 12396
rect 20717 12387 20775 12393
rect 23201 12393 23213 12396
rect 23247 12424 23259 12427
rect 27246 12424 27252 12436
rect 23247 12396 24716 12424
rect 23247 12393 23259 12396
rect 23201 12387 23259 12393
rect 19797 12291 19855 12297
rect 19797 12257 19809 12291
rect 19843 12257 19855 12291
rect 21174 12288 21180 12300
rect 21135 12260 21180 12288
rect 19797 12251 19855 12257
rect 21174 12248 21180 12260
rect 21232 12248 21238 12300
rect 23017 12291 23075 12297
rect 23017 12257 23029 12291
rect 23063 12288 23075 12291
rect 24026 12288 24032 12300
rect 23063 12260 23888 12288
rect 23987 12260 24032 12288
rect 23063 12257 23075 12260
rect 23017 12251 23075 12257
rect 17880 12192 18920 12220
rect 17773 12183 17831 12189
rect 14792 12124 16252 12152
rect 17788 12152 17816 12183
rect 18598 12152 18604 12164
rect 17788 12124 18604 12152
rect 14792 12112 14798 12124
rect 18598 12112 18604 12124
rect 18656 12112 18662 12164
rect 11054 12084 11060 12096
rect 8496 12056 11060 12084
rect 11054 12044 11060 12056
rect 11112 12044 11118 12096
rect 11330 12084 11336 12096
rect 11291 12056 11336 12084
rect 11330 12044 11336 12056
rect 11388 12044 11394 12096
rect 11606 12044 11612 12096
rect 11664 12084 11670 12096
rect 12161 12087 12219 12093
rect 12161 12084 12173 12087
rect 11664 12056 12173 12084
rect 11664 12044 11670 12056
rect 12161 12053 12173 12056
rect 12207 12084 12219 12087
rect 12250 12084 12256 12096
rect 12207 12056 12256 12084
rect 12207 12053 12219 12056
rect 12161 12047 12219 12053
rect 12250 12044 12256 12056
rect 12308 12044 12314 12096
rect 13170 12044 13176 12096
rect 13228 12084 13234 12096
rect 14553 12087 14611 12093
rect 14553 12084 14565 12087
rect 13228 12056 14565 12084
rect 13228 12044 13234 12056
rect 14553 12053 14565 12056
rect 14599 12084 14611 12087
rect 14642 12084 14648 12096
rect 14599 12056 14648 12084
rect 14599 12053 14611 12056
rect 14553 12047 14611 12053
rect 14642 12044 14648 12056
rect 14700 12044 14706 12096
rect 17310 12044 17316 12096
rect 17368 12084 17374 12096
rect 18785 12087 18843 12093
rect 18785 12084 18797 12087
rect 17368 12056 18797 12084
rect 17368 12044 17374 12056
rect 18785 12053 18797 12056
rect 18831 12053 18843 12087
rect 18892 12084 18920 12192
rect 19058 12180 19064 12232
rect 19116 12220 19122 12232
rect 19245 12223 19303 12229
rect 19245 12220 19257 12223
rect 19116 12192 19257 12220
rect 19116 12180 19122 12192
rect 19245 12189 19257 12192
rect 19291 12189 19303 12223
rect 20898 12220 20904 12232
rect 20859 12192 20904 12220
rect 19245 12183 19303 12189
rect 20898 12180 20904 12192
rect 20956 12180 20962 12232
rect 23750 12220 23756 12232
rect 23711 12192 23756 12220
rect 23750 12180 23756 12192
rect 23808 12180 23814 12232
rect 23860 12220 23888 12260
rect 24026 12248 24032 12260
rect 24084 12248 24090 12300
rect 24688 12288 24716 12396
rect 27080 12396 27252 12424
rect 27080 12365 27108 12396
rect 27246 12384 27252 12396
rect 27304 12384 27310 12436
rect 27614 12384 27620 12436
rect 27672 12424 27678 12436
rect 27982 12424 27988 12436
rect 27672 12396 27988 12424
rect 27672 12384 27678 12396
rect 27982 12384 27988 12396
rect 28040 12384 28046 12436
rect 29638 12384 29644 12436
rect 29696 12424 29702 12436
rect 30006 12424 30012 12436
rect 29696 12396 30012 12424
rect 29696 12384 29702 12396
rect 30006 12384 30012 12396
rect 30064 12384 30070 12436
rect 27065 12359 27123 12365
rect 27065 12325 27077 12359
rect 27111 12325 27123 12359
rect 27065 12319 27123 12325
rect 27433 12359 27491 12365
rect 27433 12325 27445 12359
rect 27479 12356 27491 12359
rect 28534 12356 28540 12368
rect 27479 12328 28540 12356
rect 27479 12325 27491 12328
rect 27433 12319 27491 12325
rect 28534 12316 28540 12328
rect 28592 12316 28598 12368
rect 29365 12359 29423 12365
rect 29365 12325 29377 12359
rect 29411 12356 29423 12359
rect 29454 12356 29460 12368
rect 29411 12328 29460 12356
rect 29411 12325 29423 12328
rect 29365 12319 29423 12325
rect 29454 12316 29460 12328
rect 29512 12316 29518 12368
rect 32214 12356 32220 12368
rect 29840 12328 32220 12356
rect 27249 12291 27307 12297
rect 27249 12288 27261 12291
rect 24688 12260 27261 12288
rect 27249 12257 27261 12260
rect 27295 12257 27307 12291
rect 27249 12251 27307 12257
rect 27341 12291 27399 12297
rect 27341 12257 27353 12291
rect 27387 12288 27399 12291
rect 27614 12288 27620 12300
rect 27387 12260 27620 12288
rect 27387 12257 27399 12260
rect 27341 12251 27399 12257
rect 27614 12248 27620 12260
rect 27672 12288 27678 12300
rect 27890 12288 27896 12300
rect 27672 12260 27896 12288
rect 27672 12248 27678 12260
rect 27890 12248 27896 12260
rect 27948 12248 27954 12300
rect 28810 12288 28816 12300
rect 28771 12260 28816 12288
rect 28810 12248 28816 12260
rect 28868 12248 28874 12300
rect 29086 12288 29092 12300
rect 29047 12260 29092 12288
rect 29086 12248 29092 12260
rect 29144 12248 29150 12300
rect 29840 12297 29868 12328
rect 32214 12316 32220 12328
rect 32272 12316 32278 12368
rect 32306 12316 32312 12368
rect 32364 12356 32370 12368
rect 32490 12356 32496 12368
rect 32364 12328 32409 12356
rect 32451 12328 32496 12356
rect 32364 12316 32370 12328
rect 32490 12316 32496 12328
rect 32548 12316 32554 12368
rect 29825 12291 29883 12297
rect 29825 12257 29837 12291
rect 29871 12257 29883 12291
rect 29825 12251 29883 12257
rect 30282 12248 30288 12300
rect 30340 12288 30346 12300
rect 30837 12291 30895 12297
rect 30837 12288 30849 12291
rect 30340 12260 30849 12288
rect 30340 12248 30346 12260
rect 30837 12257 30849 12260
rect 30883 12257 30895 12291
rect 30837 12251 30895 12257
rect 31294 12248 31300 12300
rect 31352 12288 31358 12300
rect 32398 12288 32404 12300
rect 31352 12260 31397 12288
rect 32359 12260 32404 12288
rect 31352 12248 31358 12260
rect 32398 12248 32404 12260
rect 32456 12248 32462 12300
rect 33962 12288 33968 12300
rect 33923 12260 33968 12288
rect 33962 12248 33968 12260
rect 34020 12248 34026 12300
rect 34333 12291 34391 12297
rect 34333 12257 34345 12291
rect 34379 12288 34391 12291
rect 34606 12288 34612 12300
rect 34379 12260 34612 12288
rect 34379 12257 34391 12260
rect 34333 12251 34391 12257
rect 34606 12248 34612 12260
rect 34664 12248 34670 12300
rect 36817 12291 36875 12297
rect 36817 12257 36829 12291
rect 36863 12288 36875 12291
rect 37734 12288 37740 12300
rect 36863 12260 37740 12288
rect 36863 12257 36875 12260
rect 36817 12251 36875 12257
rect 37734 12248 37740 12260
rect 37792 12248 37798 12300
rect 25498 12220 25504 12232
rect 23860 12192 25504 12220
rect 25498 12180 25504 12192
rect 25556 12180 25562 12232
rect 27798 12220 27804 12232
rect 27759 12192 27804 12220
rect 27798 12180 27804 12192
rect 27856 12180 27862 12232
rect 28353 12223 28411 12229
rect 28353 12189 28365 12223
rect 28399 12189 28411 12223
rect 30561 12223 30619 12229
rect 30561 12220 30573 12223
rect 28353 12183 28411 12189
rect 28460 12192 30573 12220
rect 28368 12152 28396 12183
rect 24688 12124 28396 12152
rect 20717 12087 20775 12093
rect 20717 12084 20729 12087
rect 18892 12056 20729 12084
rect 18785 12047 18843 12053
rect 20717 12053 20729 12056
rect 20763 12053 20775 12087
rect 20717 12047 20775 12053
rect 22094 12044 22100 12096
rect 22152 12084 22158 12096
rect 22281 12087 22339 12093
rect 22281 12084 22293 12087
rect 22152 12056 22293 12084
rect 22152 12044 22158 12056
rect 22281 12053 22293 12056
rect 22327 12053 22339 12087
rect 22281 12047 22339 12053
rect 23658 12044 23664 12096
rect 23716 12084 23722 12096
rect 24688 12084 24716 12124
rect 23716 12056 24716 12084
rect 25317 12087 25375 12093
rect 23716 12044 23722 12056
rect 25317 12053 25329 12087
rect 25363 12084 25375 12087
rect 25590 12084 25596 12096
rect 25363 12056 25596 12084
rect 25363 12053 25375 12056
rect 25317 12047 25375 12053
rect 25590 12044 25596 12056
rect 25648 12044 25654 12096
rect 27246 12044 27252 12096
rect 27304 12084 27310 12096
rect 28166 12084 28172 12096
rect 27304 12056 28172 12084
rect 27304 12044 27310 12056
rect 28166 12044 28172 12056
rect 28224 12084 28230 12096
rect 28460 12084 28488 12192
rect 30561 12189 30573 12192
rect 30607 12220 30619 12223
rect 31202 12220 31208 12232
rect 30607 12192 31208 12220
rect 30607 12189 30619 12192
rect 30561 12183 30619 12189
rect 31202 12180 31208 12192
rect 31260 12180 31266 12232
rect 31573 12223 31631 12229
rect 31573 12189 31585 12223
rect 31619 12220 31631 12223
rect 31754 12220 31760 12232
rect 31619 12192 31760 12220
rect 31619 12189 31631 12192
rect 31573 12183 31631 12189
rect 31754 12180 31760 12192
rect 31812 12180 31818 12232
rect 32122 12220 32128 12232
rect 32083 12192 32128 12220
rect 32122 12180 32128 12192
rect 32180 12180 32186 12232
rect 32858 12220 32864 12232
rect 32819 12192 32864 12220
rect 32858 12180 32864 12192
rect 32916 12180 32922 12232
rect 33502 12220 33508 12232
rect 33463 12192 33508 12220
rect 33502 12180 33508 12192
rect 33560 12180 33566 12232
rect 35161 12223 35219 12229
rect 35161 12189 35173 12223
rect 35207 12189 35219 12223
rect 35434 12220 35440 12232
rect 35395 12192 35440 12220
rect 35161 12183 35219 12189
rect 28718 12112 28724 12164
rect 28776 12152 28782 12164
rect 30742 12152 30748 12164
rect 28776 12124 30748 12152
rect 28776 12112 28782 12124
rect 30742 12112 30748 12124
rect 30800 12112 30806 12164
rect 34238 12152 34244 12164
rect 34199 12124 34244 12152
rect 34238 12112 34244 12124
rect 34296 12112 34302 12164
rect 28224 12056 28488 12084
rect 29917 12087 29975 12093
rect 28224 12044 28230 12056
rect 29917 12053 29929 12087
rect 29963 12084 29975 12087
rect 30006 12084 30012 12096
rect 29963 12056 30012 12084
rect 29963 12053 29975 12056
rect 29917 12047 29975 12053
rect 30006 12044 30012 12056
rect 30064 12084 30070 12096
rect 30282 12084 30288 12096
rect 30064 12056 30288 12084
rect 30064 12044 30070 12056
rect 30282 12044 30288 12056
rect 30340 12044 30346 12096
rect 35176 12084 35204 12183
rect 35434 12180 35440 12192
rect 35492 12180 35498 12232
rect 37274 12180 37280 12232
rect 37332 12220 37338 12232
rect 37829 12223 37887 12229
rect 37829 12220 37841 12223
rect 37332 12192 37841 12220
rect 37332 12180 37338 12192
rect 37829 12189 37841 12192
rect 37875 12189 37887 12223
rect 37829 12183 37887 12189
rect 35342 12084 35348 12096
rect 35176 12056 35348 12084
rect 35342 12044 35348 12056
rect 35400 12044 35406 12096
rect 1104 11994 38824 12016
rect 1104 11942 4246 11994
rect 4298 11942 4310 11994
rect 4362 11942 4374 11994
rect 4426 11942 4438 11994
rect 4490 11942 34966 11994
rect 35018 11942 35030 11994
rect 35082 11942 35094 11994
rect 35146 11942 35158 11994
rect 35210 11942 38824 11994
rect 1104 11920 38824 11942
rect 4062 11880 4068 11892
rect 2056 11852 4068 11880
rect 1762 11676 1768 11688
rect 1723 11648 1768 11676
rect 1762 11636 1768 11648
rect 1820 11636 1826 11688
rect 2056 11685 2084 11852
rect 4062 11840 4068 11852
rect 4120 11840 4126 11892
rect 4249 11883 4307 11889
rect 4249 11849 4261 11883
rect 4295 11880 4307 11883
rect 4614 11880 4620 11892
rect 4295 11852 4620 11880
rect 4295 11849 4307 11852
rect 4249 11843 4307 11849
rect 4614 11840 4620 11852
rect 4672 11880 4678 11892
rect 5258 11880 5264 11892
rect 4672 11852 5264 11880
rect 4672 11840 4678 11852
rect 5258 11840 5264 11852
rect 5316 11840 5322 11892
rect 6270 11840 6276 11892
rect 6328 11880 6334 11892
rect 8113 11883 8171 11889
rect 6328 11852 7052 11880
rect 6328 11840 6334 11852
rect 5810 11772 5816 11824
rect 5868 11812 5874 11824
rect 6917 11815 6975 11821
rect 6917 11812 6929 11815
rect 5868 11784 6929 11812
rect 5868 11772 5874 11784
rect 6917 11781 6929 11784
rect 6963 11781 6975 11815
rect 7024 11812 7052 11852
rect 8113 11849 8125 11883
rect 8159 11880 8171 11883
rect 8294 11880 8300 11892
rect 8159 11852 8300 11880
rect 8159 11849 8171 11852
rect 8113 11843 8171 11849
rect 8294 11840 8300 11852
rect 8352 11840 8358 11892
rect 14734 11880 14740 11892
rect 12820 11852 14740 11880
rect 10686 11812 10692 11824
rect 7024 11784 10692 11812
rect 6917 11775 6975 11781
rect 10686 11772 10692 11784
rect 10744 11772 10750 11824
rect 10870 11812 10876 11824
rect 10831 11784 10876 11812
rect 10870 11772 10876 11784
rect 10928 11772 10934 11824
rect 12820 11821 12848 11852
rect 14734 11840 14740 11852
rect 14792 11840 14798 11892
rect 16132 11852 18184 11880
rect 12805 11815 12863 11821
rect 10980 11784 11284 11812
rect 2958 11744 2964 11756
rect 2919 11716 2964 11744
rect 2958 11704 2964 11716
rect 3016 11704 3022 11756
rect 6270 11744 6276 11756
rect 5276 11716 6276 11744
rect 5276 11688 5304 11716
rect 6270 11704 6276 11716
rect 6328 11704 6334 11756
rect 6454 11704 6460 11756
rect 6512 11744 6518 11756
rect 8938 11744 8944 11756
rect 6512 11716 8340 11744
rect 8899 11716 8944 11744
rect 6512 11704 6518 11716
rect 2041 11679 2099 11685
rect 2041 11645 2053 11679
rect 2087 11645 2099 11679
rect 2041 11639 2099 11645
rect 2685 11679 2743 11685
rect 2685 11645 2697 11679
rect 2731 11645 2743 11679
rect 4798 11676 4804 11688
rect 4759 11648 4804 11676
rect 2685 11639 2743 11645
rect 1854 11568 1860 11620
rect 1912 11608 1918 11620
rect 2700 11608 2728 11639
rect 4798 11636 4804 11648
rect 4856 11636 4862 11688
rect 5258 11676 5264 11688
rect 5171 11648 5264 11676
rect 5258 11636 5264 11648
rect 5316 11636 5322 11688
rect 5350 11636 5356 11688
rect 5408 11676 5414 11688
rect 5537 11679 5595 11685
rect 5537 11676 5549 11679
rect 5408 11648 5549 11676
rect 5408 11636 5414 11648
rect 5537 11645 5549 11648
rect 5583 11645 5595 11679
rect 7098 11676 7104 11688
rect 7059 11648 7104 11676
rect 5537 11639 5595 11645
rect 7098 11636 7104 11648
rect 7156 11636 7162 11688
rect 7374 11676 7380 11688
rect 7335 11648 7380 11676
rect 7374 11636 7380 11648
rect 7432 11636 7438 11688
rect 8312 11685 8340 11716
rect 8938 11704 8944 11716
rect 8996 11704 9002 11756
rect 9858 11704 9864 11756
rect 9916 11744 9922 11756
rect 10980 11744 11008 11784
rect 9916 11716 11008 11744
rect 9916 11704 9922 11716
rect 11146 11704 11152 11756
rect 11204 11704 11210 11756
rect 11256 11744 11284 11784
rect 12805 11781 12817 11815
rect 12851 11781 12863 11815
rect 15378 11812 15384 11824
rect 12805 11775 12863 11781
rect 14292 11784 15384 11812
rect 11256 11716 13216 11744
rect 8297 11679 8355 11685
rect 8297 11645 8309 11679
rect 8343 11645 8355 11679
rect 8297 11639 8355 11645
rect 8386 11636 8392 11688
rect 8444 11676 8450 11688
rect 8444 11648 8489 11676
rect 8444 11636 8450 11648
rect 8570 11636 8576 11688
rect 8628 11676 8634 11688
rect 8757 11679 8815 11685
rect 8757 11676 8769 11679
rect 8628 11648 8769 11676
rect 8628 11636 8634 11648
rect 8757 11645 8769 11648
rect 8803 11645 8815 11679
rect 9122 11676 9128 11688
rect 9083 11648 9128 11676
rect 8757 11639 8815 11645
rect 9122 11636 9128 11648
rect 9180 11636 9186 11688
rect 9950 11636 9956 11688
rect 10008 11676 10014 11688
rect 10045 11679 10103 11685
rect 10045 11676 10057 11679
rect 10008 11648 10057 11676
rect 10008 11636 10014 11648
rect 10045 11645 10057 11648
rect 10091 11676 10103 11679
rect 10226 11676 10232 11688
rect 10091 11648 10232 11676
rect 10091 11645 10103 11648
rect 10045 11639 10103 11645
rect 10226 11636 10232 11648
rect 10284 11636 10290 11688
rect 10318 11636 10324 11688
rect 10376 11676 10382 11688
rect 10413 11679 10471 11685
rect 10413 11676 10425 11679
rect 10376 11648 10425 11676
rect 10376 11636 10382 11648
rect 10413 11645 10425 11648
rect 10459 11645 10471 11679
rect 10413 11639 10471 11645
rect 10965 11679 11023 11685
rect 10965 11645 10977 11679
rect 11011 11676 11023 11679
rect 11164 11676 11192 11704
rect 11011 11648 11192 11676
rect 11609 11679 11667 11685
rect 11011 11645 11023 11648
rect 10965 11639 11023 11645
rect 11609 11645 11621 11679
rect 11655 11676 11667 11679
rect 12986 11676 12992 11688
rect 11655 11648 12992 11676
rect 11655 11645 11667 11648
rect 11609 11639 11667 11645
rect 12986 11636 12992 11648
rect 13044 11636 13050 11688
rect 13188 11685 13216 11716
rect 13173 11679 13231 11685
rect 13173 11645 13185 11679
rect 13219 11645 13231 11679
rect 13354 11676 13360 11688
rect 13315 11648 13360 11676
rect 13173 11639 13231 11645
rect 13354 11636 13360 11648
rect 13412 11636 13418 11688
rect 14292 11685 14320 11784
rect 15378 11772 15384 11784
rect 15436 11772 15442 11824
rect 15562 11772 15568 11824
rect 15620 11812 15626 11824
rect 16132 11812 16160 11852
rect 15620 11784 16160 11812
rect 16577 11815 16635 11821
rect 15620 11772 15626 11784
rect 16577 11781 16589 11815
rect 16623 11812 16635 11815
rect 17402 11812 17408 11824
rect 16623 11784 17408 11812
rect 16623 11781 16635 11784
rect 16577 11775 16635 11781
rect 17402 11772 17408 11784
rect 17460 11772 17466 11824
rect 14458 11744 14464 11756
rect 14419 11716 14464 11744
rect 14458 11704 14464 11716
rect 14516 11704 14522 11756
rect 17310 11744 17316 11756
rect 17271 11716 17316 11744
rect 17310 11704 17316 11716
rect 17368 11704 17374 11756
rect 14277 11679 14335 11685
rect 14277 11645 14289 11679
rect 14323 11645 14335 11679
rect 14642 11676 14648 11688
rect 14603 11648 14648 11676
rect 14277 11639 14335 11645
rect 14642 11636 14648 11648
rect 14700 11636 14706 11688
rect 15105 11679 15163 11685
rect 15105 11645 15117 11679
rect 15151 11676 15163 11679
rect 15378 11676 15384 11688
rect 15151 11648 15384 11676
rect 15151 11645 15163 11648
rect 15105 11639 15163 11645
rect 15378 11636 15384 11648
rect 15436 11636 15442 11688
rect 15470 11636 15476 11688
rect 15528 11676 15534 11688
rect 15930 11676 15936 11688
rect 15528 11648 15936 11676
rect 15528 11636 15534 11648
rect 15930 11636 15936 11648
rect 15988 11636 15994 11688
rect 16390 11676 16396 11688
rect 16351 11648 16396 11676
rect 16390 11636 16396 11648
rect 16448 11636 16454 11688
rect 16853 11679 16911 11685
rect 16853 11645 16865 11679
rect 16899 11645 16911 11679
rect 18046 11676 18052 11688
rect 18007 11648 18052 11676
rect 16853 11639 16911 11645
rect 1912 11580 2728 11608
rect 5997 11611 6055 11617
rect 1912 11568 1918 11580
rect 5997 11577 6009 11611
rect 6043 11608 6055 11611
rect 6043 11580 12204 11608
rect 6043 11577 6055 11580
rect 5997 11571 6055 11577
rect 1581 11543 1639 11549
rect 1581 11509 1593 11543
rect 1627 11540 1639 11543
rect 1670 11540 1676 11552
rect 1627 11512 1676 11540
rect 1627 11509 1639 11512
rect 1581 11503 1639 11509
rect 1670 11500 1676 11512
rect 1728 11500 1734 11552
rect 4890 11500 4896 11552
rect 4948 11540 4954 11552
rect 8110 11540 8116 11552
rect 4948 11512 8116 11540
rect 4948 11500 4954 11512
rect 8110 11500 8116 11512
rect 8168 11500 8174 11552
rect 10134 11500 10140 11552
rect 10192 11540 10198 11552
rect 11793 11543 11851 11549
rect 11793 11540 11805 11543
rect 10192 11512 11805 11540
rect 10192 11500 10198 11512
rect 11793 11509 11805 11512
rect 11839 11509 11851 11543
rect 12176 11540 12204 11580
rect 12894 11568 12900 11620
rect 12952 11608 12958 11620
rect 16868 11608 16896 11639
rect 18046 11636 18052 11648
rect 18104 11636 18110 11688
rect 12952 11580 16896 11608
rect 18156 11608 18184 11852
rect 18598 11840 18604 11892
rect 18656 11880 18662 11892
rect 18877 11883 18935 11889
rect 18877 11880 18889 11883
rect 18656 11852 18889 11880
rect 18656 11840 18662 11852
rect 18877 11849 18889 11852
rect 18923 11880 18935 11883
rect 19058 11880 19064 11892
rect 18923 11852 19064 11880
rect 18923 11849 18935 11852
rect 18877 11843 18935 11849
rect 19058 11840 19064 11852
rect 19116 11840 19122 11892
rect 19702 11840 19708 11892
rect 19760 11880 19766 11892
rect 20901 11883 20959 11889
rect 20901 11880 20913 11883
rect 19760 11852 20913 11880
rect 19760 11840 19766 11852
rect 20901 11849 20913 11852
rect 20947 11849 20959 11883
rect 20901 11843 20959 11849
rect 24210 11840 24216 11892
rect 24268 11880 24274 11892
rect 27706 11880 27712 11892
rect 24268 11852 27712 11880
rect 24268 11840 24274 11852
rect 27706 11840 27712 11852
rect 27764 11840 27770 11892
rect 27982 11840 27988 11892
rect 28040 11880 28046 11892
rect 29822 11880 29828 11892
rect 28040 11852 29828 11880
rect 28040 11840 28046 11852
rect 29822 11840 29828 11852
rect 29880 11840 29886 11892
rect 30116 11852 31248 11880
rect 25498 11812 25504 11824
rect 24228 11784 25504 11812
rect 19797 11747 19855 11753
rect 19797 11713 19809 11747
rect 19843 11744 19855 11747
rect 19886 11744 19892 11756
rect 19843 11716 19892 11744
rect 19843 11713 19855 11716
rect 19797 11707 19855 11713
rect 19886 11704 19892 11716
rect 19944 11704 19950 11756
rect 21266 11704 21272 11756
rect 21324 11744 21330 11756
rect 22005 11747 22063 11753
rect 22005 11744 22017 11747
rect 21324 11716 22017 11744
rect 21324 11704 21330 11716
rect 22005 11713 22017 11716
rect 22051 11713 22063 11747
rect 22005 11707 22063 11713
rect 18782 11676 18788 11688
rect 18743 11648 18788 11676
rect 18782 11636 18788 11648
rect 18840 11636 18846 11688
rect 19521 11679 19579 11685
rect 19521 11645 19533 11679
rect 19567 11676 19579 11679
rect 20254 11676 20260 11688
rect 19567 11648 20260 11676
rect 19567 11645 19579 11648
rect 19521 11639 19579 11645
rect 20254 11636 20260 11648
rect 20312 11636 20318 11688
rect 20898 11636 20904 11688
rect 20956 11676 20962 11688
rect 21450 11676 21456 11688
rect 20956 11648 21456 11676
rect 20956 11636 20962 11648
rect 21450 11636 21456 11648
rect 21508 11636 21514 11688
rect 22094 11636 22100 11688
rect 22152 11676 22158 11688
rect 22152 11648 22197 11676
rect 22152 11636 22158 11648
rect 22462 11636 22468 11688
rect 22520 11676 22526 11688
rect 24121 11679 24179 11685
rect 24121 11676 24133 11679
rect 22520 11648 24133 11676
rect 22520 11636 22526 11648
rect 24121 11645 24133 11648
rect 24167 11676 24179 11679
rect 24228 11676 24256 11784
rect 25498 11772 25504 11784
rect 25556 11772 25562 11824
rect 30116 11812 30144 11852
rect 29104 11784 30144 11812
rect 24581 11747 24639 11753
rect 24581 11713 24593 11747
rect 24627 11744 24639 11747
rect 24670 11744 24676 11756
rect 24627 11716 24676 11744
rect 24627 11713 24639 11716
rect 24581 11707 24639 11713
rect 24670 11704 24676 11716
rect 24728 11704 24734 11756
rect 25225 11747 25283 11753
rect 25225 11713 25237 11747
rect 25271 11744 25283 11747
rect 26142 11744 26148 11756
rect 25271 11716 26148 11744
rect 25271 11713 25283 11716
rect 25225 11707 25283 11713
rect 26142 11704 26148 11716
rect 26200 11744 26206 11756
rect 26200 11716 27384 11744
rect 26200 11704 26206 11716
rect 24167 11648 24256 11676
rect 24397 11679 24455 11685
rect 24167 11645 24179 11648
rect 24121 11639 24179 11645
rect 24397 11645 24409 11679
rect 24443 11676 24455 11679
rect 24443 11648 25636 11676
rect 24443 11645 24455 11648
rect 24397 11639 24455 11645
rect 25608 11620 25636 11648
rect 26418 11636 26424 11688
rect 26476 11676 26482 11688
rect 26697 11679 26755 11685
rect 26697 11676 26709 11679
rect 26476 11648 26709 11676
rect 26476 11636 26482 11648
rect 26697 11645 26709 11648
rect 26743 11676 26755 11679
rect 26970 11676 26976 11688
rect 26743 11648 26976 11676
rect 26743 11645 26755 11648
rect 26697 11639 26755 11645
rect 26970 11636 26976 11648
rect 27028 11636 27034 11688
rect 27157 11679 27215 11685
rect 27157 11645 27169 11679
rect 27203 11676 27215 11679
rect 27246 11676 27252 11688
rect 27203 11648 27252 11676
rect 27203 11645 27215 11648
rect 27157 11639 27215 11645
rect 27246 11636 27252 11648
rect 27304 11636 27310 11688
rect 27356 11685 27384 11716
rect 27614 11704 27620 11756
rect 27672 11744 27678 11756
rect 27672 11716 28120 11744
rect 27672 11704 27678 11716
rect 27341 11679 27399 11685
rect 27341 11645 27353 11679
rect 27387 11645 27399 11679
rect 27706 11676 27712 11688
rect 27667 11648 27712 11676
rect 27341 11639 27399 11645
rect 27706 11636 27712 11648
rect 27764 11636 27770 11688
rect 28092 11685 28120 11716
rect 29104 11685 29132 11784
rect 30190 11772 30196 11824
rect 30248 11772 30254 11824
rect 31220 11812 31248 11852
rect 31294 11840 31300 11892
rect 31352 11880 31358 11892
rect 37458 11880 37464 11892
rect 31352 11852 37464 11880
rect 31352 11840 31358 11852
rect 37458 11840 37464 11852
rect 37516 11840 37522 11892
rect 37826 11880 37832 11892
rect 37787 11852 37832 11880
rect 37826 11840 37832 11852
rect 37884 11840 37890 11892
rect 31938 11812 31944 11824
rect 31220 11784 31944 11812
rect 31938 11772 31944 11784
rect 31996 11772 32002 11824
rect 32769 11815 32827 11821
rect 32769 11812 32781 11815
rect 32048 11784 32781 11812
rect 30208 11744 30236 11772
rect 32048 11744 32076 11784
rect 32769 11781 32781 11784
rect 32815 11781 32827 11815
rect 32769 11775 32827 11781
rect 33137 11815 33195 11821
rect 33137 11781 33149 11815
rect 33183 11812 33195 11815
rect 33962 11812 33968 11824
rect 33183 11784 33968 11812
rect 33183 11781 33195 11784
rect 33137 11775 33195 11781
rect 33962 11772 33968 11784
rect 34020 11772 34026 11824
rect 29840 11716 32076 11744
rect 28077 11679 28135 11685
rect 28077 11645 28089 11679
rect 28123 11645 28135 11679
rect 28077 11639 28135 11645
rect 29089 11679 29147 11685
rect 29089 11645 29101 11679
rect 29135 11645 29147 11679
rect 29089 11639 29147 11645
rect 29178 11636 29184 11688
rect 29236 11636 29242 11688
rect 29840 11685 29868 11716
rect 32214 11704 32220 11756
rect 32272 11744 32278 11756
rect 33778 11744 33784 11756
rect 32272 11716 33784 11744
rect 32272 11704 32278 11716
rect 33778 11704 33784 11716
rect 33836 11704 33842 11756
rect 34514 11704 34520 11756
rect 34572 11744 34578 11756
rect 34790 11744 34796 11756
rect 34572 11716 34796 11744
rect 34572 11704 34578 11716
rect 34790 11704 34796 11716
rect 34848 11744 34854 11756
rect 35713 11747 35771 11753
rect 35713 11744 35725 11747
rect 34848 11716 35725 11744
rect 34848 11704 34854 11716
rect 35713 11713 35725 11716
rect 35759 11713 35771 11747
rect 35713 11707 35771 11713
rect 29825 11679 29883 11685
rect 29825 11645 29837 11679
rect 29871 11645 29883 11679
rect 29825 11639 29883 11645
rect 30009 11679 30067 11685
rect 30009 11645 30021 11679
rect 30055 11645 30067 11679
rect 30190 11676 30196 11688
rect 30151 11648 30196 11676
rect 30009 11639 30067 11645
rect 22554 11608 22560 11620
rect 18156 11580 19564 11608
rect 22515 11580 22560 11608
rect 12952 11568 12958 11580
rect 14366 11540 14372 11552
rect 12176 11512 14372 11540
rect 11793 11503 11851 11509
rect 14366 11500 14372 11512
rect 14424 11500 14430 11552
rect 14642 11500 14648 11552
rect 14700 11540 14706 11552
rect 18233 11543 18291 11549
rect 18233 11540 18245 11543
rect 14700 11512 18245 11540
rect 14700 11500 14706 11512
rect 18233 11509 18245 11512
rect 18279 11540 18291 11543
rect 19426 11540 19432 11552
rect 18279 11512 19432 11540
rect 18279 11509 18291 11512
rect 18233 11503 18291 11509
rect 19426 11500 19432 11512
rect 19484 11500 19490 11552
rect 19536 11540 19564 11580
rect 22554 11568 22560 11580
rect 22612 11568 22618 11620
rect 25314 11608 25320 11620
rect 25240 11580 25320 11608
rect 20070 11540 20076 11552
rect 19536 11512 20076 11540
rect 20070 11500 20076 11512
rect 20128 11500 20134 11552
rect 22278 11500 22284 11552
rect 22336 11540 22342 11552
rect 25240 11540 25268 11580
rect 25314 11568 25320 11580
rect 25372 11568 25378 11620
rect 25590 11608 25596 11620
rect 25551 11580 25596 11608
rect 25590 11568 25596 11580
rect 25648 11568 25654 11620
rect 25958 11608 25964 11620
rect 25919 11580 25964 11608
rect 25958 11568 25964 11580
rect 26016 11568 26022 11620
rect 26789 11611 26847 11617
rect 26789 11577 26801 11611
rect 26835 11608 26847 11611
rect 29196 11608 29224 11636
rect 26835 11580 29224 11608
rect 29273 11611 29331 11617
rect 26835 11577 26847 11580
rect 26789 11571 26847 11577
rect 29273 11577 29285 11611
rect 29319 11608 29331 11611
rect 29730 11608 29736 11620
rect 29319 11580 29736 11608
rect 29319 11577 29331 11580
rect 29273 11571 29331 11577
rect 29730 11568 29736 11580
rect 29788 11568 29794 11620
rect 30024 11608 30052 11639
rect 30190 11636 30196 11648
rect 30248 11636 30254 11688
rect 30377 11679 30435 11685
rect 30377 11645 30389 11679
rect 30423 11645 30435 11679
rect 30377 11639 30435 11645
rect 29840 11580 30052 11608
rect 30392 11608 30420 11639
rect 30466 11636 30472 11688
rect 30524 11676 30530 11688
rect 30653 11679 30711 11685
rect 30653 11676 30665 11679
rect 30524 11648 30665 11676
rect 30524 11636 30530 11648
rect 30653 11645 30665 11648
rect 30699 11645 30711 11679
rect 31202 11676 31208 11688
rect 31163 11648 31208 11676
rect 30653 11639 30711 11645
rect 31202 11636 31208 11648
rect 31260 11636 31266 11688
rect 31570 11676 31576 11688
rect 31531 11648 31576 11676
rect 31570 11636 31576 11648
rect 31628 11636 31634 11688
rect 31938 11636 31944 11688
rect 31996 11685 32002 11688
rect 31996 11679 32045 11685
rect 31996 11645 31999 11679
rect 32033 11645 32045 11679
rect 32490 11676 32496 11688
rect 31996 11639 32045 11645
rect 32140 11648 32496 11676
rect 31996 11636 32002 11639
rect 31662 11608 31668 11620
rect 30392 11580 31668 11608
rect 29840 11552 29868 11580
rect 31662 11568 31668 11580
rect 31720 11608 31726 11620
rect 32140 11608 32168 11648
rect 32490 11636 32496 11648
rect 32548 11636 32554 11688
rect 32769 11679 32827 11685
rect 32769 11645 32781 11679
rect 32815 11676 32827 11679
rect 32861 11679 32919 11685
rect 32861 11676 32873 11679
rect 32815 11648 32873 11676
rect 32815 11645 32827 11648
rect 32769 11639 32827 11645
rect 32861 11645 32873 11648
rect 32907 11645 32919 11679
rect 32861 11639 32919 11645
rect 33318 11636 33324 11688
rect 33376 11676 33382 11688
rect 33413 11679 33471 11685
rect 33413 11676 33425 11679
rect 33376 11648 33425 11676
rect 33376 11636 33382 11648
rect 33413 11645 33425 11648
rect 33459 11645 33471 11679
rect 33413 11639 33471 11645
rect 34054 11636 34060 11688
rect 34112 11676 34118 11688
rect 34885 11679 34943 11685
rect 34885 11676 34897 11679
rect 34112 11648 34897 11676
rect 34112 11636 34118 11648
rect 34885 11645 34897 11648
rect 34931 11645 34943 11679
rect 34885 11639 34943 11645
rect 35621 11679 35679 11685
rect 35621 11645 35633 11679
rect 35667 11676 35679 11679
rect 35802 11676 35808 11688
rect 35667 11648 35808 11676
rect 35667 11645 35679 11648
rect 35621 11639 35679 11645
rect 35802 11636 35808 11648
rect 35860 11636 35866 11688
rect 36446 11676 36452 11688
rect 36407 11648 36452 11676
rect 36446 11636 36452 11648
rect 36504 11636 36510 11688
rect 36722 11676 36728 11688
rect 36683 11648 36728 11676
rect 36722 11636 36728 11648
rect 36780 11636 36786 11688
rect 31720 11580 32168 11608
rect 32309 11611 32367 11617
rect 31720 11568 31726 11580
rect 32309 11577 32321 11611
rect 32355 11608 32367 11611
rect 32674 11608 32680 11620
rect 32355 11580 32680 11608
rect 32355 11577 32367 11580
rect 32309 11571 32367 11577
rect 32674 11568 32680 11580
rect 32732 11568 32738 11620
rect 25406 11540 25412 11552
rect 22336 11512 25268 11540
rect 25367 11512 25412 11540
rect 22336 11500 22342 11512
rect 25406 11500 25412 11512
rect 25464 11500 25470 11552
rect 25498 11500 25504 11552
rect 25556 11540 25562 11552
rect 28905 11543 28963 11549
rect 25556 11512 25601 11540
rect 25556 11500 25562 11512
rect 28905 11509 28917 11543
rect 28951 11540 28963 11543
rect 28994 11540 29000 11552
rect 28951 11512 29000 11540
rect 28951 11509 28963 11512
rect 28905 11503 28963 11509
rect 28994 11500 29000 11512
rect 29052 11540 29058 11552
rect 29454 11540 29460 11552
rect 29052 11512 29460 11540
rect 29052 11500 29058 11512
rect 29454 11500 29460 11512
rect 29512 11500 29518 11552
rect 29822 11500 29828 11552
rect 29880 11500 29886 11552
rect 33042 11500 33048 11552
rect 33100 11540 33106 11552
rect 34977 11543 35035 11549
rect 34977 11540 34989 11543
rect 33100 11512 34989 11540
rect 33100 11500 33106 11512
rect 34977 11509 34989 11512
rect 35023 11509 35035 11543
rect 34977 11503 35035 11509
rect 1104 11450 38824 11472
rect 1104 11398 19606 11450
rect 19658 11398 19670 11450
rect 19722 11398 19734 11450
rect 19786 11398 19798 11450
rect 19850 11398 38824 11450
rect 1104 11376 38824 11398
rect 5074 11296 5080 11348
rect 5132 11336 5138 11348
rect 5261 11339 5319 11345
rect 5261 11336 5273 11339
rect 5132 11308 5273 11336
rect 5132 11296 5138 11308
rect 5261 11305 5273 11308
rect 5307 11305 5319 11339
rect 7098 11336 7104 11348
rect 5261 11299 5319 11305
rect 5368 11308 7104 11336
rect 5368 11268 5396 11308
rect 7098 11296 7104 11308
rect 7156 11296 7162 11348
rect 7561 11339 7619 11345
rect 7561 11305 7573 11339
rect 7607 11336 7619 11339
rect 7926 11336 7932 11348
rect 7607 11308 7932 11336
rect 7607 11305 7619 11308
rect 7561 11299 7619 11305
rect 7926 11296 7932 11308
rect 7984 11296 7990 11348
rect 8110 11296 8116 11348
rect 8168 11336 8174 11348
rect 11514 11336 11520 11348
rect 8168 11308 10824 11336
rect 8168 11296 8174 11308
rect 6454 11268 6460 11280
rect 4356 11240 5396 11268
rect 5460 11240 6460 11268
rect 2406 11200 2412 11212
rect 2367 11172 2412 11200
rect 2406 11160 2412 11172
rect 2464 11160 2470 11212
rect 4356 11209 4384 11240
rect 4341 11203 4399 11209
rect 4341 11169 4353 11203
rect 4387 11169 4399 11203
rect 4614 11200 4620 11212
rect 4575 11172 4620 11200
rect 4341 11163 4399 11169
rect 4614 11160 4620 11172
rect 4672 11160 4678 11212
rect 5460 11209 5488 11240
rect 6454 11228 6460 11240
rect 6512 11228 6518 11280
rect 10134 11268 10140 11280
rect 8588 11240 10140 11268
rect 5445 11203 5503 11209
rect 5445 11169 5457 11203
rect 5491 11169 5503 11203
rect 5810 11200 5816 11212
rect 5771 11172 5816 11200
rect 5445 11163 5503 11169
rect 5810 11160 5816 11172
rect 5868 11160 5874 11212
rect 6089 11203 6147 11209
rect 6089 11169 6101 11203
rect 6135 11200 6147 11203
rect 6270 11200 6276 11212
rect 6135 11172 6276 11200
rect 6135 11169 6147 11172
rect 6089 11163 6147 11169
rect 6270 11160 6276 11172
rect 6328 11160 6334 11212
rect 6549 11203 6607 11209
rect 6549 11169 6561 11203
rect 6595 11200 6607 11203
rect 6914 11200 6920 11212
rect 6595 11172 6920 11200
rect 6595 11169 6607 11172
rect 6549 11163 6607 11169
rect 6914 11160 6920 11172
rect 6972 11160 6978 11212
rect 7377 11203 7435 11209
rect 7377 11169 7389 11203
rect 7423 11200 7435 11203
rect 7558 11200 7564 11212
rect 7423 11172 7564 11200
rect 7423 11169 7435 11172
rect 7377 11163 7435 11169
rect 7558 11160 7564 11172
rect 7616 11160 7622 11212
rect 8588 11209 8616 11240
rect 10134 11228 10140 11240
rect 10192 11228 10198 11280
rect 8573 11203 8631 11209
rect 8573 11169 8585 11203
rect 8619 11169 8631 11203
rect 8573 11163 8631 11169
rect 8757 11203 8815 11209
rect 8757 11169 8769 11203
rect 8803 11169 8815 11203
rect 8938 11200 8944 11212
rect 8899 11172 8944 11200
rect 8757 11163 8815 11169
rect 2130 11092 2136 11144
rect 2188 11132 2194 11144
rect 2317 11135 2375 11141
rect 2317 11132 2329 11135
rect 2188 11104 2329 11132
rect 2188 11092 2194 11104
rect 2317 11101 2329 11104
rect 2363 11101 2375 11135
rect 2866 11132 2872 11144
rect 2827 11104 2872 11132
rect 2317 11095 2375 11101
rect 2866 11092 2872 11104
rect 2924 11092 2930 11144
rect 4433 11135 4491 11141
rect 4433 11101 4445 11135
rect 4479 11132 4491 11135
rect 4479 11104 4660 11132
rect 4479 11101 4491 11104
rect 4433 11095 4491 11101
rect 4632 11076 4660 11104
rect 6178 11092 6184 11144
rect 6236 11132 6242 11144
rect 8772 11132 8800 11163
rect 8938 11160 8944 11172
rect 8996 11160 9002 11212
rect 10594 11200 10600 11212
rect 10555 11172 10600 11200
rect 10594 11160 10600 11172
rect 10652 11160 10658 11212
rect 10686 11132 10692 11144
rect 6236 11104 8800 11132
rect 10647 11104 10692 11132
rect 6236 11092 6242 11104
rect 10686 11092 10692 11104
rect 10744 11092 10750 11144
rect 10796 11132 10824 11308
rect 11072 11308 11520 11336
rect 10962 11200 10968 11212
rect 10923 11172 10968 11200
rect 10962 11160 10968 11172
rect 11020 11160 11026 11212
rect 11072 11209 11100 11308
rect 11514 11296 11520 11308
rect 11572 11336 11578 11348
rect 14642 11336 14648 11348
rect 11572 11308 14648 11336
rect 11572 11296 11578 11308
rect 14642 11296 14648 11308
rect 14700 11296 14706 11348
rect 15473 11339 15531 11345
rect 15473 11305 15485 11339
rect 15519 11336 15531 11339
rect 16206 11336 16212 11348
rect 15519 11308 16212 11336
rect 15519 11305 15531 11308
rect 15473 11299 15531 11305
rect 16206 11296 16212 11308
rect 16264 11296 16270 11348
rect 18230 11296 18236 11348
rect 18288 11336 18294 11348
rect 19521 11339 19579 11345
rect 19521 11336 19533 11339
rect 18288 11308 19533 11336
rect 18288 11296 18294 11308
rect 19521 11305 19533 11308
rect 19567 11305 19579 11339
rect 22370 11336 22376 11348
rect 19521 11299 19579 11305
rect 19996 11308 22376 11336
rect 12986 11228 12992 11280
rect 13044 11268 13050 11280
rect 14734 11268 14740 11280
rect 13044 11240 14740 11268
rect 13044 11228 13050 11240
rect 11057 11203 11115 11209
rect 11057 11169 11069 11203
rect 11103 11169 11115 11203
rect 11057 11163 11115 11169
rect 12713 11203 12771 11209
rect 12713 11169 12725 11203
rect 12759 11200 12771 11203
rect 12802 11200 12808 11212
rect 12759 11172 12808 11200
rect 12759 11169 12771 11172
rect 12713 11163 12771 11169
rect 12802 11160 12808 11172
rect 12860 11160 12866 11212
rect 13078 11200 13084 11212
rect 13039 11172 13084 11200
rect 13078 11160 13084 11172
rect 13136 11160 13142 11212
rect 14200 11209 14228 11240
rect 14734 11228 14740 11240
rect 14792 11228 14798 11280
rect 17773 11271 17831 11277
rect 17773 11237 17785 11271
rect 17819 11268 17831 11271
rect 17954 11268 17960 11280
rect 17819 11240 17960 11268
rect 17819 11237 17831 11240
rect 17773 11231 17831 11237
rect 17954 11228 17960 11240
rect 18012 11228 18018 11280
rect 14185 11203 14243 11209
rect 14185 11169 14197 11203
rect 14231 11169 14243 11203
rect 14366 11200 14372 11212
rect 14327 11172 14372 11200
rect 14185 11163 14243 11169
rect 14366 11160 14372 11172
rect 14424 11160 14430 11212
rect 14458 11160 14464 11212
rect 14516 11200 14522 11212
rect 14553 11203 14611 11209
rect 14553 11200 14565 11203
rect 14516 11172 14565 11200
rect 14516 11160 14522 11172
rect 14553 11169 14565 11172
rect 14599 11169 14611 11203
rect 14553 11163 14611 11169
rect 15562 11160 15568 11212
rect 15620 11200 15626 11212
rect 16022 11200 16028 11212
rect 15620 11172 15665 11200
rect 15983 11172 16028 11200
rect 15620 11160 15626 11172
rect 16022 11160 16028 11172
rect 16080 11160 16086 11212
rect 17037 11203 17095 11209
rect 17037 11200 17049 11203
rect 16132 11172 17049 11200
rect 12253 11135 12311 11141
rect 12253 11132 12265 11135
rect 10796 11104 12265 11132
rect 12253 11101 12265 11104
rect 12299 11101 12311 11135
rect 12253 11095 12311 11101
rect 15838 11092 15844 11144
rect 15896 11132 15902 11144
rect 16132 11132 16160 11172
rect 17037 11169 17049 11172
rect 17083 11200 17095 11203
rect 18046 11200 18052 11212
rect 17083 11172 18052 11200
rect 17083 11169 17095 11172
rect 17037 11163 17095 11169
rect 18046 11160 18052 11172
rect 18104 11160 18110 11212
rect 18414 11200 18420 11212
rect 18375 11172 18420 11200
rect 18414 11160 18420 11172
rect 18472 11160 18478 11212
rect 18509 11203 18567 11209
rect 18509 11169 18521 11203
rect 18555 11200 18567 11203
rect 18598 11200 18604 11212
rect 18555 11172 18604 11200
rect 18555 11169 18567 11172
rect 18509 11163 18567 11169
rect 18598 11160 18604 11172
rect 18656 11160 18662 11212
rect 18785 11203 18843 11209
rect 18785 11169 18797 11203
rect 18831 11200 18843 11203
rect 19150 11200 19156 11212
rect 18831 11172 19156 11200
rect 18831 11169 18843 11172
rect 18785 11163 18843 11169
rect 19150 11160 19156 11172
rect 19208 11160 19214 11212
rect 19426 11200 19432 11212
rect 19387 11172 19432 11200
rect 19426 11160 19432 11172
rect 19484 11160 19490 11212
rect 19996 11209 20024 11308
rect 22370 11296 22376 11308
rect 22428 11296 22434 11348
rect 22649 11339 22707 11345
rect 22649 11305 22661 11339
rect 22695 11305 22707 11339
rect 22649 11299 22707 11305
rect 23569 11339 23627 11345
rect 23569 11305 23581 11339
rect 23615 11336 23627 11339
rect 24210 11336 24216 11348
rect 23615 11308 24216 11336
rect 23615 11305 23627 11308
rect 23569 11299 23627 11305
rect 20070 11228 20076 11280
rect 20128 11268 20134 11280
rect 22664 11268 22692 11299
rect 24210 11296 24216 11308
rect 24268 11296 24274 11348
rect 24854 11336 24860 11348
rect 24320 11308 24860 11336
rect 20128 11240 22692 11268
rect 20128 11228 20134 11240
rect 19981 11203 20039 11209
rect 19981 11169 19993 11203
rect 20027 11169 20039 11203
rect 19981 11163 20039 11169
rect 21177 11203 21235 11209
rect 21177 11169 21189 11203
rect 21223 11169 21235 11203
rect 21177 11163 21235 11169
rect 21821 11203 21879 11209
rect 21821 11169 21833 11203
rect 21867 11200 21879 11203
rect 22278 11200 22284 11212
rect 21867 11172 22284 11200
rect 21867 11169 21879 11172
rect 21821 11163 21879 11169
rect 15896 11104 16160 11132
rect 16393 11135 16451 11141
rect 15896 11092 15902 11104
rect 16393 11101 16405 11135
rect 16439 11132 16451 11135
rect 16666 11132 16672 11144
rect 16439 11104 16672 11132
rect 16439 11101 16451 11104
rect 16393 11095 16451 11101
rect 16666 11092 16672 11104
rect 16724 11092 16730 11144
rect 18877 11135 18935 11141
rect 18877 11132 18889 11135
rect 17236 11104 18889 11132
rect 4614 11024 4620 11076
rect 4672 11024 4678 11076
rect 8389 11067 8447 11073
rect 8389 11033 8401 11067
rect 8435 11064 8447 11067
rect 12894 11064 12900 11076
rect 8435 11036 12900 11064
rect 8435 11033 8447 11036
rect 8389 11027 8447 11033
rect 12894 11024 12900 11036
rect 12952 11024 12958 11076
rect 13081 11067 13139 11073
rect 13081 11033 13093 11067
rect 13127 11033 13139 11067
rect 13081 11027 13139 11033
rect 14001 11067 14059 11073
rect 14001 11033 14013 11067
rect 14047 11064 14059 11067
rect 15286 11064 15292 11076
rect 14047 11036 15292 11064
rect 14047 11033 14059 11036
rect 14001 11027 14059 11033
rect 5629 10999 5687 11005
rect 5629 10965 5641 10999
rect 5675 10996 5687 10999
rect 9858 10996 9864 11008
rect 5675 10968 9864 10996
rect 5675 10965 5687 10968
rect 5629 10959 5687 10965
rect 9858 10956 9864 10968
rect 9916 10956 9922 11008
rect 10045 10999 10103 11005
rect 10045 10965 10057 10999
rect 10091 10996 10103 10999
rect 10502 10996 10508 11008
rect 10091 10968 10508 10996
rect 10091 10965 10103 10968
rect 10045 10959 10103 10965
rect 10502 10956 10508 10968
rect 10560 10956 10566 11008
rect 13096 10996 13124 11027
rect 15286 11024 15292 11036
rect 15344 11024 15350 11076
rect 17236 11073 17264 11104
rect 18877 11101 18889 11104
rect 18923 11132 18935 11135
rect 18966 11132 18972 11144
rect 18923 11104 18972 11132
rect 18923 11101 18935 11104
rect 18877 11095 18935 11101
rect 18966 11092 18972 11104
rect 19024 11092 19030 11144
rect 21192 11132 21220 11163
rect 22278 11160 22284 11172
rect 22336 11160 22342 11212
rect 22462 11200 22468 11212
rect 22423 11172 22468 11200
rect 22462 11160 22468 11172
rect 22520 11160 22526 11212
rect 22664 11200 22692 11240
rect 24320 11209 24348 11308
rect 24854 11296 24860 11308
rect 24912 11296 24918 11348
rect 25593 11339 25651 11345
rect 25593 11305 25605 11339
rect 25639 11336 25651 11339
rect 27614 11336 27620 11348
rect 25639 11308 27620 11336
rect 25639 11305 25651 11308
rect 25593 11299 25651 11305
rect 27614 11296 27620 11308
rect 27672 11296 27678 11348
rect 27706 11296 27712 11348
rect 27764 11336 27770 11348
rect 30466 11336 30472 11348
rect 27764 11308 30472 11336
rect 27764 11296 27770 11308
rect 30466 11296 30472 11308
rect 30524 11296 30530 11348
rect 30742 11296 30748 11348
rect 30800 11336 30806 11348
rect 36998 11336 37004 11348
rect 30800 11308 34468 11336
rect 36959 11308 37004 11336
rect 30800 11296 30806 11308
rect 25958 11268 25964 11280
rect 24688 11240 25964 11268
rect 24688 11209 24716 11240
rect 25958 11228 25964 11240
rect 26016 11228 26022 11280
rect 31938 11268 31944 11280
rect 28920 11240 31248 11268
rect 23385 11203 23443 11209
rect 23385 11200 23397 11203
rect 22664 11172 23397 11200
rect 23385 11169 23397 11172
rect 23431 11169 23443 11203
rect 23385 11163 23443 11169
rect 24305 11203 24363 11209
rect 24305 11169 24317 11203
rect 24351 11169 24363 11203
rect 24305 11163 24363 11169
rect 24673 11203 24731 11209
rect 24673 11169 24685 11203
rect 24719 11169 24731 11203
rect 24673 11163 24731 11169
rect 25409 11203 25467 11209
rect 25409 11169 25421 11203
rect 25455 11200 25467 11203
rect 25590 11200 25596 11212
rect 25455 11172 25596 11200
rect 25455 11169 25467 11172
rect 25409 11163 25467 11169
rect 25590 11160 25596 11172
rect 25648 11160 25654 11212
rect 26513 11203 26571 11209
rect 26513 11169 26525 11203
rect 26559 11200 26571 11203
rect 27154 11200 27160 11212
rect 26559 11172 27160 11200
rect 26559 11169 26571 11172
rect 26513 11163 26571 11169
rect 27154 11160 27160 11172
rect 27212 11160 27218 11212
rect 28626 11200 28632 11212
rect 28587 11172 28632 11200
rect 28626 11160 28632 11172
rect 28684 11160 28690 11212
rect 22480 11132 22508 11160
rect 21192 11104 22508 11132
rect 26789 11135 26847 11141
rect 26789 11101 26801 11135
rect 26835 11132 26847 11135
rect 28920 11132 28948 11240
rect 29178 11200 29184 11212
rect 29139 11172 29184 11200
rect 29178 11160 29184 11172
rect 29236 11160 29242 11212
rect 29365 11203 29423 11209
rect 29365 11169 29377 11203
rect 29411 11169 29423 11203
rect 29365 11163 29423 11169
rect 29086 11132 29092 11144
rect 26835 11104 28948 11132
rect 29047 11104 29092 11132
rect 26835 11101 26847 11104
rect 26789 11095 26847 11101
rect 29086 11092 29092 11104
rect 29144 11092 29150 11144
rect 17221 11067 17279 11073
rect 17221 11033 17233 11067
rect 17267 11033 17279 11067
rect 17221 11027 17279 11033
rect 18322 11024 18328 11076
rect 18380 11064 18386 11076
rect 20714 11064 20720 11076
rect 18380 11036 20720 11064
rect 18380 11024 18386 11036
rect 20714 11024 20720 11036
rect 20772 11064 20778 11076
rect 21269 11067 21327 11073
rect 21269 11064 21281 11067
rect 20772 11036 21281 11064
rect 20772 11024 20778 11036
rect 21269 11033 21281 11036
rect 21315 11033 21327 11067
rect 21269 11027 21327 11033
rect 21450 11024 21456 11076
rect 21508 11064 21514 11076
rect 24121 11067 24179 11073
rect 24121 11064 24133 11067
rect 21508 11036 24133 11064
rect 21508 11024 21514 11036
rect 24121 11033 24133 11036
rect 24167 11033 24179 11067
rect 24121 11027 24179 11033
rect 24857 11067 24915 11073
rect 24857 11033 24869 11067
rect 24903 11064 24915 11067
rect 26510 11064 26516 11076
rect 24903 11036 26516 11064
rect 24903 11033 24915 11036
rect 24857 11027 24915 11033
rect 26510 11024 26516 11036
rect 26568 11024 26574 11076
rect 27893 11067 27951 11073
rect 27893 11064 27905 11067
rect 27448 11036 27905 11064
rect 13814 10996 13820 11008
rect 13096 10968 13820 10996
rect 13814 10956 13820 10968
rect 13872 10956 13878 11008
rect 21910 10996 21916 11008
rect 21871 10968 21916 10996
rect 21910 10956 21916 10968
rect 21968 10956 21974 11008
rect 26142 10956 26148 11008
rect 26200 10996 26206 11008
rect 27448 10996 27476 11036
rect 27893 11033 27905 11036
rect 27939 11033 27951 11067
rect 27893 11027 27951 11033
rect 28074 11024 28080 11076
rect 28132 11064 28138 11076
rect 29380 11064 29408 11163
rect 29822 11160 29828 11212
rect 29880 11200 29886 11212
rect 29917 11203 29975 11209
rect 29917 11200 29929 11203
rect 29880 11172 29929 11200
rect 29880 11160 29886 11172
rect 29917 11169 29929 11172
rect 29963 11169 29975 11203
rect 29917 11163 29975 11169
rect 30558 11132 30564 11144
rect 30519 11104 30564 11132
rect 30558 11092 30564 11104
rect 30616 11092 30622 11144
rect 31113 11135 31171 11141
rect 31113 11101 31125 11135
rect 31159 11101 31171 11135
rect 31220 11132 31248 11240
rect 31588 11240 31944 11268
rect 31294 11160 31300 11212
rect 31352 11200 31358 11212
rect 31588 11209 31616 11240
rect 31938 11228 31944 11240
rect 31996 11268 32002 11280
rect 33134 11268 33140 11280
rect 31996 11240 33140 11268
rect 31996 11228 32002 11240
rect 33134 11228 33140 11240
rect 33192 11228 33198 11280
rect 31435 11203 31493 11209
rect 31435 11200 31447 11203
rect 31352 11172 31447 11200
rect 31352 11160 31358 11172
rect 31435 11169 31447 11172
rect 31481 11169 31493 11203
rect 31435 11163 31493 11169
rect 31573 11203 31631 11209
rect 31573 11169 31585 11203
rect 31619 11169 31631 11203
rect 31573 11163 31631 11169
rect 31754 11160 31760 11212
rect 31812 11200 31818 11212
rect 32125 11203 32183 11209
rect 32125 11200 32137 11203
rect 31812 11172 32137 11200
rect 31812 11160 31818 11172
rect 32125 11169 32137 11172
rect 32171 11169 32183 11203
rect 32674 11200 32680 11212
rect 32635 11172 32680 11200
rect 32125 11163 32183 11169
rect 32674 11160 32680 11172
rect 32732 11160 32738 11212
rect 33042 11200 33048 11212
rect 33003 11172 33048 11200
rect 33042 11160 33048 11172
rect 33100 11160 33106 11212
rect 34054 11200 34060 11212
rect 34015 11172 34060 11200
rect 34054 11160 34060 11172
rect 34112 11160 34118 11212
rect 34440 11209 34468 11308
rect 36998 11296 37004 11308
rect 37056 11296 37062 11348
rect 34425 11203 34483 11209
rect 34425 11169 34437 11203
rect 34471 11169 34483 11203
rect 34425 11163 34483 11169
rect 31220 11104 32260 11132
rect 31113 11095 31171 11101
rect 28132 11036 29408 11064
rect 31128 11064 31156 11095
rect 31754 11064 31760 11076
rect 31128 11036 31760 11064
rect 28132 11024 28138 11036
rect 31754 11024 31760 11036
rect 31812 11024 31818 11076
rect 32232 11073 32260 11104
rect 33594 11092 33600 11144
rect 33652 11132 33658 11144
rect 34238 11132 34244 11144
rect 33652 11104 34244 11132
rect 33652 11092 33658 11104
rect 34238 11092 34244 11104
rect 34296 11132 34302 11144
rect 34701 11135 34759 11141
rect 34701 11132 34713 11135
rect 34296 11104 34713 11132
rect 34296 11092 34302 11104
rect 34701 11101 34713 11104
rect 34747 11101 34759 11135
rect 34701 11095 34759 11101
rect 35342 11092 35348 11144
rect 35400 11132 35406 11144
rect 35437 11135 35495 11141
rect 35437 11132 35449 11135
rect 35400 11104 35449 11132
rect 35400 11092 35406 11104
rect 35437 11101 35449 11104
rect 35483 11101 35495 11135
rect 35710 11132 35716 11144
rect 35671 11104 35716 11132
rect 35437 11095 35495 11101
rect 35710 11092 35716 11104
rect 35768 11092 35774 11144
rect 32217 11067 32275 11073
rect 32217 11033 32229 11067
rect 32263 11033 32275 11067
rect 32217 11027 32275 11033
rect 34149 11067 34207 11073
rect 34149 11033 34161 11067
rect 34195 11064 34207 11067
rect 34195 11036 35480 11064
rect 34195 11033 34207 11036
rect 34149 11027 34207 11033
rect 26200 10968 27476 10996
rect 26200 10956 26206 10968
rect 27522 10956 27528 11008
rect 27580 10996 27586 11008
rect 33870 10996 33876 11008
rect 27580 10968 33876 10996
rect 27580 10956 27586 10968
rect 33870 10956 33876 10968
rect 33928 10956 33934 11008
rect 35452 10996 35480 11036
rect 35894 10996 35900 11008
rect 35452 10968 35900 10996
rect 35894 10956 35900 10968
rect 35952 10956 35958 11008
rect 1104 10906 38824 10928
rect 1104 10854 4246 10906
rect 4298 10854 4310 10906
rect 4362 10854 4374 10906
rect 4426 10854 4438 10906
rect 4490 10854 34966 10906
rect 35018 10854 35030 10906
rect 35082 10854 35094 10906
rect 35146 10854 35158 10906
rect 35210 10854 38824 10906
rect 1104 10832 38824 10854
rect 8662 10752 8668 10804
rect 8720 10792 8726 10804
rect 15838 10792 15844 10804
rect 8720 10764 15608 10792
rect 15799 10764 15844 10792
rect 8720 10752 8726 10764
rect 10318 10684 10324 10736
rect 10376 10724 10382 10736
rect 13170 10724 13176 10736
rect 10376 10696 13176 10724
rect 10376 10684 10382 10696
rect 13170 10684 13176 10696
rect 13228 10684 13234 10736
rect 15580 10724 15608 10764
rect 15838 10752 15844 10764
rect 15896 10752 15902 10804
rect 16850 10792 16856 10804
rect 16592 10764 16856 10792
rect 16592 10736 16620 10764
rect 16850 10752 16856 10764
rect 16908 10752 16914 10804
rect 22554 10752 22560 10804
rect 22612 10792 22618 10804
rect 22612 10764 35848 10792
rect 22612 10752 22618 10764
rect 16574 10724 16580 10736
rect 13280 10696 14320 10724
rect 4614 10656 4620 10668
rect 4356 10628 4620 10656
rect 2133 10591 2191 10597
rect 2133 10557 2145 10591
rect 2179 10588 2191 10591
rect 2222 10588 2228 10600
rect 2179 10560 2228 10588
rect 2179 10557 2191 10560
rect 2133 10551 2191 10557
rect 2222 10548 2228 10560
rect 2280 10548 2286 10600
rect 2958 10548 2964 10600
rect 3016 10588 3022 10600
rect 3053 10591 3111 10597
rect 3053 10588 3065 10591
rect 3016 10560 3065 10588
rect 3016 10548 3022 10560
rect 3053 10557 3065 10560
rect 3099 10557 3111 10591
rect 3053 10551 3111 10557
rect 3142 10548 3148 10600
rect 3200 10588 3206 10600
rect 4356 10597 4384 10628
rect 4614 10616 4620 10628
rect 4672 10616 4678 10668
rect 5261 10659 5319 10665
rect 5261 10625 5273 10659
rect 5307 10656 5319 10659
rect 6178 10656 6184 10668
rect 5307 10628 6184 10656
rect 5307 10625 5319 10628
rect 5261 10619 5319 10625
rect 6178 10616 6184 10628
rect 6236 10616 6242 10668
rect 6273 10659 6331 10665
rect 6273 10625 6285 10659
rect 6319 10656 6331 10659
rect 6730 10656 6736 10668
rect 6319 10628 6736 10656
rect 6319 10625 6331 10628
rect 6273 10619 6331 10625
rect 6730 10616 6736 10628
rect 6788 10616 6794 10668
rect 9493 10659 9551 10665
rect 9493 10625 9505 10659
rect 9539 10656 9551 10659
rect 13280 10656 13308 10696
rect 9539 10628 13308 10656
rect 9539 10625 9551 10628
rect 9493 10619 9551 10625
rect 14090 10616 14096 10668
rect 14148 10656 14154 10668
rect 14185 10659 14243 10665
rect 14185 10656 14197 10659
rect 14148 10628 14197 10656
rect 14148 10616 14154 10628
rect 14185 10625 14197 10628
rect 14231 10625 14243 10659
rect 14292 10656 14320 10696
rect 15580 10696 16580 10724
rect 15580 10656 15608 10696
rect 16574 10684 16580 10696
rect 16632 10684 16638 10736
rect 16669 10727 16727 10733
rect 16669 10693 16681 10727
rect 16715 10724 16727 10727
rect 17218 10724 17224 10736
rect 16715 10696 17224 10724
rect 16715 10693 16727 10696
rect 16669 10687 16727 10693
rect 17218 10684 17224 10696
rect 17276 10684 17282 10736
rect 18141 10727 18199 10733
rect 18141 10693 18153 10727
rect 18187 10693 18199 10727
rect 18141 10687 18199 10693
rect 21177 10727 21235 10733
rect 21177 10693 21189 10727
rect 21223 10724 21235 10727
rect 22094 10724 22100 10736
rect 21223 10696 22100 10724
rect 21223 10693 21235 10696
rect 21177 10687 21235 10693
rect 18156 10656 18184 10687
rect 22094 10684 22100 10696
rect 22152 10684 22158 10736
rect 22830 10684 22836 10736
rect 22888 10684 22894 10736
rect 23658 10684 23664 10736
rect 23716 10724 23722 10736
rect 23753 10727 23811 10733
rect 23753 10724 23765 10727
rect 23716 10696 23765 10724
rect 23716 10684 23722 10696
rect 23753 10693 23765 10696
rect 23799 10693 23811 10727
rect 23753 10687 23811 10693
rect 23934 10684 23940 10736
rect 23992 10724 23998 10736
rect 27522 10724 27528 10736
rect 23992 10696 27528 10724
rect 23992 10684 23998 10696
rect 27522 10684 27528 10696
rect 27580 10684 27586 10736
rect 27706 10684 27712 10736
rect 27764 10724 27770 10736
rect 27764 10696 28212 10724
rect 27764 10684 27770 10696
rect 14292 10628 14780 10656
rect 15580 10628 15700 10656
rect 14185 10619 14243 10625
rect 4341 10591 4399 10597
rect 3200 10560 3245 10588
rect 3200 10548 3206 10560
rect 4341 10557 4353 10591
rect 4387 10557 4399 10591
rect 4341 10551 4399 10557
rect 4525 10591 4583 10597
rect 4525 10557 4537 10591
rect 4571 10557 4583 10591
rect 4798 10588 4804 10600
rect 4759 10560 4804 10588
rect 4525 10551 4583 10557
rect 3602 10520 3608 10532
rect 3563 10492 3608 10520
rect 3602 10480 3608 10492
rect 3660 10480 3666 10532
rect 4540 10520 4568 10551
rect 4798 10548 4804 10560
rect 4856 10548 4862 10600
rect 5721 10591 5779 10597
rect 5721 10557 5733 10591
rect 5767 10557 5779 10591
rect 5721 10551 5779 10557
rect 5258 10520 5264 10532
rect 4540 10492 5264 10520
rect 5258 10480 5264 10492
rect 5316 10480 5322 10532
rect 5736 10520 5764 10551
rect 5810 10548 5816 10600
rect 5868 10588 5874 10600
rect 5868 10560 5913 10588
rect 5868 10548 5874 10560
rect 6638 10548 6644 10600
rect 6696 10588 6702 10600
rect 7469 10591 7527 10597
rect 7469 10588 7481 10591
rect 6696 10560 7481 10588
rect 6696 10548 6702 10560
rect 7469 10557 7481 10560
rect 7515 10557 7527 10591
rect 7469 10551 7527 10557
rect 8021 10591 8079 10597
rect 8021 10557 8033 10591
rect 8067 10557 8079 10591
rect 8294 10588 8300 10600
rect 8255 10560 8300 10588
rect 8021 10551 8079 10557
rect 7282 10520 7288 10532
rect 5736 10492 7288 10520
rect 7282 10480 7288 10492
rect 7340 10480 7346 10532
rect 8036 10520 8064 10551
rect 8294 10548 8300 10560
rect 8352 10548 8358 10600
rect 9401 10591 9459 10597
rect 9401 10557 9413 10591
rect 9447 10588 9459 10591
rect 9674 10588 9680 10600
rect 9447 10560 9680 10588
rect 9447 10557 9459 10560
rect 9401 10551 9459 10557
rect 9674 10548 9680 10560
rect 9732 10548 9738 10600
rect 9861 10591 9919 10597
rect 9861 10557 9873 10591
rect 9907 10588 9919 10591
rect 10321 10591 10379 10597
rect 10321 10588 10333 10591
rect 9907 10560 10333 10588
rect 9907 10557 9919 10560
rect 9861 10551 9919 10557
rect 10321 10557 10333 10560
rect 10367 10557 10379 10591
rect 10962 10588 10968 10600
rect 10923 10560 10968 10588
rect 10321 10551 10379 10557
rect 10962 10548 10968 10560
rect 11020 10548 11026 10600
rect 11057 10591 11115 10597
rect 11057 10557 11069 10591
rect 11103 10557 11115 10591
rect 11330 10588 11336 10600
rect 11291 10560 11336 10588
rect 11057 10551 11115 10557
rect 8386 10520 8392 10532
rect 8036 10492 8392 10520
rect 8386 10480 8392 10492
rect 8444 10480 8450 10532
rect 8573 10523 8631 10529
rect 8573 10489 8585 10523
rect 8619 10520 8631 10523
rect 10226 10520 10232 10532
rect 8619 10492 10232 10520
rect 8619 10489 8631 10492
rect 8573 10483 8631 10489
rect 10226 10480 10232 10492
rect 10284 10480 10290 10532
rect 10686 10480 10692 10532
rect 10744 10520 10750 10532
rect 11072 10520 11100 10551
rect 11330 10548 11336 10560
rect 11388 10548 11394 10600
rect 11514 10588 11520 10600
rect 11475 10560 11520 10588
rect 11514 10548 11520 10560
rect 11572 10548 11578 10600
rect 11790 10548 11796 10600
rect 11848 10588 11854 10600
rect 12437 10591 12495 10597
rect 12437 10588 12449 10591
rect 11848 10560 12449 10588
rect 11848 10548 11854 10560
rect 12437 10557 12449 10560
rect 12483 10557 12495 10591
rect 12986 10588 12992 10600
rect 12947 10560 12992 10588
rect 12437 10551 12495 10557
rect 12986 10548 12992 10560
rect 13044 10548 13050 10600
rect 13262 10588 13268 10600
rect 13223 10560 13268 10588
rect 13262 10548 13268 10560
rect 13320 10548 13326 10600
rect 14645 10591 14703 10597
rect 14645 10557 14657 10591
rect 14691 10557 14703 10591
rect 14645 10551 14703 10557
rect 13541 10523 13599 10529
rect 10744 10492 11836 10520
rect 10744 10480 10750 10492
rect 11808 10464 11836 10492
rect 13541 10489 13553 10523
rect 13587 10520 13599 10523
rect 13998 10520 14004 10532
rect 13587 10492 14004 10520
rect 13587 10489 13599 10492
rect 13541 10483 13599 10489
rect 13998 10480 14004 10492
rect 14056 10480 14062 10532
rect 2314 10452 2320 10464
rect 2275 10424 2320 10452
rect 2314 10412 2320 10424
rect 2372 10412 2378 10464
rect 11790 10412 11796 10464
rect 11848 10412 11854 10464
rect 14660 10452 14688 10551
rect 14752 10520 14780 10628
rect 15010 10588 15016 10600
rect 14971 10560 15016 10588
rect 15010 10548 15016 10560
rect 15068 10548 15074 10600
rect 15105 10591 15163 10597
rect 15105 10557 15117 10591
rect 15151 10588 15163 10591
rect 15562 10588 15568 10600
rect 15151 10560 15568 10588
rect 15151 10557 15163 10560
rect 15105 10551 15163 10557
rect 15562 10548 15568 10560
rect 15620 10548 15626 10600
rect 15672 10597 15700 10628
rect 16500 10628 18184 10656
rect 16500 10597 16528 10628
rect 15657 10591 15715 10597
rect 15657 10557 15669 10591
rect 15703 10557 15715 10591
rect 15657 10551 15715 10557
rect 16485 10591 16543 10597
rect 16485 10557 16497 10591
rect 16531 10557 16543 10591
rect 16485 10551 16543 10557
rect 16945 10591 17003 10597
rect 16945 10557 16957 10591
rect 16991 10557 17003 10591
rect 17402 10588 17408 10600
rect 17363 10560 17408 10588
rect 16945 10551 17003 10557
rect 16960 10520 16988 10551
rect 17402 10548 17408 10560
rect 17460 10548 17466 10600
rect 18322 10588 18328 10600
rect 18283 10560 18328 10588
rect 18322 10548 18328 10560
rect 18380 10548 18386 10600
rect 18598 10588 18604 10600
rect 18559 10560 18604 10588
rect 18598 10548 18604 10560
rect 18656 10548 18662 10600
rect 19426 10588 19432 10600
rect 19387 10560 19432 10588
rect 19426 10548 19432 10560
rect 19484 10548 19490 10600
rect 19981 10591 20039 10597
rect 19981 10557 19993 10591
rect 20027 10557 20039 10591
rect 19981 10551 20039 10557
rect 21085 10591 21143 10597
rect 21085 10557 21097 10591
rect 21131 10557 21143 10591
rect 21085 10551 21143 10557
rect 14752 10492 16988 10520
rect 15470 10452 15476 10464
rect 14660 10424 15476 10452
rect 15470 10412 15476 10424
rect 15528 10412 15534 10464
rect 19334 10412 19340 10464
rect 19392 10452 19398 10464
rect 19521 10455 19579 10461
rect 19521 10452 19533 10455
rect 19392 10424 19533 10452
rect 19392 10412 19398 10424
rect 19521 10421 19533 10424
rect 19567 10421 19579 10455
rect 19996 10452 20024 10551
rect 21100 10520 21128 10551
rect 21818 10548 21824 10600
rect 21876 10597 21882 10600
rect 21876 10591 21925 10597
rect 21876 10557 21879 10591
rect 21913 10557 21925 10591
rect 22002 10588 22008 10600
rect 21963 10560 22008 10588
rect 21876 10551 21925 10557
rect 21876 10548 21882 10551
rect 22002 10548 22008 10560
rect 22060 10548 22066 10600
rect 22370 10588 22376 10600
rect 22331 10560 22376 10588
rect 22370 10548 22376 10560
rect 22428 10548 22434 10600
rect 22462 10548 22468 10600
rect 22520 10588 22526 10600
rect 22848 10588 22876 10684
rect 26789 10659 26847 10665
rect 26789 10625 26801 10659
rect 26835 10656 26847 10659
rect 27798 10656 27804 10668
rect 26835 10628 27804 10656
rect 26835 10625 26847 10628
rect 26789 10619 26847 10625
rect 27798 10616 27804 10628
rect 27856 10616 27862 10668
rect 27982 10656 27988 10668
rect 27943 10628 27988 10656
rect 27982 10616 27988 10628
rect 28040 10616 28046 10668
rect 28184 10656 28212 10696
rect 28534 10684 28540 10736
rect 28592 10724 28598 10736
rect 28902 10724 28908 10736
rect 28592 10696 28908 10724
rect 28592 10684 28598 10696
rect 28902 10684 28908 10696
rect 28960 10684 28966 10736
rect 29641 10727 29699 10733
rect 29641 10693 29653 10727
rect 29687 10724 29699 10727
rect 30098 10724 30104 10736
rect 29687 10696 30104 10724
rect 29687 10693 29699 10696
rect 29641 10687 29699 10693
rect 30098 10684 30104 10696
rect 30156 10684 30162 10736
rect 31205 10727 31263 10733
rect 31205 10693 31217 10727
rect 31251 10724 31263 10727
rect 32214 10724 32220 10736
rect 31251 10696 32220 10724
rect 31251 10693 31263 10696
rect 31205 10687 31263 10693
rect 32214 10684 32220 10696
rect 32272 10684 32278 10736
rect 32968 10696 35756 10724
rect 28184 10628 28304 10656
rect 23658 10588 23664 10600
rect 22520 10560 22876 10588
rect 23619 10560 23664 10588
rect 22520 10548 22526 10560
rect 23658 10548 23664 10560
rect 23716 10548 23722 10600
rect 24946 10588 24952 10600
rect 24907 10560 24952 10588
rect 24946 10548 24952 10560
rect 25004 10548 25010 10600
rect 25406 10548 25412 10600
rect 25464 10588 25470 10600
rect 25685 10591 25743 10597
rect 25685 10588 25697 10591
rect 25464 10560 25697 10588
rect 25464 10548 25470 10560
rect 25685 10557 25697 10560
rect 25731 10588 25743 10591
rect 26142 10588 26148 10600
rect 25731 10560 26148 10588
rect 25731 10557 25743 10560
rect 25685 10551 25743 10557
rect 26142 10548 26148 10560
rect 26200 10548 26206 10600
rect 26510 10548 26516 10600
rect 26568 10588 26574 10600
rect 28166 10588 28172 10600
rect 26568 10560 28028 10588
rect 28127 10560 28172 10588
rect 26568 10548 26574 10560
rect 28000 10532 28028 10560
rect 28166 10548 28172 10560
rect 28224 10548 28230 10600
rect 28276 10597 28304 10628
rect 29730 10616 29736 10668
rect 29788 10656 29794 10668
rect 29788 10628 30236 10656
rect 29788 10616 29794 10628
rect 30208 10600 30236 10628
rect 31662 10616 31668 10668
rect 31720 10656 31726 10668
rect 31757 10659 31815 10665
rect 31757 10656 31769 10659
rect 31720 10628 31769 10656
rect 31720 10616 31726 10628
rect 31757 10625 31769 10628
rect 31803 10625 31815 10659
rect 32858 10656 32864 10668
rect 31757 10619 31815 10625
rect 31864 10628 32864 10656
rect 28261 10591 28319 10597
rect 28261 10557 28273 10591
rect 28307 10557 28319 10591
rect 29822 10588 29828 10600
rect 29783 10560 29828 10588
rect 28261 10551 28319 10557
rect 29822 10548 29828 10560
rect 29880 10548 29886 10600
rect 30006 10588 30012 10600
rect 29967 10560 30012 10588
rect 30006 10548 30012 10560
rect 30064 10548 30070 10600
rect 30190 10548 30196 10600
rect 30248 10588 30254 10600
rect 31021 10591 31079 10597
rect 30248 10560 30341 10588
rect 30248 10548 30254 10560
rect 31021 10557 31033 10591
rect 31067 10588 31079 10591
rect 31864 10588 31892 10628
rect 32858 10616 32864 10628
rect 32916 10616 32922 10668
rect 32263 10591 32321 10597
rect 32263 10588 32275 10591
rect 31067 10560 31892 10588
rect 31956 10560 32275 10588
rect 31067 10557 31079 10560
rect 31021 10551 31079 10557
rect 22830 10520 22836 10532
rect 21100 10492 22836 10520
rect 22830 10480 22836 10492
rect 22888 10480 22894 10532
rect 23017 10523 23075 10529
rect 23017 10489 23029 10523
rect 23063 10520 23075 10523
rect 23290 10520 23296 10532
rect 23063 10492 23296 10520
rect 23063 10489 23075 10492
rect 23017 10483 23075 10489
rect 23290 10480 23296 10492
rect 23348 10480 23354 10532
rect 26234 10520 26240 10532
rect 26195 10492 26240 10520
rect 26234 10480 26240 10492
rect 26292 10480 26298 10532
rect 27062 10520 27068 10532
rect 27023 10492 27068 10520
rect 27062 10480 27068 10492
rect 27120 10480 27126 10532
rect 27154 10480 27160 10532
rect 27212 10520 27218 10532
rect 27522 10520 27528 10532
rect 27212 10492 27257 10520
rect 27483 10492 27528 10520
rect 27212 10480 27218 10492
rect 27522 10480 27528 10492
rect 27580 10480 27586 10532
rect 27982 10480 27988 10532
rect 28040 10480 28046 10532
rect 28353 10523 28411 10529
rect 28353 10489 28365 10523
rect 28399 10520 28411 10523
rect 28721 10523 28779 10529
rect 28399 10492 28672 10520
rect 28399 10489 28411 10492
rect 28353 10483 28411 10489
rect 21634 10452 21640 10464
rect 19996 10424 21640 10452
rect 19521 10415 19579 10421
rect 21634 10412 21640 10424
rect 21692 10412 21698 10464
rect 21726 10412 21732 10464
rect 21784 10452 21790 10464
rect 26326 10452 26332 10464
rect 21784 10424 26332 10452
rect 21784 10412 21790 10424
rect 26326 10412 26332 10424
rect 26384 10412 26390 10464
rect 26973 10455 27031 10461
rect 26973 10421 26985 10455
rect 27019 10452 27031 10455
rect 27614 10452 27620 10464
rect 27019 10424 27620 10452
rect 27019 10421 27031 10424
rect 26973 10415 27031 10421
rect 27614 10412 27620 10424
rect 27672 10452 27678 10464
rect 28442 10452 28448 10464
rect 27672 10424 28448 10452
rect 27672 10412 27678 10424
rect 28442 10412 28448 10424
rect 28500 10412 28506 10464
rect 28644 10452 28672 10492
rect 28721 10489 28733 10523
rect 28767 10520 28779 10523
rect 28810 10520 28816 10532
rect 28767 10492 28816 10520
rect 28767 10489 28779 10492
rect 28721 10483 28779 10489
rect 28810 10480 28816 10492
rect 28868 10480 28874 10532
rect 31110 10480 31116 10532
rect 31168 10520 31174 10532
rect 31956 10520 31984 10560
rect 32263 10557 32275 10560
rect 32309 10557 32321 10591
rect 32582 10588 32588 10600
rect 32543 10560 32588 10588
rect 32263 10551 32321 10557
rect 32582 10548 32588 10560
rect 32640 10548 32646 10600
rect 32769 10591 32827 10597
rect 32769 10557 32781 10591
rect 32815 10588 32827 10591
rect 32968 10588 32996 10696
rect 32815 10560 32996 10588
rect 32815 10557 32827 10560
rect 32769 10551 32827 10557
rect 33042 10548 33048 10600
rect 33100 10588 33106 10600
rect 33229 10591 33287 10597
rect 33229 10588 33241 10591
rect 33100 10560 33241 10588
rect 33100 10548 33106 10560
rect 33229 10557 33241 10560
rect 33275 10557 33287 10591
rect 33594 10588 33600 10600
rect 33555 10560 33600 10588
rect 33229 10551 33287 10557
rect 33594 10548 33600 10560
rect 33652 10548 33658 10600
rect 33962 10548 33968 10600
rect 34020 10588 34026 10600
rect 34057 10591 34115 10597
rect 34057 10588 34069 10591
rect 34020 10560 34069 10588
rect 34020 10548 34026 10560
rect 34057 10557 34069 10560
rect 34103 10557 34115 10591
rect 34057 10551 34115 10557
rect 34146 10548 34152 10600
rect 34204 10588 34210 10600
rect 34885 10591 34943 10597
rect 34885 10588 34897 10591
rect 34204 10560 34897 10588
rect 34204 10548 34210 10560
rect 34885 10557 34897 10560
rect 34931 10557 34943 10591
rect 34885 10551 34943 10557
rect 35437 10591 35495 10597
rect 35437 10557 35449 10591
rect 35483 10557 35495 10591
rect 35437 10551 35495 10557
rect 31168 10492 31984 10520
rect 34333 10523 34391 10529
rect 31168 10480 31174 10492
rect 34333 10489 34345 10523
rect 34379 10520 34391 10523
rect 35452 10520 35480 10551
rect 34379 10492 35480 10520
rect 35728 10520 35756 10696
rect 35820 10588 35848 10764
rect 35894 10616 35900 10668
rect 35952 10656 35958 10668
rect 36446 10656 36452 10668
rect 35952 10628 35997 10656
rect 36407 10628 36452 10656
rect 35952 10616 35958 10628
rect 36446 10616 36452 10628
rect 36504 10616 36510 10668
rect 36725 10591 36783 10597
rect 36725 10588 36737 10591
rect 35820 10560 36737 10588
rect 36725 10557 36737 10560
rect 36771 10557 36783 10591
rect 36725 10551 36783 10557
rect 36078 10520 36084 10532
rect 35728 10492 36084 10520
rect 34379 10489 34391 10492
rect 34333 10483 34391 10489
rect 36078 10480 36084 10492
rect 36136 10480 36142 10532
rect 38102 10520 38108 10532
rect 38063 10492 38108 10520
rect 38102 10480 38108 10492
rect 38160 10480 38166 10532
rect 32122 10452 32128 10464
rect 28644 10424 32128 10452
rect 32122 10412 32128 10424
rect 32180 10412 32186 10464
rect 34698 10412 34704 10464
rect 34756 10452 34762 10464
rect 34977 10455 35035 10461
rect 34977 10452 34989 10455
rect 34756 10424 34989 10452
rect 34756 10412 34762 10424
rect 34977 10421 34989 10424
rect 35023 10421 35035 10455
rect 36096 10452 36124 10480
rect 37182 10452 37188 10464
rect 36096 10424 37188 10452
rect 34977 10415 35035 10421
rect 37182 10412 37188 10424
rect 37240 10412 37246 10464
rect 1104 10362 38824 10384
rect 1104 10310 19606 10362
rect 19658 10310 19670 10362
rect 19722 10310 19734 10362
rect 19786 10310 19798 10362
rect 19850 10310 38824 10362
rect 1104 10288 38824 10310
rect 3142 10248 3148 10260
rect 3103 10220 3148 10248
rect 3142 10208 3148 10220
rect 3200 10208 3206 10260
rect 5810 10208 5816 10260
rect 5868 10248 5874 10260
rect 6917 10251 6975 10257
rect 6917 10248 6929 10251
rect 5868 10220 6929 10248
rect 5868 10208 5874 10220
rect 6917 10217 6929 10220
rect 6963 10217 6975 10251
rect 6917 10211 6975 10217
rect 7837 10251 7895 10257
rect 7837 10217 7849 10251
rect 7883 10248 7895 10251
rect 8294 10248 8300 10260
rect 7883 10220 8300 10248
rect 7883 10217 7895 10220
rect 7837 10211 7895 10217
rect 8294 10208 8300 10220
rect 8352 10208 8358 10260
rect 8570 10208 8576 10260
rect 8628 10248 8634 10260
rect 10318 10248 10324 10260
rect 8628 10220 10324 10248
rect 8628 10208 8634 10220
rect 10318 10208 10324 10220
rect 10376 10208 10382 10260
rect 21726 10248 21732 10260
rect 11900 10220 21732 10248
rect 4801 10183 4859 10189
rect 4801 10149 4813 10183
rect 4847 10180 4859 10183
rect 11900 10180 11928 10220
rect 21726 10208 21732 10220
rect 21784 10208 21790 10260
rect 35802 10248 35808 10260
rect 22756 10220 35808 10248
rect 4847 10152 5672 10180
rect 4847 10149 4859 10152
rect 4801 10143 4859 10149
rect 2958 10072 2964 10124
rect 3016 10112 3022 10124
rect 4249 10115 4307 10121
rect 4249 10112 4261 10115
rect 3016 10084 4261 10112
rect 3016 10072 3022 10084
rect 4249 10081 4261 10084
rect 4295 10081 4307 10115
rect 4249 10075 4307 10081
rect 4341 10115 4399 10121
rect 4341 10081 4353 10115
rect 4387 10112 4399 10115
rect 4614 10112 4620 10124
rect 4387 10084 4620 10112
rect 4387 10081 4399 10084
rect 4341 10075 4399 10081
rect 4614 10072 4620 10084
rect 4672 10072 4678 10124
rect 5074 10072 5080 10124
rect 5132 10112 5138 10124
rect 5445 10115 5503 10121
rect 5445 10112 5457 10115
rect 5132 10084 5457 10112
rect 5132 10072 5138 10084
rect 5445 10081 5457 10084
rect 5491 10081 5503 10115
rect 5644 10112 5672 10152
rect 7852 10152 11928 10180
rect 7852 10112 7880 10152
rect 12618 10140 12624 10192
rect 12676 10180 12682 10192
rect 16666 10180 16672 10192
rect 12676 10152 12756 10180
rect 16627 10152 16672 10180
rect 12676 10140 12682 10152
rect 5644 10084 7880 10112
rect 7929 10115 7987 10121
rect 5445 10075 5503 10081
rect 7929 10081 7941 10115
rect 7975 10081 7987 10115
rect 7929 10075 7987 10081
rect 8481 10115 8539 10121
rect 8481 10081 8493 10115
rect 8527 10112 8539 10115
rect 8938 10112 8944 10124
rect 8527 10084 8944 10112
rect 8527 10081 8539 10084
rect 8481 10075 8539 10081
rect 1765 10047 1823 10053
rect 1765 10013 1777 10047
rect 1811 10013 1823 10047
rect 1765 10007 1823 10013
rect 2041 10047 2099 10053
rect 2041 10013 2053 10047
rect 2087 10044 2099 10047
rect 3602 10044 3608 10056
rect 2087 10016 3608 10044
rect 2087 10013 2099 10016
rect 2041 10007 2099 10013
rect 1394 9868 1400 9920
rect 1452 9908 1458 9920
rect 1780 9908 1808 10007
rect 3602 10004 3608 10016
rect 3660 10004 3666 10056
rect 5537 10047 5595 10053
rect 5537 10044 5549 10047
rect 5276 10016 5549 10044
rect 5276 9917 5304 10016
rect 5537 10013 5549 10016
rect 5583 10013 5595 10047
rect 5810 10044 5816 10056
rect 5771 10016 5816 10044
rect 5537 10007 5595 10013
rect 5810 10004 5816 10016
rect 5868 10004 5874 10056
rect 7944 10044 7972 10075
rect 8938 10072 8944 10084
rect 8996 10072 9002 10124
rect 9490 10112 9496 10124
rect 9451 10084 9496 10112
rect 9490 10072 9496 10084
rect 9548 10072 9554 10124
rect 9677 10115 9735 10121
rect 9677 10081 9689 10115
rect 9723 10112 9735 10115
rect 9858 10112 9864 10124
rect 9723 10084 9864 10112
rect 9723 10081 9735 10084
rect 9677 10075 9735 10081
rect 9858 10072 9864 10084
rect 9916 10072 9922 10124
rect 10134 10112 10140 10124
rect 10095 10084 10140 10112
rect 10134 10072 10140 10084
rect 10192 10072 10198 10124
rect 10226 10072 10232 10124
rect 10284 10112 10290 10124
rect 10321 10115 10379 10121
rect 10321 10112 10333 10115
rect 10284 10084 10333 10112
rect 10284 10072 10290 10084
rect 10321 10081 10333 10084
rect 10367 10081 10379 10115
rect 10502 10112 10508 10124
rect 10463 10084 10508 10112
rect 10321 10075 10379 10081
rect 10502 10072 10508 10084
rect 10560 10072 10566 10124
rect 11882 10072 11888 10124
rect 11940 10112 11946 10124
rect 12161 10115 12219 10121
rect 12161 10112 12173 10115
rect 11940 10084 12173 10112
rect 11940 10072 11946 10084
rect 12161 10081 12173 10084
rect 12207 10081 12219 10115
rect 12526 10112 12532 10124
rect 12487 10084 12532 10112
rect 12161 10075 12219 10081
rect 12526 10072 12532 10084
rect 12584 10072 12590 10124
rect 12728 10121 12756 10152
rect 16666 10140 16672 10152
rect 16724 10140 16730 10192
rect 18230 10180 18236 10192
rect 17328 10152 18236 10180
rect 12713 10115 12771 10121
rect 12713 10081 12725 10115
rect 12759 10081 12771 10115
rect 12713 10075 12771 10081
rect 13633 10115 13691 10121
rect 13633 10081 13645 10115
rect 13679 10081 13691 10115
rect 13814 10112 13820 10124
rect 13775 10084 13820 10112
rect 13633 10075 13691 10081
rect 8570 10044 8576 10056
rect 7944 10016 8576 10044
rect 8570 10004 8576 10016
rect 8628 10004 8634 10056
rect 8665 10047 8723 10053
rect 8665 10013 8677 10047
rect 8711 10013 8723 10047
rect 10152 10044 10180 10072
rect 11330 10044 11336 10056
rect 10152 10016 11336 10044
rect 8665 10007 8723 10013
rect 6730 9936 6736 9988
rect 6788 9976 6794 9988
rect 8680 9976 8708 10007
rect 11330 10004 11336 10016
rect 11388 10004 11394 10056
rect 12066 10044 12072 10056
rect 12027 10016 12072 10044
rect 12066 10004 12072 10016
rect 12124 10004 12130 10056
rect 12250 10004 12256 10056
rect 12308 10044 12314 10056
rect 13648 10044 13676 10075
rect 13814 10072 13820 10084
rect 13872 10072 13878 10124
rect 13998 10112 14004 10124
rect 13959 10084 14004 10112
rect 13998 10072 14004 10084
rect 14056 10072 14062 10124
rect 15746 10112 15752 10124
rect 15707 10084 15752 10112
rect 15746 10072 15752 10084
rect 15804 10072 15810 10124
rect 16206 10112 16212 10124
rect 16167 10084 16212 10112
rect 16206 10072 16212 10084
rect 16264 10072 16270 10124
rect 17328 10121 17356 10152
rect 18230 10140 18236 10152
rect 18288 10140 18294 10192
rect 18325 10183 18383 10189
rect 18325 10149 18337 10183
rect 18371 10180 18383 10183
rect 18598 10180 18604 10192
rect 18371 10152 18604 10180
rect 18371 10149 18383 10152
rect 18325 10143 18383 10149
rect 18598 10140 18604 10152
rect 18656 10140 18662 10192
rect 19058 10140 19064 10192
rect 19116 10180 19122 10192
rect 19116 10152 20024 10180
rect 19116 10140 19122 10152
rect 17313 10115 17371 10121
rect 17313 10081 17325 10115
rect 17359 10081 17371 10115
rect 17313 10075 17371 10081
rect 17402 10072 17408 10124
rect 17460 10112 17466 10124
rect 17460 10084 17505 10112
rect 17460 10072 17466 10084
rect 17586 10072 17592 10124
rect 17644 10112 17650 10124
rect 17681 10115 17739 10121
rect 17681 10112 17693 10115
rect 17644 10084 17693 10112
rect 17644 10072 17650 10084
rect 17681 10081 17693 10084
rect 17727 10081 17739 10115
rect 17681 10075 17739 10081
rect 18969 10115 19027 10121
rect 18969 10081 18981 10115
rect 19015 10112 19027 10115
rect 19150 10112 19156 10124
rect 19015 10084 19156 10112
rect 19015 10081 19027 10084
rect 18969 10075 19027 10081
rect 19150 10072 19156 10084
rect 19208 10072 19214 10124
rect 19334 10112 19340 10124
rect 19295 10084 19340 10112
rect 19334 10072 19340 10084
rect 19392 10072 19398 10124
rect 19426 10072 19432 10124
rect 19484 10112 19490 10124
rect 19996 10121 20024 10152
rect 19981 10115 20039 10121
rect 19484 10084 19529 10112
rect 19484 10072 19490 10084
rect 19981 10081 19993 10115
rect 20027 10081 20039 10115
rect 19981 10075 20039 10081
rect 20070 10072 20076 10124
rect 20128 10112 20134 10124
rect 20622 10112 20628 10124
rect 20128 10084 20628 10112
rect 20128 10072 20134 10084
rect 20622 10072 20628 10084
rect 20680 10072 20686 10124
rect 20806 10072 20812 10124
rect 20864 10112 20870 10124
rect 20901 10115 20959 10121
rect 20901 10112 20913 10115
rect 20864 10084 20913 10112
rect 20864 10072 20870 10084
rect 20901 10081 20913 10084
rect 20947 10081 20959 10115
rect 21266 10112 21272 10124
rect 21227 10084 21272 10112
rect 20901 10075 20959 10081
rect 21266 10072 21272 10084
rect 21324 10072 21330 10124
rect 21637 10115 21695 10121
rect 21637 10112 21649 10115
rect 21468 10084 21649 10112
rect 12308 10016 13676 10044
rect 12308 10004 12314 10016
rect 14090 10004 14096 10056
rect 14148 10044 14154 10056
rect 15657 10047 15715 10053
rect 15657 10044 15669 10047
rect 14148 10016 15669 10044
rect 14148 10004 14154 10016
rect 15657 10013 15669 10016
rect 15703 10013 15715 10047
rect 15657 10007 15715 10013
rect 6788 9948 8708 9976
rect 13449 9979 13507 9985
rect 6788 9936 6794 9948
rect 13449 9945 13461 9979
rect 13495 9976 13507 9979
rect 16022 9976 16028 9988
rect 13495 9948 16028 9976
rect 13495 9945 13507 9948
rect 13449 9939 13507 9945
rect 16022 9936 16028 9948
rect 16080 9936 16086 9988
rect 5261 9911 5319 9917
rect 5261 9908 5273 9911
rect 1452 9880 5273 9908
rect 1452 9868 1458 9880
rect 5261 9877 5273 9880
rect 5307 9877 5319 9911
rect 9306 9908 9312 9920
rect 9267 9880 9312 9908
rect 5261 9871 5319 9877
rect 9306 9868 9312 9880
rect 9364 9868 9370 9920
rect 11609 9911 11667 9917
rect 11609 9877 11621 9911
rect 11655 9908 11667 9911
rect 11698 9908 11704 9920
rect 11655 9880 11704 9908
rect 11655 9877 11667 9880
rect 11609 9871 11667 9877
rect 11698 9868 11704 9880
rect 11756 9868 11762 9920
rect 17420 9908 17448 10072
rect 17773 10047 17831 10053
rect 17773 10013 17785 10047
rect 17819 10013 17831 10047
rect 19058 10044 19064 10056
rect 19019 10016 19064 10044
rect 17773 10007 17831 10013
rect 17788 9976 17816 10007
rect 19058 10004 19064 10016
rect 19116 10004 19122 10056
rect 19242 10004 19248 10056
rect 19300 10044 19306 10056
rect 20530 10044 20536 10056
rect 19300 10016 20536 10044
rect 19300 10004 19306 10016
rect 20530 10004 20536 10016
rect 20588 10044 20594 10056
rect 21468 10044 21496 10084
rect 21637 10081 21649 10084
rect 21683 10081 21695 10115
rect 21637 10075 21695 10081
rect 22278 10072 22284 10124
rect 22336 10112 22342 10124
rect 22554 10112 22560 10124
rect 22336 10084 22560 10112
rect 22336 10072 22342 10084
rect 22554 10072 22560 10084
rect 22612 10072 22618 10124
rect 21726 10044 21732 10056
rect 20588 10016 21496 10044
rect 21687 10016 21732 10044
rect 20588 10004 20594 10016
rect 21726 10004 21732 10016
rect 21784 10004 21790 10056
rect 20254 9976 20260 9988
rect 17788 9948 20260 9976
rect 20254 9936 20260 9948
rect 20312 9936 20318 9988
rect 21082 9936 21088 9988
rect 21140 9976 21146 9988
rect 22002 9976 22008 9988
rect 21140 9948 22008 9976
rect 21140 9936 21146 9948
rect 22002 9936 22008 9948
rect 22060 9976 22066 9988
rect 22756 9976 22784 10220
rect 35802 10208 35808 10220
rect 35860 10208 35866 10260
rect 36630 10208 36636 10260
rect 36688 10248 36694 10260
rect 37829 10251 37887 10257
rect 37829 10248 37841 10251
rect 36688 10220 37841 10248
rect 36688 10208 36694 10220
rect 37829 10217 37841 10220
rect 37875 10217 37887 10251
rect 37829 10211 37887 10217
rect 27062 10140 27068 10192
rect 27120 10180 27126 10192
rect 27120 10152 28488 10180
rect 27120 10140 27126 10152
rect 23290 10112 23296 10124
rect 23251 10084 23296 10112
rect 23290 10072 23296 10084
rect 23348 10072 23354 10124
rect 25498 10112 25504 10124
rect 25459 10084 25504 10112
rect 25498 10072 25504 10084
rect 25556 10072 25562 10124
rect 25682 10112 25688 10124
rect 25643 10084 25688 10112
rect 25682 10072 25688 10084
rect 25740 10072 25746 10124
rect 26142 10072 26148 10124
rect 26200 10112 26206 10124
rect 26697 10115 26755 10121
rect 26697 10112 26709 10115
rect 26200 10084 26709 10112
rect 26200 10072 26206 10084
rect 26697 10081 26709 10084
rect 26743 10081 26755 10115
rect 26697 10075 26755 10081
rect 26970 10072 26976 10124
rect 27028 10112 27034 10124
rect 27617 10115 27675 10121
rect 27617 10112 27629 10115
rect 27028 10084 27629 10112
rect 27028 10072 27034 10084
rect 27617 10081 27629 10084
rect 27663 10081 27675 10115
rect 27890 10112 27896 10124
rect 27851 10084 27896 10112
rect 27617 10075 27675 10081
rect 23017 10047 23075 10053
rect 23017 10013 23029 10047
rect 23063 10044 23075 10047
rect 23198 10044 23204 10056
rect 23063 10016 23204 10044
rect 23063 10013 23075 10016
rect 23017 10007 23075 10013
rect 23198 10004 23204 10016
rect 23256 10004 23262 10056
rect 25961 10047 26019 10053
rect 25961 10013 25973 10047
rect 26007 10044 26019 10047
rect 27338 10044 27344 10056
rect 26007 10016 27344 10044
rect 26007 10013 26019 10016
rect 25961 10007 26019 10013
rect 27338 10004 27344 10016
rect 27396 10004 27402 10056
rect 22060 9948 22784 9976
rect 27632 9976 27660 10075
rect 27890 10072 27896 10084
rect 27948 10072 27954 10124
rect 27982 10072 27988 10124
rect 28040 10112 28046 10124
rect 28350 10112 28356 10124
rect 28040 10084 28356 10112
rect 28040 10072 28046 10084
rect 28350 10072 28356 10084
rect 28408 10072 28414 10124
rect 27798 10044 27804 10056
rect 27759 10016 27804 10044
rect 27798 10004 27804 10016
rect 27856 10004 27862 10056
rect 28460 10044 28488 10152
rect 28810 10140 28816 10192
rect 28868 10180 28874 10192
rect 28868 10152 30696 10180
rect 28868 10140 28874 10152
rect 28905 10115 28963 10121
rect 28905 10081 28917 10115
rect 28951 10112 28963 10115
rect 28994 10112 29000 10124
rect 28951 10084 29000 10112
rect 28951 10081 28963 10084
rect 28905 10075 28963 10081
rect 28994 10072 29000 10084
rect 29052 10072 29058 10124
rect 29178 10112 29184 10124
rect 29104 10084 29184 10112
rect 29104 10044 29132 10084
rect 29178 10072 29184 10084
rect 29236 10072 29242 10124
rect 29454 10072 29460 10124
rect 29512 10112 29518 10124
rect 30668 10121 30696 10152
rect 31202 10140 31208 10192
rect 31260 10180 31266 10192
rect 31938 10180 31944 10192
rect 31260 10152 31944 10180
rect 31260 10140 31266 10152
rect 31938 10140 31944 10152
rect 31996 10140 32002 10192
rect 33689 10183 33747 10189
rect 33689 10149 33701 10183
rect 33735 10180 33747 10183
rect 34146 10180 34152 10192
rect 33735 10152 34152 10180
rect 33735 10149 33747 10152
rect 33689 10143 33747 10149
rect 34146 10140 34152 10152
rect 34204 10140 34210 10192
rect 30009 10115 30067 10121
rect 30009 10112 30021 10115
rect 29512 10084 30021 10112
rect 29512 10072 29518 10084
rect 30009 10081 30021 10084
rect 30055 10081 30067 10115
rect 30009 10075 30067 10081
rect 30653 10115 30711 10121
rect 30653 10081 30665 10115
rect 30699 10081 30711 10115
rect 31110 10112 31116 10124
rect 31071 10084 31116 10112
rect 30653 10075 30711 10081
rect 31110 10072 31116 10084
rect 31168 10072 31174 10124
rect 32950 10112 32956 10124
rect 32911 10084 32956 10112
rect 32950 10072 32956 10084
rect 33008 10072 33014 10124
rect 33410 10112 33416 10124
rect 33371 10084 33416 10112
rect 33410 10072 33416 10084
rect 33468 10072 33474 10124
rect 33778 10072 33784 10124
rect 33836 10112 33842 10124
rect 34333 10115 34391 10121
rect 34333 10112 34345 10115
rect 33836 10084 34345 10112
rect 33836 10072 33842 10084
rect 34333 10081 34345 10084
rect 34379 10081 34391 10115
rect 34698 10112 34704 10124
rect 34659 10084 34704 10112
rect 34333 10075 34391 10081
rect 34698 10072 34704 10084
rect 34756 10072 34762 10124
rect 36541 10115 36599 10121
rect 36541 10081 36553 10115
rect 36587 10112 36599 10115
rect 36998 10112 37004 10124
rect 36587 10084 37004 10112
rect 36587 10081 36599 10084
rect 36541 10075 36599 10081
rect 36998 10072 37004 10084
rect 37056 10072 37062 10124
rect 37734 10112 37740 10124
rect 37695 10084 37740 10112
rect 37734 10072 37740 10084
rect 37792 10072 37798 10124
rect 28460 10016 29132 10044
rect 30374 10004 30380 10056
rect 30432 10004 30438 10056
rect 30469 10047 30527 10053
rect 30469 10013 30481 10047
rect 30515 10044 30527 10047
rect 30834 10044 30840 10056
rect 30515 10016 30840 10044
rect 30515 10013 30527 10016
rect 30469 10007 30527 10013
rect 30834 10004 30840 10016
rect 30892 10004 30898 10056
rect 31938 10004 31944 10056
rect 31996 10044 32002 10056
rect 32306 10044 32312 10056
rect 31996 10016 32312 10044
rect 31996 10004 32002 10016
rect 32306 10004 32312 10016
rect 32364 10044 32370 10056
rect 32769 10047 32827 10053
rect 32769 10044 32781 10047
rect 32364 10016 32781 10044
rect 32364 10004 32370 10016
rect 32769 10013 32781 10016
rect 32815 10044 32827 10047
rect 33042 10044 33048 10056
rect 32815 10016 33048 10044
rect 32815 10013 32827 10016
rect 32769 10007 32827 10013
rect 33042 10004 33048 10016
rect 33100 10004 33106 10056
rect 34425 10047 34483 10053
rect 34425 10044 34437 10047
rect 34164 10016 34437 10044
rect 27982 9976 27988 9988
rect 27632 9948 27988 9976
rect 22060 9936 22066 9948
rect 27982 9936 27988 9948
rect 28040 9936 28046 9988
rect 29730 9976 29736 9988
rect 28092 9948 29736 9976
rect 19242 9908 19248 9920
rect 17420 9880 19248 9908
rect 19242 9868 19248 9880
rect 19300 9908 19306 9920
rect 20165 9911 20223 9917
rect 20165 9908 20177 9911
rect 19300 9880 20177 9908
rect 19300 9868 19306 9880
rect 20165 9877 20177 9880
rect 20211 9877 20223 9911
rect 20165 9871 20223 9877
rect 22370 9868 22376 9920
rect 22428 9908 22434 9920
rect 22738 9908 22744 9920
rect 22428 9880 22744 9908
rect 22428 9868 22434 9880
rect 22738 9868 22744 9880
rect 22796 9868 22802 9920
rect 23290 9868 23296 9920
rect 23348 9908 23354 9920
rect 24397 9911 24455 9917
rect 24397 9908 24409 9911
rect 23348 9880 24409 9908
rect 23348 9868 23354 9880
rect 24397 9877 24409 9880
rect 24443 9908 24455 9911
rect 24946 9908 24952 9920
rect 24443 9880 24952 9908
rect 24443 9877 24455 9880
rect 24397 9871 24455 9877
rect 24946 9868 24952 9880
rect 25004 9868 25010 9920
rect 26881 9911 26939 9917
rect 26881 9877 26893 9911
rect 26927 9908 26939 9911
rect 27154 9908 27160 9920
rect 26927 9880 27160 9908
rect 26927 9877 26939 9880
rect 26881 9871 26939 9877
rect 27154 9868 27160 9880
rect 27212 9908 27218 9920
rect 28092 9908 28120 9948
rect 29730 9936 29736 9948
rect 29788 9936 29794 9988
rect 30006 9936 30012 9988
rect 30064 9976 30070 9988
rect 30392 9976 30420 10004
rect 30064 9948 30420 9976
rect 31205 9979 31263 9985
rect 30064 9936 30070 9948
rect 31205 9945 31217 9979
rect 31251 9976 31263 9979
rect 32858 9976 32864 9988
rect 31251 9948 32864 9976
rect 31251 9945 31263 9948
rect 31205 9939 31263 9945
rect 32858 9936 32864 9948
rect 32916 9936 32922 9988
rect 34164 9985 34192 10016
rect 34425 10013 34437 10016
rect 34471 10044 34483 10047
rect 34790 10044 34796 10056
rect 34471 10016 34796 10044
rect 34471 10013 34483 10016
rect 34425 10007 34483 10013
rect 34790 10004 34796 10016
rect 34848 10044 34854 10056
rect 35342 10044 35348 10056
rect 34848 10016 35348 10044
rect 34848 10004 34854 10016
rect 35342 10004 35348 10016
rect 35400 10004 35406 10056
rect 35802 10004 35808 10056
rect 35860 10004 35866 10056
rect 34149 9979 34207 9985
rect 34149 9945 34161 9979
rect 34195 9945 34207 9979
rect 35820 9976 35848 10004
rect 36725 9979 36783 9985
rect 36725 9976 36737 9979
rect 35820 9948 36737 9976
rect 34149 9939 34207 9945
rect 36725 9945 36737 9948
rect 36771 9945 36783 9979
rect 36725 9939 36783 9945
rect 27212 9880 28120 9908
rect 27212 9868 27218 9880
rect 28442 9868 28448 9920
rect 28500 9908 28506 9920
rect 28994 9908 29000 9920
rect 28500 9880 29000 9908
rect 28500 9868 28506 9880
rect 28994 9868 29000 9880
rect 29052 9868 29058 9920
rect 29454 9868 29460 9920
rect 29512 9908 29518 9920
rect 29825 9911 29883 9917
rect 29825 9908 29837 9911
rect 29512 9880 29837 9908
rect 29512 9868 29518 9880
rect 29825 9877 29837 9880
rect 29871 9877 29883 9911
rect 29825 9871 29883 9877
rect 30374 9868 30380 9920
rect 30432 9908 30438 9920
rect 31018 9908 31024 9920
rect 30432 9880 31024 9908
rect 30432 9868 30438 9880
rect 31018 9868 31024 9880
rect 31076 9868 31082 9920
rect 31386 9868 31392 9920
rect 31444 9908 31450 9920
rect 32582 9908 32588 9920
rect 31444 9880 32588 9908
rect 31444 9868 31450 9880
rect 32582 9868 32588 9880
rect 32640 9868 32646 9920
rect 33042 9868 33048 9920
rect 33100 9908 33106 9920
rect 35805 9911 35863 9917
rect 35805 9908 35817 9911
rect 33100 9880 35817 9908
rect 33100 9868 33106 9880
rect 35805 9877 35817 9880
rect 35851 9877 35863 9911
rect 35805 9871 35863 9877
rect 1104 9818 38824 9840
rect 1104 9766 4246 9818
rect 4298 9766 4310 9818
rect 4362 9766 4374 9818
rect 4426 9766 4438 9818
rect 4490 9766 34966 9818
rect 35018 9766 35030 9818
rect 35082 9766 35094 9818
rect 35146 9766 35158 9818
rect 35210 9766 38824 9818
rect 1104 9744 38824 9766
rect 2774 9664 2780 9716
rect 2832 9704 2838 9716
rect 2832 9676 2877 9704
rect 2832 9664 2838 9676
rect 7282 9664 7288 9716
rect 7340 9704 7346 9716
rect 14090 9704 14096 9716
rect 7340 9676 14096 9704
rect 7340 9664 7346 9676
rect 14090 9664 14096 9676
rect 14148 9664 14154 9716
rect 15746 9704 15752 9716
rect 15707 9676 15752 9704
rect 15746 9664 15752 9676
rect 15804 9664 15810 9716
rect 20806 9664 20812 9716
rect 20864 9704 20870 9716
rect 22005 9707 22063 9713
rect 22005 9704 22017 9707
rect 20864 9676 22017 9704
rect 20864 9664 20870 9676
rect 22005 9673 22017 9676
rect 22051 9673 22063 9707
rect 23934 9704 23940 9716
rect 22005 9667 22063 9673
rect 22940 9676 23940 9704
rect 7006 9596 7012 9648
rect 7064 9636 7070 9648
rect 7064 9608 7880 9636
rect 7064 9596 7070 9608
rect 1394 9568 1400 9580
rect 1355 9540 1400 9568
rect 1394 9528 1400 9540
rect 1452 9528 1458 9580
rect 6546 9528 6552 9580
rect 6604 9568 6610 9580
rect 6604 9540 7328 9568
rect 6604 9528 6610 9540
rect 1673 9503 1731 9509
rect 1673 9469 1685 9503
rect 1719 9500 1731 9503
rect 1762 9500 1768 9512
rect 1719 9472 1768 9500
rect 1719 9469 1731 9472
rect 1673 9463 1731 9469
rect 1762 9460 1768 9472
rect 1820 9460 1826 9512
rect 2314 9460 2320 9512
rect 2372 9500 2378 9512
rect 3513 9503 3571 9509
rect 3513 9500 3525 9503
rect 2372 9472 3525 9500
rect 2372 9460 2378 9472
rect 3513 9469 3525 9472
rect 3559 9469 3571 9503
rect 3513 9463 3571 9469
rect 4065 9503 4123 9509
rect 4065 9469 4077 9503
rect 4111 9469 4123 9503
rect 4890 9500 4896 9512
rect 4851 9472 4896 9500
rect 4065 9463 4123 9469
rect 4080 9432 4108 9463
rect 4890 9460 4896 9472
rect 4948 9460 4954 9512
rect 5813 9503 5871 9509
rect 5813 9469 5825 9503
rect 5859 9469 5871 9503
rect 5813 9463 5871 9469
rect 6089 9503 6147 9509
rect 6089 9469 6101 9503
rect 6135 9500 6147 9503
rect 6638 9500 6644 9512
rect 6135 9472 6644 9500
rect 6135 9469 6147 9472
rect 6089 9463 6147 9469
rect 5828 9432 5856 9463
rect 6638 9460 6644 9472
rect 6696 9460 6702 9512
rect 7300 9509 7328 9540
rect 7852 9512 7880 9608
rect 7926 9596 7932 9648
rect 7984 9636 7990 9648
rect 11146 9636 11152 9648
rect 7984 9608 9168 9636
rect 11107 9608 11152 9636
rect 7984 9596 7990 9608
rect 9030 9568 9036 9580
rect 8991 9540 9036 9568
rect 9030 9528 9036 9540
rect 9088 9528 9094 9580
rect 6825 9503 6883 9509
rect 6825 9469 6837 9503
rect 6871 9469 6883 9503
rect 6825 9463 6883 9469
rect 7285 9503 7343 9509
rect 7285 9469 7297 9503
rect 7331 9469 7343 9503
rect 7285 9463 7343 9469
rect 6840 9432 6868 9463
rect 7834 9460 7840 9512
rect 7892 9500 7898 9512
rect 8021 9503 8079 9509
rect 8021 9500 8033 9503
rect 7892 9472 8033 9500
rect 7892 9460 7898 9472
rect 8021 9469 8033 9472
rect 8067 9469 8079 9503
rect 8021 9463 8079 9469
rect 8665 9503 8723 9509
rect 8665 9469 8677 9503
rect 8711 9469 8723 9503
rect 8846 9500 8852 9512
rect 8807 9472 8852 9500
rect 8665 9463 8723 9469
rect 8680 9432 8708 9463
rect 8846 9460 8852 9472
rect 8904 9460 8910 9512
rect 9140 9500 9168 9608
rect 11146 9596 11152 9608
rect 11204 9596 11210 9648
rect 12710 9636 12716 9648
rect 11256 9608 12716 9636
rect 10502 9528 10508 9580
rect 10560 9568 10566 9580
rect 11256 9568 11284 9608
rect 12710 9596 12716 9608
rect 12768 9596 12774 9648
rect 13081 9639 13139 9645
rect 13081 9605 13093 9639
rect 13127 9636 13139 9639
rect 13262 9636 13268 9648
rect 13127 9608 13268 9636
rect 13127 9605 13139 9608
rect 13081 9599 13139 9605
rect 13262 9596 13268 9608
rect 13320 9596 13326 9648
rect 16574 9596 16580 9648
rect 16632 9636 16638 9648
rect 20073 9639 20131 9645
rect 16632 9608 18092 9636
rect 16632 9596 16638 9608
rect 12250 9568 12256 9580
rect 10560 9540 11284 9568
rect 11348 9540 12256 9568
rect 10560 9528 10566 9540
rect 11348 9512 11376 9540
rect 12250 9528 12256 9540
rect 12308 9528 12314 9580
rect 14090 9568 14096 9580
rect 13556 9540 14096 9568
rect 9217 9503 9275 9509
rect 9217 9500 9229 9503
rect 9140 9472 9229 9500
rect 9217 9469 9229 9472
rect 9263 9469 9275 9503
rect 9950 9500 9956 9512
rect 9911 9472 9956 9500
rect 9217 9463 9275 9469
rect 9950 9460 9956 9472
rect 10008 9460 10014 9512
rect 11330 9500 11336 9512
rect 11291 9472 11336 9500
rect 11330 9460 11336 9472
rect 11388 9460 11394 9512
rect 11514 9500 11520 9512
rect 11475 9472 11520 9500
rect 11514 9460 11520 9472
rect 11572 9460 11578 9512
rect 11698 9500 11704 9512
rect 11659 9472 11704 9500
rect 11698 9460 11704 9472
rect 11756 9460 11762 9512
rect 12158 9460 12164 9512
rect 12216 9500 12222 9512
rect 13556 9509 13584 9540
rect 14090 9528 14096 9540
rect 14148 9528 14154 9580
rect 17494 9568 17500 9580
rect 14292 9540 17264 9568
rect 17455 9540 17500 9568
rect 12805 9503 12863 9509
rect 12805 9500 12817 9503
rect 12216 9472 12817 9500
rect 12216 9460 12222 9472
rect 12805 9469 12817 9472
rect 12851 9469 12863 9503
rect 12805 9463 12863 9469
rect 13541 9503 13599 9509
rect 13541 9469 13553 9503
rect 13587 9469 13599 9503
rect 13541 9463 13599 9469
rect 13817 9503 13875 9509
rect 13817 9469 13829 9503
rect 13863 9500 13875 9503
rect 14292 9500 14320 9540
rect 13863 9472 14320 9500
rect 14369 9503 14427 9509
rect 13863 9469 13875 9472
rect 13817 9463 13875 9469
rect 14369 9469 14381 9503
rect 14415 9469 14427 9503
rect 14369 9463 14427 9469
rect 12066 9432 12072 9444
rect 4080 9404 5028 9432
rect 5828 9404 8616 9432
rect 8680 9404 12072 9432
rect 3602 9364 3608 9376
rect 3563 9336 3608 9364
rect 3602 9324 3608 9336
rect 3660 9324 3666 9376
rect 5000 9373 5028 9404
rect 4985 9367 5043 9373
rect 4985 9333 4997 9367
rect 5031 9364 5043 9367
rect 5534 9364 5540 9376
rect 5031 9336 5540 9364
rect 5031 9333 5043 9336
rect 4985 9327 5043 9333
rect 5534 9324 5540 9336
rect 5592 9324 5598 9376
rect 5810 9364 5816 9376
rect 5771 9336 5816 9364
rect 5810 9324 5816 9336
rect 5868 9324 5874 9376
rect 7098 9364 7104 9376
rect 7059 9336 7104 9364
rect 7098 9324 7104 9336
rect 7156 9324 7162 9376
rect 8588 9364 8616 9404
rect 12066 9392 12072 9404
rect 12124 9392 12130 9444
rect 14384 9432 14412 9463
rect 14458 9460 14464 9512
rect 14516 9500 14522 9512
rect 14645 9503 14703 9509
rect 14645 9500 14657 9503
rect 14516 9472 14657 9500
rect 14516 9460 14522 9472
rect 14645 9469 14657 9472
rect 14691 9469 14703 9503
rect 14645 9463 14703 9469
rect 16761 9503 16819 9509
rect 16761 9469 16773 9503
rect 16807 9469 16819 9503
rect 16761 9463 16819 9469
rect 12176 9404 14412 9432
rect 9490 9364 9496 9376
rect 8588 9336 9496 9364
rect 9490 9324 9496 9336
rect 9548 9324 9554 9376
rect 10410 9324 10416 9376
rect 10468 9364 10474 9376
rect 12176 9364 12204 9404
rect 10468 9336 12204 9364
rect 10468 9324 10474 9336
rect 12618 9324 12624 9376
rect 12676 9364 12682 9376
rect 13998 9364 14004 9376
rect 12676 9336 14004 9364
rect 12676 9324 12682 9336
rect 13998 9324 14004 9336
rect 14056 9364 14062 9376
rect 16776 9364 16804 9463
rect 17034 9364 17040 9376
rect 14056 9336 17040 9364
rect 14056 9324 14062 9336
rect 17034 9324 17040 9336
rect 17092 9324 17098 9376
rect 17236 9364 17264 9540
rect 17494 9528 17500 9540
rect 17552 9528 17558 9580
rect 18064 9509 18092 9608
rect 20073 9605 20085 9639
rect 20119 9636 20131 9639
rect 20162 9636 20168 9648
rect 20119 9608 20168 9636
rect 20119 9605 20131 9608
rect 20073 9599 20131 9605
rect 20162 9596 20168 9608
rect 20220 9596 20226 9648
rect 21910 9596 21916 9648
rect 21968 9636 21974 9648
rect 22940 9645 22968 9676
rect 23934 9664 23940 9676
rect 23992 9664 23998 9716
rect 25498 9664 25504 9716
rect 25556 9704 25562 9716
rect 32398 9704 32404 9716
rect 25556 9676 32404 9704
rect 25556 9664 25562 9676
rect 32398 9664 32404 9676
rect 32456 9664 32462 9716
rect 22925 9639 22983 9645
rect 22925 9636 22937 9639
rect 21968 9608 22937 9636
rect 21968 9596 21974 9608
rect 22925 9605 22937 9608
rect 22971 9605 22983 9639
rect 25682 9636 25688 9648
rect 22925 9599 22983 9605
rect 23860 9608 25688 9636
rect 19886 9528 19892 9580
rect 19944 9568 19950 9580
rect 22094 9568 22100 9580
rect 19944 9540 22100 9568
rect 19944 9528 19950 9540
rect 22094 9528 22100 9540
rect 22152 9528 22158 9580
rect 23198 9568 23204 9580
rect 22388 9540 23204 9568
rect 17313 9503 17371 9509
rect 17313 9469 17325 9503
rect 17359 9469 17371 9503
rect 17313 9463 17371 9469
rect 18049 9503 18107 9509
rect 18049 9469 18061 9503
rect 18095 9469 18107 9503
rect 18049 9463 18107 9469
rect 17328 9432 17356 9463
rect 18598 9460 18604 9512
rect 18656 9500 18662 9512
rect 18785 9503 18843 9509
rect 18785 9500 18797 9503
rect 18656 9472 18797 9500
rect 18656 9460 18662 9472
rect 18785 9469 18797 9472
rect 18831 9500 18843 9503
rect 18966 9500 18972 9512
rect 18831 9472 18972 9500
rect 18831 9469 18843 9472
rect 18785 9463 18843 9469
rect 18966 9460 18972 9472
rect 19024 9460 19030 9512
rect 19337 9503 19395 9509
rect 19337 9469 19349 9503
rect 19383 9500 19395 9503
rect 19978 9500 19984 9512
rect 19383 9472 19840 9500
rect 19939 9472 19984 9500
rect 19383 9469 19395 9472
rect 19337 9463 19395 9469
rect 19426 9432 19432 9444
rect 17328 9404 19432 9432
rect 19426 9392 19432 9404
rect 19484 9392 19490 9444
rect 17954 9364 17960 9376
rect 17236 9336 17960 9364
rect 17954 9324 17960 9336
rect 18012 9324 18018 9376
rect 18233 9367 18291 9373
rect 18233 9333 18245 9367
rect 18279 9364 18291 9367
rect 18322 9364 18328 9376
rect 18279 9336 18328 9364
rect 18279 9333 18291 9336
rect 18233 9327 18291 9333
rect 18322 9324 18328 9336
rect 18380 9324 18386 9376
rect 18874 9364 18880 9376
rect 18835 9336 18880 9364
rect 18874 9324 18880 9336
rect 18932 9324 18938 9376
rect 19812 9364 19840 9472
rect 19978 9460 19984 9472
rect 20036 9460 20042 9512
rect 20162 9460 20168 9512
rect 20220 9500 20226 9512
rect 20625 9503 20683 9509
rect 20625 9500 20637 9503
rect 20220 9472 20637 9500
rect 20220 9460 20226 9472
rect 20625 9469 20637 9472
rect 20671 9469 20683 9503
rect 20898 9500 20904 9512
rect 20859 9472 20904 9500
rect 20625 9463 20683 9469
rect 20898 9460 20904 9472
rect 20956 9460 20962 9512
rect 21266 9460 21272 9512
rect 21324 9500 21330 9512
rect 21910 9500 21916 9512
rect 21324 9472 21916 9500
rect 21324 9460 21330 9472
rect 21910 9460 21916 9472
rect 21968 9460 21974 9512
rect 22002 9460 22008 9512
rect 22060 9500 22066 9512
rect 22388 9500 22416 9540
rect 23198 9528 23204 9540
rect 23256 9528 23262 9580
rect 22060 9472 22416 9500
rect 22741 9503 22799 9509
rect 22060 9460 22066 9472
rect 22741 9469 22753 9503
rect 22787 9500 22799 9503
rect 22922 9500 22928 9512
rect 22787 9472 22928 9500
rect 22787 9469 22799 9472
rect 22741 9463 22799 9469
rect 22922 9460 22928 9472
rect 22980 9460 22986 9512
rect 23860 9364 23888 9608
rect 25682 9596 25688 9608
rect 25740 9596 25746 9648
rect 29270 9596 29276 9648
rect 29328 9636 29334 9648
rect 30374 9636 30380 9648
rect 29328 9608 30380 9636
rect 29328 9596 29334 9608
rect 30374 9596 30380 9608
rect 30432 9596 30438 9648
rect 31110 9596 31116 9648
rect 31168 9596 31174 9648
rect 34238 9636 34244 9648
rect 34199 9608 34244 9636
rect 34238 9596 34244 9608
rect 34296 9596 34302 9648
rect 26234 9528 26240 9580
rect 26292 9568 26298 9580
rect 30282 9568 30288 9580
rect 26292 9540 27200 9568
rect 26292 9528 26298 9540
rect 23937 9503 23995 9509
rect 23937 9469 23949 9503
rect 23983 9500 23995 9503
rect 24210 9500 24216 9512
rect 23983 9472 24216 9500
rect 23983 9469 23995 9472
rect 23937 9463 23995 9469
rect 24210 9460 24216 9472
rect 24268 9460 24274 9512
rect 25498 9500 25504 9512
rect 25459 9472 25504 9500
rect 25498 9460 25504 9472
rect 25556 9460 25562 9512
rect 25958 9500 25964 9512
rect 25919 9472 25964 9500
rect 25958 9460 25964 9472
rect 26016 9460 26022 9512
rect 27172 9509 27200 9540
rect 27724 9540 30288 9568
rect 26513 9503 26571 9509
rect 26513 9469 26525 9503
rect 26559 9500 26571 9503
rect 26973 9503 27031 9509
rect 26973 9500 26985 9503
rect 26559 9472 26985 9500
rect 26559 9469 26571 9472
rect 26513 9463 26571 9469
rect 26973 9469 26985 9472
rect 27019 9469 27031 9503
rect 26973 9463 27031 9469
rect 27157 9503 27215 9509
rect 27157 9469 27169 9503
rect 27203 9469 27215 9503
rect 27157 9463 27215 9469
rect 27338 9460 27344 9512
rect 27396 9500 27402 9512
rect 27724 9509 27752 9540
rect 30282 9528 30288 9540
rect 30340 9528 30346 9580
rect 30469 9571 30527 9577
rect 30469 9537 30481 9571
rect 30515 9568 30527 9571
rect 31128 9568 31156 9596
rect 37829 9571 37887 9577
rect 37829 9568 37841 9571
rect 30515 9540 31156 9568
rect 31404 9540 32352 9568
rect 30515 9537 30527 9540
rect 30469 9531 30527 9537
rect 27525 9503 27583 9509
rect 27525 9500 27537 9503
rect 27396 9472 27537 9500
rect 27396 9460 27402 9472
rect 27525 9469 27537 9472
rect 27571 9469 27583 9503
rect 27525 9463 27583 9469
rect 27709 9503 27767 9509
rect 27709 9469 27721 9503
rect 27755 9469 27767 9503
rect 27709 9463 27767 9469
rect 27893 9503 27951 9509
rect 27893 9469 27905 9503
rect 27939 9469 27951 9503
rect 28442 9500 28448 9512
rect 28403 9472 28448 9500
rect 27893 9463 27951 9469
rect 26878 9392 26884 9444
rect 26936 9432 26942 9444
rect 27724 9432 27752 9463
rect 26936 9404 27752 9432
rect 26936 9392 26942 9404
rect 24026 9364 24032 9376
rect 19812 9336 23888 9364
rect 23939 9336 24032 9364
rect 24026 9324 24032 9336
rect 24084 9364 24090 9376
rect 27908 9364 27936 9463
rect 28442 9460 28448 9472
rect 28500 9460 28506 9512
rect 29365 9503 29423 9509
rect 29365 9469 29377 9503
rect 29411 9500 29423 9503
rect 29730 9500 29736 9512
rect 29411 9472 29736 9500
rect 29411 9469 29423 9472
rect 29365 9463 29423 9469
rect 29730 9460 29736 9472
rect 29788 9460 29794 9512
rect 30101 9503 30159 9509
rect 30101 9469 30113 9503
rect 30147 9469 30159 9503
rect 30834 9500 30840 9512
rect 30747 9472 30840 9500
rect 30101 9463 30159 9469
rect 27982 9392 27988 9444
rect 28040 9432 28046 9444
rect 30116 9432 30144 9463
rect 30834 9460 30840 9472
rect 30892 9460 30898 9512
rect 31205 9503 31263 9509
rect 31205 9469 31217 9503
rect 31251 9500 31263 9503
rect 31294 9500 31300 9512
rect 31251 9472 31300 9500
rect 31251 9469 31263 9472
rect 31205 9463 31263 9469
rect 31294 9460 31300 9472
rect 31352 9460 31358 9512
rect 28040 9404 30144 9432
rect 30852 9432 30880 9460
rect 31404 9432 31432 9540
rect 32324 9512 32352 9540
rect 35682 9540 37841 9568
rect 35682 9512 35710 9540
rect 37829 9537 37841 9540
rect 37875 9537 37887 9571
rect 37829 9531 37887 9537
rect 31481 9503 31539 9509
rect 31481 9469 31493 9503
rect 31527 9469 31539 9503
rect 31481 9463 31539 9469
rect 32033 9503 32091 9509
rect 32033 9469 32045 9503
rect 32079 9500 32091 9503
rect 32122 9500 32128 9512
rect 32079 9472 32128 9500
rect 32079 9469 32091 9472
rect 32033 9463 32091 9469
rect 30852 9404 31432 9432
rect 28040 9392 28046 9404
rect 24084 9336 27936 9364
rect 24084 9324 24090 9336
rect 28166 9324 28172 9376
rect 28224 9364 28230 9376
rect 29549 9367 29607 9373
rect 29549 9364 29561 9367
rect 28224 9336 29561 9364
rect 28224 9324 28230 9336
rect 29549 9333 29561 9336
rect 29595 9364 29607 9367
rect 31496 9364 31524 9463
rect 32122 9460 32128 9472
rect 32180 9460 32186 9512
rect 32306 9460 32312 9512
rect 32364 9500 32370 9512
rect 32493 9503 32551 9509
rect 32493 9500 32505 9503
rect 32364 9472 32505 9500
rect 32364 9460 32370 9472
rect 32493 9469 32505 9472
rect 32539 9469 32551 9503
rect 32950 9500 32956 9512
rect 32911 9472 32956 9500
rect 32493 9463 32551 9469
rect 32950 9460 32956 9472
rect 33008 9460 33014 9512
rect 33410 9500 33416 9512
rect 33371 9472 33416 9500
rect 33410 9460 33416 9472
rect 33468 9460 33474 9512
rect 34057 9503 34115 9509
rect 34057 9469 34069 9503
rect 34103 9500 34115 9503
rect 34514 9500 34520 9512
rect 34103 9472 34520 9500
rect 34103 9469 34115 9472
rect 34057 9463 34115 9469
rect 34514 9460 34520 9472
rect 34572 9460 34578 9512
rect 35526 9500 35532 9512
rect 35487 9472 35532 9500
rect 35526 9460 35532 9472
rect 35584 9460 35590 9512
rect 35618 9460 35624 9512
rect 35676 9509 35710 9512
rect 35676 9503 35725 9509
rect 35676 9469 35679 9503
rect 35713 9469 35725 9503
rect 35676 9463 35725 9469
rect 35676 9460 35682 9463
rect 35802 9460 35808 9512
rect 35860 9500 35866 9512
rect 35860 9472 35905 9500
rect 35860 9460 35866 9472
rect 35986 9460 35992 9512
rect 36044 9500 36050 9512
rect 36449 9503 36507 9509
rect 36449 9500 36461 9503
rect 36044 9472 36461 9500
rect 36044 9460 36050 9472
rect 36449 9469 36461 9472
rect 36495 9469 36507 9503
rect 36449 9463 36507 9469
rect 36725 9503 36783 9509
rect 36725 9469 36737 9503
rect 36771 9500 36783 9503
rect 38010 9500 38016 9512
rect 36771 9472 38016 9500
rect 36771 9469 36783 9472
rect 36725 9463 36783 9469
rect 38010 9460 38016 9472
rect 38068 9460 38074 9512
rect 32766 9392 32772 9444
rect 32824 9432 32830 9444
rect 33597 9435 33655 9441
rect 33597 9432 33609 9435
rect 32824 9404 33609 9432
rect 32824 9392 32830 9404
rect 33597 9401 33609 9404
rect 33643 9401 33655 9435
rect 33597 9395 33655 9401
rect 34977 9435 35035 9441
rect 34977 9401 34989 9435
rect 35023 9432 35035 9435
rect 35342 9432 35348 9444
rect 35023 9404 35348 9432
rect 35023 9401 35035 9404
rect 34977 9395 35035 9401
rect 35342 9392 35348 9404
rect 35400 9392 35406 9444
rect 29595 9336 31524 9364
rect 29595 9333 29607 9336
rect 29549 9327 29607 9333
rect 31570 9324 31576 9376
rect 31628 9364 31634 9376
rect 36262 9364 36268 9376
rect 31628 9336 36268 9364
rect 31628 9324 31634 9336
rect 36262 9324 36268 9336
rect 36320 9324 36326 9376
rect 1104 9274 38824 9296
rect 1104 9222 19606 9274
rect 19658 9222 19670 9274
rect 19722 9222 19734 9274
rect 19786 9222 19798 9274
rect 19850 9222 38824 9274
rect 1104 9200 38824 9222
rect 8021 9163 8079 9169
rect 8021 9129 8033 9163
rect 8067 9160 8079 9163
rect 8570 9160 8576 9172
rect 8067 9132 8576 9160
rect 8067 9129 8079 9132
rect 8021 9123 8079 9129
rect 8570 9120 8576 9132
rect 8628 9160 8634 9172
rect 9766 9160 9772 9172
rect 8628 9132 9772 9160
rect 8628 9120 8634 9132
rect 9766 9120 9772 9132
rect 9824 9120 9830 9172
rect 15381 9163 15439 9169
rect 11808 9132 14596 9160
rect 3513 9095 3571 9101
rect 3513 9061 3525 9095
rect 3559 9092 3571 9095
rect 4614 9092 4620 9104
rect 3559 9064 4620 9092
rect 3559 9061 3571 9064
rect 3513 9055 3571 9061
rect 4614 9052 4620 9064
rect 4672 9052 4678 9104
rect 4816 9064 8616 9092
rect 1394 8984 1400 9036
rect 1452 9024 1458 9036
rect 4816 9033 4844 9064
rect 1857 9027 1915 9033
rect 1857 9024 1869 9027
rect 1452 8996 1869 9024
rect 1452 8984 1458 8996
rect 1857 8993 1869 8996
rect 1903 8993 1915 9027
rect 1857 8987 1915 8993
rect 4801 9027 4859 9033
rect 4801 8993 4813 9027
rect 4847 8993 4859 9027
rect 4801 8987 4859 8993
rect 5445 9027 5503 9033
rect 5445 8993 5457 9027
rect 5491 8993 5503 9027
rect 5445 8987 5503 8993
rect 2130 8956 2136 8968
rect 2091 8928 2136 8956
rect 2130 8916 2136 8928
rect 2188 8916 2194 8968
rect 5460 8956 5488 8987
rect 5534 8984 5540 9036
rect 5592 9024 5598 9036
rect 5905 9027 5963 9033
rect 5905 9024 5917 9027
rect 5592 8996 5917 9024
rect 5592 8984 5598 8996
rect 5905 8993 5917 8996
rect 5951 8993 5963 9027
rect 6454 9024 6460 9036
rect 6415 8996 6460 9024
rect 5905 8987 5963 8993
rect 6454 8984 6460 8996
rect 6512 8984 6518 9036
rect 6822 9024 6828 9036
rect 6783 8996 6828 9024
rect 6822 8984 6828 8996
rect 6880 8984 6886 9036
rect 7006 8984 7012 9036
rect 7064 9024 7070 9036
rect 7101 9027 7159 9033
rect 7101 9024 7113 9027
rect 7064 8996 7113 9024
rect 7064 8984 7070 8996
rect 7101 8993 7113 8996
rect 7147 8993 7159 9027
rect 7101 8987 7159 8993
rect 8205 9027 8263 9033
rect 8205 8993 8217 9027
rect 8251 9024 8263 9027
rect 8294 9024 8300 9036
rect 8251 8996 8300 9024
rect 8251 8993 8263 8996
rect 8205 8987 8263 8993
rect 8294 8984 8300 8996
rect 8352 8984 8358 9036
rect 5994 8956 6000 8968
rect 5460 8928 6000 8956
rect 5994 8916 6000 8928
rect 6052 8916 6058 8968
rect 4706 8848 4712 8900
rect 4764 8888 4770 8900
rect 5537 8891 5595 8897
rect 5537 8888 5549 8891
rect 4764 8860 5549 8888
rect 4764 8848 4770 8860
rect 5537 8857 5549 8860
rect 5583 8857 5595 8891
rect 5537 8851 5595 8857
rect 4893 8823 4951 8829
rect 4893 8789 4905 8823
rect 4939 8820 4951 8823
rect 7374 8820 7380 8832
rect 4939 8792 7380 8820
rect 4939 8789 4951 8792
rect 4893 8783 4951 8789
rect 7374 8780 7380 8792
rect 7432 8780 7438 8832
rect 8588 8820 8616 9064
rect 9674 9052 9680 9104
rect 9732 9092 9738 9104
rect 9953 9095 10011 9101
rect 9953 9092 9965 9095
rect 9732 9064 9965 9092
rect 9732 9052 9738 9064
rect 9953 9061 9965 9064
rect 9999 9061 10011 9095
rect 9953 9055 10011 9061
rect 10428 9064 11652 9092
rect 8665 9027 8723 9033
rect 8665 8993 8677 9027
rect 8711 8993 8723 9027
rect 8665 8987 8723 8993
rect 9033 9027 9091 9033
rect 9033 8993 9045 9027
rect 9079 9024 9091 9027
rect 9214 9024 9220 9036
rect 9079 8996 9220 9024
rect 9079 8993 9091 8996
rect 9033 8987 9091 8993
rect 8680 8888 8708 8987
rect 9214 8984 9220 8996
rect 9272 8984 9278 9036
rect 9490 8984 9496 9036
rect 9548 9024 9554 9036
rect 10428 9024 10456 9064
rect 10594 9024 10600 9036
rect 9548 8996 10456 9024
rect 10555 8996 10600 9024
rect 9548 8984 9554 8996
rect 10594 8984 10600 8996
rect 10652 8984 10658 9036
rect 10778 8984 10784 9036
rect 10836 9024 10842 9036
rect 11624 9033 11652 9064
rect 10965 9027 11023 9033
rect 10965 9024 10977 9027
rect 10836 8996 10977 9024
rect 10836 8984 10842 8996
rect 10965 8993 10977 8996
rect 11011 9024 11023 9027
rect 11609 9027 11667 9033
rect 11011 8996 11192 9024
rect 11011 8993 11023 8996
rect 10965 8987 11023 8993
rect 8757 8959 8815 8965
rect 8757 8925 8769 8959
rect 8803 8956 8815 8959
rect 9122 8956 9128 8968
rect 8803 8928 9128 8956
rect 8803 8925 8815 8928
rect 8757 8919 8815 8925
rect 9122 8916 9128 8928
rect 9180 8916 9186 8968
rect 10318 8916 10324 8968
rect 10376 8956 10382 8968
rect 10505 8959 10563 8965
rect 10505 8956 10517 8959
rect 10376 8928 10517 8956
rect 10376 8916 10382 8928
rect 10505 8925 10517 8928
rect 10551 8925 10563 8959
rect 10505 8919 10563 8925
rect 11057 8959 11115 8965
rect 11057 8925 11069 8959
rect 11103 8925 11115 8959
rect 11164 8956 11192 8996
rect 11609 8993 11621 9027
rect 11655 8993 11667 9027
rect 11609 8987 11667 8993
rect 11808 8956 11836 9132
rect 12345 9095 12403 9101
rect 12345 9061 12357 9095
rect 12391 9092 12403 9095
rect 14458 9092 14464 9104
rect 12391 9064 14464 9092
rect 12391 9061 12403 9064
rect 12345 9055 12403 9061
rect 14458 9052 14464 9064
rect 14516 9052 14522 9104
rect 12066 9024 12072 9036
rect 12027 8996 12072 9024
rect 12066 8984 12072 8996
rect 12124 8984 12130 9036
rect 13541 9027 13599 9033
rect 13541 8993 13553 9027
rect 13587 9024 13599 9027
rect 13906 9024 13912 9036
rect 13587 8996 13768 9024
rect 13867 8996 13912 9024
rect 13587 8993 13599 8996
rect 13541 8987 13599 8993
rect 11164 8928 11836 8956
rect 11057 8919 11115 8925
rect 9766 8888 9772 8900
rect 8680 8860 9772 8888
rect 9766 8848 9772 8860
rect 9824 8848 9830 8900
rect 8662 8820 8668 8832
rect 8588 8792 8668 8820
rect 8662 8780 8668 8792
rect 8720 8780 8726 8832
rect 11072 8820 11100 8919
rect 12084 8888 12112 8984
rect 12158 8916 12164 8968
rect 12216 8956 12222 8968
rect 13446 8956 13452 8968
rect 12216 8928 13452 8956
rect 12216 8916 12222 8928
rect 13446 8916 13452 8928
rect 13504 8916 13510 8968
rect 13740 8956 13768 8996
rect 13906 8984 13912 8996
rect 13964 8984 13970 9036
rect 13998 8984 14004 9036
rect 14056 9024 14062 9036
rect 14568 9033 14596 9132
rect 15381 9129 15393 9163
rect 15427 9160 15439 9163
rect 15654 9160 15660 9172
rect 15427 9132 15660 9160
rect 15427 9129 15439 9132
rect 15381 9123 15439 9129
rect 15654 9120 15660 9132
rect 15712 9120 15718 9172
rect 17034 9160 17040 9172
rect 16995 9132 17040 9160
rect 17034 9120 17040 9132
rect 17092 9120 17098 9172
rect 19978 9120 19984 9172
rect 20036 9160 20042 9172
rect 21082 9160 21088 9172
rect 20036 9132 21088 9160
rect 20036 9120 20042 9132
rect 21082 9120 21088 9132
rect 21140 9120 21146 9172
rect 22830 9120 22836 9172
rect 22888 9160 22894 9172
rect 24581 9163 24639 9169
rect 24581 9160 24593 9163
rect 22888 9132 24593 9160
rect 22888 9120 22894 9132
rect 24581 9129 24593 9132
rect 24627 9129 24639 9163
rect 24581 9123 24639 9129
rect 25869 9163 25927 9169
rect 25869 9129 25881 9163
rect 25915 9160 25927 9163
rect 27062 9160 27068 9172
rect 25915 9132 27068 9160
rect 25915 9129 25927 9132
rect 25869 9123 25927 9129
rect 27062 9120 27068 9132
rect 27120 9120 27126 9172
rect 28350 9120 28356 9172
rect 28408 9160 28414 9172
rect 28408 9132 28764 9160
rect 28408 9120 28414 9132
rect 19153 9095 19211 9101
rect 19153 9092 19165 9095
rect 16316 9064 19165 9092
rect 14553 9027 14611 9033
rect 14056 8996 14101 9024
rect 14056 8984 14062 8996
rect 14553 8993 14565 9027
rect 14599 8993 14611 9027
rect 15470 9024 15476 9036
rect 15431 8996 15476 9024
rect 14553 8987 14611 8993
rect 15470 8984 15476 8996
rect 15528 8984 15534 9036
rect 15838 9024 15844 9036
rect 15799 8996 15844 9024
rect 15838 8984 15844 8996
rect 15896 8984 15902 9036
rect 16316 9033 16344 9064
rect 19153 9061 19165 9064
rect 19199 9061 19211 9095
rect 19153 9055 19211 9061
rect 20622 9052 20628 9104
rect 20680 9092 20686 9104
rect 22278 9092 22284 9104
rect 20680 9064 22284 9092
rect 20680 9052 20686 9064
rect 22278 9052 22284 9064
rect 22336 9052 22342 9104
rect 27080 9092 27108 9120
rect 28736 9092 28764 9132
rect 28810 9120 28816 9172
rect 28868 9160 28874 9172
rect 28868 9132 30512 9160
rect 28868 9120 28874 9132
rect 27080 9064 28672 9092
rect 28736 9064 29684 9092
rect 16301 9027 16359 9033
rect 16301 8993 16313 9027
rect 16347 8993 16359 9027
rect 16301 8987 16359 8993
rect 16574 8984 16580 9036
rect 16632 9024 16638 9036
rect 16853 9027 16911 9033
rect 16853 9024 16865 9027
rect 16632 8996 16865 9024
rect 16632 8984 16638 8996
rect 16853 8993 16865 8996
rect 16899 8993 16911 9027
rect 16853 8987 16911 8993
rect 17034 8984 17040 9036
rect 17092 9024 17098 9036
rect 17773 9027 17831 9033
rect 17773 9024 17785 9027
rect 17092 8996 17785 9024
rect 17092 8984 17098 8996
rect 17773 8993 17785 8996
rect 17819 8993 17831 9027
rect 17773 8987 17831 8993
rect 18325 9027 18383 9033
rect 18325 8993 18337 9027
rect 18371 9024 18383 9027
rect 18371 8996 19012 9024
rect 18371 8993 18383 8996
rect 18325 8987 18383 8993
rect 13814 8956 13820 8968
rect 13740 8928 13820 8956
rect 13814 8916 13820 8928
rect 13872 8916 13878 8968
rect 18414 8956 18420 8968
rect 18375 8928 18420 8956
rect 18414 8916 18420 8928
rect 18472 8916 18478 8968
rect 14645 8891 14703 8897
rect 14645 8888 14657 8891
rect 12084 8860 14657 8888
rect 14645 8857 14657 8860
rect 14691 8857 14703 8891
rect 18984 8888 19012 8996
rect 19058 8984 19064 9036
rect 19116 9024 19122 9036
rect 19797 9027 19855 9033
rect 19797 9024 19809 9027
rect 19116 8996 19809 9024
rect 19116 8984 19122 8996
rect 19797 8993 19809 8996
rect 19843 8993 19855 9027
rect 19797 8987 19855 8993
rect 20165 9027 20223 9033
rect 20165 8993 20177 9027
rect 20211 9024 20223 9027
rect 20806 9024 20812 9036
rect 20211 8996 20812 9024
rect 20211 8993 20223 8996
rect 20165 8987 20223 8993
rect 20806 8984 20812 8996
rect 20864 8984 20870 9036
rect 21453 9027 21511 9033
rect 21453 8993 21465 9027
rect 21499 8993 21511 9027
rect 21726 9024 21732 9036
rect 21687 8996 21732 9024
rect 21453 8987 21511 8993
rect 19242 8916 19248 8968
rect 19300 8956 19306 8968
rect 19705 8959 19763 8965
rect 19705 8956 19717 8959
rect 19300 8928 19717 8956
rect 19300 8916 19306 8928
rect 19705 8925 19717 8928
rect 19751 8925 19763 8959
rect 20254 8956 20260 8968
rect 20215 8928 20260 8956
rect 19705 8919 19763 8925
rect 20254 8916 20260 8928
rect 20312 8916 20318 8968
rect 20993 8959 21051 8965
rect 20993 8956 21005 8959
rect 20732 8928 21005 8956
rect 19886 8888 19892 8900
rect 18984 8860 19892 8888
rect 14645 8851 14703 8857
rect 19886 8848 19892 8860
rect 19944 8848 19950 8900
rect 20346 8848 20352 8900
rect 20404 8888 20410 8900
rect 20732 8888 20760 8928
rect 20993 8925 21005 8928
rect 21039 8925 21051 8959
rect 21468 8956 21496 8987
rect 21726 8984 21732 8996
rect 21784 8984 21790 9036
rect 21818 8984 21824 9036
rect 21876 9024 21882 9036
rect 22465 9027 22523 9033
rect 22465 9024 22477 9027
rect 21876 8996 22477 9024
rect 21876 8984 21882 8996
rect 22465 8993 22477 8996
rect 22511 8993 22523 9027
rect 22465 8987 22523 8993
rect 25685 9027 25743 9033
rect 25685 8993 25697 9027
rect 25731 9024 25743 9027
rect 26878 9024 26884 9036
rect 25731 8996 26884 9024
rect 25731 8993 25743 8996
rect 25685 8987 25743 8993
rect 26878 8984 26884 8996
rect 26936 8984 26942 9036
rect 27522 9024 27528 9036
rect 27483 8996 27528 9024
rect 27522 8984 27528 8996
rect 27580 8984 27586 9036
rect 27798 8984 27804 9036
rect 27856 9024 27862 9036
rect 28644 9033 28672 9064
rect 27893 9027 27951 9033
rect 27893 9024 27905 9027
rect 27856 8996 27905 9024
rect 27856 8984 27862 8996
rect 27893 8993 27905 8996
rect 27939 8993 27951 9027
rect 27893 8987 27951 8993
rect 28629 9027 28687 9033
rect 28629 8993 28641 9027
rect 28675 8993 28687 9027
rect 29178 9024 29184 9036
rect 29139 8996 29184 9024
rect 28629 8987 28687 8993
rect 29178 8984 29184 8996
rect 29236 8984 29242 9036
rect 29656 9033 29684 9064
rect 29641 9027 29699 9033
rect 29641 8993 29653 9027
rect 29687 9024 29699 9027
rect 29730 9024 29736 9036
rect 29687 8996 29736 9024
rect 29687 8993 29699 8996
rect 29641 8987 29699 8993
rect 29730 8984 29736 8996
rect 29788 8984 29794 9036
rect 29917 9027 29975 9033
rect 29917 8993 29929 9027
rect 29963 8993 29975 9027
rect 30484 9024 30512 9132
rect 31294 9120 31300 9172
rect 31352 9160 31358 9172
rect 31662 9160 31668 9172
rect 31352 9132 31668 9160
rect 31352 9120 31358 9132
rect 31662 9120 31668 9132
rect 31720 9120 31726 9172
rect 32398 9120 32404 9172
rect 32456 9160 32462 9172
rect 34149 9163 34207 9169
rect 34149 9160 34161 9163
rect 32456 9132 34161 9160
rect 32456 9120 32462 9132
rect 34149 9129 34161 9132
rect 34195 9129 34207 9163
rect 34149 9123 34207 9129
rect 30561 9095 30619 9101
rect 30561 9061 30573 9095
rect 30607 9092 30619 9095
rect 31570 9092 31576 9104
rect 30607 9064 31576 9092
rect 30607 9061 30619 9064
rect 30561 9055 30619 9061
rect 31570 9052 31576 9064
rect 31628 9052 31634 9104
rect 35345 9095 35403 9101
rect 35345 9061 35357 9095
rect 35391 9092 35403 9095
rect 35434 9092 35440 9104
rect 35391 9064 35440 9092
rect 35391 9061 35403 9064
rect 35345 9055 35403 9061
rect 35434 9052 35440 9064
rect 35492 9052 35498 9104
rect 31386 9024 31392 9036
rect 30484 8996 31392 9024
rect 29917 8987 29975 8993
rect 22278 8956 22284 8968
rect 21468 8928 22284 8956
rect 20993 8919 21051 8925
rect 22278 8916 22284 8928
rect 22336 8916 22342 8968
rect 23198 8956 23204 8968
rect 23159 8928 23204 8956
rect 23198 8916 23204 8928
rect 23256 8916 23262 8968
rect 23474 8956 23480 8968
rect 23435 8928 23480 8956
rect 23474 8916 23480 8928
rect 23532 8916 23538 8968
rect 27249 8959 27307 8965
rect 27249 8925 27261 8959
rect 27295 8925 27307 8959
rect 28166 8956 28172 8968
rect 28127 8928 28172 8956
rect 27249 8919 27307 8925
rect 20404 8860 20760 8888
rect 20404 8848 20410 8860
rect 20898 8848 20904 8900
rect 20956 8888 20962 8900
rect 21729 8891 21787 8897
rect 21729 8888 21741 8891
rect 20956 8860 21741 8888
rect 20956 8848 20962 8860
rect 21729 8857 21741 8860
rect 21775 8857 21787 8891
rect 21729 8851 21787 8857
rect 26970 8848 26976 8900
rect 27028 8888 27034 8900
rect 27264 8888 27292 8919
rect 28166 8916 28172 8928
rect 28224 8916 28230 8968
rect 28718 8916 28724 8968
rect 28776 8956 28782 8968
rect 29932 8956 29960 8987
rect 31386 8984 31392 8996
rect 31444 8984 31450 9036
rect 31754 8984 31760 9036
rect 31812 9024 31818 9036
rect 32125 9027 32183 9033
rect 32125 9024 32137 9027
rect 31812 8996 32137 9024
rect 31812 8984 31818 8996
rect 32125 8993 32137 8996
rect 32171 8993 32183 9027
rect 33042 9024 33048 9036
rect 33003 8996 33048 9024
rect 32125 8987 32183 8993
rect 33042 8984 33048 8996
rect 33100 8984 33106 9036
rect 36173 9027 36231 9033
rect 36173 8993 36185 9027
rect 36219 8993 36231 9027
rect 36814 9024 36820 9036
rect 36775 8996 36820 9024
rect 36173 8987 36231 8993
rect 28776 8928 29960 8956
rect 28776 8916 28782 8928
rect 30006 8916 30012 8968
rect 30064 8956 30070 8968
rect 30064 8928 30109 8956
rect 30064 8916 30070 8928
rect 31018 8916 31024 8968
rect 31076 8956 31082 8968
rect 31113 8959 31171 8965
rect 31113 8956 31125 8959
rect 31076 8928 31125 8956
rect 31076 8916 31082 8928
rect 31113 8925 31125 8928
rect 31159 8925 31171 8959
rect 31113 8919 31171 8925
rect 31294 8916 31300 8968
rect 31352 8956 31358 8968
rect 31573 8959 31631 8965
rect 31573 8956 31585 8959
rect 31352 8928 31585 8956
rect 31352 8916 31358 8928
rect 31573 8925 31585 8928
rect 31619 8956 31631 8959
rect 32769 8959 32827 8965
rect 31619 8928 32720 8956
rect 31619 8925 31631 8928
rect 31573 8919 31631 8925
rect 27890 8888 27896 8900
rect 27028 8860 27896 8888
rect 27028 8848 27034 8860
rect 27890 8848 27896 8860
rect 27948 8888 27954 8900
rect 28736 8888 28764 8916
rect 27948 8860 28764 8888
rect 27948 8848 27954 8860
rect 29822 8848 29828 8900
rect 29880 8888 29886 8900
rect 32217 8891 32275 8897
rect 32217 8888 32229 8891
rect 29880 8860 32229 8888
rect 29880 8848 29886 8860
rect 32217 8857 32229 8860
rect 32263 8857 32275 8891
rect 32217 8851 32275 8857
rect 12618 8820 12624 8832
rect 11072 8792 12624 8820
rect 12618 8780 12624 8792
rect 12676 8780 12682 8832
rect 12989 8823 13047 8829
rect 12989 8789 13001 8823
rect 13035 8820 13047 8823
rect 13262 8820 13268 8832
rect 13035 8792 13268 8820
rect 13035 8789 13047 8792
rect 12989 8783 13047 8789
rect 13262 8780 13268 8792
rect 13320 8780 13326 8832
rect 15930 8780 15936 8832
rect 15988 8820 15994 8832
rect 20162 8820 20168 8832
rect 15988 8792 20168 8820
rect 15988 8780 15994 8792
rect 20162 8780 20168 8792
rect 20220 8820 20226 8832
rect 22002 8820 22008 8832
rect 20220 8792 22008 8820
rect 20220 8780 20226 8792
rect 22002 8780 22008 8792
rect 22060 8780 22066 8832
rect 22649 8823 22707 8829
rect 22649 8789 22661 8823
rect 22695 8820 22707 8823
rect 23842 8820 23848 8832
rect 22695 8792 23848 8820
rect 22695 8789 22707 8792
rect 22649 8783 22707 8789
rect 23842 8780 23848 8792
rect 23900 8780 23906 8832
rect 25958 8780 25964 8832
rect 26016 8820 26022 8832
rect 31938 8820 31944 8832
rect 26016 8792 31944 8820
rect 26016 8780 26022 8792
rect 31938 8780 31944 8792
rect 31996 8780 32002 8832
rect 32692 8820 32720 8928
rect 32769 8925 32781 8959
rect 32815 8956 32827 8959
rect 34698 8956 34704 8968
rect 32815 8928 34704 8956
rect 32815 8925 32827 8928
rect 32769 8919 32827 8925
rect 34698 8916 34704 8928
rect 34756 8956 34762 8968
rect 35434 8956 35440 8968
rect 34756 8928 35440 8956
rect 34756 8916 34762 8928
rect 35434 8916 35440 8928
rect 35492 8916 35498 8968
rect 35894 8956 35900 8968
rect 35855 8928 35900 8956
rect 35894 8916 35900 8928
rect 35952 8916 35958 8968
rect 36188 8888 36216 8987
rect 36814 8984 36820 8996
rect 36872 8984 36878 9036
rect 36354 8956 36360 8968
rect 36315 8928 36360 8956
rect 36354 8916 36360 8928
rect 36412 8916 36418 8968
rect 37826 8888 37832 8900
rect 35452 8860 37832 8888
rect 35452 8820 35480 8860
rect 37826 8848 37832 8860
rect 37884 8848 37890 8900
rect 32692 8792 35480 8820
rect 35526 8780 35532 8832
rect 35584 8820 35590 8832
rect 37001 8823 37059 8829
rect 37001 8820 37013 8823
rect 35584 8792 37013 8820
rect 35584 8780 35590 8792
rect 37001 8789 37013 8792
rect 37047 8789 37059 8823
rect 37001 8783 37059 8789
rect 1104 8730 38824 8752
rect 1104 8678 4246 8730
rect 4298 8678 4310 8730
rect 4362 8678 4374 8730
rect 4426 8678 4438 8730
rect 4490 8678 34966 8730
rect 35018 8678 35030 8730
rect 35082 8678 35094 8730
rect 35146 8678 35158 8730
rect 35210 8678 38824 8730
rect 1104 8656 38824 8678
rect 1762 8616 1768 8628
rect 1723 8588 1768 8616
rect 1762 8576 1768 8588
rect 1820 8576 1826 8628
rect 4890 8576 4896 8628
rect 4948 8616 4954 8628
rect 5813 8619 5871 8625
rect 5813 8616 5825 8619
rect 4948 8588 5825 8616
rect 4948 8576 4954 8588
rect 5813 8585 5825 8588
rect 5859 8585 5871 8619
rect 6914 8616 6920 8628
rect 6875 8588 6920 8616
rect 5813 8579 5871 8585
rect 2958 8548 2964 8560
rect 1504 8520 2964 8548
rect 1504 8489 1532 8520
rect 2958 8508 2964 8520
rect 3016 8508 3022 8560
rect 1489 8483 1547 8489
rect 1489 8449 1501 8483
rect 1535 8449 1547 8483
rect 1489 8443 1547 8449
rect 2130 8440 2136 8492
rect 2188 8480 2194 8492
rect 3053 8483 3111 8489
rect 3053 8480 3065 8483
rect 2188 8452 3065 8480
rect 2188 8440 2194 8452
rect 3053 8449 3065 8452
rect 3099 8449 3111 8483
rect 4706 8480 4712 8492
rect 4667 8452 4712 8480
rect 3053 8443 3111 8449
rect 4706 8440 4712 8452
rect 4764 8440 4770 8492
rect 1581 8415 1639 8421
rect 1581 8381 1593 8415
rect 1627 8381 1639 8415
rect 1581 8375 1639 8381
rect 1596 8344 1624 8375
rect 1854 8372 1860 8424
rect 1912 8412 1918 8424
rect 2314 8412 2320 8424
rect 1912 8384 2320 8412
rect 1912 8372 1918 8384
rect 2314 8372 2320 8384
rect 2372 8412 2378 8424
rect 2501 8415 2559 8421
rect 2501 8412 2513 8415
rect 2372 8384 2513 8412
rect 2372 8372 2378 8384
rect 2501 8381 2513 8384
rect 2547 8381 2559 8415
rect 2501 8375 2559 8381
rect 2961 8415 3019 8421
rect 2961 8381 2973 8415
rect 3007 8381 3019 8415
rect 2961 8375 3019 8381
rect 3789 8415 3847 8421
rect 3789 8381 3801 8415
rect 3835 8412 3847 8415
rect 4154 8412 4160 8424
rect 3835 8384 4160 8412
rect 3835 8381 3847 8384
rect 3789 8375 3847 8381
rect 2774 8344 2780 8356
rect 1596 8316 2780 8344
rect 2774 8304 2780 8316
rect 2832 8304 2838 8356
rect 2976 8344 3004 8375
rect 4154 8372 4160 8384
rect 4212 8372 4218 8424
rect 4433 8415 4491 8421
rect 4433 8381 4445 8415
rect 4479 8412 4491 8415
rect 5534 8412 5540 8424
rect 4479 8384 5540 8412
rect 4479 8381 4491 8384
rect 4433 8375 4491 8381
rect 5534 8372 5540 8384
rect 5592 8372 5598 8424
rect 5828 8412 5856 8579
rect 6914 8576 6920 8588
rect 6972 8576 6978 8628
rect 10137 8619 10195 8625
rect 7024 8588 9536 8616
rect 5994 8508 6000 8560
rect 6052 8548 6058 8560
rect 7024 8548 7052 8588
rect 8294 8548 8300 8560
rect 6052 8520 7052 8548
rect 8255 8520 8300 8548
rect 6052 8508 6058 8520
rect 8294 8508 8300 8520
rect 8352 8508 8358 8560
rect 9508 8548 9536 8588
rect 10137 8585 10149 8619
rect 10183 8616 10195 8619
rect 10778 8616 10784 8628
rect 10183 8588 10784 8616
rect 10183 8585 10195 8588
rect 10137 8579 10195 8585
rect 10778 8576 10784 8588
rect 10836 8576 10842 8628
rect 13446 8576 13452 8628
rect 13504 8616 13510 8628
rect 14001 8619 14059 8625
rect 14001 8616 14013 8619
rect 13504 8588 14013 8616
rect 13504 8576 13510 8588
rect 14001 8585 14013 8588
rect 14047 8585 14059 8619
rect 15838 8616 15844 8628
rect 14001 8579 14059 8585
rect 14108 8588 15844 8616
rect 12250 8548 12256 8560
rect 9508 8520 12256 8548
rect 12250 8508 12256 8520
rect 12308 8508 12314 8560
rect 12713 8551 12771 8557
rect 12713 8517 12725 8551
rect 12759 8548 12771 8551
rect 14108 8548 14136 8588
rect 15838 8576 15844 8588
rect 15896 8576 15902 8628
rect 16114 8576 16120 8628
rect 16172 8616 16178 8628
rect 16209 8619 16267 8625
rect 16209 8616 16221 8619
rect 16172 8588 16221 8616
rect 16172 8576 16178 8588
rect 16209 8585 16221 8588
rect 16255 8585 16267 8619
rect 23014 8616 23020 8628
rect 16209 8579 16267 8585
rect 18892 8588 23020 8616
rect 12759 8520 14136 8548
rect 14829 8551 14887 8557
rect 12759 8517 12771 8520
rect 12713 8511 12771 8517
rect 14829 8517 14841 8551
rect 14875 8548 14887 8551
rect 15194 8548 15200 8560
rect 14875 8520 15200 8548
rect 14875 8517 14887 8520
rect 14829 8511 14887 8517
rect 15194 8508 15200 8520
rect 15252 8508 15258 8560
rect 8849 8483 8907 8489
rect 8496 8452 8800 8480
rect 6825 8415 6883 8421
rect 6825 8412 6837 8415
rect 5828 8384 6837 8412
rect 6825 8381 6837 8384
rect 6871 8381 6883 8415
rect 7374 8412 7380 8424
rect 7335 8384 7380 8412
rect 6825 8375 6883 8381
rect 7374 8372 7380 8384
rect 7432 8372 7438 8424
rect 8496 8421 8524 8452
rect 8481 8415 8539 8421
rect 8481 8381 8493 8415
rect 8527 8381 8539 8415
rect 8481 8375 8539 8381
rect 8570 8372 8576 8424
rect 8628 8412 8634 8424
rect 8772 8412 8800 8452
rect 8849 8449 8861 8483
rect 8895 8480 8907 8483
rect 9030 8480 9036 8492
rect 8895 8452 9036 8480
rect 8895 8449 8907 8452
rect 8849 8443 8907 8449
rect 9030 8440 9036 8452
rect 9088 8440 9094 8492
rect 11882 8480 11888 8492
rect 11843 8452 11888 8480
rect 11882 8440 11888 8452
rect 11940 8440 11946 8492
rect 15470 8480 15476 8492
rect 14752 8452 15476 8480
rect 10410 8412 10416 8424
rect 8628 8384 8673 8412
rect 8772 8384 10416 8412
rect 8628 8372 8634 8384
rect 10410 8372 10416 8384
rect 10468 8372 10474 8424
rect 11330 8412 11336 8424
rect 11291 8384 11336 8412
rect 11330 8372 11336 8384
rect 11388 8372 11394 8424
rect 11701 8415 11759 8421
rect 11701 8381 11713 8415
rect 11747 8412 11759 8415
rect 12618 8412 12624 8424
rect 11747 8384 12624 8412
rect 11747 8381 11759 8384
rect 11701 8375 11759 8381
rect 12618 8372 12624 8384
rect 12676 8372 12682 8424
rect 12894 8412 12900 8424
rect 12855 8384 12900 8412
rect 12894 8372 12900 8384
rect 12952 8372 12958 8424
rect 13262 8412 13268 8424
rect 13223 8384 13268 8412
rect 13262 8372 13268 8384
rect 13320 8372 13326 8424
rect 13354 8372 13360 8424
rect 13412 8412 13418 8424
rect 13906 8412 13912 8424
rect 13412 8384 13457 8412
rect 13819 8384 13912 8412
rect 13412 8372 13418 8384
rect 13906 8372 13912 8384
rect 13964 8412 13970 8424
rect 14274 8412 14280 8424
rect 13964 8384 14280 8412
rect 13964 8372 13970 8384
rect 14274 8372 14280 8384
rect 14332 8372 14338 8424
rect 14752 8421 14780 8452
rect 15470 8440 15476 8452
rect 15528 8440 15534 8492
rect 14737 8415 14795 8421
rect 14737 8381 14749 8415
rect 14783 8381 14795 8415
rect 14737 8375 14795 8381
rect 15105 8415 15163 8421
rect 15105 8381 15117 8415
rect 15151 8381 15163 8415
rect 15105 8375 15163 8381
rect 15565 8415 15623 8421
rect 15565 8381 15577 8415
rect 15611 8381 15623 8415
rect 16206 8412 16212 8424
rect 16167 8384 16212 8412
rect 15565 8375 15623 8381
rect 3881 8347 3939 8353
rect 3881 8344 3893 8347
rect 2976 8316 3893 8344
rect 3881 8313 3893 8316
rect 3927 8344 3939 8347
rect 4522 8344 4528 8356
rect 3927 8316 4528 8344
rect 3927 8313 3939 8316
rect 3881 8307 3939 8313
rect 4522 8304 4528 8316
rect 4580 8304 4586 8356
rect 5626 8304 5632 8356
rect 5684 8344 5690 8356
rect 5902 8344 5908 8356
rect 5684 8316 5908 8344
rect 5684 8304 5690 8316
rect 5902 8304 5908 8316
rect 5960 8304 5966 8356
rect 11146 8304 11152 8356
rect 11204 8344 11210 8356
rect 15120 8344 15148 8375
rect 11204 8316 15148 8344
rect 15580 8344 15608 8375
rect 16206 8372 16212 8384
rect 16264 8372 16270 8424
rect 16574 8372 16580 8424
rect 16632 8412 16638 8424
rect 16669 8415 16727 8421
rect 16669 8412 16681 8415
rect 16632 8384 16681 8412
rect 16632 8372 16638 8384
rect 16669 8381 16681 8384
rect 16715 8381 16727 8415
rect 17310 8412 17316 8424
rect 17271 8384 17316 8412
rect 16669 8375 16727 8381
rect 17310 8372 17316 8384
rect 17368 8372 17374 8424
rect 18598 8412 18604 8424
rect 18559 8384 18604 8412
rect 18598 8372 18604 8384
rect 18656 8372 18662 8424
rect 18892 8421 18920 8588
rect 23014 8576 23020 8588
rect 23072 8576 23078 8628
rect 24394 8576 24400 8628
rect 24452 8616 24458 8628
rect 34885 8619 34943 8625
rect 34885 8616 34897 8619
rect 24452 8588 34897 8616
rect 24452 8576 24458 8588
rect 34885 8585 34897 8588
rect 34931 8585 34943 8619
rect 34885 8579 34943 8585
rect 35434 8576 35440 8628
rect 35492 8616 35498 8628
rect 35986 8616 35992 8628
rect 35492 8588 35992 8616
rect 35492 8576 35498 8588
rect 35986 8576 35992 8588
rect 36044 8576 36050 8628
rect 36078 8576 36084 8628
rect 36136 8616 36142 8628
rect 37829 8619 37887 8625
rect 37829 8616 37841 8619
rect 36136 8588 37841 8616
rect 36136 8576 36142 8588
rect 37829 8585 37841 8588
rect 37875 8585 37887 8619
rect 37829 8579 37887 8585
rect 18966 8508 18972 8560
rect 19024 8548 19030 8560
rect 19613 8551 19671 8557
rect 19613 8548 19625 8551
rect 19024 8520 19625 8548
rect 19024 8508 19030 8520
rect 19613 8517 19625 8520
rect 19659 8517 19671 8551
rect 21358 8548 21364 8560
rect 19613 8511 19671 8517
rect 19720 8520 21364 8548
rect 19058 8480 19064 8492
rect 19019 8452 19064 8480
rect 19058 8440 19064 8452
rect 19116 8440 19122 8492
rect 18877 8415 18935 8421
rect 18877 8381 18889 8415
rect 18923 8381 18935 8415
rect 18877 8375 18935 8381
rect 18966 8372 18972 8424
rect 19024 8412 19030 8424
rect 19720 8412 19748 8520
rect 21358 8508 21364 8520
rect 21416 8508 21422 8560
rect 22370 8508 22376 8560
rect 22428 8548 22434 8560
rect 24026 8548 24032 8560
rect 22428 8520 24032 8548
rect 22428 8508 22434 8520
rect 24026 8508 24032 8520
rect 24084 8508 24090 8560
rect 28629 8551 28687 8557
rect 28629 8517 28641 8551
rect 28675 8548 28687 8551
rect 28718 8548 28724 8560
rect 28675 8520 28724 8548
rect 28675 8517 28687 8520
rect 28629 8511 28687 8517
rect 28718 8508 28724 8520
rect 28776 8508 28782 8560
rect 29825 8551 29883 8557
rect 29825 8517 29837 8551
rect 29871 8548 29883 8551
rect 32861 8551 32919 8557
rect 29871 8520 31064 8548
rect 29871 8517 29883 8520
rect 29825 8511 29883 8517
rect 20073 8483 20131 8489
rect 20073 8480 20085 8483
rect 19024 8384 19748 8412
rect 19812 8452 20085 8480
rect 19024 8372 19030 8384
rect 18230 8344 18236 8356
rect 15580 8316 18236 8344
rect 11204 8304 11210 8316
rect 18230 8304 18236 8316
rect 18288 8304 18294 8356
rect 19058 8304 19064 8356
rect 19116 8344 19122 8356
rect 19242 8344 19248 8356
rect 19116 8316 19248 8344
rect 19116 8304 19122 8316
rect 19242 8304 19248 8316
rect 19300 8344 19306 8356
rect 19812 8344 19840 8452
rect 20073 8449 20085 8452
rect 20119 8449 20131 8483
rect 20898 8480 20904 8492
rect 20073 8443 20131 8449
rect 20732 8452 20904 8480
rect 20165 8415 20223 8421
rect 20165 8381 20177 8415
rect 20211 8381 20223 8415
rect 20165 8375 20223 8381
rect 19300 8316 19840 8344
rect 20180 8344 20208 8375
rect 20254 8372 20260 8424
rect 20312 8412 20318 8424
rect 20732 8421 20760 8452
rect 20898 8440 20904 8452
rect 20956 8440 20962 8492
rect 23017 8483 23075 8489
rect 23017 8449 23029 8483
rect 23063 8480 23075 8483
rect 24397 8483 24455 8489
rect 24397 8480 24409 8483
rect 23063 8452 24409 8480
rect 23063 8449 23075 8452
rect 23017 8443 23075 8449
rect 24397 8449 24409 8452
rect 24443 8449 24455 8483
rect 26786 8480 26792 8492
rect 26747 8452 26792 8480
rect 24397 8443 24455 8449
rect 26786 8440 26792 8452
rect 26844 8440 26850 8492
rect 30926 8480 30932 8492
rect 28460 8452 30932 8480
rect 20533 8415 20591 8421
rect 20533 8412 20545 8415
rect 20312 8384 20545 8412
rect 20312 8372 20318 8384
rect 20533 8381 20545 8384
rect 20579 8381 20591 8415
rect 20533 8375 20591 8381
rect 20717 8415 20775 8421
rect 20717 8381 20729 8415
rect 20763 8381 20775 8415
rect 20717 8375 20775 8381
rect 20806 8372 20812 8424
rect 20864 8412 20870 8424
rect 21174 8412 21180 8424
rect 20864 8384 21180 8412
rect 20864 8372 20870 8384
rect 21174 8372 21180 8384
rect 21232 8372 21238 8424
rect 21818 8372 21824 8424
rect 21876 8412 21882 8424
rect 21913 8415 21971 8421
rect 21913 8412 21925 8415
rect 21876 8384 21925 8412
rect 21876 8372 21882 8384
rect 21913 8381 21925 8384
rect 21959 8381 21971 8415
rect 21913 8375 21971 8381
rect 22005 8415 22063 8421
rect 22005 8381 22017 8415
rect 22051 8381 22063 8415
rect 22370 8412 22376 8424
rect 22331 8384 22376 8412
rect 22005 8375 22063 8381
rect 20898 8344 20904 8356
rect 20180 8316 20904 8344
rect 19300 8304 19306 8316
rect 20898 8304 20904 8316
rect 20956 8304 20962 8356
rect 22020 8344 22048 8375
rect 22370 8372 22376 8384
rect 22428 8372 22434 8424
rect 22462 8372 22468 8424
rect 22520 8412 22526 8424
rect 22922 8412 22928 8424
rect 22520 8384 22928 8412
rect 22520 8372 22526 8384
rect 22922 8372 22928 8384
rect 22980 8372 22986 8424
rect 23198 8372 23204 8424
rect 23256 8412 23262 8424
rect 23382 8412 23388 8424
rect 23256 8384 23388 8412
rect 23256 8372 23262 8384
rect 23382 8372 23388 8384
rect 23440 8412 23446 8424
rect 24121 8415 24179 8421
rect 24121 8412 24133 8415
rect 23440 8384 24133 8412
rect 23440 8372 23446 8384
rect 24121 8381 24133 8384
rect 24167 8381 24179 8415
rect 24121 8375 24179 8381
rect 24210 8372 24216 8424
rect 24268 8412 24274 8424
rect 24268 8384 25820 8412
rect 24268 8372 24274 8384
rect 25792 8353 25820 8384
rect 26326 8372 26332 8424
rect 26384 8412 26390 8424
rect 27062 8412 27068 8424
rect 26384 8384 27068 8412
rect 26384 8372 26390 8384
rect 27062 8372 27068 8384
rect 27120 8372 27126 8424
rect 27246 8412 27252 8424
rect 27207 8384 27252 8412
rect 27246 8372 27252 8384
rect 27304 8372 27310 8424
rect 27338 8372 27344 8424
rect 27396 8412 27402 8424
rect 27617 8415 27675 8421
rect 27617 8412 27629 8415
rect 27396 8384 27629 8412
rect 27396 8372 27402 8384
rect 27617 8381 27629 8384
rect 27663 8381 27675 8415
rect 27617 8375 27675 8381
rect 27801 8415 27859 8421
rect 27801 8381 27813 8415
rect 27847 8412 27859 8415
rect 27890 8412 27896 8424
rect 27847 8384 27896 8412
rect 27847 8381 27859 8384
rect 27801 8375 27859 8381
rect 27890 8372 27896 8384
rect 27948 8412 27954 8424
rect 28460 8421 28488 8452
rect 30926 8440 30932 8452
rect 30984 8440 30990 8492
rect 31036 8480 31064 8520
rect 32861 8517 32873 8551
rect 32907 8548 32919 8551
rect 33042 8548 33048 8560
rect 32907 8520 33048 8548
rect 32907 8517 32919 8520
rect 32861 8511 32919 8517
rect 33042 8508 33048 8520
rect 33100 8508 33106 8560
rect 34330 8508 34336 8560
rect 34388 8548 34394 8560
rect 34388 8520 36032 8548
rect 34388 8508 34394 8520
rect 34977 8483 35035 8489
rect 31036 8452 31616 8480
rect 28445 8415 28503 8421
rect 27948 8384 28396 8412
rect 27948 8372 27954 8384
rect 25777 8347 25835 8353
rect 22020 8316 24256 8344
rect 9214 8236 9220 8288
rect 9272 8276 9278 8288
rect 15838 8276 15844 8288
rect 9272 8248 15844 8276
rect 9272 8236 9278 8248
rect 15838 8236 15844 8248
rect 15896 8276 15902 8288
rect 16482 8276 16488 8288
rect 15896 8248 16488 8276
rect 15896 8236 15902 8248
rect 16482 8236 16488 8248
rect 16540 8236 16546 8288
rect 16942 8236 16948 8288
rect 17000 8276 17006 8288
rect 17405 8279 17463 8285
rect 17405 8276 17417 8279
rect 17000 8248 17417 8276
rect 17000 8236 17006 8248
rect 17405 8245 17417 8248
rect 17451 8245 17463 8279
rect 17405 8239 17463 8245
rect 17494 8236 17500 8288
rect 17552 8276 17558 8288
rect 21082 8276 21088 8288
rect 17552 8248 21088 8276
rect 17552 8236 17558 8248
rect 21082 8236 21088 8248
rect 21140 8236 21146 8288
rect 24228 8276 24256 8316
rect 25777 8313 25789 8347
rect 25823 8344 25835 8347
rect 27982 8344 27988 8356
rect 25823 8316 27988 8344
rect 25823 8313 25835 8316
rect 25777 8307 25835 8313
rect 27982 8304 27988 8316
rect 28040 8304 28046 8356
rect 24394 8276 24400 8288
rect 24228 8248 24400 8276
rect 24394 8236 24400 8248
rect 24452 8236 24458 8288
rect 28368 8276 28396 8384
rect 28445 8381 28457 8415
rect 28491 8381 28503 8415
rect 28445 8375 28503 8381
rect 30009 8415 30067 8421
rect 30009 8381 30021 8415
rect 30055 8412 30067 8415
rect 30190 8412 30196 8424
rect 30055 8384 30196 8412
rect 30055 8381 30067 8384
rect 30009 8375 30067 8381
rect 30190 8372 30196 8384
rect 30248 8372 30254 8424
rect 30377 8415 30435 8421
rect 30377 8381 30389 8415
rect 30423 8381 30435 8415
rect 30377 8375 30435 8381
rect 30392 8344 30420 8375
rect 30466 8372 30472 8424
rect 30524 8412 30530 8424
rect 31018 8412 31024 8424
rect 30524 8384 30569 8412
rect 30979 8384 31024 8412
rect 30524 8372 30530 8384
rect 31018 8372 31024 8384
rect 31076 8372 31082 8424
rect 31588 8421 31616 8452
rect 34977 8449 34989 8483
rect 35023 8480 35035 8483
rect 35894 8480 35900 8492
rect 35023 8452 35900 8480
rect 35023 8449 35035 8452
rect 34977 8443 35035 8449
rect 35894 8440 35900 8452
rect 35952 8440 35958 8492
rect 36004 8480 36032 8520
rect 36725 8483 36783 8489
rect 36725 8480 36737 8483
rect 36004 8452 36737 8480
rect 36725 8449 36737 8452
rect 36771 8449 36783 8483
rect 36725 8443 36783 8449
rect 31573 8415 31631 8421
rect 31573 8381 31585 8415
rect 31619 8381 31631 8415
rect 31573 8375 31631 8381
rect 32033 8415 32091 8421
rect 32033 8381 32045 8415
rect 32079 8412 32091 8415
rect 32490 8412 32496 8424
rect 32079 8384 32496 8412
rect 32079 8381 32091 8384
rect 32033 8375 32091 8381
rect 32490 8372 32496 8384
rect 32548 8372 32554 8424
rect 32766 8412 32772 8424
rect 32727 8384 32772 8412
rect 32766 8372 32772 8384
rect 32824 8372 32830 8424
rect 32858 8372 32864 8424
rect 32916 8412 32922 8424
rect 33137 8415 33195 8421
rect 33137 8412 33149 8415
rect 32916 8384 33149 8412
rect 32916 8372 32922 8384
rect 33137 8381 33149 8384
rect 33183 8381 33195 8415
rect 33410 8412 33416 8424
rect 33371 8384 33416 8412
rect 33137 8375 33195 8381
rect 33410 8372 33416 8384
rect 33468 8372 33474 8424
rect 34146 8412 34152 8424
rect 34107 8384 34152 8412
rect 34146 8372 34152 8384
rect 34204 8372 34210 8424
rect 35526 8412 35532 8424
rect 35487 8384 35532 8412
rect 35526 8372 35532 8384
rect 35584 8372 35590 8424
rect 35618 8372 35624 8424
rect 35676 8421 35682 8424
rect 35676 8415 35725 8421
rect 35676 8381 35679 8415
rect 35713 8381 35725 8415
rect 35676 8375 35725 8381
rect 35805 8415 35863 8421
rect 35805 8381 35817 8415
rect 35851 8381 35863 8415
rect 35805 8375 35863 8381
rect 35676 8372 35682 8375
rect 34241 8347 34299 8353
rect 34241 8344 34253 8347
rect 30392 8316 34253 8344
rect 34241 8313 34253 8316
rect 34287 8313 34299 8347
rect 34241 8307 34299 8313
rect 34885 8347 34943 8353
rect 34885 8313 34897 8347
rect 34931 8344 34943 8347
rect 35250 8344 35256 8356
rect 34931 8316 35256 8344
rect 34931 8313 34943 8316
rect 34885 8307 34943 8313
rect 35250 8304 35256 8316
rect 35308 8344 35314 8356
rect 35820 8344 35848 8375
rect 35986 8372 35992 8424
rect 36044 8412 36050 8424
rect 36262 8412 36268 8424
rect 36044 8384 36268 8412
rect 36044 8372 36050 8384
rect 36262 8372 36268 8384
rect 36320 8412 36326 8424
rect 36449 8415 36507 8421
rect 36449 8412 36461 8415
rect 36320 8384 36461 8412
rect 36320 8372 36326 8384
rect 36449 8381 36461 8384
rect 36495 8381 36507 8415
rect 36449 8375 36507 8381
rect 35308 8316 35848 8344
rect 35308 8304 35314 8316
rect 30650 8276 30656 8288
rect 28368 8248 30656 8276
rect 30650 8236 30656 8248
rect 30708 8236 30714 8288
rect 31110 8276 31116 8288
rect 31071 8248 31116 8276
rect 31110 8236 31116 8248
rect 31168 8236 31174 8288
rect 1104 8186 38824 8208
rect 1104 8134 19606 8186
rect 19658 8134 19670 8186
rect 19722 8134 19734 8186
rect 19786 8134 19798 8186
rect 19850 8134 38824 8186
rect 1104 8112 38824 8134
rect 2774 8032 2780 8084
rect 2832 8072 2838 8084
rect 7834 8072 7840 8084
rect 2832 8044 2877 8072
rect 6656 8044 7840 8072
rect 2832 8032 2838 8044
rect 6656 8004 6684 8044
rect 7834 8032 7840 8044
rect 7892 8032 7898 8084
rect 8386 8032 8392 8084
rect 8444 8072 8450 8084
rect 8941 8075 8999 8081
rect 8941 8072 8953 8075
rect 8444 8044 8953 8072
rect 8444 8032 8450 8044
rect 8941 8041 8953 8044
rect 8987 8072 8999 8075
rect 9493 8075 9551 8081
rect 9493 8072 9505 8075
rect 8987 8044 9505 8072
rect 8987 8041 8999 8044
rect 8941 8035 8999 8041
rect 9493 8041 9505 8044
rect 9539 8041 9551 8075
rect 9493 8035 9551 8041
rect 11701 8075 11759 8081
rect 11701 8041 11713 8075
rect 11747 8072 11759 8075
rect 11790 8072 11796 8084
rect 11747 8044 11796 8072
rect 11747 8041 11759 8044
rect 11701 8035 11759 8041
rect 11790 8032 11796 8044
rect 11848 8032 11854 8084
rect 13814 8032 13820 8084
rect 13872 8072 13878 8084
rect 14093 8075 14151 8081
rect 14093 8072 14105 8075
rect 13872 8044 14105 8072
rect 13872 8032 13878 8044
rect 14093 8041 14105 8044
rect 14139 8041 14151 8075
rect 14093 8035 14151 8041
rect 15194 8032 15200 8084
rect 15252 8072 15258 8084
rect 15746 8072 15752 8084
rect 15252 8044 15752 8072
rect 15252 8032 15258 8044
rect 15746 8032 15752 8044
rect 15804 8032 15810 8084
rect 16022 8032 16028 8084
rect 16080 8072 16086 8084
rect 20073 8075 20131 8081
rect 16080 8044 18368 8072
rect 16080 8032 16086 8044
rect 9398 8004 9404 8016
rect 6564 7976 6684 8004
rect 6932 7976 9404 8004
rect 1394 7936 1400 7948
rect 1355 7908 1400 7936
rect 1394 7896 1400 7908
rect 1452 7896 1458 7948
rect 4154 7896 4160 7948
rect 4212 7936 4218 7948
rect 4525 7939 4583 7945
rect 4525 7936 4537 7939
rect 4212 7908 4537 7936
rect 4212 7896 4218 7908
rect 4525 7905 4537 7908
rect 4571 7936 4583 7939
rect 4614 7936 4620 7948
rect 4571 7908 4620 7936
rect 4571 7905 4583 7908
rect 4525 7899 4583 7905
rect 4614 7896 4620 7908
rect 4672 7896 4678 7948
rect 4982 7936 4988 7948
rect 4943 7908 4988 7936
rect 4982 7896 4988 7908
rect 5040 7896 5046 7948
rect 5629 7939 5687 7945
rect 5629 7905 5641 7939
rect 5675 7936 5687 7939
rect 6086 7936 6092 7948
rect 5675 7908 6092 7936
rect 5675 7905 5687 7908
rect 5629 7899 5687 7905
rect 6086 7896 6092 7908
rect 6144 7896 6150 7948
rect 6564 7945 6592 7976
rect 6549 7939 6607 7945
rect 6549 7905 6561 7939
rect 6595 7905 6607 7939
rect 6549 7899 6607 7905
rect 6638 7896 6644 7948
rect 6696 7936 6702 7948
rect 6932 7945 6960 7976
rect 9398 7964 9404 7976
rect 9456 7964 9462 8016
rect 18230 8004 18236 8016
rect 10520 7976 18092 8004
rect 18191 7976 18236 8004
rect 6917 7939 6975 7945
rect 6917 7936 6929 7939
rect 6696 7908 6929 7936
rect 6696 7896 6702 7908
rect 6917 7905 6929 7908
rect 6963 7905 6975 7939
rect 6917 7899 6975 7905
rect 7285 7939 7343 7945
rect 7285 7905 7297 7939
rect 7331 7905 7343 7939
rect 7742 7936 7748 7948
rect 7703 7908 7748 7936
rect 7285 7899 7343 7905
rect 1670 7868 1676 7880
rect 1631 7840 1676 7868
rect 1670 7828 1676 7840
rect 1728 7828 1734 7880
rect 6730 7868 6736 7880
rect 6691 7840 6736 7868
rect 6730 7828 6736 7840
rect 6788 7828 6794 7880
rect 4341 7803 4399 7809
rect 4341 7769 4353 7803
rect 4387 7800 4399 7803
rect 4798 7800 4804 7812
rect 4387 7772 4804 7800
rect 4387 7769 4399 7772
rect 4341 7763 4399 7769
rect 4798 7760 4804 7772
rect 4856 7760 4862 7812
rect 5813 7803 5871 7809
rect 5813 7769 5825 7803
rect 5859 7800 5871 7803
rect 6454 7800 6460 7812
rect 5859 7772 6460 7800
rect 5859 7769 5871 7772
rect 5813 7763 5871 7769
rect 6454 7760 6460 7772
rect 6512 7800 6518 7812
rect 7300 7800 7328 7899
rect 7742 7896 7748 7908
rect 7800 7936 7806 7948
rect 7926 7936 7932 7948
rect 7800 7908 7932 7936
rect 7800 7896 7806 7908
rect 7926 7896 7932 7908
rect 7984 7896 7990 7948
rect 8297 7939 8355 7945
rect 8297 7905 8309 7939
rect 8343 7936 8355 7939
rect 8570 7936 8576 7948
rect 8343 7908 8576 7936
rect 8343 7905 8355 7908
rect 8297 7899 8355 7905
rect 8570 7896 8576 7908
rect 8628 7896 8634 7948
rect 8754 7936 8760 7948
rect 8715 7908 8760 7936
rect 8754 7896 8760 7908
rect 8812 7896 8818 7948
rect 10134 7896 10140 7948
rect 10192 7936 10198 7948
rect 10520 7945 10548 7976
rect 10505 7939 10563 7945
rect 10505 7936 10517 7939
rect 10192 7908 10517 7936
rect 10192 7896 10198 7908
rect 10505 7905 10517 7908
rect 10551 7905 10563 7939
rect 10686 7936 10692 7948
rect 10647 7908 10692 7936
rect 10505 7899 10563 7905
rect 10686 7896 10692 7908
rect 10744 7896 10750 7948
rect 10778 7896 10784 7948
rect 10836 7936 10842 7948
rect 10965 7939 11023 7945
rect 10965 7936 10977 7939
rect 10836 7908 10977 7936
rect 10836 7896 10842 7908
rect 10965 7905 10977 7908
rect 11011 7905 11023 7939
rect 10965 7899 11023 7905
rect 11517 7939 11575 7945
rect 11517 7905 11529 7939
rect 11563 7936 11575 7939
rect 12158 7936 12164 7948
rect 11563 7908 12164 7936
rect 11563 7905 11575 7908
rect 11517 7899 11575 7905
rect 12158 7896 12164 7908
rect 12216 7896 12222 7948
rect 12986 7936 12992 7948
rect 12947 7908 12992 7936
rect 12986 7896 12992 7908
rect 13044 7896 13050 7948
rect 13265 7939 13323 7945
rect 13265 7905 13277 7939
rect 13311 7936 13323 7939
rect 13630 7936 13636 7948
rect 13311 7908 13636 7936
rect 13311 7905 13323 7908
rect 13265 7899 13323 7905
rect 13630 7896 13636 7908
rect 13688 7896 13694 7948
rect 14185 7939 14243 7945
rect 14185 7905 14197 7939
rect 14231 7905 14243 7939
rect 14185 7899 14243 7905
rect 7374 7828 7380 7880
rect 7432 7868 7438 7880
rect 8386 7868 8392 7880
rect 7432 7840 8392 7868
rect 7432 7828 7438 7840
rect 8386 7828 8392 7840
rect 8444 7828 8450 7880
rect 11974 7828 11980 7880
rect 12032 7868 12038 7880
rect 12529 7871 12587 7877
rect 12529 7868 12541 7871
rect 12032 7840 12541 7868
rect 12032 7828 12038 7840
rect 12529 7837 12541 7840
rect 12575 7837 12587 7871
rect 13354 7868 13360 7880
rect 13315 7840 13360 7868
rect 12529 7831 12587 7837
rect 13354 7828 13360 7840
rect 13412 7828 13418 7880
rect 14200 7868 14228 7899
rect 14274 7896 14280 7948
rect 14332 7936 14338 7948
rect 14461 7939 14519 7945
rect 14461 7936 14473 7939
rect 14332 7908 14473 7936
rect 14332 7896 14338 7908
rect 14461 7905 14473 7908
rect 14507 7905 14519 7939
rect 14461 7899 14519 7905
rect 15654 7896 15660 7948
rect 15712 7936 15718 7948
rect 15841 7939 15899 7945
rect 15841 7936 15853 7939
rect 15712 7908 15853 7936
rect 15712 7896 15718 7908
rect 15841 7905 15853 7908
rect 15887 7936 15899 7939
rect 16022 7936 16028 7948
rect 15887 7908 16028 7936
rect 15887 7905 15899 7908
rect 15841 7899 15899 7905
rect 16022 7896 16028 7908
rect 16080 7896 16086 7948
rect 16301 7939 16359 7945
rect 16301 7905 16313 7939
rect 16347 7905 16359 7939
rect 16301 7899 16359 7905
rect 16485 7939 16543 7945
rect 16485 7905 16497 7939
rect 16531 7936 16543 7939
rect 16574 7936 16580 7948
rect 16531 7908 16580 7936
rect 16531 7905 16543 7908
rect 16485 7899 16543 7905
rect 14918 7868 14924 7880
rect 14200 7840 14924 7868
rect 8846 7800 8852 7812
rect 6512 7772 8852 7800
rect 6512 7760 6518 7772
rect 8846 7760 8852 7772
rect 8904 7800 8910 7812
rect 11146 7800 11152 7812
rect 8904 7772 11152 7800
rect 8904 7760 8910 7772
rect 11146 7760 11152 7772
rect 11204 7760 11210 7812
rect 11330 7760 11336 7812
rect 11388 7800 11394 7812
rect 14200 7800 14228 7840
rect 14918 7828 14924 7840
rect 14976 7828 14982 7880
rect 16316 7868 16344 7899
rect 16574 7896 16580 7908
rect 16632 7896 16638 7948
rect 16758 7896 16764 7948
rect 16816 7936 16822 7948
rect 16853 7939 16911 7945
rect 16853 7936 16865 7939
rect 16816 7908 16865 7936
rect 16816 7896 16822 7908
rect 16853 7905 16865 7908
rect 16899 7936 16911 7939
rect 17494 7936 17500 7948
rect 16899 7908 17500 7936
rect 16899 7905 16911 7908
rect 16853 7899 16911 7905
rect 17494 7896 17500 7908
rect 17552 7896 17558 7948
rect 17589 7939 17647 7945
rect 17589 7905 17601 7939
rect 17635 7936 17647 7939
rect 17678 7936 17684 7948
rect 17635 7908 17684 7936
rect 17635 7905 17647 7908
rect 17589 7899 17647 7905
rect 17678 7896 17684 7908
rect 17736 7936 17742 7948
rect 18064 7936 18092 7976
rect 18230 7964 18236 7976
rect 18288 7964 18294 8016
rect 18340 8004 18368 8044
rect 20073 8041 20085 8075
rect 20119 8072 20131 8075
rect 20162 8072 20168 8084
rect 20119 8044 20168 8072
rect 20119 8041 20131 8044
rect 20073 8035 20131 8041
rect 20162 8032 20168 8044
rect 20220 8032 20226 8084
rect 20898 8032 20904 8084
rect 20956 8072 20962 8084
rect 20993 8075 21051 8081
rect 20993 8072 21005 8075
rect 20956 8044 21005 8072
rect 20956 8032 20962 8044
rect 20993 8041 21005 8044
rect 21039 8041 21051 8075
rect 20993 8035 21051 8041
rect 22094 8032 22100 8084
rect 22152 8072 22158 8084
rect 23198 8072 23204 8084
rect 22152 8044 23204 8072
rect 22152 8032 22158 8044
rect 23198 8032 23204 8044
rect 23256 8032 23262 8084
rect 23474 8072 23480 8084
rect 23435 8044 23480 8072
rect 23474 8032 23480 8044
rect 23532 8032 23538 8084
rect 27062 8032 27068 8084
rect 27120 8072 27126 8084
rect 30098 8072 30104 8084
rect 27120 8044 30104 8072
rect 27120 8032 27126 8044
rect 30098 8032 30104 8044
rect 30156 8032 30162 8084
rect 30926 8032 30932 8084
rect 30984 8072 30990 8084
rect 31021 8075 31079 8081
rect 31021 8072 31033 8075
rect 30984 8044 31033 8072
rect 30984 8032 30990 8044
rect 31021 8041 31033 8044
rect 31067 8041 31079 8075
rect 31021 8035 31079 8041
rect 31113 8075 31171 8081
rect 31113 8041 31125 8075
rect 31159 8072 31171 8075
rect 32122 8072 32128 8084
rect 31159 8044 31340 8072
rect 31159 8041 31171 8044
rect 31113 8035 31171 8041
rect 20806 8004 20812 8016
rect 18340 7976 20812 8004
rect 20806 7964 20812 7976
rect 20864 7964 20870 8016
rect 23750 8004 23756 8016
rect 21008 7976 23756 8004
rect 18414 7936 18420 7948
rect 17736 7908 18000 7936
rect 18064 7908 18420 7936
rect 17736 7896 17742 7908
rect 16942 7868 16948 7880
rect 16316 7840 16948 7868
rect 16942 7828 16948 7840
rect 17000 7828 17006 7880
rect 11388 7772 14228 7800
rect 11388 7760 11394 7772
rect 15562 7760 15568 7812
rect 15620 7800 15626 7812
rect 15749 7803 15807 7809
rect 15749 7800 15761 7803
rect 15620 7772 15761 7800
rect 15620 7760 15626 7772
rect 15749 7769 15761 7772
rect 15795 7769 15807 7803
rect 15749 7763 15807 7769
rect 8386 7692 8392 7744
rect 8444 7732 8450 7744
rect 8754 7732 8760 7744
rect 8444 7704 8760 7732
rect 8444 7692 8450 7704
rect 8754 7692 8760 7704
rect 8812 7692 8818 7744
rect 9493 7735 9551 7741
rect 9493 7701 9505 7735
rect 9539 7732 9551 7735
rect 11422 7732 11428 7744
rect 9539 7704 11428 7732
rect 9539 7701 9551 7704
rect 9493 7695 9551 7701
rect 11422 7692 11428 7704
rect 11480 7692 11486 7744
rect 12250 7692 12256 7744
rect 12308 7732 12314 7744
rect 16850 7732 16856 7744
rect 12308 7704 16856 7732
rect 12308 7692 12314 7704
rect 16850 7692 16856 7704
rect 16908 7692 16914 7744
rect 17972 7732 18000 7908
rect 18414 7896 18420 7908
rect 18472 7896 18478 7948
rect 18874 7936 18880 7948
rect 18835 7908 18880 7936
rect 18874 7896 18880 7908
rect 18932 7896 18938 7948
rect 18969 7939 19027 7945
rect 18969 7905 18981 7939
rect 19015 7936 19027 7939
rect 19058 7936 19064 7948
rect 19015 7908 19064 7936
rect 19015 7905 19027 7908
rect 18969 7899 19027 7905
rect 19058 7896 19064 7908
rect 19116 7896 19122 7948
rect 19245 7939 19303 7945
rect 19245 7905 19257 7939
rect 19291 7936 19303 7939
rect 19426 7936 19432 7948
rect 19291 7908 19432 7936
rect 19291 7905 19303 7908
rect 19245 7899 19303 7905
rect 19426 7896 19432 7908
rect 19484 7896 19490 7948
rect 19886 7936 19892 7948
rect 19847 7908 19892 7936
rect 19886 7896 19892 7908
rect 19944 7896 19950 7948
rect 20162 7896 20168 7948
rect 20220 7936 20226 7948
rect 20901 7939 20959 7945
rect 20901 7936 20913 7939
rect 20220 7908 20913 7936
rect 20220 7896 20226 7908
rect 20901 7905 20913 7908
rect 20947 7905 20959 7939
rect 20901 7899 20959 7905
rect 19337 7871 19395 7877
rect 19337 7837 19349 7871
rect 19383 7868 19395 7871
rect 20180 7868 20208 7896
rect 19383 7840 20208 7868
rect 19383 7837 19395 7840
rect 19337 7831 19395 7837
rect 18414 7760 18420 7812
rect 18472 7800 18478 7812
rect 19886 7800 19892 7812
rect 18472 7772 19892 7800
rect 18472 7760 18478 7772
rect 19886 7760 19892 7772
rect 19944 7760 19950 7812
rect 21008 7732 21036 7976
rect 23750 7964 23756 7976
rect 23808 7964 23814 8016
rect 24302 7964 24308 8016
rect 24360 8004 24366 8016
rect 26970 8004 26976 8016
rect 24360 7976 24532 8004
rect 24360 7964 24366 7976
rect 21453 7939 21511 7945
rect 21453 7905 21465 7939
rect 21499 7905 21511 7939
rect 21453 7899 21511 7905
rect 21468 7800 21496 7899
rect 21818 7896 21824 7948
rect 21876 7936 21882 7948
rect 22465 7939 22523 7945
rect 22465 7936 22477 7939
rect 21876 7908 22477 7936
rect 21876 7896 21882 7908
rect 22465 7905 22477 7908
rect 22511 7905 22523 7939
rect 22465 7899 22523 7905
rect 22922 7896 22928 7948
rect 22980 7936 22986 7948
rect 23017 7939 23075 7945
rect 23017 7936 23029 7939
rect 22980 7908 23029 7936
rect 22980 7896 22986 7908
rect 23017 7905 23029 7908
rect 23063 7905 23075 7939
rect 23198 7936 23204 7948
rect 23159 7908 23204 7936
rect 23017 7899 23075 7905
rect 23198 7896 23204 7908
rect 23256 7936 23262 7948
rect 24394 7936 24400 7948
rect 23256 7908 24256 7936
rect 24355 7908 24400 7936
rect 23256 7896 23262 7908
rect 22002 7828 22008 7880
rect 22060 7868 22066 7880
rect 22281 7871 22339 7877
rect 22281 7868 22293 7871
rect 22060 7840 22293 7868
rect 22060 7828 22066 7840
rect 22281 7837 22293 7840
rect 22327 7837 22339 7871
rect 24228 7868 24256 7908
rect 24394 7896 24400 7908
rect 24452 7896 24458 7948
rect 24504 7945 24532 7976
rect 25792 7976 26976 8004
rect 24489 7939 24547 7945
rect 24489 7905 24501 7939
rect 24535 7905 24547 7939
rect 25130 7936 25136 7948
rect 25091 7908 25136 7936
rect 24489 7899 24547 7905
rect 25130 7896 25136 7908
rect 25188 7896 25194 7948
rect 25792 7945 25820 7976
rect 26970 7964 26976 7976
rect 27028 7964 27034 8016
rect 27816 7976 28856 8004
rect 25777 7939 25835 7945
rect 25777 7905 25789 7939
rect 25823 7905 25835 7939
rect 25777 7899 25835 7905
rect 26789 7939 26847 7945
rect 26789 7905 26801 7939
rect 26835 7936 26847 7939
rect 27246 7936 27252 7948
rect 26835 7908 27252 7936
rect 26835 7905 26847 7908
rect 26789 7899 26847 7905
rect 26804 7868 26832 7899
rect 27246 7896 27252 7908
rect 27304 7896 27310 7948
rect 27430 7936 27436 7948
rect 27391 7908 27436 7936
rect 27430 7896 27436 7908
rect 27488 7896 27494 7948
rect 27816 7945 27844 7976
rect 27801 7939 27859 7945
rect 27801 7905 27813 7939
rect 27847 7905 27859 7939
rect 27982 7936 27988 7948
rect 27943 7908 27988 7936
rect 27801 7899 27859 7905
rect 27982 7896 27988 7908
rect 28040 7896 28046 7948
rect 27154 7868 27160 7880
rect 24228 7840 26832 7868
rect 27115 7840 27160 7868
rect 22281 7831 22339 7837
rect 27154 7828 27160 7840
rect 27212 7828 27218 7880
rect 28721 7871 28779 7877
rect 28721 7837 28733 7871
rect 28767 7837 28779 7871
rect 28828 7868 28856 7976
rect 30650 7964 30656 8016
rect 30708 8004 30714 8016
rect 30837 8007 30895 8013
rect 30837 8004 30849 8007
rect 30708 7976 30849 8004
rect 30708 7964 30714 7976
rect 30837 7973 30849 7976
rect 30883 7973 30895 8007
rect 30837 7967 30895 7973
rect 31205 8007 31263 8013
rect 31205 7973 31217 8007
rect 31251 7973 31263 8007
rect 31205 7967 31263 7973
rect 28997 7939 29055 7945
rect 28997 7905 29009 7939
rect 29043 7936 29055 7939
rect 29362 7936 29368 7948
rect 29043 7908 29368 7936
rect 29043 7905 29055 7908
rect 28997 7899 29055 7905
rect 29362 7896 29368 7908
rect 29420 7896 29426 7948
rect 30282 7896 30288 7948
rect 30340 7936 30346 7948
rect 31220 7936 31248 7967
rect 30340 7908 30696 7936
rect 30340 7896 30346 7908
rect 30466 7868 30472 7880
rect 28828 7840 30472 7868
rect 28721 7831 28779 7837
rect 27246 7800 27252 7812
rect 21468 7772 27252 7800
rect 27246 7760 27252 7772
rect 27304 7760 27310 7812
rect 17972 7704 21036 7732
rect 21082 7692 21088 7744
rect 21140 7732 21146 7744
rect 24213 7735 24271 7741
rect 24213 7732 24225 7735
rect 21140 7704 24225 7732
rect 21140 7692 21146 7704
rect 24213 7701 24225 7704
rect 24259 7701 24271 7735
rect 24213 7695 24271 7701
rect 25869 7735 25927 7741
rect 25869 7701 25881 7735
rect 25915 7732 25927 7735
rect 27338 7732 27344 7744
rect 25915 7704 27344 7732
rect 25915 7701 25927 7704
rect 25869 7695 25927 7701
rect 27338 7692 27344 7704
rect 27396 7692 27402 7744
rect 28736 7732 28764 7831
rect 30466 7828 30472 7840
rect 30524 7828 30530 7880
rect 30668 7868 30696 7908
rect 30944 7908 31248 7936
rect 30944 7868 30972 7908
rect 30668 7840 30972 7868
rect 30098 7760 30104 7812
rect 30156 7800 30162 7812
rect 31312 7800 31340 8044
rect 31588 8044 32128 8072
rect 31588 8013 31616 8044
rect 32122 8032 32128 8044
rect 32180 8032 32186 8084
rect 32306 8072 32312 8084
rect 32267 8044 32312 8072
rect 32306 8032 32312 8044
rect 32364 8032 32370 8084
rect 32490 8032 32496 8084
rect 32548 8072 32554 8084
rect 34885 8075 34943 8081
rect 34885 8072 34897 8075
rect 32548 8044 34897 8072
rect 32548 8032 32554 8044
rect 34885 8041 34897 8044
rect 34931 8041 34943 8075
rect 34885 8035 34943 8041
rect 31573 8007 31631 8013
rect 31573 7973 31585 8007
rect 31619 7973 31631 8007
rect 34054 8004 34060 8016
rect 31573 7967 31631 7973
rect 33428 7976 34060 8004
rect 32125 7939 32183 7945
rect 32125 7905 32137 7939
rect 32171 7936 32183 7939
rect 32398 7936 32404 7948
rect 32171 7908 32404 7936
rect 32171 7905 32183 7908
rect 32125 7899 32183 7905
rect 32398 7896 32404 7908
rect 32456 7896 32462 7948
rect 33318 7896 33324 7948
rect 33376 7936 33382 7948
rect 33428 7945 33456 7976
rect 34054 7964 34060 7976
rect 34112 8004 34118 8016
rect 34112 7976 34836 8004
rect 34112 7964 34118 7976
rect 33413 7939 33471 7945
rect 33413 7936 33425 7939
rect 33376 7908 33425 7936
rect 33376 7896 33382 7908
rect 33413 7905 33425 7908
rect 33459 7905 33471 7939
rect 33870 7936 33876 7948
rect 33831 7908 33876 7936
rect 33413 7899 33471 7905
rect 33870 7896 33876 7908
rect 33928 7896 33934 7948
rect 34238 7936 34244 7948
rect 34199 7908 34244 7936
rect 34238 7896 34244 7908
rect 34296 7896 34302 7948
rect 34808 7945 34836 7976
rect 34793 7939 34851 7945
rect 34793 7905 34805 7939
rect 34839 7905 34851 7939
rect 34793 7899 34851 7905
rect 35250 7896 35256 7948
rect 35308 7936 35314 7948
rect 35345 7939 35403 7945
rect 35345 7936 35357 7939
rect 35308 7908 35357 7936
rect 35308 7896 35314 7908
rect 35345 7905 35357 7908
rect 35391 7905 35403 7939
rect 35345 7899 35403 7905
rect 35434 7896 35440 7948
rect 35492 7936 35498 7948
rect 36357 7939 36415 7945
rect 36357 7936 36369 7939
rect 35492 7908 36369 7936
rect 35492 7896 35498 7908
rect 36357 7905 36369 7908
rect 36403 7905 36415 7939
rect 36357 7899 36415 7905
rect 34514 7828 34520 7880
rect 34572 7868 34578 7880
rect 35621 7871 35679 7877
rect 35621 7868 35633 7871
rect 34572 7840 35633 7868
rect 34572 7828 34578 7840
rect 35621 7837 35633 7840
rect 35667 7837 35679 7871
rect 35621 7831 35679 7837
rect 30156 7772 31340 7800
rect 30156 7760 30162 7772
rect 32214 7760 32220 7812
rect 32272 7800 32278 7812
rect 33321 7803 33379 7809
rect 33321 7800 33333 7803
rect 32272 7772 33333 7800
rect 32272 7760 32278 7772
rect 33321 7769 33333 7772
rect 33367 7769 33379 7803
rect 33321 7763 33379 7769
rect 29178 7732 29184 7744
rect 28736 7704 29184 7732
rect 29178 7692 29184 7704
rect 29236 7732 29242 7744
rect 29454 7732 29460 7744
rect 29236 7704 29460 7732
rect 29236 7692 29242 7704
rect 29454 7692 29460 7704
rect 29512 7692 29518 7744
rect 30466 7692 30472 7744
rect 30524 7732 30530 7744
rect 31478 7732 31484 7744
rect 30524 7704 31484 7732
rect 30524 7692 30530 7704
rect 31478 7692 31484 7704
rect 31536 7732 31542 7744
rect 36449 7735 36507 7741
rect 36449 7732 36461 7735
rect 31536 7704 36461 7732
rect 31536 7692 31542 7704
rect 36449 7701 36461 7704
rect 36495 7701 36507 7735
rect 36449 7695 36507 7701
rect 1104 7642 38824 7664
rect 1104 7590 4246 7642
rect 4298 7590 4310 7642
rect 4362 7590 4374 7642
rect 4426 7590 4438 7642
rect 4490 7590 34966 7642
rect 35018 7590 35030 7642
rect 35082 7590 35094 7642
rect 35146 7590 35158 7642
rect 35210 7590 38824 7642
rect 1104 7568 38824 7590
rect 4157 7531 4215 7537
rect 4157 7497 4169 7531
rect 4203 7528 4215 7531
rect 4614 7528 4620 7540
rect 4203 7500 4620 7528
rect 4203 7497 4215 7500
rect 4157 7491 4215 7497
rect 4614 7488 4620 7500
rect 4672 7488 4678 7540
rect 7285 7531 7343 7537
rect 7285 7497 7297 7531
rect 7331 7528 7343 7531
rect 9214 7528 9220 7540
rect 7331 7500 9220 7528
rect 7331 7497 7343 7500
rect 7285 7491 7343 7497
rect 5077 7395 5135 7401
rect 5077 7361 5089 7395
rect 5123 7392 5135 7395
rect 5350 7392 5356 7404
rect 5123 7364 5356 7392
rect 5123 7361 5135 7364
rect 5077 7355 5135 7361
rect 5350 7352 5356 7364
rect 5408 7352 5414 7404
rect 7300 7392 7328 7491
rect 9214 7488 9220 7500
rect 9272 7488 9278 7540
rect 14182 7528 14188 7540
rect 11256 7500 14188 7528
rect 7742 7420 7748 7472
rect 7800 7460 7806 7472
rect 10410 7460 10416 7472
rect 7800 7432 9076 7460
rect 10371 7432 10416 7460
rect 7800 7420 7806 7432
rect 7926 7392 7932 7404
rect 5644 7364 7328 7392
rect 7887 7364 7932 7392
rect 2590 7324 2596 7336
rect 2551 7296 2596 7324
rect 2590 7284 2596 7296
rect 2648 7284 2654 7336
rect 2869 7327 2927 7333
rect 2869 7293 2881 7327
rect 2915 7324 2927 7327
rect 4154 7324 4160 7336
rect 2915 7296 4160 7324
rect 2915 7293 2927 7296
rect 2869 7287 2927 7293
rect 4154 7284 4160 7296
rect 4212 7284 4218 7336
rect 4798 7324 4804 7336
rect 4759 7296 4804 7324
rect 4798 7284 4804 7296
rect 4856 7284 4862 7336
rect 4982 7284 4988 7336
rect 5040 7324 5046 7336
rect 5445 7327 5503 7333
rect 5445 7324 5457 7327
rect 5040 7296 5457 7324
rect 5040 7284 5046 7296
rect 5445 7293 5457 7296
rect 5491 7324 5503 7327
rect 5644 7324 5672 7364
rect 7926 7352 7932 7364
rect 7984 7352 7990 7404
rect 5491 7296 5672 7324
rect 5997 7327 6055 7333
rect 5491 7293 5503 7296
rect 5445 7287 5503 7293
rect 5997 7293 6009 7327
rect 6043 7324 6055 7327
rect 6086 7324 6092 7336
rect 6043 7296 6092 7324
rect 6043 7293 6055 7296
rect 5997 7287 6055 7293
rect 6086 7284 6092 7296
rect 6144 7284 6150 7336
rect 7101 7327 7159 7333
rect 7101 7293 7113 7327
rect 7147 7324 7159 7327
rect 7374 7324 7380 7336
rect 7147 7296 7380 7324
rect 7147 7293 7159 7296
rect 7101 7287 7159 7293
rect 7374 7284 7380 7296
rect 7432 7284 7438 7336
rect 7834 7324 7840 7336
rect 7795 7296 7840 7324
rect 7834 7284 7840 7296
rect 7892 7284 7898 7336
rect 8481 7327 8539 7333
rect 8481 7293 8493 7327
rect 8527 7293 8539 7327
rect 8846 7324 8852 7336
rect 8807 7296 8852 7324
rect 8481 7287 8539 7293
rect 8496 7256 8524 7287
rect 8846 7284 8852 7296
rect 8904 7284 8910 7336
rect 9048 7333 9076 7432
rect 10410 7420 10416 7432
rect 10468 7420 10474 7472
rect 9398 7352 9404 7404
rect 9456 7392 9462 7404
rect 10873 7395 10931 7401
rect 10873 7392 10885 7395
rect 9456 7364 10885 7392
rect 9456 7352 9462 7364
rect 10873 7361 10885 7364
rect 10919 7392 10931 7395
rect 11054 7392 11060 7404
rect 10919 7364 11060 7392
rect 10919 7361 10931 7364
rect 10873 7355 10931 7361
rect 11054 7352 11060 7364
rect 11112 7352 11118 7404
rect 9033 7327 9091 7333
rect 9033 7293 9045 7327
rect 9079 7293 9091 7327
rect 9033 7287 9091 7293
rect 9585 7327 9643 7333
rect 9585 7293 9597 7327
rect 9631 7324 9643 7327
rect 10502 7324 10508 7336
rect 9631 7296 10508 7324
rect 9631 7293 9643 7296
rect 9585 7287 9643 7293
rect 10502 7284 10508 7296
rect 10560 7284 10566 7336
rect 10597 7327 10655 7333
rect 10597 7293 10609 7327
rect 10643 7324 10655 7327
rect 11256 7324 11284 7500
rect 14182 7488 14188 7500
rect 14240 7488 14246 7540
rect 15930 7528 15936 7540
rect 15304 7500 15936 7528
rect 13630 7460 13636 7472
rect 13591 7432 13636 7460
rect 13630 7420 13636 7432
rect 13688 7420 13694 7472
rect 11790 7392 11796 7404
rect 11751 7364 11796 7392
rect 11790 7352 11796 7364
rect 11848 7352 11854 7404
rect 14550 7392 14556 7404
rect 14511 7364 14556 7392
rect 14550 7352 14556 7364
rect 14608 7352 14614 7404
rect 15304 7401 15332 7500
rect 15930 7488 15936 7500
rect 15988 7488 15994 7540
rect 16853 7531 16911 7537
rect 16853 7497 16865 7531
rect 16899 7528 16911 7531
rect 17310 7528 17316 7540
rect 16899 7500 17316 7528
rect 16899 7497 16911 7500
rect 16853 7491 16911 7497
rect 17310 7488 17316 7500
rect 17368 7488 17374 7540
rect 20622 7528 20628 7540
rect 18340 7500 20628 7528
rect 15289 7395 15347 7401
rect 15289 7361 15301 7395
rect 15335 7361 15347 7395
rect 15562 7392 15568 7404
rect 15523 7364 15568 7392
rect 15289 7355 15347 7361
rect 15562 7352 15568 7364
rect 15620 7352 15626 7404
rect 15746 7352 15752 7404
rect 15804 7392 15810 7404
rect 16482 7392 16488 7404
rect 15804 7364 16488 7392
rect 15804 7352 15810 7364
rect 16482 7352 16488 7364
rect 16540 7352 16546 7404
rect 10643 7296 11284 7324
rect 11333 7327 11391 7333
rect 10643 7293 10655 7296
rect 10597 7287 10655 7293
rect 11333 7293 11345 7327
rect 11379 7324 11391 7327
rect 11422 7324 11428 7336
rect 11379 7296 11428 7324
rect 11379 7293 11391 7296
rect 11333 7287 11391 7293
rect 11422 7284 11428 7296
rect 11480 7284 11486 7336
rect 11698 7324 11704 7336
rect 11659 7296 11704 7324
rect 11698 7284 11704 7296
rect 11756 7284 11762 7336
rect 12897 7327 12955 7333
rect 12897 7293 12909 7327
rect 12943 7293 12955 7327
rect 12897 7287 12955 7293
rect 13725 7327 13783 7333
rect 13725 7293 13737 7327
rect 13771 7324 13783 7327
rect 13906 7324 13912 7336
rect 13771 7296 13912 7324
rect 13771 7293 13783 7296
rect 13725 7287 13783 7293
rect 8496 7228 8616 7256
rect 6178 7188 6184 7200
rect 6139 7160 6184 7188
rect 6178 7148 6184 7160
rect 6236 7148 6242 7200
rect 8588 7188 8616 7228
rect 10410 7216 10416 7268
rect 10468 7256 10474 7268
rect 12710 7256 12716 7268
rect 10468 7228 12716 7256
rect 10468 7216 10474 7228
rect 12710 7216 12716 7228
rect 12768 7216 12774 7268
rect 12912 7256 12940 7287
rect 13906 7284 13912 7296
rect 13964 7284 13970 7336
rect 14090 7324 14096 7336
rect 14051 7296 14096 7324
rect 14090 7284 14096 7296
rect 14148 7284 14154 7336
rect 18340 7324 18368 7500
rect 20622 7488 20628 7500
rect 20680 7488 20686 7540
rect 22830 7488 22836 7540
rect 22888 7528 22894 7540
rect 25869 7531 25927 7537
rect 22888 7500 25176 7528
rect 22888 7488 22894 7500
rect 25148 7472 25176 7500
rect 25869 7497 25881 7531
rect 25915 7528 25927 7531
rect 27430 7528 27436 7540
rect 25915 7500 27436 7528
rect 25915 7497 25927 7500
rect 25869 7491 25927 7497
rect 27430 7488 27436 7500
rect 27488 7488 27494 7540
rect 30282 7488 30288 7540
rect 30340 7528 30346 7540
rect 32493 7531 32551 7537
rect 32493 7528 32505 7531
rect 30340 7500 32505 7528
rect 30340 7488 30346 7500
rect 32493 7497 32505 7500
rect 32539 7528 32551 7531
rect 35434 7528 35440 7540
rect 32539 7500 35440 7528
rect 32539 7497 32551 7500
rect 32493 7491 32551 7497
rect 35434 7488 35440 7500
rect 35492 7488 35498 7540
rect 37826 7528 37832 7540
rect 37787 7500 37832 7528
rect 37826 7488 37832 7500
rect 37884 7488 37890 7540
rect 21726 7460 21732 7472
rect 18984 7432 21732 7460
rect 15396 7296 18368 7324
rect 15396 7256 15424 7296
rect 18414 7284 18420 7336
rect 18472 7324 18478 7336
rect 18984 7333 19012 7432
rect 21726 7420 21732 7432
rect 21784 7420 21790 7472
rect 24302 7460 24308 7472
rect 22388 7432 24308 7460
rect 19150 7392 19156 7404
rect 19111 7364 19156 7392
rect 19150 7352 19156 7364
rect 19208 7352 19214 7404
rect 19886 7392 19892 7404
rect 19847 7364 19892 7392
rect 19886 7352 19892 7364
rect 19944 7352 19950 7404
rect 22186 7392 22192 7404
rect 22147 7364 22192 7392
rect 22186 7352 22192 7364
rect 22244 7352 22250 7404
rect 18969 7327 19027 7333
rect 18472 7296 18517 7324
rect 18472 7284 18478 7296
rect 18969 7293 18981 7327
rect 19015 7293 19027 7327
rect 18969 7287 19027 7293
rect 19334 7284 19340 7336
rect 19392 7324 19398 7336
rect 19613 7327 19671 7333
rect 19613 7324 19625 7327
rect 19392 7296 19625 7324
rect 19392 7284 19398 7296
rect 19613 7293 19625 7296
rect 19659 7293 19671 7327
rect 19613 7287 19671 7293
rect 20257 7327 20315 7333
rect 20257 7293 20269 7327
rect 20303 7293 20315 7327
rect 20530 7324 20536 7336
rect 20491 7296 20536 7324
rect 20257 7287 20315 7293
rect 12912 7228 15424 7256
rect 19628 7256 19656 7287
rect 20162 7256 20168 7268
rect 19628 7228 20168 7256
rect 20162 7216 20168 7228
rect 20220 7216 20226 7268
rect 20272 7256 20300 7287
rect 20530 7284 20536 7296
rect 20588 7284 20594 7336
rect 21910 7324 21916 7336
rect 21871 7296 21916 7324
rect 21910 7284 21916 7296
rect 21968 7284 21974 7336
rect 22094 7284 22100 7336
rect 22152 7324 22158 7336
rect 22388 7333 22416 7432
rect 24302 7420 24308 7432
rect 24360 7420 24366 7472
rect 25130 7420 25136 7472
rect 25188 7460 25194 7472
rect 29270 7460 29276 7472
rect 25188 7432 29276 7460
rect 25188 7420 25194 7432
rect 29270 7420 29276 7432
rect 29328 7420 29334 7472
rect 29454 7420 29460 7472
rect 29512 7460 29518 7472
rect 33410 7460 33416 7472
rect 29512 7432 30972 7460
rect 33371 7432 33416 7460
rect 29512 7420 29518 7432
rect 26878 7392 26884 7404
rect 26839 7364 26884 7392
rect 26878 7352 26884 7364
rect 26936 7352 26942 7404
rect 27338 7352 27344 7404
rect 27396 7392 27402 7404
rect 30944 7401 30972 7432
rect 33410 7420 33416 7432
rect 33468 7420 33474 7472
rect 36170 7420 36176 7472
rect 36228 7460 36234 7472
rect 36228 7432 36492 7460
rect 36228 7420 36234 7432
rect 30929 7395 30987 7401
rect 27396 7364 29960 7392
rect 27396 7352 27402 7364
rect 22373 7327 22431 7333
rect 22373 7324 22385 7327
rect 22152 7296 22385 7324
rect 22152 7284 22158 7296
rect 22373 7293 22385 7296
rect 22419 7293 22431 7327
rect 22373 7287 22431 7293
rect 22741 7327 22799 7333
rect 22741 7293 22753 7327
rect 22787 7324 22799 7327
rect 22830 7324 22836 7336
rect 22787 7296 22836 7324
rect 22787 7293 22799 7296
rect 22741 7287 22799 7293
rect 22830 7284 22836 7296
rect 22888 7284 22894 7336
rect 23842 7324 23848 7336
rect 23803 7296 23848 7324
rect 23842 7284 23848 7296
rect 23900 7284 23906 7336
rect 23937 7327 23995 7333
rect 23937 7293 23949 7327
rect 23983 7324 23995 7327
rect 23983 7296 24348 7324
rect 23983 7293 23995 7296
rect 23937 7287 23995 7293
rect 20806 7256 20812 7268
rect 20272 7228 20812 7256
rect 20806 7216 20812 7228
rect 20864 7256 20870 7268
rect 21266 7256 21272 7268
rect 20864 7228 21272 7256
rect 20864 7216 20870 7228
rect 21266 7216 21272 7228
rect 21324 7216 21330 7268
rect 22278 7256 22284 7268
rect 21376 7228 22284 7256
rect 11974 7188 11980 7200
rect 8588 7160 11980 7188
rect 11974 7148 11980 7160
rect 12032 7148 12038 7200
rect 12158 7148 12164 7200
rect 12216 7188 12222 7200
rect 12989 7191 13047 7197
rect 12989 7188 13001 7191
rect 12216 7160 13001 7188
rect 12216 7148 12222 7160
rect 12989 7157 13001 7160
rect 13035 7188 13047 7191
rect 15562 7188 15568 7200
rect 13035 7160 15568 7188
rect 13035 7157 13047 7160
rect 12989 7151 13047 7157
rect 15562 7148 15568 7160
rect 15620 7148 15626 7200
rect 16482 7148 16488 7200
rect 16540 7188 16546 7200
rect 21376 7188 21404 7228
rect 22278 7216 22284 7228
rect 22336 7216 22342 7268
rect 24320 7256 24348 7296
rect 24394 7284 24400 7336
rect 24452 7324 24458 7336
rect 24578 7324 24584 7336
rect 24452 7296 24497 7324
rect 24539 7296 24584 7324
rect 24452 7284 24458 7296
rect 24578 7284 24584 7296
rect 24636 7324 24642 7336
rect 25590 7324 25596 7336
rect 24636 7296 25596 7324
rect 24636 7284 24642 7296
rect 25590 7284 25596 7296
rect 25648 7284 25654 7336
rect 25685 7327 25743 7333
rect 25685 7293 25697 7327
rect 25731 7324 25743 7327
rect 26326 7324 26332 7336
rect 25731 7296 26332 7324
rect 25731 7293 25743 7296
rect 25685 7287 25743 7293
rect 26326 7284 26332 7296
rect 26384 7284 26390 7336
rect 26697 7327 26755 7333
rect 26697 7293 26709 7327
rect 26743 7293 26755 7327
rect 26970 7324 26976 7336
rect 26931 7296 26976 7324
rect 26697 7287 26755 7293
rect 26712 7256 26740 7287
rect 26970 7284 26976 7296
rect 27028 7284 27034 7336
rect 27246 7324 27252 7336
rect 27207 7296 27252 7324
rect 27246 7284 27252 7296
rect 27304 7284 27310 7336
rect 27890 7324 27896 7336
rect 27851 7296 27896 7324
rect 27890 7284 27896 7296
rect 27948 7284 27954 7336
rect 28258 7284 28264 7336
rect 28316 7324 28322 7336
rect 28353 7327 28411 7333
rect 28353 7324 28365 7327
rect 28316 7296 28365 7324
rect 28316 7284 28322 7296
rect 28353 7293 28365 7296
rect 28399 7293 28411 7327
rect 28353 7287 28411 7293
rect 29546 7284 29552 7336
rect 29604 7324 29610 7336
rect 29932 7333 29960 7364
rect 30929 7361 30941 7395
rect 30975 7361 30987 7395
rect 30929 7355 30987 7361
rect 31110 7352 31116 7404
rect 31168 7392 31174 7404
rect 31205 7395 31263 7401
rect 31205 7392 31217 7395
rect 31168 7364 31217 7392
rect 31168 7352 31174 7364
rect 31205 7361 31217 7364
rect 31251 7361 31263 7395
rect 33318 7392 33324 7404
rect 31205 7355 31263 7361
rect 33152 7364 33324 7392
rect 29733 7327 29791 7333
rect 29733 7324 29745 7327
rect 29604 7296 29745 7324
rect 29604 7284 29610 7296
rect 29733 7293 29745 7296
rect 29779 7293 29791 7327
rect 29733 7287 29791 7293
rect 29917 7327 29975 7333
rect 29917 7293 29929 7327
rect 29963 7293 29975 7327
rect 29917 7287 29975 7293
rect 30101 7327 30159 7333
rect 30101 7293 30113 7327
rect 30147 7324 30159 7327
rect 30834 7324 30840 7336
rect 30147 7296 30840 7324
rect 30147 7293 30159 7296
rect 30101 7287 30159 7293
rect 30834 7284 30840 7296
rect 30892 7284 30898 7336
rect 33152 7333 33180 7364
rect 33318 7352 33324 7364
rect 33376 7352 33382 7404
rect 34149 7395 34207 7401
rect 34149 7361 34161 7395
rect 34195 7392 34207 7395
rect 34238 7392 34244 7404
rect 34195 7364 34244 7392
rect 34195 7361 34207 7364
rect 34149 7355 34207 7361
rect 34238 7352 34244 7364
rect 34296 7352 34302 7404
rect 35342 7352 35348 7404
rect 35400 7392 35406 7404
rect 35529 7395 35587 7401
rect 35529 7392 35541 7395
rect 35400 7364 35541 7392
rect 35400 7352 35406 7364
rect 35529 7361 35541 7364
rect 35575 7361 35587 7395
rect 35529 7355 35587 7361
rect 35989 7395 36047 7401
rect 35989 7361 36001 7395
rect 36035 7392 36047 7395
rect 36354 7392 36360 7404
rect 36035 7364 36360 7392
rect 36035 7361 36047 7364
rect 35989 7355 36047 7361
rect 36354 7352 36360 7364
rect 36412 7352 36418 7404
rect 36464 7392 36492 7432
rect 36725 7395 36783 7401
rect 36725 7392 36737 7395
rect 36464 7364 36737 7392
rect 36725 7361 36737 7364
rect 36771 7361 36783 7395
rect 36725 7355 36783 7361
rect 33137 7327 33195 7333
rect 33137 7293 33149 7327
rect 33183 7293 33195 7327
rect 33137 7287 33195 7293
rect 33226 7284 33232 7336
rect 33284 7324 33290 7336
rect 33689 7327 33747 7333
rect 33689 7324 33701 7327
rect 33284 7296 33701 7324
rect 33284 7284 33290 7296
rect 33689 7293 33701 7296
rect 33735 7293 33747 7327
rect 33689 7287 33747 7293
rect 34977 7327 35035 7333
rect 34977 7293 34989 7327
rect 35023 7324 35035 7327
rect 35710 7324 35716 7336
rect 35023 7296 35716 7324
rect 35023 7293 35035 7296
rect 34977 7287 35035 7293
rect 35710 7284 35716 7296
rect 35768 7284 35774 7336
rect 35805 7327 35863 7333
rect 35805 7293 35817 7327
rect 35851 7324 35863 7327
rect 36078 7324 36084 7336
rect 35851 7296 36084 7324
rect 35851 7293 35863 7296
rect 35805 7287 35863 7293
rect 36078 7284 36084 7296
rect 36136 7284 36142 7336
rect 36170 7284 36176 7336
rect 36228 7324 36234 7336
rect 36449 7327 36507 7333
rect 36449 7324 36461 7327
rect 36228 7296 36461 7324
rect 36228 7284 36234 7296
rect 36449 7293 36461 7296
rect 36495 7293 36507 7327
rect 36449 7287 36507 7293
rect 27522 7256 27528 7268
rect 24320 7228 26648 7256
rect 26712 7228 27528 7256
rect 16540 7160 21404 7188
rect 16540 7148 16546 7160
rect 21818 7148 21824 7200
rect 21876 7188 21882 7200
rect 24394 7188 24400 7200
rect 21876 7160 24400 7188
rect 21876 7148 21882 7160
rect 24394 7148 24400 7160
rect 24452 7148 24458 7200
rect 24854 7188 24860 7200
rect 24815 7160 24860 7188
rect 24854 7148 24860 7160
rect 24912 7148 24918 7200
rect 26620 7188 26648 7228
rect 27522 7216 27528 7228
rect 27580 7216 27586 7268
rect 28994 7216 29000 7268
rect 29052 7256 29058 7268
rect 29273 7259 29331 7265
rect 29273 7256 29285 7259
rect 29052 7228 29285 7256
rect 29052 7216 29058 7228
rect 29273 7225 29285 7228
rect 29319 7225 29331 7259
rect 29273 7219 29331 7225
rect 28537 7191 28595 7197
rect 28537 7188 28549 7191
rect 26620 7160 28549 7188
rect 28537 7157 28549 7160
rect 28583 7188 28595 7191
rect 30742 7188 30748 7200
rect 28583 7160 30748 7188
rect 28583 7157 28595 7160
rect 28537 7151 28595 7157
rect 30742 7148 30748 7160
rect 30800 7148 30806 7200
rect 1104 7098 38824 7120
rect 1104 7046 19606 7098
rect 19658 7046 19670 7098
rect 19722 7046 19734 7098
rect 19786 7046 19798 7098
rect 19850 7046 38824 7098
rect 1104 7024 38824 7046
rect 7006 6944 7012 6996
rect 7064 6984 7070 6996
rect 7064 6956 11100 6984
rect 7064 6944 7070 6956
rect 5736 6888 6040 6916
rect 1857 6851 1915 6857
rect 1857 6817 1869 6851
rect 1903 6848 1915 6851
rect 2590 6848 2596 6860
rect 1903 6820 2596 6848
rect 1903 6817 1915 6820
rect 1857 6811 1915 6817
rect 2590 6808 2596 6820
rect 2648 6848 2654 6860
rect 4249 6851 4307 6857
rect 2648 6820 4016 6848
rect 2648 6808 2654 6820
rect 2130 6780 2136 6792
rect 2091 6752 2136 6780
rect 2130 6740 2136 6752
rect 2188 6740 2194 6792
rect 3418 6644 3424 6656
rect 3379 6616 3424 6644
rect 3418 6604 3424 6616
rect 3476 6604 3482 6656
rect 3988 6644 4016 6820
rect 4249 6817 4261 6851
rect 4295 6817 4307 6851
rect 4706 6848 4712 6860
rect 4667 6820 4712 6848
rect 4249 6811 4307 6817
rect 4154 6780 4160 6792
rect 4115 6752 4160 6780
rect 4154 6740 4160 6752
rect 4212 6740 4218 6792
rect 4264 6712 4292 6811
rect 4706 6808 4712 6820
rect 4764 6808 4770 6860
rect 5077 6851 5135 6857
rect 5077 6817 5089 6851
rect 5123 6817 5135 6851
rect 5077 6811 5135 6817
rect 5445 6851 5503 6857
rect 5445 6817 5457 6851
rect 5491 6848 5503 6851
rect 5736 6848 5764 6888
rect 5902 6848 5908 6860
rect 5491 6820 5764 6848
rect 5863 6820 5908 6848
rect 5491 6817 5503 6820
rect 5445 6811 5503 6817
rect 4614 6740 4620 6792
rect 4672 6780 4678 6792
rect 5092 6780 5120 6811
rect 5902 6808 5908 6820
rect 5960 6808 5966 6860
rect 6012 6848 6040 6888
rect 7466 6876 7472 6928
rect 7524 6916 7530 6928
rect 10873 6919 10931 6925
rect 7524 6888 8616 6916
rect 7524 6876 7530 6888
rect 6730 6848 6736 6860
rect 6012 6820 6592 6848
rect 6691 6820 6736 6848
rect 6178 6780 6184 6792
rect 4672 6752 6184 6780
rect 4672 6740 4678 6752
rect 6178 6740 6184 6752
rect 6236 6740 6242 6792
rect 6454 6780 6460 6792
rect 6415 6752 6460 6780
rect 6454 6740 6460 6752
rect 6512 6740 6518 6792
rect 6564 6780 6592 6820
rect 6730 6808 6736 6820
rect 6788 6808 6794 6860
rect 8588 6857 8616 6888
rect 10873 6885 10885 6919
rect 10919 6916 10931 6919
rect 10962 6916 10968 6928
rect 10919 6888 10968 6916
rect 10919 6885 10931 6888
rect 10873 6879 10931 6885
rect 10962 6876 10968 6888
rect 11020 6876 11026 6928
rect 11072 6916 11100 6956
rect 11698 6944 11704 6996
rect 11756 6984 11762 6996
rect 11793 6987 11851 6993
rect 11793 6984 11805 6987
rect 11756 6956 11805 6984
rect 11756 6944 11762 6956
rect 11793 6953 11805 6956
rect 11839 6953 11851 6987
rect 11793 6947 11851 6953
rect 15930 6944 15936 6996
rect 15988 6984 15994 6996
rect 16485 6987 16543 6993
rect 16485 6984 16497 6987
rect 15988 6956 16497 6984
rect 15988 6944 15994 6956
rect 16485 6953 16497 6956
rect 16531 6953 16543 6987
rect 16485 6947 16543 6953
rect 20254 6944 20260 6996
rect 20312 6984 20318 6996
rect 21542 6984 21548 6996
rect 20312 6956 21548 6984
rect 20312 6944 20318 6956
rect 21542 6944 21548 6956
rect 21600 6944 21606 6996
rect 21910 6944 21916 6996
rect 21968 6984 21974 6996
rect 23658 6984 23664 6996
rect 21968 6956 23664 6984
rect 21968 6944 21974 6956
rect 23658 6944 23664 6956
rect 23716 6984 23722 6996
rect 31938 6984 31944 6996
rect 23716 6956 31944 6984
rect 23716 6944 23722 6956
rect 31938 6944 31944 6956
rect 31996 6944 32002 6996
rect 32122 6944 32128 6996
rect 32180 6944 32186 6996
rect 36354 6944 36360 6996
rect 36412 6984 36418 6996
rect 36449 6987 36507 6993
rect 36449 6984 36461 6987
rect 36412 6956 36461 6984
rect 36412 6944 36418 6956
rect 36449 6953 36461 6956
rect 36495 6953 36507 6987
rect 36449 6947 36507 6953
rect 12158 6916 12164 6928
rect 11072 6888 12164 6916
rect 12158 6876 12164 6888
rect 12216 6876 12222 6928
rect 15562 6876 15568 6928
rect 15620 6916 15626 6928
rect 19978 6916 19984 6928
rect 15620 6888 17632 6916
rect 15620 6876 15626 6888
rect 8579 6851 8637 6857
rect 8579 6817 8591 6851
rect 8625 6817 8637 6851
rect 10134 6848 10140 6860
rect 10095 6820 10140 6848
rect 8579 6811 8637 6817
rect 10134 6808 10140 6820
rect 10192 6808 10198 6860
rect 10226 6808 10232 6860
rect 10284 6848 10290 6860
rect 10597 6851 10655 6857
rect 10597 6848 10609 6851
rect 10284 6820 10609 6848
rect 10284 6808 10290 6820
rect 10597 6817 10609 6820
rect 10643 6817 10655 6851
rect 10597 6811 10655 6817
rect 11885 6851 11943 6857
rect 11885 6817 11897 6851
rect 11931 6817 11943 6851
rect 11885 6811 11943 6817
rect 12253 6851 12311 6857
rect 12253 6817 12265 6851
rect 12299 6817 12311 6851
rect 12253 6811 12311 6817
rect 11900 6780 11928 6811
rect 12158 6780 12164 6792
rect 6564 6752 8616 6780
rect 11900 6752 12164 6780
rect 5258 6712 5264 6724
rect 4264 6684 5264 6712
rect 5258 6672 5264 6684
rect 5316 6672 5322 6724
rect 4982 6644 4988 6656
rect 3988 6616 4988 6644
rect 4982 6604 4988 6616
rect 5040 6604 5046 6656
rect 5074 6604 5080 6656
rect 5132 6644 5138 6656
rect 7837 6647 7895 6653
rect 7837 6644 7849 6647
rect 5132 6616 7849 6644
rect 5132 6604 5138 6616
rect 7837 6613 7849 6616
rect 7883 6613 7895 6647
rect 8588 6644 8616 6752
rect 12158 6740 12164 6752
rect 12216 6740 12222 6792
rect 8757 6715 8815 6721
rect 8757 6681 8769 6715
rect 8803 6712 8815 6715
rect 8938 6712 8944 6724
rect 8803 6684 8944 6712
rect 8803 6681 8815 6684
rect 8757 6675 8815 6681
rect 8938 6672 8944 6684
rect 8996 6712 9002 6724
rect 12268 6712 12296 6811
rect 12434 6808 12440 6860
rect 12492 6848 12498 6860
rect 13633 6851 13691 6857
rect 13633 6848 13645 6851
rect 12492 6820 13645 6848
rect 12492 6808 12498 6820
rect 13633 6817 13645 6820
rect 13679 6848 13691 6851
rect 13906 6848 13912 6860
rect 13679 6820 13912 6848
rect 13679 6817 13691 6820
rect 13633 6811 13691 6817
rect 13906 6808 13912 6820
rect 13964 6808 13970 6860
rect 14001 6851 14059 6857
rect 14001 6817 14013 6851
rect 14047 6848 14059 6851
rect 14090 6848 14096 6860
rect 14047 6820 14096 6848
rect 14047 6817 14059 6820
rect 14001 6811 14059 6817
rect 12526 6780 12532 6792
rect 12487 6752 12532 6780
rect 12526 6740 12532 6752
rect 12584 6740 12590 6792
rect 14016 6780 14044 6811
rect 14090 6808 14096 6820
rect 14148 6808 14154 6860
rect 15470 6848 15476 6860
rect 15431 6820 15476 6848
rect 15470 6808 15476 6820
rect 15528 6808 15534 6860
rect 15838 6848 15844 6860
rect 15799 6820 15844 6848
rect 15838 6808 15844 6820
rect 15896 6808 15902 6860
rect 16669 6851 16727 6857
rect 16669 6817 16681 6851
rect 16715 6817 16727 6851
rect 16850 6848 16856 6860
rect 16811 6820 16856 6848
rect 16669 6811 16727 6817
rect 14458 6780 14464 6792
rect 13004 6752 14044 6780
rect 14419 6752 14464 6780
rect 13004 6712 13032 6752
rect 14458 6740 14464 6752
rect 14516 6740 14522 6792
rect 15562 6740 15568 6792
rect 15620 6780 15626 6792
rect 16684 6780 16712 6811
rect 16850 6808 16856 6820
rect 16908 6808 16914 6860
rect 17310 6848 17316 6860
rect 17271 6820 17316 6848
rect 17310 6808 17316 6820
rect 17368 6808 17374 6860
rect 17494 6848 17500 6860
rect 17455 6820 17500 6848
rect 17494 6808 17500 6820
rect 17552 6808 17558 6860
rect 17604 6848 17632 6888
rect 18064 6888 18276 6916
rect 18064 6848 18092 6888
rect 17604 6820 18092 6848
rect 18141 6851 18199 6857
rect 18141 6817 18153 6851
rect 18187 6817 18199 6851
rect 18248 6848 18276 6888
rect 19720 6888 19984 6916
rect 18417 6851 18475 6857
rect 18417 6848 18429 6851
rect 18248 6820 18429 6848
rect 18141 6811 18199 6817
rect 18417 6817 18429 6820
rect 18463 6817 18475 6851
rect 18417 6811 18475 6817
rect 19429 6851 19487 6857
rect 19429 6817 19441 6851
rect 19475 6848 19487 6851
rect 19720 6848 19748 6888
rect 19978 6876 19984 6888
rect 20036 6876 20042 6928
rect 22002 6916 22008 6928
rect 20088 6888 22008 6916
rect 19475 6820 19748 6848
rect 19797 6851 19855 6857
rect 19475 6817 19487 6820
rect 19429 6811 19487 6817
rect 19797 6817 19809 6851
rect 19843 6848 19855 6851
rect 20088 6848 20116 6888
rect 22002 6876 22008 6888
rect 22060 6876 22066 6928
rect 29730 6916 29736 6928
rect 29472 6888 29736 6916
rect 19843 6820 20116 6848
rect 20165 6851 20223 6857
rect 19843 6817 19855 6820
rect 19797 6811 19855 6817
rect 20165 6817 20177 6851
rect 20211 6817 20223 6851
rect 20165 6811 20223 6817
rect 20901 6851 20959 6857
rect 20901 6817 20913 6851
rect 20947 6848 20959 6851
rect 21634 6848 21640 6860
rect 20947 6820 21640 6848
rect 20947 6817 20959 6820
rect 20901 6811 20959 6817
rect 18156 6780 18184 6811
rect 18230 6780 18236 6792
rect 15620 6752 16712 6780
rect 18143 6752 18236 6780
rect 15620 6740 15626 6752
rect 18230 6740 18236 6752
rect 18288 6780 18294 6792
rect 19245 6783 19303 6789
rect 19245 6780 19257 6783
rect 18288 6752 19257 6780
rect 18288 6740 18294 6752
rect 19245 6749 19257 6752
rect 19291 6749 19303 6783
rect 20180 6780 20208 6811
rect 21634 6808 21640 6820
rect 21692 6808 21698 6860
rect 21729 6851 21787 6857
rect 21729 6817 21741 6851
rect 21775 6848 21787 6851
rect 22462 6848 22468 6860
rect 21775 6820 22468 6848
rect 21775 6817 21787 6820
rect 21729 6811 21787 6817
rect 22462 6808 22468 6820
rect 22520 6808 22526 6860
rect 22557 6851 22615 6857
rect 22557 6817 22569 6851
rect 22603 6817 22615 6851
rect 22557 6811 22615 6817
rect 22094 6780 22100 6792
rect 20180 6752 22100 6780
rect 19245 6743 19303 6749
rect 22094 6740 22100 6752
rect 22152 6740 22158 6792
rect 22572 6780 22600 6811
rect 22646 6808 22652 6860
rect 22704 6848 22710 6860
rect 22833 6851 22891 6857
rect 22833 6848 22845 6851
rect 22704 6820 22845 6848
rect 22704 6808 22710 6820
rect 22833 6817 22845 6820
rect 22879 6817 22891 6851
rect 22833 6811 22891 6817
rect 23106 6808 23112 6860
rect 23164 6848 23170 6860
rect 23201 6851 23259 6857
rect 23201 6848 23213 6851
rect 23164 6820 23213 6848
rect 23164 6808 23170 6820
rect 23201 6817 23213 6820
rect 23247 6817 23259 6851
rect 23201 6811 23259 6817
rect 23382 6808 23388 6860
rect 23440 6848 23446 6860
rect 24213 6851 24271 6857
rect 24213 6848 24225 6851
rect 23440 6820 24225 6848
rect 23440 6808 23446 6820
rect 24213 6817 24225 6820
rect 24259 6817 24271 6851
rect 24213 6811 24271 6817
rect 24489 6851 24547 6857
rect 24489 6817 24501 6851
rect 24535 6848 24547 6851
rect 24854 6848 24860 6860
rect 24535 6820 24860 6848
rect 24535 6817 24547 6820
rect 24489 6811 24547 6817
rect 24854 6808 24860 6820
rect 24912 6808 24918 6860
rect 25682 6808 25688 6860
rect 25740 6848 25746 6860
rect 26605 6851 26663 6857
rect 26605 6848 26617 6851
rect 25740 6820 26617 6848
rect 25740 6808 25746 6820
rect 26605 6817 26617 6820
rect 26651 6817 26663 6851
rect 26605 6811 26663 6817
rect 27249 6851 27307 6857
rect 27249 6817 27261 6851
rect 27295 6817 27307 6851
rect 27249 6811 27307 6817
rect 24578 6780 24584 6792
rect 22572 6752 24584 6780
rect 24578 6740 24584 6752
rect 24636 6740 24642 6792
rect 25498 6740 25504 6792
rect 25556 6780 25562 6792
rect 25593 6783 25651 6789
rect 25593 6780 25605 6783
rect 25556 6752 25605 6780
rect 25556 6740 25562 6752
rect 25593 6749 25605 6752
rect 25639 6749 25651 6783
rect 27062 6780 27068 6792
rect 27023 6752 27068 6780
rect 25593 6743 25651 6749
rect 27062 6740 27068 6752
rect 27120 6740 27126 6792
rect 27264 6780 27292 6811
rect 27338 6808 27344 6860
rect 27396 6848 27402 6860
rect 27525 6851 27583 6857
rect 27525 6848 27537 6851
rect 27396 6820 27537 6848
rect 27396 6808 27402 6820
rect 27525 6817 27537 6820
rect 27571 6817 27583 6851
rect 27890 6848 27896 6860
rect 27851 6820 27896 6848
rect 27525 6811 27583 6817
rect 27890 6808 27896 6820
rect 27948 6808 27954 6860
rect 28813 6851 28871 6857
rect 28813 6817 28825 6851
rect 28859 6848 28871 6851
rect 28994 6848 29000 6860
rect 28859 6820 29000 6848
rect 28859 6817 28871 6820
rect 28813 6811 28871 6817
rect 28994 6808 29000 6820
rect 29052 6808 29058 6860
rect 29472 6857 29500 6888
rect 29730 6876 29736 6888
rect 29788 6876 29794 6928
rect 30834 6876 30840 6928
rect 30892 6916 30898 6928
rect 32140 6916 32168 6944
rect 32493 6919 32551 6925
rect 32493 6916 32505 6919
rect 30892 6888 31432 6916
rect 32140 6888 32505 6916
rect 30892 6876 30898 6888
rect 29181 6851 29239 6857
rect 29181 6817 29193 6851
rect 29227 6817 29239 6851
rect 29181 6811 29239 6817
rect 29457 6851 29515 6857
rect 29457 6817 29469 6851
rect 29503 6817 29515 6851
rect 29457 6811 29515 6817
rect 27430 6780 27436 6792
rect 27264 6752 27436 6780
rect 27430 6740 27436 6752
rect 27488 6740 27494 6792
rect 28166 6740 28172 6792
rect 28224 6780 28230 6792
rect 29196 6780 29224 6811
rect 29546 6808 29552 6860
rect 29604 6848 29610 6860
rect 31404 6857 31432 6888
rect 32493 6885 32505 6888
rect 32539 6885 32551 6919
rect 32493 6879 32551 6885
rect 33042 6876 33048 6928
rect 33100 6916 33106 6928
rect 36372 6916 36400 6944
rect 33100 6888 35756 6916
rect 33100 6876 33106 6888
rect 31021 6851 31079 6857
rect 31021 6848 31033 6851
rect 29604 6820 31033 6848
rect 29604 6808 29610 6820
rect 31021 6817 31033 6820
rect 31067 6817 31079 6851
rect 31021 6811 31079 6817
rect 31389 6851 31447 6857
rect 31389 6817 31401 6851
rect 31435 6817 31447 6851
rect 31389 6811 31447 6817
rect 28224 6752 29224 6780
rect 28224 6740 28230 6752
rect 29270 6740 29276 6792
rect 29328 6780 29334 6792
rect 31294 6780 31300 6792
rect 29328 6752 31300 6780
rect 29328 6740 29334 6752
rect 31294 6740 31300 6752
rect 31352 6740 31358 6792
rect 8996 6684 13032 6712
rect 8996 6672 9002 6684
rect 13078 6672 13084 6724
rect 13136 6712 13142 6724
rect 13541 6715 13599 6721
rect 13541 6712 13553 6715
rect 13136 6684 13553 6712
rect 13136 6672 13142 6684
rect 13541 6681 13553 6684
rect 13587 6681 13599 6715
rect 15378 6712 15384 6724
rect 15339 6684 15384 6712
rect 13541 6675 13599 6681
rect 15378 6672 15384 6684
rect 15436 6672 15442 6724
rect 16114 6672 16120 6724
rect 16172 6712 16178 6724
rect 16853 6715 16911 6721
rect 16853 6712 16865 6715
rect 16172 6684 16865 6712
rect 16172 6672 16178 6684
rect 16853 6681 16865 6684
rect 16899 6681 16911 6715
rect 16853 6675 16911 6681
rect 21818 6672 21824 6724
rect 21876 6712 21882 6724
rect 21913 6715 21971 6721
rect 21913 6712 21925 6715
rect 21876 6684 21925 6712
rect 21876 6672 21882 6684
rect 21913 6681 21925 6684
rect 21959 6681 21971 6715
rect 21913 6675 21971 6681
rect 28905 6715 28963 6721
rect 28905 6681 28917 6715
rect 28951 6681 28963 6715
rect 28905 6675 28963 6681
rect 30837 6715 30895 6721
rect 30837 6681 30849 6715
rect 30883 6712 30895 6715
rect 31018 6712 31024 6724
rect 30883 6684 31024 6712
rect 30883 6681 30895 6684
rect 30837 6675 30895 6681
rect 10502 6644 10508 6656
rect 8588 6616 10508 6644
rect 7837 6607 7895 6613
rect 10502 6604 10508 6616
rect 10560 6644 10566 6656
rect 15286 6644 15292 6656
rect 10560 6616 15292 6644
rect 10560 6604 10566 6616
rect 15286 6604 15292 6616
rect 15344 6604 15350 6656
rect 20530 6604 20536 6656
rect 20588 6644 20594 6656
rect 21085 6647 21143 6653
rect 21085 6644 21097 6647
rect 20588 6616 21097 6644
rect 20588 6604 20594 6616
rect 21085 6613 21097 6616
rect 21131 6613 21143 6647
rect 22554 6644 22560 6656
rect 22515 6616 22560 6644
rect 21085 6607 21143 6613
rect 22554 6604 22560 6616
rect 22612 6604 22618 6656
rect 28920 6644 28948 6675
rect 31018 6672 31024 6684
rect 31076 6672 31082 6724
rect 31404 6712 31432 6811
rect 31478 6808 31484 6860
rect 31536 6848 31542 6860
rect 31536 6820 31581 6848
rect 31536 6808 31542 6820
rect 31662 6808 31668 6860
rect 31720 6848 31726 6860
rect 32125 6851 32183 6857
rect 32125 6848 32137 6851
rect 31720 6820 32137 6848
rect 31720 6808 31726 6820
rect 32125 6817 32137 6820
rect 32171 6817 32183 6851
rect 32306 6848 32312 6860
rect 32267 6820 32312 6848
rect 32125 6811 32183 6817
rect 32306 6808 32312 6820
rect 32364 6808 32370 6860
rect 32401 6851 32459 6857
rect 32401 6817 32413 6851
rect 32447 6817 32459 6851
rect 32401 6811 32459 6817
rect 32861 6851 32919 6857
rect 32861 6817 32873 6851
rect 32907 6848 32919 6851
rect 33594 6848 33600 6860
rect 32907 6820 33600 6848
rect 32907 6817 32919 6820
rect 32861 6811 32919 6817
rect 31570 6740 31576 6792
rect 31628 6780 31634 6792
rect 32416 6780 32444 6811
rect 33594 6808 33600 6820
rect 33652 6808 33658 6860
rect 34238 6848 34244 6860
rect 34199 6820 34244 6848
rect 34238 6808 34244 6820
rect 34296 6808 34302 6860
rect 35728 6857 35756 6888
rect 35912 6888 36400 6916
rect 35713 6851 35771 6857
rect 35713 6817 35725 6851
rect 35759 6817 35771 6851
rect 35713 6811 35771 6817
rect 31628 6752 32444 6780
rect 31628 6740 31634 6752
rect 32490 6740 32496 6792
rect 32548 6780 32554 6792
rect 33413 6783 33471 6789
rect 33413 6780 33425 6783
rect 32548 6752 33425 6780
rect 32548 6740 32554 6752
rect 33413 6749 33425 6752
rect 33459 6749 33471 6783
rect 33962 6780 33968 6792
rect 33923 6752 33968 6780
rect 33413 6743 33471 6749
rect 33962 6740 33968 6752
rect 34020 6740 34026 6792
rect 34425 6783 34483 6789
rect 34425 6749 34437 6783
rect 34471 6780 34483 6783
rect 34514 6780 34520 6792
rect 34471 6752 34520 6780
rect 34471 6749 34483 6752
rect 34425 6743 34483 6749
rect 34514 6740 34520 6752
rect 34572 6740 34578 6792
rect 34698 6740 34704 6792
rect 34756 6780 34762 6792
rect 34885 6783 34943 6789
rect 34885 6780 34897 6783
rect 34756 6752 34897 6780
rect 34756 6740 34762 6752
rect 34885 6749 34897 6752
rect 34931 6749 34943 6783
rect 35434 6780 35440 6792
rect 35395 6752 35440 6780
rect 34885 6743 34943 6749
rect 35434 6740 35440 6752
rect 35492 6740 35498 6792
rect 35728 6780 35756 6811
rect 35802 6808 35808 6860
rect 35860 6848 35866 6860
rect 35912 6857 35940 6888
rect 35897 6851 35955 6857
rect 35897 6848 35909 6851
rect 35860 6820 35909 6848
rect 35860 6808 35866 6820
rect 35897 6817 35909 6820
rect 35943 6817 35955 6851
rect 35897 6811 35955 6817
rect 35986 6808 35992 6860
rect 36044 6848 36050 6860
rect 36357 6851 36415 6857
rect 36357 6848 36369 6851
rect 36044 6820 36369 6848
rect 36044 6808 36050 6820
rect 36357 6817 36369 6820
rect 36403 6817 36415 6851
rect 36357 6811 36415 6817
rect 37366 6780 37372 6792
rect 35728 6752 37372 6780
rect 37366 6740 37372 6752
rect 37424 6740 37430 6792
rect 31404 6684 32812 6712
rect 29546 6644 29552 6656
rect 28920 6616 29552 6644
rect 29546 6604 29552 6616
rect 29604 6604 29610 6656
rect 29730 6604 29736 6656
rect 29788 6644 29794 6656
rect 32214 6644 32220 6656
rect 29788 6616 32220 6644
rect 29788 6604 29794 6616
rect 32214 6604 32220 6616
rect 32272 6604 32278 6656
rect 32784 6644 32812 6684
rect 33226 6644 33232 6656
rect 32784 6616 33232 6644
rect 33226 6604 33232 6616
rect 33284 6644 33290 6656
rect 33686 6644 33692 6656
rect 33284 6616 33692 6644
rect 33284 6604 33290 6616
rect 33686 6604 33692 6616
rect 33744 6604 33750 6656
rect 1104 6554 38824 6576
rect 1104 6502 4246 6554
rect 4298 6502 4310 6554
rect 4362 6502 4374 6554
rect 4426 6502 4438 6554
rect 4490 6502 34966 6554
rect 35018 6502 35030 6554
rect 35082 6502 35094 6554
rect 35146 6502 35158 6554
rect 35210 6502 38824 6554
rect 1104 6480 38824 6502
rect 4908 6412 8524 6440
rect 2130 6332 2136 6384
rect 2188 6372 2194 6384
rect 3513 6375 3571 6381
rect 3513 6372 3525 6375
rect 2188 6344 3525 6372
rect 2188 6332 2194 6344
rect 3513 6341 3525 6344
rect 3559 6341 3571 6375
rect 3513 6335 3571 6341
rect 2332 6276 3924 6304
rect 1854 6236 1860 6248
rect 1815 6208 1860 6236
rect 1854 6196 1860 6208
rect 1912 6196 1918 6248
rect 2332 6245 2360 6276
rect 3896 6245 3924 6276
rect 2317 6239 2375 6245
rect 2317 6205 2329 6239
rect 2363 6205 2375 6239
rect 2317 6199 2375 6205
rect 3605 6239 3663 6245
rect 3605 6205 3617 6239
rect 3651 6205 3663 6239
rect 3605 6199 3663 6205
rect 3881 6239 3939 6245
rect 3881 6205 3893 6239
rect 3927 6236 3939 6239
rect 4062 6236 4068 6248
rect 3927 6208 4068 6236
rect 3927 6205 3939 6208
rect 3881 6199 3939 6205
rect 3620 6168 3648 6199
rect 4062 6196 4068 6208
rect 4120 6196 4126 6248
rect 4433 6239 4491 6245
rect 4433 6205 4445 6239
rect 4479 6236 4491 6239
rect 4614 6236 4620 6248
rect 4479 6208 4620 6236
rect 4479 6205 4491 6208
rect 4433 6199 4491 6205
rect 4614 6196 4620 6208
rect 4672 6196 4678 6248
rect 4801 6239 4859 6245
rect 4801 6205 4813 6239
rect 4847 6236 4859 6239
rect 4908 6236 4936 6412
rect 8496 6372 8524 6412
rect 8570 6400 8576 6452
rect 8628 6440 8634 6452
rect 12526 6440 12532 6452
rect 8628 6412 12532 6440
rect 8628 6400 8634 6412
rect 12526 6400 12532 6412
rect 12584 6400 12590 6452
rect 15286 6400 15292 6452
rect 15344 6440 15350 6452
rect 21453 6443 21511 6449
rect 21453 6440 21465 6443
rect 15344 6412 21465 6440
rect 15344 6400 15350 6412
rect 21453 6409 21465 6412
rect 21499 6409 21511 6443
rect 21453 6403 21511 6409
rect 24673 6443 24731 6449
rect 24673 6409 24685 6443
rect 24719 6440 24731 6443
rect 25130 6440 25136 6452
rect 24719 6412 25136 6440
rect 24719 6409 24731 6412
rect 24673 6403 24731 6409
rect 25130 6400 25136 6412
rect 25188 6400 25194 6452
rect 27430 6400 27436 6452
rect 27488 6440 27494 6452
rect 30837 6443 30895 6449
rect 27488 6412 30788 6440
rect 27488 6400 27494 6412
rect 13262 6372 13268 6384
rect 8496 6344 13268 6372
rect 13262 6332 13268 6344
rect 13320 6332 13326 6384
rect 14734 6372 14740 6384
rect 14384 6344 14740 6372
rect 4982 6264 4988 6316
rect 5040 6304 5046 6316
rect 5534 6304 5540 6316
rect 5040 6276 5540 6304
rect 5040 6264 5046 6276
rect 5534 6264 5540 6276
rect 5592 6304 5598 6316
rect 6454 6304 6460 6316
rect 5592 6276 6460 6304
rect 5592 6264 5598 6276
rect 6454 6264 6460 6276
rect 6512 6304 6518 6316
rect 7837 6307 7895 6313
rect 6512 6276 7512 6304
rect 6512 6264 6518 6276
rect 7484 6248 7512 6276
rect 7837 6273 7849 6307
rect 7883 6304 7895 6307
rect 7926 6304 7932 6316
rect 7883 6276 7932 6304
rect 7883 6273 7895 6276
rect 7837 6267 7895 6273
rect 7926 6264 7932 6276
rect 7984 6264 7990 6316
rect 9490 6264 9496 6316
rect 9548 6304 9554 6316
rect 13357 6307 13415 6313
rect 9548 6276 10548 6304
rect 9548 6264 9554 6276
rect 4847 6208 4936 6236
rect 5353 6239 5411 6245
rect 4847 6205 4859 6208
rect 4801 6199 4859 6205
rect 5353 6205 5365 6239
rect 5399 6205 5411 6239
rect 5353 6199 5411 6205
rect 5813 6239 5871 6245
rect 5813 6205 5825 6239
rect 5859 6236 5871 6239
rect 5994 6236 6000 6248
rect 5859 6208 6000 6236
rect 5859 6205 5871 6208
rect 5813 6199 5871 6205
rect 5258 6168 5264 6180
rect 3620 6140 5264 6168
rect 5258 6128 5264 6140
rect 5316 6128 5322 6180
rect 5368 6168 5396 6199
rect 5994 6196 6000 6208
rect 6052 6196 6058 6248
rect 6825 6239 6883 6245
rect 6825 6205 6837 6239
rect 6871 6236 6883 6239
rect 7006 6236 7012 6248
rect 6871 6208 7012 6236
rect 6871 6205 6883 6208
rect 6825 6199 6883 6205
rect 7006 6196 7012 6208
rect 7064 6196 7070 6248
rect 7466 6196 7472 6248
rect 7524 6236 7530 6248
rect 7561 6239 7619 6245
rect 7561 6236 7573 6239
rect 7524 6208 7573 6236
rect 7524 6196 7530 6208
rect 7561 6205 7573 6208
rect 7607 6205 7619 6239
rect 10134 6236 10140 6248
rect 10095 6208 10140 6236
rect 7561 6199 7619 6205
rect 10134 6196 10140 6208
rect 10192 6196 10198 6248
rect 10413 6239 10471 6245
rect 10413 6205 10425 6239
rect 10459 6205 10471 6239
rect 10520 6236 10548 6276
rect 13357 6273 13369 6307
rect 13403 6304 13415 6307
rect 14384 6304 14412 6344
rect 14734 6332 14740 6344
rect 14792 6332 14798 6384
rect 20162 6372 20168 6384
rect 20123 6344 20168 6372
rect 20162 6332 20168 6344
rect 20220 6332 20226 6384
rect 29270 6332 29276 6384
rect 29328 6332 29334 6384
rect 30760 6372 30788 6412
rect 30837 6409 30849 6443
rect 30883 6440 30895 6443
rect 30926 6440 30932 6452
rect 30883 6412 30932 6440
rect 30883 6409 30895 6412
rect 30837 6403 30895 6409
rect 30926 6400 30932 6412
rect 30984 6400 30990 6452
rect 31202 6400 31208 6452
rect 31260 6440 31266 6452
rect 37734 6440 37740 6452
rect 31260 6412 37740 6440
rect 31260 6400 31266 6412
rect 37734 6400 37740 6412
rect 37792 6440 37798 6452
rect 38013 6443 38071 6449
rect 38013 6440 38025 6443
rect 37792 6412 38025 6440
rect 37792 6400 37798 6412
rect 38013 6409 38025 6412
rect 38059 6409 38071 6443
rect 38013 6403 38071 6409
rect 32306 6372 32312 6384
rect 30760 6344 32312 6372
rect 32306 6332 32312 6344
rect 32364 6332 32370 6384
rect 32490 6372 32496 6384
rect 32416 6344 32496 6372
rect 13403 6276 14412 6304
rect 13403 6273 13415 6276
rect 13357 6267 13415 6273
rect 14458 6264 14464 6316
rect 14516 6304 14522 6316
rect 16114 6304 16120 6316
rect 14516 6276 15976 6304
rect 16075 6276 16120 6304
rect 14516 6264 14522 6276
rect 11149 6239 11207 6245
rect 11149 6236 11161 6239
rect 10520 6208 11161 6236
rect 10413 6199 10471 6205
rect 11149 6205 11161 6208
rect 11195 6205 11207 6239
rect 11149 6199 11207 6205
rect 5902 6168 5908 6180
rect 5368 6140 5908 6168
rect 5902 6128 5908 6140
rect 5960 6168 5966 6180
rect 10428 6168 10456 6199
rect 11238 6196 11244 6248
rect 11296 6236 11302 6248
rect 11701 6239 11759 6245
rect 11701 6236 11713 6239
rect 11296 6208 11713 6236
rect 11296 6196 11302 6208
rect 11701 6205 11713 6208
rect 11747 6236 11759 6239
rect 11974 6236 11980 6248
rect 11747 6208 11980 6236
rect 11747 6205 11759 6208
rect 11701 6199 11759 6205
rect 11974 6196 11980 6208
rect 12032 6196 12038 6248
rect 12434 6196 12440 6248
rect 12492 6236 12498 6248
rect 12492 6208 12537 6236
rect 12492 6196 12498 6208
rect 12710 6196 12716 6248
rect 12768 6236 12774 6248
rect 13265 6239 13323 6245
rect 13265 6236 13277 6239
rect 12768 6208 13277 6236
rect 12768 6196 12774 6208
rect 13265 6205 13277 6208
rect 13311 6205 13323 6239
rect 13265 6199 13323 6205
rect 13633 6239 13691 6245
rect 13633 6205 13645 6239
rect 13679 6236 13691 6239
rect 13906 6236 13912 6248
rect 13679 6208 13912 6236
rect 13679 6205 13691 6208
rect 13633 6199 13691 6205
rect 13906 6196 13912 6208
rect 13964 6196 13970 6248
rect 15562 6236 15568 6248
rect 14476 6208 15568 6236
rect 5960 6140 6868 6168
rect 5960 6128 5966 6140
rect 6840 6112 6868 6140
rect 8496 6140 10456 6168
rect 1670 6060 1676 6112
rect 1728 6100 1734 6112
rect 1857 6103 1915 6109
rect 1857 6100 1869 6103
rect 1728 6072 1869 6100
rect 1728 6060 1734 6072
rect 1857 6069 1869 6072
rect 1903 6069 1915 6103
rect 5994 6100 6000 6112
rect 5955 6072 6000 6100
rect 1857 6063 1915 6069
rect 5994 6060 6000 6072
rect 6052 6060 6058 6112
rect 6822 6060 6828 6112
rect 6880 6100 6886 6112
rect 7009 6103 7067 6109
rect 7009 6100 7021 6103
rect 6880 6072 7021 6100
rect 6880 6060 6886 6072
rect 7009 6069 7021 6072
rect 7055 6069 7067 6103
rect 7009 6063 7067 6069
rect 7282 6060 7288 6112
rect 7340 6100 7346 6112
rect 8496 6100 8524 6140
rect 10594 6128 10600 6180
rect 10652 6168 10658 6180
rect 10689 6171 10747 6177
rect 10689 6168 10701 6171
rect 10652 6140 10701 6168
rect 10652 6128 10658 6140
rect 10689 6137 10701 6140
rect 10735 6137 10747 6171
rect 10689 6131 10747 6137
rect 11885 6171 11943 6177
rect 11885 6137 11897 6171
rect 11931 6168 11943 6171
rect 12802 6168 12808 6180
rect 11931 6140 12808 6168
rect 11931 6137 11943 6140
rect 11885 6131 11943 6137
rect 12802 6128 12808 6140
rect 12860 6128 12866 6180
rect 7340 6072 8524 6100
rect 9125 6103 9183 6109
rect 7340 6060 7346 6072
rect 9125 6069 9137 6103
rect 9171 6100 9183 6103
rect 9674 6100 9680 6112
rect 9171 6072 9680 6100
rect 9171 6069 9183 6072
rect 9125 6063 9183 6069
rect 9674 6060 9680 6072
rect 9732 6060 9738 6112
rect 10226 6060 10232 6112
rect 10284 6100 10290 6112
rect 12529 6103 12587 6109
rect 12529 6100 12541 6103
rect 10284 6072 12541 6100
rect 10284 6060 10290 6072
rect 12529 6069 12541 6072
rect 12575 6069 12587 6103
rect 12529 6063 12587 6069
rect 13081 6103 13139 6109
rect 13081 6069 13093 6103
rect 13127 6100 13139 6103
rect 14476 6100 14504 6208
rect 15562 6196 15568 6208
rect 15620 6236 15626 6248
rect 15657 6239 15715 6245
rect 15657 6236 15669 6239
rect 15620 6208 15669 6236
rect 15620 6196 15626 6208
rect 15657 6205 15669 6208
rect 15703 6205 15715 6239
rect 15657 6199 15715 6205
rect 15749 6239 15807 6245
rect 15749 6205 15761 6239
rect 15795 6236 15807 6239
rect 15841 6239 15899 6245
rect 15841 6236 15853 6239
rect 15795 6208 15853 6236
rect 15795 6205 15807 6208
rect 15749 6199 15807 6205
rect 15841 6205 15853 6208
rect 15887 6205 15899 6239
rect 15948 6236 15976 6276
rect 16114 6264 16120 6276
rect 16172 6264 16178 6316
rect 17221 6307 17279 6313
rect 17221 6273 17233 6307
rect 17267 6273 17279 6307
rect 17221 6267 17279 6273
rect 28721 6307 28779 6313
rect 28721 6273 28733 6307
rect 28767 6304 28779 6307
rect 29288 6304 29316 6332
rect 29546 6304 29552 6316
rect 28767 6276 29316 6304
rect 29507 6276 29552 6304
rect 28767 6273 28779 6276
rect 28721 6267 28779 6273
rect 17236 6236 17264 6267
rect 29546 6264 29552 6276
rect 29604 6264 29610 6316
rect 30190 6264 30196 6316
rect 30248 6304 30254 6316
rect 31202 6304 31208 6316
rect 30248 6276 31208 6304
rect 30248 6264 30254 6276
rect 31202 6264 31208 6276
rect 31260 6264 31266 6316
rect 31849 6307 31907 6313
rect 31849 6273 31861 6307
rect 31895 6304 31907 6307
rect 32214 6304 32220 6316
rect 31895 6276 32220 6304
rect 31895 6273 31907 6276
rect 31849 6267 31907 6273
rect 32214 6264 32220 6276
rect 32272 6264 32278 6316
rect 32416 6313 32444 6344
rect 32490 6332 32496 6344
rect 32548 6332 32554 6384
rect 34514 6372 34520 6384
rect 34348 6344 34520 6372
rect 32401 6307 32459 6313
rect 32401 6273 32413 6307
rect 32447 6273 32459 6307
rect 32861 6307 32919 6313
rect 32861 6304 32873 6307
rect 32401 6267 32459 6273
rect 32508 6276 32873 6304
rect 18049 6239 18107 6245
rect 18049 6236 18061 6239
rect 15948 6208 18061 6236
rect 15841 6199 15899 6205
rect 18049 6205 18061 6208
rect 18095 6205 18107 6239
rect 18049 6199 18107 6205
rect 18785 6239 18843 6245
rect 18785 6205 18797 6239
rect 18831 6205 18843 6239
rect 18785 6199 18843 6205
rect 19061 6239 19119 6245
rect 19061 6205 19073 6239
rect 19107 6236 19119 6239
rect 19150 6236 19156 6248
rect 19107 6208 19156 6236
rect 19107 6205 19119 6208
rect 19061 6199 19119 6205
rect 18800 6168 18828 6199
rect 19150 6196 19156 6208
rect 19208 6196 19214 6248
rect 21358 6236 21364 6248
rect 21319 6208 21364 6236
rect 21358 6196 21364 6208
rect 21416 6196 21422 6248
rect 22002 6236 22008 6248
rect 21963 6208 22008 6236
rect 22002 6196 22008 6208
rect 22060 6196 22066 6248
rect 22373 6239 22431 6245
rect 22373 6205 22385 6239
rect 22419 6236 22431 6239
rect 22830 6236 22836 6248
rect 22419 6208 22836 6236
rect 22419 6205 22431 6208
rect 22373 6199 22431 6205
rect 22830 6196 22836 6208
rect 22888 6196 22894 6248
rect 23566 6196 23572 6248
rect 23624 6236 23630 6248
rect 23661 6239 23719 6245
rect 23661 6236 23673 6239
rect 23624 6208 23673 6236
rect 23624 6196 23630 6208
rect 23661 6205 23673 6208
rect 23707 6205 23719 6239
rect 24489 6239 24547 6245
rect 24489 6236 24501 6239
rect 23661 6199 23719 6205
rect 23860 6208 24501 6236
rect 17236 6140 18828 6168
rect 13127 6072 14504 6100
rect 13127 6069 13139 6072
rect 13081 6063 13139 6069
rect 14550 6060 14556 6112
rect 14608 6100 14614 6112
rect 14737 6103 14795 6109
rect 14737 6100 14749 6103
rect 14608 6072 14749 6100
rect 14608 6060 14614 6072
rect 14737 6069 14749 6072
rect 14783 6069 14795 6103
rect 14737 6063 14795 6069
rect 14826 6060 14832 6112
rect 14884 6100 14890 6112
rect 15473 6103 15531 6109
rect 15473 6100 15485 6103
rect 14884 6072 15485 6100
rect 14884 6060 14890 6072
rect 15473 6069 15485 6072
rect 15519 6100 15531 6103
rect 15749 6103 15807 6109
rect 15749 6100 15761 6103
rect 15519 6072 15761 6100
rect 15519 6069 15531 6072
rect 15473 6063 15531 6069
rect 15749 6069 15761 6072
rect 15795 6100 15807 6103
rect 17236 6100 17264 6140
rect 15795 6072 17264 6100
rect 15795 6069 15807 6072
rect 15749 6063 15807 6069
rect 17310 6060 17316 6112
rect 17368 6100 17374 6112
rect 18141 6103 18199 6109
rect 18141 6100 18153 6103
rect 17368 6072 18153 6100
rect 17368 6060 17374 6072
rect 18141 6069 18153 6072
rect 18187 6069 18199 6103
rect 18141 6063 18199 6069
rect 23658 6060 23664 6112
rect 23716 6100 23722 6112
rect 23860 6109 23888 6208
rect 24489 6205 24501 6208
rect 24535 6205 24547 6239
rect 24489 6199 24547 6205
rect 25130 6196 25136 6248
rect 25188 6236 25194 6248
rect 25225 6239 25283 6245
rect 25225 6236 25237 6239
rect 25188 6208 25237 6236
rect 25188 6196 25194 6208
rect 25225 6205 25237 6208
rect 25271 6205 25283 6239
rect 25225 6199 25283 6205
rect 25314 6196 25320 6248
rect 25372 6236 25378 6248
rect 25501 6239 25559 6245
rect 25501 6236 25513 6239
rect 25372 6208 25513 6236
rect 25372 6196 25378 6208
rect 25501 6205 25513 6208
rect 25547 6205 25559 6239
rect 25501 6199 25559 6205
rect 26881 6239 26939 6245
rect 26881 6205 26893 6239
rect 26927 6236 26939 6239
rect 27890 6236 27896 6248
rect 26927 6208 27896 6236
rect 26927 6205 26939 6208
rect 26881 6199 26939 6205
rect 27890 6196 27896 6208
rect 27948 6196 27954 6248
rect 27982 6196 27988 6248
rect 28040 6236 28046 6248
rect 28261 6239 28319 6245
rect 28261 6236 28273 6239
rect 28040 6208 28273 6236
rect 28040 6196 28046 6208
rect 28261 6205 28273 6208
rect 28307 6205 28319 6239
rect 28534 6236 28540 6248
rect 28495 6208 28540 6236
rect 28261 6199 28319 6205
rect 28534 6196 28540 6208
rect 28592 6196 28598 6248
rect 29178 6196 29184 6248
rect 29236 6236 29242 6248
rect 29273 6239 29331 6245
rect 29273 6236 29285 6239
rect 29236 6208 29285 6236
rect 29236 6196 29242 6208
rect 29273 6205 29285 6208
rect 29319 6205 29331 6239
rect 30558 6236 30564 6248
rect 29273 6199 29331 6205
rect 29380 6208 30564 6236
rect 27706 6168 27712 6180
rect 27667 6140 27712 6168
rect 27706 6128 27712 6140
rect 27764 6128 27770 6180
rect 27798 6128 27804 6180
rect 27856 6168 27862 6180
rect 29380 6168 29408 6208
rect 30558 6196 30564 6208
rect 30616 6196 30622 6248
rect 31938 6196 31944 6248
rect 31996 6236 32002 6248
rect 32508 6236 32536 6276
rect 32861 6273 32873 6276
rect 32907 6304 32919 6307
rect 33042 6304 33048 6316
rect 32907 6276 33048 6304
rect 32907 6273 32919 6276
rect 32861 6267 32919 6273
rect 33042 6264 33048 6276
rect 33100 6264 33106 6316
rect 34348 6313 34376 6344
rect 34514 6332 34520 6344
rect 34572 6372 34578 6384
rect 35710 6372 35716 6384
rect 34572 6344 35716 6372
rect 34572 6332 34578 6344
rect 35710 6332 35716 6344
rect 35768 6332 35774 6384
rect 34333 6307 34391 6313
rect 33796 6276 34192 6304
rect 31996 6208 32536 6236
rect 32677 6239 32735 6245
rect 31996 6196 32002 6208
rect 32677 6205 32689 6239
rect 32723 6205 32735 6239
rect 33796 6236 33824 6276
rect 34164 6248 34192 6276
rect 34333 6273 34345 6307
rect 34379 6273 34391 6307
rect 34333 6267 34391 6273
rect 34977 6307 35035 6313
rect 34977 6273 34989 6307
rect 35023 6304 35035 6307
rect 35434 6304 35440 6316
rect 35023 6276 35440 6304
rect 35023 6273 35035 6276
rect 34977 6267 35035 6273
rect 35434 6264 35440 6276
rect 35492 6264 35498 6316
rect 35894 6264 35900 6316
rect 35952 6304 35958 6316
rect 35989 6307 36047 6313
rect 35989 6304 36001 6307
rect 35952 6276 36001 6304
rect 35952 6264 35958 6276
rect 35989 6273 36001 6276
rect 36035 6273 36047 6307
rect 35989 6267 36047 6273
rect 32677 6199 32735 6205
rect 33152 6208 33824 6236
rect 33873 6239 33931 6245
rect 27856 6140 29408 6168
rect 32692 6168 32720 6199
rect 33152 6168 33180 6208
rect 33873 6205 33885 6239
rect 33919 6205 33931 6239
rect 34146 6236 34152 6248
rect 34059 6208 34152 6236
rect 33873 6199 33931 6205
rect 33318 6168 33324 6180
rect 32692 6140 33180 6168
rect 33279 6140 33324 6168
rect 27856 6128 27862 6140
rect 33318 6128 33324 6140
rect 33376 6128 33382 6180
rect 33888 6168 33916 6199
rect 34146 6196 34152 6208
rect 34204 6196 34210 6248
rect 34514 6196 34520 6248
rect 34572 6236 34578 6248
rect 35526 6236 35532 6248
rect 34572 6208 35532 6236
rect 34572 6196 34578 6208
rect 35526 6196 35532 6208
rect 35584 6196 35590 6248
rect 35618 6196 35624 6248
rect 35676 6236 35682 6248
rect 35805 6239 35863 6245
rect 35805 6236 35817 6239
rect 35676 6208 35817 6236
rect 35676 6196 35682 6208
rect 35805 6205 35817 6208
rect 35851 6236 35863 6239
rect 36078 6236 36084 6248
rect 35851 6208 36084 6236
rect 35851 6205 35863 6208
rect 35805 6199 35863 6205
rect 36078 6196 36084 6208
rect 36136 6196 36142 6248
rect 36998 6236 37004 6248
rect 36959 6208 37004 6236
rect 36998 6196 37004 6208
rect 37056 6196 37062 6248
rect 37274 6236 37280 6248
rect 37235 6208 37280 6236
rect 37274 6196 37280 6208
rect 37332 6196 37338 6248
rect 37458 6236 37464 6248
rect 37419 6208 37464 6236
rect 37458 6196 37464 6208
rect 37516 6196 37522 6248
rect 37550 6196 37556 6248
rect 37608 6236 37614 6248
rect 37921 6239 37979 6245
rect 37921 6236 37933 6239
rect 37608 6208 37933 6236
rect 37608 6196 37614 6208
rect 37921 6205 37933 6208
rect 37967 6205 37979 6239
rect 37921 6199 37979 6205
rect 36449 6171 36507 6177
rect 36449 6168 36461 6171
rect 33888 6140 36461 6168
rect 36449 6137 36461 6140
rect 36495 6137 36507 6171
rect 36449 6131 36507 6137
rect 23845 6103 23903 6109
rect 23845 6100 23857 6103
rect 23716 6072 23857 6100
rect 23716 6060 23722 6072
rect 23845 6069 23857 6072
rect 23891 6069 23903 6103
rect 23845 6063 23903 6069
rect 29086 6060 29092 6112
rect 29144 6100 29150 6112
rect 29638 6100 29644 6112
rect 29144 6072 29644 6100
rect 29144 6060 29150 6072
rect 29638 6060 29644 6072
rect 29696 6100 29702 6112
rect 30466 6100 30472 6112
rect 29696 6072 30472 6100
rect 29696 6060 29702 6072
rect 30466 6060 30472 6072
rect 30524 6060 30530 6112
rect 32214 6060 32220 6112
rect 32272 6100 32278 6112
rect 35618 6100 35624 6112
rect 32272 6072 35624 6100
rect 32272 6060 32278 6072
rect 35618 6060 35624 6072
rect 35676 6060 35682 6112
rect 1104 6010 38824 6032
rect 1104 5958 19606 6010
rect 19658 5958 19670 6010
rect 19722 5958 19734 6010
rect 19786 5958 19798 6010
rect 19850 5958 38824 6010
rect 1104 5936 38824 5958
rect 2774 5856 2780 5908
rect 2832 5896 2838 5908
rect 2832 5868 2877 5896
rect 2832 5856 2838 5868
rect 4062 5856 4068 5908
rect 4120 5896 4126 5908
rect 4249 5899 4307 5905
rect 4249 5896 4261 5899
rect 4120 5868 4261 5896
rect 4120 5856 4126 5868
rect 4249 5865 4261 5868
rect 4295 5865 4307 5899
rect 8570 5896 8576 5908
rect 4249 5859 4307 5865
rect 4356 5868 8576 5896
rect 3418 5720 3424 5772
rect 3476 5760 3482 5772
rect 4157 5763 4215 5769
rect 4157 5760 4169 5763
rect 3476 5732 4169 5760
rect 3476 5720 3482 5732
rect 4157 5729 4169 5732
rect 4203 5760 4215 5763
rect 4356 5760 4384 5868
rect 8570 5856 8576 5868
rect 8628 5856 8634 5908
rect 9769 5899 9827 5905
rect 9769 5865 9781 5899
rect 9815 5896 9827 5899
rect 11238 5896 11244 5908
rect 9815 5868 11244 5896
rect 9815 5865 9827 5868
rect 9769 5859 9827 5865
rect 11238 5856 11244 5868
rect 11296 5856 11302 5908
rect 13262 5896 13268 5908
rect 13175 5868 13268 5896
rect 13262 5856 13268 5868
rect 13320 5896 13326 5908
rect 13320 5868 15700 5896
rect 13320 5856 13326 5868
rect 6178 5788 6184 5840
rect 6236 5828 6242 5840
rect 6236 5800 6500 5828
rect 6236 5788 6242 5800
rect 5074 5760 5080 5772
rect 4203 5732 4384 5760
rect 5035 5732 5080 5760
rect 4203 5729 4215 5732
rect 4157 5723 4215 5729
rect 5074 5720 5080 5732
rect 5132 5720 5138 5772
rect 5258 5720 5264 5772
rect 5316 5760 5322 5772
rect 5905 5763 5963 5769
rect 5905 5760 5917 5763
rect 5316 5732 5917 5760
rect 5316 5720 5322 5732
rect 5905 5729 5917 5732
rect 5951 5760 5963 5763
rect 5994 5760 6000 5772
rect 5951 5732 6000 5760
rect 5951 5729 5963 5732
rect 5905 5723 5963 5729
rect 5994 5720 6000 5732
rect 6052 5720 6058 5772
rect 6472 5769 6500 5800
rect 6822 5788 6828 5840
rect 6880 5828 6886 5840
rect 6880 5800 7420 5828
rect 6880 5788 6886 5800
rect 7392 5769 7420 5800
rect 9490 5788 9496 5840
rect 9548 5828 9554 5840
rect 11333 5831 11391 5837
rect 9548 5800 10640 5828
rect 9548 5788 9554 5800
rect 6365 5763 6423 5769
rect 6365 5729 6377 5763
rect 6411 5729 6423 5763
rect 6365 5723 6423 5729
rect 6457 5763 6515 5769
rect 6457 5729 6469 5763
rect 6503 5729 6515 5763
rect 6457 5723 6515 5729
rect 7101 5763 7159 5769
rect 7101 5729 7113 5763
rect 7147 5760 7159 5763
rect 7377 5763 7435 5769
rect 7147 5732 7328 5760
rect 7147 5729 7159 5732
rect 7101 5723 7159 5729
rect 1394 5692 1400 5704
rect 1355 5664 1400 5692
rect 1394 5652 1400 5664
rect 1452 5652 1458 5704
rect 1670 5692 1676 5704
rect 1631 5664 1676 5692
rect 1670 5652 1676 5664
rect 1728 5652 1734 5704
rect 6380 5624 6408 5723
rect 6733 5695 6791 5701
rect 6733 5661 6745 5695
rect 6779 5692 6791 5695
rect 7190 5692 7196 5704
rect 6779 5664 7196 5692
rect 6779 5661 6791 5664
rect 6733 5655 6791 5661
rect 7190 5652 7196 5664
rect 7248 5652 7254 5704
rect 7300 5692 7328 5732
rect 7377 5729 7389 5763
rect 7423 5729 7435 5763
rect 8294 5760 8300 5772
rect 8255 5732 8300 5760
rect 7377 5723 7435 5729
rect 8294 5720 8300 5732
rect 8352 5720 8358 5772
rect 8389 5763 8447 5769
rect 8389 5729 8401 5763
rect 8435 5760 8447 5763
rect 8478 5760 8484 5772
rect 8435 5732 8484 5760
rect 8435 5729 8447 5732
rect 8389 5723 8447 5729
rect 8478 5720 8484 5732
rect 8536 5760 8542 5772
rect 9030 5760 9036 5772
rect 8536 5732 9036 5760
rect 8536 5720 8542 5732
rect 9030 5720 9036 5732
rect 9088 5720 9094 5772
rect 9674 5760 9680 5772
rect 9635 5732 9680 5760
rect 9674 5720 9680 5732
rect 9732 5720 9738 5772
rect 10612 5769 10640 5800
rect 11333 5797 11345 5831
rect 11379 5828 11391 5831
rect 12526 5828 12532 5840
rect 11379 5800 12532 5828
rect 11379 5797 11391 5800
rect 11333 5791 11391 5797
rect 12526 5788 12532 5800
rect 12584 5788 12590 5840
rect 10597 5763 10655 5769
rect 10597 5729 10609 5763
rect 10643 5729 10655 5763
rect 11054 5760 11060 5772
rect 11015 5732 11060 5760
rect 10597 5723 10655 5729
rect 11054 5720 11060 5732
rect 11112 5720 11118 5772
rect 11974 5760 11980 5772
rect 11935 5732 11980 5760
rect 11974 5720 11980 5732
rect 12032 5720 12038 5772
rect 12345 5763 12403 5769
rect 12345 5729 12357 5763
rect 12391 5760 12403 5763
rect 12618 5760 12624 5772
rect 12391 5732 12624 5760
rect 12391 5729 12403 5732
rect 12345 5723 12403 5729
rect 12618 5720 12624 5732
rect 12676 5720 12682 5772
rect 12805 5763 12863 5769
rect 12805 5729 12817 5763
rect 12851 5729 12863 5763
rect 12805 5723 12863 5729
rect 13173 5763 13231 5769
rect 13173 5729 13185 5763
rect 13219 5760 13231 5763
rect 13280 5760 13308 5856
rect 15562 5828 15568 5840
rect 13740 5800 15568 5828
rect 13740 5772 13768 5800
rect 15562 5788 15568 5800
rect 15620 5788 15626 5840
rect 15672 5828 15700 5868
rect 16666 5856 16672 5908
rect 16724 5896 16730 5908
rect 22186 5896 22192 5908
rect 16724 5868 22192 5896
rect 16724 5856 16730 5868
rect 22186 5856 22192 5868
rect 22244 5856 22250 5908
rect 27062 5896 27068 5908
rect 27023 5868 27068 5896
rect 27062 5856 27068 5868
rect 27120 5856 27126 5908
rect 27706 5856 27712 5908
rect 27764 5896 27770 5908
rect 36630 5896 36636 5908
rect 27764 5868 36636 5896
rect 27764 5856 27770 5868
rect 36630 5856 36636 5868
rect 36688 5856 36694 5908
rect 19978 5828 19984 5840
rect 15672 5800 19984 5828
rect 19978 5788 19984 5800
rect 20036 5788 20042 5840
rect 20714 5788 20720 5840
rect 20772 5828 20778 5840
rect 20772 5800 21588 5828
rect 20772 5788 20778 5800
rect 13722 5760 13728 5772
rect 13219 5732 13308 5760
rect 13635 5732 13728 5760
rect 13219 5729 13231 5732
rect 13173 5723 13231 5729
rect 10962 5692 10968 5704
rect 7300 5664 10968 5692
rect 10962 5652 10968 5664
rect 11020 5652 11026 5704
rect 12710 5692 12716 5704
rect 12671 5664 12716 5692
rect 12710 5652 12716 5664
rect 12768 5652 12774 5704
rect 12820 5692 12848 5723
rect 13722 5720 13728 5732
rect 13780 5720 13786 5772
rect 14461 5763 14519 5769
rect 14461 5729 14473 5763
rect 14507 5760 14519 5763
rect 15473 5763 15531 5769
rect 14507 5732 14780 5760
rect 14507 5729 14519 5732
rect 14461 5723 14519 5729
rect 12986 5692 12992 5704
rect 12820 5664 12992 5692
rect 12986 5652 12992 5664
rect 13044 5692 13050 5704
rect 14752 5692 14780 5732
rect 15473 5729 15485 5763
rect 15519 5760 15531 5763
rect 15654 5760 15660 5772
rect 15519 5732 15660 5760
rect 15519 5729 15531 5732
rect 15473 5723 15531 5729
rect 15654 5720 15660 5732
rect 15712 5720 15718 5772
rect 15838 5760 15844 5772
rect 15799 5732 15844 5760
rect 15838 5720 15844 5732
rect 15896 5720 15902 5772
rect 16301 5763 16359 5769
rect 16301 5729 16313 5763
rect 16347 5729 16359 5763
rect 16666 5760 16672 5772
rect 16627 5732 16672 5760
rect 16301 5723 16359 5729
rect 16316 5692 16344 5723
rect 16666 5720 16672 5732
rect 16724 5720 16730 5772
rect 17221 5763 17279 5769
rect 17221 5729 17233 5763
rect 17267 5760 17279 5763
rect 17678 5760 17684 5772
rect 17267 5732 17684 5760
rect 17267 5729 17279 5732
rect 17221 5723 17279 5729
rect 17678 5720 17684 5732
rect 17736 5760 17742 5772
rect 18506 5760 18512 5772
rect 17736 5732 18512 5760
rect 17736 5720 17742 5732
rect 18506 5720 18512 5732
rect 18564 5720 18570 5772
rect 19334 5760 19340 5772
rect 19295 5732 19340 5760
rect 19334 5720 19340 5732
rect 19392 5720 19398 5772
rect 19886 5760 19892 5772
rect 19847 5732 19892 5760
rect 19886 5720 19892 5732
rect 19944 5720 19950 5772
rect 20901 5763 20959 5769
rect 20901 5729 20913 5763
rect 20947 5729 20959 5763
rect 20901 5723 20959 5729
rect 16574 5692 16580 5704
rect 13044 5664 14688 5692
rect 14752 5664 16580 5692
rect 13044 5652 13050 5664
rect 7282 5624 7288 5636
rect 6380 5596 7288 5624
rect 7282 5584 7288 5596
rect 7340 5584 7346 5636
rect 8573 5627 8631 5633
rect 8573 5593 8585 5627
rect 8619 5624 8631 5627
rect 9490 5624 9496 5636
rect 8619 5596 9496 5624
rect 8619 5593 8631 5596
rect 8573 5587 8631 5593
rect 9490 5584 9496 5596
rect 9548 5584 9554 5636
rect 14660 5568 14688 5664
rect 16574 5652 16580 5664
rect 16632 5692 16638 5704
rect 17862 5692 17868 5704
rect 16632 5664 17868 5692
rect 16632 5652 16638 5664
rect 17862 5652 17868 5664
rect 17920 5652 17926 5704
rect 19061 5695 19119 5701
rect 19061 5661 19073 5695
rect 19107 5661 19119 5695
rect 19061 5655 19119 5661
rect 15010 5584 15016 5636
rect 15068 5624 15074 5636
rect 15381 5627 15439 5633
rect 15381 5624 15393 5627
rect 15068 5596 15393 5624
rect 15068 5584 15074 5596
rect 15381 5593 15393 5596
rect 15427 5593 15439 5627
rect 19076 5624 19104 5655
rect 19150 5652 19156 5704
rect 19208 5692 19214 5704
rect 19797 5695 19855 5701
rect 19797 5692 19809 5695
rect 19208 5664 19809 5692
rect 19208 5652 19214 5664
rect 19797 5661 19809 5664
rect 19843 5661 19855 5695
rect 19797 5655 19855 5661
rect 19886 5624 19892 5636
rect 19076 5596 19892 5624
rect 15381 5587 15439 5593
rect 19886 5584 19892 5596
rect 19944 5624 19950 5636
rect 20254 5624 20260 5636
rect 19944 5596 20260 5624
rect 19944 5584 19950 5596
rect 20254 5584 20260 5596
rect 20312 5584 20318 5636
rect 20916 5624 20944 5723
rect 20990 5720 20996 5772
rect 21048 5760 21054 5772
rect 21560 5769 21588 5800
rect 21726 5788 21732 5840
rect 21784 5828 21790 5840
rect 25314 5828 25320 5840
rect 21784 5800 24992 5828
rect 25275 5800 25320 5828
rect 21784 5788 21790 5800
rect 21545 5763 21603 5769
rect 21048 5732 21093 5760
rect 21048 5720 21054 5732
rect 21545 5729 21557 5763
rect 21591 5729 21603 5763
rect 22462 5760 22468 5772
rect 22423 5732 22468 5760
rect 21545 5723 21603 5729
rect 22462 5720 22468 5732
rect 22520 5720 22526 5772
rect 22646 5760 22652 5772
rect 22607 5732 22652 5760
rect 22646 5720 22652 5732
rect 22704 5720 22710 5772
rect 23106 5760 23112 5772
rect 23067 5732 23112 5760
rect 23106 5720 23112 5732
rect 23164 5720 23170 5772
rect 23842 5720 23848 5772
rect 23900 5760 23906 5772
rect 24118 5760 24124 5772
rect 23900 5732 24124 5760
rect 23900 5720 23906 5732
rect 24118 5720 24124 5732
rect 24176 5760 24182 5772
rect 24213 5763 24271 5769
rect 24213 5760 24225 5763
rect 24176 5732 24225 5760
rect 24176 5720 24182 5732
rect 24213 5729 24225 5732
rect 24259 5729 24271 5763
rect 24213 5723 24271 5729
rect 24302 5720 24308 5772
rect 24360 5760 24366 5772
rect 24670 5760 24676 5772
rect 24360 5732 24676 5760
rect 24360 5720 24366 5732
rect 24670 5720 24676 5732
rect 24728 5760 24734 5772
rect 24964 5769 24992 5800
rect 25314 5788 25320 5800
rect 25372 5788 25378 5840
rect 26786 5828 26792 5840
rect 26747 5800 26792 5828
rect 26786 5788 26792 5800
rect 26844 5788 26850 5840
rect 26878 5788 26884 5840
rect 26936 5828 26942 5840
rect 26973 5831 27031 5837
rect 26973 5828 26985 5831
rect 26936 5800 26985 5828
rect 26936 5788 26942 5800
rect 26973 5797 26985 5800
rect 27019 5797 27031 5831
rect 27154 5828 27160 5840
rect 27115 5800 27160 5828
rect 26973 5791 27031 5797
rect 27154 5788 27160 5800
rect 27212 5788 27218 5840
rect 27525 5831 27583 5837
rect 27525 5797 27537 5831
rect 27571 5828 27583 5831
rect 27798 5828 27804 5840
rect 27571 5800 27804 5828
rect 27571 5797 27583 5800
rect 27525 5791 27583 5797
rect 27798 5788 27804 5800
rect 27856 5788 27862 5840
rect 27982 5828 27988 5840
rect 27943 5800 27988 5828
rect 27982 5788 27988 5800
rect 28040 5788 28046 5840
rect 28534 5788 28540 5840
rect 28592 5828 28598 5840
rect 30190 5828 30196 5840
rect 28592 5800 30196 5828
rect 28592 5788 28598 5800
rect 30190 5788 30196 5800
rect 30248 5788 30254 5840
rect 32214 5828 32220 5840
rect 30300 5800 32220 5828
rect 24765 5763 24823 5769
rect 24765 5760 24777 5763
rect 24728 5732 24777 5760
rect 24728 5720 24734 5732
rect 24765 5729 24777 5732
rect 24811 5729 24823 5763
rect 24765 5723 24823 5729
rect 24949 5763 25007 5769
rect 24949 5729 24961 5763
rect 24995 5760 25007 5763
rect 27430 5760 27436 5772
rect 24995 5732 27436 5760
rect 24995 5729 25007 5732
rect 24949 5723 25007 5729
rect 27430 5720 27436 5732
rect 27488 5720 27494 5772
rect 28810 5760 28816 5772
rect 28771 5732 28816 5760
rect 28810 5720 28816 5732
rect 28868 5720 28874 5772
rect 28902 5720 28908 5772
rect 28960 5760 28966 5772
rect 30300 5769 30328 5800
rect 32214 5788 32220 5800
rect 32272 5788 32278 5840
rect 36078 5828 36084 5840
rect 36039 5800 36084 5828
rect 36078 5788 36084 5800
rect 36136 5788 36142 5840
rect 29457 5763 29515 5769
rect 29457 5760 29469 5763
rect 28960 5732 29469 5760
rect 28960 5720 28966 5732
rect 29457 5729 29469 5732
rect 29503 5729 29515 5763
rect 29457 5723 29515 5729
rect 30285 5763 30343 5769
rect 30285 5729 30297 5763
rect 30331 5729 30343 5763
rect 30285 5723 30343 5729
rect 31297 5763 31355 5769
rect 31297 5729 31309 5763
rect 31343 5729 31355 5763
rect 31297 5723 31355 5729
rect 22278 5692 22284 5704
rect 22239 5664 22284 5692
rect 22278 5652 22284 5664
rect 22336 5652 22342 5704
rect 24029 5695 24087 5701
rect 24029 5661 24041 5695
rect 24075 5661 24087 5695
rect 24029 5655 24087 5661
rect 28537 5695 28595 5701
rect 28537 5661 28549 5695
rect 28583 5661 28595 5695
rect 28537 5655 28595 5661
rect 28997 5695 29055 5701
rect 28997 5661 29009 5695
rect 29043 5692 29055 5695
rect 30006 5692 30012 5704
rect 29043 5664 29868 5692
rect 29967 5664 30012 5692
rect 29043 5661 29055 5664
rect 28997 5655 29055 5661
rect 21358 5624 21364 5636
rect 20916 5596 21364 5624
rect 21358 5584 21364 5596
rect 21416 5624 21422 5636
rect 24044 5624 24072 5655
rect 26234 5624 26240 5636
rect 21416 5596 26240 5624
rect 21416 5584 21422 5596
rect 26234 5584 26240 5596
rect 26292 5584 26298 5636
rect 28552 5624 28580 5655
rect 29840 5624 29868 5664
rect 30006 5652 30012 5664
rect 30064 5652 30070 5704
rect 30466 5652 30472 5704
rect 30524 5692 30530 5704
rect 31202 5692 31208 5704
rect 30524 5664 31208 5692
rect 30524 5652 30530 5664
rect 31202 5652 31208 5664
rect 31260 5652 31266 5704
rect 31312 5692 31340 5723
rect 32766 5720 32772 5772
rect 32824 5760 32830 5772
rect 34698 5760 34704 5772
rect 32824 5732 34560 5760
rect 34659 5732 34704 5760
rect 32824 5720 32830 5732
rect 32030 5692 32036 5704
rect 31312 5664 32036 5692
rect 32030 5652 32036 5664
rect 32088 5652 32094 5704
rect 32122 5652 32128 5704
rect 32180 5692 32186 5704
rect 32398 5692 32404 5704
rect 32180 5664 32225 5692
rect 32359 5664 32404 5692
rect 32180 5652 32186 5664
rect 32398 5652 32404 5664
rect 32456 5652 32462 5704
rect 32490 5652 32496 5704
rect 32548 5692 32554 5704
rect 33505 5695 33563 5701
rect 33505 5692 33517 5695
rect 32548 5664 33517 5692
rect 32548 5652 32554 5664
rect 33505 5661 33517 5664
rect 33551 5661 33563 5695
rect 33505 5655 33563 5661
rect 34425 5695 34483 5701
rect 34425 5661 34437 5695
rect 34471 5661 34483 5695
rect 34532 5692 34560 5732
rect 34698 5720 34704 5732
rect 34756 5720 34762 5772
rect 35802 5720 35808 5772
rect 35860 5760 35866 5772
rect 36541 5763 36599 5769
rect 36541 5760 36553 5763
rect 35860 5732 36553 5760
rect 35860 5720 35866 5732
rect 36541 5729 36553 5732
rect 36587 5729 36599 5763
rect 36541 5723 36599 5729
rect 36722 5720 36728 5772
rect 36780 5760 36786 5772
rect 37737 5763 37795 5769
rect 37737 5760 37749 5763
rect 36780 5732 37749 5760
rect 36780 5720 36786 5732
rect 37737 5729 37749 5732
rect 37783 5729 37795 5763
rect 37737 5723 37795 5729
rect 34532 5664 36768 5692
rect 34425 5655 34483 5661
rect 31938 5624 31944 5636
rect 28552 5596 29040 5624
rect 29840 5596 31944 5624
rect 29012 5568 29040 5596
rect 31938 5584 31944 5596
rect 31996 5584 32002 5636
rect 5169 5559 5227 5565
rect 5169 5525 5181 5559
rect 5215 5556 5227 5559
rect 6638 5556 6644 5568
rect 5215 5528 6644 5556
rect 5215 5525 5227 5528
rect 5169 5519 5227 5525
rect 6638 5516 6644 5528
rect 6696 5516 6702 5568
rect 7466 5516 7472 5568
rect 7524 5556 7530 5568
rect 8113 5559 8171 5565
rect 8113 5556 8125 5559
rect 7524 5528 8125 5556
rect 7524 5516 7530 5528
rect 8113 5525 8125 5528
rect 8159 5525 8171 5559
rect 8113 5519 8171 5525
rect 11514 5516 11520 5568
rect 11572 5556 11578 5568
rect 13722 5556 13728 5568
rect 11572 5528 13728 5556
rect 11572 5516 11578 5528
rect 13722 5516 13728 5528
rect 13780 5516 13786 5568
rect 14642 5556 14648 5568
rect 14603 5528 14648 5556
rect 14642 5516 14648 5528
rect 14700 5516 14706 5568
rect 15562 5516 15568 5568
rect 15620 5556 15626 5568
rect 17865 5559 17923 5565
rect 17865 5556 17877 5559
rect 15620 5528 17877 5556
rect 15620 5516 15626 5528
rect 17865 5525 17877 5528
rect 17911 5525 17923 5559
rect 21634 5556 21640 5568
rect 21595 5528 21640 5556
rect 17865 5519 17923 5525
rect 21634 5516 21640 5528
rect 21692 5516 21698 5568
rect 28994 5516 29000 5568
rect 29052 5516 29058 5568
rect 30926 5516 30932 5568
rect 30984 5556 30990 5568
rect 31481 5559 31539 5565
rect 31481 5556 31493 5559
rect 30984 5528 31493 5556
rect 30984 5516 30990 5528
rect 31481 5525 31493 5528
rect 31527 5525 31539 5559
rect 34440 5556 34468 5655
rect 36740 5633 36768 5664
rect 36725 5627 36783 5633
rect 36725 5593 36737 5627
rect 36771 5593 36783 5627
rect 37918 5624 37924 5636
rect 37879 5596 37924 5624
rect 36725 5587 36783 5593
rect 37918 5584 37924 5596
rect 37976 5584 37982 5636
rect 36078 5556 36084 5568
rect 34440 5528 36084 5556
rect 31481 5519 31539 5525
rect 36078 5516 36084 5528
rect 36136 5516 36142 5568
rect 1104 5466 38824 5488
rect 1104 5414 4246 5466
rect 4298 5414 4310 5466
rect 4362 5414 4374 5466
rect 4426 5414 4438 5466
rect 4490 5414 34966 5466
rect 35018 5414 35030 5466
rect 35082 5414 35094 5466
rect 35146 5414 35158 5466
rect 35210 5414 38824 5466
rect 1104 5392 38824 5414
rect 1670 5312 1676 5364
rect 1728 5352 1734 5364
rect 2225 5355 2283 5361
rect 2225 5352 2237 5355
rect 1728 5324 2237 5352
rect 1728 5312 1734 5324
rect 2225 5321 2237 5324
rect 2271 5321 2283 5355
rect 16666 5352 16672 5364
rect 2225 5315 2283 5321
rect 4816 5324 16672 5352
rect 3234 5176 3240 5228
rect 3292 5216 3298 5228
rect 3421 5219 3479 5225
rect 3421 5216 3433 5219
rect 3292 5188 3433 5216
rect 3292 5176 3298 5188
rect 3421 5185 3433 5188
rect 3467 5185 3479 5219
rect 3421 5179 3479 5185
rect 1949 5151 2007 5157
rect 1949 5117 1961 5151
rect 1995 5117 2007 5151
rect 1949 5111 2007 5117
rect 1964 5012 1992 5111
rect 2038 5108 2044 5160
rect 2096 5148 2102 5160
rect 3513 5151 3571 5157
rect 2096 5120 2141 5148
rect 2096 5108 2102 5120
rect 3513 5117 3525 5151
rect 3559 5117 3571 5151
rect 3786 5148 3792 5160
rect 3747 5120 3792 5148
rect 3513 5111 3571 5117
rect 2958 5012 2964 5024
rect 1964 4984 2964 5012
rect 2958 4972 2964 4984
rect 3016 5012 3022 5024
rect 3418 5012 3424 5024
rect 3016 4984 3424 5012
rect 3016 4972 3022 4984
rect 3418 4972 3424 4984
rect 3476 4972 3482 5024
rect 3528 5012 3556 5111
rect 3786 5108 3792 5120
rect 3844 5108 3850 5160
rect 4341 5151 4399 5157
rect 4341 5117 4353 5151
rect 4387 5148 4399 5151
rect 4614 5148 4620 5160
rect 4387 5120 4620 5148
rect 4387 5117 4399 5120
rect 4341 5111 4399 5117
rect 4614 5108 4620 5120
rect 4672 5108 4678 5160
rect 4709 5151 4767 5157
rect 4709 5117 4721 5151
rect 4755 5148 4767 5151
rect 4816 5148 4844 5324
rect 16666 5312 16672 5324
rect 16724 5312 16730 5364
rect 20254 5312 20260 5364
rect 20312 5352 20318 5364
rect 21361 5355 21419 5361
rect 21361 5352 21373 5355
rect 20312 5324 21373 5352
rect 20312 5312 20318 5324
rect 21361 5321 21373 5324
rect 21407 5321 21419 5355
rect 21361 5315 21419 5321
rect 23106 5312 23112 5364
rect 23164 5352 23170 5364
rect 23845 5355 23903 5361
rect 23845 5352 23857 5355
rect 23164 5324 23857 5352
rect 23164 5312 23170 5324
rect 23845 5321 23857 5324
rect 23891 5321 23903 5355
rect 23845 5315 23903 5321
rect 26878 5312 26884 5364
rect 26936 5352 26942 5364
rect 28445 5355 28503 5361
rect 28445 5352 28457 5355
rect 26936 5324 28457 5352
rect 26936 5312 26942 5324
rect 28445 5321 28457 5324
rect 28491 5321 28503 5355
rect 28445 5315 28503 5321
rect 30926 5312 30932 5364
rect 30984 5352 30990 5364
rect 32858 5352 32864 5364
rect 30984 5324 32864 5352
rect 30984 5312 30990 5324
rect 32858 5312 32864 5324
rect 32916 5312 32922 5364
rect 33502 5312 33508 5364
rect 33560 5352 33566 5364
rect 33597 5355 33655 5361
rect 33597 5352 33609 5355
rect 33560 5324 33609 5352
rect 33560 5312 33566 5324
rect 33597 5321 33609 5324
rect 33643 5321 33655 5355
rect 33597 5315 33655 5321
rect 37366 5312 37372 5364
rect 37424 5352 37430 5364
rect 37737 5355 37795 5361
rect 37737 5352 37749 5355
rect 37424 5324 37749 5352
rect 37424 5312 37430 5324
rect 37737 5321 37749 5324
rect 37783 5321 37795 5355
rect 37737 5315 37795 5321
rect 6181 5287 6239 5293
rect 6181 5253 6193 5287
rect 6227 5253 6239 5287
rect 6181 5247 6239 5253
rect 6917 5287 6975 5293
rect 6917 5253 6929 5287
rect 6963 5284 6975 5287
rect 7282 5284 7288 5296
rect 6963 5256 7288 5284
rect 6963 5253 6975 5256
rect 6917 5247 6975 5253
rect 6196 5216 6224 5247
rect 7282 5244 7288 5256
rect 7340 5244 7346 5296
rect 9033 5287 9091 5293
rect 9033 5253 9045 5287
rect 9079 5284 9091 5287
rect 12434 5284 12440 5296
rect 9079 5256 12440 5284
rect 9079 5253 9091 5256
rect 9033 5247 9091 5253
rect 12434 5244 12440 5256
rect 12492 5244 12498 5296
rect 12805 5287 12863 5293
rect 12805 5253 12817 5287
rect 12851 5284 12863 5287
rect 13081 5287 13139 5293
rect 13081 5284 13093 5287
rect 12851 5256 13093 5284
rect 12851 5253 12863 5256
rect 12805 5247 12863 5253
rect 13081 5253 13093 5256
rect 13127 5284 13139 5287
rect 13906 5284 13912 5296
rect 13127 5256 13676 5284
rect 13867 5256 13912 5284
rect 13127 5253 13139 5256
rect 13081 5247 13139 5253
rect 7374 5216 7380 5228
rect 6196 5188 7380 5216
rect 7374 5176 7380 5188
rect 7432 5176 7438 5228
rect 7745 5219 7803 5225
rect 7745 5185 7757 5219
rect 7791 5216 7803 5219
rect 9677 5219 9735 5225
rect 9677 5216 9689 5219
rect 7791 5188 9689 5216
rect 7791 5185 7803 5188
rect 7745 5179 7803 5185
rect 9677 5185 9689 5188
rect 9723 5185 9735 5219
rect 10870 5216 10876 5228
rect 9677 5179 9735 5185
rect 10612 5188 10876 5216
rect 4755 5120 4844 5148
rect 5261 5151 5319 5157
rect 4755 5117 4767 5120
rect 4709 5111 4767 5117
rect 5261 5117 5273 5151
rect 5307 5117 5319 5151
rect 5261 5111 5319 5117
rect 5276 5080 5304 5111
rect 5810 5108 5816 5160
rect 5868 5148 5874 5160
rect 5997 5151 6055 5157
rect 5997 5148 6009 5151
rect 5868 5120 6009 5148
rect 5868 5108 5874 5120
rect 5997 5117 6009 5120
rect 6043 5117 6055 5151
rect 5997 5111 6055 5117
rect 6825 5151 6883 5157
rect 6825 5117 6837 5151
rect 6871 5148 6883 5151
rect 7006 5148 7012 5160
rect 6871 5120 7012 5148
rect 6871 5117 6883 5120
rect 6825 5111 6883 5117
rect 7006 5108 7012 5120
rect 7064 5108 7070 5160
rect 7466 5148 7472 5160
rect 7427 5120 7472 5148
rect 7466 5108 7472 5120
rect 7524 5108 7530 5160
rect 9769 5151 9827 5157
rect 9769 5117 9781 5151
rect 9815 5117 9827 5151
rect 10226 5148 10232 5160
rect 10187 5120 10232 5148
rect 9769 5111 9827 5117
rect 5276 5052 6868 5080
rect 6840 5024 6868 5052
rect 5258 5012 5264 5024
rect 3528 4984 5264 5012
rect 5258 4972 5264 4984
rect 5316 4972 5322 5024
rect 6822 4972 6828 5024
rect 6880 4972 6886 5024
rect 9784 5012 9812 5111
rect 10226 5108 10232 5120
rect 10284 5108 10290 5160
rect 10612 5157 10640 5188
rect 10870 5176 10876 5188
rect 10928 5216 10934 5228
rect 12986 5216 12992 5228
rect 10928 5188 12992 5216
rect 10928 5176 10934 5188
rect 12986 5176 12992 5188
rect 13044 5176 13050 5228
rect 10597 5151 10655 5157
rect 10597 5117 10609 5151
rect 10643 5117 10655 5151
rect 10962 5148 10968 5160
rect 10923 5120 10968 5148
rect 10597 5111 10655 5117
rect 10962 5108 10968 5120
rect 11020 5108 11026 5160
rect 11514 5148 11520 5160
rect 11475 5120 11520 5148
rect 11514 5108 11520 5120
rect 11572 5108 11578 5160
rect 13648 5157 13676 5256
rect 13906 5244 13912 5256
rect 13964 5244 13970 5296
rect 22005 5287 22063 5293
rect 22005 5284 22017 5287
rect 19352 5256 22017 5284
rect 19352 5228 19380 5256
rect 22005 5253 22017 5256
rect 22051 5253 22063 5287
rect 22005 5247 22063 5253
rect 22646 5244 22652 5296
rect 22704 5244 22710 5296
rect 31110 5244 31116 5296
rect 31168 5284 31174 5296
rect 34422 5284 34428 5296
rect 31168 5256 34428 5284
rect 31168 5244 31174 5256
rect 13722 5176 13728 5228
rect 13780 5216 13786 5228
rect 19334 5216 19340 5228
rect 13780 5188 19340 5216
rect 13780 5176 13786 5188
rect 19334 5176 19340 5188
rect 19392 5176 19398 5228
rect 20806 5216 20812 5228
rect 20456 5188 20812 5216
rect 12897 5151 12955 5157
rect 12897 5117 12909 5151
rect 12943 5117 12955 5151
rect 12897 5111 12955 5117
rect 13633 5151 13691 5157
rect 13633 5117 13645 5151
rect 13679 5117 13691 5151
rect 14274 5148 14280 5160
rect 14235 5120 14280 5148
rect 13633 5111 13691 5117
rect 12912 5080 12940 5111
rect 14274 5108 14280 5120
rect 14332 5108 14338 5160
rect 14642 5148 14648 5160
rect 14603 5120 14648 5148
rect 14642 5108 14648 5120
rect 14700 5108 14706 5160
rect 15013 5151 15071 5157
rect 15013 5117 15025 5151
rect 15059 5148 15071 5151
rect 15194 5148 15200 5160
rect 15059 5120 15200 5148
rect 15059 5117 15071 5120
rect 15013 5111 15071 5117
rect 15194 5108 15200 5120
rect 15252 5108 15258 5160
rect 15562 5148 15568 5160
rect 15523 5120 15568 5148
rect 15562 5108 15568 5120
rect 15620 5108 15626 5160
rect 16482 5148 16488 5160
rect 16443 5120 16488 5148
rect 16482 5108 16488 5120
rect 16540 5108 16546 5160
rect 16942 5148 16948 5160
rect 16903 5120 16948 5148
rect 16942 5108 16948 5120
rect 17000 5108 17006 5160
rect 18049 5151 18107 5157
rect 18049 5148 18061 5151
rect 17052 5120 18061 5148
rect 15930 5080 15936 5092
rect 12912 5052 15936 5080
rect 15930 5040 15936 5052
rect 15988 5040 15994 5092
rect 16500 5080 16528 5108
rect 17052 5080 17080 5120
rect 18049 5117 18061 5120
rect 18095 5117 18107 5151
rect 18598 5148 18604 5160
rect 18559 5120 18604 5148
rect 18049 5111 18107 5117
rect 18598 5108 18604 5120
rect 18656 5108 18662 5160
rect 19426 5108 19432 5160
rect 19484 5148 19490 5160
rect 19521 5151 19579 5157
rect 19521 5148 19533 5151
rect 19484 5120 19533 5148
rect 19484 5108 19490 5120
rect 19521 5117 19533 5120
rect 19567 5117 19579 5151
rect 19521 5111 19579 5117
rect 20073 5151 20131 5157
rect 20073 5117 20085 5151
rect 20119 5148 20131 5151
rect 20456 5148 20484 5188
rect 20806 5176 20812 5188
rect 20864 5216 20870 5228
rect 21266 5216 21272 5228
rect 20864 5188 21272 5216
rect 20864 5176 20870 5188
rect 21266 5176 21272 5188
rect 21324 5176 21330 5228
rect 22664 5216 22692 5244
rect 22572 5188 22692 5216
rect 20119 5120 20484 5148
rect 20533 5151 20591 5157
rect 20119 5117 20131 5120
rect 20073 5111 20131 5117
rect 20533 5117 20545 5151
rect 20579 5148 20591 5151
rect 21177 5151 21235 5157
rect 21177 5148 21189 5151
rect 20579 5120 21189 5148
rect 20579 5117 20591 5120
rect 20533 5111 20591 5117
rect 21177 5117 21189 5120
rect 21223 5148 21235 5151
rect 21634 5148 21640 5160
rect 21223 5120 21640 5148
rect 21223 5117 21235 5120
rect 21177 5111 21235 5117
rect 21634 5108 21640 5120
rect 21692 5108 21698 5160
rect 22572 5157 22600 5188
rect 24854 5176 24860 5228
rect 24912 5216 24918 5228
rect 24949 5219 25007 5225
rect 24949 5216 24961 5219
rect 24912 5188 24961 5216
rect 24912 5176 24918 5188
rect 24949 5185 24961 5188
rect 24995 5216 25007 5219
rect 25130 5216 25136 5228
rect 24995 5188 25136 5216
rect 24995 5185 25007 5188
rect 24949 5179 25007 5185
rect 25130 5176 25136 5188
rect 25188 5216 25194 5228
rect 26786 5216 26792 5228
rect 25188 5188 26792 5216
rect 25188 5176 25194 5188
rect 26786 5176 26792 5188
rect 26844 5216 26850 5228
rect 27065 5219 27123 5225
rect 27065 5216 27077 5219
rect 26844 5188 27077 5216
rect 26844 5176 26850 5188
rect 27065 5185 27077 5188
rect 27111 5216 27123 5219
rect 29178 5216 29184 5228
rect 27111 5188 29184 5216
rect 27111 5185 27123 5188
rect 27065 5179 27123 5185
rect 29178 5176 29184 5188
rect 29236 5176 29242 5228
rect 29825 5219 29883 5225
rect 29825 5185 29837 5219
rect 29871 5216 29883 5219
rect 30006 5216 30012 5228
rect 29871 5188 30012 5216
rect 29871 5185 29883 5188
rect 29825 5179 29883 5185
rect 30006 5176 30012 5188
rect 30064 5176 30070 5228
rect 32508 5225 32536 5256
rect 34422 5244 34428 5256
rect 34480 5244 34486 5296
rect 32493 5219 32551 5225
rect 30116 5188 32444 5216
rect 22189 5151 22247 5157
rect 22189 5117 22201 5151
rect 22235 5117 22247 5151
rect 22189 5111 22247 5117
rect 22557 5151 22615 5157
rect 22557 5117 22569 5151
rect 22603 5117 22615 5151
rect 22922 5148 22928 5160
rect 22883 5120 22928 5148
rect 22557 5111 22615 5117
rect 16500 5052 17080 5080
rect 17221 5083 17279 5089
rect 17221 5049 17233 5083
rect 17267 5080 17279 5083
rect 18322 5080 18328 5092
rect 17267 5052 18328 5080
rect 17267 5049 17279 5052
rect 17221 5043 17279 5049
rect 18322 5040 18328 5052
rect 18380 5040 18386 5092
rect 18785 5083 18843 5089
rect 18785 5049 18797 5083
rect 18831 5080 18843 5083
rect 20622 5080 20628 5092
rect 18831 5052 20628 5080
rect 18831 5049 18843 5052
rect 18785 5043 18843 5049
rect 20622 5040 20628 5052
rect 20680 5040 20686 5092
rect 20714 5040 20720 5092
rect 20772 5080 20778 5092
rect 20772 5052 20817 5080
rect 20772 5040 20778 5052
rect 10226 5012 10232 5024
rect 9784 4984 10232 5012
rect 10226 4972 10232 4984
rect 10284 5012 10290 5024
rect 11974 5012 11980 5024
rect 10284 4984 11980 5012
rect 10284 4972 10290 4984
rect 11974 4972 11980 4984
rect 12032 5012 12038 5024
rect 12805 5015 12863 5021
rect 12805 5012 12817 5015
rect 12032 4984 12817 5012
rect 12032 4972 12038 4984
rect 12805 4981 12817 4984
rect 12851 4981 12863 5015
rect 12805 4975 12863 4981
rect 17954 4972 17960 5024
rect 18012 5012 18018 5024
rect 20898 5012 20904 5024
rect 18012 4984 20904 5012
rect 18012 4972 18018 4984
rect 20898 4972 20904 4984
rect 20956 4972 20962 5024
rect 22204 5012 22232 5111
rect 22922 5108 22928 5120
rect 22980 5108 22986 5160
rect 23658 5148 23664 5160
rect 23619 5120 23664 5148
rect 23658 5108 23664 5120
rect 23716 5108 23722 5160
rect 25222 5148 25228 5160
rect 25183 5120 25228 5148
rect 25222 5108 25228 5120
rect 25280 5108 25286 5160
rect 27341 5151 27399 5157
rect 27341 5117 27353 5151
rect 27387 5148 27399 5151
rect 30116 5148 30144 5188
rect 27387 5120 30144 5148
rect 30377 5151 30435 5157
rect 27387 5117 27399 5120
rect 27341 5111 27399 5117
rect 30377 5117 30389 5151
rect 30423 5117 30435 5151
rect 30650 5148 30656 5160
rect 30611 5120 30656 5148
rect 30377 5111 30435 5117
rect 26605 5083 26663 5089
rect 26605 5049 26617 5083
rect 26651 5080 26663 5083
rect 27154 5080 27160 5092
rect 26651 5052 27160 5080
rect 26651 5049 26663 5052
rect 26605 5043 26663 5049
rect 27154 5040 27160 5052
rect 27212 5040 27218 5092
rect 30392 5080 30420 5111
rect 30650 5108 30656 5120
rect 30708 5108 30714 5160
rect 30834 5148 30840 5160
rect 30795 5120 30840 5148
rect 30834 5108 30840 5120
rect 30892 5148 30898 5160
rect 31754 5148 31760 5160
rect 30892 5120 31760 5148
rect 30892 5108 30898 5120
rect 31754 5108 31760 5120
rect 31812 5108 31818 5160
rect 32416 5148 32444 5188
rect 32493 5185 32505 5219
rect 32539 5185 32551 5219
rect 34885 5219 34943 5225
rect 34885 5216 34897 5219
rect 32493 5179 32551 5185
rect 32692 5188 34897 5216
rect 32692 5148 32720 5188
rect 34885 5185 34897 5188
rect 34931 5185 34943 5219
rect 34885 5179 34943 5185
rect 35802 5176 35808 5228
rect 35860 5216 35866 5228
rect 35897 5219 35955 5225
rect 35897 5216 35909 5219
rect 35860 5188 35909 5216
rect 35860 5176 35866 5188
rect 35897 5185 35909 5188
rect 35943 5185 35955 5219
rect 36630 5216 36636 5228
rect 36591 5188 36636 5216
rect 35897 5179 35955 5185
rect 36630 5176 36636 5188
rect 36688 5176 36694 5228
rect 32416 5120 32720 5148
rect 32769 5151 32827 5157
rect 32769 5117 32781 5151
rect 32815 5148 32827 5151
rect 32858 5148 32864 5160
rect 32815 5120 32864 5148
rect 32815 5117 32827 5120
rect 32769 5111 32827 5117
rect 32858 5108 32864 5120
rect 32916 5108 32922 5160
rect 32953 5151 33011 5157
rect 32953 5117 32965 5151
rect 32999 5117 33011 5151
rect 32953 5111 33011 5117
rect 31110 5080 31116 5092
rect 30392 5052 31116 5080
rect 31110 5040 31116 5052
rect 31168 5040 31174 5092
rect 31941 5083 31999 5089
rect 31941 5049 31953 5083
rect 31987 5080 31999 5083
rect 32674 5080 32680 5092
rect 31987 5052 32680 5080
rect 31987 5049 31999 5052
rect 31941 5043 31999 5049
rect 32674 5040 32680 5052
rect 32732 5040 32738 5092
rect 32968 5024 32996 5111
rect 33226 5108 33232 5160
rect 33284 5148 33290 5160
rect 33413 5151 33471 5157
rect 33413 5148 33425 5151
rect 33284 5120 33425 5148
rect 33284 5108 33290 5120
rect 33413 5117 33425 5120
rect 33459 5117 33471 5151
rect 33413 5111 33471 5117
rect 33594 5108 33600 5160
rect 33652 5148 33658 5160
rect 35437 5151 35495 5157
rect 35437 5148 35449 5151
rect 33652 5120 35449 5148
rect 33652 5108 33658 5120
rect 35437 5117 35449 5120
rect 35483 5117 35495 5151
rect 35710 5148 35716 5160
rect 35671 5120 35716 5148
rect 35437 5111 35495 5117
rect 35710 5108 35716 5120
rect 35768 5108 35774 5160
rect 36078 5108 36084 5160
rect 36136 5148 36142 5160
rect 36357 5151 36415 5157
rect 36357 5148 36369 5151
rect 36136 5120 36369 5148
rect 36136 5108 36142 5120
rect 36357 5117 36369 5120
rect 36403 5117 36415 5151
rect 36357 5111 36415 5117
rect 28166 5012 28172 5024
rect 22204 4984 28172 5012
rect 28166 4972 28172 4984
rect 28224 4972 28230 5024
rect 31754 4972 31760 5024
rect 31812 5012 31818 5024
rect 32950 5012 32956 5024
rect 31812 4984 32956 5012
rect 31812 4972 31818 4984
rect 32950 4972 32956 4984
rect 33008 4972 33014 5024
rect 1104 4922 38824 4944
rect 1104 4870 19606 4922
rect 19658 4870 19670 4922
rect 19722 4870 19734 4922
rect 19786 4870 19798 4922
rect 19850 4870 38824 4922
rect 1104 4848 38824 4870
rect 2038 4768 2044 4820
rect 2096 4808 2102 4820
rect 2777 4811 2835 4817
rect 2777 4808 2789 4811
rect 2096 4780 2789 4808
rect 2096 4768 2102 4780
rect 2777 4777 2789 4780
rect 2823 4777 2835 4811
rect 2777 4771 2835 4777
rect 6472 4780 11192 4808
rect 6362 4740 6368 4752
rect 4448 4712 6368 4740
rect 4448 4681 4476 4712
rect 6362 4700 6368 4712
rect 6420 4700 6426 4752
rect 4433 4675 4491 4681
rect 4433 4641 4445 4675
rect 4479 4641 4491 4675
rect 5258 4672 5264 4684
rect 5219 4644 5264 4672
rect 4433 4635 4491 4641
rect 5258 4632 5264 4644
rect 5316 4632 5322 4684
rect 5537 4675 5595 4681
rect 5537 4641 5549 4675
rect 5583 4641 5595 4675
rect 5537 4635 5595 4641
rect 6089 4675 6147 4681
rect 6089 4641 6101 4675
rect 6135 4672 6147 4675
rect 6178 4672 6184 4684
rect 6135 4644 6184 4672
rect 6135 4641 6147 4644
rect 6089 4635 6147 4641
rect 1394 4604 1400 4616
rect 1355 4576 1400 4604
rect 1394 4564 1400 4576
rect 1452 4564 1458 4616
rect 1670 4604 1676 4616
rect 1631 4576 1676 4604
rect 1670 4564 1676 4576
rect 1728 4564 1734 4616
rect 5442 4604 5448 4616
rect 5403 4576 5448 4604
rect 5442 4564 5448 4576
rect 5500 4564 5506 4616
rect 5552 4536 5580 4635
rect 6178 4632 6184 4644
rect 6236 4632 6242 4684
rect 6472 4681 6500 4780
rect 9125 4743 9183 4749
rect 9125 4709 9137 4743
rect 9171 4740 9183 4743
rect 9766 4740 9772 4752
rect 9171 4712 9772 4740
rect 9171 4709 9183 4712
rect 9125 4703 9183 4709
rect 9766 4700 9772 4712
rect 9824 4700 9830 4752
rect 6457 4675 6515 4681
rect 6457 4641 6469 4675
rect 6503 4641 6515 4675
rect 6822 4672 6828 4684
rect 6783 4644 6828 4672
rect 6457 4635 6515 4641
rect 6822 4632 6828 4644
rect 6880 4632 6886 4684
rect 7466 4672 7472 4684
rect 7379 4644 7472 4672
rect 7466 4632 7472 4644
rect 7524 4672 7530 4684
rect 7834 4672 7840 4684
rect 7524 4644 7840 4672
rect 7524 4632 7530 4644
rect 7834 4632 7840 4644
rect 7892 4632 7898 4684
rect 10226 4672 10232 4684
rect 10187 4644 10232 4672
rect 10226 4632 10232 4644
rect 10284 4632 10290 4684
rect 10686 4672 10692 4684
rect 10647 4644 10692 4672
rect 10686 4632 10692 4644
rect 10744 4632 10750 4684
rect 10870 4672 10876 4684
rect 10831 4644 10876 4672
rect 10870 4632 10876 4644
rect 10928 4632 10934 4684
rect 11164 4672 11192 4780
rect 12066 4768 12072 4820
rect 12124 4808 12130 4820
rect 12124 4780 14228 4808
rect 12124 4768 12130 4780
rect 14200 4740 14228 4780
rect 14274 4768 14280 4820
rect 14332 4808 14338 4820
rect 14645 4811 14703 4817
rect 14645 4808 14657 4811
rect 14332 4780 14657 4808
rect 14332 4768 14338 4780
rect 14645 4777 14657 4780
rect 14691 4777 14703 4811
rect 14645 4771 14703 4777
rect 18598 4768 18604 4820
rect 18656 4808 18662 4820
rect 20993 4811 21051 4817
rect 20993 4808 21005 4811
rect 18656 4780 21005 4808
rect 18656 4768 18662 4780
rect 20993 4777 21005 4780
rect 21039 4777 21051 4811
rect 20993 4771 21051 4777
rect 22738 4768 22744 4820
rect 22796 4808 22802 4820
rect 23385 4811 23443 4817
rect 23385 4808 23397 4811
rect 22796 4780 23397 4808
rect 22796 4768 22802 4780
rect 23385 4777 23397 4780
rect 23431 4777 23443 4811
rect 30926 4808 30932 4820
rect 23385 4771 23443 4777
rect 24228 4780 30932 4808
rect 22646 4740 22652 4752
rect 14200 4712 22140 4740
rect 11238 4672 11244 4684
rect 11151 4644 11244 4672
rect 11238 4632 11244 4644
rect 11296 4632 11302 4684
rect 11514 4632 11520 4684
rect 11572 4672 11578 4684
rect 11701 4675 11759 4681
rect 11701 4672 11713 4675
rect 11572 4644 11713 4672
rect 11572 4632 11578 4644
rect 11701 4641 11713 4644
rect 11747 4641 11759 4675
rect 12710 4672 12716 4684
rect 12671 4644 12716 4672
rect 11701 4635 11759 4641
rect 12710 4632 12716 4644
rect 12768 4632 12774 4684
rect 14550 4672 14556 4684
rect 14511 4644 14556 4672
rect 14550 4632 14556 4644
rect 14608 4632 14614 4684
rect 15746 4672 15752 4684
rect 15707 4644 15752 4672
rect 15746 4632 15752 4644
rect 15804 4632 15810 4684
rect 15930 4632 15936 4684
rect 15988 4672 15994 4684
rect 16853 4675 16911 4681
rect 16853 4672 16865 4675
rect 15988 4644 16865 4672
rect 15988 4632 15994 4644
rect 16853 4641 16865 4644
rect 16899 4641 16911 4675
rect 16853 4635 16911 4641
rect 16942 4632 16948 4684
rect 17000 4632 17006 4684
rect 17497 4675 17555 4681
rect 17497 4641 17509 4675
rect 17543 4641 17555 4675
rect 17862 4672 17868 4684
rect 17823 4644 17868 4672
rect 17497 4635 17555 4641
rect 7745 4607 7803 4613
rect 7745 4573 7757 4607
rect 7791 4604 7803 4607
rect 9490 4604 9496 4616
rect 7791 4576 9496 4604
rect 7791 4573 7803 4576
rect 7745 4567 7803 4573
rect 9490 4564 9496 4576
rect 9548 4564 9554 4616
rect 12437 4607 12495 4613
rect 12437 4573 12449 4607
rect 12483 4604 12495 4607
rect 14734 4604 14740 4616
rect 12483 4576 14740 4604
rect 12483 4573 12495 4576
rect 12437 4567 12495 4573
rect 14734 4564 14740 4576
rect 14792 4564 14798 4616
rect 15657 4607 15715 4613
rect 15657 4573 15669 4607
rect 15703 4604 15715 4607
rect 16960 4604 16988 4632
rect 15703 4576 16988 4604
rect 17512 4604 17540 4635
rect 17862 4632 17868 4644
rect 17920 4632 17926 4684
rect 18230 4672 18236 4684
rect 18191 4644 18236 4672
rect 18230 4632 18236 4644
rect 18288 4632 18294 4684
rect 18506 4672 18512 4684
rect 18467 4644 18512 4672
rect 18506 4632 18512 4644
rect 18564 4632 18570 4684
rect 19797 4675 19855 4681
rect 19797 4641 19809 4675
rect 19843 4641 19855 4675
rect 19797 4635 19855 4641
rect 20165 4675 20223 4681
rect 20165 4641 20177 4675
rect 20211 4672 20223 4675
rect 20714 4672 20720 4684
rect 20211 4644 20720 4672
rect 20211 4641 20223 4644
rect 20165 4635 20223 4641
rect 18598 4604 18604 4616
rect 17512 4576 18604 4604
rect 15703 4573 15715 4576
rect 15657 4567 15715 4573
rect 10134 4536 10140 4548
rect 4632 4508 5580 4536
rect 10095 4508 10140 4536
rect 4632 4480 4660 4508
rect 10134 4496 10140 4508
rect 10192 4496 10198 4548
rect 13446 4496 13452 4548
rect 13504 4536 13510 4548
rect 15672 4536 15700 4567
rect 18598 4564 18604 4576
rect 18656 4564 18662 4616
rect 19429 4607 19487 4613
rect 19429 4573 19441 4607
rect 19475 4573 19487 4607
rect 19812 4604 19840 4635
rect 20714 4632 20720 4644
rect 20772 4632 20778 4684
rect 20898 4672 20904 4684
rect 20859 4644 20904 4672
rect 20898 4632 20904 4644
rect 20956 4632 20962 4684
rect 21928 4681 21956 4712
rect 21913 4675 21971 4681
rect 21913 4641 21925 4675
rect 21959 4641 21971 4675
rect 21913 4635 21971 4641
rect 19978 4604 19984 4616
rect 19812 4576 19984 4604
rect 19429 4567 19487 4573
rect 13504 4508 15700 4536
rect 13504 4496 13510 4508
rect 16850 4496 16856 4548
rect 16908 4536 16914 4548
rect 16945 4539 17003 4545
rect 16945 4536 16957 4539
rect 16908 4508 16957 4536
rect 16908 4496 16914 4508
rect 16945 4505 16957 4508
rect 16991 4505 17003 4539
rect 16945 4499 17003 4505
rect 18138 4496 18144 4548
rect 18196 4536 18202 4548
rect 18966 4536 18972 4548
rect 18196 4508 18972 4536
rect 18196 4496 18202 4508
rect 18966 4496 18972 4508
rect 19024 4496 19030 4548
rect 19444 4536 19472 4567
rect 19978 4564 19984 4576
rect 20036 4604 20042 4616
rect 21729 4607 21787 4613
rect 21729 4604 21741 4607
rect 20036 4576 21741 4604
rect 20036 4564 20042 4576
rect 21729 4573 21741 4576
rect 21775 4573 21787 4607
rect 22112 4604 22140 4712
rect 22296 4712 22652 4740
rect 22296 4681 22324 4712
rect 22646 4700 22652 4712
rect 22704 4700 22710 4752
rect 22281 4675 22339 4681
rect 22281 4641 22293 4675
rect 22327 4641 22339 4675
rect 22281 4635 22339 4641
rect 22557 4675 22615 4681
rect 22557 4641 22569 4675
rect 22603 4672 22615 4675
rect 22922 4672 22928 4684
rect 22603 4644 22928 4672
rect 22603 4641 22615 4644
rect 22557 4635 22615 4641
rect 22922 4632 22928 4644
rect 22980 4632 22986 4684
rect 23290 4672 23296 4684
rect 23251 4644 23296 4672
rect 23290 4632 23296 4644
rect 23348 4632 23354 4684
rect 24118 4672 24124 4684
rect 24079 4644 24124 4672
rect 24118 4632 24124 4644
rect 24176 4632 24182 4684
rect 24228 4681 24256 4780
rect 30926 4768 30932 4780
rect 30984 4768 30990 4820
rect 31110 4808 31116 4820
rect 31071 4780 31116 4808
rect 31110 4768 31116 4780
rect 31168 4768 31174 4820
rect 31202 4768 31208 4820
rect 31260 4808 31266 4820
rect 32766 4808 32772 4820
rect 31260 4780 32772 4808
rect 31260 4768 31266 4780
rect 32766 4768 32772 4780
rect 32824 4768 32830 4820
rect 32950 4768 32956 4820
rect 33008 4808 33014 4820
rect 33008 4780 34468 4808
rect 33008 4768 33014 4780
rect 25222 4740 25228 4752
rect 25183 4712 25228 4740
rect 25222 4700 25228 4712
rect 25280 4700 25286 4752
rect 25590 4700 25596 4752
rect 25648 4740 25654 4752
rect 25869 4743 25927 4749
rect 25869 4740 25881 4743
rect 25648 4712 25881 4740
rect 25648 4700 25654 4712
rect 25869 4709 25881 4712
rect 25915 4709 25927 4743
rect 30374 4740 30380 4752
rect 25869 4703 25927 4709
rect 30024 4712 30380 4740
rect 24213 4675 24271 4681
rect 24213 4641 24225 4675
rect 24259 4641 24271 4675
rect 24670 4672 24676 4684
rect 24631 4644 24676 4672
rect 24213 4635 24271 4641
rect 24228 4604 24256 4635
rect 24670 4632 24676 4644
rect 24728 4632 24734 4684
rect 24857 4675 24915 4681
rect 24857 4641 24869 4675
rect 24903 4672 24915 4675
rect 24903 4644 25084 4672
rect 24903 4641 24915 4644
rect 24857 4635 24915 4641
rect 22112 4576 24256 4604
rect 25056 4604 25084 4644
rect 25498 4632 25504 4684
rect 25556 4672 25562 4684
rect 25777 4675 25835 4681
rect 25777 4672 25789 4675
rect 25556 4644 25789 4672
rect 25556 4632 25562 4644
rect 25777 4641 25789 4644
rect 25823 4641 25835 4675
rect 26786 4672 26792 4684
rect 26747 4644 26792 4672
rect 25777 4635 25835 4641
rect 26786 4632 26792 4644
rect 26844 4632 26850 4684
rect 27065 4675 27123 4681
rect 27065 4641 27077 4675
rect 27111 4672 27123 4675
rect 28902 4672 28908 4684
rect 27111 4644 28908 4672
rect 27111 4641 27123 4644
rect 27065 4635 27123 4641
rect 28902 4632 28908 4644
rect 28960 4632 28966 4684
rect 30024 4681 30052 4712
rect 30374 4700 30380 4712
rect 30432 4740 30438 4752
rect 31128 4740 31156 4768
rect 30432 4712 31156 4740
rect 32125 4743 32183 4749
rect 30432 4700 30438 4712
rect 32125 4709 32137 4743
rect 32171 4740 32183 4743
rect 32398 4740 32404 4752
rect 32171 4712 32404 4740
rect 32171 4709 32183 4712
rect 32125 4703 32183 4709
rect 32398 4700 32404 4712
rect 32456 4700 32462 4752
rect 32784 4740 32812 4768
rect 33594 4740 33600 4752
rect 32784 4712 32858 4740
rect 33555 4712 33600 4740
rect 30009 4675 30067 4681
rect 30009 4641 30021 4675
rect 30055 4641 30067 4675
rect 30009 4635 30067 4641
rect 30285 4675 30343 4681
rect 30285 4641 30297 4675
rect 30331 4641 30343 4675
rect 30285 4635 30343 4641
rect 30469 4675 30527 4681
rect 30469 4641 30481 4675
rect 30515 4672 30527 4675
rect 30834 4672 30840 4684
rect 30515 4644 30840 4672
rect 30515 4641 30527 4644
rect 30469 4635 30527 4641
rect 25682 4604 25688 4616
rect 25056 4576 25688 4604
rect 21729 4567 21787 4573
rect 25682 4564 25688 4576
rect 25740 4564 25746 4616
rect 28166 4604 28172 4616
rect 25792 4576 27752 4604
rect 28127 4576 28172 4604
rect 19886 4536 19892 4548
rect 19444 4508 19892 4536
rect 19886 4496 19892 4508
rect 19944 4496 19950 4548
rect 20070 4536 20076 4548
rect 20031 4508 20076 4536
rect 20070 4496 20076 4508
rect 20128 4496 20134 4548
rect 22462 4496 22468 4548
rect 22520 4536 22526 4548
rect 22738 4536 22744 4548
rect 22520 4508 22744 4536
rect 22520 4496 22526 4508
rect 22738 4496 22744 4508
rect 22796 4536 22802 4548
rect 25792 4536 25820 4576
rect 22796 4508 25820 4536
rect 27724 4536 27752 4576
rect 28166 4564 28172 4576
rect 28224 4564 28230 4616
rect 29457 4607 29515 4613
rect 29457 4573 29469 4607
rect 29503 4604 29515 4607
rect 29822 4604 29828 4616
rect 29503 4576 29828 4604
rect 29503 4573 29515 4576
rect 29457 4567 29515 4573
rect 29822 4564 29828 4576
rect 29880 4564 29886 4616
rect 30300 4604 30328 4635
rect 30834 4632 30840 4644
rect 30892 4632 30898 4684
rect 30926 4632 30932 4684
rect 30984 4672 30990 4684
rect 32674 4672 32680 4684
rect 30984 4644 31077 4672
rect 32635 4644 32680 4672
rect 30984 4632 30990 4644
rect 32674 4632 32680 4644
rect 32732 4632 32738 4684
rect 32830 4681 32858 4712
rect 33594 4700 33600 4712
rect 33652 4700 33658 4752
rect 33870 4700 33876 4752
rect 33928 4740 33934 4752
rect 34440 4740 34468 4780
rect 37274 4740 37280 4752
rect 33928 4712 34376 4740
rect 34440 4712 34652 4740
rect 33928 4700 33934 4712
rect 32815 4675 32873 4681
rect 32815 4641 32827 4675
rect 32861 4641 32873 4675
rect 32815 4635 32873 4641
rect 32953 4675 33011 4681
rect 32953 4641 32965 4675
rect 32999 4672 33011 4675
rect 34348 4672 34376 4712
rect 34624 4684 34652 4712
rect 35912 4712 37280 4740
rect 34425 4675 34483 4681
rect 34425 4672 34437 4675
rect 32999 4644 34284 4672
rect 34348 4644 34437 4672
rect 32999 4641 33011 4644
rect 32953 4635 33011 4641
rect 30650 4604 30656 4616
rect 30300 4576 30656 4604
rect 30300 4536 30328 4576
rect 30650 4564 30656 4576
rect 30708 4564 30714 4616
rect 30944 4604 30972 4632
rect 30852 4576 30972 4604
rect 27724 4508 30328 4536
rect 22796 4496 22802 4508
rect 4525 4471 4583 4477
rect 4525 4437 4537 4471
rect 4571 4468 4583 4471
rect 4614 4468 4620 4480
rect 4571 4440 4620 4468
rect 4571 4437 4583 4440
rect 4525 4431 4583 4437
rect 4614 4428 4620 4440
rect 4672 4428 4678 4480
rect 13814 4468 13820 4480
rect 13775 4440 13820 4468
rect 13814 4428 13820 4440
rect 13872 4428 13878 4480
rect 15930 4468 15936 4480
rect 15891 4440 15936 4468
rect 15930 4428 15936 4440
rect 15988 4428 15994 4480
rect 19334 4428 19340 4480
rect 19392 4468 19398 4480
rect 22554 4468 22560 4480
rect 19392 4440 22560 4468
rect 19392 4428 19398 4440
rect 22554 4428 22560 4440
rect 22612 4428 22618 4480
rect 23658 4428 23664 4480
rect 23716 4468 23722 4480
rect 30852 4468 30880 4576
rect 31018 4564 31024 4616
rect 31076 4604 31082 4616
rect 33870 4604 33876 4616
rect 31076 4576 33876 4604
rect 31076 4564 31082 4576
rect 33870 4564 33876 4576
rect 33928 4564 33934 4616
rect 34149 4607 34207 4613
rect 34149 4573 34161 4607
rect 34195 4573 34207 4607
rect 34256 4604 34284 4644
rect 34425 4641 34437 4644
rect 34471 4641 34483 4675
rect 34606 4672 34612 4684
rect 34519 4644 34612 4672
rect 34425 4635 34483 4641
rect 34606 4632 34612 4644
rect 34664 4632 34670 4684
rect 35434 4632 35440 4684
rect 35492 4672 35498 4684
rect 35912 4681 35940 4712
rect 37274 4700 37280 4712
rect 37332 4700 37338 4752
rect 35621 4675 35679 4681
rect 35621 4672 35633 4675
rect 35492 4644 35633 4672
rect 35492 4632 35498 4644
rect 35621 4641 35633 4644
rect 35667 4641 35679 4675
rect 35621 4635 35679 4641
rect 35897 4675 35955 4681
rect 35897 4641 35909 4675
rect 35943 4641 35955 4675
rect 36538 4672 36544 4684
rect 36499 4644 36544 4672
rect 35897 4635 35955 4641
rect 36538 4632 36544 4644
rect 36596 4632 36602 4684
rect 37734 4672 37740 4684
rect 37695 4644 37740 4672
rect 37734 4632 37740 4644
rect 37792 4632 37798 4684
rect 34514 4604 34520 4616
rect 34256 4576 34520 4604
rect 34149 4567 34207 4573
rect 32398 4496 32404 4548
rect 32456 4536 32462 4548
rect 34164 4536 34192 4567
rect 34514 4564 34520 4576
rect 34572 4564 34578 4616
rect 35069 4607 35127 4613
rect 35069 4573 35081 4607
rect 35115 4604 35127 4607
rect 35526 4604 35532 4616
rect 35115 4576 35532 4604
rect 35115 4573 35127 4576
rect 35069 4567 35127 4573
rect 35526 4564 35532 4576
rect 35584 4564 35590 4616
rect 36081 4607 36139 4613
rect 36081 4573 36093 4607
rect 36127 4573 36139 4607
rect 36081 4567 36139 4573
rect 34422 4536 34428 4548
rect 32456 4508 34428 4536
rect 32456 4496 32462 4508
rect 34422 4496 34428 4508
rect 34480 4496 34486 4548
rect 34532 4536 34560 4564
rect 36096 4536 36124 4567
rect 34532 4508 36124 4536
rect 23716 4440 30880 4468
rect 23716 4428 23722 4440
rect 33962 4428 33968 4480
rect 34020 4468 34026 4480
rect 35434 4468 35440 4480
rect 34020 4440 35440 4468
rect 34020 4428 34026 4440
rect 35434 4428 35440 4440
rect 35492 4468 35498 4480
rect 36725 4471 36783 4477
rect 36725 4468 36737 4471
rect 35492 4440 36737 4468
rect 35492 4428 35498 4440
rect 36725 4437 36737 4440
rect 36771 4468 36783 4471
rect 36998 4468 37004 4480
rect 36771 4440 37004 4468
rect 36771 4437 36783 4440
rect 36725 4431 36783 4437
rect 36998 4428 37004 4440
rect 37056 4428 37062 4480
rect 37918 4468 37924 4480
rect 37879 4440 37924 4468
rect 37918 4428 37924 4440
rect 37976 4428 37982 4480
rect 1104 4378 38824 4400
rect 1104 4326 4246 4378
rect 4298 4326 4310 4378
rect 4362 4326 4374 4378
rect 4426 4326 4438 4378
rect 4490 4326 34966 4378
rect 35018 4326 35030 4378
rect 35082 4326 35094 4378
rect 35146 4326 35158 4378
rect 35210 4326 38824 4378
rect 1104 4304 38824 4326
rect 7006 4224 7012 4276
rect 7064 4264 7070 4276
rect 8205 4267 8263 4273
rect 8205 4264 8217 4267
rect 7064 4236 8217 4264
rect 7064 4224 7070 4236
rect 8205 4233 8217 4236
rect 8251 4233 8263 4267
rect 8205 4227 8263 4233
rect 11238 4224 11244 4276
rect 11296 4264 11302 4276
rect 19426 4264 19432 4276
rect 11296 4236 19288 4264
rect 19387 4236 19432 4264
rect 11296 4224 11302 4236
rect 9490 4196 9496 4208
rect 9451 4168 9496 4196
rect 9490 4156 9496 4168
rect 9548 4156 9554 4208
rect 10686 4156 10692 4208
rect 10744 4196 10750 4208
rect 10744 4168 11652 4196
rect 10744 4156 10750 4168
rect 3234 4128 3240 4140
rect 3195 4100 3240 4128
rect 3234 4088 3240 4100
rect 3292 4088 3298 4140
rect 4614 4128 4620 4140
rect 3804 4100 4620 4128
rect 1854 4020 1860 4072
rect 1912 4060 1918 4072
rect 1949 4063 2007 4069
rect 1949 4060 1961 4063
rect 1912 4032 1961 4060
rect 1912 4020 1918 4032
rect 1949 4029 1961 4032
rect 1995 4029 2007 4063
rect 1949 4023 2007 4029
rect 2225 4063 2283 4069
rect 2225 4029 2237 4063
rect 2271 4029 2283 4063
rect 2958 4060 2964 4072
rect 2919 4032 2964 4060
rect 2225 4023 2283 4029
rect 1670 3884 1676 3936
rect 1728 3924 1734 3936
rect 1765 3927 1823 3933
rect 1765 3924 1777 3927
rect 1728 3896 1777 3924
rect 1728 3884 1734 3896
rect 1765 3893 1777 3896
rect 1811 3893 1823 3927
rect 1964 3924 1992 4023
rect 2240 3992 2268 4023
rect 2958 4020 2964 4032
rect 3016 4020 3022 4072
rect 3804 4060 3832 4100
rect 4614 4088 4620 4100
rect 4672 4088 4678 4140
rect 7101 4131 7159 4137
rect 7101 4097 7113 4131
rect 7147 4128 7159 4131
rect 7190 4128 7196 4140
rect 7147 4100 7196 4128
rect 7147 4097 7159 4100
rect 7101 4091 7159 4097
rect 7190 4088 7196 4100
rect 7248 4088 7254 4140
rect 10226 4128 10232 4140
rect 9600 4100 10232 4128
rect 5077 4063 5135 4069
rect 5077 4060 5089 4063
rect 3068 4032 3832 4060
rect 3896 4032 5089 4060
rect 3068 3992 3096 4032
rect 2240 3964 3096 3992
rect 3896 3924 3924 4032
rect 5077 4029 5089 4032
rect 5123 4029 5135 4063
rect 5077 4023 5135 4029
rect 5537 4063 5595 4069
rect 5537 4029 5549 4063
rect 5583 4029 5595 4063
rect 5537 4023 5595 4029
rect 6825 4063 6883 4069
rect 6825 4029 6837 4063
rect 6871 4060 6883 4063
rect 6914 4060 6920 4072
rect 6871 4032 6920 4060
rect 6871 4029 6883 4032
rect 6825 4023 6883 4029
rect 3970 3952 3976 4004
rect 4028 3992 4034 4004
rect 5552 3992 5580 4023
rect 6914 4020 6920 4032
rect 6972 4060 6978 4072
rect 7834 4060 7840 4072
rect 6972 4032 7840 4060
rect 6972 4020 6978 4032
rect 7834 4020 7840 4032
rect 7892 4020 7898 4072
rect 9600 4069 9628 4100
rect 10226 4088 10232 4100
rect 10284 4088 10290 4140
rect 10870 4128 10876 4140
rect 10428 4100 10876 4128
rect 9585 4063 9643 4069
rect 9585 4029 9597 4063
rect 9631 4029 9643 4063
rect 9858 4060 9864 4072
rect 9819 4032 9864 4060
rect 9585 4023 9643 4029
rect 9858 4020 9864 4032
rect 9916 4020 9922 4072
rect 10428 4069 10456 4100
rect 10870 4088 10876 4100
rect 10928 4088 10934 4140
rect 11514 4128 11520 4140
rect 11348 4100 11520 4128
rect 10413 4063 10471 4069
rect 10413 4029 10425 4063
rect 10459 4029 10471 4063
rect 10413 4023 10471 4029
rect 10502 4020 10508 4072
rect 10560 4060 10566 4072
rect 11348 4069 11376 4100
rect 11514 4088 11520 4100
rect 11572 4088 11578 4140
rect 11624 4128 11652 4168
rect 13814 4156 13820 4208
rect 13872 4156 13878 4208
rect 19260 4196 19288 4236
rect 19426 4224 19432 4236
rect 19484 4224 19490 4276
rect 21542 4264 21548 4276
rect 21503 4236 21548 4264
rect 21542 4224 21548 4236
rect 21600 4224 21606 4276
rect 26234 4224 26240 4276
rect 26292 4264 26298 4276
rect 27157 4267 27215 4273
rect 27157 4264 27169 4267
rect 26292 4236 27169 4264
rect 26292 4224 26298 4236
rect 27157 4233 27169 4236
rect 27203 4264 27215 4267
rect 31018 4264 31024 4276
rect 27203 4236 31024 4264
rect 27203 4233 27215 4236
rect 27157 4227 27215 4233
rect 31018 4224 31024 4236
rect 31076 4224 31082 4276
rect 32214 4224 32220 4276
rect 32272 4264 32278 4276
rect 37274 4264 37280 4276
rect 32272 4236 34192 4264
rect 32272 4224 32278 4236
rect 19334 4196 19340 4208
rect 19260 4168 19340 4196
rect 19334 4156 19340 4168
rect 19392 4156 19398 4208
rect 22094 4156 22100 4208
rect 22152 4196 22158 4208
rect 30650 4196 30656 4208
rect 22152 4168 23796 4196
rect 30611 4168 30656 4196
rect 22152 4156 22158 4168
rect 12529 4131 12587 4137
rect 12529 4128 12541 4131
rect 11624 4100 12541 4128
rect 12529 4097 12541 4100
rect 12575 4097 12587 4131
rect 13832 4128 13860 4156
rect 15010 4128 15016 4140
rect 12529 4091 12587 4097
rect 13096 4100 13860 4128
rect 14971 4100 15016 4128
rect 10597 4063 10655 4069
rect 10597 4060 10609 4063
rect 10560 4032 10609 4060
rect 10560 4020 10566 4032
rect 10597 4029 10609 4032
rect 10643 4029 10655 4063
rect 10597 4023 10655 4029
rect 11333 4063 11391 4069
rect 11333 4029 11345 4063
rect 11379 4029 11391 4063
rect 11333 4023 11391 4029
rect 11422 4020 11428 4072
rect 11480 4060 11486 4072
rect 13096 4069 13124 4100
rect 15010 4088 15016 4100
rect 15068 4088 15074 4140
rect 15470 4088 15476 4140
rect 15528 4128 15534 4140
rect 16117 4131 16175 4137
rect 16117 4128 16129 4131
rect 15528 4100 16129 4128
rect 15528 4088 15534 4100
rect 16117 4097 16129 4100
rect 16163 4097 16175 4131
rect 16117 4091 16175 4097
rect 18325 4131 18383 4137
rect 18325 4097 18337 4131
rect 18371 4128 18383 4131
rect 20070 4128 20076 4140
rect 18371 4100 20076 4128
rect 18371 4097 18383 4100
rect 18325 4091 18383 4097
rect 20070 4088 20076 4100
rect 20128 4088 20134 4140
rect 23661 4131 23719 4137
rect 23661 4097 23673 4131
rect 23707 4128 23719 4131
rect 23768 4128 23796 4168
rect 30650 4156 30656 4168
rect 30708 4156 30714 4208
rect 33962 4196 33968 4208
rect 33704 4168 33968 4196
rect 24854 4128 24860 4140
rect 23707 4100 23796 4128
rect 24815 4100 24860 4128
rect 23707 4097 23719 4100
rect 23661 4091 23719 4097
rect 24854 4088 24860 4100
rect 24912 4088 24918 4140
rect 28721 4131 28779 4137
rect 24964 4100 28672 4128
rect 12437 4063 12495 4069
rect 12437 4060 12449 4063
rect 11480 4032 12449 4060
rect 11480 4020 11486 4032
rect 12437 4029 12449 4032
rect 12483 4029 12495 4063
rect 12437 4023 12495 4029
rect 13081 4063 13139 4069
rect 13081 4029 13093 4063
rect 13127 4029 13139 4063
rect 13081 4023 13139 4029
rect 13725 4063 13783 4069
rect 13725 4029 13737 4063
rect 13771 4029 13783 4063
rect 13725 4023 13783 4029
rect 13858 4063 13916 4069
rect 13858 4029 13870 4063
rect 13904 4060 13916 4063
rect 13998 4060 14004 4072
rect 13904 4032 14004 4060
rect 13904 4029 13916 4032
rect 13858 4023 13916 4029
rect 13740 3992 13768 4023
rect 13998 4020 14004 4032
rect 14056 4020 14062 4072
rect 14734 4060 14740 4072
rect 14695 4032 14740 4060
rect 14734 4020 14740 4032
rect 14792 4020 14798 4072
rect 16942 4060 16948 4072
rect 16903 4032 16948 4060
rect 16942 4020 16948 4032
rect 17000 4020 17006 4072
rect 17034 4020 17040 4072
rect 17092 4060 17098 4072
rect 18046 4060 18052 4072
rect 17092 4032 17137 4060
rect 18007 4032 18052 4060
rect 17092 4020 17098 4032
rect 18046 4020 18052 4032
rect 18104 4020 18110 4072
rect 20162 4060 20168 4072
rect 20123 4032 20168 4060
rect 20162 4020 20168 4032
rect 20220 4020 20226 4072
rect 20438 4060 20444 4072
rect 20399 4032 20444 4060
rect 20438 4020 20444 4032
rect 20496 4020 20502 4072
rect 22094 4020 22100 4072
rect 22152 4060 22158 4072
rect 22281 4063 22339 4069
rect 22281 4060 22293 4063
rect 22152 4032 22293 4060
rect 22152 4020 22158 4032
rect 22281 4029 22293 4032
rect 22327 4029 22339 4063
rect 22281 4023 22339 4029
rect 22370 4020 22376 4072
rect 22428 4060 22434 4072
rect 22428 4032 22473 4060
rect 22428 4020 22434 4032
rect 22554 4020 22560 4072
rect 22612 4060 22618 4072
rect 23753 4063 23811 4069
rect 23753 4060 23765 4063
rect 22612 4032 23765 4060
rect 22612 4020 22618 4032
rect 23753 4029 23765 4032
rect 23799 4029 23811 4063
rect 23753 4023 23811 4029
rect 24578 4020 24584 4072
rect 24636 4060 24642 4072
rect 24964 4060 24992 4100
rect 24636 4032 24992 4060
rect 25133 4063 25191 4069
rect 24636 4020 24642 4032
rect 25133 4029 25145 4063
rect 25179 4060 25191 4063
rect 25774 4060 25780 4072
rect 25179 4032 25780 4060
rect 25179 4029 25191 4032
rect 25133 4023 25191 4029
rect 25774 4020 25780 4032
rect 25832 4020 25838 4072
rect 26878 4020 26884 4072
rect 26936 4060 26942 4072
rect 26973 4063 27031 4069
rect 26973 4060 26985 4063
rect 26936 4032 26985 4060
rect 26936 4020 26942 4032
rect 26973 4029 26985 4032
rect 27019 4029 27031 4063
rect 26973 4023 27031 4029
rect 28261 4063 28319 4069
rect 28261 4029 28273 4063
rect 28307 4060 28319 4063
rect 28442 4060 28448 4072
rect 28307 4032 28448 4060
rect 28307 4029 28319 4032
rect 28261 4023 28319 4029
rect 28442 4020 28448 4032
rect 28500 4020 28506 4072
rect 28537 4063 28595 4069
rect 28537 4029 28549 4063
rect 28583 4029 28595 4063
rect 28644 4060 28672 4100
rect 28721 4097 28733 4131
rect 28767 4128 28779 4131
rect 29086 4128 29092 4140
rect 28767 4100 29092 4128
rect 28767 4097 28779 4100
rect 28721 4091 28779 4097
rect 29086 4088 29092 4100
rect 29144 4088 29150 4140
rect 29178 4088 29184 4140
rect 29236 4128 29242 4140
rect 29273 4131 29331 4137
rect 29273 4128 29285 4131
rect 29236 4100 29285 4128
rect 29236 4088 29242 4100
rect 29273 4097 29285 4100
rect 29319 4128 29331 4131
rect 30282 4128 30288 4140
rect 29319 4100 30288 4128
rect 29319 4097 29331 4100
rect 29273 4091 29331 4097
rect 30282 4088 30288 4100
rect 30340 4088 30346 4140
rect 32217 4131 32275 4137
rect 32217 4097 32229 4131
rect 32263 4128 32275 4131
rect 32398 4128 32404 4140
rect 32263 4100 32404 4128
rect 32263 4097 32275 4100
rect 32217 4091 32275 4097
rect 32398 4088 32404 4100
rect 32456 4088 32462 4140
rect 32674 4128 32680 4140
rect 32635 4100 32680 4128
rect 32674 4088 32680 4100
rect 32732 4088 32738 4140
rect 33704 4137 33732 4168
rect 33962 4156 33968 4168
rect 34020 4156 34026 4208
rect 34164 4137 34192 4236
rect 35912 4236 37280 4264
rect 35912 4196 35940 4236
rect 37274 4224 37280 4236
rect 37332 4224 37338 4276
rect 34532 4168 35940 4196
rect 33689 4131 33747 4137
rect 33689 4097 33701 4131
rect 33735 4097 33747 4131
rect 33689 4091 33747 4097
rect 34149 4131 34207 4137
rect 34149 4097 34161 4131
rect 34195 4128 34207 4131
rect 34330 4128 34336 4140
rect 34195 4100 34336 4128
rect 34195 4097 34207 4100
rect 34149 4091 34207 4097
rect 34330 4088 34336 4100
rect 34388 4088 34394 4140
rect 34532 4128 34560 4168
rect 34440 4100 34560 4128
rect 29362 4060 29368 4072
rect 28644 4032 29368 4060
rect 28537 4023 28595 4029
rect 14182 3992 14188 4004
rect 4028 3964 5580 3992
rect 12544 3964 14188 3992
rect 4028 3952 4034 3964
rect 1964 3896 3924 3924
rect 4525 3927 4583 3933
rect 1765 3887 1823 3893
rect 4525 3893 4537 3927
rect 4571 3924 4583 3927
rect 4798 3924 4804 3936
rect 4571 3896 4804 3924
rect 4571 3893 4583 3896
rect 4525 3887 4583 3893
rect 4798 3884 4804 3896
rect 4856 3884 4862 3936
rect 5166 3924 5172 3936
rect 5127 3896 5172 3924
rect 5166 3884 5172 3896
rect 5224 3884 5230 3936
rect 7374 3884 7380 3936
rect 7432 3924 7438 3936
rect 12544 3924 12572 3964
rect 14182 3952 14188 3964
rect 14240 3952 14246 4004
rect 14277 3995 14335 4001
rect 14277 3961 14289 3995
rect 14323 3961 14335 3995
rect 14277 3955 14335 3961
rect 17497 3995 17555 4001
rect 17497 3961 17509 3995
rect 17543 3961 17555 3995
rect 17497 3955 17555 3961
rect 7432 3896 12572 3924
rect 7432 3884 7438 3896
rect 12618 3884 12624 3936
rect 12676 3924 12682 3936
rect 13173 3927 13231 3933
rect 13173 3924 13185 3927
rect 12676 3896 13185 3924
rect 12676 3884 12682 3896
rect 13173 3893 13185 3896
rect 13219 3893 13231 3927
rect 14292 3924 14320 3955
rect 16022 3924 16028 3936
rect 14292 3896 16028 3924
rect 13173 3887 13231 3893
rect 16022 3884 16028 3896
rect 16080 3884 16086 3936
rect 17512 3924 17540 3955
rect 19058 3952 19064 4004
rect 19116 3992 19122 4004
rect 20070 3992 20076 4004
rect 19116 3964 20076 3992
rect 19116 3952 19122 3964
rect 20070 3952 20076 3964
rect 20128 3952 20134 4004
rect 22833 3995 22891 4001
rect 22833 3961 22845 3995
rect 22879 3992 22891 3995
rect 24118 3992 24124 4004
rect 22879 3964 24124 3992
rect 22879 3961 22891 3964
rect 22833 3955 22891 3961
rect 24118 3952 24124 3964
rect 24176 3952 24182 4004
rect 24213 3995 24271 4001
rect 24213 3961 24225 3995
rect 24259 3992 24271 3995
rect 24854 3992 24860 4004
rect 24259 3964 24860 3992
rect 24259 3961 24271 3964
rect 24213 3955 24271 3961
rect 24854 3952 24860 3964
rect 24912 3952 24918 4004
rect 26510 3992 26516 4004
rect 26471 3964 26516 3992
rect 26510 3952 26516 3964
rect 26568 3952 26574 4004
rect 27709 3995 27767 4001
rect 27709 3961 27721 3995
rect 27755 3992 27767 3995
rect 28074 3992 28080 4004
rect 27755 3964 28080 3992
rect 27755 3961 27767 3964
rect 27709 3955 27767 3961
rect 28074 3952 28080 3964
rect 28132 3952 28138 4004
rect 19242 3924 19248 3936
rect 17512 3896 19248 3924
rect 19242 3884 19248 3896
rect 19300 3884 19306 3936
rect 19426 3884 19432 3936
rect 19484 3924 19490 3936
rect 22002 3924 22008 3936
rect 19484 3896 22008 3924
rect 19484 3884 19490 3896
rect 22002 3884 22008 3896
rect 22060 3884 22066 3936
rect 28552 3924 28580 4023
rect 29362 4020 29368 4032
rect 29420 4020 29426 4072
rect 29546 4060 29552 4072
rect 29507 4032 29552 4060
rect 29546 4020 29552 4032
rect 29604 4020 29610 4072
rect 32493 4063 32551 4069
rect 32493 4029 32505 4063
rect 32539 4060 32551 4063
rect 33965 4063 34023 4069
rect 33965 4060 33977 4063
rect 32539 4032 33977 4060
rect 32539 4029 32551 4032
rect 32493 4023 32551 4029
rect 33965 4029 33977 4032
rect 34011 4060 34023 4063
rect 34238 4060 34244 4072
rect 34011 4032 34244 4060
rect 34011 4029 34023 4032
rect 33965 4023 34023 4029
rect 34238 4020 34244 4032
rect 34296 4060 34302 4072
rect 34440 4060 34468 4100
rect 35710 4088 35716 4140
rect 35768 4128 35774 4140
rect 37461 4131 37519 4137
rect 37461 4128 37473 4131
rect 35768 4100 37473 4128
rect 35768 4088 35774 4100
rect 37461 4097 37473 4100
rect 37507 4097 37519 4131
rect 37461 4091 37519 4097
rect 34296 4032 34468 4060
rect 34977 4063 35035 4069
rect 34296 4020 34302 4032
rect 34977 4029 34989 4063
rect 35023 4060 35035 4063
rect 35894 4060 35900 4072
rect 35023 4032 35900 4060
rect 35023 4029 35035 4032
rect 34977 4023 35035 4029
rect 35894 4020 35900 4032
rect 35952 4020 35958 4072
rect 36078 4060 36084 4072
rect 36039 4032 36084 4060
rect 36078 4020 36084 4032
rect 36136 4020 36142 4072
rect 36357 4063 36415 4069
rect 36357 4060 36369 4063
rect 36188 4032 36369 4060
rect 31665 3995 31723 4001
rect 31665 3961 31677 3995
rect 31711 3961 31723 3995
rect 31665 3955 31723 3961
rect 33137 3995 33195 4001
rect 33137 3961 33149 3995
rect 33183 3992 33195 3995
rect 35434 3992 35440 4004
rect 33183 3964 35440 3992
rect 33183 3961 33195 3964
rect 33137 3955 33195 3961
rect 30190 3924 30196 3936
rect 28552 3896 30196 3924
rect 30190 3884 30196 3896
rect 30248 3884 30254 3936
rect 31680 3924 31708 3955
rect 35434 3952 35440 3964
rect 35492 3952 35498 4004
rect 35618 3952 35624 4004
rect 35676 3992 35682 4004
rect 36188 3992 36216 4032
rect 36357 4029 36369 4032
rect 36403 4029 36415 4063
rect 36357 4023 36415 4029
rect 35676 3964 36216 3992
rect 35676 3952 35682 3964
rect 33870 3924 33876 3936
rect 31680 3896 33876 3924
rect 33870 3884 33876 3896
rect 33928 3884 33934 3936
rect 34606 3884 34612 3936
rect 34664 3924 34670 3936
rect 35161 3927 35219 3933
rect 35161 3924 35173 3927
rect 34664 3896 35173 3924
rect 34664 3884 34670 3896
rect 35161 3893 35173 3896
rect 35207 3893 35219 3927
rect 35161 3887 35219 3893
rect 1104 3834 38824 3856
rect 1104 3782 19606 3834
rect 19658 3782 19670 3834
rect 19722 3782 19734 3834
rect 19786 3782 19798 3834
rect 19850 3782 38824 3834
rect 1104 3760 38824 3782
rect 2958 3680 2964 3732
rect 3016 3720 3022 3732
rect 6546 3720 6552 3732
rect 3016 3692 5304 3720
rect 6507 3692 6552 3720
rect 3016 3680 3022 3692
rect 5166 3652 5172 3664
rect 3436 3624 5172 3652
rect 2133 3587 2191 3593
rect 2133 3553 2145 3587
rect 2179 3584 2191 3587
rect 3436 3584 3464 3624
rect 5166 3612 5172 3624
rect 5224 3612 5230 3664
rect 2179 3556 3464 3584
rect 3513 3587 3571 3593
rect 2179 3553 2191 3556
rect 2133 3547 2191 3553
rect 3513 3553 3525 3587
rect 3559 3584 3571 3587
rect 4249 3587 4307 3593
rect 4249 3584 4261 3587
rect 3559 3556 4261 3584
rect 3559 3553 3571 3556
rect 3513 3547 3571 3553
rect 4249 3553 4261 3556
rect 4295 3553 4307 3587
rect 4249 3547 4307 3553
rect 1394 3476 1400 3528
rect 1452 3516 1458 3528
rect 1857 3519 1915 3525
rect 1857 3516 1869 3519
rect 1452 3488 1869 3516
rect 1452 3476 1458 3488
rect 1857 3485 1869 3488
rect 1903 3516 1915 3519
rect 2590 3516 2596 3528
rect 1903 3488 2596 3516
rect 1903 3485 1915 3488
rect 1857 3479 1915 3485
rect 2590 3476 2596 3488
rect 2648 3476 2654 3528
rect 3418 3476 3424 3528
rect 3476 3516 3482 3528
rect 4062 3516 4068 3528
rect 3476 3488 4068 3516
rect 3476 3476 3482 3488
rect 4062 3476 4068 3488
rect 4120 3516 4126 3528
rect 4157 3519 4215 3525
rect 4157 3516 4169 3519
rect 4120 3488 4169 3516
rect 4120 3476 4126 3488
rect 4157 3485 4169 3488
rect 4203 3485 4215 3519
rect 4706 3516 4712 3528
rect 4667 3488 4712 3516
rect 4157 3479 4215 3485
rect 4706 3476 4712 3488
rect 4764 3476 4770 3528
rect 5169 3519 5227 3525
rect 5169 3485 5181 3519
rect 5215 3516 5227 3519
rect 5276 3516 5304 3692
rect 6546 3680 6552 3692
rect 6604 3680 6610 3732
rect 11977 3723 12035 3729
rect 7300 3692 11836 3720
rect 5442 3584 5448 3596
rect 5403 3556 5448 3584
rect 5442 3544 5448 3556
rect 5500 3544 5506 3596
rect 5810 3544 5816 3596
rect 5868 3584 5874 3596
rect 7300 3584 7328 3692
rect 9766 3652 9772 3664
rect 8956 3624 9772 3652
rect 7466 3584 7472 3596
rect 5868 3556 7328 3584
rect 7427 3556 7472 3584
rect 5868 3544 5874 3556
rect 7466 3544 7472 3556
rect 7524 3544 7530 3596
rect 8662 3584 8668 3596
rect 8623 3556 8668 3584
rect 8662 3544 8668 3556
rect 8720 3544 8726 3596
rect 8956 3593 8984 3624
rect 9766 3612 9772 3624
rect 9824 3612 9830 3664
rect 11808 3593 11836 3692
rect 11977 3689 11989 3723
rect 12023 3720 12035 3723
rect 12618 3720 12624 3732
rect 12023 3692 12624 3720
rect 12023 3689 12035 3692
rect 11977 3683 12035 3689
rect 12618 3680 12624 3692
rect 12676 3720 12682 3732
rect 13446 3720 13452 3732
rect 12676 3692 13452 3720
rect 12676 3680 12682 3692
rect 13446 3680 13452 3692
rect 13504 3680 13510 3732
rect 14826 3680 14832 3732
rect 14884 3720 14890 3732
rect 15381 3723 15439 3729
rect 15381 3720 15393 3723
rect 14884 3692 15393 3720
rect 14884 3680 14890 3692
rect 15381 3689 15393 3692
rect 15427 3689 15439 3723
rect 15381 3683 15439 3689
rect 16022 3680 16028 3732
rect 16080 3720 16086 3732
rect 25590 3720 25596 3732
rect 16080 3692 25596 3720
rect 16080 3680 16086 3692
rect 25590 3680 25596 3692
rect 25648 3680 25654 3732
rect 25774 3720 25780 3732
rect 25735 3692 25780 3720
rect 25774 3680 25780 3692
rect 25832 3680 25838 3732
rect 26605 3723 26663 3729
rect 26605 3689 26617 3723
rect 26651 3720 26663 3723
rect 27246 3720 27252 3732
rect 26651 3692 27252 3720
rect 26651 3689 26663 3692
rect 26605 3683 26663 3689
rect 19334 3612 19340 3664
rect 19392 3652 19398 3664
rect 20349 3655 20407 3661
rect 19392 3624 19656 3652
rect 19392 3612 19398 3624
rect 8941 3587 8999 3593
rect 8941 3553 8953 3587
rect 8987 3553 8999 3587
rect 8941 3547 8999 3553
rect 9125 3587 9183 3593
rect 9125 3553 9137 3587
rect 9171 3584 9183 3587
rect 9953 3587 10011 3593
rect 9953 3584 9965 3587
rect 9171 3556 9965 3584
rect 9171 3553 9183 3556
rect 9125 3547 9183 3553
rect 9953 3553 9965 3556
rect 9999 3553 10011 3587
rect 9953 3547 10011 3553
rect 11793 3587 11851 3593
rect 11793 3553 11805 3587
rect 11839 3553 11851 3587
rect 11793 3547 11851 3553
rect 12250 3544 12256 3596
rect 12308 3584 12314 3596
rect 12802 3584 12808 3596
rect 12308 3556 12664 3584
rect 12763 3556 12808 3584
rect 12308 3544 12314 3556
rect 6914 3516 6920 3528
rect 5215 3488 6920 3516
rect 5215 3485 5227 3488
rect 5169 3479 5227 3485
rect 6914 3476 6920 3488
rect 6972 3476 6978 3528
rect 7374 3516 7380 3528
rect 7335 3488 7380 3516
rect 7374 3476 7380 3488
rect 7432 3476 7438 3528
rect 7926 3516 7932 3528
rect 7887 3488 7932 3516
rect 7926 3476 7932 3488
rect 7984 3476 7990 3528
rect 9306 3476 9312 3528
rect 9364 3516 9370 3528
rect 9677 3519 9735 3525
rect 9677 3516 9689 3519
rect 9364 3488 9689 3516
rect 9364 3476 9370 3488
rect 9677 3485 9689 3488
rect 9723 3516 9735 3519
rect 11333 3519 11391 3525
rect 9723 3488 11284 3516
rect 9723 3485 9735 3488
rect 9677 3479 9735 3485
rect 6822 3408 6828 3460
rect 6880 3448 6886 3460
rect 9324 3448 9352 3476
rect 6880 3420 9352 3448
rect 11256 3448 11284 3488
rect 11333 3485 11345 3519
rect 11379 3516 11391 3519
rect 12434 3516 12440 3528
rect 11379 3488 12440 3516
rect 11379 3485 11391 3488
rect 11333 3479 11391 3485
rect 12434 3476 12440 3488
rect 12492 3476 12498 3528
rect 12529 3519 12587 3525
rect 12529 3485 12541 3519
rect 12575 3485 12587 3519
rect 12636 3516 12664 3556
rect 12802 3544 12808 3556
rect 12860 3544 12866 3596
rect 15286 3584 15292 3596
rect 14660 3556 15292 3584
rect 14660 3516 14688 3556
rect 15286 3544 15292 3556
rect 15344 3544 15350 3596
rect 15562 3544 15568 3596
rect 15620 3584 15626 3596
rect 15838 3584 15844 3596
rect 15620 3556 15844 3584
rect 15620 3544 15626 3556
rect 15838 3544 15844 3556
rect 15896 3544 15902 3596
rect 16850 3584 16856 3596
rect 16811 3556 16856 3584
rect 16850 3544 16856 3556
rect 16908 3544 16914 3596
rect 16942 3544 16948 3596
rect 17000 3584 17006 3596
rect 19426 3584 19432 3596
rect 17000 3556 19432 3584
rect 17000 3544 17006 3556
rect 19426 3544 19432 3556
rect 19484 3544 19490 3596
rect 19628 3593 19656 3624
rect 20349 3621 20361 3655
rect 20395 3652 20407 3655
rect 20438 3652 20444 3664
rect 20395 3624 20444 3652
rect 20395 3621 20407 3624
rect 20349 3615 20407 3621
rect 20438 3612 20444 3624
rect 20496 3612 20502 3664
rect 21542 3652 21548 3664
rect 21192 3624 21548 3652
rect 21192 3593 21220 3624
rect 21542 3612 21548 3624
rect 21600 3612 21606 3664
rect 24026 3652 24032 3664
rect 22940 3624 24032 3652
rect 19613 3587 19671 3593
rect 19613 3553 19625 3587
rect 19659 3553 19671 3587
rect 19613 3547 19671 3553
rect 20165 3587 20223 3593
rect 20165 3553 20177 3587
rect 20211 3553 20223 3587
rect 20165 3547 20223 3553
rect 21177 3587 21235 3593
rect 21177 3553 21189 3587
rect 21223 3553 21235 3587
rect 21177 3547 21235 3553
rect 12636 3488 14688 3516
rect 12529 3479 12587 3485
rect 12342 3448 12348 3460
rect 11256 3420 12348 3448
rect 6880 3408 6886 3420
rect 12342 3408 12348 3420
rect 12400 3448 12406 3460
rect 12544 3448 12572 3479
rect 14734 3476 14740 3528
rect 14792 3516 14798 3528
rect 16577 3519 16635 3525
rect 16577 3516 16589 3519
rect 14792 3488 16589 3516
rect 14792 3476 14798 3488
rect 16577 3485 16589 3488
rect 16623 3516 16635 3519
rect 19337 3519 19395 3525
rect 16623 3488 18092 3516
rect 16623 3485 16635 3488
rect 16577 3479 16635 3485
rect 18064 3460 18092 3488
rect 19337 3485 19349 3519
rect 19383 3516 19395 3519
rect 19886 3516 19892 3528
rect 19383 3488 19892 3516
rect 19383 3485 19395 3488
rect 19337 3479 19395 3485
rect 19886 3476 19892 3488
rect 19944 3476 19950 3528
rect 20180 3516 20208 3547
rect 21266 3544 21272 3596
rect 21324 3584 21330 3596
rect 21634 3584 21640 3596
rect 21324 3556 21369 3584
rect 21595 3556 21640 3584
rect 21324 3544 21330 3556
rect 21634 3544 21640 3556
rect 21692 3544 21698 3596
rect 22738 3584 22744 3596
rect 22699 3556 22744 3584
rect 22738 3544 22744 3556
rect 22796 3544 22802 3596
rect 22940 3593 22968 3624
rect 24026 3612 24032 3624
rect 24084 3652 24090 3664
rect 26620 3652 26648 3683
rect 27246 3680 27252 3692
rect 27304 3680 27310 3732
rect 28442 3680 28448 3732
rect 28500 3720 28506 3732
rect 28500 3692 29960 3720
rect 28500 3680 28506 3692
rect 24084 3624 24808 3652
rect 24084 3612 24090 3624
rect 22925 3587 22983 3593
rect 22925 3553 22937 3587
rect 22971 3553 22983 3587
rect 22925 3547 22983 3553
rect 23014 3544 23020 3596
rect 23072 3584 23078 3596
rect 23385 3587 23443 3593
rect 23385 3584 23397 3587
rect 23072 3556 23397 3584
rect 23072 3544 23078 3556
rect 23385 3553 23397 3556
rect 23431 3553 23443 3587
rect 23385 3547 23443 3553
rect 23477 3587 23535 3593
rect 23477 3553 23489 3587
rect 23523 3584 23535 3587
rect 24670 3584 24676 3596
rect 23523 3556 24676 3584
rect 23523 3553 23535 3556
rect 23477 3547 23535 3553
rect 24670 3544 24676 3556
rect 24728 3544 24734 3596
rect 24780 3593 24808 3624
rect 25516 3624 26648 3652
rect 25516 3593 25544 3624
rect 29362 3612 29368 3664
rect 29420 3652 29426 3664
rect 29932 3661 29960 3692
rect 30190 3680 30196 3732
rect 30248 3720 30254 3732
rect 36265 3723 36323 3729
rect 36265 3720 36277 3723
rect 30248 3692 36277 3720
rect 30248 3680 30254 3692
rect 36265 3689 36277 3692
rect 36311 3689 36323 3723
rect 36265 3683 36323 3689
rect 29457 3655 29515 3661
rect 29457 3652 29469 3655
rect 29420 3624 29469 3652
rect 29420 3612 29426 3624
rect 29457 3621 29469 3624
rect 29503 3621 29515 3655
rect 29457 3615 29515 3621
rect 29917 3655 29975 3661
rect 29917 3621 29929 3655
rect 29963 3621 29975 3655
rect 29917 3615 29975 3621
rect 34425 3655 34483 3661
rect 34425 3621 34437 3655
rect 34471 3652 34483 3655
rect 34514 3652 34520 3664
rect 34471 3624 34520 3652
rect 34471 3621 34483 3624
rect 34425 3615 34483 3621
rect 24765 3587 24823 3593
rect 24765 3553 24777 3587
rect 24811 3553 24823 3587
rect 25317 3587 25375 3593
rect 25317 3584 25329 3587
rect 24765 3547 24823 3553
rect 24872 3556 25329 3584
rect 20993 3519 21051 3525
rect 20993 3516 21005 3519
rect 20180 3488 21005 3516
rect 20993 3485 21005 3488
rect 21039 3485 21051 3519
rect 24578 3516 24584 3528
rect 24539 3488 24584 3516
rect 20993 3479 21051 3485
rect 24578 3476 24584 3488
rect 24636 3476 24642 3528
rect 24688 3516 24716 3544
rect 24872 3516 24900 3556
rect 25317 3553 25329 3556
rect 25363 3553 25375 3587
rect 25317 3547 25375 3553
rect 25501 3587 25559 3593
rect 25501 3553 25513 3587
rect 25547 3553 25559 3587
rect 26510 3584 26516 3596
rect 26471 3556 26516 3584
rect 25501 3547 25559 3553
rect 26510 3544 26516 3556
rect 26568 3544 26574 3596
rect 27154 3584 27160 3596
rect 27115 3556 27160 3584
rect 27154 3544 27160 3556
rect 27212 3544 27218 3596
rect 28074 3584 28080 3596
rect 28035 3556 28080 3584
rect 28074 3544 28080 3556
rect 28132 3544 28138 3596
rect 24688 3488 24900 3516
rect 27801 3519 27859 3525
rect 27801 3485 27813 3519
rect 27847 3516 27859 3519
rect 29178 3516 29184 3528
rect 27847 3488 29184 3516
rect 27847 3485 27859 3488
rect 27801 3479 27859 3485
rect 29178 3476 29184 3488
rect 29236 3476 29242 3528
rect 29472 3516 29500 3615
rect 34514 3612 34520 3624
rect 34572 3612 34578 3664
rect 36280 3652 36308 3683
rect 37274 3680 37280 3732
rect 37332 3720 37338 3732
rect 37921 3723 37979 3729
rect 37921 3720 37933 3723
rect 37332 3692 37933 3720
rect 37332 3680 37338 3692
rect 37921 3689 37933 3692
rect 37967 3689 37979 3723
rect 37921 3683 37979 3689
rect 37458 3652 37464 3664
rect 36280 3624 37464 3652
rect 37458 3612 37464 3624
rect 37516 3612 37522 3664
rect 30374 3544 30380 3596
rect 30432 3584 30438 3596
rect 30469 3587 30527 3593
rect 30469 3584 30481 3587
rect 30432 3556 30481 3584
rect 30432 3544 30438 3556
rect 30469 3553 30481 3556
rect 30515 3553 30527 3587
rect 30469 3547 30527 3553
rect 30745 3587 30803 3593
rect 30745 3553 30757 3587
rect 30791 3553 30803 3587
rect 30745 3547 30803 3553
rect 30760 3516 30788 3547
rect 33318 3544 33324 3596
rect 33376 3584 33382 3596
rect 35161 3587 35219 3593
rect 35161 3584 35173 3587
rect 33376 3556 35173 3584
rect 33376 3544 33382 3556
rect 35161 3553 35173 3556
rect 35207 3553 35219 3587
rect 35161 3547 35219 3553
rect 37550 3544 37556 3596
rect 37608 3584 37614 3596
rect 37737 3587 37795 3593
rect 37737 3584 37749 3587
rect 37608 3556 37749 3584
rect 37608 3544 37614 3556
rect 37737 3553 37749 3556
rect 37783 3553 37795 3587
rect 37737 3547 37795 3553
rect 29472 3488 30788 3516
rect 30929 3519 30987 3525
rect 30929 3485 30941 3519
rect 30975 3516 30987 3519
rect 31754 3516 31760 3528
rect 30975 3488 31760 3516
rect 30975 3485 30987 3488
rect 30929 3479 30987 3485
rect 31754 3476 31760 3488
rect 31812 3476 31818 3528
rect 32122 3476 32128 3528
rect 32180 3516 32186 3528
rect 32766 3516 32772 3528
rect 32180 3488 32772 3516
rect 32180 3476 32186 3488
rect 32766 3476 32772 3488
rect 32824 3476 32830 3528
rect 33045 3519 33103 3525
rect 33045 3485 33057 3519
rect 33091 3516 33103 3519
rect 34422 3516 34428 3528
rect 33091 3488 34428 3516
rect 33091 3485 33103 3488
rect 33045 3479 33103 3485
rect 34422 3476 34428 3488
rect 34480 3476 34486 3528
rect 34698 3476 34704 3528
rect 34756 3516 34762 3528
rect 34885 3519 34943 3525
rect 34885 3516 34897 3519
rect 34756 3488 34897 3516
rect 34756 3476 34762 3488
rect 34885 3485 34897 3488
rect 34931 3516 34943 3519
rect 36078 3516 36084 3528
rect 34931 3488 36084 3516
rect 34931 3485 34943 3488
rect 34885 3479 34943 3485
rect 36078 3476 36084 3488
rect 36136 3476 36142 3528
rect 17954 3448 17960 3460
rect 12400 3420 12572 3448
rect 17915 3420 17960 3448
rect 12400 3408 12406 3420
rect 17954 3408 17960 3420
rect 18012 3408 18018 3460
rect 18046 3408 18052 3460
rect 18104 3448 18110 3460
rect 20162 3448 20168 3460
rect 18104 3420 20168 3448
rect 18104 3408 18110 3420
rect 20162 3408 20168 3420
rect 20220 3408 20226 3460
rect 22830 3408 22836 3460
rect 22888 3448 22894 3460
rect 34790 3448 34796 3460
rect 22888 3420 27384 3448
rect 22888 3408 22894 3420
rect 14093 3383 14151 3389
rect 14093 3349 14105 3383
rect 14139 3380 14151 3383
rect 14458 3380 14464 3392
rect 14139 3352 14464 3380
rect 14139 3349 14151 3352
rect 14093 3343 14151 3349
rect 14458 3340 14464 3352
rect 14516 3340 14522 3392
rect 14918 3340 14924 3392
rect 14976 3380 14982 3392
rect 20254 3380 20260 3392
rect 14976 3352 20260 3380
rect 14976 3340 14982 3352
rect 20254 3340 20260 3352
rect 20312 3340 20318 3392
rect 23934 3380 23940 3392
rect 23895 3352 23940 3380
rect 23934 3340 23940 3352
rect 23992 3340 23998 3392
rect 25682 3340 25688 3392
rect 25740 3380 25746 3392
rect 27249 3383 27307 3389
rect 27249 3380 27261 3383
rect 25740 3352 27261 3380
rect 25740 3340 25746 3352
rect 27249 3349 27261 3352
rect 27295 3349 27307 3383
rect 27356 3380 27384 3420
rect 34072 3420 34796 3448
rect 34072 3380 34100 3420
rect 34790 3408 34796 3420
rect 34848 3408 34854 3460
rect 27356 3352 34100 3380
rect 27249 3343 27307 3349
rect 1104 3290 38824 3312
rect 1104 3238 4246 3290
rect 4298 3238 4310 3290
rect 4362 3238 4374 3290
rect 4426 3238 4438 3290
rect 4490 3238 34966 3290
rect 35018 3238 35030 3290
rect 35082 3238 35094 3290
rect 35146 3238 35158 3290
rect 35210 3238 38824 3290
rect 1104 3216 38824 3238
rect 2041 3179 2099 3185
rect 2041 3145 2053 3179
rect 2087 3176 2099 3179
rect 3786 3176 3792 3188
rect 2087 3148 3792 3176
rect 2087 3145 2099 3148
rect 2041 3139 2099 3145
rect 3786 3136 3792 3148
rect 3844 3136 3850 3188
rect 4062 3136 4068 3188
rect 4120 3176 4126 3188
rect 4893 3179 4951 3185
rect 4893 3176 4905 3179
rect 4120 3148 4905 3176
rect 4120 3136 4126 3148
rect 4893 3145 4905 3148
rect 4939 3145 4951 3179
rect 4893 3139 4951 3145
rect 7466 3136 7472 3188
rect 7524 3176 7530 3188
rect 8205 3179 8263 3185
rect 8205 3176 8217 3179
rect 7524 3148 8217 3176
rect 7524 3136 7530 3148
rect 8205 3145 8217 3148
rect 8251 3145 8263 3179
rect 8205 3139 8263 3145
rect 8662 3136 8668 3188
rect 8720 3176 8726 3188
rect 9217 3179 9275 3185
rect 9217 3176 9229 3179
rect 8720 3148 9229 3176
rect 8720 3136 8726 3148
rect 9217 3145 9229 3148
rect 9263 3176 9275 3179
rect 11422 3176 11428 3188
rect 9263 3148 11284 3176
rect 11383 3148 11428 3176
rect 9263 3145 9275 3148
rect 9217 3139 9275 3145
rect 7834 3068 7840 3120
rect 7892 3108 7898 3120
rect 9769 3111 9827 3117
rect 9769 3108 9781 3111
rect 7892 3080 9781 3108
rect 7892 3068 7898 3080
rect 9769 3077 9781 3080
rect 9815 3077 9827 3111
rect 11256 3108 11284 3148
rect 11422 3136 11428 3148
rect 11480 3136 11486 3188
rect 13998 3176 14004 3188
rect 13959 3148 14004 3176
rect 13998 3136 14004 3148
rect 14056 3136 14062 3188
rect 15746 3136 15752 3188
rect 15804 3176 15810 3188
rect 15933 3179 15991 3185
rect 15933 3176 15945 3179
rect 15804 3148 15945 3176
rect 15804 3136 15810 3148
rect 15933 3145 15945 3148
rect 15979 3145 15991 3179
rect 15933 3139 15991 3145
rect 17034 3136 17040 3188
rect 17092 3176 17098 3188
rect 19429 3179 19487 3185
rect 19429 3176 19441 3179
rect 17092 3148 19441 3176
rect 17092 3136 17098 3148
rect 19429 3145 19441 3148
rect 19475 3145 19487 3179
rect 19429 3139 19487 3145
rect 20162 3136 20168 3188
rect 20220 3176 20226 3188
rect 20220 3148 23704 3176
rect 20220 3136 20226 3148
rect 12250 3108 12256 3120
rect 11256 3080 12256 3108
rect 9769 3071 9827 3077
rect 12250 3068 12256 3080
rect 12308 3068 12314 3120
rect 22189 3111 22247 3117
rect 22189 3077 22201 3111
rect 22235 3108 22247 3111
rect 22554 3108 22560 3120
rect 22235 3080 22560 3108
rect 22235 3077 22247 3080
rect 22189 3071 22247 3077
rect 22554 3068 22560 3080
rect 22612 3068 22618 3120
rect 23014 3108 23020 3120
rect 22975 3080 23020 3108
rect 23014 3068 23020 3080
rect 23072 3068 23078 3120
rect 2866 3040 2872 3052
rect 2827 3012 2872 3040
rect 2866 3000 2872 3012
rect 2924 3000 2930 3052
rect 6273 3043 6331 3049
rect 6273 3009 6285 3043
rect 6319 3040 6331 3043
rect 7558 3040 7564 3052
rect 6319 3012 7564 3040
rect 6319 3009 6331 3012
rect 6273 3003 6331 3009
rect 7558 3000 7564 3012
rect 7616 3000 7622 3052
rect 10042 3040 10048 3052
rect 8956 3012 10048 3040
rect 1949 2975 2007 2981
rect 1949 2941 1961 2975
rect 1995 2941 2007 2975
rect 2590 2972 2596 2984
rect 2551 2944 2596 2972
rect 1949 2935 2007 2941
rect 1964 2836 1992 2935
rect 2590 2932 2596 2944
rect 2648 2932 2654 2984
rect 4709 2975 4767 2981
rect 4709 2941 4721 2975
rect 4755 2972 4767 2975
rect 5718 2972 5724 2984
rect 4755 2944 5724 2972
rect 4755 2941 4767 2944
rect 4709 2935 4767 2941
rect 5718 2932 5724 2944
rect 5776 2932 5782 2984
rect 5813 2975 5871 2981
rect 5813 2941 5825 2975
rect 5859 2972 5871 2975
rect 6089 2975 6147 2981
rect 5859 2944 6040 2972
rect 5859 2941 5871 2944
rect 5813 2935 5871 2941
rect 4249 2907 4307 2913
rect 4249 2873 4261 2907
rect 4295 2904 4307 2907
rect 4614 2904 4620 2916
rect 4295 2876 4620 2904
rect 4295 2873 4307 2876
rect 4249 2867 4307 2873
rect 4614 2864 4620 2876
rect 4672 2864 4678 2916
rect 4798 2836 4804 2848
rect 1964 2808 4804 2836
rect 4798 2796 4804 2808
rect 4856 2796 4862 2848
rect 6012 2836 6040 2944
rect 6089 2941 6101 2975
rect 6135 2972 6147 2975
rect 6638 2972 6644 2984
rect 6135 2944 6644 2972
rect 6135 2941 6147 2944
rect 6089 2935 6147 2941
rect 6638 2932 6644 2944
rect 6696 2932 6702 2984
rect 6822 2972 6828 2984
rect 6783 2944 6828 2972
rect 6822 2932 6828 2944
rect 6880 2932 6886 2984
rect 7098 2972 7104 2984
rect 7059 2944 7104 2972
rect 7098 2932 7104 2944
rect 7156 2932 7162 2984
rect 7190 2932 7196 2984
rect 7248 2972 7254 2984
rect 8956 2972 8984 3012
rect 10042 3000 10048 3012
rect 10100 3000 10106 3052
rect 12342 3000 12348 3052
rect 12400 3040 12406 3052
rect 12437 3043 12495 3049
rect 12437 3040 12449 3043
rect 12400 3012 12449 3040
rect 12400 3000 12406 3012
rect 12437 3009 12449 3012
rect 12483 3040 12495 3043
rect 14826 3040 14832 3052
rect 12483 3012 14596 3040
rect 14787 3012 14832 3040
rect 12483 3009 12495 3012
rect 12437 3003 12495 3009
rect 7248 2944 8984 2972
rect 7248 2932 7254 2944
rect 9030 2932 9036 2984
rect 9088 2972 9094 2984
rect 9769 2975 9827 2981
rect 9088 2944 9133 2972
rect 9088 2932 9094 2944
rect 9769 2941 9781 2975
rect 9815 2972 9827 2975
rect 9861 2975 9919 2981
rect 9861 2972 9873 2975
rect 9815 2944 9873 2972
rect 9815 2941 9827 2944
rect 9769 2935 9827 2941
rect 9861 2941 9873 2944
rect 9907 2941 9919 2975
rect 10134 2972 10140 2984
rect 10095 2944 10140 2972
rect 9861 2935 9919 2941
rect 10134 2932 10140 2944
rect 10192 2932 10198 2984
rect 12526 2932 12532 2984
rect 12584 2972 12590 2984
rect 14568 2981 14596 3012
rect 14826 3000 14832 3012
rect 14884 3000 14890 3052
rect 15286 3000 15292 3052
rect 15344 3040 15350 3052
rect 16482 3040 16488 3052
rect 15344 3012 16488 3040
rect 15344 3000 15350 3012
rect 16482 3000 16488 3012
rect 16540 3040 16546 3052
rect 16540 3012 16804 3040
rect 16540 3000 16546 3012
rect 16776 2981 16804 3012
rect 16850 3000 16856 3052
rect 16908 3040 16914 3052
rect 22830 3040 22836 3052
rect 16908 3012 22836 3040
rect 16908 3000 16914 3012
rect 22830 3000 22836 3012
rect 22888 3000 22894 3052
rect 23676 3049 23704 3148
rect 25590 3136 25596 3188
rect 25648 3176 25654 3188
rect 25648 3148 35572 3176
rect 25648 3136 25654 3148
rect 27525 3111 27583 3117
rect 27525 3077 27537 3111
rect 27571 3108 27583 3111
rect 27571 3080 31156 3108
rect 27571 3077 27583 3080
rect 27525 3071 27583 3077
rect 23661 3043 23719 3049
rect 22940 3012 23152 3040
rect 12713 2975 12771 2981
rect 12713 2972 12725 2975
rect 12584 2944 12725 2972
rect 12584 2932 12590 2944
rect 12713 2941 12725 2944
rect 12759 2941 12771 2975
rect 12713 2935 12771 2941
rect 14553 2975 14611 2981
rect 14553 2941 14565 2975
rect 14599 2972 14611 2975
rect 16761 2975 16819 2981
rect 14599 2944 15700 2972
rect 14599 2941 14611 2944
rect 14553 2935 14611 2941
rect 15672 2916 15700 2944
rect 16761 2941 16773 2975
rect 16807 2941 16819 2975
rect 17310 2972 17316 2984
rect 17271 2944 17316 2972
rect 16761 2935 16819 2941
rect 17310 2932 17316 2944
rect 17368 2932 17374 2984
rect 18049 2975 18107 2981
rect 18049 2972 18061 2975
rect 17420 2944 18061 2972
rect 7760 2876 9352 2904
rect 7190 2836 7196 2848
rect 6012 2808 7196 2836
rect 7190 2796 7196 2808
rect 7248 2796 7254 2848
rect 7466 2796 7472 2848
rect 7524 2836 7530 2848
rect 7760 2836 7788 2876
rect 7524 2808 7788 2836
rect 9324 2836 9352 2876
rect 15654 2864 15660 2916
rect 15712 2904 15718 2916
rect 17420 2904 17448 2944
rect 18049 2941 18061 2944
rect 18095 2941 18107 2975
rect 18322 2972 18328 2984
rect 18283 2944 18328 2972
rect 18049 2935 18107 2941
rect 18322 2932 18328 2944
rect 18380 2932 18386 2984
rect 20622 2972 20628 2984
rect 20583 2944 20628 2972
rect 20622 2932 20628 2944
rect 20680 2932 20686 2984
rect 20898 2972 20904 2984
rect 20859 2944 20904 2972
rect 20898 2932 20904 2944
rect 20956 2932 20962 2984
rect 22940 2981 22968 3012
rect 22925 2975 22983 2981
rect 22925 2941 22937 2975
rect 22971 2941 22983 2975
rect 23124 2972 23152 3012
rect 23661 3009 23673 3043
rect 23707 3009 23719 3043
rect 23934 3040 23940 3052
rect 23895 3012 23940 3040
rect 23661 3003 23719 3009
rect 23934 3000 23940 3012
rect 23992 3000 23998 3052
rect 25041 3043 25099 3049
rect 25041 3009 25053 3043
rect 25087 3009 25099 3043
rect 25041 3003 25099 3009
rect 25056 2972 25084 3003
rect 25866 3000 25872 3052
rect 25924 3040 25930 3052
rect 25961 3043 26019 3049
rect 25961 3040 25973 3043
rect 25924 3012 25973 3040
rect 25924 3000 25930 3012
rect 25961 3009 25973 3012
rect 26007 3040 26019 3043
rect 26878 3040 26884 3052
rect 26007 3012 26884 3040
rect 26007 3009 26019 3012
rect 25961 3003 26019 3009
rect 26878 3000 26884 3012
rect 26936 3000 26942 3052
rect 29273 3043 29331 3049
rect 29273 3009 29285 3043
rect 29319 3040 29331 3043
rect 29546 3040 29552 3052
rect 29319 3012 29552 3040
rect 29319 3009 29331 3012
rect 29273 3003 29331 3009
rect 29546 3000 29552 3012
rect 29604 3000 29610 3052
rect 29822 3040 29828 3052
rect 29783 3012 29828 3040
rect 29822 3000 29828 3012
rect 29880 3000 29886 3052
rect 30285 3043 30343 3049
rect 30285 3040 30297 3043
rect 30024 3012 30297 3040
rect 26234 2972 26240 2984
rect 23124 2944 25084 2972
rect 26195 2944 26240 2972
rect 22925 2935 22983 2941
rect 26234 2932 26240 2944
rect 26292 2932 26298 2984
rect 27890 2932 27896 2984
rect 27948 2972 27954 2984
rect 28077 2975 28135 2981
rect 28077 2972 28089 2975
rect 27948 2944 28089 2972
rect 27948 2932 27954 2944
rect 28077 2941 28089 2944
rect 28123 2941 28135 2975
rect 28077 2935 28135 2941
rect 29086 2932 29092 2984
rect 29144 2972 29150 2984
rect 30024 2972 30052 3012
rect 30285 3009 30297 3012
rect 30331 3009 30343 3043
rect 31128 3040 31156 3080
rect 32214 3068 32220 3120
rect 32272 3108 32278 3120
rect 32585 3111 32643 3117
rect 32585 3108 32597 3111
rect 32272 3080 32597 3108
rect 32272 3068 32278 3080
rect 32585 3077 32597 3080
rect 32631 3077 32643 3111
rect 32585 3071 32643 3077
rect 33336 3080 34928 3108
rect 33226 3040 33232 3052
rect 31128 3012 33232 3040
rect 30285 3003 30343 3009
rect 33226 3000 33232 3012
rect 33284 3000 33290 3052
rect 29144 2944 30052 2972
rect 30101 2975 30159 2981
rect 29144 2932 29150 2944
rect 30101 2941 30113 2975
rect 30147 2941 30159 2975
rect 30101 2935 30159 2941
rect 15712 2876 17448 2904
rect 17497 2907 17555 2913
rect 15712 2864 15718 2876
rect 17497 2873 17509 2907
rect 17543 2904 17555 2907
rect 17954 2904 17960 2916
rect 17543 2876 17960 2904
rect 17543 2873 17555 2876
rect 17497 2867 17555 2873
rect 17954 2864 17960 2876
rect 18012 2864 18018 2916
rect 27522 2864 27528 2916
rect 27580 2904 27586 2916
rect 28169 2907 28227 2913
rect 28169 2904 28181 2907
rect 27580 2876 28181 2904
rect 27580 2864 27586 2876
rect 28169 2873 28181 2876
rect 28215 2873 28227 2907
rect 28169 2867 28227 2873
rect 10594 2836 10600 2848
rect 9324 2808 10600 2836
rect 7524 2796 7530 2808
rect 10594 2796 10600 2808
rect 10652 2796 10658 2848
rect 18690 2796 18696 2848
rect 18748 2836 18754 2848
rect 23014 2836 23020 2848
rect 18748 2808 23020 2836
rect 18748 2796 18754 2808
rect 23014 2796 23020 2808
rect 23072 2796 23078 2848
rect 30116 2836 30144 2935
rect 30374 2932 30380 2984
rect 30432 2972 30438 2984
rect 31205 2975 31263 2981
rect 31205 2972 31217 2975
rect 30432 2944 31217 2972
rect 30432 2932 30438 2944
rect 31205 2941 31217 2944
rect 31251 2941 31263 2975
rect 31205 2935 31263 2941
rect 31481 2975 31539 2981
rect 31481 2941 31493 2975
rect 31527 2972 31539 2975
rect 33336 2972 33364 3080
rect 34330 3040 34336 3052
rect 34291 3012 34336 3040
rect 34330 3000 34336 3012
rect 34388 3000 34394 3052
rect 34900 3049 34928 3080
rect 34885 3043 34943 3049
rect 34885 3009 34897 3043
rect 34931 3009 34943 3043
rect 35434 3040 35440 3052
rect 35395 3012 35440 3040
rect 34885 3003 34943 3009
rect 35434 3000 35440 3012
rect 35492 3000 35498 3052
rect 35544 3040 35572 3148
rect 36725 3043 36783 3049
rect 36725 3040 36737 3043
rect 35544 3012 36737 3040
rect 36725 3009 36737 3012
rect 36771 3009 36783 3043
rect 36725 3003 36783 3009
rect 33870 2972 33876 2984
rect 31527 2944 33364 2972
rect 33831 2944 33876 2972
rect 31527 2941 31539 2944
rect 31481 2935 31539 2941
rect 33870 2932 33876 2944
rect 33928 2932 33934 2984
rect 34146 2972 34152 2984
rect 34107 2944 34152 2972
rect 34146 2932 34152 2944
rect 34204 2932 34210 2984
rect 34514 2932 34520 2984
rect 34572 2972 34578 2984
rect 35575 2975 35633 2981
rect 35575 2972 35587 2975
rect 34572 2944 35587 2972
rect 34572 2932 34578 2944
rect 35575 2941 35587 2944
rect 35621 2941 35633 2975
rect 35575 2935 35633 2941
rect 35713 2975 35771 2981
rect 35713 2941 35725 2975
rect 35759 2941 35771 2975
rect 36446 2972 36452 2984
rect 36407 2944 36452 2972
rect 35713 2935 35771 2941
rect 32214 2864 32220 2916
rect 32272 2904 32278 2916
rect 33321 2907 33379 2913
rect 33321 2904 33333 2907
rect 32272 2876 33333 2904
rect 32272 2864 32278 2876
rect 33321 2873 33333 2876
rect 33367 2873 33379 2907
rect 34164 2904 34192 2932
rect 35728 2904 35756 2935
rect 36446 2932 36452 2944
rect 36504 2932 36510 2984
rect 36262 2904 36268 2916
rect 34164 2876 36268 2904
rect 33321 2867 33379 2873
rect 36262 2864 36268 2876
rect 36320 2864 36326 2916
rect 38102 2904 38108 2916
rect 38063 2876 38108 2904
rect 38102 2864 38108 2876
rect 38160 2864 38166 2916
rect 32122 2836 32128 2848
rect 30116 2808 32128 2836
rect 32122 2796 32128 2808
rect 32180 2836 32186 2848
rect 32674 2836 32680 2848
rect 32180 2808 32680 2836
rect 32180 2796 32186 2808
rect 32674 2796 32680 2808
rect 32732 2796 32738 2848
rect 32766 2796 32772 2848
rect 32824 2836 32830 2848
rect 34698 2836 34704 2848
rect 32824 2808 34704 2836
rect 32824 2796 32830 2808
rect 34698 2796 34704 2808
rect 34756 2796 34762 2848
rect 1104 2746 38824 2768
rect 1104 2694 19606 2746
rect 19658 2694 19670 2746
rect 19722 2694 19734 2746
rect 19786 2694 19798 2746
rect 19850 2694 38824 2746
rect 1104 2672 38824 2694
rect 6638 2592 6644 2644
rect 6696 2632 6702 2644
rect 9858 2632 9864 2644
rect 6696 2604 7604 2632
rect 9819 2604 9864 2632
rect 6696 2592 6702 2604
rect 6273 2567 6331 2573
rect 6273 2533 6285 2567
rect 6319 2564 6331 2567
rect 7466 2564 7472 2576
rect 6319 2536 7472 2564
rect 6319 2533 6331 2536
rect 6273 2527 6331 2533
rect 7466 2524 7472 2536
rect 7524 2524 7530 2576
rect 7576 2564 7604 2604
rect 9858 2592 9864 2604
rect 9916 2592 9922 2644
rect 14936 2604 22324 2632
rect 12069 2567 12127 2573
rect 7576 2536 8432 2564
rect 1673 2499 1731 2505
rect 1673 2465 1685 2499
rect 1719 2496 1731 2499
rect 1946 2496 1952 2508
rect 1719 2468 1952 2496
rect 1719 2465 1731 2468
rect 1673 2459 1731 2465
rect 1946 2456 1952 2468
rect 2004 2456 2010 2508
rect 2590 2456 2596 2508
rect 2648 2496 2654 2508
rect 4617 2499 4675 2505
rect 4617 2496 4629 2499
rect 2648 2468 4629 2496
rect 2648 2456 2654 2468
rect 4617 2465 4629 2468
rect 4663 2465 4675 2499
rect 4617 2459 4675 2465
rect 4706 2456 4712 2508
rect 4764 2496 4770 2508
rect 4893 2499 4951 2505
rect 4893 2496 4905 2499
rect 4764 2468 4905 2496
rect 4764 2456 4770 2468
rect 4893 2465 4905 2468
rect 4939 2465 4951 2499
rect 6914 2496 6920 2508
rect 6875 2468 6920 2496
rect 4893 2459 4951 2465
rect 6914 2456 6920 2468
rect 6972 2456 6978 2508
rect 7558 2496 7564 2508
rect 7519 2468 7564 2496
rect 7558 2456 7564 2468
rect 7616 2456 7622 2508
rect 8404 2505 8432 2536
rect 12069 2533 12081 2567
rect 12115 2564 12127 2567
rect 12894 2564 12900 2576
rect 12115 2536 12900 2564
rect 12115 2533 12127 2536
rect 12069 2527 12127 2533
rect 12894 2524 12900 2536
rect 12952 2524 12958 2576
rect 14936 2573 14964 2604
rect 14921 2567 14979 2573
rect 13740 2536 14872 2564
rect 8113 2499 8171 2505
rect 8113 2465 8125 2499
rect 8159 2465 8171 2499
rect 8113 2459 8171 2465
rect 8389 2499 8447 2505
rect 8389 2465 8401 2499
rect 8435 2465 8447 2499
rect 8389 2459 8447 2465
rect 1397 2431 1455 2437
rect 1397 2397 1409 2431
rect 1443 2428 1455 2431
rect 2608 2428 2636 2456
rect 1443 2400 2636 2428
rect 7009 2431 7067 2437
rect 1443 2397 1455 2400
rect 1397 2391 1455 2397
rect 7009 2397 7021 2431
rect 7055 2428 7067 2431
rect 8128 2428 8156 2459
rect 9674 2456 9680 2508
rect 9732 2496 9738 2508
rect 9769 2499 9827 2505
rect 9769 2496 9781 2499
rect 9732 2468 9781 2496
rect 9732 2456 9738 2468
rect 9769 2465 9781 2468
rect 9815 2465 9827 2499
rect 9769 2459 9827 2465
rect 10689 2499 10747 2505
rect 10689 2465 10701 2499
rect 10735 2496 10747 2499
rect 10735 2468 12388 2496
rect 10735 2465 10747 2468
rect 10689 2459 10747 2465
rect 7055 2400 8156 2428
rect 7055 2397 7067 2400
rect 7009 2391 7067 2397
rect 9306 2388 9312 2440
rect 9364 2428 9370 2440
rect 10413 2431 10471 2437
rect 10413 2428 10425 2431
rect 9364 2400 10425 2428
rect 9364 2388 9370 2400
rect 10413 2397 10425 2400
rect 10459 2397 10471 2431
rect 10413 2391 10471 2397
rect 7745 2363 7803 2369
rect 7745 2329 7757 2363
rect 7791 2329 7803 2363
rect 7745 2323 7803 2329
rect 2590 2252 2596 2304
rect 2648 2292 2654 2304
rect 2777 2295 2835 2301
rect 2777 2292 2789 2295
rect 2648 2264 2789 2292
rect 2648 2252 2654 2264
rect 2777 2261 2789 2264
rect 2823 2261 2835 2295
rect 2777 2255 2835 2261
rect 7650 2252 7656 2304
rect 7708 2292 7714 2304
rect 7760 2292 7788 2323
rect 7708 2264 7788 2292
rect 12360 2292 12388 2468
rect 12434 2456 12440 2508
rect 12492 2496 12498 2508
rect 13740 2505 13768 2536
rect 12713 2499 12771 2505
rect 12713 2496 12725 2499
rect 12492 2468 12725 2496
rect 12492 2456 12498 2468
rect 12713 2465 12725 2468
rect 12759 2465 12771 2499
rect 12713 2459 12771 2465
rect 13725 2499 13783 2505
rect 13725 2465 13737 2499
rect 13771 2465 13783 2499
rect 14458 2496 14464 2508
rect 14419 2468 14464 2496
rect 13725 2459 13783 2465
rect 14458 2456 14464 2468
rect 14516 2456 14522 2508
rect 14844 2496 14872 2536
rect 14921 2533 14933 2567
rect 14967 2533 14979 2567
rect 14921 2527 14979 2533
rect 17954 2524 17960 2576
rect 18012 2564 18018 2576
rect 22296 2564 22324 2604
rect 22370 2592 22376 2644
rect 22428 2632 22434 2644
rect 22557 2635 22615 2641
rect 22557 2632 22569 2635
rect 22428 2604 22569 2632
rect 22428 2592 22434 2604
rect 22557 2601 22569 2604
rect 22603 2601 22615 2635
rect 26234 2632 26240 2644
rect 22557 2595 22615 2601
rect 22664 2604 26240 2632
rect 22664 2564 22692 2604
rect 26234 2592 26240 2604
rect 26292 2592 26298 2644
rect 36262 2592 36268 2644
rect 36320 2632 36326 2644
rect 37918 2632 37924 2644
rect 36320 2604 37924 2632
rect 36320 2592 36326 2604
rect 37918 2592 37924 2604
rect 37976 2592 37982 2644
rect 32030 2564 32036 2576
rect 18012 2536 18460 2564
rect 22296 2536 22692 2564
rect 31991 2536 32036 2564
rect 18012 2524 18018 2536
rect 15470 2496 15476 2508
rect 14844 2468 15476 2496
rect 15470 2456 15476 2468
rect 15528 2456 15534 2508
rect 15654 2496 15660 2508
rect 15615 2468 15660 2496
rect 15654 2456 15660 2468
rect 15712 2456 15718 2508
rect 15930 2496 15936 2508
rect 15891 2468 15936 2496
rect 15930 2456 15936 2468
rect 15988 2456 15994 2508
rect 18325 2499 18383 2505
rect 18325 2465 18337 2499
rect 18371 2465 18383 2499
rect 18432 2496 18460 2536
rect 32030 2524 32036 2536
rect 32088 2524 32094 2576
rect 34422 2524 34428 2576
rect 34480 2564 34486 2576
rect 35437 2567 35495 2573
rect 35437 2564 35449 2567
rect 34480 2536 35449 2564
rect 34480 2524 34486 2536
rect 35437 2533 35449 2536
rect 35483 2533 35495 2567
rect 35437 2527 35495 2533
rect 21453 2499 21511 2505
rect 21453 2496 21465 2499
rect 18432 2468 21465 2496
rect 18325 2459 18383 2465
rect 21453 2465 21465 2468
rect 21499 2465 21511 2499
rect 21453 2459 21511 2465
rect 12618 2428 12624 2440
rect 12579 2400 12624 2428
rect 12618 2388 12624 2400
rect 12676 2388 12682 2440
rect 14182 2388 14188 2440
rect 14240 2428 14246 2440
rect 14369 2431 14427 2437
rect 14369 2428 14381 2431
rect 14240 2400 14381 2428
rect 14240 2388 14246 2400
rect 14369 2397 14381 2400
rect 14415 2397 14427 2431
rect 14369 2391 14427 2397
rect 13817 2363 13875 2369
rect 13817 2329 13829 2363
rect 13863 2360 13875 2363
rect 15562 2360 15568 2372
rect 13863 2332 15568 2360
rect 13863 2329 13875 2332
rect 13817 2323 13875 2329
rect 15562 2320 15568 2332
rect 15620 2320 15626 2372
rect 18340 2360 18368 2459
rect 24118 2456 24124 2508
rect 24176 2496 24182 2508
rect 24854 2496 24860 2508
rect 24176 2468 24716 2496
rect 24815 2468 24860 2496
rect 24176 2456 24182 2468
rect 18874 2388 18880 2440
rect 18932 2428 18938 2440
rect 18969 2431 19027 2437
rect 18969 2428 18981 2431
rect 18932 2400 18981 2428
rect 18932 2388 18938 2400
rect 18969 2397 18981 2400
rect 19015 2397 19027 2431
rect 19242 2428 19248 2440
rect 19203 2400 19248 2428
rect 18969 2391 19027 2397
rect 19242 2388 19248 2400
rect 19300 2388 19306 2440
rect 20622 2388 20628 2440
rect 20680 2428 20686 2440
rect 21177 2431 21235 2437
rect 21177 2428 21189 2431
rect 20680 2400 21189 2428
rect 20680 2388 20686 2400
rect 21177 2397 21189 2400
rect 21223 2428 21235 2431
rect 21358 2428 21364 2440
rect 21223 2400 21364 2428
rect 21223 2397 21235 2400
rect 21177 2391 21235 2397
rect 21358 2388 21364 2400
rect 21416 2428 21422 2440
rect 24581 2431 24639 2437
rect 24581 2428 24593 2431
rect 21416 2400 24593 2428
rect 21416 2388 21422 2400
rect 24581 2397 24593 2400
rect 24627 2397 24639 2431
rect 24688 2428 24716 2468
rect 24854 2456 24860 2468
rect 24912 2456 24918 2508
rect 27157 2499 27215 2505
rect 27157 2496 27169 2499
rect 26804 2468 27169 2496
rect 26804 2428 26832 2468
rect 27157 2465 27169 2468
rect 27203 2465 27215 2499
rect 27157 2459 27215 2465
rect 28368 2468 30236 2496
rect 24688 2400 26832 2428
rect 24581 2391 24639 2397
rect 26878 2388 26884 2440
rect 26936 2428 26942 2440
rect 28368 2428 28396 2468
rect 26936 2400 28396 2428
rect 26936 2388 26942 2400
rect 29270 2388 29276 2440
rect 29328 2428 29334 2440
rect 29733 2431 29791 2437
rect 29733 2428 29745 2431
rect 29328 2400 29745 2428
rect 29328 2388 29334 2400
rect 29733 2397 29745 2400
rect 29779 2397 29791 2431
rect 30208 2428 30236 2468
rect 30282 2456 30288 2508
rect 30340 2496 30346 2508
rect 30377 2499 30435 2505
rect 30377 2496 30389 2499
rect 30340 2468 30389 2496
rect 30340 2456 30346 2468
rect 30377 2465 30389 2468
rect 30423 2465 30435 2499
rect 30377 2459 30435 2465
rect 30653 2499 30711 2505
rect 30653 2465 30665 2499
rect 30699 2496 30711 2499
rect 32214 2496 32220 2508
rect 30699 2468 32220 2496
rect 30699 2465 30711 2468
rect 30653 2459 30711 2465
rect 32214 2456 32220 2468
rect 32272 2456 32278 2508
rect 33134 2456 33140 2508
rect 33192 2496 33198 2508
rect 33505 2499 33563 2505
rect 33505 2496 33517 2499
rect 33192 2468 33517 2496
rect 33192 2456 33198 2468
rect 33505 2465 33517 2468
rect 33551 2465 33563 2499
rect 33505 2459 33563 2465
rect 35526 2456 35532 2508
rect 35584 2496 35590 2508
rect 36280 2505 36308 2592
rect 35989 2499 36047 2505
rect 35989 2496 36001 2499
rect 35584 2468 36001 2496
rect 35584 2456 35590 2468
rect 35989 2465 36001 2468
rect 36035 2465 36047 2499
rect 35989 2459 36047 2465
rect 36265 2499 36323 2505
rect 36265 2465 36277 2499
rect 36311 2465 36323 2499
rect 36265 2459 36323 2465
rect 36449 2499 36507 2505
rect 36449 2465 36461 2499
rect 36495 2496 36507 2499
rect 37458 2496 37464 2508
rect 36495 2468 37464 2496
rect 36495 2465 36507 2468
rect 36449 2459 36507 2465
rect 37458 2456 37464 2468
rect 37516 2456 37522 2508
rect 33229 2431 33287 2437
rect 33229 2428 33241 2431
rect 30208 2400 33241 2428
rect 29733 2391 29791 2397
rect 33229 2397 33241 2400
rect 33275 2428 33287 2431
rect 36354 2428 36360 2440
rect 33275 2400 36360 2428
rect 33275 2397 33287 2400
rect 33229 2391 33287 2397
rect 36354 2388 36360 2400
rect 36412 2388 36418 2440
rect 18340 2332 19012 2360
rect 12897 2295 12955 2301
rect 12897 2292 12909 2295
rect 12360 2264 12909 2292
rect 7708 2252 7714 2264
rect 12897 2261 12909 2264
rect 12943 2261 12955 2295
rect 12897 2255 12955 2261
rect 16942 2252 16948 2304
rect 17000 2292 17006 2304
rect 17037 2295 17095 2301
rect 17037 2292 17049 2295
rect 17000 2264 17049 2292
rect 17000 2252 17006 2264
rect 17037 2261 17049 2264
rect 17083 2261 17095 2295
rect 17037 2255 17095 2261
rect 17862 2252 17868 2304
rect 17920 2292 17926 2304
rect 18417 2295 18475 2301
rect 18417 2292 18429 2295
rect 17920 2264 18429 2292
rect 17920 2252 17926 2264
rect 18417 2261 18429 2264
rect 18463 2261 18475 2295
rect 18984 2292 19012 2332
rect 20346 2292 20352 2304
rect 18984 2264 20352 2292
rect 18417 2255 18475 2261
rect 20346 2252 20352 2264
rect 20404 2252 20410 2304
rect 20533 2295 20591 2301
rect 20533 2261 20545 2295
rect 20579 2292 20591 2295
rect 20990 2292 20996 2304
rect 20579 2264 20996 2292
rect 20579 2261 20591 2264
rect 20533 2255 20591 2261
rect 20990 2252 20996 2264
rect 21048 2252 21054 2304
rect 26145 2295 26203 2301
rect 26145 2261 26157 2295
rect 26191 2292 26203 2295
rect 27246 2292 27252 2304
rect 26191 2264 27252 2292
rect 26191 2261 26203 2264
rect 26145 2255 26203 2261
rect 27246 2252 27252 2264
rect 27304 2252 27310 2304
rect 28445 2295 28503 2301
rect 28445 2261 28457 2295
rect 28491 2292 28503 2295
rect 31294 2292 31300 2304
rect 28491 2264 31300 2292
rect 28491 2261 28503 2264
rect 28445 2255 28503 2261
rect 31294 2252 31300 2264
rect 31352 2252 31358 2304
rect 33134 2292 33140 2304
rect 33095 2264 33140 2292
rect 33134 2252 33140 2264
rect 33192 2252 33198 2304
rect 34793 2295 34851 2301
rect 34793 2261 34805 2295
rect 34839 2292 34851 2295
rect 35342 2292 35348 2304
rect 34839 2264 35348 2292
rect 34839 2261 34851 2264
rect 34793 2255 34851 2261
rect 35342 2252 35348 2264
rect 35400 2252 35406 2304
rect 37550 2292 37556 2304
rect 37511 2264 37556 2292
rect 37550 2252 37556 2264
rect 37608 2252 37614 2304
rect 1104 2202 38824 2224
rect 1104 2150 4246 2202
rect 4298 2150 4310 2202
rect 4362 2150 4374 2202
rect 4426 2150 4438 2202
rect 4490 2150 34966 2202
rect 35018 2150 35030 2202
rect 35082 2150 35094 2202
rect 35146 2150 35158 2202
rect 35210 2150 38824 2202
rect 1104 2128 38824 2150
rect 7926 2048 7932 2100
rect 7984 2088 7990 2100
rect 33134 2088 33140 2100
rect 7984 2060 33140 2088
rect 7984 2048 7990 2060
rect 33134 2048 33140 2060
rect 33192 2048 33198 2100
rect 6914 1980 6920 2032
rect 6972 2020 6978 2032
rect 8662 2020 8668 2032
rect 6972 1992 8668 2020
rect 6972 1980 6978 1992
rect 8662 1980 8668 1992
rect 8720 1980 8726 2032
rect 18874 1980 18880 2032
rect 18932 2020 18938 2032
rect 20622 2020 20628 2032
rect 18932 1992 20628 2020
rect 18932 1980 18938 1992
rect 20622 1980 20628 1992
rect 20680 1980 20686 2032
rect 20070 1912 20076 1964
rect 20128 1952 20134 1964
rect 25222 1952 25228 1964
rect 20128 1924 25228 1952
rect 20128 1912 20134 1924
rect 25222 1912 25228 1924
rect 25280 1912 25286 1964
<< via1 >>
rect 21916 39108 21968 39160
rect 23756 39108 23808 39160
rect 19606 37510 19658 37562
rect 19670 37510 19722 37562
rect 19734 37510 19786 37562
rect 19798 37510 19850 37562
rect 5448 37340 5500 37392
rect 9404 37340 9456 37392
rect 4712 37272 4764 37324
rect 6920 37272 6972 37324
rect 7564 37315 7616 37324
rect 7564 37281 7573 37315
rect 7573 37281 7607 37315
rect 7607 37281 7616 37315
rect 7564 37272 7616 37281
rect 7840 37315 7892 37324
rect 7840 37281 7849 37315
rect 7849 37281 7883 37315
rect 7883 37281 7892 37315
rect 7840 37272 7892 37281
rect 7932 37272 7984 37324
rect 9680 37272 9732 37324
rect 9864 37272 9916 37324
rect 11704 37315 11756 37324
rect 11704 37281 11713 37315
rect 11713 37281 11747 37315
rect 11747 37281 11756 37315
rect 11704 37272 11756 37281
rect 21272 37272 21324 37324
rect 24952 37315 25004 37324
rect 24952 37281 24961 37315
rect 24961 37281 24995 37315
rect 24995 37281 25004 37315
rect 24952 37272 25004 37281
rect 5632 37204 5684 37256
rect 15476 37247 15528 37256
rect 15476 37213 15485 37247
rect 15485 37213 15519 37247
rect 15519 37213 15528 37247
rect 15476 37204 15528 37213
rect 15752 37247 15804 37256
rect 15752 37213 15761 37247
rect 15761 37213 15795 37247
rect 15795 37213 15804 37247
rect 15752 37204 15804 37213
rect 1308 37136 1360 37188
rect 7472 37136 7524 37188
rect 9680 37136 9732 37188
rect 4804 37068 4856 37120
rect 5724 37111 5776 37120
rect 5724 37077 5733 37111
rect 5733 37077 5767 37111
rect 5767 37077 5776 37111
rect 5724 37068 5776 37077
rect 9864 37111 9916 37120
rect 9864 37077 9873 37111
rect 9873 37077 9907 37111
rect 9907 37077 9916 37111
rect 9864 37068 9916 37077
rect 12256 37068 12308 37120
rect 32036 37340 32088 37392
rect 36452 37340 36504 37392
rect 29184 37272 29236 37324
rect 33140 37272 33192 37324
rect 35900 37315 35952 37324
rect 29000 37204 29052 37256
rect 30012 37247 30064 37256
rect 30012 37213 30021 37247
rect 30021 37213 30055 37247
rect 30055 37213 30064 37247
rect 30012 37204 30064 37213
rect 33508 37204 33560 37256
rect 35900 37281 35909 37315
rect 35909 37281 35943 37315
rect 35943 37281 35952 37315
rect 35900 37272 35952 37281
rect 35532 37204 35584 37256
rect 37004 37272 37056 37324
rect 37188 37315 37240 37324
rect 37188 37281 37197 37315
rect 37197 37281 37231 37315
rect 37231 37281 37240 37315
rect 37188 37272 37240 37281
rect 16856 37111 16908 37120
rect 16856 37077 16865 37111
rect 16865 37077 16899 37111
rect 16899 37077 16908 37111
rect 16856 37068 16908 37077
rect 26240 37111 26292 37120
rect 26240 37077 26249 37111
rect 26249 37077 26283 37111
rect 26283 37077 26292 37111
rect 26240 37068 26292 37077
rect 36728 37136 36780 37188
rect 37096 37136 37148 37188
rect 31024 37068 31076 37120
rect 37004 37068 37056 37120
rect 4246 36966 4298 37018
rect 4310 36966 4362 37018
rect 4374 36966 4426 37018
rect 4438 36966 4490 37018
rect 34966 36966 35018 37018
rect 35030 36966 35082 37018
rect 35094 36966 35146 37018
rect 35158 36966 35210 37018
rect 2780 36864 2832 36916
rect 2504 36796 2556 36848
rect 6828 36796 6880 36848
rect 7472 36864 7524 36916
rect 7932 36796 7984 36848
rect 13820 36839 13872 36848
rect 13820 36805 13829 36839
rect 13829 36805 13863 36839
rect 13863 36805 13872 36839
rect 13820 36796 13872 36805
rect 15752 36796 15804 36848
rect 2504 36703 2556 36712
rect 2504 36669 2513 36703
rect 2513 36669 2547 36703
rect 2547 36669 2556 36703
rect 2504 36660 2556 36669
rect 3332 36703 3384 36712
rect 3332 36669 3341 36703
rect 3341 36669 3375 36703
rect 3375 36669 3384 36703
rect 3332 36660 3384 36669
rect 3976 36703 4028 36712
rect 3976 36669 3985 36703
rect 3985 36669 4019 36703
rect 4019 36669 4028 36703
rect 3976 36660 4028 36669
rect 5816 36660 5868 36712
rect 5632 36635 5684 36644
rect 5632 36601 5641 36635
rect 5641 36601 5675 36635
rect 5675 36601 5684 36635
rect 7472 36660 7524 36712
rect 8208 36660 8260 36712
rect 9864 36660 9916 36712
rect 11060 36703 11112 36712
rect 11060 36669 11069 36703
rect 11069 36669 11103 36703
rect 11103 36669 11112 36703
rect 11060 36660 11112 36669
rect 11520 36660 11572 36712
rect 12440 36703 12492 36712
rect 12440 36669 12449 36703
rect 12449 36669 12483 36703
rect 12483 36669 12492 36703
rect 12440 36660 12492 36669
rect 12808 36660 12860 36712
rect 16856 36728 16908 36780
rect 15476 36660 15528 36712
rect 15752 36703 15804 36712
rect 15752 36669 15761 36703
rect 15761 36669 15795 36703
rect 15795 36669 15804 36703
rect 15752 36660 15804 36669
rect 23848 36728 23900 36780
rect 18328 36703 18380 36712
rect 5632 36592 5684 36601
rect 18328 36669 18337 36703
rect 18337 36669 18371 36703
rect 18371 36669 18380 36703
rect 18328 36660 18380 36669
rect 20812 36660 20864 36712
rect 21272 36703 21324 36712
rect 21272 36669 21281 36703
rect 21281 36669 21315 36703
rect 21315 36669 21324 36703
rect 21272 36660 21324 36669
rect 21548 36703 21600 36712
rect 21548 36669 21557 36703
rect 21557 36669 21591 36703
rect 21591 36669 21600 36703
rect 21548 36660 21600 36669
rect 23020 36660 23072 36712
rect 23940 36703 23992 36712
rect 23940 36669 23949 36703
rect 23949 36669 23983 36703
rect 23983 36669 23992 36703
rect 23940 36660 23992 36669
rect 26516 36660 26568 36712
rect 27160 36703 27212 36712
rect 27160 36669 27169 36703
rect 27169 36669 27203 36703
rect 27203 36669 27212 36703
rect 27160 36660 27212 36669
rect 30012 36728 30064 36780
rect 30288 36728 30340 36780
rect 37188 36864 37240 36916
rect 35992 36796 36044 36848
rect 37096 36796 37148 36848
rect 30840 36703 30892 36712
rect 1952 36567 2004 36576
rect 1952 36533 1961 36567
rect 1961 36533 1995 36567
rect 1995 36533 2004 36567
rect 1952 36524 2004 36533
rect 6920 36524 6972 36576
rect 10048 36567 10100 36576
rect 10048 36533 10057 36567
rect 10057 36533 10091 36567
rect 10091 36533 10100 36567
rect 10048 36524 10100 36533
rect 11428 36524 11480 36576
rect 11796 36567 11848 36576
rect 11796 36533 11805 36567
rect 11805 36533 11839 36567
rect 11839 36533 11848 36567
rect 11796 36524 11848 36533
rect 17040 36524 17092 36576
rect 18052 36524 18104 36576
rect 23296 36592 23348 36644
rect 28908 36592 28960 36644
rect 30840 36669 30849 36703
rect 30849 36669 30883 36703
rect 30883 36669 30892 36703
rect 30840 36660 30892 36669
rect 30104 36592 30156 36644
rect 36176 36728 36228 36780
rect 37004 36728 37056 36780
rect 32956 36703 33008 36712
rect 32956 36669 32965 36703
rect 32965 36669 32999 36703
rect 32999 36669 33008 36703
rect 32956 36660 33008 36669
rect 35532 36660 35584 36712
rect 35992 36703 36044 36712
rect 35992 36669 36001 36703
rect 36001 36669 36035 36703
rect 36035 36669 36044 36703
rect 35992 36660 36044 36669
rect 35348 36592 35400 36644
rect 36084 36592 36136 36644
rect 19432 36567 19484 36576
rect 19432 36533 19441 36567
rect 19441 36533 19475 36567
rect 19475 36533 19484 36567
rect 19432 36524 19484 36533
rect 20076 36524 20128 36576
rect 25044 36567 25096 36576
rect 25044 36533 25053 36567
rect 25053 36533 25087 36567
rect 25087 36533 25096 36567
rect 25044 36524 25096 36533
rect 29368 36567 29420 36576
rect 29368 36533 29377 36567
rect 29377 36533 29411 36567
rect 29411 36533 29420 36567
rect 29368 36524 29420 36533
rect 35900 36524 35952 36576
rect 19606 36422 19658 36474
rect 19670 36422 19722 36474
rect 19734 36422 19786 36474
rect 19798 36422 19850 36474
rect 3976 36320 4028 36372
rect 7380 36320 7432 36372
rect 2688 36227 2740 36236
rect 2688 36193 2697 36227
rect 2697 36193 2731 36227
rect 2731 36193 2740 36227
rect 2688 36184 2740 36193
rect 4804 36227 4856 36236
rect 2872 36116 2924 36168
rect 3056 36091 3108 36100
rect 3056 36057 3065 36091
rect 3065 36057 3099 36091
rect 3099 36057 3108 36091
rect 3056 36048 3108 36057
rect 3332 36116 3384 36168
rect 4804 36193 4813 36227
rect 4813 36193 4847 36227
rect 4847 36193 4856 36227
rect 4804 36184 4856 36193
rect 10140 36320 10192 36372
rect 21548 36320 21600 36372
rect 23940 36320 23992 36372
rect 27160 36320 27212 36372
rect 8208 36252 8260 36304
rect 8392 36227 8444 36236
rect 8392 36193 8401 36227
rect 8401 36193 8435 36227
rect 8435 36193 8444 36227
rect 8392 36184 8444 36193
rect 10140 36227 10192 36236
rect 4896 36116 4948 36168
rect 6736 36116 6788 36168
rect 9772 36159 9824 36168
rect 9772 36125 9781 36159
rect 9781 36125 9815 36159
rect 9815 36125 9824 36159
rect 9772 36116 9824 36125
rect 10140 36193 10149 36227
rect 10149 36193 10183 36227
rect 10183 36193 10192 36227
rect 10140 36184 10192 36193
rect 10416 36227 10468 36236
rect 10416 36193 10425 36227
rect 10425 36193 10459 36227
rect 10459 36193 10468 36227
rect 10416 36184 10468 36193
rect 11152 36116 11204 36168
rect 6276 36048 6328 36100
rect 10048 36048 10100 36100
rect 18328 36252 18380 36304
rect 12256 36227 12308 36236
rect 12256 36193 12265 36227
rect 12265 36193 12299 36227
rect 12299 36193 12308 36227
rect 12256 36184 12308 36193
rect 13544 36184 13596 36236
rect 15476 36227 15528 36236
rect 15476 36193 15485 36227
rect 15485 36193 15519 36227
rect 15519 36193 15528 36227
rect 15476 36184 15528 36193
rect 15568 36227 15620 36236
rect 15568 36193 15577 36227
rect 15577 36193 15611 36227
rect 15611 36193 15620 36227
rect 15568 36184 15620 36193
rect 15752 36184 15804 36236
rect 18052 36184 18104 36236
rect 19432 36227 19484 36236
rect 19432 36193 19441 36227
rect 19441 36193 19475 36227
rect 19475 36193 19484 36227
rect 19432 36184 19484 36193
rect 20076 36227 20128 36236
rect 20076 36193 20085 36227
rect 20085 36193 20119 36227
rect 20119 36193 20128 36227
rect 20076 36184 20128 36193
rect 20812 36184 20864 36236
rect 23296 36227 23348 36236
rect 23296 36193 23305 36227
rect 23305 36193 23339 36227
rect 23339 36193 23348 36227
rect 23296 36184 23348 36193
rect 26240 36184 26292 36236
rect 28908 36227 28960 36236
rect 28908 36193 28917 36227
rect 28917 36193 28951 36227
rect 28951 36193 28960 36227
rect 28908 36184 28960 36193
rect 12440 36116 12492 36168
rect 14188 36116 14240 36168
rect 17040 36116 17092 36168
rect 19156 36116 19208 36168
rect 23020 36159 23072 36168
rect 23020 36125 23029 36159
rect 23029 36125 23063 36159
rect 23063 36125 23072 36159
rect 23020 36116 23072 36125
rect 26516 36159 26568 36168
rect 26516 36125 26525 36159
rect 26525 36125 26559 36159
rect 26559 36125 26568 36159
rect 26516 36116 26568 36125
rect 29000 36116 29052 36168
rect 8484 36023 8536 36032
rect 8484 35989 8493 36023
rect 8493 35989 8527 36023
rect 8527 35989 8536 36023
rect 8484 35980 8536 35989
rect 9680 35980 9732 36032
rect 13912 35980 13964 36032
rect 14280 35980 14332 36032
rect 15752 36023 15804 36032
rect 15752 35989 15761 36023
rect 15761 35989 15795 36023
rect 15795 35989 15804 36023
rect 15752 35980 15804 35989
rect 32312 36184 32364 36236
rect 32956 36252 33008 36304
rect 33140 36184 33192 36236
rect 34704 36184 34756 36236
rect 35348 36227 35400 36236
rect 33508 36159 33560 36168
rect 33508 36125 33517 36159
rect 33517 36125 33551 36159
rect 33551 36125 33560 36159
rect 33508 36116 33560 36125
rect 35348 36193 35357 36227
rect 35357 36193 35391 36227
rect 35391 36193 35400 36227
rect 35348 36184 35400 36193
rect 35532 36227 35584 36236
rect 35532 36193 35541 36227
rect 35541 36193 35575 36227
rect 35575 36193 35584 36227
rect 35532 36184 35584 36193
rect 35624 36184 35676 36236
rect 36728 36227 36780 36236
rect 36728 36193 36737 36227
rect 36737 36193 36771 36227
rect 36771 36193 36780 36227
rect 36728 36184 36780 36193
rect 35900 36116 35952 36168
rect 36452 36159 36504 36168
rect 36452 36125 36461 36159
rect 36461 36125 36495 36159
rect 36495 36125 36504 36159
rect 36452 36116 36504 36125
rect 33416 36091 33468 36100
rect 33416 36057 33425 36091
rect 33425 36057 33459 36091
rect 33459 36057 33468 36091
rect 33416 36048 33468 36057
rect 34520 36048 34572 36100
rect 30012 36023 30064 36032
rect 30012 35989 30021 36023
rect 30021 35989 30055 36023
rect 30055 35989 30064 36023
rect 30012 35980 30064 35989
rect 30380 35980 30432 36032
rect 37096 35980 37148 36032
rect 4246 35878 4298 35930
rect 4310 35878 4362 35930
rect 4374 35878 4426 35930
rect 4438 35878 4490 35930
rect 34966 35878 35018 35930
rect 35030 35878 35082 35930
rect 35094 35878 35146 35930
rect 35158 35878 35210 35930
rect 20812 35819 20864 35828
rect 20812 35785 20821 35819
rect 20821 35785 20855 35819
rect 20855 35785 20864 35819
rect 20812 35776 20864 35785
rect 21272 35776 21324 35828
rect 24952 35776 25004 35828
rect 3976 35640 4028 35692
rect 2228 35572 2280 35624
rect 5632 35708 5684 35760
rect 23020 35708 23072 35760
rect 5448 35640 5500 35692
rect 6920 35615 6972 35624
rect 5540 35504 5592 35556
rect 6920 35581 6929 35615
rect 6929 35581 6963 35615
rect 6963 35581 6972 35615
rect 6920 35572 6972 35581
rect 8484 35640 8536 35692
rect 10416 35640 10468 35692
rect 11152 35683 11204 35692
rect 11152 35649 11161 35683
rect 11161 35649 11195 35683
rect 11195 35649 11204 35683
rect 11152 35640 11204 35649
rect 15752 35640 15804 35692
rect 6460 35504 6512 35556
rect 9956 35572 10008 35624
rect 10048 35572 10100 35624
rect 10876 35615 10928 35624
rect 10876 35581 10885 35615
rect 10885 35581 10919 35615
rect 10919 35581 10928 35615
rect 10876 35572 10928 35581
rect 11060 35615 11112 35624
rect 11060 35581 11069 35615
rect 11069 35581 11103 35615
rect 11103 35581 11112 35615
rect 11060 35572 11112 35581
rect 11520 35615 11572 35624
rect 11520 35581 11529 35615
rect 11529 35581 11563 35615
rect 11563 35581 11572 35615
rect 11520 35572 11572 35581
rect 9680 35504 9732 35556
rect 12532 35615 12584 35624
rect 12532 35581 12541 35615
rect 12541 35581 12575 35615
rect 12575 35581 12584 35615
rect 12532 35572 12584 35581
rect 13544 35615 13596 35624
rect 13544 35581 13553 35615
rect 13553 35581 13587 35615
rect 13587 35581 13596 35615
rect 13544 35572 13596 35581
rect 14004 35572 14056 35624
rect 15844 35572 15896 35624
rect 16488 35615 16540 35624
rect 16488 35581 16497 35615
rect 16497 35581 16531 35615
rect 16531 35581 16540 35615
rect 16488 35572 16540 35581
rect 17868 35572 17920 35624
rect 19156 35572 19208 35624
rect 19432 35640 19484 35692
rect 21548 35615 21600 35624
rect 21548 35581 21557 35615
rect 21557 35581 21591 35615
rect 21591 35581 21600 35615
rect 21548 35572 21600 35581
rect 25044 35640 25096 35692
rect 27988 35776 28040 35828
rect 29000 35776 29052 35828
rect 29920 35776 29972 35828
rect 38292 35776 38344 35828
rect 26516 35640 26568 35692
rect 28908 35640 28960 35692
rect 30012 35640 30064 35692
rect 34244 35708 34296 35760
rect 34704 35708 34756 35760
rect 26332 35615 26384 35624
rect 13820 35547 13872 35556
rect 13820 35513 13829 35547
rect 13829 35513 13863 35547
rect 13863 35513 13872 35547
rect 13820 35504 13872 35513
rect 16120 35504 16172 35556
rect 18972 35504 19024 35556
rect 20812 35504 20864 35556
rect 4712 35436 4764 35488
rect 5264 35436 5316 35488
rect 5356 35436 5408 35488
rect 7748 35436 7800 35488
rect 8024 35479 8076 35488
rect 8024 35445 8033 35479
rect 8033 35445 8067 35479
rect 8067 35445 8076 35479
rect 8024 35436 8076 35445
rect 13360 35436 13412 35488
rect 26332 35581 26341 35615
rect 26341 35581 26375 35615
rect 26375 35581 26384 35615
rect 26332 35572 26384 35581
rect 29092 35615 29144 35624
rect 29092 35581 29101 35615
rect 29101 35581 29135 35615
rect 29135 35581 29144 35615
rect 29092 35572 29144 35581
rect 22652 35547 22704 35556
rect 22652 35513 22661 35547
rect 22661 35513 22695 35547
rect 22695 35513 22704 35547
rect 22652 35504 22704 35513
rect 30288 35572 30340 35624
rect 30656 35479 30708 35488
rect 30656 35445 30665 35479
rect 30665 35445 30699 35479
rect 30699 35445 30708 35479
rect 30656 35436 30708 35445
rect 31116 35436 31168 35488
rect 33784 35572 33836 35624
rect 35992 35640 36044 35692
rect 37096 35640 37148 35692
rect 34152 35615 34204 35624
rect 34152 35581 34161 35615
rect 34161 35581 34195 35615
rect 34195 35581 34204 35615
rect 34152 35572 34204 35581
rect 35624 35615 35676 35624
rect 35624 35581 35633 35615
rect 35633 35581 35667 35615
rect 35667 35581 35676 35615
rect 35624 35572 35676 35581
rect 35808 35436 35860 35488
rect 19606 35334 19658 35386
rect 19670 35334 19722 35386
rect 19734 35334 19786 35386
rect 19798 35334 19850 35386
rect 2228 35275 2280 35284
rect 2228 35241 2237 35275
rect 2237 35241 2271 35275
rect 2271 35241 2280 35275
rect 2228 35232 2280 35241
rect 3424 35232 3476 35284
rect 3056 35164 3108 35216
rect 5264 35164 5316 35216
rect 8392 35232 8444 35284
rect 2872 35139 2924 35148
rect 2872 35105 2881 35139
rect 2881 35105 2915 35139
rect 2915 35105 2924 35139
rect 2872 35096 2924 35105
rect 2688 35028 2740 35080
rect 4712 35096 4764 35148
rect 5448 35096 5500 35148
rect 5632 35096 5684 35148
rect 6460 35139 6512 35148
rect 6460 35105 6469 35139
rect 6469 35105 6503 35139
rect 6503 35105 6512 35139
rect 6460 35096 6512 35105
rect 1676 34892 1728 34944
rect 2688 34892 2740 34944
rect 4712 34960 4764 35012
rect 4896 35003 4948 35012
rect 4896 34969 4905 35003
rect 4905 34969 4939 35003
rect 4939 34969 4948 35003
rect 4896 34960 4948 34969
rect 3792 34892 3844 34944
rect 7012 35028 7064 35080
rect 10048 35164 10100 35216
rect 7380 35096 7432 35148
rect 9680 35139 9732 35148
rect 9680 35105 9689 35139
rect 9689 35105 9723 35139
rect 9723 35105 9732 35139
rect 9680 35096 9732 35105
rect 7564 35071 7616 35080
rect 7564 35037 7573 35071
rect 7573 35037 7607 35071
rect 7607 35037 7616 35071
rect 7564 35028 7616 35037
rect 7748 35028 7800 35080
rect 16488 35232 16540 35284
rect 10232 35164 10284 35216
rect 10876 35164 10928 35216
rect 10324 35096 10376 35148
rect 10784 35096 10836 35148
rect 11428 35139 11480 35148
rect 11428 35105 11437 35139
rect 11437 35105 11471 35139
rect 11471 35105 11480 35139
rect 11428 35096 11480 35105
rect 11520 35096 11572 35148
rect 12624 35096 12676 35148
rect 13360 35164 13412 35216
rect 11704 35071 11756 35080
rect 11704 35037 11713 35071
rect 11713 35037 11747 35071
rect 11747 35037 11756 35071
rect 11704 35028 11756 35037
rect 9680 34960 9732 35012
rect 11888 34960 11940 35012
rect 13544 34960 13596 35012
rect 8300 34892 8352 34944
rect 9864 34935 9916 34944
rect 9864 34901 9873 34935
rect 9873 34901 9907 34935
rect 9907 34901 9916 34935
rect 9864 34892 9916 34901
rect 9956 34892 10008 34944
rect 15568 35164 15620 35216
rect 13820 35139 13872 35148
rect 13820 35105 13829 35139
rect 13829 35105 13863 35139
rect 13863 35105 13872 35139
rect 13820 35096 13872 35105
rect 14188 35139 14240 35148
rect 14188 35105 14197 35139
rect 14197 35105 14231 35139
rect 14231 35105 14240 35139
rect 14188 35096 14240 35105
rect 17132 35096 17184 35148
rect 18880 35232 18932 35284
rect 19156 35232 19208 35284
rect 17592 35096 17644 35148
rect 21548 35232 21600 35284
rect 20996 35139 21048 35148
rect 20996 35105 21005 35139
rect 21005 35105 21039 35139
rect 21039 35105 21048 35139
rect 20996 35096 21048 35105
rect 22652 35139 22704 35148
rect 22652 35105 22661 35139
rect 22661 35105 22695 35139
rect 22695 35105 22704 35139
rect 22652 35096 22704 35105
rect 24768 35096 24820 35148
rect 15568 35028 15620 35080
rect 15844 35071 15896 35080
rect 15844 35037 15853 35071
rect 15853 35037 15887 35071
rect 15887 35037 15896 35071
rect 15844 35028 15896 35037
rect 16488 35028 16540 35080
rect 20812 35028 20864 35080
rect 22376 35071 22428 35080
rect 22376 35037 22385 35071
rect 22385 35037 22419 35071
rect 22419 35037 22428 35071
rect 22376 35028 22428 35037
rect 23388 35028 23440 35080
rect 26516 35071 26568 35080
rect 26516 35037 26525 35071
rect 26525 35037 26559 35071
rect 26559 35037 26568 35071
rect 26516 35028 26568 35037
rect 29092 35232 29144 35284
rect 33784 35275 33836 35284
rect 30656 35164 30708 35216
rect 29368 35139 29420 35148
rect 29368 35105 29377 35139
rect 29377 35105 29411 35139
rect 29411 35105 29420 35139
rect 29368 35096 29420 35105
rect 30104 35096 30156 35148
rect 30380 35096 30432 35148
rect 33784 35241 33793 35275
rect 33793 35241 33827 35275
rect 33827 35241 33836 35275
rect 33784 35232 33836 35241
rect 31024 35164 31076 35216
rect 31024 35071 31076 35080
rect 31024 35037 31033 35071
rect 31033 35037 31067 35071
rect 31067 35037 31076 35071
rect 31024 35028 31076 35037
rect 31852 35028 31904 35080
rect 32220 35071 32272 35080
rect 32220 35037 32229 35071
rect 32229 35037 32263 35071
rect 32263 35037 32272 35071
rect 32220 35028 32272 35037
rect 33416 35096 33468 35148
rect 34152 35164 34204 35216
rect 35900 35232 35952 35284
rect 35532 35164 35584 35216
rect 35808 35164 35860 35216
rect 36084 35139 36136 35148
rect 36084 35105 36093 35139
rect 36093 35105 36127 35139
rect 36127 35105 36136 35139
rect 36084 35096 36136 35105
rect 19064 34892 19116 34944
rect 21180 34935 21232 34944
rect 21180 34901 21189 34935
rect 21189 34901 21223 34935
rect 21223 34901 21232 34935
rect 21180 34892 21232 34901
rect 24400 34892 24452 34944
rect 25964 34892 26016 34944
rect 30748 35003 30800 35012
rect 30748 34969 30757 35003
rect 30757 34969 30791 35003
rect 30791 34969 30800 35003
rect 36912 35028 36964 35080
rect 30748 34960 30800 34969
rect 35256 34960 35308 35012
rect 27528 34892 27580 34944
rect 35440 34935 35492 34944
rect 35440 34901 35449 34935
rect 35449 34901 35483 34935
rect 35483 34901 35492 34935
rect 35440 34892 35492 34901
rect 4246 34790 4298 34842
rect 4310 34790 4362 34842
rect 4374 34790 4426 34842
rect 4438 34790 4490 34842
rect 34966 34790 35018 34842
rect 35030 34790 35082 34842
rect 35094 34790 35146 34842
rect 35158 34790 35210 34842
rect 2228 34688 2280 34740
rect 6920 34688 6972 34740
rect 4160 34552 4212 34604
rect 2228 34484 2280 34536
rect 2688 34527 2740 34536
rect 2688 34493 2697 34527
rect 2697 34493 2731 34527
rect 2731 34493 2740 34527
rect 2688 34484 2740 34493
rect 3240 34527 3292 34536
rect 3240 34493 3249 34527
rect 3249 34493 3283 34527
rect 3283 34493 3292 34527
rect 3240 34484 3292 34493
rect 3608 34527 3660 34536
rect 3608 34493 3617 34527
rect 3617 34493 3651 34527
rect 3651 34493 3660 34527
rect 3608 34484 3660 34493
rect 3792 34527 3844 34536
rect 3792 34493 3801 34527
rect 3801 34493 3835 34527
rect 3835 34493 3844 34527
rect 3792 34484 3844 34493
rect 4620 34484 4672 34536
rect 5540 34620 5592 34672
rect 8576 34620 8628 34672
rect 1584 34459 1636 34468
rect 1584 34425 1593 34459
rect 1593 34425 1627 34459
rect 1627 34425 1636 34459
rect 1584 34416 1636 34425
rect 5632 34527 5684 34536
rect 5632 34493 5641 34527
rect 5641 34493 5675 34527
rect 5675 34493 5684 34527
rect 5632 34484 5684 34493
rect 5724 34484 5776 34536
rect 6828 34552 6880 34604
rect 7932 34595 7984 34604
rect 7932 34561 7941 34595
rect 7941 34561 7975 34595
rect 7975 34561 7984 34595
rect 7932 34552 7984 34561
rect 10784 34620 10836 34672
rect 10324 34595 10376 34604
rect 10324 34561 10333 34595
rect 10333 34561 10367 34595
rect 10367 34561 10376 34595
rect 10324 34552 10376 34561
rect 7288 34527 7340 34536
rect 7288 34493 7297 34527
rect 7297 34493 7331 34527
rect 7331 34493 7340 34527
rect 7288 34484 7340 34493
rect 6000 34416 6052 34468
rect 7012 34416 7064 34468
rect 9864 34484 9916 34536
rect 11520 34552 11572 34604
rect 17592 34688 17644 34740
rect 10784 34527 10836 34536
rect 10784 34493 10793 34527
rect 10793 34493 10827 34527
rect 10827 34493 10836 34527
rect 10784 34484 10836 34493
rect 11888 34484 11940 34536
rect 11152 34416 11204 34468
rect 16856 34620 16908 34672
rect 14280 34552 14332 34604
rect 15016 34552 15068 34604
rect 16120 34595 16172 34604
rect 16120 34561 16129 34595
rect 16129 34561 16163 34595
rect 16163 34561 16172 34595
rect 16120 34552 16172 34561
rect 17684 34552 17736 34604
rect 19248 34552 19300 34604
rect 12532 34484 12584 34536
rect 13360 34484 13412 34536
rect 13820 34527 13872 34536
rect 13820 34493 13829 34527
rect 13829 34493 13863 34527
rect 13863 34493 13872 34527
rect 13820 34484 13872 34493
rect 14004 34527 14056 34536
rect 14004 34493 14013 34527
rect 14013 34493 14047 34527
rect 14047 34493 14056 34527
rect 14004 34484 14056 34493
rect 14188 34527 14240 34536
rect 14188 34493 14197 34527
rect 14197 34493 14231 34527
rect 14231 34493 14240 34527
rect 14188 34484 14240 34493
rect 14464 34527 14516 34536
rect 14464 34493 14473 34527
rect 14473 34493 14507 34527
rect 14507 34493 14516 34527
rect 14464 34484 14516 34493
rect 18052 34527 18104 34536
rect 18052 34493 18061 34527
rect 18061 34493 18095 34527
rect 18095 34493 18104 34527
rect 18052 34484 18104 34493
rect 18144 34484 18196 34536
rect 18696 34416 18748 34468
rect 21180 34552 21232 34604
rect 32312 34688 32364 34740
rect 33140 34688 33192 34740
rect 36360 34688 36412 34740
rect 22376 34552 22428 34604
rect 24400 34595 24452 34604
rect 24400 34561 24409 34595
rect 24409 34561 24443 34595
rect 24443 34561 24452 34595
rect 24400 34552 24452 34561
rect 25504 34595 25556 34604
rect 25504 34561 25513 34595
rect 25513 34561 25547 34595
rect 25547 34561 25556 34595
rect 25504 34552 25556 34561
rect 27528 34552 27580 34604
rect 21364 34484 21416 34536
rect 21732 34527 21784 34536
rect 21732 34493 21741 34527
rect 21741 34493 21775 34527
rect 21775 34493 21784 34527
rect 21732 34484 21784 34493
rect 23848 34484 23900 34536
rect 24216 34484 24268 34536
rect 26516 34484 26568 34536
rect 28908 34484 28960 34536
rect 29552 34527 29604 34536
rect 29552 34493 29561 34527
rect 29561 34493 29595 34527
rect 29595 34493 29604 34527
rect 29552 34484 29604 34493
rect 31392 34527 31444 34536
rect 31392 34493 31401 34527
rect 31401 34493 31435 34527
rect 31435 34493 31444 34527
rect 31392 34484 31444 34493
rect 31668 34527 31720 34536
rect 31668 34493 31677 34527
rect 31677 34493 31711 34527
rect 31711 34493 31720 34527
rect 31668 34484 31720 34493
rect 33508 34484 33560 34536
rect 35808 34620 35860 34672
rect 34520 34552 34572 34604
rect 37280 34595 37332 34604
rect 37280 34561 37289 34595
rect 37289 34561 37323 34595
rect 37323 34561 37332 34595
rect 37280 34552 37332 34561
rect 35440 34484 35492 34536
rect 37188 34484 37240 34536
rect 7656 34348 7708 34400
rect 11060 34391 11112 34400
rect 11060 34357 11069 34391
rect 11069 34357 11103 34391
rect 11103 34357 11112 34391
rect 11060 34348 11112 34357
rect 28448 34391 28500 34400
rect 28448 34357 28457 34391
rect 28457 34357 28491 34391
rect 28491 34357 28500 34391
rect 28448 34348 28500 34357
rect 30656 34391 30708 34400
rect 30656 34357 30665 34391
rect 30665 34357 30699 34391
rect 30699 34357 30708 34391
rect 30656 34348 30708 34357
rect 19606 34246 19658 34298
rect 19670 34246 19722 34298
rect 19734 34246 19786 34298
rect 19798 34246 19850 34298
rect 2688 34144 2740 34196
rect 6000 34187 6052 34196
rect 6000 34153 6009 34187
rect 6009 34153 6043 34187
rect 6043 34153 6052 34187
rect 6000 34144 6052 34153
rect 4160 34008 4212 34060
rect 8576 34144 8628 34196
rect 11244 34144 11296 34196
rect 12624 34144 12676 34196
rect 14464 34144 14516 34196
rect 29552 34187 29604 34196
rect 29552 34153 29561 34187
rect 29561 34153 29595 34187
rect 29595 34153 29604 34187
rect 29552 34144 29604 34153
rect 7012 34076 7064 34128
rect 7288 34051 7340 34060
rect 7288 34017 7297 34051
rect 7297 34017 7331 34051
rect 7331 34017 7340 34051
rect 7288 34008 7340 34017
rect 9772 34076 9824 34128
rect 7932 34008 7984 34060
rect 8392 34008 8444 34060
rect 8760 34008 8812 34060
rect 10140 34076 10192 34128
rect 10876 34076 10928 34128
rect 11060 34051 11112 34060
rect 11060 34017 11069 34051
rect 11069 34017 11103 34051
rect 11103 34017 11112 34051
rect 11060 34008 11112 34017
rect 11520 34051 11572 34060
rect 11520 34017 11529 34051
rect 11529 34017 11563 34051
rect 11563 34017 11572 34051
rect 11520 34008 11572 34017
rect 11796 34051 11848 34060
rect 11796 34017 11805 34051
rect 11805 34017 11839 34051
rect 11839 34017 11848 34051
rect 11796 34008 11848 34017
rect 20996 34076 21048 34128
rect 21732 34119 21784 34128
rect 21732 34085 21741 34119
rect 21741 34085 21775 34119
rect 21775 34085 21784 34119
rect 21732 34076 21784 34085
rect 1400 33983 1452 33992
rect 1400 33949 1409 33983
rect 1409 33949 1443 33983
rect 1443 33949 1452 33983
rect 1400 33940 1452 33949
rect 1860 33940 1912 33992
rect 3976 33940 4028 33992
rect 5080 33940 5132 33992
rect 6920 33983 6972 33992
rect 6920 33949 6929 33983
rect 6929 33949 6963 33983
rect 6963 33949 6972 33983
rect 6920 33940 6972 33949
rect 8300 33940 8352 33992
rect 13360 34008 13412 34060
rect 16856 34008 16908 34060
rect 18696 34051 18748 34060
rect 18696 34017 18705 34051
rect 18705 34017 18739 34051
rect 18739 34017 18748 34051
rect 18696 34008 18748 34017
rect 18972 34051 19024 34060
rect 18972 34017 18981 34051
rect 18981 34017 19015 34051
rect 19015 34017 19024 34051
rect 18972 34008 19024 34017
rect 19248 34008 19300 34060
rect 13268 33983 13320 33992
rect 12440 33872 12492 33924
rect 13268 33949 13277 33983
rect 13277 33949 13311 33983
rect 13311 33949 13320 33983
rect 13268 33940 13320 33949
rect 15292 33940 15344 33992
rect 16396 33940 16448 33992
rect 23388 34008 23440 34060
rect 28448 34051 28500 34060
rect 28448 34017 28457 34051
rect 28457 34017 28491 34051
rect 28491 34017 28500 34051
rect 28448 34008 28500 34017
rect 29276 34008 29328 34060
rect 31668 34076 31720 34128
rect 31944 34008 31996 34060
rect 32220 34144 32272 34196
rect 36452 34144 36504 34196
rect 33048 34008 33100 34060
rect 35532 34008 35584 34060
rect 37004 34051 37056 34060
rect 37004 34017 37013 34051
rect 37013 34017 37047 34051
rect 37047 34017 37056 34051
rect 37004 34008 37056 34017
rect 17592 33804 17644 33856
rect 18420 33804 18472 33856
rect 21640 33804 21692 33856
rect 23940 33940 23992 33992
rect 24216 33940 24268 33992
rect 24952 33940 25004 33992
rect 22376 33804 22428 33856
rect 24216 33804 24268 33856
rect 24676 33804 24728 33856
rect 25872 33847 25924 33856
rect 25872 33813 25881 33847
rect 25881 33813 25915 33847
rect 25915 33813 25924 33847
rect 25872 33804 25924 33813
rect 25964 33804 26016 33856
rect 28908 33940 28960 33992
rect 31024 33983 31076 33992
rect 31024 33949 31033 33983
rect 31033 33949 31067 33983
rect 31067 33949 31076 33983
rect 31024 33940 31076 33949
rect 33692 33940 33744 33992
rect 36176 33983 36228 33992
rect 36176 33949 36185 33983
rect 36185 33949 36219 33983
rect 36219 33949 36228 33983
rect 36176 33940 36228 33949
rect 36636 33940 36688 33992
rect 37188 33983 37240 33992
rect 37188 33949 37197 33983
rect 37197 33949 37231 33983
rect 37231 33949 37240 33983
rect 37188 33940 37240 33949
rect 29092 33804 29144 33856
rect 30472 33847 30524 33856
rect 30472 33813 30481 33847
rect 30481 33813 30515 33847
rect 30515 33813 30524 33847
rect 30472 33804 30524 33813
rect 35348 33804 35400 33856
rect 4246 33702 4298 33754
rect 4310 33702 4362 33754
rect 4374 33702 4426 33754
rect 4438 33702 4490 33754
rect 34966 33702 35018 33754
rect 35030 33702 35082 33754
rect 35094 33702 35146 33754
rect 35158 33702 35210 33754
rect 1860 33643 1912 33652
rect 1860 33609 1869 33643
rect 1869 33609 1903 33643
rect 1903 33609 1912 33643
rect 1860 33600 1912 33609
rect 4620 33600 4672 33652
rect 1400 33464 1452 33516
rect 3976 33464 4028 33516
rect 1492 33439 1544 33448
rect 1492 33405 1501 33439
rect 1501 33405 1535 33439
rect 1535 33405 1544 33439
rect 1492 33396 1544 33405
rect 1676 33439 1728 33448
rect 1676 33405 1685 33439
rect 1685 33405 1719 33439
rect 1719 33405 1728 33439
rect 1676 33396 1728 33405
rect 4160 33396 4212 33448
rect 1584 33371 1636 33380
rect 1584 33337 1593 33371
rect 1593 33337 1627 33371
rect 1627 33337 1636 33371
rect 1584 33328 1636 33337
rect 6092 33532 6144 33584
rect 7012 33600 7064 33652
rect 9680 33600 9732 33652
rect 13268 33600 13320 33652
rect 16396 33600 16448 33652
rect 16580 33600 16632 33652
rect 18052 33600 18104 33652
rect 22376 33600 22428 33652
rect 23940 33643 23992 33652
rect 23940 33609 23949 33643
rect 23949 33609 23983 33643
rect 23983 33609 23992 33643
rect 23940 33600 23992 33609
rect 24952 33643 25004 33652
rect 24952 33609 24961 33643
rect 24961 33609 24995 33643
rect 24995 33609 25004 33643
rect 24952 33600 25004 33609
rect 33048 33600 33100 33652
rect 37188 33600 37240 33652
rect 7564 33575 7616 33584
rect 7564 33541 7573 33575
rect 7573 33541 7607 33575
rect 7607 33541 7616 33575
rect 7564 33532 7616 33541
rect 7932 33532 7984 33584
rect 4620 33396 4672 33448
rect 6644 33464 6696 33516
rect 5724 33439 5776 33448
rect 5724 33405 5733 33439
rect 5733 33405 5767 33439
rect 5767 33405 5776 33439
rect 5724 33396 5776 33405
rect 5540 33371 5592 33380
rect 5540 33337 5549 33371
rect 5549 33337 5583 33371
rect 5583 33337 5592 33371
rect 5540 33328 5592 33337
rect 6920 33396 6972 33448
rect 7472 33439 7524 33448
rect 7472 33405 7481 33439
rect 7481 33405 7515 33439
rect 7515 33405 7524 33439
rect 7472 33396 7524 33405
rect 7656 33439 7708 33448
rect 7656 33405 7665 33439
rect 7665 33405 7699 33439
rect 7699 33405 7708 33439
rect 7656 33396 7708 33405
rect 7932 33396 7984 33448
rect 8760 33396 8812 33448
rect 9128 33439 9180 33448
rect 8668 33328 8720 33380
rect 4620 33260 4672 33312
rect 7288 33260 7340 33312
rect 8484 33260 8536 33312
rect 9128 33405 9137 33439
rect 9137 33405 9171 33439
rect 9171 33405 9180 33439
rect 9128 33396 9180 33405
rect 9772 33439 9824 33448
rect 9772 33405 9781 33439
rect 9781 33405 9815 33439
rect 9815 33405 9824 33439
rect 9772 33396 9824 33405
rect 11244 33439 11296 33448
rect 11244 33405 11253 33439
rect 11253 33405 11287 33439
rect 11287 33405 11296 33439
rect 11244 33396 11296 33405
rect 12624 33464 12676 33516
rect 12992 33439 13044 33448
rect 12992 33405 13001 33439
rect 13001 33405 13035 33439
rect 13035 33405 13044 33439
rect 12992 33396 13044 33405
rect 13360 33439 13412 33448
rect 13360 33405 13369 33439
rect 13369 33405 13403 33439
rect 13403 33405 13412 33439
rect 13360 33396 13412 33405
rect 14004 33396 14056 33448
rect 14188 33439 14240 33448
rect 14188 33405 14197 33439
rect 14197 33405 14231 33439
rect 14231 33405 14240 33439
rect 14188 33396 14240 33405
rect 16396 33464 16448 33516
rect 11244 33260 11296 33312
rect 17132 33439 17184 33448
rect 17132 33405 17141 33439
rect 17141 33405 17175 33439
rect 17175 33405 17184 33439
rect 17132 33396 17184 33405
rect 18420 33439 18472 33448
rect 18420 33405 18429 33439
rect 18429 33405 18463 33439
rect 18463 33405 18472 33439
rect 18420 33396 18472 33405
rect 19340 33439 19392 33448
rect 17224 33328 17276 33380
rect 19340 33405 19349 33439
rect 19349 33405 19383 33439
rect 19383 33405 19392 33439
rect 19340 33396 19392 33405
rect 19432 33396 19484 33448
rect 23020 33464 23072 33516
rect 23848 33464 23900 33516
rect 20352 33439 20404 33448
rect 20352 33405 20361 33439
rect 20361 33405 20395 33439
rect 20395 33405 20404 33439
rect 20352 33396 20404 33405
rect 19984 33328 20036 33380
rect 20076 33260 20128 33312
rect 20628 33260 20680 33312
rect 22652 33396 22704 33448
rect 23388 33396 23440 33448
rect 23756 33439 23808 33448
rect 23756 33405 23765 33439
rect 23765 33405 23799 33439
rect 23799 33405 23808 33439
rect 24676 33439 24728 33448
rect 23756 33396 23808 33405
rect 24676 33405 24685 33439
rect 24685 33405 24719 33439
rect 24719 33405 24728 33439
rect 24676 33396 24728 33405
rect 30656 33464 30708 33516
rect 31852 33464 31904 33516
rect 36636 33464 36688 33516
rect 25780 33439 25832 33448
rect 25780 33405 25789 33439
rect 25789 33405 25823 33439
rect 25823 33405 25832 33439
rect 25780 33396 25832 33405
rect 23020 33328 23072 33380
rect 23388 33260 23440 33312
rect 27160 33303 27212 33312
rect 27160 33269 27169 33303
rect 27169 33269 27203 33303
rect 27203 33269 27212 33303
rect 27160 33260 27212 33269
rect 28356 33439 28408 33448
rect 28356 33405 28365 33439
rect 28365 33405 28399 33439
rect 28399 33405 28408 33439
rect 28356 33396 28408 33405
rect 28540 33439 28592 33448
rect 28540 33405 28549 33439
rect 28549 33405 28583 33439
rect 28583 33405 28592 33439
rect 28540 33396 28592 33405
rect 28908 33396 28960 33448
rect 30748 33396 30800 33448
rect 31392 33396 31444 33448
rect 35532 33439 35584 33448
rect 35532 33405 35541 33439
rect 35541 33405 35575 33439
rect 35575 33405 35584 33439
rect 35532 33396 35584 33405
rect 36452 33439 36504 33448
rect 29368 33328 29420 33380
rect 36452 33405 36461 33439
rect 36461 33405 36495 33439
rect 36495 33405 36504 33439
rect 36452 33396 36504 33405
rect 36728 33439 36780 33448
rect 36728 33405 36737 33439
rect 36737 33405 36771 33439
rect 36771 33405 36780 33439
rect 36728 33396 36780 33405
rect 36268 33260 36320 33312
rect 19606 33158 19658 33210
rect 19670 33158 19722 33210
rect 19734 33158 19786 33210
rect 19798 33158 19850 33210
rect 5632 33099 5684 33108
rect 5632 33065 5641 33099
rect 5641 33065 5675 33099
rect 5675 33065 5684 33099
rect 5632 33056 5684 33065
rect 6368 33056 6420 33108
rect 11244 33099 11296 33108
rect 1492 32988 1544 33040
rect 4160 32988 4212 33040
rect 4712 32988 4764 33040
rect 2596 32963 2648 32972
rect 2596 32929 2605 32963
rect 2605 32929 2639 32963
rect 2639 32929 2648 32963
rect 2596 32920 2648 32929
rect 2780 32963 2832 32972
rect 2780 32929 2789 32963
rect 2789 32929 2823 32963
rect 2823 32929 2832 32963
rect 2964 32963 3016 32972
rect 2780 32920 2832 32929
rect 2964 32929 2973 32963
rect 2973 32929 3007 32963
rect 3007 32929 3016 32963
rect 2964 32920 3016 32929
rect 3148 32963 3200 32972
rect 3148 32929 3157 32963
rect 3157 32929 3191 32963
rect 3191 32929 3200 32963
rect 3148 32920 3200 32929
rect 3240 32920 3292 32972
rect 3608 32920 3660 32972
rect 6276 32920 6328 32972
rect 8484 32988 8536 33040
rect 11244 33065 11253 33099
rect 11253 33065 11287 33099
rect 11287 33065 11296 33099
rect 11244 33056 11296 33065
rect 12992 33056 13044 33108
rect 15292 33056 15344 33108
rect 11336 32988 11388 33040
rect 14004 32988 14056 33040
rect 8392 32963 8444 32972
rect 8392 32929 8401 32963
rect 8401 32929 8435 32963
rect 8435 32929 8444 32963
rect 8392 32920 8444 32929
rect 8576 32963 8628 32972
rect 8576 32929 8585 32963
rect 8585 32929 8619 32963
rect 8619 32929 8628 32963
rect 8576 32920 8628 32929
rect 8760 32963 8812 32972
rect 8760 32929 8769 32963
rect 8769 32929 8803 32963
rect 8803 32929 8812 32963
rect 8760 32920 8812 32929
rect 8852 32920 8904 32972
rect 11152 32920 11204 32972
rect 12348 32920 12400 32972
rect 15568 32963 15620 32972
rect 4068 32852 4120 32904
rect 4712 32852 4764 32904
rect 6184 32895 6236 32904
rect 6184 32861 6193 32895
rect 6193 32861 6227 32895
rect 6227 32861 6236 32895
rect 6184 32852 6236 32861
rect 6828 32852 6880 32904
rect 9588 32852 9640 32904
rect 9956 32895 10008 32904
rect 9956 32861 9965 32895
rect 9965 32861 9999 32895
rect 9999 32861 10008 32895
rect 9956 32852 10008 32861
rect 12256 32895 12308 32904
rect 12256 32861 12265 32895
rect 12265 32861 12299 32895
rect 12299 32861 12308 32895
rect 12256 32852 12308 32861
rect 15292 32895 15344 32904
rect 15292 32861 15301 32895
rect 15301 32861 15335 32895
rect 15335 32861 15344 32895
rect 15292 32852 15344 32861
rect 15568 32929 15577 32963
rect 15577 32929 15611 32963
rect 15611 32929 15620 32963
rect 15568 32920 15620 32929
rect 19156 33056 19208 33108
rect 36728 33056 36780 33108
rect 29092 32988 29144 33040
rect 16948 32852 17000 32904
rect 7564 32784 7616 32836
rect 7380 32716 7432 32768
rect 9220 32716 9272 32768
rect 16304 32716 16356 32768
rect 16856 32759 16908 32768
rect 16856 32725 16865 32759
rect 16865 32725 16899 32759
rect 16899 32725 16908 32759
rect 16856 32716 16908 32725
rect 19984 32920 20036 32972
rect 20536 32920 20588 32972
rect 21640 32963 21692 32972
rect 21640 32929 21649 32963
rect 21649 32929 21683 32963
rect 21683 32929 21692 32963
rect 21640 32920 21692 32929
rect 22376 32920 22428 32972
rect 25964 32920 26016 32972
rect 27160 32920 27212 32972
rect 28632 32963 28684 32972
rect 28632 32929 28641 32963
rect 28641 32929 28675 32963
rect 28675 32929 28684 32963
rect 28632 32920 28684 32929
rect 29828 32920 29880 32972
rect 30564 32963 30616 32972
rect 30564 32929 30573 32963
rect 30573 32929 30607 32963
rect 30607 32929 30616 32963
rect 30564 32920 30616 32929
rect 33232 32963 33284 32972
rect 17684 32852 17736 32904
rect 23848 32852 23900 32904
rect 24216 32852 24268 32904
rect 17500 32784 17552 32836
rect 25780 32784 25832 32836
rect 25964 32784 26016 32836
rect 31760 32852 31812 32904
rect 32772 32895 32824 32904
rect 32772 32861 32781 32895
rect 32781 32861 32815 32895
rect 32815 32861 32824 32895
rect 32772 32852 32824 32861
rect 33232 32929 33241 32963
rect 33241 32929 33275 32963
rect 33275 32929 33284 32963
rect 33232 32920 33284 32929
rect 33600 32963 33652 32972
rect 33600 32929 33609 32963
rect 33609 32929 33643 32963
rect 33643 32929 33652 32963
rect 33600 32920 33652 32929
rect 35348 32963 35400 32972
rect 30748 32827 30800 32836
rect 30748 32793 30757 32827
rect 30757 32793 30791 32827
rect 30791 32793 30800 32827
rect 30748 32784 30800 32793
rect 34796 32895 34848 32904
rect 34796 32861 34805 32895
rect 34805 32861 34839 32895
rect 34839 32861 34848 32895
rect 34796 32852 34848 32861
rect 35348 32929 35357 32963
rect 35357 32929 35391 32963
rect 35391 32929 35400 32963
rect 35348 32920 35400 32929
rect 36360 32963 36412 32972
rect 36360 32929 36369 32963
rect 36369 32929 36403 32963
rect 36403 32929 36412 32963
rect 36360 32920 36412 32929
rect 37280 32920 37332 32972
rect 35716 32852 35768 32904
rect 35440 32784 35492 32836
rect 18512 32716 18564 32768
rect 18788 32716 18840 32768
rect 19340 32716 19392 32768
rect 21088 32759 21140 32768
rect 21088 32725 21097 32759
rect 21097 32725 21131 32759
rect 21131 32725 21140 32759
rect 21088 32716 21140 32725
rect 23756 32716 23808 32768
rect 24308 32716 24360 32768
rect 27804 32716 27856 32768
rect 27988 32716 28040 32768
rect 35624 32716 35676 32768
rect 4246 32614 4298 32666
rect 4310 32614 4362 32666
rect 4374 32614 4426 32666
rect 4438 32614 4490 32666
rect 34966 32614 35018 32666
rect 35030 32614 35082 32666
rect 35094 32614 35146 32666
rect 35158 32614 35210 32666
rect 6092 32512 6144 32564
rect 7932 32512 7984 32564
rect 2964 32444 3016 32496
rect 3976 32444 4028 32496
rect 4068 32376 4120 32428
rect 1860 32308 1912 32360
rect 2228 32351 2280 32360
rect 2228 32317 2237 32351
rect 2237 32317 2271 32351
rect 2271 32317 2280 32351
rect 2228 32308 2280 32317
rect 2872 32308 2924 32360
rect 3700 32351 3752 32360
rect 3700 32317 3709 32351
rect 3709 32317 3743 32351
rect 3743 32317 3752 32351
rect 3700 32308 3752 32317
rect 3884 32351 3936 32360
rect 3884 32317 3893 32351
rect 3893 32317 3927 32351
rect 3927 32317 3936 32351
rect 3884 32308 3936 32317
rect 4620 32351 4672 32360
rect 4620 32317 4629 32351
rect 4629 32317 4663 32351
rect 4663 32317 4672 32351
rect 4620 32308 4672 32317
rect 8024 32444 8076 32496
rect 12256 32444 12308 32496
rect 5540 32419 5592 32428
rect 5540 32385 5549 32419
rect 5549 32385 5583 32419
rect 5583 32385 5592 32419
rect 5540 32376 5592 32385
rect 6276 32419 6328 32428
rect 6276 32385 6285 32419
rect 6285 32385 6319 32419
rect 6319 32385 6328 32419
rect 6276 32376 6328 32385
rect 5724 32351 5776 32360
rect 5724 32317 5733 32351
rect 5733 32317 5767 32351
rect 5767 32317 5776 32351
rect 5724 32308 5776 32317
rect 8576 32376 8628 32428
rect 8852 32376 8904 32428
rect 8208 32351 8260 32360
rect 8208 32317 8217 32351
rect 8217 32317 8251 32351
rect 8251 32317 8260 32351
rect 8208 32308 8260 32317
rect 8300 32308 8352 32360
rect 8760 32308 8812 32360
rect 10876 32351 10928 32360
rect 6000 32240 6052 32292
rect 7656 32240 7708 32292
rect 8392 32240 8444 32292
rect 9772 32240 9824 32292
rect 10876 32317 10885 32351
rect 10885 32317 10919 32351
rect 10919 32317 10928 32351
rect 10876 32308 10928 32317
rect 11336 32351 11388 32360
rect 11336 32317 11345 32351
rect 11345 32317 11379 32351
rect 11379 32317 11388 32351
rect 11336 32308 11388 32317
rect 14280 32444 14332 32496
rect 14924 32351 14976 32360
rect 11060 32240 11112 32292
rect 14924 32317 14933 32351
rect 14933 32317 14967 32351
rect 14967 32317 14976 32351
rect 14924 32308 14976 32317
rect 17224 32512 17276 32564
rect 18420 32512 18472 32564
rect 32772 32555 32824 32564
rect 16304 32444 16356 32496
rect 17132 32444 17184 32496
rect 20352 32487 20404 32496
rect 15568 32308 15620 32360
rect 16580 32376 16632 32428
rect 16304 32308 16356 32360
rect 16672 32308 16724 32360
rect 16948 32308 17000 32360
rect 16764 32283 16816 32292
rect 16764 32249 16773 32283
rect 16773 32249 16807 32283
rect 16807 32249 16816 32283
rect 16764 32240 16816 32249
rect 18144 32376 18196 32428
rect 18788 32376 18840 32428
rect 20352 32453 20361 32487
rect 20361 32453 20395 32487
rect 20395 32453 20404 32487
rect 20352 32444 20404 32453
rect 22192 32444 22244 32496
rect 25504 32444 25556 32496
rect 30564 32487 30616 32496
rect 21088 32376 21140 32428
rect 23388 32376 23440 32428
rect 17776 32308 17828 32360
rect 18604 32351 18656 32360
rect 18604 32317 18613 32351
rect 18613 32317 18647 32351
rect 18647 32317 18656 32351
rect 18604 32308 18656 32317
rect 19892 32308 19944 32360
rect 20076 32308 20128 32360
rect 20352 32351 20404 32360
rect 20352 32317 20361 32351
rect 20361 32317 20395 32351
rect 20395 32317 20404 32351
rect 20352 32308 20404 32317
rect 22008 32351 22060 32360
rect 22008 32317 22017 32351
rect 22017 32317 22051 32351
rect 22051 32317 22060 32351
rect 22008 32308 22060 32317
rect 22376 32351 22428 32360
rect 1676 32215 1728 32224
rect 1676 32181 1685 32215
rect 1685 32181 1719 32215
rect 1719 32181 1728 32215
rect 1676 32172 1728 32181
rect 7288 32172 7340 32224
rect 8208 32172 8260 32224
rect 17224 32172 17276 32224
rect 21824 32240 21876 32292
rect 22376 32317 22385 32351
rect 22385 32317 22419 32351
rect 22419 32317 22428 32351
rect 22376 32308 22428 32317
rect 23756 32351 23808 32360
rect 23756 32317 23765 32351
rect 23765 32317 23799 32351
rect 23799 32317 23808 32351
rect 23756 32308 23808 32317
rect 25320 32308 25372 32360
rect 25964 32351 26016 32360
rect 25964 32317 25973 32351
rect 25973 32317 26007 32351
rect 26007 32317 26016 32351
rect 25964 32308 26016 32317
rect 29736 32376 29788 32428
rect 30564 32453 30573 32487
rect 30573 32453 30607 32487
rect 30607 32453 30616 32487
rect 30564 32444 30616 32453
rect 32772 32521 32781 32555
rect 32781 32521 32815 32555
rect 32815 32521 32824 32555
rect 32772 32512 32824 32521
rect 33600 32512 33652 32564
rect 36636 32512 36688 32564
rect 24032 32240 24084 32292
rect 18236 32172 18288 32224
rect 25228 32215 25280 32224
rect 25228 32181 25237 32215
rect 25237 32181 25271 32215
rect 25271 32181 25280 32215
rect 25228 32172 25280 32181
rect 29460 32308 29512 32360
rect 30288 32308 30340 32360
rect 30472 32351 30524 32360
rect 30472 32317 30481 32351
rect 30481 32317 30515 32351
rect 30515 32317 30524 32351
rect 30748 32376 30800 32428
rect 34796 32376 34848 32428
rect 30472 32308 30524 32317
rect 31024 32308 31076 32360
rect 31208 32351 31260 32360
rect 31208 32317 31217 32351
rect 31217 32317 31251 32351
rect 31251 32317 31260 32351
rect 31208 32308 31260 32317
rect 34888 32308 34940 32360
rect 35256 32308 35308 32360
rect 38108 32376 38160 32428
rect 30932 32240 30984 32292
rect 33416 32240 33468 32292
rect 37924 32308 37976 32360
rect 35808 32172 35860 32224
rect 37556 32172 37608 32224
rect 19606 32070 19658 32122
rect 19670 32070 19722 32122
rect 19734 32070 19786 32122
rect 19798 32070 19850 32122
rect 7104 31968 7156 32020
rect 8852 31968 8904 32020
rect 9220 32011 9272 32020
rect 9220 31977 9229 32011
rect 9229 31977 9263 32011
rect 9263 31977 9272 32011
rect 9220 31968 9272 31977
rect 15844 31968 15896 32020
rect 3240 31900 3292 31952
rect 4436 31900 4488 31952
rect 5080 31900 5132 31952
rect 6828 31943 6880 31952
rect 6828 31909 6837 31943
rect 6837 31909 6871 31943
rect 6871 31909 6880 31943
rect 6828 31900 6880 31909
rect 1676 31875 1728 31884
rect 1676 31841 1685 31875
rect 1685 31841 1719 31875
rect 1719 31841 1728 31875
rect 1676 31832 1728 31841
rect 4988 31832 5040 31884
rect 1400 31807 1452 31816
rect 1400 31773 1409 31807
rect 1409 31773 1443 31807
rect 1443 31773 1452 31807
rect 1400 31764 1452 31773
rect 4436 31764 4488 31816
rect 5172 31807 5224 31816
rect 5172 31773 5181 31807
rect 5181 31773 5215 31807
rect 5215 31773 5224 31807
rect 5172 31764 5224 31773
rect 5540 31764 5592 31816
rect 6460 31696 6512 31748
rect 7656 31875 7708 31884
rect 7656 31841 7665 31875
rect 7665 31841 7699 31875
rect 7699 31841 7708 31875
rect 7656 31832 7708 31841
rect 8116 31875 8168 31884
rect 8116 31841 8125 31875
rect 8125 31841 8159 31875
rect 8159 31841 8168 31875
rect 8116 31832 8168 31841
rect 8208 31832 8260 31884
rect 8852 31832 8904 31884
rect 9588 31832 9640 31884
rect 7932 31764 7984 31816
rect 10876 31832 10928 31884
rect 11244 31875 11296 31884
rect 11244 31841 11253 31875
rect 11253 31841 11287 31875
rect 11287 31841 11296 31875
rect 11244 31832 11296 31841
rect 14280 31875 14332 31884
rect 11428 31696 11480 31748
rect 5816 31628 5868 31680
rect 9956 31628 10008 31680
rect 10784 31628 10836 31680
rect 14280 31841 14289 31875
rect 14289 31841 14323 31875
rect 14323 31841 14332 31875
rect 14280 31832 14332 31841
rect 14372 31832 14424 31884
rect 16764 31900 16816 31952
rect 20076 31968 20128 32020
rect 18328 31943 18380 31952
rect 18328 31909 18337 31943
rect 18337 31909 18371 31943
rect 18371 31909 18380 31943
rect 18328 31900 18380 31909
rect 18512 31900 18564 31952
rect 20628 31968 20680 32020
rect 23388 31968 23440 32020
rect 20352 31943 20404 31952
rect 15568 31832 15620 31884
rect 12072 31807 12124 31816
rect 12072 31773 12081 31807
rect 12081 31773 12115 31807
rect 12115 31773 12124 31807
rect 12072 31764 12124 31773
rect 12716 31764 12768 31816
rect 13820 31764 13872 31816
rect 14924 31764 14976 31816
rect 16580 31832 16632 31884
rect 16856 31875 16908 31884
rect 16856 31841 16865 31875
rect 16865 31841 16899 31875
rect 16899 31841 16908 31875
rect 16856 31832 16908 31841
rect 17592 31832 17644 31884
rect 18236 31875 18288 31884
rect 18236 31841 18245 31875
rect 18245 31841 18279 31875
rect 18279 31841 18288 31875
rect 20352 31909 20361 31943
rect 20361 31909 20395 31943
rect 20395 31909 20404 31943
rect 20352 31900 20404 31909
rect 18236 31832 18288 31841
rect 20076 31875 20128 31884
rect 20076 31841 20085 31875
rect 20085 31841 20119 31875
rect 20119 31841 20128 31875
rect 20076 31832 20128 31841
rect 16212 31807 16264 31816
rect 16212 31773 16221 31807
rect 16221 31773 16255 31807
rect 16255 31773 16264 31807
rect 16212 31764 16264 31773
rect 18328 31764 18380 31816
rect 18604 31764 18656 31816
rect 21824 31875 21876 31884
rect 21824 31841 21833 31875
rect 21833 31841 21867 31875
rect 21867 31841 21876 31875
rect 21824 31832 21876 31841
rect 22008 31900 22060 31952
rect 23204 31832 23256 31884
rect 29276 31968 29328 32020
rect 29460 32011 29512 32020
rect 29460 31977 29469 32011
rect 29469 31977 29503 32011
rect 29503 31977 29512 32011
rect 29460 31968 29512 31977
rect 29736 31968 29788 32020
rect 33416 31900 33468 31952
rect 34888 31968 34940 32020
rect 23848 31832 23900 31884
rect 24032 31875 24084 31884
rect 24032 31841 24041 31875
rect 24041 31841 24075 31875
rect 24075 31841 24084 31875
rect 24032 31832 24084 31841
rect 24860 31832 24912 31884
rect 27988 31832 28040 31884
rect 28356 31875 28408 31884
rect 28356 31841 28365 31875
rect 28365 31841 28399 31875
rect 28399 31841 28408 31875
rect 28356 31832 28408 31841
rect 30656 31875 30708 31884
rect 30656 31841 30665 31875
rect 30665 31841 30699 31875
rect 30699 31841 30708 31875
rect 30656 31832 30708 31841
rect 32496 31832 32548 31884
rect 32772 31875 32824 31884
rect 32772 31841 32781 31875
rect 32781 31841 32815 31875
rect 32815 31841 32824 31875
rect 32772 31832 32824 31841
rect 33600 31875 33652 31884
rect 33600 31841 33609 31875
rect 33609 31841 33643 31875
rect 33643 31841 33652 31875
rect 33600 31832 33652 31841
rect 22376 31764 22428 31816
rect 25320 31807 25372 31816
rect 25320 31773 25329 31807
rect 25329 31773 25363 31807
rect 25363 31773 25372 31807
rect 25320 31764 25372 31773
rect 26608 31807 26660 31816
rect 26608 31773 26617 31807
rect 26617 31773 26651 31807
rect 26651 31773 26660 31807
rect 26608 31764 26660 31773
rect 27712 31764 27764 31816
rect 31760 31764 31812 31816
rect 32036 31764 32088 31816
rect 33968 31832 34020 31884
rect 35808 31875 35860 31884
rect 35808 31841 35817 31875
rect 35817 31841 35851 31875
rect 35851 31841 35860 31875
rect 35808 31832 35860 31841
rect 36728 31875 36780 31884
rect 36728 31841 36737 31875
rect 36737 31841 36771 31875
rect 36771 31841 36780 31875
rect 36728 31832 36780 31841
rect 37464 31832 37516 31884
rect 33876 31807 33928 31816
rect 33876 31773 33885 31807
rect 33885 31773 33919 31807
rect 33919 31773 33928 31807
rect 33876 31764 33928 31773
rect 35716 31807 35768 31816
rect 35716 31773 35725 31807
rect 35725 31773 35759 31807
rect 35759 31773 35768 31807
rect 35716 31764 35768 31773
rect 37280 31764 37332 31816
rect 19156 31696 19208 31748
rect 20352 31696 20404 31748
rect 20812 31696 20864 31748
rect 27252 31696 27304 31748
rect 30748 31739 30800 31748
rect 30748 31705 30757 31739
rect 30757 31705 30791 31739
rect 30791 31705 30800 31739
rect 30748 31696 30800 31705
rect 12532 31628 12584 31680
rect 16672 31628 16724 31680
rect 17592 31628 17644 31680
rect 36912 31628 36964 31680
rect 4246 31526 4298 31578
rect 4310 31526 4362 31578
rect 4374 31526 4426 31578
rect 4438 31526 4490 31578
rect 34966 31526 35018 31578
rect 35030 31526 35082 31578
rect 35094 31526 35146 31578
rect 35158 31526 35210 31578
rect 3516 31424 3568 31476
rect 3976 31424 4028 31476
rect 2872 31399 2924 31408
rect 2228 31288 2280 31340
rect 2872 31365 2881 31399
rect 2881 31365 2915 31399
rect 2915 31365 2924 31399
rect 2872 31356 2924 31365
rect 2780 31288 2832 31340
rect 3332 31288 3384 31340
rect 2136 31220 2188 31272
rect 3240 31220 3292 31272
rect 3700 31220 3752 31272
rect 3884 31263 3936 31272
rect 3884 31229 3893 31263
rect 3893 31229 3927 31263
rect 3927 31229 3936 31263
rect 3884 31220 3936 31229
rect 7104 31424 7156 31476
rect 9772 31424 9824 31476
rect 5632 31399 5684 31408
rect 5632 31365 5641 31399
rect 5641 31365 5675 31399
rect 5675 31365 5684 31399
rect 5632 31356 5684 31365
rect 11244 31356 11296 31408
rect 7380 31288 7432 31340
rect 10784 31331 10836 31340
rect 10784 31297 10793 31331
rect 10793 31297 10827 31331
rect 10827 31297 10836 31331
rect 10784 31288 10836 31297
rect 4436 31263 4488 31272
rect 4436 31229 4445 31263
rect 4445 31229 4479 31263
rect 4479 31229 4488 31263
rect 4436 31220 4488 31229
rect 5816 31263 5868 31272
rect 5816 31229 5825 31263
rect 5825 31229 5859 31263
rect 5859 31229 5868 31263
rect 5816 31220 5868 31229
rect 6184 31263 6236 31272
rect 6184 31229 6193 31263
rect 6193 31229 6227 31263
rect 6227 31229 6236 31263
rect 6184 31220 6236 31229
rect 7012 31220 7064 31272
rect 8116 31263 8168 31272
rect 8116 31229 8125 31263
rect 8125 31229 8159 31263
rect 8159 31229 8168 31263
rect 8116 31220 8168 31229
rect 9956 31263 10008 31272
rect 9956 31229 9965 31263
rect 9965 31229 9999 31263
rect 9999 31229 10008 31263
rect 9956 31220 10008 31229
rect 10048 31127 10100 31136
rect 10048 31093 10057 31127
rect 10057 31093 10091 31127
rect 10091 31093 10100 31127
rect 10048 31084 10100 31093
rect 11336 31220 11388 31272
rect 13084 31220 13136 31272
rect 23020 31467 23072 31476
rect 23020 31433 23029 31467
rect 23029 31433 23063 31467
rect 23063 31433 23072 31467
rect 23020 31424 23072 31433
rect 25964 31424 26016 31476
rect 27712 31424 27764 31476
rect 20260 31356 20312 31408
rect 20444 31356 20496 31408
rect 21824 31356 21876 31408
rect 13820 31331 13872 31340
rect 13820 31297 13829 31331
rect 13829 31297 13863 31331
rect 13863 31297 13872 31331
rect 13820 31288 13872 31297
rect 16856 31288 16908 31340
rect 20168 31288 20220 31340
rect 15292 31220 15344 31272
rect 16304 31263 16356 31272
rect 15200 31195 15252 31204
rect 15200 31161 15209 31195
rect 15209 31161 15243 31195
rect 15243 31161 15252 31195
rect 15200 31152 15252 31161
rect 12072 31084 12124 31136
rect 12900 31084 12952 31136
rect 14648 31084 14700 31136
rect 16304 31229 16313 31263
rect 16313 31229 16347 31263
rect 16347 31229 16356 31263
rect 16304 31220 16356 31229
rect 18604 31220 18656 31272
rect 18788 31263 18840 31272
rect 18788 31229 18797 31263
rect 18797 31229 18831 31263
rect 18831 31229 18840 31263
rect 18788 31220 18840 31229
rect 19984 31220 20036 31272
rect 20260 31152 20312 31204
rect 20996 31220 21048 31272
rect 21548 31263 21600 31272
rect 21548 31229 21557 31263
rect 21557 31229 21591 31263
rect 21591 31229 21600 31263
rect 21548 31220 21600 31229
rect 22836 31263 22888 31272
rect 20812 31152 20864 31204
rect 22836 31229 22845 31263
rect 22845 31229 22879 31263
rect 22879 31229 22888 31263
rect 22836 31220 22888 31229
rect 23204 31220 23256 31272
rect 25228 31356 25280 31408
rect 32496 31356 32548 31408
rect 25872 31288 25924 31340
rect 27252 31331 27304 31340
rect 27252 31297 27261 31331
rect 27261 31297 27295 31331
rect 27295 31297 27304 31331
rect 27252 31288 27304 31297
rect 30748 31288 30800 31340
rect 34244 31288 34296 31340
rect 36636 31288 36688 31340
rect 24308 31263 24360 31272
rect 24308 31229 24317 31263
rect 24317 31229 24351 31263
rect 24351 31229 24360 31263
rect 24308 31220 24360 31229
rect 25412 31263 25464 31272
rect 25412 31229 25421 31263
rect 25421 31229 25455 31263
rect 25455 31229 25464 31263
rect 25412 31220 25464 31229
rect 25596 31263 25648 31272
rect 25596 31229 25605 31263
rect 25605 31229 25639 31263
rect 25639 31229 25648 31263
rect 25596 31220 25648 31229
rect 25780 31263 25832 31272
rect 25780 31229 25789 31263
rect 25789 31229 25823 31263
rect 25823 31229 25832 31263
rect 25780 31220 25832 31229
rect 26884 31220 26936 31272
rect 26976 31263 27028 31272
rect 26976 31229 26985 31263
rect 26985 31229 27019 31263
rect 27019 31229 27028 31263
rect 28632 31263 28684 31272
rect 26976 31220 27028 31229
rect 28632 31229 28641 31263
rect 28641 31229 28675 31263
rect 28675 31229 28684 31263
rect 28632 31220 28684 31229
rect 30288 31220 30340 31272
rect 30472 31220 30524 31272
rect 30932 31220 30984 31272
rect 30564 31195 30616 31204
rect 30564 31161 30573 31195
rect 30573 31161 30607 31195
rect 30607 31161 30616 31195
rect 30564 31152 30616 31161
rect 16764 31084 16816 31136
rect 20536 31127 20588 31136
rect 20536 31093 20545 31127
rect 20545 31093 20579 31127
rect 20579 31093 20588 31127
rect 20536 31084 20588 31093
rect 24492 31127 24544 31136
rect 24492 31093 24501 31127
rect 24501 31093 24535 31127
rect 24535 31093 24544 31127
rect 24492 31084 24544 31093
rect 30196 31084 30248 31136
rect 33232 31220 33284 31272
rect 33968 31263 34020 31272
rect 33968 31229 33977 31263
rect 33977 31229 34011 31263
rect 34011 31229 34020 31263
rect 33968 31220 34020 31229
rect 34796 31220 34848 31272
rect 35348 31220 35400 31272
rect 36452 31263 36504 31272
rect 36452 31229 36461 31263
rect 36461 31229 36495 31263
rect 36495 31229 36504 31263
rect 36452 31220 36504 31229
rect 35440 31152 35492 31204
rect 32772 31084 32824 31136
rect 19606 30982 19658 31034
rect 19670 30982 19722 31034
rect 19734 30982 19786 31034
rect 19798 30982 19850 31034
rect 3608 30880 3660 30932
rect 5540 30880 5592 30932
rect 14648 30923 14700 30932
rect 14648 30889 14657 30923
rect 14657 30889 14691 30923
rect 14691 30889 14700 30923
rect 14648 30880 14700 30889
rect 16304 30880 16356 30932
rect 8116 30812 8168 30864
rect 16764 30855 16816 30864
rect 16764 30821 16773 30855
rect 16773 30821 16807 30855
rect 16807 30821 16816 30855
rect 16764 30812 16816 30821
rect 20260 30880 20312 30932
rect 22008 30880 22060 30932
rect 22376 30880 22428 30932
rect 24860 30880 24912 30932
rect 26608 30880 26660 30932
rect 33876 30880 33928 30932
rect 36728 30923 36780 30932
rect 36728 30889 36737 30923
rect 36737 30889 36771 30923
rect 36771 30889 36780 30923
rect 36728 30880 36780 30889
rect 19156 30812 19208 30864
rect 1860 30744 1912 30796
rect 2964 30787 3016 30796
rect 2964 30753 2973 30787
rect 2973 30753 3007 30787
rect 3007 30753 3016 30787
rect 2964 30744 3016 30753
rect 3608 30744 3660 30796
rect 5632 30787 5684 30796
rect 5632 30753 5641 30787
rect 5641 30753 5675 30787
rect 5675 30753 5684 30787
rect 5632 30744 5684 30753
rect 6828 30787 6880 30796
rect 6828 30753 6837 30787
rect 6837 30753 6871 30787
rect 6871 30753 6880 30787
rect 6828 30744 6880 30753
rect 7012 30787 7064 30796
rect 7012 30753 7021 30787
rect 7021 30753 7055 30787
rect 7055 30753 7064 30787
rect 7012 30744 7064 30753
rect 7656 30744 7708 30796
rect 8392 30787 8444 30796
rect 8392 30753 8401 30787
rect 8401 30753 8435 30787
rect 8435 30753 8444 30787
rect 8392 30744 8444 30753
rect 8668 30787 8720 30796
rect 8668 30753 8677 30787
rect 8677 30753 8711 30787
rect 8711 30753 8720 30787
rect 8668 30744 8720 30753
rect 8944 30744 8996 30796
rect 10324 30787 10376 30796
rect 10324 30753 10333 30787
rect 10333 30753 10367 30787
rect 10367 30753 10376 30787
rect 10324 30744 10376 30753
rect 11152 30787 11204 30796
rect 11152 30753 11161 30787
rect 11161 30753 11195 30787
rect 11195 30753 11204 30787
rect 11152 30744 11204 30753
rect 3148 30651 3200 30660
rect 3148 30617 3157 30651
rect 3157 30617 3191 30651
rect 3191 30617 3200 30651
rect 3148 30608 3200 30617
rect 6552 30676 6604 30728
rect 9772 30676 9824 30728
rect 11428 30719 11480 30728
rect 11428 30685 11437 30719
rect 11437 30685 11471 30719
rect 11471 30685 11480 30719
rect 11428 30676 11480 30685
rect 6460 30608 6512 30660
rect 13728 30744 13780 30796
rect 14464 30676 14516 30728
rect 15200 30744 15252 30796
rect 16396 30744 16448 30796
rect 13820 30608 13872 30660
rect 16764 30676 16816 30728
rect 17592 30744 17644 30796
rect 17960 30787 18012 30796
rect 17960 30753 17969 30787
rect 17969 30753 18003 30787
rect 18003 30753 18012 30787
rect 17960 30744 18012 30753
rect 18512 30787 18564 30796
rect 18512 30753 18521 30787
rect 18521 30753 18555 30787
rect 18555 30753 18564 30787
rect 18512 30744 18564 30753
rect 19432 30744 19484 30796
rect 20628 30744 20680 30796
rect 23572 30744 23624 30796
rect 25136 30812 25188 30864
rect 17316 30676 17368 30728
rect 20812 30676 20864 30728
rect 21088 30676 21140 30728
rect 22284 30719 22336 30728
rect 22284 30685 22293 30719
rect 22293 30685 22327 30719
rect 22327 30685 22336 30719
rect 22284 30676 22336 30685
rect 5632 30540 5684 30592
rect 9220 30540 9272 30592
rect 10416 30583 10468 30592
rect 10416 30549 10425 30583
rect 10425 30549 10459 30583
rect 10459 30549 10468 30583
rect 10416 30540 10468 30549
rect 12716 30583 12768 30592
rect 12716 30549 12725 30583
rect 12725 30549 12759 30583
rect 12759 30549 12768 30583
rect 12716 30540 12768 30549
rect 14740 30540 14792 30592
rect 16948 30540 17000 30592
rect 24952 30719 25004 30728
rect 24952 30685 24961 30719
rect 24961 30685 24995 30719
rect 24995 30685 25004 30719
rect 24952 30676 25004 30685
rect 26700 30744 26752 30796
rect 27160 30787 27212 30796
rect 27160 30753 27169 30787
rect 27169 30753 27203 30787
rect 27203 30753 27212 30787
rect 27160 30744 27212 30753
rect 27712 30787 27764 30796
rect 27712 30753 27721 30787
rect 27721 30753 27755 30787
rect 27755 30753 27764 30787
rect 27712 30744 27764 30753
rect 30564 30812 30616 30864
rect 30288 30787 30340 30796
rect 30288 30753 30297 30787
rect 30297 30753 30331 30787
rect 30331 30753 30340 30787
rect 30288 30744 30340 30753
rect 30472 30744 30524 30796
rect 32772 30744 32824 30796
rect 33692 30812 33744 30864
rect 35256 30812 35308 30864
rect 34244 30787 34296 30796
rect 34244 30753 34253 30787
rect 34253 30753 34287 30787
rect 34287 30753 34296 30787
rect 34244 30744 34296 30753
rect 35624 30787 35676 30796
rect 35624 30753 35633 30787
rect 35633 30753 35667 30787
rect 35667 30753 35676 30787
rect 35624 30744 35676 30753
rect 37740 30787 37792 30796
rect 37740 30753 37749 30787
rect 37749 30753 37783 30787
rect 37783 30753 37792 30787
rect 37740 30744 37792 30753
rect 27988 30719 28040 30728
rect 25412 30608 25464 30660
rect 27988 30685 27997 30719
rect 27997 30685 28031 30719
rect 28031 30685 28040 30719
rect 27988 30676 28040 30685
rect 31024 30676 31076 30728
rect 33140 30676 33192 30728
rect 30656 30651 30708 30660
rect 30656 30617 30665 30651
rect 30665 30617 30699 30651
rect 30699 30617 30708 30651
rect 30656 30608 30708 30617
rect 32036 30608 32088 30660
rect 27896 30540 27948 30592
rect 29276 30583 29328 30592
rect 29276 30549 29285 30583
rect 29285 30549 29319 30583
rect 29319 30549 29328 30583
rect 29276 30540 29328 30549
rect 36820 30540 36872 30592
rect 4246 30438 4298 30490
rect 4310 30438 4362 30490
rect 4374 30438 4426 30490
rect 4438 30438 4490 30490
rect 34966 30438 35018 30490
rect 35030 30438 35082 30490
rect 35094 30438 35146 30490
rect 35158 30438 35210 30490
rect 6644 30336 6696 30388
rect 13820 30336 13872 30388
rect 26700 30379 26752 30388
rect 26700 30345 26709 30379
rect 26709 30345 26743 30379
rect 26743 30345 26752 30379
rect 26700 30336 26752 30345
rect 30932 30336 30984 30388
rect 31392 30336 31444 30388
rect 33600 30336 33652 30388
rect 3608 30311 3660 30320
rect 3608 30277 3617 30311
rect 3617 30277 3651 30311
rect 3651 30277 3660 30311
rect 3608 30268 3660 30277
rect 8852 30268 8904 30320
rect 12624 30268 12676 30320
rect 17040 30268 17092 30320
rect 21548 30268 21600 30320
rect 3148 30200 3200 30252
rect 3700 30200 3752 30252
rect 4712 30200 4764 30252
rect 1400 30175 1452 30184
rect 1400 30141 1409 30175
rect 1409 30141 1443 30175
rect 1443 30141 1452 30175
rect 3516 30175 3568 30184
rect 1400 30132 1452 30141
rect 3516 30141 3525 30175
rect 3525 30141 3559 30175
rect 3559 30141 3568 30175
rect 3516 30132 3568 30141
rect 3884 30132 3936 30184
rect 7288 30200 7340 30252
rect 5908 30132 5960 30184
rect 7012 30175 7064 30184
rect 5172 30064 5224 30116
rect 7012 30141 7021 30175
rect 7021 30141 7055 30175
rect 7055 30141 7064 30175
rect 7012 30132 7064 30141
rect 7380 30175 7432 30184
rect 7380 30141 7389 30175
rect 7389 30141 7423 30175
rect 7423 30141 7432 30175
rect 7380 30132 7432 30141
rect 7564 30132 7616 30184
rect 8392 30175 8444 30184
rect 7932 30107 7984 30116
rect 7932 30073 7941 30107
rect 7941 30073 7975 30107
rect 7975 30073 7984 30107
rect 7932 30064 7984 30073
rect 8392 30141 8401 30175
rect 8401 30141 8435 30175
rect 8435 30141 8444 30175
rect 8392 30132 8444 30141
rect 10048 30200 10100 30252
rect 9404 30175 9456 30184
rect 9404 30141 9413 30175
rect 9413 30141 9447 30175
rect 9447 30141 9456 30175
rect 12992 30200 13044 30252
rect 9404 30132 9456 30141
rect 11612 30132 11664 30184
rect 12532 30175 12584 30184
rect 12532 30141 12541 30175
rect 12541 30141 12575 30175
rect 12575 30141 12584 30175
rect 12532 30132 12584 30141
rect 12900 30175 12952 30184
rect 12900 30141 12909 30175
rect 12909 30141 12943 30175
rect 12943 30141 12952 30175
rect 12900 30132 12952 30141
rect 14648 30200 14700 30252
rect 18512 30200 18564 30252
rect 20812 30243 20864 30252
rect 20812 30209 20821 30243
rect 20821 30209 20855 30243
rect 20855 30209 20864 30243
rect 20812 30200 20864 30209
rect 24952 30268 25004 30320
rect 27988 30268 28040 30320
rect 29368 30311 29420 30320
rect 29368 30277 29377 30311
rect 29377 30277 29411 30311
rect 29411 30277 29420 30311
rect 29368 30268 29420 30277
rect 35256 30268 35308 30320
rect 14280 30175 14332 30184
rect 14280 30141 14289 30175
rect 14289 30141 14323 30175
rect 14323 30141 14332 30175
rect 14280 30132 14332 30141
rect 14372 30132 14424 30184
rect 9128 30064 9180 30116
rect 11060 30107 11112 30116
rect 11060 30073 11069 30107
rect 11069 30073 11103 30107
rect 11103 30073 11112 30107
rect 11060 30064 11112 30073
rect 14556 30132 14608 30184
rect 15200 30132 15252 30184
rect 17040 30175 17092 30184
rect 17040 30141 17049 30175
rect 17049 30141 17083 30175
rect 17083 30141 17092 30175
rect 17040 30132 17092 30141
rect 17316 30175 17368 30184
rect 17316 30141 17325 30175
rect 17325 30141 17359 30175
rect 17359 30141 17368 30175
rect 17316 30132 17368 30141
rect 2872 29996 2924 30048
rect 4988 29996 5040 30048
rect 5264 29996 5316 30048
rect 5448 30039 5500 30048
rect 5448 30005 5457 30039
rect 5457 30005 5491 30039
rect 5491 30005 5500 30039
rect 5448 29996 5500 30005
rect 7196 29996 7248 30048
rect 11612 30039 11664 30048
rect 11612 30005 11621 30039
rect 11621 30005 11655 30039
rect 11655 30005 11664 30039
rect 11612 29996 11664 30005
rect 12348 29996 12400 30048
rect 17408 30064 17460 30116
rect 15660 29996 15712 30048
rect 15752 30039 15804 30048
rect 15752 30005 15761 30039
rect 15761 30005 15795 30039
rect 15795 30005 15804 30039
rect 15752 29996 15804 30005
rect 16028 29996 16080 30048
rect 16396 29996 16448 30048
rect 18052 30132 18104 30184
rect 19432 30132 19484 30184
rect 19984 30175 20036 30184
rect 19984 30141 19993 30175
rect 19993 30141 20027 30175
rect 20027 30141 20036 30175
rect 19984 30132 20036 30141
rect 20628 30132 20680 30184
rect 20996 30132 21048 30184
rect 22468 30132 22520 30184
rect 22652 30175 22704 30184
rect 22652 30141 22661 30175
rect 22661 30141 22695 30175
rect 22695 30141 22704 30175
rect 22652 30132 22704 30141
rect 25596 30243 25648 30252
rect 25596 30209 25605 30243
rect 25605 30209 25639 30243
rect 25639 30209 25648 30243
rect 25596 30200 25648 30209
rect 33140 30200 33192 30252
rect 36452 30243 36504 30252
rect 23480 30132 23532 30184
rect 23848 30175 23900 30184
rect 23848 30141 23857 30175
rect 23857 30141 23891 30175
rect 23891 30141 23900 30175
rect 23848 30132 23900 30141
rect 24216 30175 24268 30184
rect 24216 30141 24225 30175
rect 24225 30141 24259 30175
rect 24259 30141 24268 30175
rect 24216 30132 24268 30141
rect 19340 30064 19392 30116
rect 25044 30064 25096 30116
rect 18972 29996 19024 30048
rect 20076 29996 20128 30048
rect 27160 30132 27212 30184
rect 26424 30064 26476 30116
rect 29000 30132 29052 30184
rect 29460 30175 29512 30184
rect 29460 30141 29469 30175
rect 29469 30141 29503 30175
rect 29503 30141 29512 30175
rect 29460 30132 29512 30141
rect 29644 30132 29696 30184
rect 29828 30175 29880 30184
rect 29828 30141 29837 30175
rect 29837 30141 29871 30175
rect 29871 30141 29880 30175
rect 29828 30132 29880 30141
rect 30932 30132 30984 30184
rect 31852 30175 31904 30184
rect 31852 30141 31861 30175
rect 31861 30141 31895 30175
rect 31895 30141 31904 30175
rect 31852 30132 31904 30141
rect 32036 30175 32088 30184
rect 32036 30141 32045 30175
rect 32045 30141 32079 30175
rect 32079 30141 32088 30175
rect 32036 30132 32088 30141
rect 32956 30132 33008 30184
rect 33416 30132 33468 30184
rect 34520 30132 34572 30184
rect 35624 30175 35676 30184
rect 34244 30064 34296 30116
rect 35624 30141 35633 30175
rect 35633 30141 35667 30175
rect 35667 30141 35676 30175
rect 35624 30132 35676 30141
rect 35900 30064 35952 30116
rect 26976 29996 27028 30048
rect 27436 29996 27488 30048
rect 31668 29996 31720 30048
rect 32772 29996 32824 30048
rect 34612 29996 34664 30048
rect 36452 30209 36461 30243
rect 36461 30209 36495 30243
rect 36495 30209 36504 30243
rect 36452 30200 36504 30209
rect 37372 30132 37424 30184
rect 37556 30132 37608 30184
rect 37188 29996 37240 30048
rect 37556 29996 37608 30048
rect 19606 29894 19658 29946
rect 19670 29894 19722 29946
rect 19734 29894 19786 29946
rect 19798 29894 19850 29946
rect 3516 29792 3568 29844
rect 3884 29792 3936 29844
rect 4620 29792 4672 29844
rect 4804 29792 4856 29844
rect 5264 29792 5316 29844
rect 5172 29724 5224 29776
rect 2872 29699 2924 29708
rect 2872 29665 2881 29699
rect 2881 29665 2915 29699
rect 2915 29665 2924 29699
rect 2872 29656 2924 29665
rect 4068 29699 4120 29708
rect 4068 29665 4077 29699
rect 4077 29665 4111 29699
rect 4111 29665 4120 29699
rect 4068 29656 4120 29665
rect 5264 29656 5316 29708
rect 7380 29724 7432 29776
rect 5632 29699 5684 29708
rect 5632 29665 5641 29699
rect 5641 29665 5675 29699
rect 5675 29665 5684 29699
rect 5632 29656 5684 29665
rect 6552 29656 6604 29708
rect 7932 29699 7984 29708
rect 7932 29665 7941 29699
rect 7941 29665 7975 29699
rect 7975 29665 7984 29699
rect 7932 29656 7984 29665
rect 7012 29631 7064 29640
rect 7012 29597 7021 29631
rect 7021 29597 7055 29631
rect 7055 29597 7064 29631
rect 8392 29656 8444 29708
rect 12624 29792 12676 29844
rect 13728 29792 13780 29844
rect 14556 29835 14608 29844
rect 12348 29699 12400 29708
rect 7012 29588 7064 29597
rect 9036 29588 9088 29640
rect 12348 29665 12357 29699
rect 12357 29665 12391 29699
rect 12391 29665 12400 29699
rect 12348 29656 12400 29665
rect 12992 29699 13044 29708
rect 12992 29665 13001 29699
rect 13001 29665 13035 29699
rect 13035 29665 13044 29699
rect 12992 29656 13044 29665
rect 14556 29801 14565 29835
rect 14565 29801 14599 29835
rect 14599 29801 14608 29835
rect 14556 29792 14608 29801
rect 15660 29792 15712 29844
rect 21180 29792 21232 29844
rect 17960 29724 18012 29776
rect 19156 29724 19208 29776
rect 25780 29792 25832 29844
rect 11336 29588 11388 29640
rect 14464 29656 14516 29708
rect 15752 29656 15804 29708
rect 16028 29656 16080 29708
rect 17500 29656 17552 29708
rect 20168 29699 20220 29708
rect 20168 29665 20177 29699
rect 20177 29665 20211 29699
rect 20211 29665 20220 29699
rect 20168 29656 20220 29665
rect 23204 29724 23256 29776
rect 24216 29724 24268 29776
rect 22928 29699 22980 29708
rect 16764 29588 16816 29640
rect 18236 29588 18288 29640
rect 20076 29588 20128 29640
rect 20536 29588 20588 29640
rect 22928 29665 22937 29699
rect 22937 29665 22971 29699
rect 22971 29665 22980 29699
rect 22928 29656 22980 29665
rect 23296 29699 23348 29708
rect 23296 29665 23305 29699
rect 23305 29665 23339 29699
rect 23339 29665 23348 29699
rect 23296 29656 23348 29665
rect 23572 29699 23624 29708
rect 23572 29665 23581 29699
rect 23581 29665 23615 29699
rect 23615 29665 23624 29699
rect 23572 29656 23624 29665
rect 24768 29699 24820 29708
rect 24768 29665 24777 29699
rect 24777 29665 24811 29699
rect 24811 29665 24820 29699
rect 24768 29656 24820 29665
rect 25044 29699 25096 29708
rect 25044 29665 25053 29699
rect 25053 29665 25087 29699
rect 25087 29665 25096 29699
rect 25044 29656 25096 29665
rect 25504 29699 25556 29708
rect 25504 29665 25513 29699
rect 25513 29665 25547 29699
rect 25547 29665 25556 29699
rect 25504 29656 25556 29665
rect 26056 29656 26108 29708
rect 29920 29792 29972 29844
rect 32772 29792 32824 29844
rect 31852 29724 31904 29776
rect 7564 29520 7616 29572
rect 10600 29563 10652 29572
rect 10600 29529 10609 29563
rect 10609 29529 10643 29563
rect 10643 29529 10652 29563
rect 10600 29520 10652 29529
rect 2964 29452 3016 29504
rect 8484 29452 8536 29504
rect 9036 29495 9088 29504
rect 9036 29461 9045 29495
rect 9045 29461 9079 29495
rect 9079 29461 9088 29495
rect 9036 29452 9088 29461
rect 9128 29452 9180 29504
rect 17960 29520 18012 29572
rect 17132 29452 17184 29504
rect 19708 29520 19760 29572
rect 19800 29520 19852 29572
rect 21088 29520 21140 29572
rect 26424 29588 26476 29640
rect 27620 29588 27672 29640
rect 28080 29631 28132 29640
rect 27436 29520 27488 29572
rect 28080 29597 28089 29631
rect 28089 29597 28123 29631
rect 28123 29597 28132 29631
rect 28080 29588 28132 29597
rect 29276 29656 29328 29708
rect 30288 29699 30340 29708
rect 30288 29665 30297 29699
rect 30297 29665 30331 29699
rect 30331 29665 30340 29699
rect 30288 29656 30340 29665
rect 30472 29656 30524 29708
rect 31024 29656 31076 29708
rect 32864 29699 32916 29708
rect 32864 29665 32873 29699
rect 32873 29665 32907 29699
rect 32907 29665 32916 29699
rect 32864 29656 32916 29665
rect 33140 29699 33192 29708
rect 33140 29665 33149 29699
rect 33149 29665 33183 29699
rect 33183 29665 33192 29699
rect 33140 29656 33192 29665
rect 33600 29656 33652 29708
rect 35624 29656 35676 29708
rect 36820 29699 36872 29708
rect 36820 29665 36829 29699
rect 36829 29665 36863 29699
rect 36863 29665 36872 29699
rect 36820 29656 36872 29665
rect 37648 29656 37700 29708
rect 29644 29588 29696 29640
rect 31760 29588 31812 29640
rect 32956 29588 33008 29640
rect 34152 29631 34204 29640
rect 34152 29597 34161 29631
rect 34161 29597 34195 29631
rect 34195 29597 34204 29631
rect 34152 29588 34204 29597
rect 37096 29631 37148 29640
rect 37096 29597 37105 29631
rect 37105 29597 37139 29631
rect 37139 29597 37148 29631
rect 37096 29588 37148 29597
rect 32772 29520 32824 29572
rect 36728 29520 36780 29572
rect 19432 29452 19484 29504
rect 20168 29452 20220 29504
rect 35256 29495 35308 29504
rect 35256 29461 35265 29495
rect 35265 29461 35299 29495
rect 35299 29461 35308 29495
rect 35256 29452 35308 29461
rect 36820 29452 36872 29504
rect 4246 29350 4298 29402
rect 4310 29350 4362 29402
rect 4374 29350 4426 29402
rect 4438 29350 4490 29402
rect 34966 29350 35018 29402
rect 35030 29350 35082 29402
rect 35094 29350 35146 29402
rect 35158 29350 35210 29402
rect 4068 29248 4120 29300
rect 9956 29248 10008 29300
rect 18236 29248 18288 29300
rect 19800 29248 19852 29300
rect 20444 29248 20496 29300
rect 21732 29248 21784 29300
rect 26424 29248 26476 29300
rect 26884 29291 26936 29300
rect 26884 29257 26893 29291
rect 26893 29257 26927 29291
rect 26927 29257 26936 29291
rect 26884 29248 26936 29257
rect 6092 29180 6144 29232
rect 2780 29044 2832 29096
rect 2964 29087 3016 29096
rect 2964 29053 2973 29087
rect 2973 29053 3007 29087
rect 3007 29053 3016 29087
rect 2964 29044 3016 29053
rect 3240 29044 3292 29096
rect 4712 29112 4764 29164
rect 5908 29112 5960 29164
rect 6828 29112 6880 29164
rect 4068 29044 4120 29096
rect 4620 29044 4672 29096
rect 7012 29087 7064 29096
rect 4804 28976 4856 29028
rect 5172 28976 5224 29028
rect 7012 29053 7021 29087
rect 7021 29053 7055 29087
rect 7055 29053 7064 29087
rect 7012 29044 7064 29053
rect 10416 29112 10468 29164
rect 8668 29044 8720 29096
rect 9404 29044 9456 29096
rect 12164 29112 12216 29164
rect 6920 28976 6972 29028
rect 10692 29044 10744 29096
rect 12716 29180 12768 29232
rect 14280 29180 14332 29232
rect 15844 29180 15896 29232
rect 12716 29044 12768 29096
rect 14556 29112 14608 29164
rect 16028 29112 16080 29164
rect 19432 29180 19484 29232
rect 21180 29180 21232 29232
rect 28080 29223 28132 29232
rect 14372 29087 14424 29096
rect 14372 29053 14381 29087
rect 14381 29053 14415 29087
rect 14415 29053 14424 29087
rect 14372 29044 14424 29053
rect 14924 29087 14976 29096
rect 14924 29053 14933 29087
rect 14933 29053 14967 29087
rect 14967 29053 14976 29087
rect 14924 29044 14976 29053
rect 2872 28908 2924 28960
rect 2964 28908 3016 28960
rect 4896 28908 4948 28960
rect 7564 28908 7616 28960
rect 13360 28976 13412 29028
rect 9680 28951 9732 28960
rect 9680 28917 9689 28951
rect 9689 28917 9723 28951
rect 9723 28917 9732 28951
rect 17040 29044 17092 29096
rect 19340 29112 19392 29164
rect 18972 29087 19024 29096
rect 18972 29053 18981 29087
rect 18981 29053 19015 29087
rect 19015 29053 19024 29087
rect 18972 29044 19024 29053
rect 19800 29044 19852 29096
rect 20260 29044 20312 29096
rect 20444 29087 20496 29096
rect 20444 29053 20453 29087
rect 20453 29053 20487 29087
rect 20487 29053 20496 29087
rect 20444 29044 20496 29053
rect 28080 29189 28089 29223
rect 28089 29189 28123 29223
rect 28123 29189 28132 29223
rect 28080 29180 28132 29189
rect 22652 29155 22704 29164
rect 22652 29121 22661 29155
rect 22661 29121 22695 29155
rect 22695 29121 22704 29155
rect 22652 29112 22704 29121
rect 22928 29112 22980 29164
rect 23848 29112 23900 29164
rect 24676 29112 24728 29164
rect 24768 29087 24820 29096
rect 19156 28976 19208 29028
rect 19984 28976 20036 29028
rect 23388 28976 23440 29028
rect 24768 29053 24777 29087
rect 24777 29053 24811 29087
rect 24811 29053 24820 29087
rect 24768 29044 24820 29053
rect 25228 29087 25280 29096
rect 25228 29053 25237 29087
rect 25237 29053 25271 29087
rect 25271 29053 25280 29087
rect 25228 29044 25280 29053
rect 25320 29044 25372 29096
rect 26056 29087 26108 29096
rect 26056 29053 26065 29087
rect 26065 29053 26099 29087
rect 26099 29053 26108 29087
rect 26056 29044 26108 29053
rect 26148 28976 26200 29028
rect 27160 29087 27212 29096
rect 27160 29053 27169 29087
rect 27169 29053 27203 29087
rect 27203 29053 27212 29087
rect 27160 29044 27212 29053
rect 27620 29044 27672 29096
rect 31024 29248 31076 29300
rect 32956 29291 33008 29300
rect 32956 29257 32965 29291
rect 32965 29257 32999 29291
rect 32999 29257 33008 29291
rect 32956 29248 33008 29257
rect 37740 29248 37792 29300
rect 34428 29180 34480 29232
rect 29920 29155 29972 29164
rect 29920 29121 29929 29155
rect 29929 29121 29963 29155
rect 29963 29121 29972 29155
rect 29920 29112 29972 29121
rect 30932 29155 30984 29164
rect 30932 29121 30941 29155
rect 30941 29121 30975 29155
rect 30975 29121 30984 29155
rect 30932 29112 30984 29121
rect 31392 29155 31444 29164
rect 31392 29121 31401 29155
rect 31401 29121 31435 29155
rect 31435 29121 31444 29155
rect 31392 29112 31444 29121
rect 31668 29155 31720 29164
rect 31668 29121 31677 29155
rect 31677 29121 31711 29155
rect 31711 29121 31720 29155
rect 31668 29112 31720 29121
rect 35348 29112 35400 29164
rect 36452 29155 36504 29164
rect 36452 29121 36461 29155
rect 36461 29121 36495 29155
rect 36495 29121 36504 29155
rect 36452 29112 36504 29121
rect 36728 29155 36780 29164
rect 36728 29121 36737 29155
rect 36737 29121 36771 29155
rect 36771 29121 36780 29155
rect 36728 29112 36780 29121
rect 29460 29044 29512 29096
rect 30380 29087 30432 29096
rect 30380 29053 30389 29087
rect 30389 29053 30423 29087
rect 30423 29053 30432 29087
rect 30380 29044 30432 29053
rect 30472 29044 30524 29096
rect 35256 29044 35308 29096
rect 35532 29044 35584 29096
rect 33508 28976 33560 29028
rect 34704 28976 34756 29028
rect 35440 28976 35492 29028
rect 9680 28908 9732 28917
rect 20168 28908 20220 28960
rect 20812 28908 20864 28960
rect 21088 28908 21140 28960
rect 36728 28908 36780 28960
rect 37924 28976 37976 29028
rect 38016 28908 38068 28960
rect 19606 28806 19658 28858
rect 19670 28806 19722 28858
rect 19734 28806 19786 28858
rect 19798 28806 19850 28858
rect 7380 28704 7432 28756
rect 11612 28704 11664 28756
rect 13268 28704 13320 28756
rect 13360 28704 13412 28756
rect 17040 28747 17092 28756
rect 17040 28713 17049 28747
rect 17049 28713 17083 28747
rect 17083 28713 17092 28747
rect 17040 28704 17092 28713
rect 20444 28704 20496 28756
rect 20628 28704 20680 28756
rect 21548 28704 21600 28756
rect 22284 28747 22336 28756
rect 22284 28713 22293 28747
rect 22293 28713 22327 28747
rect 22327 28713 22336 28747
rect 22284 28704 22336 28713
rect 5448 28636 5500 28688
rect 4620 28611 4672 28620
rect 4620 28577 4629 28611
rect 4629 28577 4663 28611
rect 4663 28577 4672 28611
rect 4620 28568 4672 28577
rect 4896 28611 4948 28620
rect 4896 28577 4905 28611
rect 4905 28577 4939 28611
rect 4939 28577 4948 28611
rect 4896 28568 4948 28577
rect 5816 28611 5868 28620
rect 5816 28577 5825 28611
rect 5825 28577 5859 28611
rect 5859 28577 5868 28611
rect 5816 28568 5868 28577
rect 11428 28636 11480 28688
rect 1400 28543 1452 28552
rect 1400 28509 1409 28543
rect 1409 28509 1443 28543
rect 1443 28509 1452 28543
rect 1400 28500 1452 28509
rect 1860 28500 1912 28552
rect 4712 28500 4764 28552
rect 5356 28500 5408 28552
rect 7932 28568 7984 28620
rect 9956 28611 10008 28620
rect 9956 28577 9965 28611
rect 9965 28577 9999 28611
rect 9999 28577 10008 28611
rect 9956 28568 10008 28577
rect 10324 28568 10376 28620
rect 10600 28568 10652 28620
rect 11612 28568 11664 28620
rect 12716 28611 12768 28620
rect 12716 28577 12725 28611
rect 12725 28577 12759 28611
rect 12759 28577 12768 28611
rect 12716 28568 12768 28577
rect 12900 28500 12952 28552
rect 13452 28568 13504 28620
rect 20536 28636 20588 28688
rect 20812 28636 20864 28688
rect 15384 28611 15436 28620
rect 15384 28577 15393 28611
rect 15393 28577 15427 28611
rect 15427 28577 15436 28611
rect 15384 28568 15436 28577
rect 15752 28611 15804 28620
rect 15752 28577 15761 28611
rect 15761 28577 15795 28611
rect 15795 28577 15804 28611
rect 15752 28568 15804 28577
rect 16212 28611 16264 28620
rect 16212 28577 16221 28611
rect 16221 28577 16255 28611
rect 16255 28577 16264 28611
rect 16212 28568 16264 28577
rect 16948 28611 17000 28620
rect 16948 28577 16957 28611
rect 16957 28577 16991 28611
rect 16991 28577 17000 28611
rect 16948 28568 17000 28577
rect 17684 28611 17736 28620
rect 17684 28577 17693 28611
rect 17693 28577 17727 28611
rect 17727 28577 17736 28611
rect 17684 28568 17736 28577
rect 16120 28500 16172 28552
rect 18328 28568 18380 28620
rect 19892 28568 19944 28620
rect 20720 28568 20772 28620
rect 21088 28568 21140 28620
rect 21732 28636 21784 28688
rect 32312 28704 32364 28756
rect 26056 28636 26108 28688
rect 22192 28611 22244 28620
rect 22192 28577 22201 28611
rect 22201 28577 22235 28611
rect 22235 28577 22244 28611
rect 22192 28568 22244 28577
rect 23020 28611 23072 28620
rect 23020 28577 23029 28611
rect 23029 28577 23063 28611
rect 23063 28577 23072 28611
rect 23020 28568 23072 28577
rect 18420 28500 18472 28552
rect 19432 28500 19484 28552
rect 20260 28500 20312 28552
rect 23664 28611 23716 28620
rect 23664 28577 23673 28611
rect 23673 28577 23707 28611
rect 23707 28577 23716 28611
rect 24860 28611 24912 28620
rect 23664 28568 23716 28577
rect 24860 28577 24869 28611
rect 24869 28577 24903 28611
rect 24903 28577 24912 28611
rect 24860 28568 24912 28577
rect 24952 28611 25004 28620
rect 24952 28577 24961 28611
rect 24961 28577 24995 28611
rect 24995 28577 25004 28611
rect 25320 28611 25372 28620
rect 24952 28568 25004 28577
rect 25320 28577 25329 28611
rect 25329 28577 25363 28611
rect 25363 28577 25372 28611
rect 25320 28568 25372 28577
rect 26516 28611 26568 28620
rect 26516 28577 26525 28611
rect 26525 28577 26559 28611
rect 26559 28577 26568 28611
rect 26516 28568 26568 28577
rect 29368 28636 29420 28688
rect 33508 28704 33560 28756
rect 34152 28704 34204 28756
rect 33140 28636 33192 28688
rect 37648 28704 37700 28756
rect 26884 28543 26936 28552
rect 2412 28432 2464 28484
rect 5724 28475 5776 28484
rect 5724 28441 5733 28475
rect 5733 28441 5767 28475
rect 5767 28441 5776 28475
rect 5724 28432 5776 28441
rect 12164 28432 12216 28484
rect 26884 28509 26893 28543
rect 26893 28509 26927 28543
rect 26927 28509 26936 28543
rect 26884 28500 26936 28509
rect 26976 28500 27028 28552
rect 29276 28568 29328 28620
rect 29644 28611 29696 28620
rect 29644 28577 29653 28611
rect 29653 28577 29687 28611
rect 29687 28577 29696 28611
rect 29644 28568 29696 28577
rect 30656 28611 30708 28620
rect 30656 28577 30665 28611
rect 30665 28577 30699 28611
rect 30699 28577 30708 28611
rect 30656 28568 30708 28577
rect 32404 28568 32456 28620
rect 27896 28500 27948 28552
rect 31484 28543 31536 28552
rect 31484 28509 31493 28543
rect 31493 28509 31527 28543
rect 31527 28509 31536 28543
rect 31484 28500 31536 28509
rect 32772 28568 32824 28620
rect 34244 28611 34296 28620
rect 34244 28577 34253 28611
rect 34253 28577 34287 28611
rect 34287 28577 34296 28611
rect 34244 28568 34296 28577
rect 33784 28500 33836 28552
rect 35532 28568 35584 28620
rect 36360 28611 36412 28620
rect 36360 28577 36369 28611
rect 36369 28577 36403 28611
rect 36403 28577 36412 28611
rect 36360 28568 36412 28577
rect 36452 28611 36504 28620
rect 36452 28577 36461 28611
rect 36461 28577 36495 28611
rect 36495 28577 36504 28611
rect 36452 28568 36504 28577
rect 37648 28568 37700 28620
rect 28540 28432 28592 28484
rect 29000 28475 29052 28484
rect 29000 28441 29009 28475
rect 29009 28441 29043 28475
rect 29043 28441 29052 28475
rect 29000 28432 29052 28441
rect 30564 28475 30616 28484
rect 30564 28441 30573 28475
rect 30573 28441 30607 28475
rect 30607 28441 30616 28475
rect 30564 28432 30616 28441
rect 32036 28432 32088 28484
rect 36544 28500 36596 28552
rect 2964 28407 3016 28416
rect 2964 28373 2973 28407
rect 2973 28373 3007 28407
rect 3007 28373 3016 28407
rect 2964 28364 3016 28373
rect 8208 28364 8260 28416
rect 37188 28364 37240 28416
rect 4246 28262 4298 28314
rect 4310 28262 4362 28314
rect 4374 28262 4426 28314
rect 4438 28262 4490 28314
rect 34966 28262 35018 28314
rect 35030 28262 35082 28314
rect 35094 28262 35146 28314
rect 35158 28262 35210 28314
rect 1860 28203 1912 28212
rect 1860 28169 1869 28203
rect 1869 28169 1903 28203
rect 1903 28169 1912 28203
rect 1860 28160 1912 28169
rect 4712 28160 4764 28212
rect 8208 28160 8260 28212
rect 3332 28135 3384 28144
rect 3332 28101 3341 28135
rect 3341 28101 3375 28135
rect 3375 28101 3384 28135
rect 3332 28092 3384 28101
rect 5816 28135 5868 28144
rect 5816 28101 5825 28135
rect 5825 28101 5859 28135
rect 5859 28101 5868 28135
rect 5816 28092 5868 28101
rect 7932 28135 7984 28144
rect 2964 28024 3016 28076
rect 2412 27956 2464 28008
rect 2780 27999 2832 28008
rect 2780 27965 2789 27999
rect 2789 27965 2823 27999
rect 2823 27965 2832 27999
rect 3240 27999 3292 28008
rect 2780 27956 2832 27965
rect 3240 27965 3249 27999
rect 3249 27965 3283 27999
rect 3283 27965 3292 27999
rect 3240 27956 3292 27965
rect 4068 27956 4120 28008
rect 5448 28024 5500 28076
rect 5356 27999 5408 28008
rect 5356 27965 5365 27999
rect 5365 27965 5399 27999
rect 5399 27965 5408 27999
rect 5356 27956 5408 27965
rect 6368 27956 6420 28008
rect 6920 27956 6972 28008
rect 7932 28101 7941 28135
rect 7941 28101 7975 28135
rect 7975 28101 7984 28135
rect 7932 28092 7984 28101
rect 8668 28135 8720 28144
rect 8668 28101 8677 28135
rect 8677 28101 8711 28135
rect 8711 28101 8720 28135
rect 8668 28092 8720 28101
rect 8484 27956 8536 28008
rect 8852 27999 8904 28008
rect 8852 27965 8861 27999
rect 8861 27965 8895 27999
rect 8895 27965 8904 27999
rect 8852 27956 8904 27965
rect 9588 28092 9640 28144
rect 9680 28092 9732 28144
rect 9956 28067 10008 28076
rect 9956 28033 9965 28067
rect 9965 28033 9999 28067
rect 9999 28033 10008 28067
rect 9956 28024 10008 28033
rect 10600 28067 10652 28076
rect 10600 28033 10609 28067
rect 10609 28033 10643 28067
rect 10643 28033 10652 28067
rect 10600 28024 10652 28033
rect 11336 28024 11388 28076
rect 12440 28092 12492 28144
rect 14372 28160 14424 28212
rect 15292 28092 15344 28144
rect 9772 27999 9824 28008
rect 9772 27965 9781 27999
rect 9781 27965 9815 27999
rect 9815 27965 9824 27999
rect 9772 27956 9824 27965
rect 11428 27999 11480 28008
rect 11428 27965 11437 27999
rect 11437 27965 11471 27999
rect 11471 27965 11480 27999
rect 11428 27956 11480 27965
rect 12072 27956 12124 28008
rect 7564 27820 7616 27872
rect 11060 27820 11112 27872
rect 13820 27956 13872 28008
rect 17132 28160 17184 28212
rect 23020 28203 23072 28212
rect 23020 28169 23029 28203
rect 23029 28169 23063 28203
rect 23063 28169 23072 28203
rect 23020 28160 23072 28169
rect 31944 28160 31996 28212
rect 32312 28160 32364 28212
rect 16212 28092 16264 28144
rect 18328 28135 18380 28144
rect 18328 28101 18337 28135
rect 18337 28101 18371 28135
rect 18371 28101 18380 28135
rect 18328 28092 18380 28101
rect 23572 28092 23624 28144
rect 24860 28092 24912 28144
rect 16120 28067 16172 28076
rect 16120 28033 16129 28067
rect 16129 28033 16163 28067
rect 16163 28033 16172 28067
rect 16120 28024 16172 28033
rect 17684 28024 17736 28076
rect 15936 27999 15988 28008
rect 14372 27888 14424 27940
rect 15936 27965 15945 27999
rect 15945 27965 15979 27999
rect 15979 27965 15988 27999
rect 15936 27956 15988 27965
rect 17500 27956 17552 28008
rect 18052 27999 18104 28008
rect 18052 27965 18061 27999
rect 18061 27965 18095 27999
rect 18095 27965 18104 27999
rect 18052 27956 18104 27965
rect 18420 27956 18472 28008
rect 20628 28024 20680 28076
rect 22008 28024 22060 28076
rect 26884 28067 26936 28076
rect 26884 28033 26893 28067
rect 26893 28033 26927 28067
rect 26927 28033 26936 28067
rect 26884 28024 26936 28033
rect 32404 28092 32456 28144
rect 33416 28160 33468 28212
rect 34520 28160 34572 28212
rect 37924 28203 37976 28212
rect 37924 28169 37933 28203
rect 37933 28169 37967 28203
rect 37967 28169 37976 28203
rect 37924 28160 37976 28169
rect 21180 27999 21232 28008
rect 14924 27888 14976 27940
rect 21180 27965 21189 27999
rect 21189 27965 21223 27999
rect 21223 27965 21232 27999
rect 21180 27956 21232 27965
rect 23296 27956 23348 28008
rect 24676 27999 24728 28008
rect 20996 27888 21048 27940
rect 21456 27888 21508 27940
rect 22744 27888 22796 27940
rect 24676 27965 24685 27999
rect 24685 27965 24719 27999
rect 24719 27965 24728 27999
rect 24676 27956 24728 27965
rect 25136 27999 25188 28008
rect 25136 27965 25145 27999
rect 25145 27965 25179 27999
rect 25179 27965 25188 27999
rect 25136 27956 25188 27965
rect 26056 27956 26108 28008
rect 26424 27956 26476 28008
rect 26240 27888 26292 27940
rect 14464 27820 14516 27872
rect 15292 27820 15344 27872
rect 17408 27820 17460 27872
rect 20260 27863 20312 27872
rect 20260 27829 20269 27863
rect 20269 27829 20303 27863
rect 20303 27829 20312 27863
rect 20260 27820 20312 27829
rect 21548 27820 21600 27872
rect 29368 27956 29420 28008
rect 30196 27956 30248 28008
rect 30288 27999 30340 28008
rect 30288 27965 30297 27999
rect 30297 27965 30331 27999
rect 30331 27965 30340 27999
rect 30288 27956 30340 27965
rect 30564 27999 30616 28008
rect 30564 27965 30573 27999
rect 30573 27965 30607 27999
rect 30607 27965 30616 27999
rect 32864 27999 32916 28008
rect 30564 27956 30616 27965
rect 32864 27965 32873 27999
rect 32873 27965 32907 27999
rect 32907 27965 32916 27999
rect 32864 27956 32916 27965
rect 28264 27931 28316 27940
rect 28264 27897 28273 27931
rect 28273 27897 28307 27931
rect 28307 27897 28316 27931
rect 28264 27888 28316 27897
rect 27344 27820 27396 27872
rect 33508 27956 33560 28008
rect 36452 28024 36504 28076
rect 37096 28067 37148 28076
rect 37096 28033 37105 28067
rect 37105 28033 37139 28067
rect 37139 28033 37148 28067
rect 37096 28024 37148 28033
rect 35256 27956 35308 28008
rect 35532 27956 35584 28008
rect 36360 27956 36412 28008
rect 36728 27999 36780 28008
rect 36728 27965 36737 27999
rect 36737 27965 36771 27999
rect 36771 27965 36780 27999
rect 36728 27956 36780 27965
rect 37004 27888 37056 27940
rect 19606 27718 19658 27770
rect 19670 27718 19722 27770
rect 19734 27718 19786 27770
rect 19798 27718 19850 27770
rect 4896 27616 4948 27668
rect 5264 27616 5316 27668
rect 11152 27616 11204 27668
rect 14280 27616 14332 27668
rect 15108 27616 15160 27668
rect 30104 27616 30156 27668
rect 36636 27616 36688 27668
rect 6828 27591 6880 27600
rect 6828 27557 6837 27591
rect 6837 27557 6871 27591
rect 6871 27557 6880 27591
rect 6828 27548 6880 27557
rect 8944 27591 8996 27600
rect 8944 27557 8953 27591
rect 8953 27557 8987 27591
rect 8987 27557 8996 27591
rect 8944 27548 8996 27557
rect 2688 27523 2740 27532
rect 2688 27489 2697 27523
rect 2697 27489 2731 27523
rect 2731 27489 2740 27523
rect 2688 27480 2740 27489
rect 3240 27480 3292 27532
rect 4068 27523 4120 27532
rect 4068 27489 4077 27523
rect 4077 27489 4111 27523
rect 4111 27489 4120 27523
rect 4068 27480 4120 27489
rect 4988 27523 5040 27532
rect 4988 27489 4997 27523
rect 4997 27489 5031 27523
rect 5031 27489 5040 27523
rect 4988 27480 5040 27489
rect 5724 27480 5776 27532
rect 7656 27480 7708 27532
rect 8116 27523 8168 27532
rect 1492 27412 1544 27464
rect 3148 27455 3200 27464
rect 3148 27421 3157 27455
rect 3157 27421 3191 27455
rect 3191 27421 3200 27455
rect 3148 27412 3200 27421
rect 4620 27276 4672 27328
rect 6368 27412 6420 27464
rect 8116 27489 8125 27523
rect 8125 27489 8159 27523
rect 8159 27489 8168 27523
rect 8116 27480 8168 27489
rect 8392 27480 8444 27532
rect 10324 27480 10376 27532
rect 12624 27548 12676 27600
rect 20076 27591 20128 27600
rect 20076 27557 20085 27591
rect 20085 27557 20119 27591
rect 20119 27557 20128 27591
rect 20076 27548 20128 27557
rect 20720 27548 20772 27600
rect 11796 27523 11848 27532
rect 7288 27387 7340 27396
rect 7288 27353 7297 27387
rect 7297 27353 7331 27387
rect 7331 27353 7340 27387
rect 7288 27344 7340 27353
rect 7932 27412 7984 27464
rect 11796 27489 11805 27523
rect 11805 27489 11839 27523
rect 11839 27489 11848 27523
rect 11796 27480 11848 27489
rect 12440 27480 12492 27532
rect 11704 27344 11756 27396
rect 13084 27480 13136 27532
rect 13820 27523 13872 27532
rect 13820 27489 13829 27523
rect 13829 27489 13863 27523
rect 13863 27489 13872 27523
rect 13820 27480 13872 27489
rect 14004 27523 14056 27532
rect 14004 27489 14013 27523
rect 14013 27489 14047 27523
rect 14047 27489 14056 27523
rect 14004 27480 14056 27489
rect 14464 27523 14516 27532
rect 14464 27489 14473 27523
rect 14473 27489 14507 27523
rect 14507 27489 14516 27523
rect 14464 27480 14516 27489
rect 14556 27480 14608 27532
rect 15844 27480 15896 27532
rect 16856 27523 16908 27532
rect 16856 27489 16865 27523
rect 16865 27489 16899 27523
rect 16899 27489 16908 27523
rect 16856 27480 16908 27489
rect 18236 27480 18288 27532
rect 19340 27480 19392 27532
rect 19524 27523 19576 27532
rect 19524 27489 19533 27523
rect 19533 27489 19567 27523
rect 19567 27489 19576 27523
rect 19524 27480 19576 27489
rect 19984 27523 20036 27532
rect 19984 27489 19993 27523
rect 19993 27489 20027 27523
rect 20027 27489 20036 27523
rect 19984 27480 20036 27489
rect 20444 27480 20496 27532
rect 22008 27523 22060 27532
rect 22008 27489 22017 27523
rect 22017 27489 22051 27523
rect 22051 27489 22060 27523
rect 22008 27480 22060 27489
rect 22376 27523 22428 27532
rect 22376 27489 22385 27523
rect 22385 27489 22419 27523
rect 22419 27489 22428 27523
rect 22376 27480 22428 27489
rect 22836 27523 22888 27532
rect 22836 27489 22845 27523
rect 22845 27489 22879 27523
rect 22879 27489 22888 27523
rect 22836 27480 22888 27489
rect 23388 27523 23440 27532
rect 23388 27489 23397 27523
rect 23397 27489 23431 27523
rect 23431 27489 23440 27523
rect 23388 27480 23440 27489
rect 23848 27523 23900 27532
rect 23848 27489 23857 27523
rect 23857 27489 23891 27523
rect 23891 27489 23900 27523
rect 23848 27480 23900 27489
rect 24124 27523 24176 27532
rect 24124 27489 24133 27523
rect 24133 27489 24167 27523
rect 24167 27489 24176 27523
rect 24124 27480 24176 27489
rect 24216 27480 24268 27532
rect 14740 27455 14792 27464
rect 14740 27421 14749 27455
rect 14749 27421 14783 27455
rect 14783 27421 14792 27455
rect 14740 27412 14792 27421
rect 8852 27276 8904 27328
rect 9772 27276 9824 27328
rect 22928 27412 22980 27464
rect 23480 27455 23532 27464
rect 23480 27421 23489 27455
rect 23489 27421 23523 27455
rect 23523 27421 23532 27455
rect 23480 27412 23532 27421
rect 15936 27276 15988 27328
rect 19432 27344 19484 27396
rect 20812 27344 20864 27396
rect 21088 27344 21140 27396
rect 26240 27480 26292 27532
rect 26792 27480 26844 27532
rect 27160 27412 27212 27464
rect 27528 27412 27580 27464
rect 28264 27480 28316 27532
rect 30380 27480 30432 27532
rect 31208 27523 31260 27532
rect 31208 27489 31217 27523
rect 31217 27489 31251 27523
rect 31251 27489 31260 27523
rect 31208 27480 31260 27489
rect 33416 27548 33468 27600
rect 34704 27523 34756 27532
rect 28448 27455 28500 27464
rect 26516 27344 26568 27396
rect 27436 27344 27488 27396
rect 28448 27421 28457 27455
rect 28457 27421 28491 27455
rect 28491 27421 28500 27455
rect 28448 27412 28500 27421
rect 32496 27455 32548 27464
rect 32496 27421 32505 27455
rect 32505 27421 32539 27455
rect 32539 27421 32548 27455
rect 32496 27412 32548 27421
rect 34336 27412 34388 27464
rect 34704 27489 34713 27523
rect 34713 27489 34747 27523
rect 34747 27489 34756 27523
rect 34704 27480 34756 27489
rect 36544 27523 36596 27532
rect 36544 27489 36553 27523
rect 36553 27489 36587 27523
rect 36587 27489 36596 27523
rect 36544 27480 36596 27489
rect 37740 27523 37792 27532
rect 30656 27344 30708 27396
rect 32956 27344 33008 27396
rect 37740 27489 37749 27523
rect 37749 27489 37783 27523
rect 37783 27489 37792 27523
rect 37740 27480 37792 27489
rect 19156 27276 19208 27328
rect 19340 27276 19392 27328
rect 20628 27276 20680 27328
rect 22284 27276 22336 27328
rect 23388 27276 23440 27328
rect 29920 27276 29972 27328
rect 33784 27276 33836 27328
rect 35532 27276 35584 27328
rect 37832 27319 37884 27328
rect 37832 27285 37841 27319
rect 37841 27285 37875 27319
rect 37875 27285 37884 27319
rect 37832 27276 37884 27285
rect 4246 27174 4298 27226
rect 4310 27174 4362 27226
rect 4374 27174 4426 27226
rect 4438 27174 4490 27226
rect 34966 27174 35018 27226
rect 35030 27174 35082 27226
rect 35094 27174 35146 27226
rect 35158 27174 35210 27226
rect 1492 27115 1544 27124
rect 1492 27081 1501 27115
rect 1501 27081 1535 27115
rect 1535 27081 1544 27115
rect 1492 27072 1544 27081
rect 1676 27072 1728 27124
rect 4068 27115 4120 27124
rect 4068 27081 4077 27115
rect 4077 27081 4111 27115
rect 4111 27081 4120 27115
rect 4068 27072 4120 27081
rect 4804 27072 4856 27124
rect 8116 27072 8168 27124
rect 14740 27072 14792 27124
rect 22928 27115 22980 27124
rect 1768 26911 1820 26920
rect 1768 26877 1777 26911
rect 1777 26877 1811 26911
rect 1811 26877 1820 26911
rect 1768 26868 1820 26877
rect 2780 26868 2832 26920
rect 3148 26868 3200 26920
rect 4068 26911 4120 26920
rect 4068 26877 4077 26911
rect 4077 26877 4111 26911
rect 4111 26877 4120 26911
rect 4068 26868 4120 26877
rect 4620 26911 4672 26920
rect 4620 26877 4629 26911
rect 4629 26877 4663 26911
rect 4663 26877 4672 26911
rect 4620 26868 4672 26877
rect 4896 26911 4948 26920
rect 4896 26877 4905 26911
rect 4905 26877 4939 26911
rect 4939 26877 4948 26911
rect 4896 26868 4948 26877
rect 4712 26800 4764 26852
rect 7380 26936 7432 26988
rect 8024 26936 8076 26988
rect 8668 26936 8720 26988
rect 9220 26979 9272 26988
rect 6920 26868 6972 26920
rect 7196 26911 7248 26920
rect 7196 26877 7205 26911
rect 7205 26877 7239 26911
rect 7239 26877 7248 26911
rect 7196 26868 7248 26877
rect 7932 26911 7984 26920
rect 7932 26877 7941 26911
rect 7941 26877 7975 26911
rect 7975 26877 7984 26911
rect 7932 26868 7984 26877
rect 9220 26945 9229 26979
rect 9229 26945 9263 26979
rect 9263 26945 9272 26979
rect 9220 26936 9272 26945
rect 9312 26936 9364 26988
rect 9680 26868 9732 26920
rect 11244 26868 11296 26920
rect 6000 26800 6052 26852
rect 7380 26775 7432 26784
rect 7380 26741 7389 26775
rect 7389 26741 7423 26775
rect 7423 26741 7432 26775
rect 7380 26732 7432 26741
rect 7472 26732 7524 26784
rect 10324 26800 10376 26852
rect 11152 26732 11204 26784
rect 11796 27004 11848 27056
rect 11704 26911 11756 26920
rect 11704 26877 11713 26911
rect 11713 26877 11747 26911
rect 11747 26877 11756 26911
rect 11704 26868 11756 26877
rect 12716 27004 12768 27056
rect 13820 27004 13872 27056
rect 17224 27004 17276 27056
rect 17684 27004 17736 27056
rect 12532 26868 12584 26920
rect 12992 26868 13044 26920
rect 13084 26868 13136 26920
rect 15844 26936 15896 26988
rect 17592 26936 17644 26988
rect 20720 27004 20772 27056
rect 22928 27081 22937 27115
rect 22937 27081 22971 27115
rect 22971 27081 22980 27115
rect 22928 27072 22980 27081
rect 23388 27004 23440 27056
rect 24124 27004 24176 27056
rect 24952 27072 25004 27124
rect 32036 27072 32088 27124
rect 33784 27115 33836 27124
rect 33784 27081 33793 27115
rect 33793 27081 33827 27115
rect 33827 27081 33836 27115
rect 33784 27072 33836 27081
rect 25320 27004 25372 27056
rect 28448 27047 28500 27056
rect 28448 27013 28457 27047
rect 28457 27013 28491 27047
rect 28491 27013 28500 27047
rect 28448 27004 28500 27013
rect 30288 27004 30340 27056
rect 15108 26868 15160 26920
rect 16396 26911 16448 26920
rect 15568 26800 15620 26852
rect 16396 26877 16405 26911
rect 16405 26877 16439 26911
rect 16439 26877 16448 26911
rect 16396 26868 16448 26877
rect 16580 26911 16632 26920
rect 16580 26877 16589 26911
rect 16589 26877 16623 26911
rect 16623 26877 16632 26911
rect 16580 26868 16632 26877
rect 16948 26800 17000 26852
rect 14372 26732 14424 26784
rect 17776 26732 17828 26784
rect 18972 26868 19024 26920
rect 19340 26936 19392 26988
rect 21180 26936 21232 26988
rect 22100 26936 22152 26988
rect 19524 26868 19576 26920
rect 19892 26868 19944 26920
rect 20444 26868 20496 26920
rect 20628 26868 20680 26920
rect 20996 26911 21048 26920
rect 20996 26877 21005 26911
rect 21005 26877 21039 26911
rect 21039 26877 21048 26911
rect 20996 26868 21048 26877
rect 21088 26868 21140 26920
rect 23572 26868 23624 26920
rect 24768 26868 24820 26920
rect 25596 26911 25648 26920
rect 25596 26877 25605 26911
rect 25605 26877 25639 26911
rect 25639 26877 25648 26911
rect 25596 26868 25648 26877
rect 25872 26911 25924 26920
rect 25872 26877 25881 26911
rect 25881 26877 25915 26911
rect 25915 26877 25924 26911
rect 25872 26868 25924 26877
rect 26056 26868 26108 26920
rect 27528 26868 27580 26920
rect 28448 26911 28500 26920
rect 28448 26877 28457 26911
rect 28457 26877 28491 26911
rect 28491 26877 28500 26911
rect 28448 26868 28500 26877
rect 29092 26868 29144 26920
rect 29920 26911 29972 26920
rect 29920 26877 29929 26911
rect 29929 26877 29963 26911
rect 29963 26877 29972 26911
rect 29920 26868 29972 26877
rect 30380 26911 30432 26920
rect 30380 26877 30389 26911
rect 30389 26877 30423 26911
rect 30423 26877 30432 26911
rect 30380 26868 30432 26877
rect 32772 26936 32824 26988
rect 34336 26936 34388 26988
rect 19984 26800 20036 26852
rect 18328 26775 18380 26784
rect 18328 26741 18337 26775
rect 18337 26741 18371 26775
rect 18371 26741 18380 26775
rect 18328 26732 18380 26741
rect 19156 26732 19208 26784
rect 23664 26800 23716 26852
rect 23848 26843 23900 26852
rect 23848 26809 23857 26843
rect 23857 26809 23891 26843
rect 23891 26809 23900 26843
rect 23848 26800 23900 26809
rect 24492 26800 24544 26852
rect 22008 26732 22060 26784
rect 22744 26732 22796 26784
rect 27988 26732 28040 26784
rect 32312 26868 32364 26920
rect 32680 26911 32732 26920
rect 32680 26877 32689 26911
rect 32689 26877 32723 26911
rect 32723 26877 32732 26911
rect 32680 26868 32732 26877
rect 34612 26868 34664 26920
rect 35716 26911 35768 26920
rect 32220 26800 32272 26852
rect 31116 26732 31168 26784
rect 35716 26877 35725 26911
rect 35725 26877 35759 26911
rect 35759 26877 35768 26911
rect 35716 26868 35768 26877
rect 36360 26868 36412 26920
rect 37832 26936 37884 26988
rect 37004 26868 37056 26920
rect 35992 26843 36044 26852
rect 35992 26809 36001 26843
rect 36001 26809 36035 26843
rect 36035 26809 36044 26843
rect 35992 26800 36044 26809
rect 36820 26732 36872 26784
rect 37004 26732 37056 26784
rect 19606 26630 19658 26682
rect 19670 26630 19722 26682
rect 19734 26630 19786 26682
rect 19798 26630 19850 26682
rect 1400 26435 1452 26444
rect 1400 26401 1409 26435
rect 1409 26401 1443 26435
rect 1443 26401 1452 26435
rect 1400 26392 1452 26401
rect 1676 26435 1728 26444
rect 1676 26401 1685 26435
rect 1685 26401 1719 26435
rect 1719 26401 1728 26435
rect 1676 26392 1728 26401
rect 4804 26435 4856 26444
rect 4804 26401 4813 26435
rect 4813 26401 4847 26435
rect 4847 26401 4856 26435
rect 4804 26392 4856 26401
rect 7196 26435 7248 26444
rect 7196 26401 7205 26435
rect 7205 26401 7239 26435
rect 7239 26401 7248 26435
rect 7196 26392 7248 26401
rect 8576 26435 8628 26444
rect 8576 26401 8585 26435
rect 8585 26401 8619 26435
rect 8619 26401 8628 26435
rect 8576 26392 8628 26401
rect 8760 26435 8812 26444
rect 8760 26401 8769 26435
rect 8769 26401 8803 26435
rect 8803 26401 8812 26435
rect 8760 26392 8812 26401
rect 8852 26392 8904 26444
rect 12440 26528 12492 26580
rect 12624 26528 12676 26580
rect 11152 26460 11204 26512
rect 4528 26367 4580 26376
rect 2688 26256 2740 26308
rect 4528 26333 4537 26367
rect 4537 26333 4571 26367
rect 4571 26333 4580 26367
rect 4528 26324 4580 26333
rect 4712 26324 4764 26376
rect 10784 26392 10836 26444
rect 11704 26435 11756 26444
rect 11704 26401 11713 26435
rect 11713 26401 11747 26435
rect 11747 26401 11756 26435
rect 11704 26392 11756 26401
rect 11888 26460 11940 26512
rect 16580 26528 16632 26580
rect 19984 26528 20036 26580
rect 20260 26528 20312 26580
rect 22376 26528 22428 26580
rect 23112 26528 23164 26580
rect 26056 26528 26108 26580
rect 29644 26528 29696 26580
rect 32680 26528 32732 26580
rect 12532 26435 12584 26444
rect 12532 26401 12541 26435
rect 12541 26401 12575 26435
rect 12575 26401 12584 26435
rect 12532 26392 12584 26401
rect 12992 26435 13044 26444
rect 12992 26401 13001 26435
rect 13001 26401 13035 26435
rect 13035 26401 13044 26435
rect 12992 26392 13044 26401
rect 13820 26392 13872 26444
rect 13084 26367 13136 26376
rect 8392 26299 8444 26308
rect 8392 26265 8401 26299
rect 8401 26265 8435 26299
rect 8435 26265 8444 26299
rect 8392 26256 8444 26265
rect 13084 26333 13093 26367
rect 13093 26333 13127 26367
rect 13127 26333 13136 26367
rect 13084 26324 13136 26333
rect 14280 26367 14332 26376
rect 14280 26333 14289 26367
rect 14289 26333 14323 26367
rect 14323 26333 14332 26367
rect 14280 26324 14332 26333
rect 15844 26392 15896 26444
rect 16120 26435 16172 26444
rect 16120 26401 16129 26435
rect 16129 26401 16163 26435
rect 16163 26401 16172 26435
rect 16120 26392 16172 26401
rect 16764 26460 16816 26512
rect 17592 26435 17644 26444
rect 17592 26401 17601 26435
rect 17601 26401 17635 26435
rect 17635 26401 17644 26435
rect 17592 26392 17644 26401
rect 18052 26392 18104 26444
rect 19340 26460 19392 26512
rect 19708 26460 19760 26512
rect 21548 26460 21600 26512
rect 22836 26460 22888 26512
rect 18972 26392 19024 26444
rect 19892 26392 19944 26444
rect 19984 26435 20036 26444
rect 19984 26401 19993 26435
rect 19993 26401 20027 26435
rect 20027 26401 20036 26435
rect 19984 26392 20036 26401
rect 20628 26392 20680 26444
rect 15108 26324 15160 26376
rect 16488 26324 16540 26376
rect 17408 26324 17460 26376
rect 17316 26256 17368 26308
rect 18420 26256 18472 26308
rect 21088 26435 21140 26444
rect 21088 26401 21097 26435
rect 21097 26401 21131 26435
rect 21131 26401 21140 26435
rect 21088 26392 21140 26401
rect 21456 26392 21508 26444
rect 22284 26435 22336 26444
rect 22284 26401 22293 26435
rect 22293 26401 22327 26435
rect 22327 26401 22336 26435
rect 22284 26392 22336 26401
rect 22744 26435 22796 26444
rect 22744 26401 22753 26435
rect 22753 26401 22787 26435
rect 22787 26401 22796 26435
rect 22744 26392 22796 26401
rect 23388 26392 23440 26444
rect 23572 26435 23624 26444
rect 23572 26401 23581 26435
rect 23581 26401 23615 26435
rect 23615 26401 23624 26435
rect 23572 26392 23624 26401
rect 25136 26460 25188 26512
rect 25320 26460 25372 26512
rect 24584 26392 24636 26444
rect 26792 26435 26844 26444
rect 26792 26401 26801 26435
rect 26801 26401 26835 26435
rect 26835 26401 26844 26435
rect 26792 26392 26844 26401
rect 29000 26460 29052 26512
rect 27620 26392 27672 26444
rect 29920 26460 29972 26512
rect 33048 26460 33100 26512
rect 29644 26435 29696 26444
rect 29644 26401 29653 26435
rect 29653 26401 29687 26435
rect 29687 26401 29696 26435
rect 29644 26392 29696 26401
rect 31024 26392 31076 26444
rect 32036 26392 32088 26444
rect 32220 26435 32272 26444
rect 32220 26401 32229 26435
rect 32229 26401 32263 26435
rect 32263 26401 32272 26435
rect 32220 26392 32272 26401
rect 32956 26435 33008 26444
rect 32956 26401 32965 26435
rect 32965 26401 32999 26435
rect 32999 26401 33008 26435
rect 32956 26392 33008 26401
rect 23664 26324 23716 26376
rect 24768 26324 24820 26376
rect 29276 26324 29328 26376
rect 30748 26324 30800 26376
rect 31484 26324 31536 26376
rect 34704 26392 34756 26444
rect 35348 26392 35400 26444
rect 35992 26392 36044 26444
rect 36820 26435 36872 26444
rect 36820 26401 36829 26435
rect 36829 26401 36863 26435
rect 36863 26401 36872 26435
rect 36820 26392 36872 26401
rect 37004 26435 37056 26444
rect 37004 26401 37013 26435
rect 37013 26401 37047 26435
rect 37047 26401 37056 26435
rect 37004 26392 37056 26401
rect 34796 26324 34848 26376
rect 21088 26256 21140 26308
rect 21272 26256 21324 26308
rect 22008 26256 22060 26308
rect 22652 26256 22704 26308
rect 22928 26256 22980 26308
rect 28172 26256 28224 26308
rect 28448 26256 28500 26308
rect 30656 26299 30708 26308
rect 30656 26265 30665 26299
rect 30665 26265 30699 26299
rect 30699 26265 30708 26299
rect 30656 26256 30708 26265
rect 37740 26256 37792 26308
rect 4804 26188 4856 26240
rect 4896 26188 4948 26240
rect 6460 26188 6512 26240
rect 9864 26188 9916 26240
rect 13084 26188 13136 26240
rect 17592 26188 17644 26240
rect 18236 26188 18288 26240
rect 20996 26188 21048 26240
rect 22192 26231 22244 26240
rect 22192 26197 22201 26231
rect 22201 26197 22235 26231
rect 22235 26197 22244 26231
rect 22192 26188 22244 26197
rect 33968 26231 34020 26240
rect 33968 26197 33977 26231
rect 33977 26197 34011 26231
rect 34011 26197 34020 26231
rect 33968 26188 34020 26197
rect 34612 26231 34664 26240
rect 34612 26197 34621 26231
rect 34621 26197 34655 26231
rect 34655 26197 34664 26231
rect 34612 26188 34664 26197
rect 4246 26086 4298 26138
rect 4310 26086 4362 26138
rect 4374 26086 4426 26138
rect 4438 26086 4490 26138
rect 34966 26086 35018 26138
rect 35030 26086 35082 26138
rect 35094 26086 35146 26138
rect 35158 26086 35210 26138
rect 3976 25984 4028 26036
rect 12624 25984 12676 26036
rect 18328 25984 18380 26036
rect 21456 25984 21508 26036
rect 1860 25916 1912 25968
rect 7748 25959 7800 25968
rect 7748 25925 7757 25959
rect 7757 25925 7791 25959
rect 7791 25925 7800 25959
rect 7748 25916 7800 25925
rect 15384 25959 15436 25968
rect 15384 25925 15393 25959
rect 15393 25925 15427 25959
rect 15427 25925 15436 25959
rect 15384 25916 15436 25925
rect 17776 25916 17828 25968
rect 1768 25848 1820 25900
rect 4620 25891 4672 25900
rect 4620 25857 4629 25891
rect 4629 25857 4663 25891
rect 4663 25857 4672 25891
rect 4620 25848 4672 25857
rect 8576 25848 8628 25900
rect 2688 25823 2740 25832
rect 2688 25789 2697 25823
rect 2697 25789 2731 25823
rect 2731 25789 2740 25823
rect 2688 25780 2740 25789
rect 3148 25823 3200 25832
rect 3148 25789 3157 25823
rect 3157 25789 3191 25823
rect 3191 25789 3200 25823
rect 3148 25780 3200 25789
rect 3240 25823 3292 25832
rect 3240 25789 3249 25823
rect 3249 25789 3283 25823
rect 3283 25789 3292 25823
rect 3240 25780 3292 25789
rect 3976 25780 4028 25832
rect 4712 25780 4764 25832
rect 5172 25823 5224 25832
rect 5172 25789 5181 25823
rect 5181 25789 5215 25823
rect 5215 25789 5224 25823
rect 5172 25780 5224 25789
rect 5632 25780 5684 25832
rect 7012 25780 7064 25832
rect 7932 25823 7984 25832
rect 7932 25789 7941 25823
rect 7941 25789 7975 25823
rect 7975 25789 7984 25823
rect 7932 25780 7984 25789
rect 8392 25823 8444 25832
rect 8392 25789 8401 25823
rect 8401 25789 8435 25823
rect 8435 25789 8444 25823
rect 8392 25780 8444 25789
rect 8852 25823 8904 25832
rect 8852 25789 8861 25823
rect 8861 25789 8895 25823
rect 8895 25789 8904 25823
rect 8852 25780 8904 25789
rect 12532 25848 12584 25900
rect 13544 25848 13596 25900
rect 14648 25891 14700 25900
rect 14648 25857 14657 25891
rect 14657 25857 14691 25891
rect 14691 25857 14700 25891
rect 14648 25848 14700 25857
rect 16948 25848 17000 25900
rect 18236 25848 18288 25900
rect 8760 25712 8812 25764
rect 9864 25780 9916 25832
rect 13820 25780 13872 25832
rect 14372 25823 14424 25832
rect 11244 25755 11296 25764
rect 6000 25687 6052 25696
rect 6000 25653 6009 25687
rect 6009 25653 6043 25687
rect 6043 25653 6052 25687
rect 6000 25644 6052 25653
rect 8392 25644 8444 25696
rect 11244 25721 11253 25755
rect 11253 25721 11287 25755
rect 11287 25721 11296 25755
rect 11244 25712 11296 25721
rect 11612 25755 11664 25764
rect 11612 25721 11621 25755
rect 11621 25721 11655 25755
rect 11655 25721 11664 25755
rect 11612 25712 11664 25721
rect 13452 25712 13504 25764
rect 14372 25789 14381 25823
rect 14381 25789 14415 25823
rect 14415 25789 14424 25823
rect 14372 25780 14424 25789
rect 11060 25687 11112 25696
rect 11060 25653 11069 25687
rect 11069 25653 11103 25687
rect 11103 25653 11112 25687
rect 11060 25644 11112 25653
rect 11152 25687 11204 25696
rect 11152 25653 11161 25687
rect 11161 25653 11195 25687
rect 11195 25653 11204 25687
rect 11152 25644 11204 25653
rect 11888 25644 11940 25696
rect 15660 25780 15712 25832
rect 16120 25780 16172 25832
rect 18420 25780 18472 25832
rect 18604 25848 18656 25900
rect 19984 25848 20036 25900
rect 19892 25823 19944 25832
rect 17408 25712 17460 25764
rect 17960 25712 18012 25764
rect 15844 25644 15896 25696
rect 16856 25644 16908 25696
rect 19892 25789 19901 25823
rect 19901 25789 19935 25823
rect 19935 25789 19944 25823
rect 19892 25780 19944 25789
rect 20260 25823 20312 25832
rect 20260 25789 20269 25823
rect 20269 25789 20303 25823
rect 20303 25789 20312 25823
rect 20260 25780 20312 25789
rect 21272 25848 21324 25900
rect 22192 25891 22244 25900
rect 22192 25857 22201 25891
rect 22201 25857 22235 25891
rect 22235 25857 22244 25891
rect 22192 25848 22244 25857
rect 20904 25823 20956 25832
rect 20904 25789 20913 25823
rect 20913 25789 20947 25823
rect 20947 25789 20956 25823
rect 20904 25780 20956 25789
rect 20996 25780 21048 25832
rect 23756 25984 23808 26036
rect 25044 25984 25096 26036
rect 25688 25984 25740 26036
rect 32036 25984 32088 26036
rect 34428 25984 34480 26036
rect 35348 26027 35400 26036
rect 35348 25993 35357 26027
rect 35357 25993 35391 26027
rect 35391 25993 35400 26027
rect 35348 25984 35400 25993
rect 26424 25916 26476 25968
rect 23664 25823 23716 25832
rect 23664 25789 23673 25823
rect 23673 25789 23707 25823
rect 23707 25789 23716 25823
rect 23664 25780 23716 25789
rect 23020 25644 23072 25696
rect 24400 25823 24452 25832
rect 24400 25789 24409 25823
rect 24409 25789 24443 25823
rect 24443 25789 24452 25823
rect 24400 25780 24452 25789
rect 24676 25823 24728 25832
rect 24676 25789 24685 25823
rect 24685 25789 24719 25823
rect 24719 25789 24728 25823
rect 24676 25780 24728 25789
rect 24768 25780 24820 25832
rect 26516 25780 26568 25832
rect 27988 25848 28040 25900
rect 30288 25848 30340 25900
rect 30656 25891 30708 25900
rect 30656 25857 30665 25891
rect 30665 25857 30699 25891
rect 30699 25857 30708 25891
rect 30656 25848 30708 25857
rect 31760 25848 31812 25900
rect 29276 25780 29328 25832
rect 32496 25823 32548 25832
rect 32496 25789 32505 25823
rect 32505 25789 32539 25823
rect 32539 25789 32548 25823
rect 32496 25780 32548 25789
rect 33968 25848 34020 25900
rect 34520 25848 34572 25900
rect 33416 25823 33468 25832
rect 33416 25789 33425 25823
rect 33425 25789 33459 25823
rect 33459 25789 33468 25823
rect 33416 25780 33468 25789
rect 34612 25780 34664 25832
rect 35532 25823 35584 25832
rect 35532 25789 35541 25823
rect 35541 25789 35575 25823
rect 35575 25789 35584 25823
rect 35532 25780 35584 25789
rect 24492 25644 24544 25696
rect 31116 25644 31168 25696
rect 36360 25780 36412 25832
rect 36544 25644 36596 25696
rect 19606 25542 19658 25594
rect 19670 25542 19722 25594
rect 19734 25542 19786 25594
rect 19798 25542 19850 25594
rect 3240 25440 3292 25492
rect 7012 25440 7064 25492
rect 11152 25440 11204 25492
rect 11244 25372 11296 25424
rect 1400 25347 1452 25356
rect 1400 25313 1409 25347
rect 1409 25313 1443 25347
rect 1443 25313 1452 25347
rect 1400 25304 1452 25313
rect 2688 25304 2740 25356
rect 4068 25347 4120 25356
rect 4068 25313 4077 25347
rect 4077 25313 4111 25347
rect 4111 25313 4120 25347
rect 4068 25304 4120 25313
rect 5632 25347 5684 25356
rect 1676 25279 1728 25288
rect 1676 25245 1685 25279
rect 1685 25245 1719 25279
rect 1719 25245 1728 25279
rect 1676 25236 1728 25245
rect 5632 25313 5641 25347
rect 5641 25313 5675 25347
rect 5675 25313 5684 25347
rect 5632 25304 5684 25313
rect 7012 25304 7064 25356
rect 11612 25304 11664 25356
rect 5540 25236 5592 25288
rect 4712 25168 4764 25220
rect 7196 25236 7248 25288
rect 9680 25279 9732 25288
rect 9680 25245 9689 25279
rect 9689 25245 9723 25279
rect 9723 25245 9732 25279
rect 9956 25279 10008 25288
rect 9680 25236 9732 25245
rect 9956 25245 9965 25279
rect 9965 25245 9999 25279
rect 9999 25245 10008 25279
rect 9956 25236 10008 25245
rect 15660 25440 15712 25492
rect 15844 25483 15896 25492
rect 15844 25449 15853 25483
rect 15853 25449 15887 25483
rect 15887 25449 15896 25483
rect 15844 25440 15896 25449
rect 12624 25347 12676 25356
rect 12624 25313 12633 25347
rect 12633 25313 12667 25347
rect 12667 25313 12676 25347
rect 12624 25304 12676 25313
rect 15200 25304 15252 25356
rect 16028 25372 16080 25424
rect 16856 25347 16908 25356
rect 16856 25313 16865 25347
rect 16865 25313 16899 25347
rect 16899 25313 16908 25347
rect 16856 25304 16908 25313
rect 18052 25440 18104 25492
rect 17316 25304 17368 25356
rect 17960 25304 18012 25356
rect 21272 25304 21324 25356
rect 22284 25440 22336 25492
rect 22008 25347 22060 25356
rect 22008 25313 22017 25347
rect 22017 25313 22051 25347
rect 22051 25313 22060 25347
rect 22008 25304 22060 25313
rect 3148 25100 3200 25152
rect 6828 25100 6880 25152
rect 8576 25100 8628 25152
rect 16672 25211 16724 25220
rect 16672 25177 16681 25211
rect 16681 25177 16715 25211
rect 16715 25177 16724 25211
rect 16672 25168 16724 25177
rect 19432 25236 19484 25288
rect 19892 25279 19944 25288
rect 19892 25245 19901 25279
rect 19901 25245 19935 25279
rect 19935 25245 19944 25279
rect 19892 25236 19944 25245
rect 22744 25372 22796 25424
rect 23112 25347 23164 25356
rect 21824 25168 21876 25220
rect 23112 25313 23121 25347
rect 23121 25313 23155 25347
rect 23155 25313 23164 25347
rect 23112 25304 23164 25313
rect 23664 25236 23716 25288
rect 11060 25100 11112 25152
rect 11612 25100 11664 25152
rect 11980 25143 12032 25152
rect 11980 25109 11989 25143
rect 11989 25109 12023 25143
rect 12023 25109 12032 25143
rect 11980 25100 12032 25109
rect 13544 25100 13596 25152
rect 14924 25100 14976 25152
rect 15568 25100 15620 25152
rect 16856 25100 16908 25152
rect 17592 25100 17644 25152
rect 21640 25100 21692 25152
rect 22008 25100 22060 25152
rect 24768 25372 24820 25424
rect 24032 25347 24084 25356
rect 24032 25313 24041 25347
rect 24041 25313 24075 25347
rect 24075 25313 24084 25347
rect 24032 25304 24084 25313
rect 24492 25304 24544 25356
rect 35440 25440 35492 25492
rect 35624 25440 35676 25492
rect 26424 25372 26476 25424
rect 26148 25304 26200 25356
rect 29920 25372 29972 25424
rect 28172 25347 28224 25356
rect 28172 25313 28181 25347
rect 28181 25313 28215 25347
rect 28215 25313 28224 25347
rect 28172 25304 28224 25313
rect 30564 25347 30616 25356
rect 30564 25313 30573 25347
rect 30573 25313 30607 25347
rect 30607 25313 30616 25347
rect 30564 25304 30616 25313
rect 30748 25347 30800 25356
rect 30748 25313 30757 25347
rect 30757 25313 30791 25347
rect 30791 25313 30800 25347
rect 30748 25304 30800 25313
rect 32772 25347 32824 25356
rect 24308 25211 24360 25220
rect 24308 25177 24317 25211
rect 24317 25177 24351 25211
rect 24351 25177 24360 25211
rect 24308 25168 24360 25177
rect 27620 25236 27672 25288
rect 24492 25168 24544 25220
rect 26516 25168 26568 25220
rect 27436 25168 27488 25220
rect 29828 25236 29880 25288
rect 32772 25313 32781 25347
rect 32781 25313 32815 25347
rect 32815 25313 32824 25347
rect 32772 25304 32824 25313
rect 33968 25304 34020 25356
rect 37372 25304 37424 25356
rect 31208 25236 31260 25288
rect 32956 25236 33008 25288
rect 34336 25236 34388 25288
rect 35716 25236 35768 25288
rect 25412 25100 25464 25152
rect 31944 25100 31996 25152
rect 33784 25100 33836 25152
rect 35532 25100 35584 25152
rect 36544 25100 36596 25152
rect 4246 24998 4298 25050
rect 4310 24998 4362 25050
rect 4374 24998 4426 25050
rect 4438 24998 4490 25050
rect 34966 24998 35018 25050
rect 35030 24998 35082 25050
rect 35094 24998 35146 25050
rect 35158 24998 35210 25050
rect 9772 24896 9824 24948
rect 12624 24896 12676 24948
rect 8668 24828 8720 24880
rect 3240 24760 3292 24812
rect 4068 24760 4120 24812
rect 5540 24803 5592 24812
rect 5540 24769 5549 24803
rect 5549 24769 5583 24803
rect 5583 24769 5592 24803
rect 5540 24760 5592 24769
rect 7196 24803 7248 24812
rect 7196 24769 7205 24803
rect 7205 24769 7239 24803
rect 7239 24769 7248 24803
rect 7196 24760 7248 24769
rect 7748 24803 7800 24812
rect 7748 24769 7757 24803
rect 7757 24769 7791 24803
rect 7791 24769 7800 24803
rect 7748 24760 7800 24769
rect 8392 24760 8444 24812
rect 11980 24828 12032 24880
rect 1860 24735 1912 24744
rect 1860 24701 1869 24735
rect 1869 24701 1903 24735
rect 1903 24701 1912 24735
rect 1860 24692 1912 24701
rect 2688 24692 2740 24744
rect 5448 24692 5500 24744
rect 6920 24692 6972 24744
rect 9220 24735 9272 24744
rect 9220 24701 9229 24735
rect 9229 24701 9263 24735
rect 9263 24701 9272 24735
rect 9220 24692 9272 24701
rect 7104 24624 7156 24676
rect 9496 24624 9548 24676
rect 6828 24556 6880 24608
rect 10048 24692 10100 24744
rect 10784 24692 10836 24744
rect 12440 24803 12492 24812
rect 12440 24769 12449 24803
rect 12449 24769 12483 24803
rect 12483 24769 12492 24803
rect 12440 24760 12492 24769
rect 13544 24760 13596 24812
rect 19432 24896 19484 24948
rect 22284 24896 22336 24948
rect 25044 24896 25096 24948
rect 27804 24896 27856 24948
rect 36268 24896 36320 24948
rect 38016 24896 38068 24948
rect 18052 24828 18104 24880
rect 18972 24828 19024 24880
rect 20076 24871 20128 24880
rect 20076 24837 20085 24871
rect 20085 24837 20119 24871
rect 20119 24837 20128 24871
rect 20076 24828 20128 24837
rect 21088 24803 21140 24812
rect 11612 24735 11664 24744
rect 11612 24701 11621 24735
rect 11621 24701 11655 24735
rect 11655 24701 11664 24735
rect 11612 24692 11664 24701
rect 12072 24692 12124 24744
rect 10692 24624 10744 24676
rect 14280 24692 14332 24744
rect 14648 24692 14700 24744
rect 14924 24735 14976 24744
rect 14924 24701 14933 24735
rect 14933 24701 14967 24735
rect 14967 24701 14976 24735
rect 14924 24692 14976 24701
rect 15660 24735 15712 24744
rect 15660 24701 15669 24735
rect 15669 24701 15703 24735
rect 15703 24701 15712 24735
rect 15660 24692 15712 24701
rect 16672 24692 16724 24744
rect 17132 24735 17184 24744
rect 17132 24701 17141 24735
rect 17141 24701 17175 24735
rect 17175 24701 17184 24735
rect 17132 24692 17184 24701
rect 16212 24624 16264 24676
rect 18788 24735 18840 24744
rect 18144 24667 18196 24676
rect 18144 24633 18153 24667
rect 18153 24633 18187 24667
rect 18187 24633 18196 24667
rect 18144 24624 18196 24633
rect 18788 24701 18797 24735
rect 18797 24701 18831 24735
rect 18831 24701 18840 24735
rect 18788 24692 18840 24701
rect 18972 24735 19024 24744
rect 18972 24701 18981 24735
rect 18981 24701 19015 24735
rect 19015 24701 19024 24735
rect 18972 24692 19024 24701
rect 19892 24735 19944 24744
rect 19892 24701 19901 24735
rect 19901 24701 19935 24735
rect 19935 24701 19944 24735
rect 19892 24692 19944 24701
rect 21088 24769 21097 24803
rect 21097 24769 21131 24803
rect 21131 24769 21140 24803
rect 21088 24760 21140 24769
rect 21272 24735 21324 24744
rect 21272 24701 21281 24735
rect 21281 24701 21315 24735
rect 21315 24701 21324 24735
rect 21640 24735 21692 24744
rect 21272 24692 21324 24701
rect 21640 24701 21649 24735
rect 21649 24701 21683 24735
rect 21683 24701 21692 24735
rect 21640 24692 21692 24701
rect 21824 24735 21876 24744
rect 21824 24701 21833 24735
rect 21833 24701 21867 24735
rect 21867 24701 21876 24735
rect 21824 24692 21876 24701
rect 19340 24624 19392 24676
rect 23664 24828 23716 24880
rect 25596 24828 25648 24880
rect 29092 24828 29144 24880
rect 22744 24760 22796 24812
rect 28264 24760 28316 24812
rect 31944 24760 31996 24812
rect 22652 24735 22704 24744
rect 22652 24701 22661 24735
rect 22661 24701 22695 24735
rect 22695 24701 22704 24735
rect 22652 24692 22704 24701
rect 23664 24735 23716 24744
rect 23664 24701 23673 24735
rect 23673 24701 23707 24735
rect 23707 24701 23716 24735
rect 23664 24692 23716 24701
rect 24216 24692 24268 24744
rect 24952 24735 25004 24744
rect 24952 24701 24961 24735
rect 24961 24701 24995 24735
rect 24995 24701 25004 24735
rect 24952 24692 25004 24701
rect 25412 24735 25464 24744
rect 25412 24701 25421 24735
rect 25421 24701 25455 24735
rect 25455 24701 25464 24735
rect 25412 24692 25464 24701
rect 26148 24735 26200 24744
rect 26148 24701 26157 24735
rect 26157 24701 26191 24735
rect 26191 24701 26200 24735
rect 26148 24692 26200 24701
rect 27712 24735 27764 24744
rect 27712 24701 27721 24735
rect 27721 24701 27755 24735
rect 27755 24701 27764 24735
rect 27712 24692 27764 24701
rect 28080 24735 28132 24744
rect 28080 24701 28089 24735
rect 28089 24701 28123 24735
rect 28123 24701 28132 24735
rect 28080 24692 28132 24701
rect 29276 24735 29328 24744
rect 29276 24701 29285 24735
rect 29285 24701 29319 24735
rect 29319 24701 29328 24735
rect 29276 24692 29328 24701
rect 29828 24735 29880 24744
rect 29828 24701 29837 24735
rect 29837 24701 29871 24735
rect 29871 24701 29880 24735
rect 29828 24692 29880 24701
rect 30472 24735 30524 24744
rect 30472 24701 30481 24735
rect 30481 24701 30515 24735
rect 30515 24701 30524 24735
rect 30472 24692 30524 24701
rect 31392 24735 31444 24744
rect 31392 24701 31401 24735
rect 31401 24701 31435 24735
rect 31435 24701 31444 24735
rect 31392 24692 31444 24701
rect 32036 24735 32088 24744
rect 32036 24701 32045 24735
rect 32045 24701 32079 24735
rect 32079 24701 32088 24735
rect 32036 24692 32088 24701
rect 33048 24692 33100 24744
rect 33968 24760 34020 24812
rect 34520 24760 34572 24812
rect 34612 24760 34664 24812
rect 11704 24556 11756 24608
rect 14924 24556 14976 24608
rect 15568 24556 15620 24608
rect 32588 24624 32640 24676
rect 33600 24667 33652 24676
rect 33600 24633 33609 24667
rect 33609 24633 33643 24667
rect 33643 24633 33652 24667
rect 33600 24624 33652 24633
rect 33968 24667 34020 24676
rect 33968 24633 33977 24667
rect 33977 24633 34011 24667
rect 34011 24633 34020 24667
rect 33968 24624 34020 24633
rect 34336 24624 34388 24676
rect 36084 24692 36136 24744
rect 36360 24692 36412 24744
rect 37188 24735 37240 24744
rect 37188 24701 37197 24735
rect 37197 24701 37231 24735
rect 37231 24701 37240 24735
rect 37188 24692 37240 24701
rect 37832 24692 37884 24744
rect 38016 24624 38068 24676
rect 22468 24556 22520 24608
rect 23572 24556 23624 24608
rect 24400 24556 24452 24608
rect 24676 24556 24728 24608
rect 29000 24556 29052 24608
rect 30656 24556 30708 24608
rect 31484 24556 31536 24608
rect 32312 24556 32364 24608
rect 32864 24556 32916 24608
rect 36820 24556 36872 24608
rect 19606 24454 19658 24506
rect 19670 24454 19722 24506
rect 19734 24454 19786 24506
rect 19798 24454 19850 24506
rect 16212 24352 16264 24404
rect 2228 24216 2280 24268
rect 4896 24284 4948 24336
rect 7012 24284 7064 24336
rect 8392 24284 8444 24336
rect 8760 24327 8812 24336
rect 8760 24293 8769 24327
rect 8769 24293 8803 24327
rect 8803 24293 8812 24327
rect 8760 24284 8812 24293
rect 2872 24216 2924 24268
rect 3240 24216 3292 24268
rect 6000 24216 6052 24268
rect 7104 24216 7156 24268
rect 7748 24259 7800 24268
rect 2780 24148 2832 24200
rect 3148 24191 3200 24200
rect 3148 24157 3157 24191
rect 3157 24157 3191 24191
rect 3191 24157 3200 24191
rect 3148 24148 3200 24157
rect 4712 24148 4764 24200
rect 7472 24191 7524 24200
rect 7472 24157 7481 24191
rect 7481 24157 7515 24191
rect 7515 24157 7524 24191
rect 7472 24148 7524 24157
rect 7748 24225 7757 24259
rect 7757 24225 7791 24259
rect 7791 24225 7800 24259
rect 7748 24216 7800 24225
rect 8668 24259 8720 24268
rect 8668 24225 8677 24259
rect 8677 24225 8711 24259
rect 8711 24225 8720 24259
rect 8668 24216 8720 24225
rect 9128 24259 9180 24268
rect 9128 24225 9137 24259
rect 9137 24225 9171 24259
rect 9171 24225 9180 24259
rect 9128 24216 9180 24225
rect 9496 24216 9548 24268
rect 8024 24148 8076 24200
rect 8852 24148 8904 24200
rect 9588 24148 9640 24200
rect 9956 24216 10008 24268
rect 10508 24259 10560 24268
rect 10508 24225 10517 24259
rect 10517 24225 10551 24259
rect 10551 24225 10560 24259
rect 10508 24216 10560 24225
rect 11060 24284 11112 24336
rect 11704 24284 11756 24336
rect 13176 24216 13228 24268
rect 13268 24259 13320 24268
rect 13268 24225 13277 24259
rect 13277 24225 13311 24259
rect 13311 24225 13320 24259
rect 14924 24284 14976 24336
rect 16764 24284 16816 24336
rect 13268 24216 13320 24225
rect 14648 24216 14700 24268
rect 15108 24216 15160 24268
rect 16488 24216 16540 24268
rect 16948 24259 17000 24268
rect 16948 24225 16957 24259
rect 16957 24225 16991 24259
rect 16991 24225 17000 24259
rect 16948 24216 17000 24225
rect 18144 24259 18196 24268
rect 18144 24225 18153 24259
rect 18153 24225 18187 24259
rect 18187 24225 18196 24259
rect 18144 24216 18196 24225
rect 19340 24284 19392 24336
rect 19984 24284 20036 24336
rect 19432 24216 19484 24268
rect 20904 24216 20956 24268
rect 21088 24259 21140 24268
rect 21088 24225 21097 24259
rect 21097 24225 21131 24259
rect 21131 24225 21140 24259
rect 21088 24216 21140 24225
rect 11704 24148 11756 24200
rect 12072 24191 12124 24200
rect 12072 24157 12081 24191
rect 12081 24157 12115 24191
rect 12115 24157 12124 24191
rect 12072 24148 12124 24157
rect 12164 24148 12216 24200
rect 2412 24123 2464 24132
rect 2412 24089 2421 24123
rect 2421 24089 2455 24123
rect 2455 24089 2464 24123
rect 2412 24080 2464 24089
rect 12532 24080 12584 24132
rect 17224 24148 17276 24200
rect 13820 24080 13872 24132
rect 24952 24352 25004 24404
rect 28080 24352 28132 24404
rect 25228 24284 25280 24336
rect 28724 24352 28776 24404
rect 34704 24352 34756 24404
rect 37832 24395 37884 24404
rect 37832 24361 37841 24395
rect 37841 24361 37875 24395
rect 37875 24361 37884 24395
rect 37832 24352 37884 24361
rect 21732 24259 21784 24268
rect 21732 24225 21741 24259
rect 21741 24225 21775 24259
rect 21775 24225 21784 24259
rect 21732 24216 21784 24225
rect 22652 24216 22704 24268
rect 23664 24259 23716 24268
rect 23664 24225 23673 24259
rect 23673 24225 23707 24259
rect 23707 24225 23716 24259
rect 23664 24216 23716 24225
rect 24032 24216 24084 24268
rect 24768 24216 24820 24268
rect 25044 24259 25096 24268
rect 25044 24225 25053 24259
rect 25053 24225 25087 24259
rect 25087 24225 25096 24259
rect 25044 24216 25096 24225
rect 25688 24259 25740 24268
rect 25688 24225 25697 24259
rect 25697 24225 25731 24259
rect 25731 24225 25740 24259
rect 25688 24216 25740 24225
rect 34796 24284 34848 24336
rect 35900 24284 35952 24336
rect 27436 24216 27488 24268
rect 28264 24259 28316 24268
rect 28264 24225 28273 24259
rect 28273 24225 28307 24259
rect 28307 24225 28316 24259
rect 28264 24216 28316 24225
rect 29000 24216 29052 24268
rect 31208 24216 31260 24268
rect 32128 24259 32180 24268
rect 24584 24148 24636 24200
rect 24676 24148 24728 24200
rect 26792 24148 26844 24200
rect 29368 24191 29420 24200
rect 29368 24157 29377 24191
rect 29377 24157 29411 24191
rect 29411 24157 29420 24191
rect 29368 24148 29420 24157
rect 9128 24012 9180 24064
rect 10508 24012 10560 24064
rect 14924 24012 14976 24064
rect 15660 24012 15712 24064
rect 19340 24012 19392 24064
rect 20260 24055 20312 24064
rect 20260 24021 20269 24055
rect 20269 24021 20303 24055
rect 20303 24021 20312 24055
rect 20260 24012 20312 24021
rect 24676 24012 24728 24064
rect 26700 24055 26752 24064
rect 26700 24021 26709 24055
rect 26709 24021 26743 24055
rect 26743 24021 26752 24055
rect 26700 24012 26752 24021
rect 27896 24012 27948 24064
rect 30472 24055 30524 24064
rect 30472 24021 30481 24055
rect 30481 24021 30515 24055
rect 30515 24021 30524 24055
rect 30472 24012 30524 24021
rect 32128 24225 32137 24259
rect 32137 24225 32171 24259
rect 32171 24225 32180 24259
rect 32128 24216 32180 24225
rect 33416 24216 33468 24268
rect 34520 24259 34572 24268
rect 34520 24225 34529 24259
rect 34529 24225 34563 24259
rect 34563 24225 34572 24259
rect 34520 24216 34572 24225
rect 34704 24259 34756 24268
rect 34704 24225 34713 24259
rect 34713 24225 34747 24259
rect 34747 24225 34756 24259
rect 34704 24216 34756 24225
rect 36268 24259 36320 24268
rect 33324 24148 33376 24200
rect 34244 24191 34296 24200
rect 34244 24157 34253 24191
rect 34253 24157 34287 24191
rect 34287 24157 34296 24191
rect 36268 24225 36277 24259
rect 36277 24225 36311 24259
rect 36311 24225 36320 24259
rect 36268 24216 36320 24225
rect 36544 24259 36596 24268
rect 36544 24225 36553 24259
rect 36553 24225 36587 24259
rect 36587 24225 36596 24259
rect 36544 24216 36596 24225
rect 36820 24259 36872 24268
rect 36820 24225 36829 24259
rect 36829 24225 36863 24259
rect 36863 24225 36872 24259
rect 36820 24216 36872 24225
rect 34244 24148 34296 24157
rect 31576 24080 31628 24132
rect 32036 24080 32088 24132
rect 36360 24080 36412 24132
rect 32588 24012 32640 24064
rect 33048 24012 33100 24064
rect 33692 24012 33744 24064
rect 4246 23910 4298 23962
rect 4310 23910 4362 23962
rect 4374 23910 4426 23962
rect 4438 23910 4490 23962
rect 34966 23910 35018 23962
rect 35030 23910 35082 23962
rect 35094 23910 35146 23962
rect 35158 23910 35210 23962
rect 7932 23808 7984 23860
rect 9220 23808 9272 23860
rect 23020 23851 23072 23860
rect 23020 23817 23029 23851
rect 23029 23817 23063 23851
rect 23063 23817 23072 23851
rect 23020 23808 23072 23817
rect 23204 23808 23256 23860
rect 24032 23808 24084 23860
rect 25044 23808 25096 23860
rect 29368 23808 29420 23860
rect 1676 23672 1728 23724
rect 2412 23715 2464 23724
rect 2412 23681 2421 23715
rect 2421 23681 2455 23715
rect 2455 23681 2464 23715
rect 2412 23672 2464 23681
rect 3148 23672 3200 23724
rect 2872 23647 2924 23656
rect 2872 23613 2881 23647
rect 2881 23613 2915 23647
rect 2915 23613 2924 23647
rect 2872 23604 2924 23613
rect 3332 23647 3384 23656
rect 3332 23613 3341 23647
rect 3341 23613 3375 23647
rect 3375 23613 3384 23647
rect 3332 23604 3384 23613
rect 6184 23672 6236 23724
rect 5448 23647 5500 23656
rect 4620 23536 4672 23588
rect 5448 23613 5457 23647
rect 5457 23613 5491 23647
rect 5491 23613 5500 23647
rect 5448 23604 5500 23613
rect 6552 23604 6604 23656
rect 7288 23604 7340 23656
rect 8116 23647 8168 23656
rect 8116 23613 8125 23647
rect 8125 23613 8159 23647
rect 8159 23613 8168 23647
rect 8116 23604 8168 23613
rect 8576 23647 8628 23656
rect 8576 23613 8585 23647
rect 8585 23613 8619 23647
rect 8619 23613 8628 23647
rect 8576 23604 8628 23613
rect 9864 23672 9916 23724
rect 10324 23672 10376 23724
rect 10692 23715 10744 23724
rect 10692 23681 10701 23715
rect 10701 23681 10735 23715
rect 10735 23681 10744 23715
rect 10692 23672 10744 23681
rect 11060 23672 11112 23724
rect 12624 23672 12676 23724
rect 14556 23740 14608 23792
rect 17132 23783 17184 23792
rect 17132 23749 17141 23783
rect 17141 23749 17175 23783
rect 17175 23749 17184 23783
rect 17132 23740 17184 23749
rect 11152 23647 11204 23656
rect 11152 23613 11161 23647
rect 11161 23613 11195 23647
rect 11195 23613 11204 23647
rect 11152 23604 11204 23613
rect 11704 23647 11756 23656
rect 11704 23613 11713 23647
rect 11713 23613 11747 23647
rect 11747 23613 11756 23647
rect 11704 23604 11756 23613
rect 12532 23647 12584 23656
rect 12532 23613 12541 23647
rect 12541 23613 12575 23647
rect 12575 23613 12584 23647
rect 12532 23604 12584 23613
rect 14648 23672 14700 23724
rect 15936 23672 15988 23724
rect 14924 23647 14976 23656
rect 6828 23536 6880 23588
rect 9956 23579 10008 23588
rect 9956 23545 9965 23579
rect 9965 23545 9999 23579
rect 9999 23545 10008 23579
rect 9956 23536 10008 23545
rect 4528 23468 4580 23520
rect 8668 23468 8720 23520
rect 10968 23468 11020 23520
rect 14924 23613 14933 23647
rect 14933 23613 14967 23647
rect 14967 23613 14976 23647
rect 14924 23604 14976 23613
rect 15476 23604 15528 23656
rect 16212 23604 16264 23656
rect 16580 23604 16632 23656
rect 17132 23647 17184 23656
rect 15384 23536 15436 23588
rect 17132 23613 17141 23647
rect 17141 23613 17175 23647
rect 17175 23613 17184 23647
rect 17132 23604 17184 23613
rect 18512 23647 18564 23656
rect 18512 23613 18521 23647
rect 18521 23613 18555 23647
rect 18555 23613 18564 23647
rect 18512 23604 18564 23613
rect 21364 23740 21416 23792
rect 22376 23740 22428 23792
rect 19340 23715 19392 23724
rect 19340 23681 19349 23715
rect 19349 23681 19383 23715
rect 19383 23681 19392 23715
rect 19340 23672 19392 23681
rect 21732 23672 21784 23724
rect 22008 23672 22060 23724
rect 19248 23647 19300 23656
rect 19248 23613 19257 23647
rect 19257 23613 19291 23647
rect 19291 23613 19300 23647
rect 19248 23604 19300 23613
rect 20628 23604 20680 23656
rect 17408 23536 17460 23588
rect 21180 23604 21232 23656
rect 22100 23647 22152 23656
rect 22100 23613 22109 23647
rect 22109 23613 22143 23647
rect 22143 23613 22152 23647
rect 22100 23604 22152 23613
rect 22744 23604 22796 23656
rect 23940 23672 23992 23724
rect 24676 23672 24728 23724
rect 26700 23672 26752 23724
rect 32128 23808 32180 23860
rect 24492 23647 24544 23656
rect 24492 23613 24501 23647
rect 24501 23613 24535 23647
rect 24535 23613 24544 23647
rect 24492 23604 24544 23613
rect 24860 23647 24912 23656
rect 15108 23468 15160 23520
rect 22652 23536 22704 23588
rect 24860 23613 24869 23647
rect 24869 23613 24903 23647
rect 24903 23613 24912 23647
rect 24860 23604 24912 23613
rect 26792 23647 26844 23656
rect 26792 23613 26801 23647
rect 26801 23613 26835 23647
rect 26835 23613 26844 23647
rect 26792 23604 26844 23613
rect 26976 23647 27028 23656
rect 26976 23613 26985 23647
rect 26985 23613 27019 23647
rect 27019 23613 27028 23647
rect 26976 23604 27028 23613
rect 25688 23536 25740 23588
rect 26608 23536 26660 23588
rect 27896 23604 27948 23656
rect 28632 23604 28684 23656
rect 29552 23536 29604 23588
rect 29920 23536 29972 23588
rect 26148 23468 26200 23520
rect 27712 23511 27764 23520
rect 27712 23477 27721 23511
rect 27721 23477 27755 23511
rect 27755 23477 27764 23511
rect 27712 23468 27764 23477
rect 29644 23468 29696 23520
rect 31024 23672 31076 23724
rect 31484 23715 31536 23724
rect 30564 23647 30616 23656
rect 30564 23613 30573 23647
rect 30573 23613 30607 23647
rect 30607 23613 30616 23647
rect 30564 23604 30616 23613
rect 31208 23647 31260 23656
rect 31208 23613 31217 23647
rect 31217 23613 31251 23647
rect 31251 23613 31260 23647
rect 31208 23604 31260 23613
rect 31484 23681 31493 23715
rect 31493 23681 31527 23715
rect 31527 23681 31536 23715
rect 31484 23672 31536 23681
rect 35716 23715 35768 23724
rect 34796 23604 34848 23656
rect 35716 23681 35725 23715
rect 35725 23681 35759 23715
rect 35759 23681 35768 23715
rect 35716 23672 35768 23681
rect 36084 23672 36136 23724
rect 35532 23604 35584 23656
rect 36820 23672 36872 23724
rect 36728 23647 36780 23656
rect 36728 23613 36737 23647
rect 36737 23613 36771 23647
rect 36771 23613 36780 23647
rect 36728 23604 36780 23613
rect 30380 23536 30432 23588
rect 34336 23579 34388 23588
rect 34336 23545 34345 23579
rect 34345 23545 34379 23579
rect 34379 23545 34388 23579
rect 34336 23536 34388 23545
rect 34244 23468 34296 23520
rect 37832 23511 37884 23520
rect 37832 23477 37841 23511
rect 37841 23477 37875 23511
rect 37875 23477 37884 23511
rect 37832 23468 37884 23477
rect 19606 23366 19658 23418
rect 19670 23366 19722 23418
rect 19734 23366 19786 23418
rect 19798 23366 19850 23418
rect 7564 23264 7616 23316
rect 8484 23264 8536 23316
rect 8668 23264 8720 23316
rect 14372 23264 14424 23316
rect 15016 23264 15068 23316
rect 17132 23307 17184 23316
rect 3608 23128 3660 23180
rect 4528 23171 4580 23180
rect 4528 23137 4537 23171
rect 4537 23137 4571 23171
rect 4571 23137 4580 23171
rect 4528 23128 4580 23137
rect 7288 23196 7340 23248
rect 9404 23196 9456 23248
rect 6828 23128 6880 23180
rect 7380 23171 7432 23180
rect 7380 23137 7389 23171
rect 7389 23137 7423 23171
rect 7423 23137 7432 23171
rect 7380 23128 7432 23137
rect 8116 23171 8168 23180
rect 4068 23060 4120 23112
rect 1400 22992 1452 23044
rect 4712 23060 4764 23112
rect 8116 23137 8125 23171
rect 8125 23137 8159 23171
rect 8159 23137 8168 23171
rect 8116 23128 8168 23137
rect 8852 23171 8904 23180
rect 8852 23137 8861 23171
rect 8861 23137 8895 23171
rect 8895 23137 8904 23171
rect 8852 23128 8904 23137
rect 9312 23128 9364 23180
rect 12532 23196 12584 23248
rect 13268 23196 13320 23248
rect 12164 23171 12216 23180
rect 10324 23060 10376 23112
rect 11152 23103 11204 23112
rect 11152 23069 11161 23103
rect 11161 23069 11195 23103
rect 11195 23069 11204 23103
rect 11152 23060 11204 23069
rect 12164 23137 12173 23171
rect 12173 23137 12207 23171
rect 12207 23137 12216 23171
rect 12164 23128 12216 23137
rect 12624 23171 12676 23180
rect 12624 23137 12633 23171
rect 12633 23137 12667 23171
rect 12667 23137 12676 23171
rect 12624 23128 12676 23137
rect 13912 23128 13964 23180
rect 15292 23128 15344 23180
rect 16672 23196 16724 23248
rect 17132 23273 17141 23307
rect 17141 23273 17175 23307
rect 17175 23273 17184 23307
rect 17132 23264 17184 23273
rect 18880 23196 18932 23248
rect 19248 23196 19300 23248
rect 19984 23264 20036 23316
rect 21548 23264 21600 23316
rect 18512 23171 18564 23180
rect 14464 23103 14516 23112
rect 6552 23035 6604 23044
rect 6552 23001 6561 23035
rect 6561 23001 6595 23035
rect 6595 23001 6604 23035
rect 6552 22992 6604 23001
rect 7380 22992 7432 23044
rect 9956 22992 10008 23044
rect 14464 23069 14473 23103
rect 14473 23069 14507 23103
rect 14507 23069 14516 23103
rect 14464 23060 14516 23069
rect 14924 23060 14976 23112
rect 14004 22992 14056 23044
rect 15108 22992 15160 23044
rect 18512 23137 18521 23171
rect 18521 23137 18555 23171
rect 18555 23137 18564 23171
rect 18512 23128 18564 23137
rect 19064 23171 19116 23180
rect 19064 23137 19073 23171
rect 19073 23137 19107 23171
rect 19107 23137 19116 23171
rect 19064 23128 19116 23137
rect 20812 23196 20864 23248
rect 22376 23196 22428 23248
rect 20076 23171 20128 23180
rect 20076 23137 20085 23171
rect 20085 23137 20119 23171
rect 20119 23137 20128 23171
rect 20076 23128 20128 23137
rect 21180 23171 21232 23180
rect 21180 23137 21189 23171
rect 21189 23137 21223 23171
rect 21223 23137 21232 23171
rect 21180 23128 21232 23137
rect 21916 23128 21968 23180
rect 24032 23196 24084 23248
rect 27712 23264 27764 23316
rect 29000 23264 29052 23316
rect 28264 23196 28316 23248
rect 30472 23264 30524 23316
rect 31392 23264 31444 23316
rect 21640 23103 21692 23112
rect 1676 22924 1728 22976
rect 5632 22967 5684 22976
rect 5632 22933 5641 22967
rect 5641 22933 5675 22967
rect 5675 22933 5684 22967
rect 5632 22924 5684 22933
rect 12716 22967 12768 22976
rect 12716 22933 12725 22967
rect 12725 22933 12759 22967
rect 12759 22933 12768 22967
rect 12716 22924 12768 22933
rect 12900 22924 12952 22976
rect 21640 23069 21649 23103
rect 21649 23069 21683 23103
rect 21683 23069 21692 23103
rect 21640 23060 21692 23069
rect 21824 23060 21876 23112
rect 23848 23128 23900 23180
rect 24216 23171 24268 23180
rect 24216 23137 24225 23171
rect 24225 23137 24259 23171
rect 24259 23137 24268 23171
rect 24216 23128 24268 23137
rect 26608 23128 26660 23180
rect 27620 23128 27672 23180
rect 24400 23060 24452 23112
rect 24860 23060 24912 23112
rect 26516 23103 26568 23112
rect 26516 23069 26525 23103
rect 26525 23069 26559 23103
rect 26559 23069 26568 23103
rect 26516 23060 26568 23069
rect 26700 23060 26752 23112
rect 29828 23060 29880 23112
rect 30012 23103 30064 23112
rect 30012 23069 30021 23103
rect 30021 23069 30055 23103
rect 30055 23069 30064 23103
rect 30012 23060 30064 23069
rect 30288 23171 30340 23180
rect 30288 23137 30297 23171
rect 30297 23137 30331 23171
rect 30331 23137 30340 23171
rect 31208 23196 31260 23248
rect 32404 23239 32456 23248
rect 32404 23205 32413 23239
rect 32413 23205 32447 23239
rect 32447 23205 32456 23239
rect 32404 23196 32456 23205
rect 32956 23239 33008 23248
rect 32956 23205 32965 23239
rect 32965 23205 32999 23239
rect 32999 23205 33008 23239
rect 32956 23196 33008 23205
rect 30288 23128 30340 23137
rect 31300 23171 31352 23180
rect 31300 23137 31309 23171
rect 31309 23137 31343 23171
rect 31343 23137 31352 23171
rect 31300 23128 31352 23137
rect 32680 23128 32732 23180
rect 34520 23264 34572 23316
rect 33692 23171 33744 23180
rect 33692 23137 33701 23171
rect 33701 23137 33735 23171
rect 33735 23137 33744 23171
rect 33692 23128 33744 23137
rect 35992 23171 36044 23180
rect 35992 23137 36001 23171
rect 36001 23137 36035 23171
rect 36035 23137 36044 23171
rect 35992 23128 36044 23137
rect 36452 23171 36504 23180
rect 36452 23137 36461 23171
rect 36461 23137 36495 23171
rect 36495 23137 36504 23171
rect 36452 23128 36504 23137
rect 37832 23128 37884 23180
rect 30380 23060 30432 23112
rect 31116 23060 31168 23112
rect 31392 23060 31444 23112
rect 35900 23060 35952 23112
rect 16580 22992 16632 23044
rect 25320 23035 25372 23044
rect 25320 23001 25329 23035
rect 25329 23001 25363 23035
rect 25363 23001 25372 23035
rect 25320 22992 25372 23001
rect 18972 22924 19024 22976
rect 22376 22924 22428 22976
rect 23388 22967 23440 22976
rect 23388 22933 23397 22967
rect 23397 22933 23431 22967
rect 23431 22933 23440 22967
rect 23388 22924 23440 22933
rect 24584 22924 24636 22976
rect 34704 22924 34756 22976
rect 35808 22924 35860 22976
rect 4246 22822 4298 22874
rect 4310 22822 4362 22874
rect 4374 22822 4426 22874
rect 4438 22822 4490 22874
rect 34966 22822 35018 22874
rect 35030 22822 35082 22874
rect 35094 22822 35146 22874
rect 35158 22822 35210 22874
rect 3148 22720 3200 22772
rect 3608 22763 3660 22772
rect 3608 22729 3617 22763
rect 3617 22729 3651 22763
rect 3651 22729 3660 22763
rect 3608 22720 3660 22729
rect 4620 22720 4672 22772
rect 7288 22652 7340 22704
rect 9680 22652 9732 22704
rect 1400 22627 1452 22636
rect 1400 22593 1409 22627
rect 1409 22593 1443 22627
rect 1443 22593 1452 22627
rect 1400 22584 1452 22593
rect 1676 22627 1728 22636
rect 1676 22593 1685 22627
rect 1685 22593 1719 22627
rect 1719 22593 1728 22627
rect 1676 22584 1728 22593
rect 3700 22559 3752 22568
rect 3700 22525 3709 22559
rect 3709 22525 3743 22559
rect 3743 22525 3752 22559
rect 3700 22516 3752 22525
rect 3332 22448 3384 22500
rect 4712 22516 4764 22568
rect 5356 22516 5408 22568
rect 5632 22584 5684 22636
rect 7380 22627 7432 22636
rect 7380 22593 7389 22627
rect 7389 22593 7423 22627
rect 7423 22593 7432 22627
rect 7380 22584 7432 22593
rect 7748 22584 7800 22636
rect 8760 22584 8812 22636
rect 13176 22627 13228 22636
rect 5540 22516 5592 22568
rect 2964 22423 3016 22432
rect 2964 22389 2973 22423
rect 2973 22389 3007 22423
rect 3007 22389 3016 22423
rect 2964 22380 3016 22389
rect 6828 22516 6880 22568
rect 8576 22516 8628 22568
rect 9404 22559 9456 22568
rect 9404 22525 9413 22559
rect 9413 22525 9447 22559
rect 9447 22525 9456 22559
rect 9404 22516 9456 22525
rect 9588 22559 9640 22568
rect 9588 22525 9597 22559
rect 9597 22525 9631 22559
rect 9631 22525 9640 22559
rect 9588 22516 9640 22525
rect 10048 22559 10100 22568
rect 10048 22525 10057 22559
rect 10057 22525 10091 22559
rect 10091 22525 10100 22559
rect 10048 22516 10100 22525
rect 10324 22559 10376 22568
rect 10324 22525 10333 22559
rect 10333 22525 10367 22559
rect 10367 22525 10376 22559
rect 10324 22516 10376 22525
rect 11336 22559 11388 22568
rect 11336 22525 11345 22559
rect 11345 22525 11379 22559
rect 11379 22525 11388 22559
rect 11336 22516 11388 22525
rect 12164 22516 12216 22568
rect 12532 22516 12584 22568
rect 7748 22491 7800 22500
rect 7748 22457 7757 22491
rect 7757 22457 7791 22491
rect 7791 22457 7800 22491
rect 7748 22448 7800 22457
rect 8116 22448 8168 22500
rect 9864 22448 9916 22500
rect 10416 22448 10468 22500
rect 13176 22593 13185 22627
rect 13185 22593 13219 22627
rect 13219 22593 13228 22627
rect 13176 22584 13228 22593
rect 14372 22559 14424 22568
rect 14372 22525 14381 22559
rect 14381 22525 14415 22559
rect 14415 22525 14424 22559
rect 14372 22516 14424 22525
rect 16672 22720 16724 22772
rect 17224 22720 17276 22772
rect 16948 22652 17000 22704
rect 19340 22720 19392 22772
rect 22744 22763 22796 22772
rect 22744 22729 22753 22763
rect 22753 22729 22787 22763
rect 22787 22729 22796 22763
rect 22744 22720 22796 22729
rect 26884 22720 26936 22772
rect 37464 22763 37516 22772
rect 15568 22516 15620 22568
rect 16672 22559 16724 22568
rect 16672 22525 16681 22559
rect 16681 22525 16715 22559
rect 16715 22525 16724 22559
rect 16672 22516 16724 22525
rect 17500 22516 17552 22568
rect 21916 22652 21968 22704
rect 19432 22559 19484 22568
rect 15108 22448 15160 22500
rect 19432 22525 19441 22559
rect 19441 22525 19475 22559
rect 19475 22525 19484 22559
rect 19432 22516 19484 22525
rect 19984 22516 20036 22568
rect 21548 22584 21600 22636
rect 8024 22380 8076 22432
rect 12532 22380 12584 22432
rect 13084 22380 13136 22432
rect 16120 22380 16172 22432
rect 16212 22380 16264 22432
rect 20444 22448 20496 22500
rect 20720 22448 20772 22500
rect 21916 22516 21968 22568
rect 22376 22516 22428 22568
rect 23388 22652 23440 22704
rect 24400 22627 24452 22636
rect 22652 22516 22704 22568
rect 23388 22516 23440 22568
rect 24124 22559 24176 22568
rect 24124 22525 24133 22559
rect 24133 22525 24167 22559
rect 24167 22525 24176 22559
rect 24124 22516 24176 22525
rect 24400 22593 24409 22627
rect 24409 22593 24443 22627
rect 24443 22593 24452 22627
rect 24400 22584 24452 22593
rect 26700 22584 26752 22636
rect 26976 22584 27028 22636
rect 24216 22448 24268 22500
rect 24952 22448 25004 22500
rect 26884 22516 26936 22568
rect 27344 22448 27396 22500
rect 27896 22627 27948 22636
rect 27896 22593 27905 22627
rect 27905 22593 27939 22627
rect 27939 22593 27948 22627
rect 27896 22584 27948 22593
rect 37464 22729 37473 22763
rect 37473 22729 37507 22763
rect 37507 22729 37516 22763
rect 37464 22720 37516 22729
rect 30012 22695 30064 22704
rect 30012 22661 30021 22695
rect 30021 22661 30055 22695
rect 30055 22661 30064 22695
rect 30012 22652 30064 22661
rect 28632 22584 28684 22636
rect 29552 22559 29604 22568
rect 29552 22525 29561 22559
rect 29561 22525 29595 22559
rect 29595 22525 29604 22559
rect 29552 22516 29604 22525
rect 30288 22516 30340 22568
rect 30840 22559 30892 22568
rect 30840 22525 30849 22559
rect 30849 22525 30883 22559
rect 30883 22525 30892 22559
rect 30840 22516 30892 22525
rect 20352 22380 20404 22432
rect 22100 22380 22152 22432
rect 31208 22584 31260 22636
rect 31760 22584 31812 22636
rect 32680 22584 32732 22636
rect 31852 22559 31904 22568
rect 31852 22525 31861 22559
rect 31861 22525 31895 22559
rect 31895 22525 31904 22559
rect 31852 22516 31904 22525
rect 33784 22559 33836 22568
rect 33784 22525 33793 22559
rect 33793 22525 33827 22559
rect 33827 22525 33836 22559
rect 33784 22516 33836 22525
rect 34612 22584 34664 22636
rect 33600 22448 33652 22500
rect 34060 22516 34112 22568
rect 35348 22516 35400 22568
rect 36084 22559 36136 22568
rect 36084 22525 36093 22559
rect 36093 22525 36127 22559
rect 36127 22525 36136 22559
rect 36084 22516 36136 22525
rect 35624 22448 35676 22500
rect 33140 22423 33192 22432
rect 33140 22389 33149 22423
rect 33149 22389 33183 22423
rect 33183 22389 33192 22423
rect 33140 22380 33192 22389
rect 19606 22278 19658 22330
rect 19670 22278 19722 22330
rect 19734 22278 19786 22330
rect 19798 22278 19850 22330
rect 6828 22176 6880 22228
rect 7472 22176 7524 22228
rect 8760 22176 8812 22228
rect 12256 22176 12308 22228
rect 17500 22219 17552 22228
rect 1768 22083 1820 22092
rect 1768 22049 1777 22083
rect 1777 22049 1811 22083
rect 1811 22049 1820 22083
rect 1768 22040 1820 22049
rect 3148 22083 3200 22092
rect 3148 22049 3157 22083
rect 3157 22049 3191 22083
rect 3191 22049 3200 22083
rect 3148 22040 3200 22049
rect 4620 22040 4672 22092
rect 4896 22040 4948 22092
rect 5632 22040 5684 22092
rect 7748 22108 7800 22160
rect 8852 22108 8904 22160
rect 3424 22015 3476 22024
rect 3424 21981 3433 22015
rect 3433 21981 3467 22015
rect 3467 21981 3476 22015
rect 3424 21972 3476 21981
rect 3700 21972 3752 22024
rect 4068 21972 4120 22024
rect 7288 22015 7340 22024
rect 7288 21981 7297 22015
rect 7297 21981 7331 22015
rect 7331 21981 7340 22015
rect 7288 21972 7340 21981
rect 8576 22083 8628 22092
rect 8576 22049 8585 22083
rect 8585 22049 8619 22083
rect 8619 22049 8628 22083
rect 9496 22083 9548 22092
rect 8576 22040 8628 22049
rect 9496 22049 9505 22083
rect 9505 22049 9539 22083
rect 9539 22049 9548 22083
rect 9496 22040 9548 22049
rect 10324 22108 10376 22160
rect 10048 22083 10100 22092
rect 10048 22049 10057 22083
rect 10057 22049 10091 22083
rect 10091 22049 10100 22083
rect 10048 22040 10100 22049
rect 10416 22083 10468 22092
rect 10416 22049 10425 22083
rect 10425 22049 10459 22083
rect 10459 22049 10468 22083
rect 10416 22040 10468 22049
rect 12624 22040 12676 22092
rect 15108 22108 15160 22160
rect 17500 22185 17509 22219
rect 17509 22185 17543 22219
rect 17543 22185 17552 22219
rect 17500 22176 17552 22185
rect 23112 22176 23164 22228
rect 23388 22176 23440 22228
rect 26792 22219 26844 22228
rect 26792 22185 26801 22219
rect 26801 22185 26835 22219
rect 26835 22185 26844 22219
rect 26792 22176 26844 22185
rect 28172 22176 28224 22228
rect 30380 22176 30432 22228
rect 33508 22176 33560 22228
rect 19984 22108 20036 22160
rect 20076 22108 20128 22160
rect 24492 22108 24544 22160
rect 10600 22015 10652 22024
rect 2320 21904 2372 21956
rect 4160 21947 4212 21956
rect 4160 21913 4169 21947
rect 4169 21913 4203 21947
rect 4203 21913 4212 21947
rect 4160 21904 4212 21913
rect 10600 21981 10609 22015
rect 10609 21981 10643 22015
rect 10643 21981 10652 22015
rect 10600 21972 10652 21981
rect 9772 21904 9824 21956
rect 12716 21972 12768 22024
rect 17040 22040 17092 22092
rect 18880 22040 18932 22092
rect 19064 22083 19116 22092
rect 19064 22049 19073 22083
rect 19073 22049 19107 22083
rect 19107 22049 19116 22083
rect 19064 22040 19116 22049
rect 19708 22083 19760 22092
rect 19708 22049 19717 22083
rect 19717 22049 19751 22083
rect 19751 22049 19760 22083
rect 19708 22040 19760 22049
rect 21732 22040 21784 22092
rect 21824 22040 21876 22092
rect 22192 22040 22244 22092
rect 22744 22083 22796 22092
rect 22744 22049 22753 22083
rect 22753 22049 22787 22083
rect 22787 22049 22796 22083
rect 22744 22040 22796 22049
rect 23388 22083 23440 22092
rect 23388 22049 23397 22083
rect 23397 22049 23431 22083
rect 23431 22049 23440 22083
rect 23388 22040 23440 22049
rect 25412 22083 25464 22092
rect 15016 21904 15068 21956
rect 17224 21972 17276 22024
rect 25412 22049 25421 22083
rect 25421 22049 25455 22083
rect 25455 22049 25464 22083
rect 25412 22040 25464 22049
rect 26884 22083 26936 22092
rect 26884 22049 26893 22083
rect 26893 22049 26927 22083
rect 26927 22049 26936 22083
rect 26884 22040 26936 22049
rect 27344 22083 27396 22092
rect 27344 22049 27353 22083
rect 27353 22049 27387 22083
rect 27387 22049 27396 22083
rect 27344 22040 27396 22049
rect 27528 22083 27580 22092
rect 27528 22049 27537 22083
rect 27537 22049 27571 22083
rect 27571 22049 27580 22083
rect 27528 22040 27580 22049
rect 29552 22108 29604 22160
rect 17776 21904 17828 21956
rect 18788 21904 18840 21956
rect 24400 21972 24452 22024
rect 24952 22015 25004 22024
rect 24952 21981 24961 22015
rect 24961 21981 24995 22015
rect 24995 21981 25004 22015
rect 24952 21972 25004 21981
rect 26976 21972 27028 22024
rect 27988 21972 28040 22024
rect 29000 22015 29052 22024
rect 29000 21981 29009 22015
rect 29009 21981 29043 22015
rect 29043 21981 29052 22015
rect 29000 21972 29052 21981
rect 29368 22040 29420 22092
rect 30656 22083 30708 22092
rect 30656 22049 30665 22083
rect 30665 22049 30699 22083
rect 30699 22049 30708 22083
rect 30656 22040 30708 22049
rect 30840 22083 30892 22092
rect 30840 22049 30849 22083
rect 30849 22049 30883 22083
rect 30883 22049 30892 22083
rect 30840 22040 30892 22049
rect 31208 22040 31260 22092
rect 32128 22083 32180 22092
rect 32128 22049 32137 22083
rect 32137 22049 32171 22083
rect 32171 22049 32180 22083
rect 32128 22040 32180 22049
rect 32680 22083 32732 22092
rect 32680 22049 32689 22083
rect 32689 22049 32723 22083
rect 32723 22049 32732 22083
rect 32680 22040 32732 22049
rect 33324 22083 33376 22092
rect 31852 21972 31904 22024
rect 33324 22049 33333 22083
rect 33333 22049 33367 22083
rect 33367 22049 33376 22083
rect 33324 22040 33376 22049
rect 34244 22108 34296 22160
rect 37280 22108 37332 22160
rect 35808 22083 35860 22092
rect 34796 22015 34848 22024
rect 34796 21981 34805 22015
rect 34805 21981 34839 22015
rect 34839 21981 34848 22015
rect 34796 21972 34848 21981
rect 35808 22049 35817 22083
rect 35817 22049 35851 22083
rect 35851 22049 35860 22083
rect 35808 22040 35860 22049
rect 37648 22040 37700 22092
rect 36452 21972 36504 22024
rect 33140 21904 33192 21956
rect 33232 21904 33284 21956
rect 34428 21904 34480 21956
rect 35532 21904 35584 21956
rect 3148 21836 3200 21888
rect 4712 21836 4764 21888
rect 7656 21836 7708 21888
rect 13912 21836 13964 21888
rect 15384 21836 15436 21888
rect 32680 21836 32732 21888
rect 33692 21836 33744 21888
rect 34244 21836 34296 21888
rect 36728 21836 36780 21888
rect 37004 21836 37056 21888
rect 4246 21734 4298 21786
rect 4310 21734 4362 21786
rect 4374 21734 4426 21786
rect 4438 21734 4490 21786
rect 34966 21734 35018 21786
rect 35030 21734 35082 21786
rect 35094 21734 35146 21786
rect 35158 21734 35210 21786
rect 7748 21632 7800 21684
rect 8576 21632 8628 21684
rect 17040 21632 17092 21684
rect 17592 21675 17644 21684
rect 17592 21641 17601 21675
rect 17601 21641 17635 21675
rect 17635 21641 17644 21675
rect 17592 21632 17644 21641
rect 20168 21632 20220 21684
rect 21640 21675 21692 21684
rect 21640 21641 21649 21675
rect 21649 21641 21683 21675
rect 21683 21641 21692 21675
rect 21640 21632 21692 21641
rect 21732 21632 21784 21684
rect 28632 21675 28684 21684
rect 28632 21641 28641 21675
rect 28641 21641 28675 21675
rect 28675 21641 28684 21675
rect 28632 21632 28684 21641
rect 30564 21632 30616 21684
rect 32496 21632 32548 21684
rect 32588 21632 32640 21684
rect 34428 21632 34480 21684
rect 37004 21632 37056 21684
rect 1768 21564 1820 21616
rect 1860 21496 1912 21548
rect 1492 21471 1544 21480
rect 1492 21437 1501 21471
rect 1501 21437 1535 21471
rect 1535 21437 1544 21471
rect 1492 21428 1544 21437
rect 2964 21496 3016 21548
rect 9404 21564 9456 21616
rect 12532 21564 12584 21616
rect 15568 21564 15620 21616
rect 16028 21564 16080 21616
rect 16488 21564 16540 21616
rect 3148 21471 3200 21480
rect 3148 21437 3157 21471
rect 3157 21437 3191 21471
rect 3191 21437 3200 21471
rect 3148 21428 3200 21437
rect 3424 21471 3476 21480
rect 3424 21437 3433 21471
rect 3433 21437 3467 21471
rect 3467 21437 3476 21471
rect 3424 21428 3476 21437
rect 4804 21428 4856 21480
rect 6184 21496 6236 21548
rect 4068 21360 4120 21412
rect 4712 21360 4764 21412
rect 5540 21428 5592 21480
rect 9680 21496 9732 21548
rect 16396 21539 16448 21548
rect 9864 21471 9916 21480
rect 1584 21335 1636 21344
rect 1584 21301 1593 21335
rect 1593 21301 1627 21335
rect 1627 21301 1636 21335
rect 1584 21292 1636 21301
rect 4620 21292 4672 21344
rect 5264 21292 5316 21344
rect 8576 21360 8628 21412
rect 9864 21437 9873 21471
rect 9873 21437 9907 21471
rect 9907 21437 9916 21471
rect 9864 21428 9916 21437
rect 10600 21471 10652 21480
rect 10600 21437 10609 21471
rect 10609 21437 10643 21471
rect 10643 21437 10652 21471
rect 10600 21428 10652 21437
rect 11336 21471 11388 21480
rect 11336 21437 11345 21471
rect 11345 21437 11379 21471
rect 11379 21437 11388 21471
rect 11336 21428 11388 21437
rect 16396 21505 16405 21539
rect 16405 21505 16439 21539
rect 16439 21505 16448 21539
rect 16396 21496 16448 21505
rect 19156 21564 19208 21616
rect 22284 21564 22336 21616
rect 13820 21428 13872 21480
rect 14004 21471 14056 21480
rect 14004 21437 14013 21471
rect 14013 21437 14047 21471
rect 14047 21437 14056 21471
rect 14004 21428 14056 21437
rect 14096 21360 14148 21412
rect 8116 21292 8168 21344
rect 12532 21335 12584 21344
rect 12532 21301 12541 21335
rect 12541 21301 12575 21335
rect 12575 21301 12584 21335
rect 12532 21292 12584 21301
rect 13728 21292 13780 21344
rect 15384 21428 15436 21480
rect 15568 21428 15620 21480
rect 16120 21471 16172 21480
rect 14372 21292 14424 21344
rect 16120 21437 16129 21471
rect 16129 21437 16163 21471
rect 16163 21437 16172 21471
rect 16120 21428 16172 21437
rect 17040 21428 17092 21480
rect 17960 21428 18012 21480
rect 18512 21428 18564 21480
rect 19340 21496 19392 21548
rect 18972 21471 19024 21480
rect 18972 21437 18981 21471
rect 18981 21437 19015 21471
rect 19015 21437 19024 21471
rect 18972 21428 19024 21437
rect 19892 21496 19944 21548
rect 24124 21496 24176 21548
rect 30380 21564 30432 21616
rect 31300 21564 31352 21616
rect 32404 21564 32456 21616
rect 26976 21496 27028 21548
rect 19800 21471 19852 21480
rect 19800 21437 19809 21471
rect 19809 21437 19843 21471
rect 19843 21437 19852 21471
rect 19800 21428 19852 21437
rect 15844 21360 15896 21412
rect 19432 21360 19484 21412
rect 20260 21428 20312 21480
rect 21180 21428 21232 21480
rect 21824 21471 21876 21480
rect 21824 21437 21833 21471
rect 21833 21437 21867 21471
rect 21867 21437 21876 21471
rect 21824 21428 21876 21437
rect 22284 21428 22336 21480
rect 22744 21428 22796 21480
rect 23572 21428 23624 21480
rect 16212 21292 16264 21344
rect 16488 21292 16540 21344
rect 20536 21292 20588 21344
rect 23664 21292 23716 21344
rect 24032 21428 24084 21480
rect 26516 21428 26568 21480
rect 27068 21428 27120 21480
rect 29368 21428 29420 21480
rect 29644 21428 29696 21480
rect 27252 21360 27304 21412
rect 27528 21360 27580 21412
rect 29920 21428 29972 21480
rect 31208 21496 31260 21548
rect 33232 21564 33284 21616
rect 32772 21539 32824 21548
rect 30932 21428 30984 21480
rect 32772 21505 32781 21539
rect 32781 21505 32815 21539
rect 32815 21505 32824 21539
rect 32772 21496 32824 21505
rect 33048 21496 33100 21548
rect 34336 21496 34388 21548
rect 37280 21496 37332 21548
rect 30472 21360 30524 21412
rect 31576 21403 31628 21412
rect 31576 21369 31585 21403
rect 31585 21369 31619 21403
rect 31619 21369 31628 21403
rect 31576 21360 31628 21369
rect 31760 21360 31812 21412
rect 32036 21360 32088 21412
rect 32220 21360 32272 21412
rect 32680 21360 32732 21412
rect 33968 21428 34020 21480
rect 35256 21428 35308 21480
rect 24400 21292 24452 21344
rect 29184 21292 29236 21344
rect 31484 21292 31536 21344
rect 36084 21428 36136 21480
rect 37648 21471 37700 21480
rect 37648 21437 37657 21471
rect 37657 21437 37691 21471
rect 37691 21437 37700 21471
rect 37648 21428 37700 21437
rect 37832 21471 37884 21480
rect 37832 21437 37841 21471
rect 37841 21437 37875 21471
rect 37875 21437 37884 21471
rect 37832 21428 37884 21437
rect 35900 21292 35952 21344
rect 37372 21292 37424 21344
rect 19606 21190 19658 21242
rect 19670 21190 19722 21242
rect 19734 21190 19786 21242
rect 19798 21190 19850 21242
rect 4068 21088 4120 21140
rect 8576 21088 8628 21140
rect 11336 21131 11388 21140
rect 11336 21097 11345 21131
rect 11345 21097 11379 21131
rect 11379 21097 11388 21131
rect 11336 21088 11388 21097
rect 14648 21131 14700 21140
rect 14648 21097 14657 21131
rect 14657 21097 14691 21131
rect 14691 21097 14700 21131
rect 14648 21088 14700 21097
rect 15384 21088 15436 21140
rect 21456 21088 21508 21140
rect 27252 21088 27304 21140
rect 29276 21088 29328 21140
rect 29552 21088 29604 21140
rect 32312 21088 32364 21140
rect 33048 21088 33100 21140
rect 1860 20995 1912 21004
rect 1860 20961 1869 20995
rect 1869 20961 1903 20995
rect 1903 20961 1912 20995
rect 1860 20952 1912 20961
rect 2320 20995 2372 21004
rect 2320 20961 2329 20995
rect 2329 20961 2363 20995
rect 2363 20961 2372 20995
rect 2320 20952 2372 20961
rect 2964 20995 3016 21004
rect 2964 20961 2973 20995
rect 2973 20961 3007 20995
rect 3007 20961 3016 20995
rect 2964 20952 3016 20961
rect 3424 20995 3476 21004
rect 3424 20961 3433 20995
rect 3433 20961 3467 20995
rect 3467 20961 3476 20995
rect 3424 20952 3476 20961
rect 5264 20952 5316 21004
rect 5540 20952 5592 21004
rect 6184 20995 6236 21004
rect 6184 20961 6193 20995
rect 6193 20961 6227 20995
rect 6227 20961 6236 20995
rect 6184 20952 6236 20961
rect 6460 20952 6512 21004
rect 8208 21020 8260 21072
rect 16764 21063 16816 21072
rect 16764 21029 16773 21063
rect 16773 21029 16807 21063
rect 16807 21029 16816 21063
rect 16764 21020 16816 21029
rect 17040 21020 17092 21072
rect 19984 21063 20036 21072
rect 7380 20995 7432 21004
rect 7380 20961 7389 20995
rect 7389 20961 7423 20995
rect 7423 20961 7432 20995
rect 7380 20952 7432 20961
rect 5908 20884 5960 20936
rect 6276 20927 6328 20936
rect 6276 20893 6285 20927
rect 6285 20893 6319 20927
rect 6319 20893 6328 20927
rect 6276 20884 6328 20893
rect 7012 20884 7064 20936
rect 8944 20995 8996 21004
rect 8944 20961 8953 20995
rect 8953 20961 8987 20995
rect 8987 20961 8996 20995
rect 8944 20952 8996 20961
rect 9772 20995 9824 21004
rect 9772 20961 9781 20995
rect 9781 20961 9815 20995
rect 9815 20961 9824 20995
rect 9772 20952 9824 20961
rect 12532 20952 12584 21004
rect 9496 20884 9548 20936
rect 1492 20816 1544 20868
rect 9036 20859 9088 20868
rect 9036 20825 9045 20859
rect 9045 20825 9079 20859
rect 9079 20825 9088 20859
rect 14464 20952 14516 21004
rect 15200 20952 15252 21004
rect 15844 20995 15896 21004
rect 15844 20961 15853 20995
rect 15853 20961 15887 20995
rect 15887 20961 15896 20995
rect 15844 20952 15896 20961
rect 17224 20995 17276 21004
rect 13820 20884 13872 20936
rect 14188 20884 14240 20936
rect 15660 20884 15712 20936
rect 9036 20816 9088 20825
rect 13544 20816 13596 20868
rect 17224 20961 17233 20995
rect 17233 20961 17267 20995
rect 17267 20961 17276 20995
rect 17224 20952 17276 20961
rect 17776 20995 17828 21004
rect 17776 20961 17785 20995
rect 17785 20961 17819 20995
rect 17819 20961 17828 20995
rect 18420 20995 18472 21004
rect 17776 20952 17828 20961
rect 18420 20961 18429 20995
rect 18429 20961 18463 20995
rect 18463 20961 18472 20995
rect 18420 20952 18472 20961
rect 19984 21029 19993 21063
rect 19993 21029 20027 21063
rect 20027 21029 20036 21063
rect 19984 21020 20036 21029
rect 20352 21063 20404 21072
rect 20352 21029 20361 21063
rect 20361 21029 20395 21063
rect 20395 21029 20404 21063
rect 20352 21020 20404 21029
rect 21364 21020 21416 21072
rect 19892 20995 19944 21004
rect 19432 20884 19484 20936
rect 19892 20961 19901 20995
rect 19901 20961 19935 20995
rect 19935 20961 19944 20995
rect 19892 20952 19944 20961
rect 20720 20952 20772 21004
rect 20536 20884 20588 20936
rect 21732 20995 21784 21004
rect 21732 20961 21741 20995
rect 21741 20961 21775 20995
rect 21775 20961 21784 20995
rect 24308 21020 24360 21072
rect 32128 21063 32180 21072
rect 21732 20952 21784 20961
rect 24032 20952 24084 21004
rect 24124 20952 24176 21004
rect 27528 20952 27580 21004
rect 32128 21029 32137 21063
rect 32137 21029 32171 21063
rect 32171 21029 32180 21063
rect 32128 21020 32180 21029
rect 32404 21020 32456 21072
rect 28908 20995 28960 21004
rect 22284 20884 22336 20936
rect 23480 20884 23532 20936
rect 23664 20884 23716 20936
rect 20444 20816 20496 20868
rect 28908 20961 28917 20995
rect 28917 20961 28951 20995
rect 28951 20961 28960 20995
rect 28908 20952 28960 20961
rect 29184 20995 29236 21004
rect 29184 20961 29193 20995
rect 29193 20961 29227 20995
rect 29227 20961 29236 20995
rect 29184 20952 29236 20961
rect 29276 20952 29328 21004
rect 30196 20952 30248 21004
rect 32036 20952 32088 21004
rect 32864 20952 32916 21004
rect 37556 21020 37608 21072
rect 33876 20995 33928 21004
rect 33876 20961 33885 20995
rect 33885 20961 33919 20995
rect 33919 20961 33928 20995
rect 33876 20952 33928 20961
rect 31760 20884 31812 20936
rect 32496 20884 32548 20936
rect 34152 20927 34204 20936
rect 34152 20893 34161 20927
rect 34161 20893 34195 20927
rect 34195 20893 34204 20927
rect 34152 20884 34204 20893
rect 34428 20952 34480 21004
rect 34704 20995 34756 21004
rect 34704 20961 34713 20995
rect 34713 20961 34747 20995
rect 34747 20961 34756 20995
rect 34704 20952 34756 20961
rect 35716 20952 35768 21004
rect 36636 20995 36688 21004
rect 36636 20961 36645 20995
rect 36645 20961 36679 20995
rect 36679 20961 36688 20995
rect 36636 20952 36688 20961
rect 37004 20995 37056 21004
rect 37004 20961 37013 20995
rect 37013 20961 37047 20995
rect 37047 20961 37056 20995
rect 37004 20952 37056 20961
rect 36820 20927 36872 20936
rect 36820 20893 36829 20927
rect 36829 20893 36863 20927
rect 36863 20893 36872 20927
rect 36820 20884 36872 20893
rect 7104 20791 7156 20800
rect 7104 20757 7113 20791
rect 7113 20757 7147 20791
rect 7147 20757 7156 20791
rect 7104 20748 7156 20757
rect 17224 20748 17276 20800
rect 22008 20748 22060 20800
rect 23020 20748 23072 20800
rect 28080 20748 28132 20800
rect 30196 20816 30248 20868
rect 30656 20748 30708 20800
rect 31668 20748 31720 20800
rect 4246 20646 4298 20698
rect 4310 20646 4362 20698
rect 4374 20646 4426 20698
rect 4438 20646 4490 20698
rect 34966 20646 35018 20698
rect 35030 20646 35082 20698
rect 35094 20646 35146 20698
rect 35158 20646 35210 20698
rect 3516 20544 3568 20596
rect 8944 20544 8996 20596
rect 14004 20587 14056 20596
rect 14004 20553 14013 20587
rect 14013 20553 14047 20587
rect 14047 20553 14056 20587
rect 14004 20544 14056 20553
rect 14556 20587 14608 20596
rect 14556 20553 14565 20587
rect 14565 20553 14599 20587
rect 14599 20553 14608 20587
rect 14556 20544 14608 20553
rect 14832 20544 14884 20596
rect 19340 20544 19392 20596
rect 20812 20544 20864 20596
rect 22928 20544 22980 20596
rect 24124 20544 24176 20596
rect 4988 20476 5040 20528
rect 7748 20476 7800 20528
rect 1584 20408 1636 20460
rect 7104 20451 7156 20460
rect 7104 20417 7113 20451
rect 7113 20417 7147 20451
rect 7147 20417 7156 20451
rect 7104 20408 7156 20417
rect 1400 20383 1452 20392
rect 1400 20349 1409 20383
rect 1409 20349 1443 20383
rect 1443 20349 1452 20383
rect 1400 20340 1452 20349
rect 3424 20340 3476 20392
rect 4712 20340 4764 20392
rect 4896 20383 4948 20392
rect 4896 20349 4905 20383
rect 4905 20349 4939 20383
rect 4939 20349 4948 20383
rect 4896 20340 4948 20349
rect 5264 20383 5316 20392
rect 5264 20349 5273 20383
rect 5273 20349 5307 20383
rect 5307 20349 5316 20383
rect 5264 20340 5316 20349
rect 5908 20383 5960 20392
rect 5908 20349 5917 20383
rect 5917 20349 5951 20383
rect 5951 20349 5960 20383
rect 5908 20340 5960 20349
rect 9036 20408 9088 20460
rect 9496 20451 9548 20460
rect 9496 20417 9505 20451
rect 9505 20417 9539 20451
rect 9539 20417 9548 20451
rect 9496 20408 9548 20417
rect 7288 20383 7340 20392
rect 7288 20349 7297 20383
rect 7297 20349 7331 20383
rect 7331 20349 7340 20383
rect 7288 20340 7340 20349
rect 8116 20383 8168 20392
rect 6368 20204 6420 20256
rect 8116 20349 8125 20383
rect 8125 20349 8159 20383
rect 8159 20349 8168 20383
rect 8116 20340 8168 20349
rect 8208 20340 8260 20392
rect 12440 20476 12492 20528
rect 15752 20519 15804 20528
rect 15752 20485 15761 20519
rect 15761 20485 15795 20519
rect 15795 20485 15804 20519
rect 15752 20476 15804 20485
rect 21272 20476 21324 20528
rect 21548 20476 21600 20528
rect 21732 20476 21784 20528
rect 20904 20408 20956 20460
rect 21364 20408 21416 20460
rect 11428 20383 11480 20392
rect 11428 20349 11437 20383
rect 11437 20349 11471 20383
rect 11471 20349 11480 20383
rect 11428 20340 11480 20349
rect 12532 20340 12584 20392
rect 14556 20340 14608 20392
rect 14740 20383 14792 20392
rect 14740 20349 14749 20383
rect 14749 20349 14783 20383
rect 14783 20349 14792 20383
rect 14740 20340 14792 20349
rect 14832 20383 14884 20392
rect 14832 20349 14841 20383
rect 14841 20349 14875 20383
rect 14875 20349 14884 20383
rect 15476 20383 15528 20392
rect 14832 20340 14884 20349
rect 15476 20349 15485 20383
rect 15485 20349 15519 20383
rect 15519 20349 15528 20383
rect 15476 20340 15528 20349
rect 16304 20383 16356 20392
rect 16304 20349 16313 20383
rect 16313 20349 16347 20383
rect 16347 20349 16356 20383
rect 16304 20340 16356 20349
rect 17040 20383 17092 20392
rect 17040 20349 17049 20383
rect 17049 20349 17083 20383
rect 17083 20349 17092 20383
rect 17040 20340 17092 20349
rect 18420 20340 18472 20392
rect 18788 20340 18840 20392
rect 19892 20340 19944 20392
rect 20444 20383 20496 20392
rect 20444 20349 20453 20383
rect 20453 20349 20487 20383
rect 20487 20349 20496 20383
rect 20444 20340 20496 20349
rect 20536 20340 20588 20392
rect 22744 20408 22796 20460
rect 27436 20544 27488 20596
rect 29644 20544 29696 20596
rect 30932 20544 30984 20596
rect 31576 20544 31628 20596
rect 37648 20587 37700 20596
rect 37648 20553 37657 20587
rect 37657 20553 37691 20587
rect 37691 20553 37700 20587
rect 37648 20544 37700 20553
rect 27804 20476 27856 20528
rect 35256 20476 35308 20528
rect 36268 20476 36320 20528
rect 27160 20408 27212 20460
rect 17684 20272 17736 20324
rect 22192 20272 22244 20324
rect 23572 20340 23624 20392
rect 23664 20383 23716 20392
rect 23664 20349 23673 20383
rect 23673 20349 23707 20383
rect 23707 20349 23716 20383
rect 23664 20340 23716 20349
rect 26056 20340 26108 20392
rect 26792 20340 26844 20392
rect 28172 20383 28224 20392
rect 28172 20349 28181 20383
rect 28181 20349 28215 20383
rect 28215 20349 28224 20383
rect 28172 20340 28224 20349
rect 28448 20383 28500 20392
rect 28448 20349 28457 20383
rect 28457 20349 28491 20383
rect 28491 20349 28500 20383
rect 28448 20340 28500 20349
rect 29276 20383 29328 20392
rect 29276 20349 29285 20383
rect 29285 20349 29319 20383
rect 29319 20349 29328 20383
rect 29276 20340 29328 20349
rect 30012 20383 30064 20392
rect 30012 20349 30021 20383
rect 30021 20349 30055 20383
rect 30055 20349 30064 20383
rect 30012 20340 30064 20349
rect 32312 20383 32364 20392
rect 32312 20349 32321 20383
rect 32321 20349 32355 20383
rect 32355 20349 32364 20383
rect 32312 20340 32364 20349
rect 30104 20272 30156 20324
rect 32128 20272 32180 20324
rect 33232 20340 33284 20392
rect 33968 20383 34020 20392
rect 33968 20349 33977 20383
rect 33977 20349 34011 20383
rect 34011 20349 34020 20383
rect 33968 20340 34020 20349
rect 35716 20383 35768 20392
rect 12440 20204 12492 20256
rect 17316 20204 17368 20256
rect 17868 20204 17920 20256
rect 18972 20204 19024 20256
rect 21456 20247 21508 20256
rect 21456 20213 21465 20247
rect 21465 20213 21499 20247
rect 21499 20213 21508 20247
rect 21456 20204 21508 20213
rect 22376 20204 22428 20256
rect 22928 20204 22980 20256
rect 23848 20204 23900 20256
rect 25872 20204 25924 20256
rect 27436 20204 27488 20256
rect 30380 20204 30432 20256
rect 32956 20204 33008 20256
rect 34428 20272 34480 20324
rect 35716 20349 35725 20383
rect 35725 20349 35759 20383
rect 35759 20349 35768 20383
rect 35716 20340 35768 20349
rect 36268 20383 36320 20392
rect 36268 20349 36277 20383
rect 36277 20349 36311 20383
rect 36311 20349 36320 20383
rect 36268 20340 36320 20349
rect 37832 20340 37884 20392
rect 34704 20204 34756 20256
rect 35348 20204 35400 20256
rect 35716 20204 35768 20256
rect 19606 20102 19658 20154
rect 19670 20102 19722 20154
rect 19734 20102 19786 20154
rect 19798 20102 19850 20154
rect 1952 19864 2004 19916
rect 2872 20000 2924 20052
rect 4620 20000 4672 20052
rect 11428 20000 11480 20052
rect 11888 20000 11940 20052
rect 12532 20000 12584 20052
rect 13452 20043 13504 20052
rect 13452 20009 13461 20043
rect 13461 20009 13495 20043
rect 13495 20009 13504 20043
rect 13452 20000 13504 20009
rect 4896 19932 4948 19984
rect 3148 19796 3200 19848
rect 4528 19864 4580 19916
rect 4712 19864 4764 19916
rect 6368 19907 6420 19916
rect 6368 19873 6377 19907
rect 6377 19873 6411 19907
rect 6411 19873 6420 19907
rect 6368 19864 6420 19873
rect 7288 19864 7340 19916
rect 8392 19932 8444 19984
rect 8944 19932 8996 19984
rect 9036 19907 9088 19916
rect 2964 19728 3016 19780
rect 7472 19796 7524 19848
rect 5264 19728 5316 19780
rect 7288 19728 7340 19780
rect 9036 19873 9045 19907
rect 9045 19873 9079 19907
rect 9079 19873 9088 19907
rect 9036 19864 9088 19873
rect 11888 19864 11940 19916
rect 12348 19907 12400 19916
rect 12348 19873 12357 19907
rect 12357 19873 12391 19907
rect 12391 19873 12400 19907
rect 12348 19864 12400 19873
rect 13544 19907 13596 19916
rect 13544 19873 13553 19907
rect 13553 19873 13587 19907
rect 13587 19873 13596 19907
rect 13544 19864 13596 19873
rect 14004 19907 14056 19916
rect 14004 19873 14013 19907
rect 14013 19873 14047 19907
rect 14047 19873 14056 19907
rect 14004 19864 14056 19873
rect 14096 19864 14148 19916
rect 17868 20000 17920 20052
rect 20260 20000 20312 20052
rect 15476 19907 15528 19916
rect 15476 19873 15485 19907
rect 15485 19873 15519 19907
rect 15519 19873 15528 19907
rect 15476 19864 15528 19873
rect 16304 19932 16356 19984
rect 20720 19932 20772 19984
rect 21180 19932 21232 19984
rect 23572 20000 23624 20052
rect 23848 20000 23900 20052
rect 16028 19864 16080 19916
rect 17592 19864 17644 19916
rect 18972 19907 19024 19916
rect 18972 19873 18981 19907
rect 18981 19873 19015 19907
rect 19015 19873 19024 19907
rect 18972 19864 19024 19873
rect 21916 19907 21968 19916
rect 21916 19873 21925 19907
rect 21925 19873 21959 19907
rect 21959 19873 21968 19907
rect 21916 19864 21968 19873
rect 22192 19864 22244 19916
rect 23940 19907 23992 19916
rect 23940 19873 23949 19907
rect 23949 19873 23983 19907
rect 23983 19873 23992 19907
rect 25136 19975 25188 19984
rect 25136 19941 25145 19975
rect 25145 19941 25179 19975
rect 25179 19941 25188 19975
rect 25136 19932 25188 19941
rect 26056 20000 26108 20052
rect 29184 20000 29236 20052
rect 29460 20000 29512 20052
rect 30380 20000 30432 20052
rect 32036 20000 32088 20052
rect 23940 19864 23992 19873
rect 27528 19932 27580 19984
rect 6276 19660 6328 19712
rect 11060 19796 11112 19848
rect 12440 19796 12492 19848
rect 18788 19796 18840 19848
rect 23112 19839 23164 19848
rect 23112 19805 23121 19839
rect 23121 19805 23155 19839
rect 23155 19805 23164 19839
rect 23112 19796 23164 19805
rect 26976 19864 27028 19916
rect 27252 19907 27304 19916
rect 27252 19873 27261 19907
rect 27261 19873 27295 19907
rect 27295 19873 27304 19907
rect 27252 19864 27304 19873
rect 27804 19907 27856 19916
rect 27804 19873 27813 19907
rect 27813 19873 27847 19907
rect 27847 19873 27856 19907
rect 27804 19864 27856 19873
rect 28080 19907 28132 19916
rect 28080 19873 28089 19907
rect 28089 19873 28123 19907
rect 28123 19873 28132 19907
rect 28080 19864 28132 19873
rect 29000 19932 29052 19984
rect 35992 20000 36044 20052
rect 20076 19728 20128 19780
rect 21456 19728 21508 19780
rect 22928 19728 22980 19780
rect 29644 19864 29696 19916
rect 32588 19932 32640 19984
rect 33416 19975 33468 19984
rect 33416 19941 33425 19975
rect 33425 19941 33459 19975
rect 33459 19941 33468 19975
rect 33416 19932 33468 19941
rect 35532 19975 35584 19984
rect 35532 19941 35541 19975
rect 35541 19941 35575 19975
rect 35575 19941 35584 19975
rect 35532 19932 35584 19941
rect 30104 19864 30156 19916
rect 31024 19864 31076 19916
rect 32772 19907 32824 19916
rect 32772 19873 32781 19907
rect 32781 19873 32815 19907
rect 32815 19873 32824 19907
rect 32772 19864 32824 19873
rect 32956 19907 33008 19916
rect 32956 19873 32965 19907
rect 32965 19873 32999 19907
rect 32999 19873 33008 19907
rect 32956 19864 33008 19873
rect 34152 19907 34204 19916
rect 34152 19873 34161 19907
rect 34161 19873 34195 19907
rect 34195 19873 34204 19907
rect 34152 19864 34204 19873
rect 36084 19907 36136 19916
rect 36084 19873 36093 19907
rect 36093 19873 36127 19907
rect 36127 19873 36136 19907
rect 36084 19864 36136 19873
rect 35256 19796 35308 19848
rect 36820 19864 36872 19916
rect 37280 19864 37332 19916
rect 9680 19660 9732 19712
rect 12532 19703 12584 19712
rect 12532 19669 12541 19703
rect 12541 19669 12575 19703
rect 12575 19669 12584 19703
rect 12532 19660 12584 19669
rect 13820 19660 13872 19712
rect 14740 19660 14792 19712
rect 16764 19660 16816 19712
rect 21180 19660 21232 19712
rect 25228 19660 25280 19712
rect 30472 19728 30524 19780
rect 36728 19728 36780 19780
rect 36912 19728 36964 19780
rect 30656 19660 30708 19712
rect 37004 19660 37056 19712
rect 4246 19558 4298 19610
rect 4310 19558 4362 19610
rect 4374 19558 4426 19610
rect 4438 19558 4490 19610
rect 34966 19558 35018 19610
rect 35030 19558 35082 19610
rect 35094 19558 35146 19610
rect 35158 19558 35210 19610
rect 4620 19499 4672 19508
rect 4620 19465 4629 19499
rect 4629 19465 4663 19499
rect 4663 19465 4672 19499
rect 4620 19456 4672 19465
rect 8208 19456 8260 19508
rect 11060 19456 11112 19508
rect 14832 19456 14884 19508
rect 25872 19456 25924 19508
rect 27160 19456 27212 19508
rect 4528 19388 4580 19440
rect 4712 19388 4764 19440
rect 6000 19388 6052 19440
rect 8024 19388 8076 19440
rect 18972 19388 19024 19440
rect 22192 19388 22244 19440
rect 7380 19363 7432 19372
rect 7380 19329 7389 19363
rect 7389 19329 7423 19363
rect 7423 19329 7432 19363
rect 7380 19320 7432 19329
rect 1400 19252 1452 19304
rect 2964 19252 3016 19304
rect 4528 19295 4580 19304
rect 4528 19261 4537 19295
rect 4537 19261 4571 19295
rect 4571 19261 4580 19295
rect 4528 19252 4580 19261
rect 5264 19295 5316 19304
rect 5264 19261 5273 19295
rect 5273 19261 5307 19295
rect 5307 19261 5316 19295
rect 5264 19252 5316 19261
rect 5448 19295 5500 19304
rect 5448 19261 5457 19295
rect 5457 19261 5491 19295
rect 5491 19261 5500 19295
rect 5448 19252 5500 19261
rect 4068 19184 4120 19236
rect 6460 19252 6512 19304
rect 7012 19295 7064 19304
rect 7012 19261 7021 19295
rect 7021 19261 7055 19295
rect 7055 19261 7064 19295
rect 7012 19252 7064 19261
rect 7288 19295 7340 19304
rect 7288 19261 7297 19295
rect 7297 19261 7331 19295
rect 7331 19261 7340 19295
rect 7288 19252 7340 19261
rect 7472 19252 7524 19304
rect 8392 19252 8444 19304
rect 8760 19252 8812 19304
rect 5908 19227 5960 19236
rect 5908 19193 5917 19227
rect 5917 19193 5951 19227
rect 5951 19193 5960 19227
rect 5908 19184 5960 19193
rect 6000 19184 6052 19236
rect 10600 19295 10652 19304
rect 10600 19261 10609 19295
rect 10609 19261 10643 19295
rect 10643 19261 10652 19295
rect 10600 19252 10652 19261
rect 13728 19320 13780 19372
rect 15936 19363 15988 19372
rect 11612 19295 11664 19304
rect 11612 19261 11621 19295
rect 11621 19261 11655 19295
rect 11655 19261 11664 19295
rect 11612 19252 11664 19261
rect 13544 19252 13596 19304
rect 14188 19295 14240 19304
rect 14188 19261 14197 19295
rect 14197 19261 14231 19295
rect 14231 19261 14240 19295
rect 14188 19252 14240 19261
rect 15200 19295 15252 19304
rect 15200 19261 15209 19295
rect 15209 19261 15243 19295
rect 15243 19261 15252 19295
rect 15200 19252 15252 19261
rect 15292 19252 15344 19304
rect 15936 19329 15945 19363
rect 15945 19329 15979 19363
rect 15979 19329 15988 19363
rect 15936 19320 15988 19329
rect 17316 19320 17368 19372
rect 20076 19320 20128 19372
rect 21180 19320 21232 19372
rect 21732 19320 21784 19372
rect 16396 19295 16448 19304
rect 16396 19261 16405 19295
rect 16405 19261 16439 19295
rect 16439 19261 16448 19295
rect 16396 19252 16448 19261
rect 16488 19295 16540 19304
rect 16488 19261 16497 19295
rect 16497 19261 16531 19295
rect 16531 19261 16540 19295
rect 17868 19295 17920 19304
rect 16488 19252 16540 19261
rect 17868 19261 17877 19295
rect 17877 19261 17911 19295
rect 17911 19261 17920 19295
rect 17868 19252 17920 19261
rect 18052 19295 18104 19304
rect 18052 19261 18061 19295
rect 18061 19261 18095 19295
rect 18095 19261 18104 19295
rect 18052 19252 18104 19261
rect 18236 19252 18288 19304
rect 20536 19252 20588 19304
rect 22008 19252 22060 19304
rect 16948 19227 17000 19236
rect 10232 19116 10284 19168
rect 16948 19193 16957 19227
rect 16957 19193 16991 19227
rect 16991 19193 17000 19227
rect 16948 19184 17000 19193
rect 17132 19184 17184 19236
rect 14280 19116 14332 19168
rect 18972 19116 19024 19168
rect 22100 19184 22152 19236
rect 28448 19456 28500 19508
rect 29184 19456 29236 19508
rect 32128 19456 32180 19508
rect 29000 19388 29052 19440
rect 30012 19388 30064 19440
rect 31024 19388 31076 19440
rect 26516 19320 26568 19372
rect 29092 19320 29144 19372
rect 29460 19320 29512 19372
rect 29644 19320 29696 19372
rect 30380 19320 30432 19372
rect 33324 19363 33376 19372
rect 33324 19329 33333 19363
rect 33333 19329 33367 19363
rect 33367 19329 33376 19363
rect 33324 19320 33376 19329
rect 36268 19320 36320 19372
rect 23296 19252 23348 19304
rect 24400 19295 24452 19304
rect 24400 19261 24409 19295
rect 24409 19261 24443 19295
rect 24443 19261 24452 19295
rect 24400 19252 24452 19261
rect 24860 19295 24912 19304
rect 24860 19261 24869 19295
rect 24869 19261 24903 19295
rect 24903 19261 24912 19295
rect 24860 19252 24912 19261
rect 25044 19295 25096 19304
rect 25044 19261 25053 19295
rect 25053 19261 25087 19295
rect 25087 19261 25096 19295
rect 25044 19252 25096 19261
rect 25136 19252 25188 19304
rect 26148 19295 26200 19304
rect 26148 19261 26157 19295
rect 26157 19261 26191 19295
rect 26191 19261 26200 19295
rect 26148 19252 26200 19261
rect 26884 19252 26936 19304
rect 27528 19295 27580 19304
rect 27528 19261 27537 19295
rect 27537 19261 27571 19295
rect 27571 19261 27580 19295
rect 27528 19252 27580 19261
rect 27896 19252 27948 19304
rect 28908 19252 28960 19304
rect 29368 19252 29420 19304
rect 24768 19184 24820 19236
rect 27252 19184 27304 19236
rect 30288 19184 30340 19236
rect 22284 19116 22336 19168
rect 22836 19116 22888 19168
rect 25964 19116 26016 19168
rect 26240 19159 26292 19168
rect 26240 19125 26249 19159
rect 26249 19125 26283 19159
rect 26283 19125 26292 19159
rect 26240 19116 26292 19125
rect 26976 19116 27028 19168
rect 27436 19116 27488 19168
rect 27712 19116 27764 19168
rect 29736 19116 29788 19168
rect 30196 19116 30248 19168
rect 31484 19295 31536 19304
rect 31484 19261 31493 19295
rect 31493 19261 31527 19295
rect 31527 19261 31536 19295
rect 31484 19252 31536 19261
rect 31760 19252 31812 19304
rect 32956 19295 33008 19304
rect 32956 19261 32965 19295
rect 32965 19261 32999 19295
rect 32999 19261 33008 19295
rect 32956 19252 33008 19261
rect 33140 19295 33192 19304
rect 33140 19261 33149 19295
rect 33149 19261 33183 19295
rect 33183 19261 33192 19295
rect 33140 19252 33192 19261
rect 33048 19184 33100 19236
rect 33600 19252 33652 19304
rect 34244 19252 34296 19304
rect 34980 19252 35032 19304
rect 35532 19252 35584 19304
rect 36544 19252 36596 19304
rect 37372 19252 37424 19304
rect 34704 19184 34756 19236
rect 32772 19116 32824 19168
rect 34796 19116 34848 19168
rect 19606 19014 19658 19066
rect 19670 19014 19722 19066
rect 19734 19014 19786 19066
rect 19798 19014 19850 19066
rect 3976 18912 4028 18964
rect 5908 18912 5960 18964
rect 6092 18912 6144 18964
rect 15476 18912 15528 18964
rect 2320 18819 2372 18828
rect 2320 18785 2329 18819
rect 2329 18785 2363 18819
rect 2363 18785 2372 18819
rect 2320 18776 2372 18785
rect 2688 18819 2740 18828
rect 2688 18785 2697 18819
rect 2697 18785 2731 18819
rect 2731 18785 2740 18819
rect 2688 18776 2740 18785
rect 3148 18776 3200 18828
rect 3424 18819 3476 18828
rect 3424 18785 3433 18819
rect 3433 18785 3467 18819
rect 3467 18785 3476 18819
rect 3424 18776 3476 18785
rect 5264 18819 5316 18828
rect 5264 18785 5273 18819
rect 5273 18785 5307 18819
rect 5307 18785 5316 18819
rect 5264 18776 5316 18785
rect 5632 18819 5684 18828
rect 5632 18785 5641 18819
rect 5641 18785 5675 18819
rect 5675 18785 5684 18819
rect 5632 18776 5684 18785
rect 5908 18776 5960 18828
rect 6184 18776 6236 18828
rect 7012 18776 7064 18828
rect 7472 18844 7524 18896
rect 13544 18887 13596 18896
rect 13544 18853 13553 18887
rect 13553 18853 13587 18887
rect 13587 18853 13596 18887
rect 13544 18844 13596 18853
rect 13728 18844 13780 18896
rect 7288 18776 7340 18828
rect 8392 18819 8444 18828
rect 8392 18785 8401 18819
rect 8401 18785 8435 18819
rect 8435 18785 8444 18819
rect 8392 18776 8444 18785
rect 9036 18776 9088 18828
rect 9680 18819 9732 18828
rect 9680 18785 9689 18819
rect 9689 18785 9723 18819
rect 9723 18785 9732 18819
rect 9680 18776 9732 18785
rect 10232 18819 10284 18828
rect 10232 18785 10241 18819
rect 10241 18785 10275 18819
rect 10275 18785 10284 18819
rect 10232 18776 10284 18785
rect 11704 18776 11756 18828
rect 11888 18819 11940 18828
rect 11888 18785 11897 18819
rect 11897 18785 11931 18819
rect 11931 18785 11940 18819
rect 11888 18776 11940 18785
rect 12532 18776 12584 18828
rect 14280 18819 14332 18828
rect 14280 18785 14289 18819
rect 14289 18785 14323 18819
rect 14323 18785 14332 18819
rect 14280 18776 14332 18785
rect 15292 18844 15344 18896
rect 16764 18844 16816 18896
rect 17960 18912 18012 18964
rect 19984 18844 20036 18896
rect 16028 18776 16080 18828
rect 17132 18819 17184 18828
rect 17132 18785 17141 18819
rect 17141 18785 17175 18819
rect 17175 18785 17184 18819
rect 17132 18776 17184 18785
rect 18880 18776 18932 18828
rect 19708 18819 19760 18828
rect 19708 18785 19717 18819
rect 19717 18785 19751 18819
rect 19751 18785 19760 18819
rect 19708 18776 19760 18785
rect 20720 18776 20772 18828
rect 22192 18912 22244 18964
rect 22284 18912 22336 18964
rect 20996 18887 21048 18896
rect 20996 18853 21005 18887
rect 21005 18853 21039 18887
rect 21039 18853 21048 18887
rect 20996 18844 21048 18853
rect 21088 18776 21140 18828
rect 21548 18819 21600 18828
rect 21548 18785 21557 18819
rect 21557 18785 21591 18819
rect 21591 18785 21600 18819
rect 21548 18776 21600 18785
rect 21916 18776 21968 18828
rect 23664 18776 23716 18828
rect 24400 18776 24452 18828
rect 24584 18844 24636 18896
rect 24860 18844 24912 18896
rect 26056 18844 26108 18896
rect 24768 18819 24820 18828
rect 24768 18785 24777 18819
rect 24777 18785 24811 18819
rect 24811 18785 24820 18819
rect 24768 18776 24820 18785
rect 25136 18819 25188 18828
rect 25136 18785 25145 18819
rect 25145 18785 25179 18819
rect 25179 18785 25188 18819
rect 25136 18776 25188 18785
rect 25872 18776 25924 18828
rect 29368 18844 29420 18896
rect 32956 18912 33008 18964
rect 29000 18776 29052 18828
rect 30196 18776 30248 18828
rect 31300 18776 31352 18828
rect 31484 18776 31536 18828
rect 2872 18751 2924 18760
rect 2872 18717 2881 18751
rect 2881 18717 2915 18751
rect 2915 18717 2924 18751
rect 2872 18708 2924 18717
rect 10600 18708 10652 18760
rect 11244 18708 11296 18760
rect 4620 18640 4672 18692
rect 11336 18640 11388 18692
rect 13912 18640 13964 18692
rect 18788 18708 18840 18760
rect 15568 18640 15620 18692
rect 17868 18640 17920 18692
rect 19248 18708 19300 18760
rect 19064 18640 19116 18692
rect 20352 18640 20404 18692
rect 22100 18708 22152 18760
rect 26976 18708 27028 18760
rect 27160 18751 27212 18760
rect 27160 18717 27169 18751
rect 27169 18717 27203 18751
rect 27203 18717 27212 18751
rect 27160 18708 27212 18717
rect 28356 18708 28408 18760
rect 29552 18751 29604 18760
rect 29552 18717 29561 18751
rect 29561 18717 29595 18751
rect 29595 18717 29604 18751
rect 29552 18708 29604 18717
rect 29644 18708 29696 18760
rect 34244 18844 34296 18896
rect 33324 18819 33376 18828
rect 33324 18785 33333 18819
rect 33333 18785 33367 18819
rect 33367 18785 33376 18819
rect 33324 18776 33376 18785
rect 33784 18776 33836 18828
rect 34980 18819 35032 18828
rect 23296 18683 23348 18692
rect 23296 18649 23305 18683
rect 23305 18649 23339 18683
rect 23339 18649 23348 18683
rect 23296 18640 23348 18649
rect 23572 18640 23624 18692
rect 30288 18640 30340 18692
rect 34152 18708 34204 18760
rect 34520 18751 34572 18760
rect 34520 18717 34529 18751
rect 34529 18717 34563 18751
rect 34563 18717 34572 18751
rect 34520 18708 34572 18717
rect 5632 18572 5684 18624
rect 7472 18572 7524 18624
rect 9772 18615 9824 18624
rect 9772 18581 9781 18615
rect 9781 18581 9815 18615
rect 9815 18581 9824 18615
rect 9772 18572 9824 18581
rect 11152 18615 11204 18624
rect 11152 18581 11161 18615
rect 11161 18581 11195 18615
rect 11195 18581 11204 18615
rect 11152 18572 11204 18581
rect 18604 18572 18656 18624
rect 19892 18615 19944 18624
rect 19892 18581 19901 18615
rect 19901 18581 19935 18615
rect 19935 18581 19944 18615
rect 19892 18572 19944 18581
rect 23204 18572 23256 18624
rect 27528 18572 27580 18624
rect 28540 18572 28592 18624
rect 28908 18572 28960 18624
rect 34704 18640 34756 18692
rect 34980 18785 34989 18819
rect 34989 18785 35023 18819
rect 35023 18785 35032 18819
rect 34980 18776 35032 18785
rect 35440 18776 35492 18828
rect 36452 18819 36504 18828
rect 36452 18785 36461 18819
rect 36461 18785 36495 18819
rect 36495 18785 36504 18819
rect 36452 18776 36504 18785
rect 37004 18819 37056 18828
rect 37004 18785 37013 18819
rect 37013 18785 37047 18819
rect 37047 18785 37056 18819
rect 37004 18776 37056 18785
rect 36268 18708 36320 18760
rect 35808 18640 35860 18692
rect 35532 18572 35584 18624
rect 35992 18572 36044 18624
rect 4246 18470 4298 18522
rect 4310 18470 4362 18522
rect 4374 18470 4426 18522
rect 4438 18470 4490 18522
rect 34966 18470 35018 18522
rect 35030 18470 35082 18522
rect 35094 18470 35146 18522
rect 35158 18470 35210 18522
rect 2688 18368 2740 18420
rect 5448 18411 5500 18420
rect 5448 18377 5457 18411
rect 5457 18377 5491 18411
rect 5491 18377 5500 18411
rect 5448 18368 5500 18377
rect 6092 18411 6144 18420
rect 6092 18377 6101 18411
rect 6101 18377 6135 18411
rect 6135 18377 6144 18411
rect 6092 18368 6144 18377
rect 6184 18368 6236 18420
rect 9036 18368 9088 18420
rect 11612 18368 11664 18420
rect 12348 18368 12400 18420
rect 12532 18368 12584 18420
rect 16396 18368 16448 18420
rect 19064 18368 19116 18420
rect 19708 18411 19760 18420
rect 19708 18377 19717 18411
rect 19717 18377 19751 18411
rect 19751 18377 19760 18411
rect 19708 18368 19760 18377
rect 22468 18368 22520 18420
rect 23204 18368 23256 18420
rect 27252 18368 27304 18420
rect 27344 18368 27396 18420
rect 36452 18368 36504 18420
rect 37740 18368 37792 18420
rect 2320 18232 2372 18284
rect 1400 18207 1452 18216
rect 1400 18173 1409 18207
rect 1409 18173 1443 18207
rect 1443 18173 1452 18207
rect 1400 18164 1452 18173
rect 3976 18164 4028 18216
rect 4712 18207 4764 18216
rect 4712 18173 4721 18207
rect 4721 18173 4755 18207
rect 4755 18173 4764 18207
rect 4712 18164 4764 18173
rect 19984 18300 20036 18352
rect 11152 18232 11204 18284
rect 11336 18232 11388 18284
rect 6276 18164 6328 18216
rect 7472 18207 7524 18216
rect 7472 18173 7481 18207
rect 7481 18173 7515 18207
rect 7515 18173 7524 18207
rect 7472 18164 7524 18173
rect 7748 18164 7800 18216
rect 8392 18207 8444 18216
rect 8392 18173 8401 18207
rect 8401 18173 8435 18207
rect 8435 18173 8444 18207
rect 8392 18164 8444 18173
rect 10140 18164 10192 18216
rect 12440 18207 12492 18216
rect 12440 18173 12449 18207
rect 12449 18173 12483 18207
rect 12483 18173 12492 18207
rect 12440 18164 12492 18173
rect 12624 18164 12676 18216
rect 13820 18207 13872 18216
rect 13820 18173 13829 18207
rect 13829 18173 13863 18207
rect 13863 18173 13872 18207
rect 13820 18164 13872 18173
rect 13912 18207 13964 18216
rect 13912 18173 13921 18207
rect 13921 18173 13955 18207
rect 13955 18173 13964 18207
rect 16120 18232 16172 18284
rect 18604 18275 18656 18284
rect 18604 18241 18613 18275
rect 18613 18241 18647 18275
rect 18647 18241 18656 18275
rect 18604 18232 18656 18241
rect 18788 18232 18840 18284
rect 20996 18232 21048 18284
rect 23204 18232 23256 18284
rect 13912 18164 13964 18173
rect 14556 18164 14608 18216
rect 16948 18164 17000 18216
rect 17132 18164 17184 18216
rect 18972 18164 19024 18216
rect 20812 18164 20864 18216
rect 22284 18164 22336 18216
rect 22744 18164 22796 18216
rect 22928 18207 22980 18216
rect 22928 18173 22937 18207
rect 22937 18173 22971 18207
rect 22971 18173 22980 18207
rect 22928 18164 22980 18173
rect 23020 18207 23072 18216
rect 23020 18173 23029 18207
rect 23029 18173 23063 18207
rect 23063 18173 23072 18207
rect 23664 18207 23716 18216
rect 23020 18164 23072 18173
rect 23664 18173 23673 18207
rect 23673 18173 23707 18207
rect 23707 18173 23716 18207
rect 23664 18164 23716 18173
rect 25504 18207 25556 18216
rect 5908 18096 5960 18148
rect 11244 18096 11296 18148
rect 6920 18071 6972 18080
rect 6920 18037 6929 18071
rect 6929 18037 6963 18071
rect 6963 18037 6972 18071
rect 6920 18028 6972 18037
rect 12716 18028 12768 18080
rect 17776 18096 17828 18148
rect 22468 18096 22520 18148
rect 22652 18096 22704 18148
rect 25504 18173 25513 18207
rect 25513 18173 25547 18207
rect 25547 18173 25556 18207
rect 25504 18164 25556 18173
rect 26240 18300 26292 18352
rect 29184 18300 29236 18352
rect 29552 18343 29604 18352
rect 29552 18309 29561 18343
rect 29561 18309 29595 18343
rect 29595 18309 29604 18343
rect 29552 18300 29604 18309
rect 30380 18300 30432 18352
rect 25872 18207 25924 18216
rect 25872 18173 25881 18207
rect 25881 18173 25915 18207
rect 25915 18173 25924 18207
rect 25872 18164 25924 18173
rect 27160 18207 27212 18216
rect 27160 18173 27169 18207
rect 27169 18173 27203 18207
rect 27203 18173 27212 18207
rect 27160 18164 27212 18173
rect 27344 18232 27396 18284
rect 28172 18232 28224 18284
rect 34152 18300 34204 18352
rect 36176 18300 36228 18352
rect 37556 18300 37608 18352
rect 27528 18164 27580 18216
rect 25044 18139 25096 18148
rect 25044 18105 25053 18139
rect 25053 18105 25087 18139
rect 25087 18105 25096 18139
rect 25044 18096 25096 18105
rect 25412 18096 25464 18148
rect 26056 18096 26108 18148
rect 34520 18232 34572 18284
rect 36728 18275 36780 18284
rect 36728 18241 36737 18275
rect 36737 18241 36771 18275
rect 36771 18241 36780 18275
rect 36728 18232 36780 18241
rect 29828 18207 29880 18216
rect 29828 18173 29837 18207
rect 29837 18173 29871 18207
rect 29871 18173 29880 18207
rect 29828 18164 29880 18173
rect 30196 18207 30248 18216
rect 30196 18173 30205 18207
rect 30205 18173 30239 18207
rect 30239 18173 30248 18207
rect 30196 18164 30248 18173
rect 32036 18207 32088 18216
rect 29736 18096 29788 18148
rect 17868 18028 17920 18080
rect 20536 18028 20588 18080
rect 21088 18071 21140 18080
rect 21088 18037 21097 18071
rect 21097 18037 21131 18071
rect 21131 18037 21140 18071
rect 21088 18028 21140 18037
rect 22100 18028 22152 18080
rect 22192 18028 22244 18080
rect 23020 18028 23072 18080
rect 23848 18071 23900 18080
rect 23848 18037 23857 18071
rect 23857 18037 23891 18071
rect 23891 18037 23900 18071
rect 23848 18028 23900 18037
rect 24492 18071 24544 18080
rect 24492 18037 24501 18071
rect 24501 18037 24535 18071
rect 24535 18037 24544 18071
rect 24492 18028 24544 18037
rect 27160 18028 27212 18080
rect 27804 18028 27856 18080
rect 32036 18173 32045 18207
rect 32045 18173 32079 18207
rect 32079 18173 32088 18207
rect 32036 18164 32088 18173
rect 32220 18207 32272 18216
rect 32220 18173 32229 18207
rect 32229 18173 32263 18207
rect 32263 18173 32272 18207
rect 32220 18164 32272 18173
rect 32312 18207 32364 18216
rect 32312 18173 32321 18207
rect 32321 18173 32355 18207
rect 32355 18173 32364 18207
rect 32312 18164 32364 18173
rect 32772 18207 32824 18216
rect 31760 18096 31812 18148
rect 32772 18173 32781 18207
rect 32781 18173 32815 18207
rect 32815 18173 32824 18207
rect 32772 18164 32824 18173
rect 33140 18164 33192 18216
rect 34704 18164 34756 18216
rect 36268 18164 36320 18216
rect 32588 18028 32640 18080
rect 34980 18071 35032 18080
rect 34980 18037 34989 18071
rect 34989 18037 35023 18071
rect 35023 18037 35032 18071
rect 34980 18028 35032 18037
rect 36268 18028 36320 18080
rect 36544 18164 36596 18216
rect 19606 17926 19658 17978
rect 19670 17926 19722 17978
rect 19734 17926 19786 17978
rect 19798 17926 19850 17978
rect 3424 17867 3476 17876
rect 3424 17833 3433 17867
rect 3433 17833 3467 17867
rect 3467 17833 3476 17867
rect 3424 17824 3476 17833
rect 8392 17824 8444 17876
rect 12624 17824 12676 17876
rect 19984 17824 20036 17876
rect 20720 17824 20772 17876
rect 24400 17824 24452 17876
rect 25964 17824 26016 17876
rect 28816 17824 28868 17876
rect 29276 17824 29328 17876
rect 30104 17824 30156 17876
rect 32036 17824 32088 17876
rect 33968 17824 34020 17876
rect 7012 17799 7064 17808
rect 7012 17765 7021 17799
rect 7021 17765 7055 17799
rect 7055 17765 7064 17799
rect 7012 17756 7064 17765
rect 4620 17688 4672 17740
rect 5448 17688 5500 17740
rect 5908 17688 5960 17740
rect 1400 17620 1452 17672
rect 2136 17663 2188 17672
rect 2136 17629 2145 17663
rect 2145 17629 2179 17663
rect 2179 17629 2188 17663
rect 2136 17620 2188 17629
rect 5356 17663 5408 17672
rect 5356 17629 5365 17663
rect 5365 17629 5399 17663
rect 5399 17629 5408 17663
rect 5356 17620 5408 17629
rect 8392 17688 8444 17740
rect 9772 17688 9824 17740
rect 12532 17731 12584 17740
rect 9680 17620 9732 17672
rect 10140 17663 10192 17672
rect 10140 17629 10149 17663
rect 10149 17629 10183 17663
rect 10183 17629 10192 17663
rect 10140 17620 10192 17629
rect 11888 17620 11940 17672
rect 12532 17697 12541 17731
rect 12541 17697 12575 17731
rect 12575 17697 12584 17731
rect 12532 17688 12584 17697
rect 15292 17688 15344 17740
rect 15660 17731 15712 17740
rect 15660 17697 15669 17731
rect 15669 17697 15703 17731
rect 15703 17697 15712 17731
rect 15660 17688 15712 17697
rect 16120 17731 16172 17740
rect 16120 17697 16129 17731
rect 16129 17697 16163 17731
rect 16163 17697 16172 17731
rect 16120 17688 16172 17697
rect 18604 17756 18656 17808
rect 17224 17731 17276 17740
rect 17224 17697 17233 17731
rect 17233 17697 17267 17731
rect 17267 17697 17276 17731
rect 17224 17688 17276 17697
rect 17316 17688 17368 17740
rect 18696 17688 18748 17740
rect 23480 17756 23532 17808
rect 27068 17799 27120 17808
rect 20444 17688 20496 17740
rect 22284 17688 22336 17740
rect 22928 17688 22980 17740
rect 23204 17731 23256 17740
rect 23204 17697 23213 17731
rect 23213 17697 23247 17731
rect 23247 17697 23256 17731
rect 23204 17688 23256 17697
rect 23664 17688 23716 17740
rect 24124 17688 24176 17740
rect 24584 17688 24636 17740
rect 24860 17731 24912 17740
rect 8944 17552 8996 17604
rect 3700 17484 3752 17536
rect 7840 17527 7892 17536
rect 7840 17493 7849 17527
rect 7849 17493 7883 17527
rect 7883 17493 7892 17527
rect 7840 17484 7892 17493
rect 12716 17484 12768 17536
rect 13820 17527 13872 17536
rect 13820 17493 13829 17527
rect 13829 17493 13863 17527
rect 13863 17493 13872 17527
rect 13820 17484 13872 17493
rect 14648 17620 14700 17672
rect 19064 17620 19116 17672
rect 23388 17620 23440 17672
rect 23848 17620 23900 17672
rect 24860 17697 24869 17731
rect 24869 17697 24903 17731
rect 24903 17697 24912 17731
rect 24860 17688 24912 17697
rect 25688 17731 25740 17740
rect 25688 17697 25697 17731
rect 25697 17697 25731 17731
rect 25731 17697 25740 17731
rect 25688 17688 25740 17697
rect 26516 17731 26568 17740
rect 26516 17697 26525 17731
rect 26525 17697 26559 17731
rect 26559 17697 26568 17731
rect 26516 17688 26568 17697
rect 27068 17765 27077 17799
rect 27077 17765 27111 17799
rect 27111 17765 27120 17799
rect 27068 17756 27120 17765
rect 27620 17688 27672 17740
rect 28632 17731 28684 17740
rect 28632 17697 28641 17731
rect 28641 17697 28675 17731
rect 28675 17697 28684 17731
rect 28632 17688 28684 17697
rect 28816 17688 28868 17740
rect 29368 17688 29420 17740
rect 30472 17731 30524 17740
rect 30472 17697 30481 17731
rect 30481 17697 30515 17731
rect 30515 17697 30524 17731
rect 30472 17688 30524 17697
rect 25780 17620 25832 17672
rect 26240 17620 26292 17672
rect 29000 17620 29052 17672
rect 31024 17731 31076 17740
rect 31024 17697 31033 17731
rect 31033 17697 31067 17731
rect 31067 17697 31076 17731
rect 31024 17688 31076 17697
rect 31208 17731 31260 17740
rect 31208 17697 31217 17731
rect 31217 17697 31251 17731
rect 31251 17697 31260 17731
rect 33048 17756 33100 17808
rect 33784 17799 33836 17808
rect 33784 17765 33793 17799
rect 33793 17765 33827 17799
rect 33827 17765 33836 17799
rect 33784 17756 33836 17765
rect 37280 17756 37332 17808
rect 31208 17688 31260 17697
rect 32772 17731 32824 17740
rect 32772 17697 32781 17731
rect 32781 17697 32815 17731
rect 32815 17697 32824 17731
rect 32772 17688 32824 17697
rect 30748 17620 30800 17672
rect 31300 17620 31352 17672
rect 34428 17688 34480 17740
rect 34796 17731 34848 17740
rect 34796 17697 34805 17731
rect 34805 17697 34839 17731
rect 34839 17697 34848 17731
rect 34796 17688 34848 17697
rect 34980 17688 35032 17740
rect 34336 17663 34388 17672
rect 34336 17629 34345 17663
rect 34345 17629 34379 17663
rect 34379 17629 34388 17663
rect 34336 17620 34388 17629
rect 15476 17552 15528 17604
rect 17684 17595 17736 17604
rect 17684 17561 17693 17595
rect 17693 17561 17727 17595
rect 17727 17561 17736 17595
rect 17684 17552 17736 17561
rect 17776 17552 17828 17604
rect 18144 17552 18196 17604
rect 21180 17552 21232 17604
rect 21732 17552 21784 17604
rect 23296 17552 23348 17604
rect 24676 17552 24728 17604
rect 34612 17552 34664 17604
rect 19892 17484 19944 17536
rect 20168 17484 20220 17536
rect 20352 17484 20404 17536
rect 20904 17484 20956 17536
rect 21272 17484 21324 17536
rect 23572 17484 23624 17536
rect 25872 17527 25924 17536
rect 25872 17493 25881 17527
rect 25881 17493 25915 17527
rect 25915 17493 25924 17527
rect 25872 17484 25924 17493
rect 27896 17484 27948 17536
rect 30380 17484 30432 17536
rect 30564 17484 30616 17536
rect 34520 17484 34572 17536
rect 35716 17620 35768 17672
rect 36268 17484 36320 17536
rect 37832 17527 37884 17536
rect 37832 17493 37841 17527
rect 37841 17493 37875 17527
rect 37875 17493 37884 17527
rect 37832 17484 37884 17493
rect 4246 17382 4298 17434
rect 4310 17382 4362 17434
rect 4374 17382 4426 17434
rect 4438 17382 4490 17434
rect 34966 17382 35018 17434
rect 35030 17382 35082 17434
rect 35094 17382 35146 17434
rect 35158 17382 35210 17434
rect 2136 17323 2188 17332
rect 2136 17289 2145 17323
rect 2145 17289 2179 17323
rect 2179 17289 2188 17323
rect 2136 17280 2188 17289
rect 6000 17280 6052 17332
rect 23572 17280 23624 17332
rect 24400 17280 24452 17332
rect 27896 17323 27948 17332
rect 2872 17119 2924 17128
rect 2872 17085 2881 17119
rect 2881 17085 2915 17119
rect 2915 17085 2924 17119
rect 2872 17076 2924 17085
rect 3700 17119 3752 17128
rect 3700 17085 3709 17119
rect 3709 17085 3743 17119
rect 3743 17085 3752 17119
rect 3700 17076 3752 17085
rect 4988 17119 5040 17128
rect 4988 17085 4997 17119
rect 4997 17085 5031 17119
rect 5031 17085 5040 17119
rect 4988 17076 5040 17085
rect 5632 17144 5684 17196
rect 5908 17144 5960 17196
rect 6920 17076 6972 17128
rect 8668 17144 8720 17196
rect 7748 17119 7800 17128
rect 7748 17085 7757 17119
rect 7757 17085 7791 17119
rect 7791 17085 7800 17119
rect 7748 17076 7800 17085
rect 8024 17119 8076 17128
rect 8024 17085 8033 17119
rect 8033 17085 8067 17119
rect 8067 17085 8076 17119
rect 8024 17076 8076 17085
rect 9864 17119 9916 17128
rect 9864 17085 9873 17119
rect 9873 17085 9907 17119
rect 9907 17085 9916 17119
rect 9864 17076 9916 17085
rect 12348 17212 12400 17264
rect 12716 17212 12768 17264
rect 16120 17212 16172 17264
rect 20444 17255 20496 17264
rect 10692 17187 10744 17196
rect 10692 17153 10701 17187
rect 10701 17153 10735 17187
rect 10735 17153 10744 17187
rect 10692 17144 10744 17153
rect 14648 17144 14700 17196
rect 15108 17187 15160 17196
rect 15108 17153 15117 17187
rect 15117 17153 15151 17187
rect 15151 17153 15160 17187
rect 15108 17144 15160 17153
rect 20444 17221 20453 17255
rect 20453 17221 20487 17255
rect 20487 17221 20496 17255
rect 20444 17212 20496 17221
rect 21088 17212 21140 17264
rect 11060 17076 11112 17128
rect 13636 17119 13688 17128
rect 5908 17051 5960 17060
rect 5908 17017 5917 17051
rect 5917 17017 5951 17051
rect 5951 17017 5960 17051
rect 5908 17008 5960 17017
rect 7196 16983 7248 16992
rect 7196 16949 7205 16983
rect 7205 16949 7239 16983
rect 7239 16949 7248 16983
rect 7196 16940 7248 16949
rect 7564 16940 7616 16992
rect 12624 17008 12676 17060
rect 13636 17085 13645 17119
rect 13645 17085 13679 17119
rect 13679 17085 13688 17119
rect 13636 17076 13688 17085
rect 13820 17119 13872 17128
rect 13820 17085 13829 17119
rect 13829 17085 13863 17119
rect 13863 17085 13872 17119
rect 13820 17076 13872 17085
rect 14188 17076 14240 17128
rect 16120 17076 16172 17128
rect 17132 17076 17184 17128
rect 17316 17076 17368 17128
rect 18052 17119 18104 17128
rect 18052 17085 18061 17119
rect 18061 17085 18095 17119
rect 18095 17085 18104 17119
rect 18052 17076 18104 17085
rect 18144 17119 18196 17128
rect 18144 17085 18153 17119
rect 18153 17085 18187 17119
rect 18187 17085 18196 17119
rect 18144 17076 18196 17085
rect 19340 17119 19392 17128
rect 9772 16940 9824 16992
rect 12440 16940 12492 16992
rect 16120 16940 16172 16992
rect 18512 17008 18564 17060
rect 18972 17008 19024 17060
rect 18144 16940 18196 16992
rect 19340 17085 19349 17119
rect 19349 17085 19383 17119
rect 19383 17085 19392 17119
rect 19340 17076 19392 17085
rect 21180 17119 21232 17128
rect 21180 17085 21189 17119
rect 21189 17085 21223 17119
rect 21223 17085 21232 17119
rect 21180 17076 21232 17085
rect 20168 16940 20220 16992
rect 20536 16940 20588 16992
rect 21824 17212 21876 17264
rect 22192 17212 22244 17264
rect 24860 17255 24912 17264
rect 24860 17221 24869 17255
rect 24869 17221 24903 17255
rect 24903 17221 24912 17255
rect 24860 17212 24912 17221
rect 26516 17212 26568 17264
rect 27896 17289 27905 17323
rect 27905 17289 27939 17323
rect 27939 17289 27948 17323
rect 27896 17280 27948 17289
rect 28356 17323 28408 17332
rect 28356 17289 28365 17323
rect 28365 17289 28399 17323
rect 28399 17289 28408 17323
rect 28356 17280 28408 17289
rect 29000 17280 29052 17332
rect 37832 17280 37884 17332
rect 30656 17212 30708 17264
rect 31116 17212 31168 17264
rect 33324 17212 33376 17264
rect 22008 17119 22060 17128
rect 22008 17085 22017 17119
rect 22017 17085 22051 17119
rect 22051 17085 22060 17119
rect 22008 17076 22060 17085
rect 22652 17076 22704 17128
rect 23756 17076 23808 17128
rect 23848 17076 23900 17128
rect 24492 17119 24544 17128
rect 24492 17085 24501 17119
rect 24501 17085 24535 17119
rect 24535 17085 24544 17119
rect 24492 17076 24544 17085
rect 24952 17076 25004 17128
rect 25780 17119 25832 17128
rect 25780 17085 25789 17119
rect 25789 17085 25823 17119
rect 25823 17085 25832 17119
rect 25780 17076 25832 17085
rect 26424 17144 26476 17196
rect 29828 17144 29880 17196
rect 26516 17119 26568 17128
rect 26516 17085 26525 17119
rect 26525 17085 26559 17119
rect 26559 17085 26568 17119
rect 26516 17076 26568 17085
rect 26700 17119 26752 17128
rect 26700 17085 26709 17119
rect 26709 17085 26743 17119
rect 26743 17085 26752 17119
rect 26700 17076 26752 17085
rect 28172 17119 28224 17128
rect 24400 17008 24452 17060
rect 28172 17085 28181 17119
rect 28181 17085 28215 17119
rect 28215 17085 28224 17119
rect 28172 17076 28224 17085
rect 28264 17076 28316 17128
rect 29644 17076 29696 17128
rect 30104 17119 30156 17128
rect 28356 17008 28408 17060
rect 23940 16940 23992 16992
rect 24584 16940 24636 16992
rect 27436 16940 27488 16992
rect 30104 17085 30113 17119
rect 30113 17085 30147 17119
rect 30147 17085 30156 17119
rect 30104 17076 30156 17085
rect 31208 17144 31260 17196
rect 30564 17076 30616 17128
rect 30656 17008 30708 17060
rect 31024 17076 31076 17128
rect 31760 17119 31812 17128
rect 31760 17085 31769 17119
rect 31769 17085 31803 17119
rect 31803 17085 31812 17119
rect 33508 17144 33560 17196
rect 31760 17076 31812 17085
rect 32956 17008 33008 17060
rect 34336 17076 34388 17128
rect 37740 17144 37792 17196
rect 34796 16940 34848 16992
rect 35992 17076 36044 17128
rect 36268 17076 36320 17128
rect 36544 17008 36596 17060
rect 36084 16940 36136 16992
rect 19606 16838 19658 16890
rect 19670 16838 19722 16890
rect 19734 16838 19786 16890
rect 19798 16838 19850 16890
rect 3056 16736 3108 16788
rect 3148 16736 3200 16788
rect 1676 16643 1728 16652
rect 1676 16609 1685 16643
rect 1685 16609 1719 16643
rect 1719 16609 1728 16643
rect 1676 16600 1728 16609
rect 4160 16643 4212 16652
rect 4160 16609 4169 16643
rect 4169 16609 4203 16643
rect 4203 16609 4212 16643
rect 4160 16600 4212 16609
rect 5632 16668 5684 16720
rect 5540 16643 5592 16652
rect 1400 16575 1452 16584
rect 1400 16541 1409 16575
rect 1409 16541 1443 16575
rect 1443 16541 1452 16575
rect 1400 16532 1452 16541
rect 5540 16609 5549 16643
rect 5549 16609 5583 16643
rect 5583 16609 5592 16643
rect 5540 16600 5592 16609
rect 5448 16575 5500 16584
rect 5448 16541 5457 16575
rect 5457 16541 5491 16575
rect 5491 16541 5500 16575
rect 5448 16532 5500 16541
rect 8024 16736 8076 16788
rect 8944 16779 8996 16788
rect 8944 16745 8953 16779
rect 8953 16745 8987 16779
rect 8987 16745 8996 16779
rect 8944 16736 8996 16745
rect 5908 16668 5960 16720
rect 12808 16736 12860 16788
rect 6000 16643 6052 16652
rect 6000 16609 6009 16643
rect 6009 16609 6043 16643
rect 6043 16609 6052 16643
rect 6000 16600 6052 16609
rect 7564 16600 7616 16652
rect 7104 16575 7156 16584
rect 7104 16541 7113 16575
rect 7113 16541 7147 16575
rect 7147 16541 7156 16575
rect 7104 16532 7156 16541
rect 9772 16643 9824 16652
rect 9772 16609 9781 16643
rect 9781 16609 9815 16643
rect 9815 16609 9824 16643
rect 9772 16600 9824 16609
rect 11244 16668 11296 16720
rect 9680 16575 9732 16584
rect 9680 16541 9689 16575
rect 9689 16541 9723 16575
rect 9723 16541 9732 16575
rect 9680 16532 9732 16541
rect 11428 16643 11480 16652
rect 11428 16609 11437 16643
rect 11437 16609 11471 16643
rect 11471 16609 11480 16643
rect 11428 16600 11480 16609
rect 12440 16600 12492 16652
rect 12716 16643 12768 16652
rect 12716 16609 12725 16643
rect 12725 16609 12759 16643
rect 12759 16609 12768 16643
rect 12716 16600 12768 16609
rect 21272 16736 21324 16788
rect 25780 16779 25832 16788
rect 25780 16745 25789 16779
rect 25789 16745 25823 16779
rect 25823 16745 25832 16779
rect 25780 16736 25832 16745
rect 26148 16736 26200 16788
rect 14372 16643 14424 16652
rect 14372 16609 14381 16643
rect 14381 16609 14415 16643
rect 14415 16609 14424 16643
rect 14372 16600 14424 16609
rect 16120 16643 16172 16652
rect 16120 16609 16129 16643
rect 16129 16609 16163 16643
rect 16163 16609 16172 16643
rect 16120 16600 16172 16609
rect 16396 16643 16448 16652
rect 16396 16609 16405 16643
rect 16405 16609 16439 16643
rect 16439 16609 16448 16643
rect 16396 16600 16448 16609
rect 16488 16600 16540 16652
rect 11060 16575 11112 16584
rect 11060 16541 11069 16575
rect 11069 16541 11103 16575
rect 11103 16541 11112 16575
rect 11060 16532 11112 16541
rect 18512 16600 18564 16652
rect 22008 16668 22060 16720
rect 23572 16668 23624 16720
rect 30840 16736 30892 16788
rect 32588 16736 32640 16788
rect 20720 16600 20772 16652
rect 21088 16643 21140 16652
rect 21088 16609 21097 16643
rect 21097 16609 21131 16643
rect 21131 16609 21140 16643
rect 21088 16600 21140 16609
rect 21180 16600 21232 16652
rect 21824 16643 21876 16652
rect 21824 16609 21833 16643
rect 21833 16609 21867 16643
rect 21867 16609 21876 16643
rect 21824 16600 21876 16609
rect 22192 16643 22244 16652
rect 11796 16464 11848 16516
rect 15292 16464 15344 16516
rect 1860 16396 1912 16448
rect 12624 16396 12676 16448
rect 16948 16396 17000 16448
rect 18052 16464 18104 16516
rect 19432 16532 19484 16584
rect 22192 16609 22201 16643
rect 22201 16609 22235 16643
rect 22235 16609 22244 16643
rect 22192 16600 22244 16609
rect 22468 16643 22520 16652
rect 22468 16609 22477 16643
rect 22477 16609 22511 16643
rect 22511 16609 22520 16643
rect 22468 16600 22520 16609
rect 23204 16643 23256 16652
rect 23204 16609 23213 16643
rect 23213 16609 23247 16643
rect 23247 16609 23256 16643
rect 23204 16600 23256 16609
rect 23664 16643 23716 16652
rect 23664 16609 23673 16643
rect 23673 16609 23707 16643
rect 23707 16609 23716 16643
rect 23664 16600 23716 16609
rect 24124 16643 24176 16652
rect 24124 16609 24133 16643
rect 24133 16609 24167 16643
rect 24167 16609 24176 16643
rect 24124 16600 24176 16609
rect 24676 16643 24728 16652
rect 24676 16609 24685 16643
rect 24685 16609 24719 16643
rect 24719 16609 24728 16643
rect 24676 16600 24728 16609
rect 24860 16643 24912 16652
rect 24860 16609 24869 16643
rect 24869 16609 24903 16643
rect 24903 16609 24912 16643
rect 24860 16600 24912 16609
rect 24952 16600 25004 16652
rect 25688 16600 25740 16652
rect 26516 16643 26568 16652
rect 26516 16609 26525 16643
rect 26525 16609 26559 16643
rect 26559 16609 26568 16643
rect 26516 16600 26568 16609
rect 30104 16668 30156 16720
rect 32036 16668 32088 16720
rect 19064 16464 19116 16516
rect 18144 16396 18196 16448
rect 18788 16396 18840 16448
rect 18972 16396 19024 16448
rect 23204 16464 23256 16516
rect 25504 16464 25556 16516
rect 27620 16600 27672 16652
rect 27804 16643 27856 16652
rect 27804 16609 27813 16643
rect 27813 16609 27847 16643
rect 27847 16609 27856 16643
rect 27804 16600 27856 16609
rect 28172 16575 28224 16584
rect 28172 16541 28181 16575
rect 28181 16541 28215 16575
rect 28215 16541 28224 16575
rect 29460 16600 29512 16652
rect 29644 16643 29696 16652
rect 29644 16609 29653 16643
rect 29653 16609 29687 16643
rect 29687 16609 29696 16643
rect 29644 16600 29696 16609
rect 31116 16643 31168 16652
rect 31116 16609 31125 16643
rect 31125 16609 31159 16643
rect 31159 16609 31168 16643
rect 31116 16600 31168 16609
rect 28172 16532 28224 16541
rect 29000 16532 29052 16584
rect 31668 16600 31720 16652
rect 35992 16736 36044 16788
rect 33048 16668 33100 16720
rect 26608 16439 26660 16448
rect 26608 16405 26617 16439
rect 26617 16405 26651 16439
rect 26651 16405 26660 16439
rect 26608 16396 26660 16405
rect 32496 16532 32548 16584
rect 33416 16600 33468 16652
rect 34520 16643 34572 16652
rect 34520 16609 34529 16643
rect 34529 16609 34563 16643
rect 34563 16609 34572 16643
rect 34520 16600 34572 16609
rect 34796 16643 34848 16652
rect 34796 16609 34805 16643
rect 34805 16609 34839 16643
rect 34839 16609 34848 16643
rect 34796 16600 34848 16609
rect 35440 16600 35492 16652
rect 33324 16575 33376 16584
rect 33324 16541 33333 16575
rect 33333 16541 33367 16575
rect 33367 16541 33376 16575
rect 33324 16532 33376 16541
rect 38108 16600 38160 16652
rect 33508 16464 33560 16516
rect 33968 16507 34020 16516
rect 33968 16473 33977 16507
rect 33977 16473 34011 16507
rect 34011 16473 34020 16507
rect 33968 16464 34020 16473
rect 29276 16396 29328 16448
rect 37924 16439 37976 16448
rect 37924 16405 37933 16439
rect 37933 16405 37967 16439
rect 37967 16405 37976 16439
rect 37924 16396 37976 16405
rect 4246 16294 4298 16346
rect 4310 16294 4362 16346
rect 4374 16294 4426 16346
rect 4438 16294 4490 16346
rect 34966 16294 35018 16346
rect 35030 16294 35082 16346
rect 35094 16294 35146 16346
rect 35158 16294 35210 16346
rect 4068 16192 4120 16244
rect 5540 16192 5592 16244
rect 8392 16235 8444 16244
rect 8392 16201 8401 16235
rect 8401 16201 8435 16235
rect 8435 16201 8444 16235
rect 8392 16192 8444 16201
rect 11244 16192 11296 16244
rect 11796 16235 11848 16244
rect 11796 16201 11805 16235
rect 11805 16201 11839 16235
rect 11839 16201 11848 16235
rect 11796 16192 11848 16201
rect 16120 16192 16172 16244
rect 18052 16192 18104 16244
rect 19248 16192 19300 16244
rect 20720 16192 20772 16244
rect 27436 16192 27488 16244
rect 1400 15988 1452 16040
rect 5356 16056 5408 16108
rect 7104 16099 7156 16108
rect 7104 16065 7113 16099
rect 7113 16065 7147 16099
rect 7147 16065 7156 16099
rect 7104 16056 7156 16065
rect 2688 15988 2740 16040
rect 4528 16031 4580 16040
rect 4528 15997 4537 16031
rect 4537 15997 4571 16031
rect 4571 15997 4580 16031
rect 4528 15988 4580 15997
rect 7748 15988 7800 16040
rect 9496 15988 9548 16040
rect 10692 16056 10744 16108
rect 10508 15988 10560 16040
rect 23112 16124 23164 16176
rect 11244 15988 11296 16040
rect 12440 15988 12492 16040
rect 12808 15988 12860 16040
rect 13912 16031 13964 16040
rect 13912 15997 13921 16031
rect 13921 15997 13955 16031
rect 13955 15997 13964 16031
rect 13912 15988 13964 15997
rect 15108 15988 15160 16040
rect 16028 16031 16080 16040
rect 16028 15997 16037 16031
rect 16037 15997 16071 16031
rect 16071 15997 16080 16031
rect 16028 15988 16080 15997
rect 17316 15988 17368 16040
rect 22652 16056 22704 16108
rect 24768 16099 24820 16108
rect 24768 16065 24777 16099
rect 24777 16065 24811 16099
rect 24811 16065 24820 16099
rect 24768 16056 24820 16065
rect 27068 16124 27120 16176
rect 27344 16124 27396 16176
rect 19064 16031 19116 16040
rect 19064 15997 19073 16031
rect 19073 15997 19107 16031
rect 19107 15997 19116 16031
rect 19064 15988 19116 15997
rect 20904 16031 20956 16040
rect 20904 15997 20913 16031
rect 20913 15997 20947 16031
rect 20947 15997 20956 16031
rect 20904 15988 20956 15997
rect 21456 16031 21508 16040
rect 9864 15852 9916 15904
rect 12348 15852 12400 15904
rect 18144 15920 18196 15972
rect 21456 15997 21465 16031
rect 21465 15997 21499 16031
rect 21499 15997 21508 16031
rect 21456 15988 21508 15997
rect 22192 15988 22244 16040
rect 24952 15988 25004 16040
rect 22100 15920 22152 15972
rect 23204 15920 23256 15972
rect 16856 15852 16908 15904
rect 19984 15852 20036 15904
rect 27344 15988 27396 16040
rect 27528 15988 27580 16040
rect 27988 15988 28040 16040
rect 30748 16192 30800 16244
rect 33048 16192 33100 16244
rect 36544 16235 36596 16244
rect 36544 16201 36553 16235
rect 36553 16201 36587 16235
rect 36587 16201 36596 16235
rect 36544 16192 36596 16201
rect 30196 16167 30248 16176
rect 30196 16133 30205 16167
rect 30205 16133 30239 16167
rect 30239 16133 30248 16167
rect 30196 16124 30248 16133
rect 31576 16056 31628 16108
rect 35716 16124 35768 16176
rect 34980 16099 35032 16108
rect 34980 16065 34989 16099
rect 34989 16065 35023 16099
rect 35023 16065 35032 16099
rect 34980 16056 35032 16065
rect 35992 16099 36044 16108
rect 29736 16031 29788 16040
rect 29736 15997 29745 16031
rect 29745 15997 29779 16031
rect 29779 15997 29788 16031
rect 29736 15988 29788 15997
rect 28540 15920 28592 15972
rect 29184 15920 29236 15972
rect 30196 15988 30248 16040
rect 31392 16031 31444 16040
rect 31392 15997 31401 16031
rect 31401 15997 31435 16031
rect 31435 15997 31444 16031
rect 31392 15988 31444 15997
rect 33324 16031 33376 16040
rect 33324 15997 33333 16031
rect 33333 15997 33367 16031
rect 33367 15997 33376 16031
rect 33324 15988 33376 15997
rect 33416 15988 33468 16040
rect 35992 16065 36001 16099
rect 36001 16065 36035 16099
rect 36035 16065 36044 16099
rect 35992 16056 36044 16065
rect 26792 15852 26844 15904
rect 27252 15895 27304 15904
rect 27252 15861 27261 15895
rect 27261 15861 27295 15895
rect 27295 15861 27304 15895
rect 27252 15852 27304 15861
rect 29368 15852 29420 15904
rect 35900 15988 35952 16040
rect 37280 16056 37332 16108
rect 37188 16031 37240 16040
rect 37188 15997 37197 16031
rect 37197 15997 37231 16031
rect 37231 15997 37240 16031
rect 37188 15988 37240 15997
rect 37372 15920 37424 15972
rect 37004 15852 37056 15904
rect 19606 15750 19658 15802
rect 19670 15750 19722 15802
rect 19734 15750 19786 15802
rect 19798 15750 19850 15802
rect 2688 15691 2740 15700
rect 2688 15657 2697 15691
rect 2697 15657 2731 15691
rect 2731 15657 2740 15691
rect 2688 15648 2740 15657
rect 4528 15648 4580 15700
rect 5632 15648 5684 15700
rect 4068 15580 4120 15632
rect 9588 15648 9640 15700
rect 10140 15648 10192 15700
rect 11428 15648 11480 15700
rect 16028 15648 16080 15700
rect 16304 15648 16356 15700
rect 19340 15648 19392 15700
rect 2964 15512 3016 15564
rect 3148 15555 3200 15564
rect 3148 15521 3157 15555
rect 3157 15521 3191 15555
rect 3191 15521 3200 15555
rect 3148 15512 3200 15521
rect 4712 15555 4764 15564
rect 1768 15444 1820 15496
rect 4712 15521 4721 15555
rect 4721 15521 4755 15555
rect 4755 15521 4764 15555
rect 4712 15512 4764 15521
rect 5632 15512 5684 15564
rect 7196 15512 7248 15564
rect 9496 15512 9548 15564
rect 5816 15444 5868 15496
rect 6276 15487 6328 15496
rect 6276 15453 6285 15487
rect 6285 15453 6319 15487
rect 6319 15453 6328 15487
rect 6276 15444 6328 15453
rect 9680 15444 9732 15496
rect 13268 15444 13320 15496
rect 14188 15555 14240 15564
rect 14188 15521 14197 15555
rect 14197 15521 14231 15555
rect 14231 15521 14240 15555
rect 14188 15512 14240 15521
rect 14004 15487 14056 15496
rect 14004 15453 14013 15487
rect 14013 15453 14047 15487
rect 14047 15453 14056 15487
rect 14004 15444 14056 15453
rect 16948 15555 17000 15564
rect 16488 15444 16540 15496
rect 16948 15521 16957 15555
rect 16957 15521 16991 15555
rect 16991 15521 17000 15555
rect 16948 15512 17000 15521
rect 17868 15555 17920 15564
rect 17132 15444 17184 15496
rect 17868 15521 17877 15555
rect 17877 15521 17911 15555
rect 17911 15521 17920 15555
rect 17868 15512 17920 15521
rect 18144 15555 18196 15564
rect 18144 15521 18153 15555
rect 18153 15521 18187 15555
rect 18187 15521 18196 15555
rect 18144 15512 18196 15521
rect 19800 15580 19852 15632
rect 18972 15555 19024 15564
rect 18972 15521 18981 15555
rect 18981 15521 19015 15555
rect 19015 15521 19024 15555
rect 18972 15512 19024 15521
rect 22836 15648 22888 15700
rect 22928 15648 22980 15700
rect 27436 15648 27488 15700
rect 29736 15691 29788 15700
rect 21180 15555 21232 15564
rect 21180 15521 21189 15555
rect 21189 15521 21223 15555
rect 21223 15521 21232 15555
rect 21180 15512 21232 15521
rect 21916 15512 21968 15564
rect 23204 15555 23256 15564
rect 23204 15521 23213 15555
rect 23213 15521 23247 15555
rect 23247 15521 23256 15555
rect 23204 15512 23256 15521
rect 24400 15512 24452 15564
rect 25504 15512 25556 15564
rect 25780 15555 25832 15564
rect 25780 15521 25789 15555
rect 25789 15521 25823 15555
rect 25823 15521 25832 15555
rect 25780 15512 25832 15521
rect 26608 15512 26660 15564
rect 27068 15555 27120 15564
rect 27068 15521 27077 15555
rect 27077 15521 27111 15555
rect 27111 15521 27120 15555
rect 27068 15512 27120 15521
rect 17960 15444 18012 15496
rect 18328 15444 18380 15496
rect 21824 15487 21876 15496
rect 16304 15376 16356 15428
rect 16580 15419 16632 15428
rect 16580 15385 16589 15419
rect 16589 15385 16623 15419
rect 16623 15385 16632 15419
rect 16580 15376 16632 15385
rect 16764 15376 16816 15428
rect 21824 15453 21833 15487
rect 21833 15453 21867 15487
rect 21867 15453 21876 15487
rect 21824 15444 21876 15453
rect 24952 15487 25004 15496
rect 24952 15453 24961 15487
rect 24961 15453 24995 15487
rect 24995 15453 25004 15487
rect 24952 15444 25004 15453
rect 26792 15444 26844 15496
rect 27528 15512 27580 15564
rect 29736 15657 29745 15691
rect 29745 15657 29779 15691
rect 29779 15657 29788 15691
rect 29736 15648 29788 15657
rect 32772 15648 32824 15700
rect 35900 15648 35952 15700
rect 28172 15580 28224 15632
rect 28540 15555 28592 15564
rect 22008 15376 22060 15428
rect 26700 15376 26752 15428
rect 28540 15521 28549 15555
rect 28549 15521 28583 15555
rect 28583 15521 28592 15555
rect 28540 15512 28592 15521
rect 29000 15555 29052 15564
rect 29000 15521 29009 15555
rect 29009 15521 29043 15555
rect 29043 15521 29052 15555
rect 29000 15512 29052 15521
rect 29368 15555 29420 15564
rect 29368 15521 29377 15555
rect 29377 15521 29411 15555
rect 29411 15521 29420 15555
rect 29368 15512 29420 15521
rect 29460 15512 29512 15564
rect 30748 15512 30800 15564
rect 30932 15580 30984 15632
rect 33416 15580 33468 15632
rect 33968 15580 34020 15632
rect 36912 15623 36964 15632
rect 30012 15444 30064 15496
rect 33048 15555 33100 15564
rect 33048 15521 33057 15555
rect 33057 15521 33091 15555
rect 33091 15521 33100 15555
rect 33048 15512 33100 15521
rect 34060 15555 34112 15564
rect 31392 15487 31444 15496
rect 31392 15453 31401 15487
rect 31401 15453 31435 15487
rect 31435 15453 31444 15487
rect 31392 15444 31444 15453
rect 32496 15444 32548 15496
rect 33324 15487 33376 15496
rect 33324 15453 33333 15487
rect 33333 15453 33367 15487
rect 33367 15453 33376 15487
rect 33324 15444 33376 15453
rect 34060 15521 34069 15555
rect 34069 15521 34103 15555
rect 34103 15521 34112 15555
rect 34060 15512 34112 15521
rect 36912 15589 36921 15623
rect 36921 15589 36955 15623
rect 36955 15589 36964 15623
rect 36912 15580 36964 15589
rect 35716 15555 35768 15564
rect 35716 15521 35725 15555
rect 35725 15521 35759 15555
rect 35759 15521 35768 15555
rect 35716 15512 35768 15521
rect 36636 15555 36688 15564
rect 35348 15444 35400 15496
rect 36636 15521 36645 15555
rect 36645 15521 36679 15555
rect 36679 15521 36688 15555
rect 36636 15512 36688 15521
rect 37280 15512 37332 15564
rect 37372 15444 37424 15496
rect 3792 15308 3844 15360
rect 11336 15308 11388 15360
rect 12532 15351 12584 15360
rect 12532 15317 12541 15351
rect 12541 15317 12575 15351
rect 12575 15317 12584 15351
rect 12532 15308 12584 15317
rect 23756 15308 23808 15360
rect 26608 15351 26660 15360
rect 26608 15317 26617 15351
rect 26617 15317 26651 15351
rect 26651 15317 26660 15351
rect 26608 15308 26660 15317
rect 35440 15308 35492 15360
rect 4246 15206 4298 15258
rect 4310 15206 4362 15258
rect 4374 15206 4426 15258
rect 4438 15206 4490 15258
rect 34966 15206 35018 15258
rect 35030 15206 35082 15258
rect 35094 15206 35146 15258
rect 35158 15206 35210 15258
rect 1676 15104 1728 15156
rect 1860 15036 1912 15088
rect 5356 15104 5408 15156
rect 14464 15104 14516 15156
rect 6000 15036 6052 15088
rect 6276 15036 6328 15088
rect 10232 15036 10284 15088
rect 2136 14943 2188 14952
rect 2136 14909 2145 14943
rect 2145 14909 2179 14943
rect 2179 14909 2188 14943
rect 2136 14900 2188 14909
rect 2780 14900 2832 14952
rect 4620 14968 4672 15020
rect 4160 14943 4212 14952
rect 4160 14909 4169 14943
rect 4169 14909 4203 14943
rect 4203 14909 4212 14943
rect 4160 14900 4212 14909
rect 7380 14968 7432 15020
rect 5632 14900 5684 14952
rect 6184 14900 6236 14952
rect 6828 14943 6880 14952
rect 6828 14909 6837 14943
rect 6837 14909 6871 14943
rect 6871 14909 6880 14943
rect 6828 14900 6880 14909
rect 7104 14900 7156 14952
rect 7564 14968 7616 15020
rect 10508 15011 10560 15020
rect 8024 14943 8076 14952
rect 6276 14832 6328 14884
rect 8024 14909 8033 14943
rect 8033 14909 8067 14943
rect 8067 14909 8076 14943
rect 8024 14900 8076 14909
rect 9036 14900 9088 14952
rect 9588 14900 9640 14952
rect 10140 14900 10192 14952
rect 10508 14977 10517 15011
rect 10517 14977 10551 15011
rect 10551 14977 10560 15011
rect 10508 14968 10560 14977
rect 12440 15036 12492 15088
rect 13268 15079 13320 15088
rect 13268 15045 13277 15079
rect 13277 15045 13311 15079
rect 13311 15045 13320 15079
rect 13268 15036 13320 15045
rect 15292 15011 15344 15020
rect 10876 14943 10928 14952
rect 10876 14909 10885 14943
rect 10885 14909 10919 14943
rect 10919 14909 10928 14943
rect 10876 14900 10928 14909
rect 7012 14807 7064 14816
rect 7012 14773 7021 14807
rect 7021 14773 7055 14807
rect 7055 14773 7064 14807
rect 7012 14764 7064 14773
rect 9772 14832 9824 14884
rect 9496 14764 9548 14816
rect 9588 14764 9640 14816
rect 12440 14900 12492 14952
rect 12808 14943 12860 14952
rect 12256 14832 12308 14884
rect 12808 14909 12817 14943
rect 12817 14909 12851 14943
rect 12851 14909 12860 14943
rect 12808 14900 12860 14909
rect 13268 14943 13320 14952
rect 13268 14909 13277 14943
rect 13277 14909 13311 14943
rect 13311 14909 13320 14943
rect 13268 14900 13320 14909
rect 15292 14977 15301 15011
rect 15301 14977 15335 15011
rect 15335 14977 15344 15011
rect 15292 14968 15344 14977
rect 16764 15104 16816 15156
rect 17040 15104 17092 15156
rect 23204 15104 23256 15156
rect 28356 15104 28408 15156
rect 34244 15104 34296 15156
rect 37372 15104 37424 15156
rect 16948 15036 17000 15088
rect 20904 15036 20956 15088
rect 21272 15036 21324 15088
rect 21824 15036 21876 15088
rect 16580 14968 16632 15020
rect 16764 14968 16816 15020
rect 19064 14968 19116 15020
rect 20352 14943 20404 14952
rect 14280 14832 14332 14884
rect 15108 14832 15160 14884
rect 17592 14832 17644 14884
rect 14188 14807 14240 14816
rect 14188 14773 14197 14807
rect 14197 14773 14231 14807
rect 14231 14773 14240 14807
rect 14188 14764 14240 14773
rect 14464 14764 14516 14816
rect 18420 14764 18472 14816
rect 19064 14832 19116 14884
rect 20352 14909 20361 14943
rect 20361 14909 20395 14943
rect 20395 14909 20404 14943
rect 20352 14900 20404 14909
rect 21640 14968 21692 15020
rect 21916 14968 21968 15020
rect 21732 14943 21784 14952
rect 21732 14909 21741 14943
rect 21741 14909 21775 14943
rect 21775 14909 21784 14943
rect 21732 14900 21784 14909
rect 19248 14832 19300 14884
rect 22100 14943 22152 14952
rect 22100 14909 22109 14943
rect 22109 14909 22143 14943
rect 22143 14909 22152 14943
rect 22468 14943 22520 14952
rect 22100 14900 22152 14909
rect 22468 14909 22477 14943
rect 22477 14909 22511 14943
rect 22511 14909 22520 14943
rect 22468 14900 22520 14909
rect 23296 14900 23348 14952
rect 23756 14900 23808 14952
rect 24400 14900 24452 14952
rect 28632 15036 28684 15088
rect 29184 15036 29236 15088
rect 29920 15036 29972 15088
rect 25964 15011 26016 15020
rect 25964 14977 25973 15011
rect 25973 14977 26007 15011
rect 26007 14977 26016 15011
rect 25964 14968 26016 14977
rect 27344 14968 27396 15020
rect 25688 14943 25740 14952
rect 22192 14832 22244 14884
rect 19432 14764 19484 14816
rect 22008 14764 22060 14816
rect 25688 14909 25697 14943
rect 25697 14909 25731 14943
rect 25731 14909 25740 14943
rect 25688 14900 25740 14909
rect 26608 14900 26660 14952
rect 26700 14900 26752 14952
rect 27436 14943 27488 14952
rect 27436 14909 27445 14943
rect 27445 14909 27479 14943
rect 27479 14909 27488 14943
rect 27436 14900 27488 14909
rect 30104 14968 30156 15020
rect 28172 14943 28224 14952
rect 28172 14909 28181 14943
rect 28181 14909 28215 14943
rect 28215 14909 28224 14943
rect 28172 14900 28224 14909
rect 29368 14900 29420 14952
rect 30196 14900 30248 14952
rect 30564 14943 30616 14952
rect 30564 14909 30573 14943
rect 30573 14909 30607 14943
rect 30607 14909 30616 14943
rect 30564 14900 30616 14909
rect 33048 14900 33100 14952
rect 33968 15036 34020 15088
rect 35532 15036 35584 15088
rect 33876 15011 33928 15020
rect 33876 14977 33885 15011
rect 33885 14977 33919 15011
rect 33919 14977 33928 15011
rect 33876 14968 33928 14977
rect 34520 14968 34572 15020
rect 35256 14968 35308 15020
rect 35992 14968 36044 15020
rect 23848 14807 23900 14816
rect 23848 14773 23857 14807
rect 23857 14773 23891 14807
rect 23891 14773 23900 14807
rect 23848 14764 23900 14773
rect 26516 14832 26568 14884
rect 27896 14832 27948 14884
rect 33968 14900 34020 14952
rect 34152 14943 34204 14952
rect 34152 14909 34161 14943
rect 34161 14909 34195 14943
rect 34195 14909 34204 14943
rect 34152 14900 34204 14909
rect 35440 14943 35492 14952
rect 35440 14909 35449 14943
rect 35449 14909 35483 14943
rect 35483 14909 35492 14943
rect 35440 14900 35492 14909
rect 35532 14900 35584 14952
rect 36268 14900 36320 14952
rect 36452 14943 36504 14952
rect 36452 14909 36461 14943
rect 36461 14909 36495 14943
rect 36495 14909 36504 14943
rect 36452 14900 36504 14909
rect 34520 14832 34572 14884
rect 27528 14764 27580 14816
rect 27620 14764 27672 14816
rect 30656 14764 30708 14816
rect 19606 14662 19658 14714
rect 19670 14662 19722 14714
rect 19734 14662 19786 14714
rect 19798 14662 19850 14714
rect 2780 14603 2832 14612
rect 2780 14569 2789 14603
rect 2789 14569 2823 14603
rect 2823 14569 2832 14603
rect 2780 14560 2832 14569
rect 1400 14399 1452 14408
rect 1400 14365 1409 14399
rect 1409 14365 1443 14399
rect 1443 14365 1452 14399
rect 1400 14356 1452 14365
rect 1676 14399 1728 14408
rect 1676 14365 1685 14399
rect 1685 14365 1719 14399
rect 1719 14365 1728 14399
rect 1676 14356 1728 14365
rect 3976 14424 4028 14476
rect 19248 14560 19300 14612
rect 4712 14424 4764 14476
rect 4988 14424 5040 14476
rect 7012 14492 7064 14544
rect 4160 14356 4212 14408
rect 5448 14356 5500 14408
rect 6920 14424 6972 14476
rect 10876 14492 10928 14544
rect 8944 14467 8996 14476
rect 7104 14356 7156 14408
rect 5080 14288 5132 14340
rect 8944 14433 8953 14467
rect 8953 14433 8987 14467
rect 8987 14433 8996 14467
rect 8944 14424 8996 14433
rect 9956 14424 10008 14476
rect 10232 14467 10284 14476
rect 10232 14433 10241 14467
rect 10241 14433 10275 14467
rect 10275 14433 10284 14467
rect 10232 14424 10284 14433
rect 10508 14467 10560 14476
rect 10508 14433 10517 14467
rect 10517 14433 10551 14467
rect 10551 14433 10560 14467
rect 10508 14424 10560 14433
rect 11336 14467 11388 14476
rect 11336 14433 11345 14467
rect 11345 14433 11379 14467
rect 11379 14433 11388 14467
rect 11336 14424 11388 14433
rect 11888 14467 11940 14476
rect 11888 14433 11897 14467
rect 11897 14433 11931 14467
rect 11931 14433 11940 14467
rect 11888 14424 11940 14433
rect 13268 14492 13320 14544
rect 14188 14492 14240 14544
rect 14004 14467 14056 14476
rect 8760 14356 8812 14408
rect 9864 14399 9916 14408
rect 9864 14365 9873 14399
rect 9873 14365 9907 14399
rect 9907 14365 9916 14399
rect 9864 14356 9916 14365
rect 13176 14399 13228 14408
rect 13176 14365 13185 14399
rect 13185 14365 13219 14399
rect 13219 14365 13228 14399
rect 13176 14356 13228 14365
rect 8484 14288 8536 14340
rect 9220 14288 9272 14340
rect 9680 14288 9732 14340
rect 11428 14288 11480 14340
rect 12348 14288 12400 14340
rect 14004 14433 14013 14467
rect 14013 14433 14047 14467
rect 14047 14433 14056 14467
rect 14004 14424 14056 14433
rect 15752 14467 15804 14476
rect 15752 14433 15761 14467
rect 15761 14433 15795 14467
rect 15795 14433 15804 14467
rect 15752 14424 15804 14433
rect 16120 14467 16172 14476
rect 16120 14433 16129 14467
rect 16129 14433 16163 14467
rect 16163 14433 16172 14467
rect 16120 14424 16172 14433
rect 18328 14492 18380 14544
rect 15844 14356 15896 14408
rect 17776 14424 17828 14476
rect 19340 14492 19392 14544
rect 19064 14467 19116 14476
rect 19064 14433 19073 14467
rect 19073 14433 19107 14467
rect 19107 14433 19116 14467
rect 19064 14424 19116 14433
rect 19156 14467 19208 14476
rect 19156 14433 19165 14467
rect 19165 14433 19199 14467
rect 19199 14433 19208 14467
rect 19800 14467 19852 14476
rect 19156 14424 19208 14433
rect 19800 14433 19809 14467
rect 19809 14433 19843 14467
rect 19843 14433 19852 14467
rect 19800 14424 19852 14433
rect 19892 14424 19944 14476
rect 22192 14560 22244 14612
rect 23388 14560 23440 14612
rect 25688 14560 25740 14612
rect 26148 14560 26200 14612
rect 27068 14560 27120 14612
rect 28632 14560 28684 14612
rect 21916 14492 21968 14544
rect 18052 14356 18104 14408
rect 19248 14356 19300 14408
rect 20444 14356 20496 14408
rect 13912 14331 13964 14340
rect 13912 14297 13921 14331
rect 13921 14297 13955 14331
rect 13955 14297 13964 14331
rect 13912 14288 13964 14297
rect 14280 14288 14332 14340
rect 17500 14288 17552 14340
rect 21824 14467 21876 14476
rect 21824 14433 21833 14467
rect 21833 14433 21867 14467
rect 21867 14433 21876 14467
rect 21824 14424 21876 14433
rect 22100 14424 22152 14476
rect 22284 14467 22336 14476
rect 22284 14433 22293 14467
rect 22293 14433 22327 14467
rect 22327 14433 22336 14467
rect 22284 14424 22336 14433
rect 22744 14424 22796 14476
rect 23388 14424 23440 14476
rect 22836 14399 22888 14408
rect 22836 14365 22845 14399
rect 22845 14365 22879 14399
rect 22879 14365 22888 14399
rect 22836 14356 22888 14365
rect 23204 14356 23256 14408
rect 23756 14424 23808 14476
rect 24124 14467 24176 14476
rect 24124 14433 24133 14467
rect 24133 14433 24167 14467
rect 24167 14433 24176 14467
rect 24124 14424 24176 14433
rect 24952 14424 25004 14476
rect 25964 14424 26016 14476
rect 27436 14492 27488 14544
rect 27344 14467 27396 14476
rect 27344 14433 27353 14467
rect 27353 14433 27387 14467
rect 27387 14433 27396 14467
rect 27344 14424 27396 14433
rect 27988 14424 28040 14476
rect 26792 14356 26844 14408
rect 30104 14560 30156 14612
rect 30564 14603 30616 14612
rect 30564 14569 30573 14603
rect 30573 14569 30607 14603
rect 30607 14569 30616 14603
rect 30564 14560 30616 14569
rect 32864 14603 32916 14612
rect 32864 14569 32873 14603
rect 32873 14569 32907 14603
rect 32907 14569 32916 14603
rect 32864 14560 32916 14569
rect 33968 14560 34020 14612
rect 29000 14424 29052 14476
rect 33508 14492 33560 14544
rect 29644 14467 29696 14476
rect 29644 14433 29653 14467
rect 29653 14433 29687 14467
rect 29687 14433 29696 14467
rect 29644 14424 29696 14433
rect 30380 14424 30432 14476
rect 30748 14467 30800 14476
rect 30748 14433 30757 14467
rect 30757 14433 30791 14467
rect 30791 14433 30800 14467
rect 30748 14424 30800 14433
rect 30932 14467 30984 14476
rect 30932 14433 30941 14467
rect 30941 14433 30975 14467
rect 30975 14433 30984 14467
rect 30932 14424 30984 14433
rect 32772 14424 32824 14476
rect 32956 14424 33008 14476
rect 34520 14492 34572 14544
rect 34796 14492 34848 14544
rect 35440 14492 35492 14544
rect 34704 14424 34756 14476
rect 35348 14424 35400 14476
rect 36268 14467 36320 14476
rect 36268 14433 36277 14467
rect 36277 14433 36311 14467
rect 36311 14433 36320 14467
rect 36268 14424 36320 14433
rect 36636 14467 36688 14476
rect 32220 14356 32272 14408
rect 34520 14356 34572 14408
rect 35716 14356 35768 14408
rect 36636 14433 36645 14467
rect 36645 14433 36679 14467
rect 36679 14433 36688 14467
rect 36636 14424 36688 14433
rect 23664 14288 23716 14340
rect 24032 14288 24084 14340
rect 27160 14288 27212 14340
rect 30472 14288 30524 14340
rect 34612 14288 34664 14340
rect 37188 14288 37240 14340
rect 1400 14220 1452 14272
rect 5816 14220 5868 14272
rect 16764 14220 16816 14272
rect 16948 14263 17000 14272
rect 16948 14229 16957 14263
rect 16957 14229 16991 14263
rect 16991 14229 17000 14263
rect 16948 14220 17000 14229
rect 17684 14220 17736 14272
rect 22928 14220 22980 14272
rect 28724 14220 28776 14272
rect 29552 14220 29604 14272
rect 32772 14220 32824 14272
rect 33508 14220 33560 14272
rect 4246 14118 4298 14170
rect 4310 14118 4362 14170
rect 4374 14118 4426 14170
rect 4438 14118 4490 14170
rect 34966 14118 35018 14170
rect 35030 14118 35082 14170
rect 35094 14118 35146 14170
rect 35158 14118 35210 14170
rect 2136 14016 2188 14068
rect 5356 14016 5408 14068
rect 1860 13923 1912 13932
rect 1860 13889 1869 13923
rect 1869 13889 1903 13923
rect 1903 13889 1912 13923
rect 1860 13880 1912 13889
rect 3976 13855 4028 13864
rect 3976 13821 3985 13855
rect 3985 13821 4019 13855
rect 4019 13821 4028 13855
rect 3976 13812 4028 13821
rect 4988 13855 5040 13864
rect 4988 13821 4997 13855
rect 4997 13821 5031 13855
rect 5031 13821 5040 13855
rect 4988 13812 5040 13821
rect 5448 13812 5500 13864
rect 5908 13855 5960 13864
rect 5908 13821 5917 13855
rect 5917 13821 5951 13855
rect 5951 13821 5960 13855
rect 5908 13812 5960 13821
rect 6920 13812 6972 13864
rect 8024 13991 8076 14000
rect 8024 13957 8033 13991
rect 8033 13957 8067 13991
rect 8067 13957 8076 13991
rect 8024 13948 8076 13957
rect 8944 14016 8996 14068
rect 16488 14016 16540 14068
rect 17132 14016 17184 14068
rect 17776 14016 17828 14068
rect 18972 14016 19024 14068
rect 21824 14016 21876 14068
rect 11428 13948 11480 14000
rect 13268 13991 13320 14000
rect 13268 13957 13277 13991
rect 13277 13957 13311 13991
rect 13311 13957 13320 13991
rect 13268 13948 13320 13957
rect 15292 13948 15344 14000
rect 19248 13948 19300 14000
rect 9772 13880 9824 13932
rect 4896 13744 4948 13796
rect 9588 13812 9640 13864
rect 10876 13880 10928 13932
rect 10692 13855 10744 13864
rect 10692 13821 10701 13855
rect 10701 13821 10735 13855
rect 10735 13821 10744 13855
rect 10692 13812 10744 13821
rect 11060 13855 11112 13864
rect 11060 13821 11069 13855
rect 11069 13821 11103 13855
rect 11103 13821 11112 13855
rect 11060 13812 11112 13821
rect 12716 13880 12768 13932
rect 14280 13923 14332 13932
rect 14280 13889 14289 13923
rect 14289 13889 14323 13923
rect 14323 13889 14332 13923
rect 14280 13880 14332 13889
rect 15108 13880 15160 13932
rect 12808 13855 12860 13864
rect 3332 13676 3384 13728
rect 12808 13821 12817 13855
rect 12817 13821 12851 13855
rect 12851 13821 12860 13855
rect 12808 13812 12860 13821
rect 13452 13812 13504 13864
rect 15016 13812 15068 13864
rect 17684 13812 17736 13864
rect 18328 13855 18380 13864
rect 18328 13821 18337 13855
rect 18337 13821 18371 13855
rect 18371 13821 18380 13855
rect 18328 13812 18380 13821
rect 18512 13880 18564 13932
rect 20444 13923 20496 13932
rect 20168 13855 20220 13864
rect 20168 13821 20177 13855
rect 20177 13821 20211 13855
rect 20211 13821 20220 13855
rect 20168 13812 20220 13821
rect 20444 13889 20453 13923
rect 20453 13889 20487 13923
rect 20487 13889 20496 13923
rect 20444 13880 20496 13889
rect 22376 13923 22428 13932
rect 22376 13889 22385 13923
rect 22385 13889 22419 13923
rect 22419 13889 22428 13923
rect 22376 13880 22428 13889
rect 23020 13880 23072 13932
rect 26240 14016 26292 14068
rect 28632 14059 28684 14068
rect 26792 13991 26844 14000
rect 26792 13957 26801 13991
rect 26801 13957 26835 13991
rect 26835 13957 26844 13991
rect 26792 13948 26844 13957
rect 28632 14025 28641 14059
rect 28641 14025 28675 14059
rect 28675 14025 28684 14059
rect 28632 14016 28684 14025
rect 29644 14016 29696 14068
rect 34336 14059 34388 14068
rect 34336 14025 34345 14059
rect 34345 14025 34379 14059
rect 34379 14025 34388 14059
rect 34336 14016 34388 14025
rect 36084 14016 36136 14068
rect 36452 14016 36504 14068
rect 23296 13812 23348 13864
rect 18144 13744 18196 13796
rect 17316 13676 17368 13728
rect 20076 13676 20128 13728
rect 21732 13676 21784 13728
rect 23480 13744 23532 13796
rect 23756 13812 23808 13864
rect 24584 13812 24636 13864
rect 25320 13812 25372 13864
rect 26240 13812 26292 13864
rect 25872 13744 25924 13796
rect 27068 13812 27120 13864
rect 28632 13812 28684 13864
rect 31392 13948 31444 14000
rect 30932 13880 30984 13932
rect 29828 13855 29880 13864
rect 29828 13821 29837 13855
rect 29837 13821 29871 13855
rect 29871 13821 29880 13855
rect 29828 13812 29880 13821
rect 30472 13855 30524 13864
rect 23572 13676 23624 13728
rect 23940 13676 23992 13728
rect 24860 13719 24912 13728
rect 24860 13685 24869 13719
rect 24869 13685 24903 13719
rect 24903 13685 24912 13719
rect 24860 13676 24912 13685
rect 25688 13676 25740 13728
rect 30472 13821 30481 13855
rect 30481 13821 30515 13855
rect 30515 13821 30524 13855
rect 30472 13812 30524 13821
rect 30288 13744 30340 13796
rect 32128 13855 32180 13864
rect 32128 13821 32137 13855
rect 32137 13821 32171 13855
rect 32171 13821 32180 13855
rect 32128 13812 32180 13821
rect 33784 13948 33836 14000
rect 36268 13948 36320 14000
rect 33232 13923 33284 13932
rect 33232 13889 33241 13923
rect 33241 13889 33275 13923
rect 33275 13889 33284 13923
rect 33232 13880 33284 13889
rect 32772 13855 32824 13864
rect 32772 13821 32781 13855
rect 32781 13821 32815 13855
rect 32815 13821 32824 13855
rect 32772 13812 32824 13821
rect 33324 13855 33376 13864
rect 33324 13821 33333 13855
rect 33333 13821 33367 13855
rect 33367 13821 33376 13855
rect 33324 13812 33376 13821
rect 33968 13880 34020 13932
rect 34244 13880 34296 13932
rect 35440 13923 35492 13932
rect 35440 13889 35449 13923
rect 35449 13889 35483 13923
rect 35483 13889 35492 13923
rect 35440 13880 35492 13889
rect 35992 13855 36044 13864
rect 35992 13821 36001 13855
rect 36001 13821 36035 13855
rect 36035 13821 36044 13855
rect 35992 13812 36044 13821
rect 36452 13855 36504 13864
rect 36452 13821 36461 13855
rect 36461 13821 36495 13855
rect 36495 13821 36504 13855
rect 36452 13812 36504 13821
rect 36544 13812 36596 13864
rect 30656 13676 30708 13728
rect 31392 13719 31444 13728
rect 31392 13685 31401 13719
rect 31401 13685 31435 13719
rect 31435 13685 31444 13719
rect 31392 13676 31444 13685
rect 31944 13719 31996 13728
rect 31944 13685 31953 13719
rect 31953 13685 31987 13719
rect 31987 13685 31996 13719
rect 31944 13676 31996 13685
rect 33692 13676 33744 13728
rect 19606 13574 19658 13626
rect 19670 13574 19722 13626
rect 19734 13574 19786 13626
rect 19798 13574 19850 13626
rect 1676 13515 1728 13524
rect 1676 13481 1685 13515
rect 1685 13481 1719 13515
rect 1719 13481 1728 13515
rect 1676 13472 1728 13481
rect 10692 13472 10744 13524
rect 10968 13472 11020 13524
rect 3976 13404 4028 13456
rect 1768 13379 1820 13388
rect 1768 13345 1777 13379
rect 1777 13345 1811 13379
rect 1811 13345 1820 13379
rect 1768 13336 1820 13345
rect 3332 13379 3384 13388
rect 3332 13345 3341 13379
rect 3341 13345 3375 13379
rect 3375 13345 3384 13379
rect 3332 13336 3384 13345
rect 4620 13336 4672 13388
rect 4896 13268 4948 13320
rect 6000 13336 6052 13388
rect 8668 13379 8720 13388
rect 6368 13311 6420 13320
rect 6368 13277 6377 13311
rect 6377 13277 6411 13311
rect 6411 13277 6420 13311
rect 6368 13268 6420 13277
rect 8668 13345 8677 13379
rect 8677 13345 8711 13379
rect 8711 13345 8720 13379
rect 8668 13336 8720 13345
rect 9680 13379 9732 13388
rect 9680 13345 9689 13379
rect 9689 13345 9723 13379
rect 9723 13345 9732 13379
rect 9680 13336 9732 13345
rect 9956 13379 10008 13388
rect 9956 13345 9965 13379
rect 9965 13345 9999 13379
rect 9999 13345 10008 13379
rect 9956 13336 10008 13345
rect 10232 13336 10284 13388
rect 19064 13515 19116 13524
rect 19064 13481 19073 13515
rect 19073 13481 19107 13515
rect 19107 13481 19116 13515
rect 19064 13472 19116 13481
rect 23480 13515 23532 13524
rect 23480 13481 23489 13515
rect 23489 13481 23523 13515
rect 23523 13481 23532 13515
rect 23480 13472 23532 13481
rect 13268 13336 13320 13388
rect 15476 13404 15528 13456
rect 14556 13379 14608 13388
rect 14556 13345 14565 13379
rect 14565 13345 14599 13379
rect 14599 13345 14608 13379
rect 14556 13336 14608 13345
rect 14924 13336 14976 13388
rect 16028 13379 16080 13388
rect 16028 13345 16037 13379
rect 16037 13345 16071 13379
rect 16071 13345 16080 13379
rect 16028 13336 16080 13345
rect 17132 13336 17184 13388
rect 17500 13404 17552 13456
rect 17960 13404 18012 13456
rect 19248 13404 19300 13456
rect 21732 13404 21784 13456
rect 17868 13379 17920 13388
rect 17868 13345 17877 13379
rect 17877 13345 17911 13379
rect 17911 13345 17920 13379
rect 17868 13336 17920 13345
rect 18144 13336 18196 13388
rect 18420 13336 18472 13388
rect 18972 13379 19024 13388
rect 18972 13345 18981 13379
rect 18981 13345 19015 13379
rect 19015 13345 19024 13379
rect 18972 13336 19024 13345
rect 19432 13336 19484 13388
rect 19984 13336 20036 13388
rect 21916 13379 21968 13388
rect 21916 13345 21925 13379
rect 21925 13345 21959 13379
rect 21959 13345 21968 13379
rect 21916 13336 21968 13345
rect 22192 13379 22244 13388
rect 22192 13345 22201 13379
rect 22201 13345 22235 13379
rect 22235 13345 22244 13379
rect 22192 13336 22244 13345
rect 23296 13379 23348 13388
rect 17316 13268 17368 13320
rect 18328 13268 18380 13320
rect 21180 13268 21232 13320
rect 21364 13311 21416 13320
rect 21364 13277 21373 13311
rect 21373 13277 21407 13311
rect 21407 13277 21416 13311
rect 21364 13268 21416 13277
rect 23296 13345 23305 13379
rect 23305 13345 23339 13379
rect 23339 13345 23348 13379
rect 23296 13336 23348 13345
rect 24308 13472 24360 13524
rect 28356 13515 28408 13524
rect 28356 13481 28365 13515
rect 28365 13481 28399 13515
rect 28399 13481 28408 13515
rect 28356 13472 28408 13481
rect 24124 13336 24176 13388
rect 25044 13379 25096 13388
rect 25044 13345 25053 13379
rect 25053 13345 25087 13379
rect 25087 13345 25096 13379
rect 25044 13336 25096 13345
rect 25688 13379 25740 13388
rect 23204 13268 23256 13320
rect 6000 13200 6052 13252
rect 11428 13200 11480 13252
rect 4620 13132 4672 13184
rect 7012 13132 7064 13184
rect 9404 13132 9456 13184
rect 14188 13200 14240 13252
rect 14464 13200 14516 13252
rect 14556 13200 14608 13252
rect 13360 13132 13412 13184
rect 13912 13132 13964 13184
rect 15384 13175 15436 13184
rect 15384 13141 15393 13175
rect 15393 13141 15427 13175
rect 15427 13141 15436 13175
rect 15384 13132 15436 13141
rect 16948 13132 17000 13184
rect 17868 13132 17920 13184
rect 19892 13132 19944 13184
rect 20536 13132 20588 13184
rect 23940 13200 23992 13252
rect 25688 13345 25697 13379
rect 25697 13345 25731 13379
rect 25731 13345 25740 13379
rect 25688 13336 25740 13345
rect 27620 13404 27672 13456
rect 27344 13379 27396 13388
rect 27344 13345 27353 13379
rect 27353 13345 27387 13379
rect 27387 13345 27396 13379
rect 27344 13336 27396 13345
rect 27528 13336 27580 13388
rect 28172 13379 28224 13388
rect 27712 13268 27764 13320
rect 28172 13345 28181 13379
rect 28181 13345 28215 13379
rect 28215 13345 28224 13379
rect 28172 13336 28224 13345
rect 28816 13336 28868 13388
rect 30196 13379 30248 13388
rect 29828 13311 29880 13320
rect 29828 13277 29837 13311
rect 29837 13277 29871 13311
rect 29871 13277 29880 13311
rect 29828 13268 29880 13277
rect 30196 13345 30205 13379
rect 30205 13345 30239 13379
rect 30239 13345 30248 13379
rect 30196 13336 30248 13345
rect 30656 13379 30708 13388
rect 30656 13345 30665 13379
rect 30665 13345 30699 13379
rect 30699 13345 30708 13379
rect 30656 13336 30708 13345
rect 30380 13268 30432 13320
rect 27804 13200 27856 13252
rect 31852 13336 31904 13388
rect 32864 13472 32916 13524
rect 34060 13472 34112 13524
rect 34336 13472 34388 13524
rect 34612 13472 34664 13524
rect 35348 13472 35400 13524
rect 33232 13336 33284 13388
rect 31944 13268 31996 13320
rect 34060 13311 34112 13320
rect 34060 13277 34069 13311
rect 34069 13277 34103 13311
rect 34103 13277 34112 13311
rect 34060 13268 34112 13277
rect 34336 13311 34388 13320
rect 34336 13277 34345 13311
rect 34345 13277 34379 13311
rect 34379 13277 34388 13311
rect 34336 13268 34388 13277
rect 32772 13200 32824 13252
rect 33140 13200 33192 13252
rect 27068 13132 27120 13184
rect 28724 13132 28776 13184
rect 31576 13132 31628 13184
rect 33324 13132 33376 13184
rect 33692 13132 33744 13184
rect 37740 13379 37792 13388
rect 37740 13345 37749 13379
rect 37749 13345 37783 13379
rect 37783 13345 37792 13379
rect 37740 13336 37792 13345
rect 36176 13311 36228 13320
rect 36176 13277 36185 13311
rect 36185 13277 36219 13311
rect 36219 13277 36228 13311
rect 36176 13268 36228 13277
rect 36268 13268 36320 13320
rect 37188 13311 37240 13320
rect 37188 13277 37197 13311
rect 37197 13277 37231 13311
rect 37231 13277 37240 13311
rect 37188 13268 37240 13277
rect 35532 13132 35584 13184
rect 4246 13030 4298 13082
rect 4310 13030 4362 13082
rect 4374 13030 4426 13082
rect 4438 13030 4490 13082
rect 34966 13030 35018 13082
rect 35030 13030 35082 13082
rect 35094 13030 35146 13082
rect 35158 13030 35210 13082
rect 6644 12928 6696 12980
rect 7656 12928 7708 12980
rect 9404 12928 9456 12980
rect 11244 12928 11296 12980
rect 11336 12928 11388 12980
rect 22008 12928 22060 12980
rect 22284 12971 22336 12980
rect 22284 12937 22293 12971
rect 22293 12937 22327 12971
rect 22327 12937 22336 12971
rect 22284 12928 22336 12937
rect 22652 12928 22704 12980
rect 28172 12928 28224 12980
rect 36820 12928 36872 12980
rect 4988 12860 5040 12912
rect 6368 12860 6420 12912
rect 1860 12792 1912 12844
rect 3976 12767 4028 12776
rect 3976 12733 3985 12767
rect 3985 12733 4019 12767
rect 4019 12733 4028 12767
rect 3976 12724 4028 12733
rect 4160 12724 4212 12776
rect 4620 12792 4672 12844
rect 13176 12860 13228 12912
rect 16672 12903 16724 12912
rect 5448 12724 5500 12776
rect 10876 12792 10928 12844
rect 11152 12835 11204 12844
rect 11152 12801 11161 12835
rect 11161 12801 11195 12835
rect 11195 12801 11204 12835
rect 11152 12792 11204 12801
rect 6644 12767 6696 12776
rect 6644 12733 6653 12767
rect 6653 12733 6687 12767
rect 6687 12733 6696 12767
rect 6644 12724 6696 12733
rect 7012 12767 7064 12776
rect 7012 12733 7021 12767
rect 7021 12733 7055 12767
rect 7055 12733 7064 12767
rect 7012 12724 7064 12733
rect 8024 12767 8076 12776
rect 4712 12656 4764 12708
rect 6000 12656 6052 12708
rect 6460 12631 6512 12640
rect 6460 12597 6469 12631
rect 6469 12597 6503 12631
rect 6503 12597 6512 12631
rect 6460 12588 6512 12597
rect 6644 12588 6696 12640
rect 6828 12588 6880 12640
rect 8024 12733 8033 12767
rect 8033 12733 8067 12767
rect 8067 12733 8076 12767
rect 8024 12724 8076 12733
rect 8760 12767 8812 12776
rect 8760 12733 8769 12767
rect 8769 12733 8803 12767
rect 8803 12733 8812 12767
rect 8760 12724 8812 12733
rect 9404 12767 9456 12776
rect 9404 12733 9413 12767
rect 9413 12733 9447 12767
rect 9447 12733 9456 12767
rect 9404 12724 9456 12733
rect 9772 12767 9824 12776
rect 9772 12733 9781 12767
rect 9781 12733 9815 12767
rect 9815 12733 9824 12767
rect 9772 12724 9824 12733
rect 8300 12656 8352 12708
rect 9496 12656 9548 12708
rect 11060 12724 11112 12776
rect 11888 12792 11940 12844
rect 13452 12835 13504 12844
rect 11428 12767 11480 12776
rect 11428 12733 11437 12767
rect 11437 12733 11471 12767
rect 11471 12733 11480 12767
rect 11428 12724 11480 12733
rect 13452 12801 13461 12835
rect 13461 12801 13495 12835
rect 13495 12801 13504 12835
rect 13452 12792 13504 12801
rect 16672 12869 16681 12903
rect 16681 12869 16715 12903
rect 16715 12869 16724 12903
rect 16672 12860 16724 12869
rect 16764 12860 16816 12912
rect 13360 12767 13412 12776
rect 11336 12656 11388 12708
rect 13360 12733 13369 12767
rect 13369 12733 13403 12767
rect 13403 12733 13412 12767
rect 13360 12724 13412 12733
rect 14648 12724 14700 12776
rect 15108 12724 15160 12776
rect 15292 12792 15344 12844
rect 16120 12792 16172 12844
rect 19892 12835 19944 12844
rect 15752 12724 15804 12776
rect 16396 12767 16448 12776
rect 16396 12733 16405 12767
rect 16405 12733 16439 12767
rect 16439 12733 16448 12767
rect 16396 12724 16448 12733
rect 13912 12656 13964 12708
rect 15292 12656 15344 12708
rect 17960 12724 18012 12776
rect 18512 12724 18564 12776
rect 19340 12767 19392 12776
rect 19340 12733 19349 12767
rect 19349 12733 19383 12767
rect 19383 12733 19392 12767
rect 19340 12724 19392 12733
rect 19892 12801 19901 12835
rect 19901 12801 19935 12835
rect 19935 12801 19944 12835
rect 19892 12792 19944 12801
rect 19984 12767 20036 12776
rect 19984 12733 19993 12767
rect 19993 12733 20027 12767
rect 20027 12733 20036 12767
rect 19984 12724 20036 12733
rect 20352 12767 20404 12776
rect 20352 12733 20361 12767
rect 20361 12733 20395 12767
rect 20395 12733 20404 12767
rect 20352 12724 20404 12733
rect 20536 12767 20588 12776
rect 20536 12733 20545 12767
rect 20545 12733 20579 12767
rect 20579 12733 20588 12767
rect 20536 12724 20588 12733
rect 20996 12767 21048 12776
rect 20996 12733 21005 12767
rect 21005 12733 21039 12767
rect 21039 12733 21048 12767
rect 20996 12724 21048 12733
rect 23480 12792 23532 12844
rect 23940 12835 23992 12844
rect 23940 12801 23949 12835
rect 23949 12801 23983 12835
rect 23983 12801 23992 12835
rect 23940 12792 23992 12801
rect 23572 12724 23624 12776
rect 19432 12656 19484 12708
rect 20260 12656 20312 12708
rect 23756 12724 23808 12776
rect 24216 12724 24268 12776
rect 24676 12724 24728 12776
rect 24860 12724 24912 12776
rect 25504 12656 25556 12708
rect 27344 12792 27396 12844
rect 26424 12724 26476 12776
rect 10416 12631 10468 12640
rect 10416 12597 10425 12631
rect 10425 12597 10459 12631
rect 10459 12597 10468 12631
rect 10416 12588 10468 12597
rect 15752 12588 15804 12640
rect 18604 12588 18656 12640
rect 20720 12588 20772 12640
rect 22928 12588 22980 12640
rect 25872 12631 25924 12640
rect 25872 12597 25881 12631
rect 25881 12597 25915 12631
rect 25915 12597 25924 12631
rect 25872 12588 25924 12597
rect 27252 12767 27304 12776
rect 27252 12733 27261 12767
rect 27261 12733 27295 12767
rect 27295 12733 27304 12767
rect 27252 12724 27304 12733
rect 27896 12724 27948 12776
rect 28540 12724 28592 12776
rect 29644 12724 29696 12776
rect 30104 12767 30156 12776
rect 30104 12733 30113 12767
rect 30113 12733 30147 12767
rect 30147 12733 30156 12767
rect 30104 12724 30156 12733
rect 31392 12860 31444 12912
rect 34336 12860 34388 12912
rect 32772 12767 32824 12776
rect 27712 12656 27764 12708
rect 29460 12656 29512 12708
rect 32772 12733 32781 12767
rect 32781 12733 32815 12767
rect 32815 12733 32824 12767
rect 32772 12724 32824 12733
rect 35440 12792 35492 12844
rect 36544 12792 36596 12844
rect 34244 12767 34296 12776
rect 32956 12656 33008 12708
rect 29184 12588 29236 12640
rect 29368 12631 29420 12640
rect 29368 12597 29377 12631
rect 29377 12597 29411 12631
rect 29411 12597 29420 12631
rect 29368 12588 29420 12597
rect 29644 12588 29696 12640
rect 29920 12588 29972 12640
rect 34244 12733 34253 12767
rect 34253 12733 34287 12767
rect 34287 12733 34296 12767
rect 34244 12724 34296 12733
rect 35256 12767 35308 12776
rect 35256 12733 35265 12767
rect 35265 12733 35299 12767
rect 35299 12733 35308 12767
rect 35256 12724 35308 12733
rect 36084 12724 36136 12776
rect 36728 12724 36780 12776
rect 37556 12631 37608 12640
rect 37556 12597 37565 12631
rect 37565 12597 37599 12631
rect 37599 12597 37608 12631
rect 37556 12588 37608 12597
rect 19606 12486 19658 12538
rect 19670 12486 19722 12538
rect 19734 12486 19786 12538
rect 19798 12486 19850 12538
rect 1400 12291 1452 12300
rect 1400 12257 1409 12291
rect 1409 12257 1443 12291
rect 1443 12257 1452 12291
rect 1400 12248 1452 12257
rect 4712 12291 4764 12300
rect 4712 12257 4721 12291
rect 4721 12257 4755 12291
rect 4755 12257 4764 12291
rect 4712 12248 4764 12257
rect 5264 12291 5316 12300
rect 5264 12257 5273 12291
rect 5273 12257 5307 12291
rect 5307 12257 5316 12291
rect 5264 12248 5316 12257
rect 7012 12316 7064 12368
rect 6552 12291 6604 12300
rect 6552 12257 6561 12291
rect 6561 12257 6595 12291
rect 6595 12257 6604 12291
rect 6552 12248 6604 12257
rect 6828 12291 6880 12300
rect 6828 12257 6837 12291
rect 6837 12257 6871 12291
rect 6871 12257 6880 12291
rect 6828 12248 6880 12257
rect 1676 12223 1728 12232
rect 1676 12189 1685 12223
rect 1685 12189 1719 12223
rect 1719 12189 1728 12223
rect 1676 12180 1728 12189
rect 4804 12180 4856 12232
rect 2964 12112 3016 12164
rect 7104 12112 7156 12164
rect 9864 12384 9916 12436
rect 10692 12384 10744 12436
rect 10876 12384 10928 12436
rect 15568 12427 15620 12436
rect 9404 12316 9456 12368
rect 9036 12291 9088 12300
rect 9036 12257 9045 12291
rect 9045 12257 9079 12291
rect 9079 12257 9088 12291
rect 9036 12248 9088 12257
rect 9680 12248 9732 12300
rect 11980 12248 12032 12300
rect 15568 12393 15577 12427
rect 15577 12393 15611 12427
rect 15611 12393 15620 12427
rect 15568 12384 15620 12393
rect 13176 12291 13228 12300
rect 13176 12257 13185 12291
rect 13185 12257 13219 12291
rect 13219 12257 13228 12291
rect 13176 12248 13228 12257
rect 14372 12291 14424 12300
rect 8024 12180 8076 12232
rect 10876 12180 10928 12232
rect 13360 12223 13412 12232
rect 13360 12189 13369 12223
rect 13369 12189 13403 12223
rect 13403 12189 13412 12223
rect 13360 12180 13412 12189
rect 14372 12257 14381 12291
rect 14381 12257 14415 12291
rect 14415 12257 14424 12291
rect 14372 12248 14424 12257
rect 16396 12316 16448 12368
rect 16120 12180 16172 12232
rect 2412 12044 2464 12096
rect 8392 12087 8444 12096
rect 8392 12053 8401 12087
rect 8401 12053 8435 12087
rect 8435 12053 8444 12087
rect 8392 12044 8444 12053
rect 14740 12112 14792 12164
rect 17500 12248 17552 12300
rect 18052 12291 18104 12300
rect 18052 12257 18061 12291
rect 18061 12257 18095 12291
rect 18095 12257 18104 12291
rect 18052 12248 18104 12257
rect 18972 12384 19024 12436
rect 19432 12316 19484 12368
rect 18604 12248 18656 12300
rect 18880 12248 18932 12300
rect 19340 12291 19392 12300
rect 19340 12257 19349 12291
rect 19349 12257 19383 12291
rect 19383 12257 19392 12291
rect 19340 12248 19392 12257
rect 19708 12291 19760 12300
rect 19708 12257 19717 12291
rect 19717 12257 19751 12291
rect 19751 12257 19760 12291
rect 19708 12248 19760 12257
rect 21180 12291 21232 12300
rect 21180 12257 21189 12291
rect 21189 12257 21223 12291
rect 21223 12257 21232 12291
rect 21180 12248 21232 12257
rect 24032 12291 24084 12300
rect 18604 12112 18656 12164
rect 11060 12044 11112 12096
rect 11336 12087 11388 12096
rect 11336 12053 11345 12087
rect 11345 12053 11379 12087
rect 11379 12053 11388 12087
rect 11336 12044 11388 12053
rect 11612 12044 11664 12096
rect 12256 12044 12308 12096
rect 13176 12044 13228 12096
rect 14648 12044 14700 12096
rect 17316 12044 17368 12096
rect 19064 12180 19116 12232
rect 20904 12223 20956 12232
rect 20904 12189 20913 12223
rect 20913 12189 20947 12223
rect 20947 12189 20956 12223
rect 20904 12180 20956 12189
rect 23756 12223 23808 12232
rect 23756 12189 23765 12223
rect 23765 12189 23799 12223
rect 23799 12189 23808 12223
rect 23756 12180 23808 12189
rect 24032 12257 24041 12291
rect 24041 12257 24075 12291
rect 24075 12257 24084 12291
rect 24032 12248 24084 12257
rect 27252 12384 27304 12436
rect 27620 12384 27672 12436
rect 27988 12384 28040 12436
rect 29644 12384 29696 12436
rect 30012 12384 30064 12436
rect 28540 12316 28592 12368
rect 29460 12316 29512 12368
rect 27620 12248 27672 12300
rect 27896 12248 27948 12300
rect 28816 12291 28868 12300
rect 28816 12257 28825 12291
rect 28825 12257 28859 12291
rect 28859 12257 28868 12291
rect 28816 12248 28868 12257
rect 29092 12291 29144 12300
rect 29092 12257 29101 12291
rect 29101 12257 29135 12291
rect 29135 12257 29144 12291
rect 29092 12248 29144 12257
rect 32220 12316 32272 12368
rect 32312 12359 32364 12368
rect 32312 12325 32321 12359
rect 32321 12325 32355 12359
rect 32355 12325 32364 12359
rect 32496 12359 32548 12368
rect 32312 12316 32364 12325
rect 32496 12325 32505 12359
rect 32505 12325 32539 12359
rect 32539 12325 32548 12359
rect 32496 12316 32548 12325
rect 30288 12248 30340 12300
rect 31300 12291 31352 12300
rect 31300 12257 31309 12291
rect 31309 12257 31343 12291
rect 31343 12257 31352 12291
rect 32404 12291 32456 12300
rect 31300 12248 31352 12257
rect 32404 12257 32413 12291
rect 32413 12257 32447 12291
rect 32447 12257 32456 12291
rect 32404 12248 32456 12257
rect 33968 12291 34020 12300
rect 33968 12257 33977 12291
rect 33977 12257 34011 12291
rect 34011 12257 34020 12291
rect 33968 12248 34020 12257
rect 34612 12248 34664 12300
rect 37740 12291 37792 12300
rect 37740 12257 37749 12291
rect 37749 12257 37783 12291
rect 37783 12257 37792 12291
rect 37740 12248 37792 12257
rect 25504 12180 25556 12232
rect 27804 12223 27856 12232
rect 27804 12189 27813 12223
rect 27813 12189 27847 12223
rect 27847 12189 27856 12223
rect 27804 12180 27856 12189
rect 22100 12044 22152 12096
rect 23664 12044 23716 12096
rect 25596 12044 25648 12096
rect 27252 12044 27304 12096
rect 28172 12044 28224 12096
rect 31208 12180 31260 12232
rect 31760 12180 31812 12232
rect 32128 12223 32180 12232
rect 32128 12189 32137 12223
rect 32137 12189 32171 12223
rect 32171 12189 32180 12223
rect 32128 12180 32180 12189
rect 32864 12223 32916 12232
rect 32864 12189 32873 12223
rect 32873 12189 32907 12223
rect 32907 12189 32916 12223
rect 32864 12180 32916 12189
rect 33508 12223 33560 12232
rect 33508 12189 33517 12223
rect 33517 12189 33551 12223
rect 33551 12189 33560 12223
rect 33508 12180 33560 12189
rect 35440 12223 35492 12232
rect 28724 12112 28776 12164
rect 30748 12112 30800 12164
rect 34244 12155 34296 12164
rect 34244 12121 34253 12155
rect 34253 12121 34287 12155
rect 34287 12121 34296 12155
rect 34244 12112 34296 12121
rect 30012 12044 30064 12096
rect 30288 12044 30340 12096
rect 35440 12189 35449 12223
rect 35449 12189 35483 12223
rect 35483 12189 35492 12223
rect 35440 12180 35492 12189
rect 37280 12180 37332 12232
rect 35348 12044 35400 12096
rect 4246 11942 4298 11994
rect 4310 11942 4362 11994
rect 4374 11942 4426 11994
rect 4438 11942 4490 11994
rect 34966 11942 35018 11994
rect 35030 11942 35082 11994
rect 35094 11942 35146 11994
rect 35158 11942 35210 11994
rect 1768 11679 1820 11688
rect 1768 11645 1777 11679
rect 1777 11645 1811 11679
rect 1811 11645 1820 11679
rect 1768 11636 1820 11645
rect 4068 11840 4120 11892
rect 4620 11840 4672 11892
rect 5264 11840 5316 11892
rect 6276 11840 6328 11892
rect 5816 11772 5868 11824
rect 8300 11840 8352 11892
rect 10692 11772 10744 11824
rect 10876 11815 10928 11824
rect 10876 11781 10885 11815
rect 10885 11781 10919 11815
rect 10919 11781 10928 11815
rect 10876 11772 10928 11781
rect 14740 11840 14792 11892
rect 2964 11747 3016 11756
rect 2964 11713 2973 11747
rect 2973 11713 3007 11747
rect 3007 11713 3016 11747
rect 2964 11704 3016 11713
rect 6276 11704 6328 11756
rect 6460 11704 6512 11756
rect 8944 11747 8996 11756
rect 4804 11679 4856 11688
rect 1860 11568 1912 11620
rect 4804 11645 4813 11679
rect 4813 11645 4847 11679
rect 4847 11645 4856 11679
rect 4804 11636 4856 11645
rect 5264 11679 5316 11688
rect 5264 11645 5273 11679
rect 5273 11645 5307 11679
rect 5307 11645 5316 11679
rect 5264 11636 5316 11645
rect 5356 11636 5408 11688
rect 7104 11679 7156 11688
rect 7104 11645 7113 11679
rect 7113 11645 7147 11679
rect 7147 11645 7156 11679
rect 7104 11636 7156 11645
rect 7380 11679 7432 11688
rect 7380 11645 7389 11679
rect 7389 11645 7423 11679
rect 7423 11645 7432 11679
rect 7380 11636 7432 11645
rect 8944 11713 8953 11747
rect 8953 11713 8987 11747
rect 8987 11713 8996 11747
rect 8944 11704 8996 11713
rect 9864 11704 9916 11756
rect 11152 11704 11204 11756
rect 8392 11679 8444 11688
rect 8392 11645 8401 11679
rect 8401 11645 8435 11679
rect 8435 11645 8444 11679
rect 8392 11636 8444 11645
rect 8576 11636 8628 11688
rect 9128 11679 9180 11688
rect 9128 11645 9137 11679
rect 9137 11645 9171 11679
rect 9171 11645 9180 11679
rect 9128 11636 9180 11645
rect 9956 11636 10008 11688
rect 10232 11636 10284 11688
rect 10324 11636 10376 11688
rect 12992 11679 13044 11688
rect 12992 11645 13001 11679
rect 13001 11645 13035 11679
rect 13035 11645 13044 11679
rect 12992 11636 13044 11645
rect 13360 11679 13412 11688
rect 13360 11645 13369 11679
rect 13369 11645 13403 11679
rect 13403 11645 13412 11679
rect 13360 11636 13412 11645
rect 15384 11772 15436 11824
rect 15568 11772 15620 11824
rect 17408 11772 17460 11824
rect 14464 11747 14516 11756
rect 14464 11713 14473 11747
rect 14473 11713 14507 11747
rect 14507 11713 14516 11747
rect 14464 11704 14516 11713
rect 17316 11747 17368 11756
rect 17316 11713 17325 11747
rect 17325 11713 17359 11747
rect 17359 11713 17368 11747
rect 17316 11704 17368 11713
rect 14648 11679 14700 11688
rect 14648 11645 14657 11679
rect 14657 11645 14691 11679
rect 14691 11645 14700 11679
rect 14648 11636 14700 11645
rect 15384 11636 15436 11688
rect 15476 11636 15528 11688
rect 15936 11636 15988 11688
rect 16396 11679 16448 11688
rect 16396 11645 16405 11679
rect 16405 11645 16439 11679
rect 16439 11645 16448 11679
rect 16396 11636 16448 11645
rect 18052 11679 18104 11688
rect 1676 11500 1728 11552
rect 4896 11500 4948 11552
rect 8116 11500 8168 11552
rect 10140 11500 10192 11552
rect 12900 11568 12952 11620
rect 18052 11645 18061 11679
rect 18061 11645 18095 11679
rect 18095 11645 18104 11679
rect 18052 11636 18104 11645
rect 18604 11840 18656 11892
rect 19064 11840 19116 11892
rect 19708 11840 19760 11892
rect 24216 11840 24268 11892
rect 27712 11840 27764 11892
rect 27988 11840 28040 11892
rect 29828 11840 29880 11892
rect 19892 11704 19944 11756
rect 21272 11704 21324 11756
rect 18788 11679 18840 11688
rect 18788 11645 18797 11679
rect 18797 11645 18831 11679
rect 18831 11645 18840 11679
rect 18788 11636 18840 11645
rect 20260 11636 20312 11688
rect 20904 11636 20956 11688
rect 21456 11636 21508 11688
rect 22100 11679 22152 11688
rect 22100 11645 22109 11679
rect 22109 11645 22143 11679
rect 22143 11645 22152 11679
rect 22100 11636 22152 11645
rect 22468 11636 22520 11688
rect 25504 11772 25556 11824
rect 24676 11704 24728 11756
rect 26148 11704 26200 11756
rect 26424 11636 26476 11688
rect 26976 11636 27028 11688
rect 27252 11636 27304 11688
rect 27620 11704 27672 11756
rect 27712 11679 27764 11688
rect 27712 11645 27721 11679
rect 27721 11645 27755 11679
rect 27755 11645 27764 11679
rect 27712 11636 27764 11645
rect 30196 11772 30248 11824
rect 31300 11840 31352 11892
rect 37464 11840 37516 11892
rect 37832 11883 37884 11892
rect 37832 11849 37841 11883
rect 37841 11849 37875 11883
rect 37875 11849 37884 11883
rect 37832 11840 37884 11849
rect 31944 11772 31996 11824
rect 33968 11772 34020 11824
rect 29184 11636 29236 11688
rect 32220 11704 32272 11756
rect 33784 11747 33836 11756
rect 33784 11713 33793 11747
rect 33793 11713 33827 11747
rect 33827 11713 33836 11747
rect 33784 11704 33836 11713
rect 34520 11704 34572 11756
rect 34796 11704 34848 11756
rect 30196 11679 30248 11688
rect 22560 11611 22612 11620
rect 14372 11500 14424 11552
rect 14648 11500 14700 11552
rect 19432 11500 19484 11552
rect 22560 11577 22569 11611
rect 22569 11577 22603 11611
rect 22603 11577 22612 11611
rect 22560 11568 22612 11577
rect 20076 11500 20128 11552
rect 22284 11500 22336 11552
rect 25320 11568 25372 11620
rect 25596 11611 25648 11620
rect 25596 11577 25605 11611
rect 25605 11577 25639 11611
rect 25639 11577 25648 11611
rect 25596 11568 25648 11577
rect 25964 11611 26016 11620
rect 25964 11577 25973 11611
rect 25973 11577 26007 11611
rect 26007 11577 26016 11611
rect 25964 11568 26016 11577
rect 29736 11568 29788 11620
rect 30196 11645 30205 11679
rect 30205 11645 30239 11679
rect 30239 11645 30248 11679
rect 30196 11636 30248 11645
rect 30472 11636 30524 11688
rect 31208 11679 31260 11688
rect 31208 11645 31217 11679
rect 31217 11645 31251 11679
rect 31251 11645 31260 11679
rect 31208 11636 31260 11645
rect 31576 11679 31628 11688
rect 31576 11645 31585 11679
rect 31585 11645 31619 11679
rect 31619 11645 31628 11679
rect 31576 11636 31628 11645
rect 31944 11636 31996 11688
rect 31668 11568 31720 11620
rect 32496 11636 32548 11688
rect 33324 11636 33376 11688
rect 34060 11636 34112 11688
rect 35808 11636 35860 11688
rect 36452 11679 36504 11688
rect 36452 11645 36461 11679
rect 36461 11645 36495 11679
rect 36495 11645 36504 11679
rect 36452 11636 36504 11645
rect 36728 11679 36780 11688
rect 36728 11645 36737 11679
rect 36737 11645 36771 11679
rect 36771 11645 36780 11679
rect 36728 11636 36780 11645
rect 32680 11568 32732 11620
rect 25412 11543 25464 11552
rect 25412 11509 25421 11543
rect 25421 11509 25455 11543
rect 25455 11509 25464 11543
rect 25412 11500 25464 11509
rect 25504 11543 25556 11552
rect 25504 11509 25513 11543
rect 25513 11509 25547 11543
rect 25547 11509 25556 11543
rect 25504 11500 25556 11509
rect 29000 11500 29052 11552
rect 29460 11500 29512 11552
rect 29828 11500 29880 11552
rect 33048 11500 33100 11552
rect 19606 11398 19658 11450
rect 19670 11398 19722 11450
rect 19734 11398 19786 11450
rect 19798 11398 19850 11450
rect 5080 11296 5132 11348
rect 7104 11296 7156 11348
rect 7932 11296 7984 11348
rect 8116 11296 8168 11348
rect 2412 11203 2464 11212
rect 2412 11169 2421 11203
rect 2421 11169 2455 11203
rect 2455 11169 2464 11203
rect 2412 11160 2464 11169
rect 4620 11203 4672 11212
rect 4620 11169 4629 11203
rect 4629 11169 4663 11203
rect 4663 11169 4672 11203
rect 4620 11160 4672 11169
rect 6460 11228 6512 11280
rect 5816 11203 5868 11212
rect 5816 11169 5825 11203
rect 5825 11169 5859 11203
rect 5859 11169 5868 11203
rect 5816 11160 5868 11169
rect 6276 11160 6328 11212
rect 6920 11160 6972 11212
rect 7564 11160 7616 11212
rect 10140 11228 10192 11280
rect 8944 11203 8996 11212
rect 2136 11092 2188 11144
rect 2872 11135 2924 11144
rect 2872 11101 2881 11135
rect 2881 11101 2915 11135
rect 2915 11101 2924 11135
rect 2872 11092 2924 11101
rect 6184 11092 6236 11144
rect 8944 11169 8953 11203
rect 8953 11169 8987 11203
rect 8987 11169 8996 11203
rect 8944 11160 8996 11169
rect 10600 11203 10652 11212
rect 10600 11169 10609 11203
rect 10609 11169 10643 11203
rect 10643 11169 10652 11203
rect 10600 11160 10652 11169
rect 10692 11135 10744 11144
rect 10692 11101 10701 11135
rect 10701 11101 10735 11135
rect 10735 11101 10744 11135
rect 10692 11092 10744 11101
rect 10968 11203 11020 11212
rect 10968 11169 10977 11203
rect 10977 11169 11011 11203
rect 11011 11169 11020 11203
rect 10968 11160 11020 11169
rect 11520 11296 11572 11348
rect 14648 11296 14700 11348
rect 16212 11296 16264 11348
rect 18236 11296 18288 11348
rect 12992 11228 13044 11280
rect 12808 11160 12860 11212
rect 13084 11203 13136 11212
rect 13084 11169 13093 11203
rect 13093 11169 13127 11203
rect 13127 11169 13136 11203
rect 13084 11160 13136 11169
rect 14740 11228 14792 11280
rect 17960 11228 18012 11280
rect 14372 11203 14424 11212
rect 14372 11169 14381 11203
rect 14381 11169 14415 11203
rect 14415 11169 14424 11203
rect 14372 11160 14424 11169
rect 14464 11160 14516 11212
rect 15568 11203 15620 11212
rect 15568 11169 15577 11203
rect 15577 11169 15611 11203
rect 15611 11169 15620 11203
rect 16028 11203 16080 11212
rect 15568 11160 15620 11169
rect 16028 11169 16037 11203
rect 16037 11169 16071 11203
rect 16071 11169 16080 11203
rect 16028 11160 16080 11169
rect 15844 11092 15896 11144
rect 18052 11160 18104 11212
rect 18420 11203 18472 11212
rect 18420 11169 18429 11203
rect 18429 11169 18463 11203
rect 18463 11169 18472 11203
rect 18420 11160 18472 11169
rect 18604 11160 18656 11212
rect 19156 11160 19208 11212
rect 19432 11203 19484 11212
rect 19432 11169 19441 11203
rect 19441 11169 19475 11203
rect 19475 11169 19484 11203
rect 19432 11160 19484 11169
rect 22376 11296 22428 11348
rect 20076 11228 20128 11280
rect 24216 11296 24268 11348
rect 16672 11092 16724 11144
rect 4620 11024 4672 11076
rect 12900 11024 12952 11076
rect 9864 10956 9916 11008
rect 10508 10956 10560 11008
rect 15292 11024 15344 11076
rect 18972 11092 19024 11144
rect 22284 11160 22336 11212
rect 22468 11203 22520 11212
rect 22468 11169 22477 11203
rect 22477 11169 22511 11203
rect 22511 11169 22520 11203
rect 22468 11160 22520 11169
rect 24860 11296 24912 11348
rect 27620 11296 27672 11348
rect 27712 11296 27764 11348
rect 30472 11296 30524 11348
rect 30748 11296 30800 11348
rect 37004 11339 37056 11348
rect 25964 11228 26016 11280
rect 25596 11160 25648 11212
rect 27160 11160 27212 11212
rect 28632 11203 28684 11212
rect 28632 11169 28641 11203
rect 28641 11169 28675 11203
rect 28675 11169 28684 11203
rect 28632 11160 28684 11169
rect 29184 11203 29236 11212
rect 29184 11169 29193 11203
rect 29193 11169 29227 11203
rect 29227 11169 29236 11203
rect 29184 11160 29236 11169
rect 29092 11135 29144 11144
rect 29092 11101 29101 11135
rect 29101 11101 29135 11135
rect 29135 11101 29144 11135
rect 29092 11092 29144 11101
rect 18328 11024 18380 11076
rect 20720 11024 20772 11076
rect 21456 11024 21508 11076
rect 26516 11024 26568 11076
rect 13820 10956 13872 11008
rect 21916 10999 21968 11008
rect 21916 10965 21925 10999
rect 21925 10965 21959 10999
rect 21959 10965 21968 10999
rect 21916 10956 21968 10965
rect 26148 10956 26200 11008
rect 28080 11024 28132 11076
rect 29828 11160 29880 11212
rect 30564 11135 30616 11144
rect 30564 11101 30573 11135
rect 30573 11101 30607 11135
rect 30607 11101 30616 11135
rect 30564 11092 30616 11101
rect 31300 11160 31352 11212
rect 31944 11228 31996 11280
rect 33140 11228 33192 11280
rect 31760 11160 31812 11212
rect 32680 11203 32732 11212
rect 32680 11169 32689 11203
rect 32689 11169 32723 11203
rect 32723 11169 32732 11203
rect 32680 11160 32732 11169
rect 33048 11203 33100 11212
rect 33048 11169 33057 11203
rect 33057 11169 33091 11203
rect 33091 11169 33100 11203
rect 33048 11160 33100 11169
rect 34060 11203 34112 11212
rect 34060 11169 34069 11203
rect 34069 11169 34103 11203
rect 34103 11169 34112 11203
rect 34060 11160 34112 11169
rect 37004 11305 37013 11339
rect 37013 11305 37047 11339
rect 37047 11305 37056 11339
rect 37004 11296 37056 11305
rect 31760 11024 31812 11076
rect 33600 11092 33652 11144
rect 34244 11092 34296 11144
rect 35348 11092 35400 11144
rect 35716 11135 35768 11144
rect 35716 11101 35725 11135
rect 35725 11101 35759 11135
rect 35759 11101 35768 11135
rect 35716 11092 35768 11101
rect 27528 10956 27580 11008
rect 33876 10956 33928 11008
rect 35900 10956 35952 11008
rect 4246 10854 4298 10906
rect 4310 10854 4362 10906
rect 4374 10854 4426 10906
rect 4438 10854 4490 10906
rect 34966 10854 35018 10906
rect 35030 10854 35082 10906
rect 35094 10854 35146 10906
rect 35158 10854 35210 10906
rect 8668 10752 8720 10804
rect 15844 10795 15896 10804
rect 10324 10684 10376 10736
rect 13176 10684 13228 10736
rect 15844 10761 15853 10795
rect 15853 10761 15887 10795
rect 15887 10761 15896 10795
rect 15844 10752 15896 10761
rect 16856 10752 16908 10804
rect 22560 10752 22612 10804
rect 2228 10548 2280 10600
rect 2964 10548 3016 10600
rect 3148 10591 3200 10600
rect 3148 10557 3157 10591
rect 3157 10557 3191 10591
rect 3191 10557 3200 10591
rect 4620 10616 4672 10668
rect 6184 10616 6236 10668
rect 6736 10616 6788 10668
rect 14096 10616 14148 10668
rect 16580 10684 16632 10736
rect 17224 10684 17276 10736
rect 22100 10684 22152 10736
rect 22836 10684 22888 10736
rect 23664 10684 23716 10736
rect 23940 10684 23992 10736
rect 27528 10684 27580 10736
rect 27712 10684 27764 10736
rect 3148 10548 3200 10557
rect 4804 10591 4856 10600
rect 3608 10523 3660 10532
rect 3608 10489 3617 10523
rect 3617 10489 3651 10523
rect 3651 10489 3660 10523
rect 3608 10480 3660 10489
rect 4804 10557 4813 10591
rect 4813 10557 4847 10591
rect 4847 10557 4856 10591
rect 4804 10548 4856 10557
rect 5264 10480 5316 10532
rect 5816 10591 5868 10600
rect 5816 10557 5825 10591
rect 5825 10557 5859 10591
rect 5859 10557 5868 10591
rect 5816 10548 5868 10557
rect 6644 10548 6696 10600
rect 8300 10591 8352 10600
rect 7288 10480 7340 10532
rect 8300 10557 8309 10591
rect 8309 10557 8343 10591
rect 8343 10557 8352 10591
rect 8300 10548 8352 10557
rect 9680 10548 9732 10600
rect 10968 10591 11020 10600
rect 10968 10557 10977 10591
rect 10977 10557 11011 10591
rect 11011 10557 11020 10591
rect 10968 10548 11020 10557
rect 11336 10591 11388 10600
rect 8392 10480 8444 10532
rect 10232 10480 10284 10532
rect 10692 10480 10744 10532
rect 11336 10557 11345 10591
rect 11345 10557 11379 10591
rect 11379 10557 11388 10591
rect 11336 10548 11388 10557
rect 11520 10591 11572 10600
rect 11520 10557 11529 10591
rect 11529 10557 11563 10591
rect 11563 10557 11572 10591
rect 11520 10548 11572 10557
rect 11796 10548 11848 10600
rect 12992 10591 13044 10600
rect 12992 10557 13001 10591
rect 13001 10557 13035 10591
rect 13035 10557 13044 10591
rect 12992 10548 13044 10557
rect 13268 10591 13320 10600
rect 13268 10557 13277 10591
rect 13277 10557 13311 10591
rect 13311 10557 13320 10591
rect 13268 10548 13320 10557
rect 14004 10480 14056 10532
rect 2320 10455 2372 10464
rect 2320 10421 2329 10455
rect 2329 10421 2363 10455
rect 2363 10421 2372 10455
rect 2320 10412 2372 10421
rect 11796 10412 11848 10464
rect 15016 10591 15068 10600
rect 15016 10557 15025 10591
rect 15025 10557 15059 10591
rect 15059 10557 15068 10591
rect 15016 10548 15068 10557
rect 15568 10548 15620 10600
rect 17408 10591 17460 10600
rect 17408 10557 17417 10591
rect 17417 10557 17451 10591
rect 17451 10557 17460 10591
rect 17408 10548 17460 10557
rect 18328 10591 18380 10600
rect 18328 10557 18337 10591
rect 18337 10557 18371 10591
rect 18371 10557 18380 10591
rect 18328 10548 18380 10557
rect 18604 10591 18656 10600
rect 18604 10557 18613 10591
rect 18613 10557 18647 10591
rect 18647 10557 18656 10591
rect 18604 10548 18656 10557
rect 19432 10591 19484 10600
rect 19432 10557 19441 10591
rect 19441 10557 19475 10591
rect 19475 10557 19484 10591
rect 19432 10548 19484 10557
rect 15476 10412 15528 10464
rect 19340 10412 19392 10464
rect 21824 10548 21876 10600
rect 22008 10591 22060 10600
rect 22008 10557 22017 10591
rect 22017 10557 22051 10591
rect 22051 10557 22060 10591
rect 22008 10548 22060 10557
rect 22376 10591 22428 10600
rect 22376 10557 22385 10591
rect 22385 10557 22419 10591
rect 22419 10557 22428 10591
rect 22376 10548 22428 10557
rect 22468 10591 22520 10600
rect 22468 10557 22477 10591
rect 22477 10557 22511 10591
rect 22511 10557 22520 10591
rect 27804 10616 27856 10668
rect 27988 10659 28040 10668
rect 27988 10625 27997 10659
rect 27997 10625 28031 10659
rect 28031 10625 28040 10659
rect 27988 10616 28040 10625
rect 28540 10684 28592 10736
rect 28908 10684 28960 10736
rect 30104 10684 30156 10736
rect 32220 10684 32272 10736
rect 23664 10591 23716 10600
rect 22468 10548 22520 10557
rect 23664 10557 23673 10591
rect 23673 10557 23707 10591
rect 23707 10557 23716 10591
rect 23664 10548 23716 10557
rect 24952 10591 25004 10600
rect 24952 10557 24961 10591
rect 24961 10557 24995 10591
rect 24995 10557 25004 10591
rect 24952 10548 25004 10557
rect 25412 10548 25464 10600
rect 26148 10548 26200 10600
rect 26516 10548 26568 10600
rect 28172 10591 28224 10600
rect 28172 10557 28181 10591
rect 28181 10557 28215 10591
rect 28215 10557 28224 10591
rect 28172 10548 28224 10557
rect 29736 10616 29788 10668
rect 31668 10616 31720 10668
rect 29828 10591 29880 10600
rect 29828 10557 29837 10591
rect 29837 10557 29871 10591
rect 29871 10557 29880 10591
rect 29828 10548 29880 10557
rect 30012 10591 30064 10600
rect 30012 10557 30021 10591
rect 30021 10557 30055 10591
rect 30055 10557 30064 10591
rect 30012 10548 30064 10557
rect 30196 10591 30248 10600
rect 30196 10557 30205 10591
rect 30205 10557 30239 10591
rect 30239 10557 30248 10591
rect 30196 10548 30248 10557
rect 32864 10616 32916 10668
rect 22836 10480 22888 10532
rect 23296 10480 23348 10532
rect 26240 10523 26292 10532
rect 26240 10489 26249 10523
rect 26249 10489 26283 10523
rect 26283 10489 26292 10523
rect 26240 10480 26292 10489
rect 27068 10523 27120 10532
rect 27068 10489 27077 10523
rect 27077 10489 27111 10523
rect 27111 10489 27120 10523
rect 27068 10480 27120 10489
rect 27160 10523 27212 10532
rect 27160 10489 27169 10523
rect 27169 10489 27203 10523
rect 27203 10489 27212 10523
rect 27528 10523 27580 10532
rect 27160 10480 27212 10489
rect 27528 10489 27537 10523
rect 27537 10489 27571 10523
rect 27571 10489 27580 10523
rect 27528 10480 27580 10489
rect 27988 10480 28040 10532
rect 21640 10412 21692 10464
rect 21732 10412 21784 10464
rect 26332 10412 26384 10464
rect 27620 10412 27672 10464
rect 28448 10412 28500 10464
rect 28816 10480 28868 10532
rect 31116 10480 31168 10532
rect 32588 10591 32640 10600
rect 32588 10557 32597 10591
rect 32597 10557 32631 10591
rect 32631 10557 32640 10591
rect 32588 10548 32640 10557
rect 33048 10548 33100 10600
rect 33600 10591 33652 10600
rect 33600 10557 33609 10591
rect 33609 10557 33643 10591
rect 33643 10557 33652 10591
rect 33600 10548 33652 10557
rect 33968 10548 34020 10600
rect 34152 10548 34204 10600
rect 35900 10659 35952 10668
rect 35900 10625 35909 10659
rect 35909 10625 35943 10659
rect 35943 10625 35952 10659
rect 36452 10659 36504 10668
rect 35900 10616 35952 10625
rect 36452 10625 36461 10659
rect 36461 10625 36495 10659
rect 36495 10625 36504 10659
rect 36452 10616 36504 10625
rect 36084 10480 36136 10532
rect 38108 10523 38160 10532
rect 38108 10489 38117 10523
rect 38117 10489 38151 10523
rect 38151 10489 38160 10523
rect 38108 10480 38160 10489
rect 32128 10412 32180 10464
rect 34704 10412 34756 10464
rect 37188 10412 37240 10464
rect 19606 10310 19658 10362
rect 19670 10310 19722 10362
rect 19734 10310 19786 10362
rect 19798 10310 19850 10362
rect 3148 10251 3200 10260
rect 3148 10217 3157 10251
rect 3157 10217 3191 10251
rect 3191 10217 3200 10251
rect 3148 10208 3200 10217
rect 5816 10208 5868 10260
rect 8300 10208 8352 10260
rect 8576 10208 8628 10260
rect 10324 10208 10376 10260
rect 21732 10208 21784 10260
rect 2964 10072 3016 10124
rect 4620 10072 4672 10124
rect 5080 10072 5132 10124
rect 12624 10140 12676 10192
rect 16672 10183 16724 10192
rect 1400 9868 1452 9920
rect 3608 10004 3660 10056
rect 5816 10047 5868 10056
rect 5816 10013 5825 10047
rect 5825 10013 5859 10047
rect 5859 10013 5868 10047
rect 5816 10004 5868 10013
rect 8944 10072 8996 10124
rect 9496 10115 9548 10124
rect 9496 10081 9505 10115
rect 9505 10081 9539 10115
rect 9539 10081 9548 10115
rect 9496 10072 9548 10081
rect 9864 10072 9916 10124
rect 10140 10115 10192 10124
rect 10140 10081 10149 10115
rect 10149 10081 10183 10115
rect 10183 10081 10192 10115
rect 10140 10072 10192 10081
rect 10232 10072 10284 10124
rect 10508 10115 10560 10124
rect 10508 10081 10517 10115
rect 10517 10081 10551 10115
rect 10551 10081 10560 10115
rect 10508 10072 10560 10081
rect 11888 10072 11940 10124
rect 12532 10115 12584 10124
rect 12532 10081 12541 10115
rect 12541 10081 12575 10115
rect 12575 10081 12584 10115
rect 12532 10072 12584 10081
rect 16672 10149 16681 10183
rect 16681 10149 16715 10183
rect 16715 10149 16724 10183
rect 16672 10140 16724 10149
rect 13820 10115 13872 10124
rect 8576 10004 8628 10056
rect 6736 9936 6788 9988
rect 11336 10004 11388 10056
rect 12072 10047 12124 10056
rect 12072 10013 12081 10047
rect 12081 10013 12115 10047
rect 12115 10013 12124 10047
rect 12072 10004 12124 10013
rect 12256 10004 12308 10056
rect 13820 10081 13829 10115
rect 13829 10081 13863 10115
rect 13863 10081 13872 10115
rect 13820 10072 13872 10081
rect 14004 10115 14056 10124
rect 14004 10081 14013 10115
rect 14013 10081 14047 10115
rect 14047 10081 14056 10115
rect 14004 10072 14056 10081
rect 15752 10115 15804 10124
rect 15752 10081 15761 10115
rect 15761 10081 15795 10115
rect 15795 10081 15804 10115
rect 15752 10072 15804 10081
rect 16212 10115 16264 10124
rect 16212 10081 16221 10115
rect 16221 10081 16255 10115
rect 16255 10081 16264 10115
rect 16212 10072 16264 10081
rect 18236 10140 18288 10192
rect 18604 10140 18656 10192
rect 19064 10140 19116 10192
rect 17408 10115 17460 10124
rect 17408 10081 17417 10115
rect 17417 10081 17451 10115
rect 17451 10081 17460 10115
rect 17408 10072 17460 10081
rect 17592 10072 17644 10124
rect 19156 10072 19208 10124
rect 19340 10115 19392 10124
rect 19340 10081 19349 10115
rect 19349 10081 19383 10115
rect 19383 10081 19392 10115
rect 19340 10072 19392 10081
rect 19432 10115 19484 10124
rect 19432 10081 19441 10115
rect 19441 10081 19475 10115
rect 19475 10081 19484 10115
rect 19432 10072 19484 10081
rect 20076 10072 20128 10124
rect 20628 10072 20680 10124
rect 20812 10072 20864 10124
rect 21272 10115 21324 10124
rect 21272 10081 21281 10115
rect 21281 10081 21315 10115
rect 21315 10081 21324 10115
rect 21272 10072 21324 10081
rect 14096 10004 14148 10056
rect 16028 9936 16080 9988
rect 9312 9911 9364 9920
rect 9312 9877 9321 9911
rect 9321 9877 9355 9911
rect 9355 9877 9364 9911
rect 9312 9868 9364 9877
rect 11704 9868 11756 9920
rect 19064 10047 19116 10056
rect 19064 10013 19073 10047
rect 19073 10013 19107 10047
rect 19107 10013 19116 10047
rect 19064 10004 19116 10013
rect 19248 10004 19300 10056
rect 20536 10004 20588 10056
rect 22284 10072 22336 10124
rect 22560 10072 22612 10124
rect 21732 10047 21784 10056
rect 21732 10013 21741 10047
rect 21741 10013 21775 10047
rect 21775 10013 21784 10047
rect 21732 10004 21784 10013
rect 20260 9936 20312 9988
rect 21088 9936 21140 9988
rect 22008 9936 22060 9988
rect 35808 10208 35860 10260
rect 36636 10208 36688 10260
rect 27068 10140 27120 10192
rect 23296 10115 23348 10124
rect 23296 10081 23305 10115
rect 23305 10081 23339 10115
rect 23339 10081 23348 10115
rect 23296 10072 23348 10081
rect 25504 10115 25556 10124
rect 25504 10081 25513 10115
rect 25513 10081 25547 10115
rect 25547 10081 25556 10115
rect 25504 10072 25556 10081
rect 25688 10115 25740 10124
rect 25688 10081 25697 10115
rect 25697 10081 25731 10115
rect 25731 10081 25740 10115
rect 25688 10072 25740 10081
rect 26148 10072 26200 10124
rect 26976 10072 27028 10124
rect 27896 10115 27948 10124
rect 23204 10004 23256 10056
rect 27344 10004 27396 10056
rect 27896 10081 27905 10115
rect 27905 10081 27939 10115
rect 27939 10081 27948 10115
rect 27896 10072 27948 10081
rect 27988 10072 28040 10124
rect 28356 10115 28408 10124
rect 28356 10081 28365 10115
rect 28365 10081 28399 10115
rect 28399 10081 28408 10115
rect 28356 10072 28408 10081
rect 27804 10047 27856 10056
rect 27804 10013 27813 10047
rect 27813 10013 27847 10047
rect 27847 10013 27856 10047
rect 27804 10004 27856 10013
rect 28816 10140 28868 10192
rect 29000 10072 29052 10124
rect 29184 10115 29236 10124
rect 29184 10081 29193 10115
rect 29193 10081 29227 10115
rect 29227 10081 29236 10115
rect 29184 10072 29236 10081
rect 29460 10072 29512 10124
rect 31208 10140 31260 10192
rect 31944 10140 31996 10192
rect 34152 10140 34204 10192
rect 31116 10115 31168 10124
rect 31116 10081 31125 10115
rect 31125 10081 31159 10115
rect 31159 10081 31168 10115
rect 31116 10072 31168 10081
rect 32956 10115 33008 10124
rect 32956 10081 32965 10115
rect 32965 10081 32999 10115
rect 32999 10081 33008 10115
rect 32956 10072 33008 10081
rect 33416 10115 33468 10124
rect 33416 10081 33425 10115
rect 33425 10081 33459 10115
rect 33459 10081 33468 10115
rect 33416 10072 33468 10081
rect 33784 10072 33836 10124
rect 34704 10115 34756 10124
rect 34704 10081 34713 10115
rect 34713 10081 34747 10115
rect 34747 10081 34756 10115
rect 34704 10072 34756 10081
rect 37004 10072 37056 10124
rect 37740 10115 37792 10124
rect 37740 10081 37749 10115
rect 37749 10081 37783 10115
rect 37783 10081 37792 10115
rect 37740 10072 37792 10081
rect 30380 10004 30432 10056
rect 30840 10004 30892 10056
rect 31944 10004 31996 10056
rect 32312 10004 32364 10056
rect 33048 10004 33100 10056
rect 27988 9936 28040 9988
rect 19248 9868 19300 9920
rect 22376 9868 22428 9920
rect 22744 9868 22796 9920
rect 23296 9868 23348 9920
rect 24952 9868 25004 9920
rect 27160 9868 27212 9920
rect 29736 9936 29788 9988
rect 30012 9936 30064 9988
rect 32864 9936 32916 9988
rect 34796 10004 34848 10056
rect 35348 10004 35400 10056
rect 35808 10004 35860 10056
rect 28448 9868 28500 9920
rect 29000 9868 29052 9920
rect 29460 9868 29512 9920
rect 30380 9868 30432 9920
rect 31024 9868 31076 9920
rect 31392 9868 31444 9920
rect 32588 9868 32640 9920
rect 33048 9868 33100 9920
rect 4246 9766 4298 9818
rect 4310 9766 4362 9818
rect 4374 9766 4426 9818
rect 4438 9766 4490 9818
rect 34966 9766 35018 9818
rect 35030 9766 35082 9818
rect 35094 9766 35146 9818
rect 35158 9766 35210 9818
rect 2780 9707 2832 9716
rect 2780 9673 2789 9707
rect 2789 9673 2823 9707
rect 2823 9673 2832 9707
rect 2780 9664 2832 9673
rect 7288 9664 7340 9716
rect 14096 9664 14148 9716
rect 15752 9707 15804 9716
rect 15752 9673 15761 9707
rect 15761 9673 15795 9707
rect 15795 9673 15804 9707
rect 15752 9664 15804 9673
rect 20812 9664 20864 9716
rect 7012 9596 7064 9648
rect 1400 9571 1452 9580
rect 1400 9537 1409 9571
rect 1409 9537 1443 9571
rect 1443 9537 1452 9571
rect 1400 9528 1452 9537
rect 6552 9528 6604 9580
rect 1768 9460 1820 9512
rect 2320 9460 2372 9512
rect 4896 9503 4948 9512
rect 4896 9469 4905 9503
rect 4905 9469 4939 9503
rect 4939 9469 4948 9503
rect 4896 9460 4948 9469
rect 6644 9460 6696 9512
rect 7932 9596 7984 9648
rect 11152 9639 11204 9648
rect 9036 9571 9088 9580
rect 9036 9537 9045 9571
rect 9045 9537 9079 9571
rect 9079 9537 9088 9571
rect 9036 9528 9088 9537
rect 7840 9460 7892 9512
rect 8852 9503 8904 9512
rect 8852 9469 8861 9503
rect 8861 9469 8895 9503
rect 8895 9469 8904 9503
rect 8852 9460 8904 9469
rect 11152 9605 11161 9639
rect 11161 9605 11195 9639
rect 11195 9605 11204 9639
rect 11152 9596 11204 9605
rect 10508 9528 10560 9580
rect 12716 9596 12768 9648
rect 13268 9596 13320 9648
rect 16580 9596 16632 9648
rect 12256 9528 12308 9580
rect 9956 9503 10008 9512
rect 9956 9469 9965 9503
rect 9965 9469 9999 9503
rect 9999 9469 10008 9503
rect 9956 9460 10008 9469
rect 11336 9503 11388 9512
rect 11336 9469 11345 9503
rect 11345 9469 11379 9503
rect 11379 9469 11388 9503
rect 11336 9460 11388 9469
rect 11520 9503 11572 9512
rect 11520 9469 11529 9503
rect 11529 9469 11563 9503
rect 11563 9469 11572 9503
rect 11520 9460 11572 9469
rect 11704 9503 11756 9512
rect 11704 9469 11713 9503
rect 11713 9469 11747 9503
rect 11747 9469 11756 9503
rect 11704 9460 11756 9469
rect 12164 9460 12216 9512
rect 14096 9528 14148 9580
rect 17500 9571 17552 9580
rect 3608 9367 3660 9376
rect 3608 9333 3617 9367
rect 3617 9333 3651 9367
rect 3651 9333 3660 9367
rect 3608 9324 3660 9333
rect 5540 9324 5592 9376
rect 5816 9367 5868 9376
rect 5816 9333 5825 9367
rect 5825 9333 5859 9367
rect 5859 9333 5868 9367
rect 5816 9324 5868 9333
rect 7104 9367 7156 9376
rect 7104 9333 7113 9367
rect 7113 9333 7147 9367
rect 7147 9333 7156 9367
rect 7104 9324 7156 9333
rect 12072 9392 12124 9444
rect 14464 9460 14516 9512
rect 9496 9324 9548 9376
rect 10416 9324 10468 9376
rect 12624 9324 12676 9376
rect 14004 9324 14056 9376
rect 17040 9324 17092 9376
rect 17500 9537 17509 9571
rect 17509 9537 17543 9571
rect 17543 9537 17552 9571
rect 17500 9528 17552 9537
rect 20168 9596 20220 9648
rect 21916 9596 21968 9648
rect 23940 9664 23992 9716
rect 25504 9664 25556 9716
rect 32404 9664 32456 9716
rect 19892 9528 19944 9580
rect 22100 9528 22152 9580
rect 18604 9460 18656 9512
rect 18972 9460 19024 9512
rect 19984 9503 20036 9512
rect 19432 9392 19484 9444
rect 17960 9324 18012 9376
rect 18328 9324 18380 9376
rect 18880 9367 18932 9376
rect 18880 9333 18889 9367
rect 18889 9333 18923 9367
rect 18923 9333 18932 9367
rect 18880 9324 18932 9333
rect 19984 9469 19993 9503
rect 19993 9469 20027 9503
rect 20027 9469 20036 9503
rect 19984 9460 20036 9469
rect 20168 9460 20220 9512
rect 20904 9503 20956 9512
rect 20904 9469 20913 9503
rect 20913 9469 20947 9503
rect 20947 9469 20956 9503
rect 20904 9460 20956 9469
rect 21272 9460 21324 9512
rect 21916 9460 21968 9512
rect 22008 9460 22060 9512
rect 23204 9528 23256 9580
rect 22928 9460 22980 9512
rect 25688 9596 25740 9648
rect 29276 9596 29328 9648
rect 30380 9596 30432 9648
rect 31116 9596 31168 9648
rect 34244 9639 34296 9648
rect 34244 9605 34253 9639
rect 34253 9605 34287 9639
rect 34287 9605 34296 9639
rect 34244 9596 34296 9605
rect 26240 9528 26292 9580
rect 24216 9460 24268 9512
rect 25504 9503 25556 9512
rect 25504 9469 25513 9503
rect 25513 9469 25547 9503
rect 25547 9469 25556 9503
rect 25504 9460 25556 9469
rect 25964 9503 26016 9512
rect 25964 9469 25973 9503
rect 25973 9469 26007 9503
rect 26007 9469 26016 9503
rect 25964 9460 26016 9469
rect 27344 9460 27396 9512
rect 30288 9528 30340 9580
rect 28448 9503 28500 9512
rect 26884 9392 26936 9444
rect 24032 9367 24084 9376
rect 24032 9333 24041 9367
rect 24041 9333 24075 9367
rect 24075 9333 24084 9367
rect 28448 9469 28457 9503
rect 28457 9469 28491 9503
rect 28491 9469 28500 9503
rect 28448 9460 28500 9469
rect 29736 9460 29788 9512
rect 30840 9503 30892 9512
rect 27988 9392 28040 9444
rect 30840 9469 30849 9503
rect 30849 9469 30883 9503
rect 30883 9469 30892 9503
rect 30840 9460 30892 9469
rect 31300 9460 31352 9512
rect 24032 9324 24084 9333
rect 28172 9324 28224 9376
rect 32128 9460 32180 9512
rect 32312 9460 32364 9512
rect 32956 9503 33008 9512
rect 32956 9469 32965 9503
rect 32965 9469 32999 9503
rect 32999 9469 33008 9503
rect 32956 9460 33008 9469
rect 33416 9503 33468 9512
rect 33416 9469 33425 9503
rect 33425 9469 33459 9503
rect 33459 9469 33468 9503
rect 33416 9460 33468 9469
rect 34520 9460 34572 9512
rect 35532 9503 35584 9512
rect 35532 9469 35541 9503
rect 35541 9469 35575 9503
rect 35575 9469 35584 9503
rect 35532 9460 35584 9469
rect 35624 9460 35676 9512
rect 35808 9503 35860 9512
rect 35808 9469 35817 9503
rect 35817 9469 35851 9503
rect 35851 9469 35860 9503
rect 35808 9460 35860 9469
rect 35992 9460 36044 9512
rect 38016 9460 38068 9512
rect 32772 9392 32824 9444
rect 35348 9392 35400 9444
rect 31576 9324 31628 9376
rect 36268 9324 36320 9376
rect 19606 9222 19658 9274
rect 19670 9222 19722 9274
rect 19734 9222 19786 9274
rect 19798 9222 19850 9274
rect 8576 9120 8628 9172
rect 9772 9120 9824 9172
rect 4620 9052 4672 9104
rect 1400 8984 1452 9036
rect 2136 8959 2188 8968
rect 2136 8925 2145 8959
rect 2145 8925 2179 8959
rect 2179 8925 2188 8959
rect 2136 8916 2188 8925
rect 5540 8984 5592 9036
rect 6460 9027 6512 9036
rect 6460 8993 6469 9027
rect 6469 8993 6503 9027
rect 6503 8993 6512 9027
rect 6460 8984 6512 8993
rect 6828 9027 6880 9036
rect 6828 8993 6837 9027
rect 6837 8993 6871 9027
rect 6871 8993 6880 9027
rect 6828 8984 6880 8993
rect 7012 8984 7064 9036
rect 8300 8984 8352 9036
rect 6000 8916 6052 8968
rect 4712 8848 4764 8900
rect 7380 8780 7432 8832
rect 9680 9052 9732 9104
rect 9220 8984 9272 9036
rect 9496 8984 9548 9036
rect 10600 9027 10652 9036
rect 10600 8993 10609 9027
rect 10609 8993 10643 9027
rect 10643 8993 10652 9027
rect 10600 8984 10652 8993
rect 10784 8984 10836 9036
rect 9128 8916 9180 8968
rect 10324 8916 10376 8968
rect 14464 9052 14516 9104
rect 12072 9027 12124 9036
rect 12072 8993 12081 9027
rect 12081 8993 12115 9027
rect 12115 8993 12124 9027
rect 12072 8984 12124 8993
rect 13912 9027 13964 9036
rect 9772 8848 9824 8900
rect 8668 8780 8720 8832
rect 12164 8916 12216 8968
rect 13452 8959 13504 8968
rect 13452 8925 13461 8959
rect 13461 8925 13495 8959
rect 13495 8925 13504 8959
rect 13452 8916 13504 8925
rect 13912 8993 13921 9027
rect 13921 8993 13955 9027
rect 13955 8993 13964 9027
rect 13912 8984 13964 8993
rect 14004 9027 14056 9036
rect 14004 8993 14013 9027
rect 14013 8993 14047 9027
rect 14047 8993 14056 9027
rect 15660 9120 15712 9172
rect 17040 9163 17092 9172
rect 17040 9129 17049 9163
rect 17049 9129 17083 9163
rect 17083 9129 17092 9163
rect 17040 9120 17092 9129
rect 19984 9120 20036 9172
rect 21088 9120 21140 9172
rect 22836 9120 22888 9172
rect 27068 9120 27120 9172
rect 28356 9120 28408 9172
rect 14004 8984 14056 8993
rect 15476 9027 15528 9036
rect 15476 8993 15485 9027
rect 15485 8993 15519 9027
rect 15519 8993 15528 9027
rect 15476 8984 15528 8993
rect 15844 9027 15896 9036
rect 15844 8993 15853 9027
rect 15853 8993 15887 9027
rect 15887 8993 15896 9027
rect 15844 8984 15896 8993
rect 20628 9052 20680 9104
rect 22284 9052 22336 9104
rect 28816 9120 28868 9172
rect 16580 8984 16632 9036
rect 17040 8984 17092 9036
rect 13820 8916 13872 8968
rect 18420 8959 18472 8968
rect 18420 8925 18429 8959
rect 18429 8925 18463 8959
rect 18463 8925 18472 8959
rect 18420 8916 18472 8925
rect 19064 8984 19116 9036
rect 20812 8984 20864 9036
rect 21732 9027 21784 9036
rect 19248 8916 19300 8968
rect 20260 8959 20312 8968
rect 20260 8925 20269 8959
rect 20269 8925 20303 8959
rect 20303 8925 20312 8959
rect 20260 8916 20312 8925
rect 19892 8848 19944 8900
rect 20352 8848 20404 8900
rect 21732 8993 21741 9027
rect 21741 8993 21775 9027
rect 21775 8993 21784 9027
rect 21732 8984 21784 8993
rect 21824 8984 21876 9036
rect 26884 8984 26936 9036
rect 27528 9027 27580 9036
rect 27528 8993 27537 9027
rect 27537 8993 27571 9027
rect 27571 8993 27580 9027
rect 27528 8984 27580 8993
rect 27804 8984 27856 9036
rect 29184 9027 29236 9036
rect 29184 8993 29193 9027
rect 29193 8993 29227 9027
rect 29227 8993 29236 9027
rect 29184 8984 29236 8993
rect 29736 8984 29788 9036
rect 31300 9120 31352 9172
rect 31668 9120 31720 9172
rect 32404 9120 32456 9172
rect 31576 9052 31628 9104
rect 35440 9052 35492 9104
rect 31392 9027 31444 9036
rect 22284 8916 22336 8968
rect 23204 8959 23256 8968
rect 23204 8925 23213 8959
rect 23213 8925 23247 8959
rect 23247 8925 23256 8959
rect 23204 8916 23256 8925
rect 23480 8959 23532 8968
rect 23480 8925 23489 8959
rect 23489 8925 23523 8959
rect 23523 8925 23532 8959
rect 23480 8916 23532 8925
rect 28172 8959 28224 8968
rect 20904 8848 20956 8900
rect 26976 8848 27028 8900
rect 28172 8925 28181 8959
rect 28181 8925 28215 8959
rect 28215 8925 28224 8959
rect 28172 8916 28224 8925
rect 28724 8916 28776 8968
rect 31392 8993 31401 9027
rect 31401 8993 31435 9027
rect 31435 8993 31444 9027
rect 31392 8984 31444 8993
rect 31760 8984 31812 9036
rect 33048 9027 33100 9036
rect 33048 8993 33057 9027
rect 33057 8993 33091 9027
rect 33091 8993 33100 9027
rect 33048 8984 33100 8993
rect 36820 9027 36872 9036
rect 30012 8959 30064 8968
rect 30012 8925 30021 8959
rect 30021 8925 30055 8959
rect 30055 8925 30064 8959
rect 30012 8916 30064 8925
rect 31024 8916 31076 8968
rect 31300 8916 31352 8968
rect 27896 8848 27948 8900
rect 29828 8848 29880 8900
rect 12624 8780 12676 8832
rect 13268 8780 13320 8832
rect 15936 8780 15988 8832
rect 20168 8780 20220 8832
rect 22008 8780 22060 8832
rect 23848 8780 23900 8832
rect 25964 8780 26016 8832
rect 31944 8780 31996 8832
rect 34704 8916 34756 8968
rect 35440 8916 35492 8968
rect 35900 8959 35952 8968
rect 35900 8925 35909 8959
rect 35909 8925 35943 8959
rect 35943 8925 35952 8959
rect 35900 8916 35952 8925
rect 36820 8993 36829 9027
rect 36829 8993 36863 9027
rect 36863 8993 36872 9027
rect 36820 8984 36872 8993
rect 36360 8959 36412 8968
rect 36360 8925 36369 8959
rect 36369 8925 36403 8959
rect 36403 8925 36412 8959
rect 36360 8916 36412 8925
rect 37832 8848 37884 8900
rect 35532 8780 35584 8832
rect 4246 8678 4298 8730
rect 4310 8678 4362 8730
rect 4374 8678 4426 8730
rect 4438 8678 4490 8730
rect 34966 8678 35018 8730
rect 35030 8678 35082 8730
rect 35094 8678 35146 8730
rect 35158 8678 35210 8730
rect 1768 8619 1820 8628
rect 1768 8585 1777 8619
rect 1777 8585 1811 8619
rect 1811 8585 1820 8619
rect 1768 8576 1820 8585
rect 4896 8576 4948 8628
rect 6920 8619 6972 8628
rect 2964 8508 3016 8560
rect 2136 8440 2188 8492
rect 4712 8483 4764 8492
rect 4712 8449 4721 8483
rect 4721 8449 4755 8483
rect 4755 8449 4764 8483
rect 4712 8440 4764 8449
rect 1860 8372 1912 8424
rect 2320 8372 2372 8424
rect 2780 8304 2832 8356
rect 4160 8372 4212 8424
rect 5540 8372 5592 8424
rect 6920 8585 6929 8619
rect 6929 8585 6963 8619
rect 6963 8585 6972 8619
rect 6920 8576 6972 8585
rect 6000 8508 6052 8560
rect 8300 8551 8352 8560
rect 8300 8517 8309 8551
rect 8309 8517 8343 8551
rect 8343 8517 8352 8551
rect 8300 8508 8352 8517
rect 10784 8576 10836 8628
rect 13452 8576 13504 8628
rect 12256 8508 12308 8560
rect 15844 8576 15896 8628
rect 16120 8576 16172 8628
rect 15200 8508 15252 8560
rect 7380 8415 7432 8424
rect 7380 8381 7389 8415
rect 7389 8381 7423 8415
rect 7423 8381 7432 8415
rect 7380 8372 7432 8381
rect 8576 8415 8628 8424
rect 8576 8381 8585 8415
rect 8585 8381 8619 8415
rect 8619 8381 8628 8415
rect 9036 8440 9088 8492
rect 11888 8483 11940 8492
rect 11888 8449 11897 8483
rect 11897 8449 11931 8483
rect 11931 8449 11940 8483
rect 11888 8440 11940 8449
rect 8576 8372 8628 8381
rect 10416 8372 10468 8424
rect 11336 8415 11388 8424
rect 11336 8381 11345 8415
rect 11345 8381 11379 8415
rect 11379 8381 11388 8415
rect 11336 8372 11388 8381
rect 12624 8372 12676 8424
rect 12900 8415 12952 8424
rect 12900 8381 12909 8415
rect 12909 8381 12943 8415
rect 12943 8381 12952 8415
rect 12900 8372 12952 8381
rect 13268 8415 13320 8424
rect 13268 8381 13277 8415
rect 13277 8381 13311 8415
rect 13311 8381 13320 8415
rect 13268 8372 13320 8381
rect 13360 8415 13412 8424
rect 13360 8381 13369 8415
rect 13369 8381 13403 8415
rect 13403 8381 13412 8415
rect 13912 8415 13964 8424
rect 13360 8372 13412 8381
rect 13912 8381 13921 8415
rect 13921 8381 13955 8415
rect 13955 8381 13964 8415
rect 13912 8372 13964 8381
rect 14280 8372 14332 8424
rect 15476 8440 15528 8492
rect 16212 8415 16264 8424
rect 4528 8304 4580 8356
rect 5632 8304 5684 8356
rect 5908 8304 5960 8356
rect 11152 8304 11204 8356
rect 16212 8381 16221 8415
rect 16221 8381 16255 8415
rect 16255 8381 16264 8415
rect 16212 8372 16264 8381
rect 16580 8372 16632 8424
rect 17316 8415 17368 8424
rect 17316 8381 17325 8415
rect 17325 8381 17359 8415
rect 17359 8381 17368 8415
rect 17316 8372 17368 8381
rect 18604 8415 18656 8424
rect 18604 8381 18613 8415
rect 18613 8381 18647 8415
rect 18647 8381 18656 8415
rect 18604 8372 18656 8381
rect 23020 8576 23072 8628
rect 24400 8576 24452 8628
rect 35440 8576 35492 8628
rect 35992 8576 36044 8628
rect 36084 8576 36136 8628
rect 18972 8508 19024 8560
rect 19064 8483 19116 8492
rect 19064 8449 19073 8483
rect 19073 8449 19107 8483
rect 19107 8449 19116 8483
rect 19064 8440 19116 8449
rect 18972 8372 19024 8424
rect 21364 8508 21416 8560
rect 22376 8508 22428 8560
rect 24032 8508 24084 8560
rect 28724 8508 28776 8560
rect 18236 8304 18288 8356
rect 19064 8304 19116 8356
rect 19248 8304 19300 8356
rect 20260 8372 20312 8424
rect 20904 8440 20956 8492
rect 26792 8483 26844 8492
rect 26792 8449 26801 8483
rect 26801 8449 26835 8483
rect 26835 8449 26844 8483
rect 26792 8440 26844 8449
rect 20812 8372 20864 8424
rect 21180 8372 21232 8424
rect 21824 8372 21876 8424
rect 22376 8415 22428 8424
rect 20904 8304 20956 8356
rect 22376 8381 22385 8415
rect 22385 8381 22419 8415
rect 22419 8381 22428 8415
rect 22376 8372 22428 8381
rect 22468 8415 22520 8424
rect 22468 8381 22477 8415
rect 22477 8381 22511 8415
rect 22511 8381 22520 8415
rect 22468 8372 22520 8381
rect 22928 8372 22980 8424
rect 23204 8372 23256 8424
rect 23388 8372 23440 8424
rect 24216 8372 24268 8424
rect 26332 8372 26384 8424
rect 27068 8415 27120 8424
rect 27068 8381 27077 8415
rect 27077 8381 27111 8415
rect 27111 8381 27120 8415
rect 27068 8372 27120 8381
rect 27252 8415 27304 8424
rect 27252 8381 27261 8415
rect 27261 8381 27295 8415
rect 27295 8381 27304 8415
rect 27252 8372 27304 8381
rect 27344 8372 27396 8424
rect 27896 8372 27948 8424
rect 30932 8440 30984 8492
rect 33048 8508 33100 8560
rect 34336 8508 34388 8560
rect 9220 8236 9272 8288
rect 15844 8236 15896 8288
rect 16488 8236 16540 8288
rect 16948 8236 17000 8288
rect 17500 8236 17552 8288
rect 21088 8236 21140 8288
rect 27988 8304 28040 8356
rect 24400 8236 24452 8288
rect 30196 8372 30248 8424
rect 30472 8415 30524 8424
rect 30472 8381 30481 8415
rect 30481 8381 30515 8415
rect 30515 8381 30524 8415
rect 31024 8415 31076 8424
rect 30472 8372 30524 8381
rect 31024 8381 31033 8415
rect 31033 8381 31067 8415
rect 31067 8381 31076 8415
rect 31024 8372 31076 8381
rect 35900 8440 35952 8492
rect 32496 8372 32548 8424
rect 32772 8415 32824 8424
rect 32772 8381 32781 8415
rect 32781 8381 32815 8415
rect 32815 8381 32824 8415
rect 32772 8372 32824 8381
rect 32864 8372 32916 8424
rect 33416 8415 33468 8424
rect 33416 8381 33425 8415
rect 33425 8381 33459 8415
rect 33459 8381 33468 8415
rect 33416 8372 33468 8381
rect 34152 8415 34204 8424
rect 34152 8381 34161 8415
rect 34161 8381 34195 8415
rect 34195 8381 34204 8415
rect 34152 8372 34204 8381
rect 35532 8415 35584 8424
rect 35532 8381 35541 8415
rect 35541 8381 35575 8415
rect 35575 8381 35584 8415
rect 35532 8372 35584 8381
rect 35624 8372 35676 8424
rect 35256 8304 35308 8356
rect 35992 8372 36044 8424
rect 36268 8372 36320 8424
rect 30656 8236 30708 8288
rect 31116 8279 31168 8288
rect 31116 8245 31125 8279
rect 31125 8245 31159 8279
rect 31159 8245 31168 8279
rect 31116 8236 31168 8245
rect 19606 8134 19658 8186
rect 19670 8134 19722 8186
rect 19734 8134 19786 8186
rect 19798 8134 19850 8186
rect 2780 8075 2832 8084
rect 2780 8041 2789 8075
rect 2789 8041 2823 8075
rect 2823 8041 2832 8075
rect 2780 8032 2832 8041
rect 7840 8032 7892 8084
rect 8392 8032 8444 8084
rect 11796 8032 11848 8084
rect 13820 8032 13872 8084
rect 15200 8032 15252 8084
rect 15752 8032 15804 8084
rect 16028 8032 16080 8084
rect 1400 7939 1452 7948
rect 1400 7905 1409 7939
rect 1409 7905 1443 7939
rect 1443 7905 1452 7939
rect 1400 7896 1452 7905
rect 4160 7896 4212 7948
rect 4620 7896 4672 7948
rect 4988 7939 5040 7948
rect 4988 7905 4997 7939
rect 4997 7905 5031 7939
rect 5031 7905 5040 7939
rect 4988 7896 5040 7905
rect 6092 7896 6144 7948
rect 6644 7896 6696 7948
rect 9404 7964 9456 8016
rect 18236 8007 18288 8016
rect 7748 7939 7800 7948
rect 1676 7871 1728 7880
rect 1676 7837 1685 7871
rect 1685 7837 1719 7871
rect 1719 7837 1728 7871
rect 1676 7828 1728 7837
rect 6736 7871 6788 7880
rect 6736 7837 6745 7871
rect 6745 7837 6779 7871
rect 6779 7837 6788 7871
rect 6736 7828 6788 7837
rect 4804 7760 4856 7812
rect 6460 7760 6512 7812
rect 7748 7905 7757 7939
rect 7757 7905 7791 7939
rect 7791 7905 7800 7939
rect 7748 7896 7800 7905
rect 7932 7896 7984 7948
rect 8576 7896 8628 7948
rect 8760 7939 8812 7948
rect 8760 7905 8769 7939
rect 8769 7905 8803 7939
rect 8803 7905 8812 7939
rect 8760 7896 8812 7905
rect 10140 7896 10192 7948
rect 10692 7939 10744 7948
rect 10692 7905 10701 7939
rect 10701 7905 10735 7939
rect 10735 7905 10744 7939
rect 10692 7896 10744 7905
rect 10784 7896 10836 7948
rect 12164 7896 12216 7948
rect 12992 7939 13044 7948
rect 12992 7905 13001 7939
rect 13001 7905 13035 7939
rect 13035 7905 13044 7939
rect 12992 7896 13044 7905
rect 13636 7896 13688 7948
rect 7380 7828 7432 7880
rect 8392 7828 8444 7880
rect 11980 7828 12032 7880
rect 13360 7871 13412 7880
rect 13360 7837 13369 7871
rect 13369 7837 13403 7871
rect 13403 7837 13412 7871
rect 13360 7828 13412 7837
rect 14280 7896 14332 7948
rect 15660 7896 15712 7948
rect 16028 7896 16080 7948
rect 8852 7760 8904 7812
rect 11152 7760 11204 7812
rect 11336 7760 11388 7812
rect 14924 7828 14976 7880
rect 16580 7896 16632 7948
rect 16764 7896 16816 7948
rect 17500 7896 17552 7948
rect 17684 7896 17736 7948
rect 18236 7973 18245 8007
rect 18245 7973 18279 8007
rect 18279 7973 18288 8007
rect 18236 7964 18288 7973
rect 20168 8032 20220 8084
rect 20904 8032 20956 8084
rect 22100 8032 22152 8084
rect 23204 8032 23256 8084
rect 23480 8075 23532 8084
rect 23480 8041 23489 8075
rect 23489 8041 23523 8075
rect 23523 8041 23532 8075
rect 23480 8032 23532 8041
rect 27068 8032 27120 8084
rect 30104 8075 30156 8084
rect 30104 8041 30113 8075
rect 30113 8041 30147 8075
rect 30147 8041 30156 8075
rect 30104 8032 30156 8041
rect 30932 8032 30984 8084
rect 20812 7964 20864 8016
rect 16948 7828 17000 7880
rect 15568 7760 15620 7812
rect 8392 7692 8444 7744
rect 8760 7692 8812 7744
rect 11428 7692 11480 7744
rect 12256 7692 12308 7744
rect 16856 7692 16908 7744
rect 18420 7896 18472 7948
rect 18880 7939 18932 7948
rect 18880 7905 18889 7939
rect 18889 7905 18923 7939
rect 18923 7905 18932 7939
rect 18880 7896 18932 7905
rect 19064 7896 19116 7948
rect 19432 7896 19484 7948
rect 19892 7939 19944 7948
rect 19892 7905 19901 7939
rect 19901 7905 19935 7939
rect 19935 7905 19944 7939
rect 19892 7896 19944 7905
rect 20168 7896 20220 7948
rect 18420 7760 18472 7812
rect 19892 7760 19944 7812
rect 23756 7964 23808 8016
rect 24308 7964 24360 8016
rect 21824 7896 21876 7948
rect 22928 7896 22980 7948
rect 23204 7939 23256 7948
rect 23204 7905 23213 7939
rect 23213 7905 23247 7939
rect 23247 7905 23256 7939
rect 24400 7939 24452 7948
rect 23204 7896 23256 7905
rect 22008 7828 22060 7880
rect 24400 7905 24409 7939
rect 24409 7905 24443 7939
rect 24443 7905 24452 7939
rect 24400 7896 24452 7905
rect 25136 7939 25188 7948
rect 25136 7905 25145 7939
rect 25145 7905 25179 7939
rect 25179 7905 25188 7939
rect 25136 7896 25188 7905
rect 26976 7964 27028 8016
rect 27252 7896 27304 7948
rect 27436 7939 27488 7948
rect 27436 7905 27445 7939
rect 27445 7905 27479 7939
rect 27479 7905 27488 7939
rect 27436 7896 27488 7905
rect 27988 7939 28040 7948
rect 27988 7905 27997 7939
rect 27997 7905 28031 7939
rect 28031 7905 28040 7939
rect 27988 7896 28040 7905
rect 27160 7871 27212 7880
rect 27160 7837 27169 7871
rect 27169 7837 27203 7871
rect 27203 7837 27212 7871
rect 27160 7828 27212 7837
rect 30656 7964 30708 8016
rect 29368 7896 29420 7948
rect 30288 7896 30340 7948
rect 27252 7760 27304 7812
rect 21088 7692 21140 7744
rect 27344 7692 27396 7744
rect 30472 7828 30524 7880
rect 30104 7760 30156 7812
rect 32128 8032 32180 8084
rect 32312 8075 32364 8084
rect 32312 8041 32321 8075
rect 32321 8041 32355 8075
rect 32355 8041 32364 8075
rect 32312 8032 32364 8041
rect 32496 8032 32548 8084
rect 32404 7896 32456 7948
rect 33324 7896 33376 7948
rect 34060 7964 34112 8016
rect 33876 7939 33928 7948
rect 33876 7905 33885 7939
rect 33885 7905 33919 7939
rect 33919 7905 33928 7939
rect 33876 7896 33928 7905
rect 34244 7939 34296 7948
rect 34244 7905 34253 7939
rect 34253 7905 34287 7939
rect 34287 7905 34296 7939
rect 34244 7896 34296 7905
rect 35256 7896 35308 7948
rect 35440 7896 35492 7948
rect 34520 7828 34572 7880
rect 32220 7760 32272 7812
rect 29184 7692 29236 7744
rect 29460 7692 29512 7744
rect 30472 7692 30524 7744
rect 31484 7692 31536 7744
rect 4246 7590 4298 7642
rect 4310 7590 4362 7642
rect 4374 7590 4426 7642
rect 4438 7590 4490 7642
rect 34966 7590 35018 7642
rect 35030 7590 35082 7642
rect 35094 7590 35146 7642
rect 35158 7590 35210 7642
rect 4620 7488 4672 7540
rect 5356 7352 5408 7404
rect 9220 7488 9272 7540
rect 7748 7420 7800 7472
rect 10416 7463 10468 7472
rect 7932 7395 7984 7404
rect 2596 7327 2648 7336
rect 2596 7293 2605 7327
rect 2605 7293 2639 7327
rect 2639 7293 2648 7327
rect 2596 7284 2648 7293
rect 4160 7284 4212 7336
rect 4804 7327 4856 7336
rect 4804 7293 4813 7327
rect 4813 7293 4847 7327
rect 4847 7293 4856 7327
rect 4804 7284 4856 7293
rect 4988 7284 5040 7336
rect 7932 7361 7941 7395
rect 7941 7361 7975 7395
rect 7975 7361 7984 7395
rect 7932 7352 7984 7361
rect 6092 7284 6144 7336
rect 7380 7284 7432 7336
rect 7840 7327 7892 7336
rect 7840 7293 7849 7327
rect 7849 7293 7883 7327
rect 7883 7293 7892 7327
rect 7840 7284 7892 7293
rect 8852 7327 8904 7336
rect 8852 7293 8861 7327
rect 8861 7293 8895 7327
rect 8895 7293 8904 7327
rect 8852 7284 8904 7293
rect 10416 7429 10425 7463
rect 10425 7429 10459 7463
rect 10459 7429 10468 7463
rect 10416 7420 10468 7429
rect 9404 7352 9456 7404
rect 11060 7352 11112 7404
rect 10508 7284 10560 7336
rect 14188 7488 14240 7540
rect 13636 7463 13688 7472
rect 13636 7429 13645 7463
rect 13645 7429 13679 7463
rect 13679 7429 13688 7463
rect 13636 7420 13688 7429
rect 11796 7395 11848 7404
rect 11796 7361 11805 7395
rect 11805 7361 11839 7395
rect 11839 7361 11848 7395
rect 11796 7352 11848 7361
rect 14556 7395 14608 7404
rect 14556 7361 14565 7395
rect 14565 7361 14599 7395
rect 14599 7361 14608 7395
rect 14556 7352 14608 7361
rect 15936 7488 15988 7540
rect 17316 7488 17368 7540
rect 15568 7395 15620 7404
rect 15568 7361 15577 7395
rect 15577 7361 15611 7395
rect 15611 7361 15620 7395
rect 15568 7352 15620 7361
rect 15752 7352 15804 7404
rect 16488 7352 16540 7404
rect 11428 7284 11480 7336
rect 11704 7327 11756 7336
rect 11704 7293 11713 7327
rect 11713 7293 11747 7327
rect 11747 7293 11756 7327
rect 11704 7284 11756 7293
rect 6184 7191 6236 7200
rect 6184 7157 6193 7191
rect 6193 7157 6227 7191
rect 6227 7157 6236 7191
rect 6184 7148 6236 7157
rect 10416 7216 10468 7268
rect 12716 7216 12768 7268
rect 13912 7284 13964 7336
rect 14096 7327 14148 7336
rect 14096 7293 14105 7327
rect 14105 7293 14139 7327
rect 14139 7293 14148 7327
rect 14096 7284 14148 7293
rect 20628 7488 20680 7540
rect 22836 7488 22888 7540
rect 27436 7488 27488 7540
rect 30288 7488 30340 7540
rect 35440 7488 35492 7540
rect 37832 7531 37884 7540
rect 37832 7497 37841 7531
rect 37841 7497 37875 7531
rect 37875 7497 37884 7531
rect 37832 7488 37884 7497
rect 18420 7327 18472 7336
rect 18420 7293 18429 7327
rect 18429 7293 18463 7327
rect 18463 7293 18472 7327
rect 21732 7420 21784 7472
rect 19156 7395 19208 7404
rect 19156 7361 19165 7395
rect 19165 7361 19199 7395
rect 19199 7361 19208 7395
rect 19156 7352 19208 7361
rect 19892 7395 19944 7404
rect 19892 7361 19901 7395
rect 19901 7361 19935 7395
rect 19935 7361 19944 7395
rect 19892 7352 19944 7361
rect 22192 7395 22244 7404
rect 22192 7361 22201 7395
rect 22201 7361 22235 7395
rect 22235 7361 22244 7395
rect 22192 7352 22244 7361
rect 18420 7284 18472 7293
rect 19340 7284 19392 7336
rect 20536 7327 20588 7336
rect 20168 7216 20220 7268
rect 20536 7293 20545 7327
rect 20545 7293 20579 7327
rect 20579 7293 20588 7327
rect 20536 7284 20588 7293
rect 21916 7327 21968 7336
rect 21916 7293 21925 7327
rect 21925 7293 21959 7327
rect 21959 7293 21968 7327
rect 21916 7284 21968 7293
rect 22100 7284 22152 7336
rect 24308 7420 24360 7472
rect 25136 7420 25188 7472
rect 29276 7420 29328 7472
rect 29460 7420 29512 7472
rect 33416 7463 33468 7472
rect 26884 7395 26936 7404
rect 26884 7361 26893 7395
rect 26893 7361 26927 7395
rect 26927 7361 26936 7395
rect 26884 7352 26936 7361
rect 27344 7352 27396 7404
rect 33416 7429 33425 7463
rect 33425 7429 33459 7463
rect 33459 7429 33468 7463
rect 33416 7420 33468 7429
rect 36176 7420 36228 7472
rect 22836 7284 22888 7336
rect 23848 7327 23900 7336
rect 23848 7293 23857 7327
rect 23857 7293 23891 7327
rect 23891 7293 23900 7327
rect 23848 7284 23900 7293
rect 20812 7216 20864 7268
rect 21272 7216 21324 7268
rect 11980 7148 12032 7200
rect 12164 7148 12216 7200
rect 15568 7148 15620 7200
rect 16488 7148 16540 7200
rect 22284 7216 22336 7268
rect 24400 7327 24452 7336
rect 24400 7293 24409 7327
rect 24409 7293 24443 7327
rect 24443 7293 24452 7327
rect 24584 7327 24636 7336
rect 24400 7284 24452 7293
rect 24584 7293 24593 7327
rect 24593 7293 24627 7327
rect 24627 7293 24636 7327
rect 24584 7284 24636 7293
rect 25596 7284 25648 7336
rect 26332 7284 26384 7336
rect 26976 7327 27028 7336
rect 26976 7293 26985 7327
rect 26985 7293 27019 7327
rect 27019 7293 27028 7327
rect 26976 7284 27028 7293
rect 27252 7327 27304 7336
rect 27252 7293 27261 7327
rect 27261 7293 27295 7327
rect 27295 7293 27304 7327
rect 27252 7284 27304 7293
rect 27896 7327 27948 7336
rect 27896 7293 27905 7327
rect 27905 7293 27939 7327
rect 27939 7293 27948 7327
rect 27896 7284 27948 7293
rect 28264 7284 28316 7336
rect 29552 7284 29604 7336
rect 31116 7352 31168 7404
rect 30840 7284 30892 7336
rect 33324 7352 33376 7404
rect 34244 7352 34296 7404
rect 35348 7352 35400 7404
rect 36360 7352 36412 7404
rect 33232 7284 33284 7336
rect 35716 7284 35768 7336
rect 36084 7284 36136 7336
rect 36176 7284 36228 7336
rect 21824 7148 21876 7200
rect 24400 7148 24452 7200
rect 24860 7191 24912 7200
rect 24860 7157 24869 7191
rect 24869 7157 24903 7191
rect 24903 7157 24912 7191
rect 24860 7148 24912 7157
rect 27528 7216 27580 7268
rect 29000 7216 29052 7268
rect 30748 7148 30800 7200
rect 19606 7046 19658 7098
rect 19670 7046 19722 7098
rect 19734 7046 19786 7098
rect 19798 7046 19850 7098
rect 7012 6944 7064 6996
rect 2596 6808 2648 6860
rect 2136 6783 2188 6792
rect 2136 6749 2145 6783
rect 2145 6749 2179 6783
rect 2179 6749 2188 6783
rect 2136 6740 2188 6749
rect 3424 6647 3476 6656
rect 3424 6613 3433 6647
rect 3433 6613 3467 6647
rect 3467 6613 3476 6647
rect 3424 6604 3476 6613
rect 4712 6851 4764 6860
rect 4160 6783 4212 6792
rect 4160 6749 4169 6783
rect 4169 6749 4203 6783
rect 4203 6749 4212 6783
rect 4160 6740 4212 6749
rect 4712 6817 4721 6851
rect 4721 6817 4755 6851
rect 4755 6817 4764 6851
rect 4712 6808 4764 6817
rect 5908 6851 5960 6860
rect 4620 6740 4672 6792
rect 5908 6817 5917 6851
rect 5917 6817 5951 6851
rect 5951 6817 5960 6851
rect 5908 6808 5960 6817
rect 7472 6876 7524 6928
rect 6736 6851 6788 6860
rect 6184 6740 6236 6792
rect 6460 6783 6512 6792
rect 6460 6749 6469 6783
rect 6469 6749 6503 6783
rect 6503 6749 6512 6783
rect 6460 6740 6512 6749
rect 6736 6817 6745 6851
rect 6745 6817 6779 6851
rect 6779 6817 6788 6851
rect 6736 6808 6788 6817
rect 10968 6876 11020 6928
rect 11704 6944 11756 6996
rect 15936 6944 15988 6996
rect 20260 6944 20312 6996
rect 21548 6944 21600 6996
rect 21916 6944 21968 6996
rect 23664 6944 23716 6996
rect 31944 6944 31996 6996
rect 32128 6944 32180 6996
rect 36360 6944 36412 6996
rect 12164 6876 12216 6928
rect 15568 6876 15620 6928
rect 10140 6851 10192 6860
rect 10140 6817 10149 6851
rect 10149 6817 10183 6851
rect 10183 6817 10192 6851
rect 10140 6808 10192 6817
rect 10232 6808 10284 6860
rect 5264 6672 5316 6724
rect 4988 6604 5040 6656
rect 5080 6604 5132 6656
rect 12164 6740 12216 6792
rect 8944 6672 8996 6724
rect 12440 6808 12492 6860
rect 13912 6808 13964 6860
rect 12532 6783 12584 6792
rect 12532 6749 12541 6783
rect 12541 6749 12575 6783
rect 12575 6749 12584 6783
rect 12532 6740 12584 6749
rect 14096 6808 14148 6860
rect 15476 6851 15528 6860
rect 15476 6817 15485 6851
rect 15485 6817 15519 6851
rect 15519 6817 15528 6851
rect 15476 6808 15528 6817
rect 15844 6851 15896 6860
rect 15844 6817 15853 6851
rect 15853 6817 15887 6851
rect 15887 6817 15896 6851
rect 15844 6808 15896 6817
rect 16856 6851 16908 6860
rect 14464 6783 14516 6792
rect 14464 6749 14473 6783
rect 14473 6749 14507 6783
rect 14507 6749 14516 6783
rect 14464 6740 14516 6749
rect 15568 6740 15620 6792
rect 16856 6817 16865 6851
rect 16865 6817 16899 6851
rect 16899 6817 16908 6851
rect 16856 6808 16908 6817
rect 17316 6851 17368 6860
rect 17316 6817 17325 6851
rect 17325 6817 17359 6851
rect 17359 6817 17368 6851
rect 17316 6808 17368 6817
rect 17500 6851 17552 6860
rect 17500 6817 17509 6851
rect 17509 6817 17543 6851
rect 17543 6817 17552 6851
rect 17500 6808 17552 6817
rect 19984 6876 20036 6928
rect 22008 6876 22060 6928
rect 18236 6740 18288 6792
rect 21640 6808 21692 6860
rect 22468 6808 22520 6860
rect 22100 6740 22152 6792
rect 22652 6808 22704 6860
rect 23112 6808 23164 6860
rect 23388 6808 23440 6860
rect 24860 6808 24912 6860
rect 25688 6808 25740 6860
rect 24584 6740 24636 6792
rect 25504 6740 25556 6792
rect 27068 6783 27120 6792
rect 27068 6749 27077 6783
rect 27077 6749 27111 6783
rect 27111 6749 27120 6783
rect 27068 6740 27120 6749
rect 27344 6808 27396 6860
rect 27896 6851 27948 6860
rect 27896 6817 27905 6851
rect 27905 6817 27939 6851
rect 27939 6817 27948 6851
rect 27896 6808 27948 6817
rect 29000 6808 29052 6860
rect 29736 6876 29788 6928
rect 30840 6876 30892 6928
rect 27436 6740 27488 6792
rect 28172 6740 28224 6792
rect 29552 6808 29604 6860
rect 33048 6876 33100 6928
rect 29276 6740 29328 6792
rect 31300 6740 31352 6792
rect 13084 6672 13136 6724
rect 15384 6715 15436 6724
rect 15384 6681 15393 6715
rect 15393 6681 15427 6715
rect 15427 6681 15436 6715
rect 15384 6672 15436 6681
rect 16120 6672 16172 6724
rect 21824 6672 21876 6724
rect 10508 6604 10560 6656
rect 15292 6604 15344 6656
rect 20536 6604 20588 6656
rect 22560 6647 22612 6656
rect 22560 6613 22569 6647
rect 22569 6613 22603 6647
rect 22603 6613 22612 6647
rect 22560 6604 22612 6613
rect 31024 6672 31076 6724
rect 31484 6851 31536 6860
rect 31484 6817 31493 6851
rect 31493 6817 31527 6851
rect 31527 6817 31536 6851
rect 31484 6808 31536 6817
rect 31668 6808 31720 6860
rect 32312 6851 32364 6860
rect 32312 6817 32321 6851
rect 32321 6817 32355 6851
rect 32355 6817 32364 6851
rect 32312 6808 32364 6817
rect 31576 6740 31628 6792
rect 33600 6808 33652 6860
rect 34244 6851 34296 6860
rect 34244 6817 34253 6851
rect 34253 6817 34287 6851
rect 34287 6817 34296 6851
rect 34244 6808 34296 6817
rect 32496 6740 32548 6792
rect 33968 6783 34020 6792
rect 33968 6749 33977 6783
rect 33977 6749 34011 6783
rect 34011 6749 34020 6783
rect 33968 6740 34020 6749
rect 34520 6740 34572 6792
rect 34704 6740 34756 6792
rect 35440 6783 35492 6792
rect 35440 6749 35449 6783
rect 35449 6749 35483 6783
rect 35483 6749 35492 6783
rect 35440 6740 35492 6749
rect 35808 6808 35860 6860
rect 35992 6808 36044 6860
rect 37372 6740 37424 6792
rect 29552 6604 29604 6656
rect 29736 6604 29788 6656
rect 32220 6604 32272 6656
rect 33232 6604 33284 6656
rect 33692 6604 33744 6656
rect 4246 6502 4298 6554
rect 4310 6502 4362 6554
rect 4374 6502 4426 6554
rect 4438 6502 4490 6554
rect 34966 6502 35018 6554
rect 35030 6502 35082 6554
rect 35094 6502 35146 6554
rect 35158 6502 35210 6554
rect 2136 6332 2188 6384
rect 1860 6239 1912 6248
rect 1860 6205 1869 6239
rect 1869 6205 1903 6239
rect 1903 6205 1912 6239
rect 1860 6196 1912 6205
rect 4068 6196 4120 6248
rect 4620 6196 4672 6248
rect 8576 6400 8628 6452
rect 12532 6400 12584 6452
rect 15292 6400 15344 6452
rect 25136 6400 25188 6452
rect 27436 6400 27488 6452
rect 13268 6332 13320 6384
rect 4988 6264 5040 6316
rect 5540 6264 5592 6316
rect 6460 6264 6512 6316
rect 7932 6264 7984 6316
rect 9496 6264 9548 6316
rect 5264 6128 5316 6180
rect 6000 6196 6052 6248
rect 7012 6196 7064 6248
rect 7472 6196 7524 6248
rect 10140 6239 10192 6248
rect 10140 6205 10149 6239
rect 10149 6205 10183 6239
rect 10183 6205 10192 6239
rect 10140 6196 10192 6205
rect 14740 6332 14792 6384
rect 20168 6375 20220 6384
rect 20168 6341 20177 6375
rect 20177 6341 20211 6375
rect 20211 6341 20220 6375
rect 20168 6332 20220 6341
rect 29276 6332 29328 6384
rect 30932 6400 30984 6452
rect 31208 6400 31260 6452
rect 37740 6400 37792 6452
rect 32312 6332 32364 6384
rect 14464 6264 14516 6316
rect 16120 6307 16172 6316
rect 5908 6128 5960 6180
rect 11244 6196 11296 6248
rect 11980 6196 12032 6248
rect 12440 6239 12492 6248
rect 12440 6205 12449 6239
rect 12449 6205 12483 6239
rect 12483 6205 12492 6239
rect 12440 6196 12492 6205
rect 12716 6196 12768 6248
rect 13912 6196 13964 6248
rect 1676 6060 1728 6112
rect 6000 6103 6052 6112
rect 6000 6069 6009 6103
rect 6009 6069 6043 6103
rect 6043 6069 6052 6103
rect 6000 6060 6052 6069
rect 6828 6060 6880 6112
rect 7288 6060 7340 6112
rect 10600 6128 10652 6180
rect 12808 6128 12860 6180
rect 9680 6060 9732 6112
rect 10232 6060 10284 6112
rect 15568 6196 15620 6248
rect 16120 6273 16129 6307
rect 16129 6273 16163 6307
rect 16163 6273 16172 6307
rect 16120 6264 16172 6273
rect 29552 6307 29604 6316
rect 29552 6273 29561 6307
rect 29561 6273 29595 6307
rect 29595 6273 29604 6307
rect 29552 6264 29604 6273
rect 30196 6264 30248 6316
rect 31208 6264 31260 6316
rect 32220 6264 32272 6316
rect 32496 6332 32548 6384
rect 19156 6196 19208 6248
rect 21364 6239 21416 6248
rect 21364 6205 21373 6239
rect 21373 6205 21407 6239
rect 21407 6205 21416 6239
rect 21364 6196 21416 6205
rect 22008 6239 22060 6248
rect 22008 6205 22017 6239
rect 22017 6205 22051 6239
rect 22051 6205 22060 6239
rect 22008 6196 22060 6205
rect 22836 6196 22888 6248
rect 23572 6196 23624 6248
rect 14556 6060 14608 6112
rect 14832 6060 14884 6112
rect 17316 6060 17368 6112
rect 23664 6060 23716 6112
rect 25136 6196 25188 6248
rect 25320 6196 25372 6248
rect 27896 6196 27948 6248
rect 27988 6196 28040 6248
rect 28540 6239 28592 6248
rect 28540 6205 28549 6239
rect 28549 6205 28583 6239
rect 28583 6205 28592 6239
rect 28540 6196 28592 6205
rect 29184 6196 29236 6248
rect 27712 6171 27764 6180
rect 27712 6137 27721 6171
rect 27721 6137 27755 6171
rect 27755 6137 27764 6171
rect 27712 6128 27764 6137
rect 27804 6128 27856 6180
rect 30564 6196 30616 6248
rect 31944 6196 31996 6248
rect 33048 6264 33100 6316
rect 34520 6332 34572 6384
rect 35716 6332 35768 6384
rect 35440 6264 35492 6316
rect 35900 6264 35952 6316
rect 34152 6239 34204 6248
rect 33324 6171 33376 6180
rect 33324 6137 33333 6171
rect 33333 6137 33367 6171
rect 33367 6137 33376 6171
rect 33324 6128 33376 6137
rect 34152 6205 34161 6239
rect 34161 6205 34195 6239
rect 34195 6205 34204 6239
rect 34152 6196 34204 6205
rect 34520 6196 34572 6248
rect 35532 6239 35584 6248
rect 35532 6205 35541 6239
rect 35541 6205 35575 6239
rect 35575 6205 35584 6239
rect 35532 6196 35584 6205
rect 35624 6196 35676 6248
rect 36084 6196 36136 6248
rect 37004 6239 37056 6248
rect 37004 6205 37013 6239
rect 37013 6205 37047 6239
rect 37047 6205 37056 6239
rect 37004 6196 37056 6205
rect 37280 6239 37332 6248
rect 37280 6205 37289 6239
rect 37289 6205 37323 6239
rect 37323 6205 37332 6239
rect 37280 6196 37332 6205
rect 37464 6239 37516 6248
rect 37464 6205 37473 6239
rect 37473 6205 37507 6239
rect 37507 6205 37516 6239
rect 37464 6196 37516 6205
rect 37556 6196 37608 6248
rect 29092 6060 29144 6112
rect 29644 6060 29696 6112
rect 30472 6060 30524 6112
rect 32220 6060 32272 6112
rect 35624 6060 35676 6112
rect 19606 5958 19658 6010
rect 19670 5958 19722 6010
rect 19734 5958 19786 6010
rect 19798 5958 19850 6010
rect 2780 5899 2832 5908
rect 2780 5865 2789 5899
rect 2789 5865 2823 5899
rect 2823 5865 2832 5899
rect 2780 5856 2832 5865
rect 4068 5856 4120 5908
rect 3424 5720 3476 5772
rect 8576 5856 8628 5908
rect 11244 5856 11296 5908
rect 13268 5856 13320 5908
rect 6184 5788 6236 5840
rect 5080 5763 5132 5772
rect 5080 5729 5089 5763
rect 5089 5729 5123 5763
rect 5123 5729 5132 5763
rect 5080 5720 5132 5729
rect 5264 5720 5316 5772
rect 6000 5720 6052 5772
rect 6828 5788 6880 5840
rect 9496 5788 9548 5840
rect 1400 5695 1452 5704
rect 1400 5661 1409 5695
rect 1409 5661 1443 5695
rect 1443 5661 1452 5695
rect 1400 5652 1452 5661
rect 1676 5695 1728 5704
rect 1676 5661 1685 5695
rect 1685 5661 1719 5695
rect 1719 5661 1728 5695
rect 1676 5652 1728 5661
rect 7196 5652 7248 5704
rect 8300 5763 8352 5772
rect 8300 5729 8309 5763
rect 8309 5729 8343 5763
rect 8343 5729 8352 5763
rect 8300 5720 8352 5729
rect 8484 5720 8536 5772
rect 9036 5720 9088 5772
rect 9680 5763 9732 5772
rect 9680 5729 9689 5763
rect 9689 5729 9723 5763
rect 9723 5729 9732 5763
rect 9680 5720 9732 5729
rect 12532 5788 12584 5840
rect 11060 5763 11112 5772
rect 11060 5729 11069 5763
rect 11069 5729 11103 5763
rect 11103 5729 11112 5763
rect 11060 5720 11112 5729
rect 11980 5763 12032 5772
rect 11980 5729 11989 5763
rect 11989 5729 12023 5763
rect 12023 5729 12032 5763
rect 11980 5720 12032 5729
rect 12624 5720 12676 5772
rect 15568 5788 15620 5840
rect 16672 5856 16724 5908
rect 22192 5856 22244 5908
rect 27068 5899 27120 5908
rect 27068 5865 27077 5899
rect 27077 5865 27111 5899
rect 27111 5865 27120 5899
rect 27068 5856 27120 5865
rect 27712 5856 27764 5908
rect 36636 5856 36688 5908
rect 19984 5788 20036 5840
rect 20720 5788 20772 5840
rect 13728 5763 13780 5772
rect 10968 5652 11020 5704
rect 12716 5695 12768 5704
rect 12716 5661 12725 5695
rect 12725 5661 12759 5695
rect 12759 5661 12768 5695
rect 12716 5652 12768 5661
rect 13728 5729 13737 5763
rect 13737 5729 13771 5763
rect 13771 5729 13780 5763
rect 13728 5720 13780 5729
rect 12992 5652 13044 5704
rect 15660 5720 15712 5772
rect 15844 5763 15896 5772
rect 15844 5729 15853 5763
rect 15853 5729 15887 5763
rect 15887 5729 15896 5763
rect 15844 5720 15896 5729
rect 16672 5763 16724 5772
rect 16672 5729 16681 5763
rect 16681 5729 16715 5763
rect 16715 5729 16724 5763
rect 16672 5720 16724 5729
rect 17684 5763 17736 5772
rect 17684 5729 17693 5763
rect 17693 5729 17727 5763
rect 17727 5729 17736 5763
rect 17684 5720 17736 5729
rect 18512 5720 18564 5772
rect 19340 5763 19392 5772
rect 19340 5729 19349 5763
rect 19349 5729 19383 5763
rect 19383 5729 19392 5763
rect 19340 5720 19392 5729
rect 19892 5763 19944 5772
rect 19892 5729 19901 5763
rect 19901 5729 19935 5763
rect 19935 5729 19944 5763
rect 19892 5720 19944 5729
rect 7288 5584 7340 5636
rect 9496 5584 9548 5636
rect 16580 5652 16632 5704
rect 17868 5652 17920 5704
rect 15016 5584 15068 5636
rect 19156 5652 19208 5704
rect 19892 5584 19944 5636
rect 20260 5584 20312 5636
rect 20996 5763 21048 5772
rect 20996 5729 21005 5763
rect 21005 5729 21039 5763
rect 21039 5729 21048 5763
rect 21732 5788 21784 5840
rect 25320 5831 25372 5840
rect 20996 5720 21048 5729
rect 22468 5763 22520 5772
rect 22468 5729 22477 5763
rect 22477 5729 22511 5763
rect 22511 5729 22520 5763
rect 22468 5720 22520 5729
rect 22652 5763 22704 5772
rect 22652 5729 22661 5763
rect 22661 5729 22695 5763
rect 22695 5729 22704 5763
rect 22652 5720 22704 5729
rect 23112 5763 23164 5772
rect 23112 5729 23121 5763
rect 23121 5729 23155 5763
rect 23155 5729 23164 5763
rect 23112 5720 23164 5729
rect 23848 5720 23900 5772
rect 24124 5720 24176 5772
rect 24308 5720 24360 5772
rect 24676 5720 24728 5772
rect 25320 5797 25329 5831
rect 25329 5797 25363 5831
rect 25363 5797 25372 5831
rect 25320 5788 25372 5797
rect 26792 5831 26844 5840
rect 26792 5797 26801 5831
rect 26801 5797 26835 5831
rect 26835 5797 26844 5831
rect 26792 5788 26844 5797
rect 26884 5788 26936 5840
rect 27160 5831 27212 5840
rect 27160 5797 27169 5831
rect 27169 5797 27203 5831
rect 27203 5797 27212 5831
rect 27160 5788 27212 5797
rect 27804 5788 27856 5840
rect 27988 5831 28040 5840
rect 27988 5797 27997 5831
rect 27997 5797 28031 5831
rect 28031 5797 28040 5831
rect 27988 5788 28040 5797
rect 28540 5788 28592 5840
rect 30196 5788 30248 5840
rect 27436 5720 27488 5772
rect 28816 5763 28868 5772
rect 28816 5729 28825 5763
rect 28825 5729 28859 5763
rect 28859 5729 28868 5763
rect 28816 5720 28868 5729
rect 28908 5720 28960 5772
rect 32220 5788 32272 5840
rect 36084 5831 36136 5840
rect 36084 5797 36093 5831
rect 36093 5797 36127 5831
rect 36127 5797 36136 5831
rect 36084 5788 36136 5797
rect 22284 5695 22336 5704
rect 22284 5661 22293 5695
rect 22293 5661 22327 5695
rect 22327 5661 22336 5695
rect 22284 5652 22336 5661
rect 30012 5695 30064 5704
rect 21364 5584 21416 5636
rect 26240 5584 26292 5636
rect 30012 5661 30021 5695
rect 30021 5661 30055 5695
rect 30055 5661 30064 5695
rect 30012 5652 30064 5661
rect 30472 5695 30524 5704
rect 30472 5661 30481 5695
rect 30481 5661 30515 5695
rect 30515 5661 30524 5695
rect 30472 5652 30524 5661
rect 31208 5652 31260 5704
rect 32772 5720 32824 5772
rect 34704 5763 34756 5772
rect 32036 5652 32088 5704
rect 32128 5695 32180 5704
rect 32128 5661 32137 5695
rect 32137 5661 32171 5695
rect 32171 5661 32180 5695
rect 32404 5695 32456 5704
rect 32128 5652 32180 5661
rect 32404 5661 32413 5695
rect 32413 5661 32447 5695
rect 32447 5661 32456 5695
rect 32404 5652 32456 5661
rect 32496 5652 32548 5704
rect 34704 5729 34713 5763
rect 34713 5729 34747 5763
rect 34747 5729 34756 5763
rect 34704 5720 34756 5729
rect 35808 5720 35860 5772
rect 36728 5720 36780 5772
rect 31944 5584 31996 5636
rect 6644 5516 6696 5568
rect 7472 5516 7524 5568
rect 11520 5516 11572 5568
rect 13728 5516 13780 5568
rect 14648 5559 14700 5568
rect 14648 5525 14657 5559
rect 14657 5525 14691 5559
rect 14691 5525 14700 5559
rect 14648 5516 14700 5525
rect 15568 5516 15620 5568
rect 21640 5559 21692 5568
rect 21640 5525 21649 5559
rect 21649 5525 21683 5559
rect 21683 5525 21692 5559
rect 21640 5516 21692 5525
rect 29000 5516 29052 5568
rect 30932 5516 30984 5568
rect 37924 5627 37976 5636
rect 37924 5593 37933 5627
rect 37933 5593 37967 5627
rect 37967 5593 37976 5627
rect 37924 5584 37976 5593
rect 36084 5516 36136 5568
rect 4246 5414 4298 5466
rect 4310 5414 4362 5466
rect 4374 5414 4426 5466
rect 4438 5414 4490 5466
rect 34966 5414 35018 5466
rect 35030 5414 35082 5466
rect 35094 5414 35146 5466
rect 35158 5414 35210 5466
rect 1676 5312 1728 5364
rect 3240 5176 3292 5228
rect 2044 5151 2096 5160
rect 2044 5117 2053 5151
rect 2053 5117 2087 5151
rect 2087 5117 2096 5151
rect 2044 5108 2096 5117
rect 3792 5151 3844 5160
rect 2964 4972 3016 5024
rect 3424 4972 3476 5024
rect 3792 5117 3801 5151
rect 3801 5117 3835 5151
rect 3835 5117 3844 5151
rect 3792 5108 3844 5117
rect 4620 5108 4672 5160
rect 16672 5312 16724 5364
rect 20260 5312 20312 5364
rect 23112 5312 23164 5364
rect 26884 5312 26936 5364
rect 30932 5312 30984 5364
rect 32864 5312 32916 5364
rect 33508 5312 33560 5364
rect 37372 5312 37424 5364
rect 7288 5244 7340 5296
rect 12440 5244 12492 5296
rect 13912 5287 13964 5296
rect 7380 5176 7432 5228
rect 5816 5108 5868 5160
rect 7012 5108 7064 5160
rect 7472 5151 7524 5160
rect 7472 5117 7481 5151
rect 7481 5117 7515 5151
rect 7515 5117 7524 5151
rect 7472 5108 7524 5117
rect 10232 5151 10284 5160
rect 5264 4972 5316 5024
rect 6828 4972 6880 5024
rect 10232 5117 10241 5151
rect 10241 5117 10275 5151
rect 10275 5117 10284 5151
rect 10232 5108 10284 5117
rect 10876 5176 10928 5228
rect 12992 5176 13044 5228
rect 10968 5151 11020 5160
rect 10968 5117 10977 5151
rect 10977 5117 11011 5151
rect 11011 5117 11020 5151
rect 10968 5108 11020 5117
rect 11520 5151 11572 5160
rect 11520 5117 11529 5151
rect 11529 5117 11563 5151
rect 11563 5117 11572 5151
rect 11520 5108 11572 5117
rect 13912 5253 13921 5287
rect 13921 5253 13955 5287
rect 13955 5253 13964 5287
rect 13912 5244 13964 5253
rect 22652 5244 22704 5296
rect 31116 5244 31168 5296
rect 13728 5176 13780 5228
rect 19340 5176 19392 5228
rect 14280 5151 14332 5160
rect 14280 5117 14289 5151
rect 14289 5117 14323 5151
rect 14323 5117 14332 5151
rect 14280 5108 14332 5117
rect 14648 5151 14700 5160
rect 14648 5117 14657 5151
rect 14657 5117 14691 5151
rect 14691 5117 14700 5151
rect 14648 5108 14700 5117
rect 15200 5108 15252 5160
rect 15568 5151 15620 5160
rect 15568 5117 15577 5151
rect 15577 5117 15611 5151
rect 15611 5117 15620 5151
rect 15568 5108 15620 5117
rect 16488 5151 16540 5160
rect 16488 5117 16497 5151
rect 16497 5117 16531 5151
rect 16531 5117 16540 5151
rect 16488 5108 16540 5117
rect 16948 5151 17000 5160
rect 16948 5117 16957 5151
rect 16957 5117 16991 5151
rect 16991 5117 17000 5151
rect 16948 5108 17000 5117
rect 15936 5040 15988 5092
rect 18604 5151 18656 5160
rect 18604 5117 18613 5151
rect 18613 5117 18647 5151
rect 18647 5117 18656 5151
rect 18604 5108 18656 5117
rect 19432 5108 19484 5160
rect 20812 5176 20864 5228
rect 21272 5176 21324 5228
rect 21640 5108 21692 5160
rect 24860 5176 24912 5228
rect 25136 5176 25188 5228
rect 26792 5176 26844 5228
rect 29184 5176 29236 5228
rect 30012 5176 30064 5228
rect 34428 5244 34480 5296
rect 22928 5151 22980 5160
rect 18328 5040 18380 5092
rect 20628 5040 20680 5092
rect 20720 5083 20772 5092
rect 20720 5049 20729 5083
rect 20729 5049 20763 5083
rect 20763 5049 20772 5083
rect 20720 5040 20772 5049
rect 10232 4972 10284 5024
rect 11980 4972 12032 5024
rect 17960 4972 18012 5024
rect 20904 4972 20956 5024
rect 22928 5117 22937 5151
rect 22937 5117 22971 5151
rect 22971 5117 22980 5151
rect 22928 5108 22980 5117
rect 23664 5151 23716 5160
rect 23664 5117 23673 5151
rect 23673 5117 23707 5151
rect 23707 5117 23716 5151
rect 23664 5108 23716 5117
rect 25228 5151 25280 5160
rect 25228 5117 25237 5151
rect 25237 5117 25271 5151
rect 25271 5117 25280 5151
rect 25228 5108 25280 5117
rect 30656 5151 30708 5160
rect 27160 5040 27212 5092
rect 30656 5117 30665 5151
rect 30665 5117 30699 5151
rect 30699 5117 30708 5151
rect 30656 5108 30708 5117
rect 30840 5151 30892 5160
rect 30840 5117 30849 5151
rect 30849 5117 30883 5151
rect 30883 5117 30892 5151
rect 30840 5108 30892 5117
rect 31760 5108 31812 5160
rect 35808 5176 35860 5228
rect 36636 5219 36688 5228
rect 36636 5185 36645 5219
rect 36645 5185 36679 5219
rect 36679 5185 36688 5219
rect 36636 5176 36688 5185
rect 32864 5108 32916 5160
rect 31116 5040 31168 5092
rect 32680 5040 32732 5092
rect 33232 5108 33284 5160
rect 33600 5108 33652 5160
rect 35716 5151 35768 5160
rect 35716 5117 35725 5151
rect 35725 5117 35759 5151
rect 35759 5117 35768 5151
rect 35716 5108 35768 5117
rect 36084 5108 36136 5160
rect 28172 4972 28224 5024
rect 31760 4972 31812 5024
rect 32956 4972 33008 5024
rect 19606 4870 19658 4922
rect 19670 4870 19722 4922
rect 19734 4870 19786 4922
rect 19798 4870 19850 4922
rect 2044 4768 2096 4820
rect 6368 4700 6420 4752
rect 5264 4675 5316 4684
rect 5264 4641 5273 4675
rect 5273 4641 5307 4675
rect 5307 4641 5316 4675
rect 5264 4632 5316 4641
rect 1400 4607 1452 4616
rect 1400 4573 1409 4607
rect 1409 4573 1443 4607
rect 1443 4573 1452 4607
rect 1400 4564 1452 4573
rect 1676 4607 1728 4616
rect 1676 4573 1685 4607
rect 1685 4573 1719 4607
rect 1719 4573 1728 4607
rect 1676 4564 1728 4573
rect 5448 4607 5500 4616
rect 5448 4573 5457 4607
rect 5457 4573 5491 4607
rect 5491 4573 5500 4607
rect 5448 4564 5500 4573
rect 6184 4632 6236 4684
rect 9772 4700 9824 4752
rect 6828 4675 6880 4684
rect 6828 4641 6837 4675
rect 6837 4641 6871 4675
rect 6871 4641 6880 4675
rect 6828 4632 6880 4641
rect 7472 4675 7524 4684
rect 7472 4641 7481 4675
rect 7481 4641 7515 4675
rect 7515 4641 7524 4675
rect 7472 4632 7524 4641
rect 7840 4632 7892 4684
rect 10232 4675 10284 4684
rect 10232 4641 10241 4675
rect 10241 4641 10275 4675
rect 10275 4641 10284 4675
rect 10232 4632 10284 4641
rect 10692 4675 10744 4684
rect 10692 4641 10701 4675
rect 10701 4641 10735 4675
rect 10735 4641 10744 4675
rect 10692 4632 10744 4641
rect 10876 4675 10928 4684
rect 10876 4641 10885 4675
rect 10885 4641 10919 4675
rect 10919 4641 10928 4675
rect 10876 4632 10928 4641
rect 12072 4768 12124 4820
rect 14280 4768 14332 4820
rect 18604 4768 18656 4820
rect 22744 4768 22796 4820
rect 11244 4675 11296 4684
rect 11244 4641 11253 4675
rect 11253 4641 11287 4675
rect 11287 4641 11296 4675
rect 11244 4632 11296 4641
rect 11520 4632 11572 4684
rect 12716 4675 12768 4684
rect 12716 4641 12725 4675
rect 12725 4641 12759 4675
rect 12759 4641 12768 4675
rect 12716 4632 12768 4641
rect 14556 4675 14608 4684
rect 14556 4641 14565 4675
rect 14565 4641 14599 4675
rect 14599 4641 14608 4675
rect 14556 4632 14608 4641
rect 15752 4675 15804 4684
rect 15752 4641 15761 4675
rect 15761 4641 15795 4675
rect 15795 4641 15804 4675
rect 15752 4632 15804 4641
rect 15936 4632 15988 4684
rect 16948 4632 17000 4684
rect 17868 4675 17920 4684
rect 9496 4564 9548 4616
rect 14740 4564 14792 4616
rect 17868 4641 17877 4675
rect 17877 4641 17911 4675
rect 17911 4641 17920 4675
rect 17868 4632 17920 4641
rect 18236 4675 18288 4684
rect 18236 4641 18245 4675
rect 18245 4641 18279 4675
rect 18279 4641 18288 4675
rect 18236 4632 18288 4641
rect 18512 4675 18564 4684
rect 18512 4641 18521 4675
rect 18521 4641 18555 4675
rect 18555 4641 18564 4675
rect 18512 4632 18564 4641
rect 10140 4539 10192 4548
rect 10140 4505 10149 4539
rect 10149 4505 10183 4539
rect 10183 4505 10192 4539
rect 10140 4496 10192 4505
rect 13452 4496 13504 4548
rect 18604 4564 18656 4616
rect 20720 4632 20772 4684
rect 20904 4675 20956 4684
rect 20904 4641 20913 4675
rect 20913 4641 20947 4675
rect 20947 4641 20956 4675
rect 20904 4632 20956 4641
rect 16856 4496 16908 4548
rect 18144 4496 18196 4548
rect 18972 4496 19024 4548
rect 19984 4564 20036 4616
rect 22652 4700 22704 4752
rect 22928 4632 22980 4684
rect 23296 4675 23348 4684
rect 23296 4641 23305 4675
rect 23305 4641 23339 4675
rect 23339 4641 23348 4675
rect 23296 4632 23348 4641
rect 24124 4675 24176 4684
rect 24124 4641 24133 4675
rect 24133 4641 24167 4675
rect 24167 4641 24176 4675
rect 24124 4632 24176 4641
rect 30932 4768 30984 4820
rect 31116 4811 31168 4820
rect 31116 4777 31125 4811
rect 31125 4777 31159 4811
rect 31159 4777 31168 4811
rect 31116 4768 31168 4777
rect 31208 4768 31260 4820
rect 32772 4768 32824 4820
rect 32956 4768 33008 4820
rect 25228 4743 25280 4752
rect 25228 4709 25237 4743
rect 25237 4709 25271 4743
rect 25271 4709 25280 4743
rect 25228 4700 25280 4709
rect 25596 4700 25648 4752
rect 24676 4675 24728 4684
rect 24676 4641 24685 4675
rect 24685 4641 24719 4675
rect 24719 4641 24728 4675
rect 24676 4632 24728 4641
rect 25504 4632 25556 4684
rect 26792 4675 26844 4684
rect 26792 4641 26801 4675
rect 26801 4641 26835 4675
rect 26835 4641 26844 4675
rect 26792 4632 26844 4641
rect 28908 4632 28960 4684
rect 30380 4700 30432 4752
rect 32404 4700 32456 4752
rect 33600 4743 33652 4752
rect 25688 4564 25740 4616
rect 28172 4607 28224 4616
rect 19892 4496 19944 4548
rect 20076 4539 20128 4548
rect 20076 4505 20085 4539
rect 20085 4505 20119 4539
rect 20119 4505 20128 4539
rect 20076 4496 20128 4505
rect 22468 4496 22520 4548
rect 22744 4496 22796 4548
rect 28172 4573 28181 4607
rect 28181 4573 28215 4607
rect 28215 4573 28224 4607
rect 28172 4564 28224 4573
rect 29828 4564 29880 4616
rect 30840 4632 30892 4684
rect 30932 4675 30984 4684
rect 30932 4641 30941 4675
rect 30941 4641 30975 4675
rect 30975 4641 30984 4675
rect 32680 4675 32732 4684
rect 30932 4632 30984 4641
rect 32680 4641 32689 4675
rect 32689 4641 32723 4675
rect 32723 4641 32732 4675
rect 32680 4632 32732 4641
rect 33600 4709 33609 4743
rect 33609 4709 33643 4743
rect 33643 4709 33652 4743
rect 33600 4700 33652 4709
rect 33876 4700 33928 4752
rect 30656 4564 30708 4616
rect 4620 4428 4672 4480
rect 13820 4471 13872 4480
rect 13820 4437 13829 4471
rect 13829 4437 13863 4471
rect 13863 4437 13872 4471
rect 13820 4428 13872 4437
rect 15936 4471 15988 4480
rect 15936 4437 15945 4471
rect 15945 4437 15979 4471
rect 15979 4437 15988 4471
rect 15936 4428 15988 4437
rect 19340 4428 19392 4480
rect 22560 4428 22612 4480
rect 23664 4428 23716 4480
rect 31024 4564 31076 4616
rect 33876 4564 33928 4616
rect 34612 4675 34664 4684
rect 34612 4641 34621 4675
rect 34621 4641 34655 4675
rect 34655 4641 34664 4675
rect 34612 4632 34664 4641
rect 35440 4632 35492 4684
rect 37280 4700 37332 4752
rect 36544 4675 36596 4684
rect 36544 4641 36553 4675
rect 36553 4641 36587 4675
rect 36587 4641 36596 4675
rect 36544 4632 36596 4641
rect 37740 4675 37792 4684
rect 37740 4641 37749 4675
rect 37749 4641 37783 4675
rect 37783 4641 37792 4675
rect 37740 4632 37792 4641
rect 32404 4496 32456 4548
rect 34520 4564 34572 4616
rect 35532 4564 35584 4616
rect 34428 4496 34480 4548
rect 33968 4428 34020 4480
rect 35440 4428 35492 4480
rect 37004 4428 37056 4480
rect 37924 4471 37976 4480
rect 37924 4437 37933 4471
rect 37933 4437 37967 4471
rect 37967 4437 37976 4471
rect 37924 4428 37976 4437
rect 4246 4326 4298 4378
rect 4310 4326 4362 4378
rect 4374 4326 4426 4378
rect 4438 4326 4490 4378
rect 34966 4326 35018 4378
rect 35030 4326 35082 4378
rect 35094 4326 35146 4378
rect 35158 4326 35210 4378
rect 7012 4224 7064 4276
rect 11244 4224 11296 4276
rect 19432 4267 19484 4276
rect 9496 4199 9548 4208
rect 9496 4165 9505 4199
rect 9505 4165 9539 4199
rect 9539 4165 9548 4199
rect 9496 4156 9548 4165
rect 10692 4156 10744 4208
rect 3240 4131 3292 4140
rect 3240 4097 3249 4131
rect 3249 4097 3283 4131
rect 3283 4097 3292 4131
rect 3240 4088 3292 4097
rect 1860 4020 1912 4072
rect 2964 4063 3016 4072
rect 1676 3884 1728 3936
rect 2964 4029 2973 4063
rect 2973 4029 3007 4063
rect 3007 4029 3016 4063
rect 2964 4020 3016 4029
rect 4620 4088 4672 4140
rect 7196 4088 7248 4140
rect 3976 3952 4028 4004
rect 6920 4020 6972 4072
rect 7840 4020 7892 4072
rect 10232 4088 10284 4140
rect 9864 4063 9916 4072
rect 9864 4029 9873 4063
rect 9873 4029 9907 4063
rect 9907 4029 9916 4063
rect 9864 4020 9916 4029
rect 10876 4088 10928 4140
rect 10508 4020 10560 4072
rect 11520 4088 11572 4140
rect 13820 4156 13872 4208
rect 19432 4233 19441 4267
rect 19441 4233 19475 4267
rect 19475 4233 19484 4267
rect 19432 4224 19484 4233
rect 21548 4267 21600 4276
rect 21548 4233 21557 4267
rect 21557 4233 21591 4267
rect 21591 4233 21600 4267
rect 21548 4224 21600 4233
rect 26240 4224 26292 4276
rect 31024 4224 31076 4276
rect 32220 4224 32272 4276
rect 19340 4156 19392 4208
rect 22100 4156 22152 4208
rect 30656 4199 30708 4208
rect 15016 4131 15068 4140
rect 11428 4020 11480 4072
rect 15016 4097 15025 4131
rect 15025 4097 15059 4131
rect 15059 4097 15068 4131
rect 15016 4088 15068 4097
rect 15476 4088 15528 4140
rect 20076 4088 20128 4140
rect 30656 4165 30665 4199
rect 30665 4165 30699 4199
rect 30699 4165 30708 4199
rect 30656 4156 30708 4165
rect 24860 4131 24912 4140
rect 24860 4097 24869 4131
rect 24869 4097 24903 4131
rect 24903 4097 24912 4131
rect 24860 4088 24912 4097
rect 14004 4020 14056 4072
rect 14740 4063 14792 4072
rect 14740 4029 14749 4063
rect 14749 4029 14783 4063
rect 14783 4029 14792 4063
rect 14740 4020 14792 4029
rect 16948 4063 17000 4072
rect 16948 4029 16957 4063
rect 16957 4029 16991 4063
rect 16991 4029 17000 4063
rect 16948 4020 17000 4029
rect 17040 4063 17092 4072
rect 17040 4029 17049 4063
rect 17049 4029 17083 4063
rect 17083 4029 17092 4063
rect 18052 4063 18104 4072
rect 17040 4020 17092 4029
rect 18052 4029 18061 4063
rect 18061 4029 18095 4063
rect 18095 4029 18104 4063
rect 18052 4020 18104 4029
rect 20168 4063 20220 4072
rect 20168 4029 20177 4063
rect 20177 4029 20211 4063
rect 20211 4029 20220 4063
rect 20168 4020 20220 4029
rect 20444 4063 20496 4072
rect 20444 4029 20453 4063
rect 20453 4029 20487 4063
rect 20487 4029 20496 4063
rect 20444 4020 20496 4029
rect 22100 4020 22152 4072
rect 22376 4063 22428 4072
rect 22376 4029 22385 4063
rect 22385 4029 22419 4063
rect 22419 4029 22428 4063
rect 22376 4020 22428 4029
rect 22560 4020 22612 4072
rect 24584 4020 24636 4072
rect 25780 4020 25832 4072
rect 26884 4020 26936 4072
rect 28448 4020 28500 4072
rect 29092 4088 29144 4140
rect 29184 4088 29236 4140
rect 30288 4088 30340 4140
rect 32404 4088 32456 4140
rect 32680 4131 32732 4140
rect 32680 4097 32689 4131
rect 32689 4097 32723 4131
rect 32723 4097 32732 4131
rect 32680 4088 32732 4097
rect 33968 4156 34020 4208
rect 37280 4224 37332 4276
rect 34336 4088 34388 4140
rect 4804 3884 4856 3936
rect 5172 3927 5224 3936
rect 5172 3893 5181 3927
rect 5181 3893 5215 3927
rect 5215 3893 5224 3927
rect 5172 3884 5224 3893
rect 7380 3884 7432 3936
rect 14188 3952 14240 4004
rect 12624 3884 12676 3936
rect 16028 3884 16080 3936
rect 19064 3952 19116 4004
rect 20076 3952 20128 4004
rect 24124 3952 24176 4004
rect 24860 3952 24912 4004
rect 26516 3995 26568 4004
rect 26516 3961 26525 3995
rect 26525 3961 26559 3995
rect 26559 3961 26568 3995
rect 26516 3952 26568 3961
rect 28080 3952 28132 4004
rect 19248 3884 19300 3936
rect 19432 3884 19484 3936
rect 22008 3884 22060 3936
rect 29368 4020 29420 4072
rect 29552 4063 29604 4072
rect 29552 4029 29561 4063
rect 29561 4029 29595 4063
rect 29595 4029 29604 4063
rect 29552 4020 29604 4029
rect 34244 4020 34296 4072
rect 35716 4088 35768 4140
rect 35900 4020 35952 4072
rect 36084 4063 36136 4072
rect 36084 4029 36093 4063
rect 36093 4029 36127 4063
rect 36127 4029 36136 4063
rect 36084 4020 36136 4029
rect 30196 3884 30248 3936
rect 35440 3952 35492 4004
rect 35624 3952 35676 4004
rect 33876 3884 33928 3936
rect 34612 3884 34664 3936
rect 19606 3782 19658 3834
rect 19670 3782 19722 3834
rect 19734 3782 19786 3834
rect 19798 3782 19850 3834
rect 2964 3680 3016 3732
rect 6552 3723 6604 3732
rect 5172 3612 5224 3664
rect 1400 3476 1452 3528
rect 2596 3476 2648 3528
rect 3424 3476 3476 3528
rect 4068 3476 4120 3528
rect 4712 3519 4764 3528
rect 4712 3485 4721 3519
rect 4721 3485 4755 3519
rect 4755 3485 4764 3519
rect 4712 3476 4764 3485
rect 6552 3689 6561 3723
rect 6561 3689 6595 3723
rect 6595 3689 6604 3723
rect 6552 3680 6604 3689
rect 5448 3587 5500 3596
rect 5448 3553 5457 3587
rect 5457 3553 5491 3587
rect 5491 3553 5500 3587
rect 5448 3544 5500 3553
rect 5816 3544 5868 3596
rect 7472 3587 7524 3596
rect 7472 3553 7481 3587
rect 7481 3553 7515 3587
rect 7515 3553 7524 3587
rect 7472 3544 7524 3553
rect 8668 3587 8720 3596
rect 8668 3553 8677 3587
rect 8677 3553 8711 3587
rect 8711 3553 8720 3587
rect 8668 3544 8720 3553
rect 9772 3612 9824 3664
rect 12624 3680 12676 3732
rect 13452 3680 13504 3732
rect 14832 3680 14884 3732
rect 16028 3680 16080 3732
rect 25596 3680 25648 3732
rect 25780 3723 25832 3732
rect 25780 3689 25789 3723
rect 25789 3689 25823 3723
rect 25823 3689 25832 3723
rect 25780 3680 25832 3689
rect 19340 3612 19392 3664
rect 12256 3544 12308 3596
rect 12808 3587 12860 3596
rect 6920 3476 6972 3528
rect 7380 3519 7432 3528
rect 7380 3485 7389 3519
rect 7389 3485 7423 3519
rect 7423 3485 7432 3519
rect 7380 3476 7432 3485
rect 7932 3519 7984 3528
rect 7932 3485 7941 3519
rect 7941 3485 7975 3519
rect 7975 3485 7984 3519
rect 7932 3476 7984 3485
rect 9312 3476 9364 3528
rect 6828 3408 6880 3460
rect 12440 3476 12492 3528
rect 12808 3553 12817 3587
rect 12817 3553 12851 3587
rect 12851 3553 12860 3587
rect 12808 3544 12860 3553
rect 15292 3587 15344 3596
rect 15292 3553 15301 3587
rect 15301 3553 15335 3587
rect 15335 3553 15344 3587
rect 15292 3544 15344 3553
rect 15568 3544 15620 3596
rect 15844 3587 15896 3596
rect 15844 3553 15853 3587
rect 15853 3553 15887 3587
rect 15887 3553 15896 3587
rect 15844 3544 15896 3553
rect 16856 3587 16908 3596
rect 16856 3553 16865 3587
rect 16865 3553 16899 3587
rect 16899 3553 16908 3587
rect 16856 3544 16908 3553
rect 16948 3544 17000 3596
rect 19432 3544 19484 3596
rect 20444 3612 20496 3664
rect 21548 3612 21600 3664
rect 12348 3408 12400 3460
rect 14740 3476 14792 3528
rect 19892 3476 19944 3528
rect 21272 3587 21324 3596
rect 21272 3553 21281 3587
rect 21281 3553 21315 3587
rect 21315 3553 21324 3587
rect 21640 3587 21692 3596
rect 21272 3544 21324 3553
rect 21640 3553 21649 3587
rect 21649 3553 21683 3587
rect 21683 3553 21692 3587
rect 21640 3544 21692 3553
rect 22744 3587 22796 3596
rect 22744 3553 22753 3587
rect 22753 3553 22787 3587
rect 22787 3553 22796 3587
rect 22744 3544 22796 3553
rect 24032 3612 24084 3664
rect 27252 3680 27304 3732
rect 28448 3680 28500 3732
rect 23020 3544 23072 3596
rect 24676 3544 24728 3596
rect 29368 3612 29420 3664
rect 30196 3680 30248 3732
rect 24584 3519 24636 3528
rect 24584 3485 24593 3519
rect 24593 3485 24627 3519
rect 24627 3485 24636 3519
rect 24584 3476 24636 3485
rect 26516 3587 26568 3596
rect 26516 3553 26525 3587
rect 26525 3553 26559 3587
rect 26559 3553 26568 3587
rect 26516 3544 26568 3553
rect 27160 3587 27212 3596
rect 27160 3553 27169 3587
rect 27169 3553 27203 3587
rect 27203 3553 27212 3587
rect 27160 3544 27212 3553
rect 28080 3587 28132 3596
rect 28080 3553 28089 3587
rect 28089 3553 28123 3587
rect 28123 3553 28132 3587
rect 28080 3544 28132 3553
rect 29184 3476 29236 3528
rect 34520 3612 34572 3664
rect 37280 3680 37332 3732
rect 37464 3612 37516 3664
rect 30380 3544 30432 3596
rect 33324 3544 33376 3596
rect 37556 3544 37608 3596
rect 31760 3476 31812 3528
rect 32128 3476 32180 3528
rect 32772 3519 32824 3528
rect 32772 3485 32781 3519
rect 32781 3485 32815 3519
rect 32815 3485 32824 3519
rect 32772 3476 32824 3485
rect 34428 3476 34480 3528
rect 34704 3476 34756 3528
rect 36084 3476 36136 3528
rect 17960 3451 18012 3460
rect 17960 3417 17969 3451
rect 17969 3417 18003 3451
rect 18003 3417 18012 3451
rect 17960 3408 18012 3417
rect 18052 3408 18104 3460
rect 20168 3408 20220 3460
rect 22836 3408 22888 3460
rect 14464 3340 14516 3392
rect 14924 3340 14976 3392
rect 20260 3340 20312 3392
rect 23940 3383 23992 3392
rect 23940 3349 23949 3383
rect 23949 3349 23983 3383
rect 23983 3349 23992 3383
rect 23940 3340 23992 3349
rect 25688 3340 25740 3392
rect 34796 3408 34848 3460
rect 4246 3238 4298 3290
rect 4310 3238 4362 3290
rect 4374 3238 4426 3290
rect 4438 3238 4490 3290
rect 34966 3238 35018 3290
rect 35030 3238 35082 3290
rect 35094 3238 35146 3290
rect 35158 3238 35210 3290
rect 3792 3136 3844 3188
rect 4068 3136 4120 3188
rect 7472 3136 7524 3188
rect 8668 3136 8720 3188
rect 11428 3179 11480 3188
rect 7840 3068 7892 3120
rect 11428 3145 11437 3179
rect 11437 3145 11471 3179
rect 11471 3145 11480 3179
rect 11428 3136 11480 3145
rect 14004 3179 14056 3188
rect 14004 3145 14013 3179
rect 14013 3145 14047 3179
rect 14047 3145 14056 3179
rect 14004 3136 14056 3145
rect 15752 3136 15804 3188
rect 17040 3136 17092 3188
rect 20168 3136 20220 3188
rect 12256 3068 12308 3120
rect 22560 3068 22612 3120
rect 23020 3111 23072 3120
rect 23020 3077 23029 3111
rect 23029 3077 23063 3111
rect 23063 3077 23072 3111
rect 23020 3068 23072 3077
rect 2872 3043 2924 3052
rect 2872 3009 2881 3043
rect 2881 3009 2915 3043
rect 2915 3009 2924 3043
rect 2872 3000 2924 3009
rect 7564 3000 7616 3052
rect 2596 2975 2648 2984
rect 2596 2941 2605 2975
rect 2605 2941 2639 2975
rect 2639 2941 2648 2975
rect 2596 2932 2648 2941
rect 5724 2932 5776 2984
rect 4620 2864 4672 2916
rect 4804 2796 4856 2848
rect 6644 2932 6696 2984
rect 6828 2975 6880 2984
rect 6828 2941 6837 2975
rect 6837 2941 6871 2975
rect 6871 2941 6880 2975
rect 6828 2932 6880 2941
rect 7104 2975 7156 2984
rect 7104 2941 7113 2975
rect 7113 2941 7147 2975
rect 7147 2941 7156 2975
rect 7104 2932 7156 2941
rect 7196 2932 7248 2984
rect 10048 3000 10100 3052
rect 12348 3000 12400 3052
rect 14832 3043 14884 3052
rect 9036 2975 9088 2984
rect 9036 2941 9045 2975
rect 9045 2941 9079 2975
rect 9079 2941 9088 2975
rect 9036 2932 9088 2941
rect 10140 2975 10192 2984
rect 10140 2941 10149 2975
rect 10149 2941 10183 2975
rect 10183 2941 10192 2975
rect 10140 2932 10192 2941
rect 12532 2932 12584 2984
rect 14832 3009 14841 3043
rect 14841 3009 14875 3043
rect 14875 3009 14884 3043
rect 14832 3000 14884 3009
rect 15292 3000 15344 3052
rect 16488 3000 16540 3052
rect 16856 3000 16908 3052
rect 22836 3000 22888 3052
rect 25596 3136 25648 3188
rect 17316 2975 17368 2984
rect 17316 2941 17325 2975
rect 17325 2941 17359 2975
rect 17359 2941 17368 2975
rect 17316 2932 17368 2941
rect 7196 2796 7248 2848
rect 7472 2796 7524 2848
rect 15660 2864 15712 2916
rect 18328 2975 18380 2984
rect 18328 2941 18337 2975
rect 18337 2941 18371 2975
rect 18371 2941 18380 2975
rect 18328 2932 18380 2941
rect 20628 2975 20680 2984
rect 20628 2941 20637 2975
rect 20637 2941 20671 2975
rect 20671 2941 20680 2975
rect 20628 2932 20680 2941
rect 20904 2975 20956 2984
rect 20904 2941 20913 2975
rect 20913 2941 20947 2975
rect 20947 2941 20956 2975
rect 20904 2932 20956 2941
rect 23940 3043 23992 3052
rect 23940 3009 23949 3043
rect 23949 3009 23983 3043
rect 23983 3009 23992 3043
rect 23940 3000 23992 3009
rect 25872 3000 25924 3052
rect 26884 3000 26936 3052
rect 29552 3000 29604 3052
rect 29828 3043 29880 3052
rect 29828 3009 29837 3043
rect 29837 3009 29871 3043
rect 29871 3009 29880 3043
rect 29828 3000 29880 3009
rect 26240 2975 26292 2984
rect 26240 2941 26249 2975
rect 26249 2941 26283 2975
rect 26283 2941 26292 2975
rect 26240 2932 26292 2941
rect 27896 2932 27948 2984
rect 29092 2932 29144 2984
rect 32220 3068 32272 3120
rect 33232 3000 33284 3052
rect 17960 2864 18012 2916
rect 27528 2864 27580 2916
rect 10600 2796 10652 2848
rect 18696 2796 18748 2848
rect 23020 2796 23072 2848
rect 30380 2932 30432 2984
rect 34336 3043 34388 3052
rect 34336 3009 34345 3043
rect 34345 3009 34379 3043
rect 34379 3009 34388 3043
rect 34336 3000 34388 3009
rect 35440 3043 35492 3052
rect 35440 3009 35449 3043
rect 35449 3009 35483 3043
rect 35483 3009 35492 3043
rect 35440 3000 35492 3009
rect 33876 2975 33928 2984
rect 33876 2941 33885 2975
rect 33885 2941 33919 2975
rect 33919 2941 33928 2975
rect 33876 2932 33928 2941
rect 34152 2975 34204 2984
rect 34152 2941 34161 2975
rect 34161 2941 34195 2975
rect 34195 2941 34204 2975
rect 34152 2932 34204 2941
rect 34520 2932 34572 2984
rect 36452 2975 36504 2984
rect 32220 2864 32272 2916
rect 36452 2941 36461 2975
rect 36461 2941 36495 2975
rect 36495 2941 36504 2975
rect 36452 2932 36504 2941
rect 36268 2864 36320 2916
rect 38108 2907 38160 2916
rect 38108 2873 38117 2907
rect 38117 2873 38151 2907
rect 38151 2873 38160 2907
rect 38108 2864 38160 2873
rect 32128 2796 32180 2848
rect 32680 2796 32732 2848
rect 32772 2796 32824 2848
rect 34704 2796 34756 2848
rect 19606 2694 19658 2746
rect 19670 2694 19722 2746
rect 19734 2694 19786 2746
rect 19798 2694 19850 2746
rect 6644 2592 6696 2644
rect 9864 2635 9916 2644
rect 7472 2524 7524 2576
rect 9864 2601 9873 2635
rect 9873 2601 9907 2635
rect 9907 2601 9916 2635
rect 9864 2592 9916 2601
rect 1952 2456 2004 2508
rect 2596 2456 2648 2508
rect 4712 2456 4764 2508
rect 6920 2499 6972 2508
rect 6920 2465 6929 2499
rect 6929 2465 6963 2499
rect 6963 2465 6972 2499
rect 6920 2456 6972 2465
rect 7564 2499 7616 2508
rect 7564 2465 7573 2499
rect 7573 2465 7607 2499
rect 7607 2465 7616 2499
rect 7564 2456 7616 2465
rect 12900 2524 12952 2576
rect 9680 2456 9732 2508
rect 9312 2388 9364 2440
rect 2596 2252 2648 2304
rect 7656 2252 7708 2304
rect 12440 2456 12492 2508
rect 14464 2499 14516 2508
rect 14464 2465 14473 2499
rect 14473 2465 14507 2499
rect 14507 2465 14516 2499
rect 14464 2456 14516 2465
rect 17960 2524 18012 2576
rect 22376 2592 22428 2644
rect 26240 2592 26292 2644
rect 36268 2592 36320 2644
rect 37924 2592 37976 2644
rect 32036 2567 32088 2576
rect 15476 2456 15528 2508
rect 15660 2499 15712 2508
rect 15660 2465 15669 2499
rect 15669 2465 15703 2499
rect 15703 2465 15712 2499
rect 15660 2456 15712 2465
rect 15936 2499 15988 2508
rect 15936 2465 15945 2499
rect 15945 2465 15979 2499
rect 15979 2465 15988 2499
rect 15936 2456 15988 2465
rect 32036 2533 32045 2567
rect 32045 2533 32079 2567
rect 32079 2533 32088 2567
rect 32036 2524 32088 2533
rect 34428 2524 34480 2576
rect 12624 2431 12676 2440
rect 12624 2397 12633 2431
rect 12633 2397 12667 2431
rect 12667 2397 12676 2431
rect 12624 2388 12676 2397
rect 14188 2388 14240 2440
rect 15568 2320 15620 2372
rect 24124 2456 24176 2508
rect 24860 2499 24912 2508
rect 18880 2388 18932 2440
rect 19248 2431 19300 2440
rect 19248 2397 19257 2431
rect 19257 2397 19291 2431
rect 19291 2397 19300 2431
rect 19248 2388 19300 2397
rect 20628 2388 20680 2440
rect 21364 2388 21416 2440
rect 24860 2465 24869 2499
rect 24869 2465 24903 2499
rect 24903 2465 24912 2499
rect 24860 2456 24912 2465
rect 26884 2431 26936 2440
rect 26884 2397 26893 2431
rect 26893 2397 26927 2431
rect 26927 2397 26936 2431
rect 26884 2388 26936 2397
rect 29276 2388 29328 2440
rect 30288 2456 30340 2508
rect 32220 2456 32272 2508
rect 33140 2456 33192 2508
rect 35532 2456 35584 2508
rect 37464 2456 37516 2508
rect 36360 2388 36412 2440
rect 16948 2252 17000 2304
rect 17868 2252 17920 2304
rect 20352 2252 20404 2304
rect 20996 2252 21048 2304
rect 27252 2252 27304 2304
rect 31300 2252 31352 2304
rect 33140 2295 33192 2304
rect 33140 2261 33149 2295
rect 33149 2261 33183 2295
rect 33183 2261 33192 2295
rect 33140 2252 33192 2261
rect 35348 2252 35400 2304
rect 37556 2295 37608 2304
rect 37556 2261 37565 2295
rect 37565 2261 37599 2295
rect 37599 2261 37608 2295
rect 37556 2252 37608 2261
rect 4246 2150 4298 2202
rect 4310 2150 4362 2202
rect 4374 2150 4426 2202
rect 4438 2150 4490 2202
rect 34966 2150 35018 2202
rect 35030 2150 35082 2202
rect 35094 2150 35146 2202
rect 35158 2150 35210 2202
rect 7932 2048 7984 2100
rect 33140 2048 33192 2100
rect 6920 1980 6972 2032
rect 8668 1980 8720 2032
rect 18880 1980 18932 2032
rect 20628 1980 20680 2032
rect 20076 1912 20128 1964
rect 25228 1912 25280 1964
<< metal2 >>
rect 1306 39200 1362 40000
rect 3330 39200 3386 40000
rect 5354 39200 5410 40000
rect 7378 39200 7434 40000
rect 9402 39200 9458 40000
rect 11610 39200 11666 40000
rect 13634 39200 13690 40000
rect 15658 39200 15714 40000
rect 17682 39200 17738 40000
rect 19706 39200 19762 40000
rect 21914 39200 21970 40000
rect 23938 39200 23994 40000
rect 25962 39200 26018 40000
rect 27986 39200 28042 40000
rect 30010 39200 30066 40000
rect 32034 39200 32090 40000
rect 34242 39200 34298 40000
rect 36266 39200 36322 40000
rect 38290 39200 38346 40000
rect 1320 37194 1348 39200
rect 2778 37360 2834 37369
rect 2778 37295 2834 37304
rect 1308 37188 1360 37194
rect 1308 37130 1360 37136
rect 2792 36922 2820 37295
rect 2780 36916 2832 36922
rect 2780 36858 2832 36864
rect 2504 36848 2556 36854
rect 2504 36790 2556 36796
rect 3344 36802 3372 39200
rect 4712 37324 4764 37330
rect 4712 37266 4764 37272
rect 4220 37020 4516 37040
rect 4276 37018 4300 37020
rect 4356 37018 4380 37020
rect 4436 37018 4460 37020
rect 4298 36966 4300 37018
rect 4362 36966 4374 37018
rect 4436 36966 4438 37018
rect 4276 36964 4300 36966
rect 4356 36964 4380 36966
rect 4436 36964 4460 36966
rect 4220 36944 4516 36964
rect 2516 36718 2544 36790
rect 3344 36774 3464 36802
rect 2504 36712 2556 36718
rect 2504 36654 2556 36660
rect 3332 36712 3384 36718
rect 3332 36654 3384 36660
rect 1952 36576 2004 36582
rect 1952 36518 2004 36524
rect 1676 34944 1728 34950
rect 1676 34886 1728 34892
rect 1584 34468 1636 34474
rect 1584 34410 1636 34416
rect 1400 33992 1452 33998
rect 1400 33934 1452 33940
rect 1412 33522 1440 33934
rect 1400 33516 1452 33522
rect 1400 33458 1452 33464
rect 1492 33448 1544 33454
rect 1492 33390 1544 33396
rect 1504 33046 1532 33390
rect 1596 33386 1624 34410
rect 1688 33454 1716 34886
rect 1860 33992 1912 33998
rect 1860 33934 1912 33940
rect 1872 33658 1900 33934
rect 1860 33652 1912 33658
rect 1860 33594 1912 33600
rect 1676 33448 1728 33454
rect 1676 33390 1728 33396
rect 1584 33380 1636 33386
rect 1584 33322 1636 33328
rect 1492 33040 1544 33046
rect 1492 32982 1544 32988
rect 1860 32360 1912 32366
rect 1860 32302 1912 32308
rect 1676 32224 1728 32230
rect 1676 32166 1728 32172
rect 1688 31890 1716 32166
rect 1676 31884 1728 31890
rect 1676 31826 1728 31832
rect 1400 31816 1452 31822
rect 1400 31758 1452 31764
rect 1412 30190 1440 31758
rect 1872 30802 1900 32302
rect 1964 31113 1992 36518
rect 2688 36236 2740 36242
rect 2688 36178 2740 36184
rect 2228 35624 2280 35630
rect 2228 35566 2280 35572
rect 2240 35290 2268 35566
rect 2228 35284 2280 35290
rect 2228 35226 2280 35232
rect 2700 35086 2728 36178
rect 3344 36174 3372 36654
rect 2872 36168 2924 36174
rect 2872 36110 2924 36116
rect 3332 36168 3384 36174
rect 3332 36110 3384 36116
rect 2884 35154 2912 36110
rect 3056 36100 3108 36106
rect 3056 36042 3108 36048
rect 3068 35222 3096 36042
rect 3436 35290 3464 36774
rect 3976 36712 4028 36718
rect 3976 36654 4028 36660
rect 3988 36378 4016 36654
rect 3976 36372 4028 36378
rect 3976 36314 4028 36320
rect 3988 35698 4016 36314
rect 4220 35932 4516 35952
rect 4276 35930 4300 35932
rect 4356 35930 4380 35932
rect 4436 35930 4460 35932
rect 4298 35878 4300 35930
rect 4362 35878 4374 35930
rect 4436 35878 4438 35930
rect 4276 35876 4300 35878
rect 4356 35876 4380 35878
rect 4436 35876 4460 35878
rect 4220 35856 4516 35876
rect 3976 35692 4028 35698
rect 3976 35634 4028 35640
rect 3424 35284 3476 35290
rect 3424 35226 3476 35232
rect 3056 35216 3108 35222
rect 3056 35158 3108 35164
rect 2872 35148 2924 35154
rect 2872 35090 2924 35096
rect 2688 35080 2740 35086
rect 2688 35022 2740 35028
rect 2700 34950 2728 35022
rect 2688 34944 2740 34950
rect 2688 34886 2740 34892
rect 3792 34944 3844 34950
rect 3792 34886 3844 34892
rect 2228 34740 2280 34746
rect 2228 34682 2280 34688
rect 2240 34542 2268 34682
rect 3804 34542 3832 34886
rect 2228 34536 2280 34542
rect 2228 34478 2280 34484
rect 2688 34536 2740 34542
rect 2688 34478 2740 34484
rect 3240 34536 3292 34542
rect 3240 34478 3292 34484
rect 3608 34536 3660 34542
rect 3608 34478 3660 34484
rect 3792 34536 3844 34542
rect 3792 34478 3844 34484
rect 2700 34202 2728 34478
rect 2688 34196 2740 34202
rect 2688 34138 2740 34144
rect 2700 33810 2728 34138
rect 2608 33782 2728 33810
rect 2608 32978 2636 33782
rect 3252 32978 3280 34478
rect 3620 32978 3648 34478
rect 3790 34096 3846 34105
rect 3790 34031 3846 34040
rect 2596 32972 2648 32978
rect 2596 32914 2648 32920
rect 2780 32972 2832 32978
rect 2780 32914 2832 32920
rect 2964 32972 3016 32978
rect 2964 32914 3016 32920
rect 3148 32972 3200 32978
rect 3148 32914 3200 32920
rect 3240 32972 3292 32978
rect 3240 32914 3292 32920
rect 3608 32972 3660 32978
rect 3608 32914 3660 32920
rect 2228 32360 2280 32366
rect 2228 32302 2280 32308
rect 2240 31346 2268 32302
rect 2792 31346 2820 32914
rect 2976 32502 3004 32914
rect 2964 32496 3016 32502
rect 2964 32438 3016 32444
rect 2872 32360 2924 32366
rect 2872 32302 2924 32308
rect 2884 31414 2912 32302
rect 2872 31408 2924 31414
rect 2872 31350 2924 31356
rect 2228 31340 2280 31346
rect 2228 31282 2280 31288
rect 2780 31340 2832 31346
rect 2780 31282 2832 31288
rect 2136 31272 2188 31278
rect 2134 31240 2136 31249
rect 3160 31249 3188 32914
rect 3252 31958 3280 32914
rect 3240 31952 3292 31958
rect 3240 31894 3292 31900
rect 3252 31278 3280 31894
rect 3516 31476 3568 31482
rect 3516 31418 3568 31424
rect 3332 31340 3384 31346
rect 3332 31282 3384 31288
rect 3240 31272 3292 31278
rect 2188 31240 2190 31249
rect 2134 31175 2190 31184
rect 3146 31240 3202 31249
rect 3240 31214 3292 31220
rect 3146 31175 3202 31184
rect 1950 31104 2006 31113
rect 1950 31039 2006 31048
rect 1860 30796 1912 30802
rect 1860 30738 1912 30744
rect 2964 30796 3016 30802
rect 2964 30738 3016 30744
rect 1400 30184 1452 30190
rect 1400 30126 1452 30132
rect 2872 30048 2924 30054
rect 2872 29990 2924 29996
rect 2884 29714 2912 29990
rect 2872 29708 2924 29714
rect 2872 29650 2924 29656
rect 2976 29594 3004 30738
rect 3148 30660 3200 30666
rect 3148 30602 3200 30608
rect 3160 30258 3188 30602
rect 3148 30252 3200 30258
rect 3148 30194 3200 30200
rect 2884 29566 3004 29594
rect 2780 29096 2832 29102
rect 2780 29038 2832 29044
rect 1400 28552 1452 28558
rect 1400 28494 1452 28500
rect 1860 28552 1912 28558
rect 1860 28494 1912 28500
rect 1412 26450 1440 28494
rect 1872 28218 1900 28494
rect 2412 28484 2464 28490
rect 2412 28426 2464 28432
rect 1860 28212 1912 28218
rect 1860 28154 1912 28160
rect 2424 28014 2452 28426
rect 2792 28014 2820 29038
rect 2884 28966 2912 29566
rect 2964 29504 3016 29510
rect 2964 29446 3016 29452
rect 2976 29102 3004 29446
rect 2964 29096 3016 29102
rect 2964 29038 3016 29044
rect 3240 29096 3292 29102
rect 3240 29038 3292 29044
rect 2872 28960 2924 28966
rect 2872 28902 2924 28908
rect 2964 28960 3016 28966
rect 2964 28902 3016 28908
rect 2976 28422 3004 28902
rect 2964 28416 3016 28422
rect 2964 28358 3016 28364
rect 2976 28082 3004 28358
rect 3054 28112 3110 28121
rect 2964 28076 3016 28082
rect 3054 28047 3110 28056
rect 2964 28018 3016 28024
rect 2412 28008 2464 28014
rect 2412 27950 2464 27956
rect 2780 28008 2832 28014
rect 2780 27950 2832 27956
rect 2688 27532 2740 27538
rect 2688 27474 2740 27480
rect 1492 27464 1544 27470
rect 1492 27406 1544 27412
rect 1504 27130 1532 27406
rect 1492 27124 1544 27130
rect 1492 27066 1544 27072
rect 1676 27124 1728 27130
rect 1676 27066 1728 27072
rect 1688 26450 1716 27066
rect 1768 26920 1820 26926
rect 1768 26862 1820 26868
rect 2700 26908 2728 27474
rect 2780 26920 2832 26926
rect 2700 26880 2780 26908
rect 1400 26444 1452 26450
rect 1400 26386 1452 26392
rect 1676 26444 1728 26450
rect 1676 26386 1728 26392
rect 1412 25362 1440 26386
rect 1780 25906 1808 26862
rect 2700 26314 2728 26880
rect 2780 26862 2832 26868
rect 2688 26308 2740 26314
rect 2688 26250 2740 26256
rect 1860 25968 1912 25974
rect 1860 25910 1912 25916
rect 1768 25900 1820 25906
rect 1768 25842 1820 25848
rect 1400 25356 1452 25362
rect 1400 25298 1452 25304
rect 1676 25288 1728 25294
rect 1676 25230 1728 25236
rect 1688 23730 1716 25230
rect 1872 24750 1900 25910
rect 2700 25838 2728 26250
rect 2688 25832 2740 25838
rect 2688 25774 2740 25780
rect 2688 25356 2740 25362
rect 2688 25298 2740 25304
rect 2700 24750 2728 25298
rect 1860 24744 1912 24750
rect 1860 24686 1912 24692
rect 2688 24744 2740 24750
rect 2688 24686 2740 24692
rect 1676 23724 1728 23730
rect 1676 23666 1728 23672
rect 1400 23044 1452 23050
rect 1400 22986 1452 22992
rect 1412 22642 1440 22986
rect 1676 22976 1728 22982
rect 1676 22918 1728 22924
rect 1688 22642 1716 22918
rect 1400 22636 1452 22642
rect 1400 22578 1452 22584
rect 1676 22636 1728 22642
rect 1676 22578 1728 22584
rect 1768 22092 1820 22098
rect 1768 22034 1820 22040
rect 1780 21622 1808 22034
rect 1872 21706 1900 24686
rect 2228 24268 2280 24274
rect 2228 24210 2280 24216
rect 2872 24268 2924 24274
rect 2872 24210 2924 24216
rect 1872 21678 1992 21706
rect 1768 21616 1820 21622
rect 1768 21558 1820 21564
rect 1860 21548 1912 21554
rect 1860 21490 1912 21496
rect 1492 21480 1544 21486
rect 1492 21422 1544 21428
rect 1504 20874 1532 21422
rect 1584 21344 1636 21350
rect 1584 21286 1636 21292
rect 1492 20868 1544 20874
rect 1492 20810 1544 20816
rect 1596 20466 1624 21286
rect 1872 21010 1900 21490
rect 1860 21004 1912 21010
rect 1860 20946 1912 20952
rect 1584 20460 1636 20466
rect 1584 20402 1636 20408
rect 1400 20392 1452 20398
rect 1400 20334 1452 20340
rect 1412 19310 1440 20334
rect 1964 19922 1992 21678
rect 1952 19916 2004 19922
rect 1952 19858 2004 19864
rect 1400 19304 1452 19310
rect 1400 19246 1452 19252
rect 1412 18222 1440 19246
rect 1400 18216 1452 18222
rect 1400 18158 1452 18164
rect 1412 17678 1440 18158
rect 1400 17672 1452 17678
rect 1400 17614 1452 17620
rect 2136 17672 2188 17678
rect 2136 17614 2188 17620
rect 1412 16590 1440 17614
rect 2148 17338 2176 17614
rect 2136 17332 2188 17338
rect 2136 17274 2188 17280
rect 1676 16652 1728 16658
rect 1676 16594 1728 16600
rect 1400 16584 1452 16590
rect 1400 16526 1452 16532
rect 1412 16046 1440 16526
rect 1400 16040 1452 16046
rect 1400 15982 1452 15988
rect 1412 14414 1440 15982
rect 1688 15162 1716 16594
rect 1860 16448 1912 16454
rect 1860 16390 1912 16396
rect 1768 15496 1820 15502
rect 1768 15438 1820 15444
rect 1676 15156 1728 15162
rect 1676 15098 1728 15104
rect 1400 14408 1452 14414
rect 1400 14350 1452 14356
rect 1676 14408 1728 14414
rect 1676 14350 1728 14356
rect 1412 14278 1440 14350
rect 1400 14272 1452 14278
rect 1400 14214 1452 14220
rect 1412 12306 1440 14214
rect 1688 13530 1716 14350
rect 1676 13524 1728 13530
rect 1676 13466 1728 13472
rect 1780 13394 1808 15438
rect 1872 15178 1900 16390
rect 1872 15150 1992 15178
rect 1860 15088 1912 15094
rect 1860 15030 1912 15036
rect 1872 13938 1900 15030
rect 1860 13932 1912 13938
rect 1860 13874 1912 13880
rect 1768 13388 1820 13394
rect 1768 13330 1820 13336
rect 1400 12300 1452 12306
rect 1400 12242 1452 12248
rect 1676 12232 1728 12238
rect 1676 12174 1728 12180
rect 1688 11558 1716 12174
rect 1780 11694 1808 13330
rect 1872 12850 1900 13874
rect 1860 12844 1912 12850
rect 1860 12786 1912 12792
rect 1768 11688 1820 11694
rect 1768 11630 1820 11636
rect 1872 11626 1900 12786
rect 1860 11620 1912 11626
rect 1860 11562 1912 11568
rect 1676 11552 1728 11558
rect 1676 11494 1728 11500
rect 1400 9920 1452 9926
rect 1400 9862 1452 9868
rect 1412 9586 1440 9862
rect 1400 9580 1452 9586
rect 1400 9522 1452 9528
rect 1412 9042 1440 9522
rect 1768 9512 1820 9518
rect 1768 9454 1820 9460
rect 1400 9036 1452 9042
rect 1400 8978 1452 8984
rect 1412 7954 1440 8978
rect 1780 8634 1808 9454
rect 1768 8628 1820 8634
rect 1768 8570 1820 8576
rect 1860 8424 1912 8430
rect 1860 8366 1912 8372
rect 1400 7948 1452 7954
rect 1400 7890 1452 7896
rect 1412 5710 1440 7890
rect 1676 7880 1728 7886
rect 1676 7822 1728 7828
rect 1688 6118 1716 7822
rect 1872 6254 1900 8366
rect 1860 6248 1912 6254
rect 1860 6190 1912 6196
rect 1676 6112 1728 6118
rect 1676 6054 1728 6060
rect 1400 5704 1452 5710
rect 1400 5646 1452 5652
rect 1676 5704 1728 5710
rect 1676 5646 1728 5652
rect 1412 4622 1440 5646
rect 1688 5370 1716 5646
rect 1676 5364 1728 5370
rect 1676 5306 1728 5312
rect 1400 4616 1452 4622
rect 1400 4558 1452 4564
rect 1676 4616 1728 4622
rect 1676 4558 1728 4564
rect 1412 3534 1440 4558
rect 1688 3942 1716 4558
rect 1872 4078 1900 6190
rect 1860 4072 1912 4078
rect 1860 4014 1912 4020
rect 1676 3936 1728 3942
rect 1676 3878 1728 3884
rect 1400 3528 1452 3534
rect 570 3496 626 3505
rect 1400 3470 1452 3476
rect 570 3431 626 3440
rect 584 800 612 3431
rect 1964 2514 1992 15150
rect 2136 14952 2188 14958
rect 2136 14894 2188 14900
rect 2148 14074 2176 14894
rect 2136 14068 2188 14074
rect 2136 14010 2188 14016
rect 2148 11150 2176 14010
rect 2136 11144 2188 11150
rect 2136 11086 2188 11092
rect 2240 10606 2268 24210
rect 2780 24200 2832 24206
rect 2780 24142 2832 24148
rect 2412 24132 2464 24138
rect 2412 24074 2464 24080
rect 2424 23730 2452 24074
rect 2412 23724 2464 23730
rect 2412 23666 2464 23672
rect 2792 22137 2820 24142
rect 2884 23662 2912 24210
rect 2872 23656 2924 23662
rect 2872 23598 2924 23604
rect 2964 22432 3016 22438
rect 2964 22374 3016 22380
rect 2778 22128 2834 22137
rect 2778 22063 2834 22072
rect 2320 21956 2372 21962
rect 2320 21898 2372 21904
rect 2332 21010 2360 21898
rect 2976 21554 3004 22374
rect 2964 21548 3016 21554
rect 2964 21490 3016 21496
rect 2976 21010 3004 21490
rect 2320 21004 2372 21010
rect 2320 20946 2372 20952
rect 2964 21004 3016 21010
rect 2964 20946 3016 20952
rect 2872 20052 2924 20058
rect 2872 19994 2924 20000
rect 2884 18850 2912 19994
rect 2964 19780 3016 19786
rect 2964 19722 3016 19728
rect 2976 19310 3004 19722
rect 2964 19304 3016 19310
rect 2964 19246 3016 19252
rect 2320 18828 2372 18834
rect 2320 18770 2372 18776
rect 2688 18828 2740 18834
rect 2884 18822 3004 18850
rect 2688 18770 2740 18776
rect 2332 18290 2360 18770
rect 2700 18426 2728 18770
rect 2872 18760 2924 18766
rect 2872 18702 2924 18708
rect 2688 18420 2740 18426
rect 2688 18362 2740 18368
rect 2320 18284 2372 18290
rect 2320 18226 2372 18232
rect 2884 17134 2912 18702
rect 2872 17128 2924 17134
rect 2872 17070 2924 17076
rect 2976 16674 3004 18822
rect 3068 16794 3096 28047
rect 3252 28014 3280 29038
rect 3344 28150 3372 31282
rect 3528 30190 3556 31418
rect 3620 30938 3648 32914
rect 3700 32360 3752 32366
rect 3700 32302 3752 32308
rect 3712 31278 3740 32302
rect 3700 31272 3752 31278
rect 3700 31214 3752 31220
rect 3608 30932 3660 30938
rect 3608 30874 3660 30880
rect 3608 30796 3660 30802
rect 3608 30738 3660 30744
rect 3620 30326 3648 30738
rect 3608 30320 3660 30326
rect 3608 30262 3660 30268
rect 3712 30258 3740 31214
rect 3700 30252 3752 30258
rect 3700 30194 3752 30200
rect 3516 30184 3568 30190
rect 3516 30126 3568 30132
rect 3528 29850 3556 30126
rect 3516 29844 3568 29850
rect 3516 29786 3568 29792
rect 3332 28144 3384 28150
rect 3332 28086 3384 28092
rect 3240 28008 3292 28014
rect 3240 27950 3292 27956
rect 3240 27532 3292 27538
rect 3240 27474 3292 27480
rect 3148 27464 3200 27470
rect 3148 27406 3200 27412
rect 3160 26926 3188 27406
rect 3148 26920 3200 26926
rect 3148 26862 3200 26868
rect 3160 25838 3188 26862
rect 3252 25838 3280 27474
rect 3148 25832 3200 25838
rect 3148 25774 3200 25780
rect 3240 25832 3292 25838
rect 3240 25774 3292 25780
rect 3160 25158 3188 25774
rect 3252 25498 3280 25774
rect 3240 25492 3292 25498
rect 3240 25434 3292 25440
rect 3148 25152 3200 25158
rect 3148 25094 3200 25100
rect 3160 24206 3188 25094
rect 3252 24818 3280 25434
rect 3240 24812 3292 24818
rect 3240 24754 3292 24760
rect 3252 24274 3280 24754
rect 3240 24268 3292 24274
rect 3240 24210 3292 24216
rect 3148 24200 3200 24206
rect 3148 24142 3200 24148
rect 3160 23730 3188 24142
rect 3148 23724 3200 23730
rect 3148 23666 3200 23672
rect 3332 23656 3384 23662
rect 3332 23598 3384 23604
rect 3148 22772 3200 22778
rect 3148 22714 3200 22720
rect 3160 22098 3188 22714
rect 3344 22506 3372 23598
rect 3608 23180 3660 23186
rect 3608 23122 3660 23128
rect 3620 22778 3648 23122
rect 3608 22772 3660 22778
rect 3608 22714 3660 22720
rect 3700 22568 3752 22574
rect 3700 22510 3752 22516
rect 3332 22500 3384 22506
rect 3332 22442 3384 22448
rect 3148 22092 3200 22098
rect 3148 22034 3200 22040
rect 3712 22030 3740 22510
rect 3424 22024 3476 22030
rect 3422 21992 3424 22001
rect 3700 22024 3752 22030
rect 3476 21992 3478 22001
rect 3478 21950 3556 21978
rect 3700 21966 3752 21972
rect 3422 21927 3478 21936
rect 3148 21888 3200 21894
rect 3148 21830 3200 21836
rect 3160 21486 3188 21830
rect 3148 21480 3200 21486
rect 3148 21422 3200 21428
rect 3424 21480 3476 21486
rect 3424 21422 3476 21428
rect 3436 21010 3464 21422
rect 3424 21004 3476 21010
rect 3424 20946 3476 20952
rect 3436 20398 3464 20946
rect 3528 20602 3556 21950
rect 3516 20596 3568 20602
rect 3516 20538 3568 20544
rect 3424 20392 3476 20398
rect 3424 20334 3476 20340
rect 3148 19848 3200 19854
rect 3148 19790 3200 19796
rect 3160 18834 3188 19790
rect 3148 18828 3200 18834
rect 3148 18770 3200 18776
rect 3424 18828 3476 18834
rect 3424 18770 3476 18776
rect 3436 17882 3464 18770
rect 3424 17876 3476 17882
rect 3424 17818 3476 17824
rect 3700 17536 3752 17542
rect 3700 17478 3752 17484
rect 3712 17134 3740 17478
rect 3700 17128 3752 17134
rect 3700 17070 3752 17076
rect 3056 16788 3108 16794
rect 3056 16730 3108 16736
rect 3148 16788 3200 16794
rect 3148 16730 3200 16736
rect 3160 16674 3188 16730
rect 2976 16646 3188 16674
rect 2688 16040 2740 16046
rect 2688 15982 2740 15988
rect 2700 15706 2728 15982
rect 2688 15700 2740 15706
rect 2688 15642 2740 15648
rect 2976 15570 3004 16646
rect 2964 15564 3016 15570
rect 2964 15506 3016 15512
rect 3148 15564 3200 15570
rect 3148 15506 3200 15512
rect 2780 14952 2832 14958
rect 2780 14894 2832 14900
rect 2792 14618 2820 14894
rect 2780 14612 2832 14618
rect 2780 14554 2832 14560
rect 3160 14385 3188 15506
rect 3804 15366 3832 34031
rect 3988 33998 4016 35634
rect 4724 35494 4752 37266
rect 4804 37120 4856 37126
rect 4804 37062 4856 37068
rect 4816 36242 4844 37062
rect 4804 36236 4856 36242
rect 4804 36178 4856 36184
rect 4896 36168 4948 36174
rect 4896 36110 4948 36116
rect 4712 35488 4764 35494
rect 4712 35430 4764 35436
rect 4712 35148 4764 35154
rect 4712 35090 4764 35096
rect 4724 35018 4752 35090
rect 4908 35018 4936 36110
rect 5368 35494 5396 39200
rect 5448 37392 5500 37398
rect 5448 37334 5500 37340
rect 5460 35698 5488 37334
rect 6920 37324 6972 37330
rect 6920 37266 6972 37272
rect 5632 37256 5684 37262
rect 5632 37198 5684 37204
rect 5644 36650 5672 37198
rect 5724 37120 5776 37126
rect 5724 37062 5776 37068
rect 5632 36644 5684 36650
rect 5632 36586 5684 36592
rect 5736 35850 5764 37062
rect 6828 36848 6880 36854
rect 6828 36790 6880 36796
rect 5816 36712 5868 36718
rect 5816 36654 5868 36660
rect 5644 35822 5764 35850
rect 5644 35766 5672 35822
rect 5632 35760 5684 35766
rect 5632 35702 5684 35708
rect 5448 35692 5500 35698
rect 5448 35634 5500 35640
rect 5264 35488 5316 35494
rect 5264 35430 5316 35436
rect 5356 35488 5408 35494
rect 5356 35430 5408 35436
rect 5276 35222 5304 35430
rect 5264 35216 5316 35222
rect 5264 35158 5316 35164
rect 5460 35154 5488 35634
rect 5540 35556 5592 35562
rect 5540 35498 5592 35504
rect 5448 35148 5500 35154
rect 5448 35090 5500 35096
rect 5552 35034 5580 35498
rect 5644 35154 5672 35702
rect 5632 35148 5684 35154
rect 5632 35090 5684 35096
rect 5828 35034 5856 36654
rect 6736 36168 6788 36174
rect 6736 36110 6788 36116
rect 6276 36100 6328 36106
rect 6276 36042 6328 36048
rect 4712 35012 4764 35018
rect 4712 34954 4764 34960
rect 4896 35012 4948 35018
rect 5552 35006 5856 35034
rect 4896 34954 4948 34960
rect 4220 34844 4516 34864
rect 4276 34842 4300 34844
rect 4356 34842 4380 34844
rect 4436 34842 4460 34844
rect 4298 34790 4300 34842
rect 4362 34790 4374 34842
rect 4436 34790 4438 34842
rect 4276 34788 4300 34790
rect 4356 34788 4380 34790
rect 4436 34788 4460 34790
rect 4220 34768 4516 34788
rect 4160 34604 4212 34610
rect 4160 34546 4212 34552
rect 4172 34066 4200 34546
rect 4620 34536 4672 34542
rect 4620 34478 4672 34484
rect 4160 34060 4212 34066
rect 4160 34002 4212 34008
rect 3976 33992 4028 33998
rect 3976 33934 4028 33940
rect 3988 33522 4016 33934
rect 4220 33756 4516 33776
rect 4276 33754 4300 33756
rect 4356 33754 4380 33756
rect 4436 33754 4460 33756
rect 4298 33702 4300 33754
rect 4362 33702 4374 33754
rect 4436 33702 4438 33754
rect 4276 33700 4300 33702
rect 4356 33700 4380 33702
rect 4436 33700 4460 33702
rect 4220 33680 4516 33700
rect 4632 33658 4660 34478
rect 4620 33652 4672 33658
rect 4620 33594 4672 33600
rect 3976 33516 4028 33522
rect 3976 33458 4028 33464
rect 4632 33454 4660 33594
rect 4160 33448 4212 33454
rect 4160 33390 4212 33396
rect 4620 33448 4672 33454
rect 4620 33390 4672 33396
rect 4172 33046 4200 33390
rect 4620 33312 4672 33318
rect 4620 33254 4672 33260
rect 4160 33040 4212 33046
rect 4160 32982 4212 32988
rect 4068 32904 4120 32910
rect 4068 32846 4120 32852
rect 4632 32892 4660 33254
rect 4724 33046 4752 34954
rect 5540 34672 5592 34678
rect 5540 34614 5592 34620
rect 5080 33992 5132 33998
rect 5080 33934 5132 33940
rect 4712 33040 4764 33046
rect 4712 32982 4764 32988
rect 4712 32904 4764 32910
rect 4632 32864 4712 32892
rect 3976 32496 4028 32502
rect 3976 32438 4028 32444
rect 3884 32360 3936 32366
rect 3884 32302 3936 32308
rect 3896 31278 3924 32302
rect 3988 31482 4016 32438
rect 4080 32434 4108 32846
rect 4220 32668 4516 32688
rect 4276 32666 4300 32668
rect 4356 32666 4380 32668
rect 4436 32666 4460 32668
rect 4298 32614 4300 32666
rect 4362 32614 4374 32666
rect 4436 32614 4438 32666
rect 4276 32612 4300 32614
rect 4356 32612 4380 32614
rect 4436 32612 4460 32614
rect 4220 32592 4516 32612
rect 4068 32428 4120 32434
rect 4068 32370 4120 32376
rect 4632 32366 4660 32864
rect 4712 32846 4764 32852
rect 4620 32360 4672 32366
rect 4620 32302 4672 32308
rect 4436 31952 4488 31958
rect 4436 31894 4488 31900
rect 4448 31822 4476 31894
rect 4436 31816 4488 31822
rect 4436 31758 4488 31764
rect 4220 31580 4516 31600
rect 4276 31578 4300 31580
rect 4356 31578 4380 31580
rect 4436 31578 4460 31580
rect 4298 31526 4300 31578
rect 4362 31526 4374 31578
rect 4436 31526 4438 31578
rect 4276 31524 4300 31526
rect 4356 31524 4380 31526
rect 4436 31524 4460 31526
rect 4220 31504 4516 31524
rect 3976 31476 4028 31482
rect 3976 31418 4028 31424
rect 3884 31272 3936 31278
rect 4436 31272 4488 31278
rect 3884 31214 3936 31220
rect 4434 31240 4436 31249
rect 4632 31260 4660 32302
rect 5092 31958 5120 33934
rect 5552 33674 5580 34614
rect 5644 34542 5672 35006
rect 5632 34536 5684 34542
rect 5632 34478 5684 34484
rect 5724 34536 5776 34542
rect 5724 34478 5776 34484
rect 5552 33646 5672 33674
rect 5540 33380 5592 33386
rect 5540 33322 5592 33328
rect 5552 32434 5580 33322
rect 5644 33114 5672 33646
rect 5736 33454 5764 34478
rect 6000 34468 6052 34474
rect 6000 34410 6052 34416
rect 6012 34202 6040 34410
rect 6000 34196 6052 34202
rect 6000 34138 6052 34144
rect 5724 33448 5776 33454
rect 5724 33390 5776 33396
rect 5632 33108 5684 33114
rect 5632 33050 5684 33056
rect 5540 32428 5592 32434
rect 5540 32370 5592 32376
rect 5736 32366 5764 33390
rect 5724 32360 5776 32366
rect 5724 32302 5776 32308
rect 6012 32298 6040 34138
rect 6092 33584 6144 33590
rect 6092 33526 6144 33532
rect 6104 32570 6132 33526
rect 6288 33130 6316 36042
rect 6460 35556 6512 35562
rect 6460 35498 6512 35504
rect 6472 35154 6500 35498
rect 6460 35148 6512 35154
rect 6460 35090 6512 35096
rect 6644 33516 6696 33522
rect 6644 33458 6696 33464
rect 6288 33114 6408 33130
rect 6288 33108 6420 33114
rect 6288 33102 6368 33108
rect 6368 33050 6420 33056
rect 6276 32972 6328 32978
rect 6276 32914 6328 32920
rect 6184 32904 6236 32910
rect 6184 32846 6236 32852
rect 6092 32564 6144 32570
rect 6092 32506 6144 32512
rect 6000 32292 6052 32298
rect 6000 32234 6052 32240
rect 5080 31952 5132 31958
rect 5080 31894 5132 31900
rect 4988 31884 5040 31890
rect 4988 31826 5040 31832
rect 4488 31240 4660 31260
rect 4490 31232 4660 31240
rect 3896 30190 3924 31214
rect 4434 31175 4490 31184
rect 4220 30492 4516 30512
rect 4276 30490 4300 30492
rect 4356 30490 4380 30492
rect 4436 30490 4460 30492
rect 4298 30438 4300 30490
rect 4362 30438 4374 30490
rect 4436 30438 4438 30490
rect 4276 30436 4300 30438
rect 4356 30436 4380 30438
rect 4436 30436 4460 30438
rect 4220 30416 4516 30436
rect 4712 30252 4764 30258
rect 4712 30194 4764 30200
rect 3884 30184 3936 30190
rect 3884 30126 3936 30132
rect 3896 29850 3924 30126
rect 3884 29844 3936 29850
rect 3884 29786 3936 29792
rect 4620 29844 4672 29850
rect 4620 29786 4672 29792
rect 4068 29708 4120 29714
rect 4068 29650 4120 29656
rect 4080 29306 4108 29650
rect 4220 29404 4516 29424
rect 4276 29402 4300 29404
rect 4356 29402 4380 29404
rect 4436 29402 4460 29404
rect 4298 29350 4300 29402
rect 4362 29350 4374 29402
rect 4436 29350 4438 29402
rect 4276 29348 4300 29350
rect 4356 29348 4380 29350
rect 4436 29348 4460 29350
rect 4220 29328 4516 29348
rect 4068 29300 4120 29306
rect 4068 29242 4120 29248
rect 4632 29102 4660 29786
rect 4724 29170 4752 30194
rect 5000 30054 5028 31826
rect 5092 31804 5120 31894
rect 5172 31816 5224 31822
rect 5092 31776 5172 31804
rect 5172 31758 5224 31764
rect 5540 31816 5592 31822
rect 5540 31758 5592 31764
rect 5184 30122 5212 31758
rect 5552 30938 5580 31758
rect 5816 31680 5868 31686
rect 5816 31622 5868 31628
rect 5632 31408 5684 31414
rect 5632 31350 5684 31356
rect 5540 30932 5592 30938
rect 5540 30874 5592 30880
rect 5644 30802 5672 31350
rect 5828 31278 5856 31622
rect 5816 31272 5868 31278
rect 5816 31214 5868 31220
rect 5632 30796 5684 30802
rect 5632 30738 5684 30744
rect 5632 30592 5684 30598
rect 5632 30534 5684 30540
rect 5172 30116 5224 30122
rect 5172 30058 5224 30064
rect 4988 30048 5040 30054
rect 4988 29990 5040 29996
rect 4804 29844 4856 29850
rect 4804 29786 4856 29792
rect 4712 29164 4764 29170
rect 4712 29106 4764 29112
rect 4068 29096 4120 29102
rect 4068 29038 4120 29044
rect 4620 29096 4672 29102
rect 4620 29038 4672 29044
rect 4080 28014 4108 29038
rect 4632 28626 4660 29038
rect 4620 28620 4672 28626
rect 4620 28562 4672 28568
rect 4724 28558 4752 29106
rect 4816 29034 4844 29786
rect 4804 29028 4856 29034
rect 4804 28970 4856 28976
rect 4896 28960 4948 28966
rect 4896 28902 4948 28908
rect 4908 28626 4936 28902
rect 4896 28620 4948 28626
rect 4896 28562 4948 28568
rect 4712 28552 4764 28558
rect 4712 28494 4764 28500
rect 4220 28316 4516 28336
rect 4276 28314 4300 28316
rect 4356 28314 4380 28316
rect 4436 28314 4460 28316
rect 4298 28262 4300 28314
rect 4362 28262 4374 28314
rect 4436 28262 4438 28314
rect 4276 28260 4300 28262
rect 4356 28260 4380 28262
rect 4436 28260 4460 28262
rect 4220 28240 4516 28260
rect 4724 28218 4752 28494
rect 4712 28212 4764 28218
rect 4712 28154 4764 28160
rect 4068 28008 4120 28014
rect 4068 27950 4120 27956
rect 4080 27538 4108 27950
rect 4896 27668 4948 27674
rect 4896 27610 4948 27616
rect 4068 27532 4120 27538
rect 4068 27474 4120 27480
rect 4080 27130 4108 27474
rect 4620 27328 4672 27334
rect 4620 27270 4672 27276
rect 4220 27228 4516 27248
rect 4276 27226 4300 27228
rect 4356 27226 4380 27228
rect 4436 27226 4460 27228
rect 4298 27174 4300 27226
rect 4362 27174 4374 27226
rect 4436 27174 4438 27226
rect 4276 27172 4300 27174
rect 4356 27172 4380 27174
rect 4436 27172 4460 27174
rect 4220 27152 4516 27172
rect 4068 27124 4120 27130
rect 4068 27066 4120 27072
rect 4632 27044 4660 27270
rect 4804 27124 4856 27130
rect 4804 27066 4856 27072
rect 4540 27016 4660 27044
rect 4068 26920 4120 26926
rect 4068 26862 4120 26868
rect 3976 26036 4028 26042
rect 3976 25978 4028 25984
rect 3988 25838 4016 25978
rect 3976 25832 4028 25838
rect 3976 25774 4028 25780
rect 4080 25362 4108 26862
rect 4540 26382 4568 27016
rect 4620 26920 4672 26926
rect 4620 26862 4672 26868
rect 4528 26376 4580 26382
rect 4528 26318 4580 26324
rect 4220 26140 4516 26160
rect 4276 26138 4300 26140
rect 4356 26138 4380 26140
rect 4436 26138 4460 26140
rect 4298 26086 4300 26138
rect 4362 26086 4374 26138
rect 4436 26086 4438 26138
rect 4276 26084 4300 26086
rect 4356 26084 4380 26086
rect 4436 26084 4460 26086
rect 4220 26064 4516 26084
rect 4632 25906 4660 26862
rect 4712 26852 4764 26858
rect 4712 26794 4764 26800
rect 4724 26382 4752 26794
rect 4816 26450 4844 27066
rect 4908 26926 4936 27610
rect 5000 27538 5028 29990
rect 5184 29782 5212 30058
rect 5264 30048 5316 30054
rect 5264 29990 5316 29996
rect 5448 30048 5500 30054
rect 5448 29990 5500 29996
rect 5276 29850 5304 29990
rect 5264 29844 5316 29850
rect 5264 29786 5316 29792
rect 5172 29776 5224 29782
rect 5172 29718 5224 29724
rect 5264 29708 5316 29714
rect 5264 29650 5316 29656
rect 5276 29594 5304 29650
rect 5276 29566 5396 29594
rect 5172 29028 5224 29034
rect 5172 28970 5224 28976
rect 4988 27532 5040 27538
rect 4988 27474 5040 27480
rect 4896 26920 4948 26926
rect 4896 26862 4948 26868
rect 4804 26444 4856 26450
rect 4804 26386 4856 26392
rect 4712 26376 4764 26382
rect 4712 26318 4764 26324
rect 4620 25900 4672 25906
rect 4620 25842 4672 25848
rect 4724 25838 4752 26318
rect 4804 26240 4856 26246
rect 4804 26182 4856 26188
rect 4896 26240 4948 26246
rect 4896 26182 4948 26188
rect 4712 25832 4764 25838
rect 4712 25774 4764 25780
rect 4816 25650 4844 26182
rect 4724 25622 4844 25650
rect 4068 25356 4120 25362
rect 4068 25298 4120 25304
rect 3974 25120 4030 25129
rect 3974 25055 4030 25064
rect 3988 19417 4016 25055
rect 4080 24818 4108 25298
rect 4724 25226 4752 25622
rect 4712 25220 4764 25226
rect 4712 25162 4764 25168
rect 4220 25052 4516 25072
rect 4276 25050 4300 25052
rect 4356 25050 4380 25052
rect 4436 25050 4460 25052
rect 4298 24998 4300 25050
rect 4362 24998 4374 25050
rect 4436 24998 4438 25050
rect 4276 24996 4300 24998
rect 4356 24996 4380 24998
rect 4436 24996 4460 24998
rect 4220 24976 4516 24996
rect 4068 24812 4120 24818
rect 4068 24754 4120 24760
rect 4724 24206 4752 25162
rect 4908 24342 4936 26182
rect 5184 25838 5212 28970
rect 5368 28558 5396 29566
rect 5460 28694 5488 29990
rect 5644 29714 5672 30534
rect 5908 30184 5960 30190
rect 5908 30126 5960 30132
rect 5632 29708 5684 29714
rect 5632 29650 5684 29656
rect 5920 29170 5948 30126
rect 6104 29238 6132 32506
rect 6196 31278 6224 32846
rect 6288 32434 6316 32914
rect 6276 32428 6328 32434
rect 6276 32370 6328 32376
rect 6184 31272 6236 31278
rect 6184 31214 6236 31220
rect 6092 29232 6144 29238
rect 6092 29174 6144 29180
rect 5908 29164 5960 29170
rect 5908 29106 5960 29112
rect 5448 28688 5500 28694
rect 5448 28630 5500 28636
rect 5356 28552 5408 28558
rect 5356 28494 5408 28500
rect 5368 28014 5396 28494
rect 5460 28082 5488 28630
rect 5816 28620 5868 28626
rect 5816 28562 5868 28568
rect 5724 28484 5776 28490
rect 5724 28426 5776 28432
rect 5448 28076 5500 28082
rect 5448 28018 5500 28024
rect 5356 28008 5408 28014
rect 5276 27968 5356 27996
rect 5276 27674 5304 27968
rect 5356 27950 5408 27956
rect 5264 27668 5316 27674
rect 5264 27610 5316 27616
rect 5736 27538 5764 28426
rect 5828 28150 5856 28562
rect 5816 28144 5868 28150
rect 5816 28086 5868 28092
rect 5724 27532 5776 27538
rect 5724 27474 5776 27480
rect 6104 26874 6132 29174
rect 6380 28014 6408 33050
rect 6460 31748 6512 31754
rect 6460 31690 6512 31696
rect 6472 30666 6500 31690
rect 6552 30728 6604 30734
rect 6552 30670 6604 30676
rect 6460 30660 6512 30666
rect 6460 30602 6512 30608
rect 6368 28008 6420 28014
rect 6368 27950 6420 27956
rect 6380 27470 6408 27950
rect 6368 27464 6420 27470
rect 6368 27406 6420 27412
rect 6012 26858 6132 26874
rect 6000 26852 6132 26858
rect 6052 26846 6132 26852
rect 6000 26794 6052 26800
rect 6472 26246 6500 30602
rect 6564 29714 6592 30670
rect 6656 30394 6684 33458
rect 6644 30388 6696 30394
rect 6644 30330 6696 30336
rect 6552 29708 6604 29714
rect 6552 29650 6604 29656
rect 6460 26240 6512 26246
rect 6460 26182 6512 26188
rect 5172 25832 5224 25838
rect 5172 25774 5224 25780
rect 5632 25832 5684 25838
rect 5632 25774 5684 25780
rect 5644 25362 5672 25774
rect 6000 25696 6052 25702
rect 6000 25638 6052 25644
rect 5632 25356 5684 25362
rect 5632 25298 5684 25304
rect 5540 25288 5592 25294
rect 5540 25230 5592 25236
rect 5552 24818 5580 25230
rect 5540 24812 5592 24818
rect 5540 24754 5592 24760
rect 5448 24744 5500 24750
rect 5448 24686 5500 24692
rect 4896 24336 4948 24342
rect 4896 24278 4948 24284
rect 4712 24200 4764 24206
rect 4712 24142 4764 24148
rect 4220 23964 4516 23984
rect 4276 23962 4300 23964
rect 4356 23962 4380 23964
rect 4436 23962 4460 23964
rect 4298 23910 4300 23962
rect 4362 23910 4374 23962
rect 4436 23910 4438 23962
rect 4276 23908 4300 23910
rect 4356 23908 4380 23910
rect 4436 23908 4460 23910
rect 4220 23888 4516 23908
rect 4620 23588 4672 23594
rect 4620 23530 4672 23536
rect 4528 23520 4580 23526
rect 4528 23462 4580 23468
rect 4540 23186 4568 23462
rect 4528 23180 4580 23186
rect 4528 23122 4580 23128
rect 4068 23112 4120 23118
rect 4068 23054 4120 23060
rect 4080 22658 4108 23054
rect 4220 22876 4516 22896
rect 4276 22874 4300 22876
rect 4356 22874 4380 22876
rect 4436 22874 4460 22876
rect 4298 22822 4300 22874
rect 4362 22822 4374 22874
rect 4436 22822 4438 22874
rect 4276 22820 4300 22822
rect 4356 22820 4380 22822
rect 4436 22820 4460 22822
rect 4220 22800 4516 22820
rect 4632 22778 4660 23530
rect 4724 23118 4752 24142
rect 5460 23662 5488 24686
rect 6012 24274 6040 25638
rect 6000 24268 6052 24274
rect 6000 24210 6052 24216
rect 6184 23724 6236 23730
rect 6184 23666 6236 23672
rect 5448 23656 5500 23662
rect 5448 23598 5500 23604
rect 4712 23112 4764 23118
rect 4712 23054 4764 23060
rect 4620 22772 4672 22778
rect 4620 22714 4672 22720
rect 4080 22630 4200 22658
rect 4068 22024 4120 22030
rect 4068 21966 4120 21972
rect 4080 21418 4108 21966
rect 4172 21962 4200 22630
rect 4632 22098 4660 22714
rect 4712 22568 4764 22574
rect 4712 22510 4764 22516
rect 5356 22568 5408 22574
rect 5460 22556 5488 23598
rect 5632 22976 5684 22982
rect 5632 22918 5684 22924
rect 5644 22642 5672 22918
rect 5632 22636 5684 22642
rect 5632 22578 5684 22584
rect 5408 22528 5488 22556
rect 5540 22568 5592 22574
rect 5356 22510 5408 22516
rect 5540 22510 5592 22516
rect 4620 22092 4672 22098
rect 4620 22034 4672 22040
rect 4160 21956 4212 21962
rect 4160 21898 4212 21904
rect 4724 21894 4752 22510
rect 4896 22092 4948 22098
rect 4896 22034 4948 22040
rect 4712 21888 4764 21894
rect 4712 21830 4764 21836
rect 4220 21788 4516 21808
rect 4276 21786 4300 21788
rect 4356 21786 4380 21788
rect 4436 21786 4460 21788
rect 4298 21734 4300 21786
rect 4362 21734 4374 21786
rect 4436 21734 4438 21786
rect 4276 21732 4300 21734
rect 4356 21732 4380 21734
rect 4436 21732 4460 21734
rect 4220 21712 4516 21732
rect 4804 21480 4856 21486
rect 4804 21422 4856 21428
rect 4068 21412 4120 21418
rect 4068 21354 4120 21360
rect 4712 21412 4764 21418
rect 4712 21354 4764 21360
rect 4080 21146 4108 21354
rect 4620 21344 4672 21350
rect 4620 21286 4672 21292
rect 4068 21140 4120 21146
rect 4068 21082 4120 21088
rect 4220 20700 4516 20720
rect 4276 20698 4300 20700
rect 4356 20698 4380 20700
rect 4436 20698 4460 20700
rect 4298 20646 4300 20698
rect 4362 20646 4374 20698
rect 4436 20646 4438 20698
rect 4276 20644 4300 20646
rect 4356 20644 4380 20646
rect 4436 20644 4460 20646
rect 4220 20624 4516 20644
rect 4632 20058 4660 21286
rect 4724 20398 4752 21354
rect 4712 20392 4764 20398
rect 4712 20334 4764 20340
rect 4620 20052 4672 20058
rect 4620 19994 4672 20000
rect 4724 19922 4752 20334
rect 4528 19916 4580 19922
rect 4712 19916 4764 19922
rect 4580 19876 4660 19904
rect 4528 19858 4580 19864
rect 4632 19802 4660 19876
rect 4712 19858 4764 19864
rect 4816 19802 4844 21422
rect 4908 20398 4936 22034
rect 5552 21486 5580 22510
rect 5644 22098 5672 22578
rect 5632 22092 5684 22098
rect 5632 22034 5684 22040
rect 6196 21554 6224 23666
rect 6552 23656 6604 23662
rect 6552 23598 6604 23604
rect 6564 23050 6592 23598
rect 6552 23044 6604 23050
rect 6552 22986 6604 22992
rect 6184 21548 6236 21554
rect 6184 21490 6236 21496
rect 5540 21480 5592 21486
rect 5540 21422 5592 21428
rect 5264 21344 5316 21350
rect 5264 21286 5316 21292
rect 5276 21010 5304 21286
rect 5552 21010 5580 21422
rect 6196 21010 6224 21490
rect 5264 21004 5316 21010
rect 5264 20946 5316 20952
rect 5540 21004 5592 21010
rect 5540 20946 5592 20952
rect 6184 21004 6236 21010
rect 6184 20946 6236 20952
rect 6460 21004 6512 21010
rect 6460 20946 6512 20952
rect 4988 20528 5040 20534
rect 4988 20470 5040 20476
rect 4896 20392 4948 20398
rect 4896 20334 4948 20340
rect 4908 19990 4936 20334
rect 4896 19984 4948 19990
rect 4896 19926 4948 19932
rect 4632 19774 4844 19802
rect 4220 19612 4516 19632
rect 4276 19610 4300 19612
rect 4356 19610 4380 19612
rect 4436 19610 4460 19612
rect 4298 19558 4300 19610
rect 4362 19558 4374 19610
rect 4436 19558 4438 19610
rect 4276 19556 4300 19558
rect 4356 19556 4380 19558
rect 4436 19556 4460 19558
rect 4220 19536 4516 19556
rect 4632 19514 4660 19774
rect 4620 19508 4672 19514
rect 4620 19450 4672 19456
rect 4528 19440 4580 19446
rect 3974 19408 4030 19417
rect 4528 19382 4580 19388
rect 4712 19440 4764 19446
rect 4712 19382 4764 19388
rect 3974 19343 4030 19352
rect 4540 19310 4568 19382
rect 4528 19304 4580 19310
rect 4528 19246 4580 19252
rect 4068 19236 4120 19242
rect 4068 19178 4120 19184
rect 4080 19145 4108 19178
rect 4066 19136 4122 19145
rect 4066 19071 4122 19080
rect 3976 18964 4028 18970
rect 3976 18906 4028 18912
rect 3988 18222 4016 18906
rect 4620 18692 4672 18698
rect 4620 18634 4672 18640
rect 4220 18524 4516 18544
rect 4276 18522 4300 18524
rect 4356 18522 4380 18524
rect 4436 18522 4460 18524
rect 4298 18470 4300 18522
rect 4362 18470 4374 18522
rect 4436 18470 4438 18522
rect 4276 18468 4300 18470
rect 4356 18468 4380 18470
rect 4436 18468 4460 18470
rect 4220 18448 4516 18468
rect 3976 18216 4028 18222
rect 3976 18158 4028 18164
rect 4632 17746 4660 18634
rect 4724 18222 4752 19382
rect 4712 18216 4764 18222
rect 4712 18158 4764 18164
rect 4620 17740 4672 17746
rect 4620 17682 4672 17688
rect 4220 17436 4516 17456
rect 4276 17434 4300 17436
rect 4356 17434 4380 17436
rect 4436 17434 4460 17436
rect 4298 17382 4300 17434
rect 4362 17382 4374 17434
rect 4436 17382 4438 17434
rect 4276 17380 4300 17382
rect 4356 17380 4380 17382
rect 4436 17380 4460 17382
rect 4220 17360 4516 17380
rect 5000 17134 5028 20470
rect 5276 20398 5304 20946
rect 5908 20936 5960 20942
rect 5908 20878 5960 20884
rect 6276 20936 6328 20942
rect 6276 20878 6328 20884
rect 5920 20398 5948 20878
rect 5264 20392 5316 20398
rect 5264 20334 5316 20340
rect 5908 20392 5960 20398
rect 5908 20334 5960 20340
rect 5276 19786 5304 20334
rect 5264 19780 5316 19786
rect 5264 19722 5316 19728
rect 6288 19718 6316 20878
rect 6368 20256 6420 20262
rect 6368 20198 6420 20204
rect 6380 19922 6408 20198
rect 6368 19916 6420 19922
rect 6368 19858 6420 19864
rect 6276 19712 6328 19718
rect 6276 19654 6328 19660
rect 6000 19440 6052 19446
rect 6000 19382 6052 19388
rect 5264 19304 5316 19310
rect 5264 19246 5316 19252
rect 5448 19304 5500 19310
rect 5448 19246 5500 19252
rect 5276 18834 5304 19246
rect 5264 18828 5316 18834
rect 5264 18770 5316 18776
rect 5460 18426 5488 19246
rect 6012 19242 6040 19382
rect 5908 19236 5960 19242
rect 5908 19178 5960 19184
rect 6000 19236 6052 19242
rect 6000 19178 6052 19184
rect 5920 18970 5948 19178
rect 5908 18964 5960 18970
rect 5908 18906 5960 18912
rect 6092 18964 6144 18970
rect 6092 18906 6144 18912
rect 5632 18828 5684 18834
rect 5632 18770 5684 18776
rect 5908 18828 5960 18834
rect 5908 18770 5960 18776
rect 5644 18630 5672 18770
rect 5632 18624 5684 18630
rect 5632 18566 5684 18572
rect 5448 18420 5500 18426
rect 5448 18362 5500 18368
rect 5460 17746 5488 18362
rect 5920 18154 5948 18770
rect 6104 18426 6132 18906
rect 6184 18828 6236 18834
rect 6184 18770 6236 18776
rect 6196 18426 6224 18770
rect 6092 18420 6144 18426
rect 6092 18362 6144 18368
rect 6184 18420 6236 18426
rect 6184 18362 6236 18368
rect 6288 18222 6316 19654
rect 6472 19310 6500 20946
rect 6460 19304 6512 19310
rect 6460 19246 6512 19252
rect 6276 18216 6328 18222
rect 6276 18158 6328 18164
rect 5908 18148 5960 18154
rect 5908 18090 5960 18096
rect 5448 17740 5500 17746
rect 5448 17682 5500 17688
rect 5908 17740 5960 17746
rect 5908 17682 5960 17688
rect 5356 17672 5408 17678
rect 5356 17614 5408 17620
rect 4988 17128 5040 17134
rect 4988 17070 5040 17076
rect 4160 16652 4212 16658
rect 4160 16594 4212 16600
rect 4172 16538 4200 16594
rect 4080 16510 4200 16538
rect 4080 16250 4108 16510
rect 4220 16348 4516 16368
rect 4276 16346 4300 16348
rect 4356 16346 4380 16348
rect 4436 16346 4460 16348
rect 4298 16294 4300 16346
rect 4362 16294 4374 16346
rect 4436 16294 4438 16346
rect 4276 16292 4300 16294
rect 4356 16292 4380 16294
rect 4436 16292 4460 16294
rect 4220 16272 4516 16292
rect 4068 16244 4120 16250
rect 4068 16186 4120 16192
rect 5368 16114 5396 17614
rect 5920 17202 5948 17682
rect 6000 17332 6052 17338
rect 6000 17274 6052 17280
rect 5632 17196 5684 17202
rect 5632 17138 5684 17144
rect 5908 17196 5960 17202
rect 5908 17138 5960 17144
rect 5644 16726 5672 17138
rect 5908 17060 5960 17066
rect 5908 17002 5960 17008
rect 5920 16726 5948 17002
rect 5632 16720 5684 16726
rect 5632 16662 5684 16668
rect 5908 16720 5960 16726
rect 5908 16662 5960 16668
rect 5540 16652 5592 16658
rect 5540 16594 5592 16600
rect 5448 16584 5500 16590
rect 5448 16526 5500 16532
rect 5356 16108 5408 16114
rect 5356 16050 5408 16056
rect 4528 16040 4580 16046
rect 4528 15982 4580 15988
rect 4066 15872 4122 15881
rect 4066 15807 4122 15816
rect 4080 15638 4108 15807
rect 4540 15706 4568 15982
rect 4528 15700 4580 15706
rect 4528 15642 4580 15648
rect 4068 15632 4120 15638
rect 5460 15586 5488 16526
rect 5552 16250 5580 16594
rect 5540 16244 5592 16250
rect 5540 16186 5592 16192
rect 5644 15706 5672 16662
rect 6012 16658 6040 17274
rect 6000 16652 6052 16658
rect 6000 16594 6052 16600
rect 5632 15700 5684 15706
rect 5632 15642 5684 15648
rect 4068 15574 4120 15580
rect 4712 15564 4764 15570
rect 4712 15506 4764 15512
rect 5368 15558 5488 15586
rect 5632 15564 5684 15570
rect 3792 15360 3844 15366
rect 3792 15302 3844 15308
rect 4220 15260 4516 15280
rect 4276 15258 4300 15260
rect 4356 15258 4380 15260
rect 4436 15258 4460 15260
rect 4298 15206 4300 15258
rect 4362 15206 4374 15258
rect 4436 15206 4438 15258
rect 4276 15204 4300 15206
rect 4356 15204 4380 15206
rect 4436 15204 4460 15206
rect 4220 15184 4516 15204
rect 4724 15042 4752 15506
rect 5368 15162 5396 15558
rect 5632 15506 5684 15512
rect 5356 15156 5408 15162
rect 5356 15098 5408 15104
rect 4632 15026 4752 15042
rect 4620 15020 4752 15026
rect 4672 15014 4752 15020
rect 4620 14962 4672 14968
rect 4160 14952 4212 14958
rect 4160 14894 4212 14900
rect 3976 14476 4028 14482
rect 3976 14418 4028 14424
rect 3146 14376 3202 14385
rect 3146 14311 3202 14320
rect 3988 13870 4016 14418
rect 4172 14414 4200 14894
rect 4724 14482 4752 15014
rect 4712 14476 4764 14482
rect 4712 14418 4764 14424
rect 4988 14476 5040 14482
rect 4988 14418 5040 14424
rect 4160 14408 4212 14414
rect 4160 14350 4212 14356
rect 4220 14172 4516 14192
rect 4276 14170 4300 14172
rect 4356 14170 4380 14172
rect 4436 14170 4460 14172
rect 4298 14118 4300 14170
rect 4362 14118 4374 14170
rect 4436 14118 4438 14170
rect 4276 14116 4300 14118
rect 4356 14116 4380 14118
rect 4436 14116 4460 14118
rect 4220 14096 4516 14116
rect 5000 13870 5028 14418
rect 5080 14340 5132 14346
rect 5080 14282 5132 14288
rect 3976 13864 4028 13870
rect 3976 13806 4028 13812
rect 4988 13864 5040 13870
rect 4988 13806 5040 13812
rect 3332 13728 3384 13734
rect 3332 13670 3384 13676
rect 2870 13424 2926 13433
rect 2700 13382 2870 13410
rect 2700 12889 2728 13382
rect 3344 13394 3372 13670
rect 3988 13462 4016 13806
rect 4896 13796 4948 13802
rect 4896 13738 4948 13744
rect 3976 13456 4028 13462
rect 3976 13398 4028 13404
rect 2870 13359 2926 13368
rect 3332 13388 3384 13394
rect 3332 13330 3384 13336
rect 2686 12880 2742 12889
rect 2686 12815 2742 12824
rect 3988 12782 4016 13398
rect 4620 13388 4672 13394
rect 4620 13330 4672 13336
rect 4632 13274 4660 13330
rect 4908 13326 4936 13738
rect 4896 13320 4948 13326
rect 4632 13246 4752 13274
rect 4896 13262 4948 13268
rect 4620 13184 4672 13190
rect 4620 13126 4672 13132
rect 4220 13084 4516 13104
rect 4276 13082 4300 13084
rect 4356 13082 4380 13084
rect 4436 13082 4460 13084
rect 4298 13030 4300 13082
rect 4362 13030 4374 13082
rect 4436 13030 4438 13082
rect 4276 13028 4300 13030
rect 4356 13028 4380 13030
rect 4436 13028 4460 13030
rect 4220 13008 4516 13028
rect 4632 12850 4660 13126
rect 4620 12844 4672 12850
rect 4620 12786 4672 12792
rect 3976 12776 4028 12782
rect 3976 12718 4028 12724
rect 4160 12776 4212 12782
rect 4160 12718 4212 12724
rect 2964 12164 3016 12170
rect 2964 12106 3016 12112
rect 2412 12096 2464 12102
rect 2412 12038 2464 12044
rect 2424 11218 2452 12038
rect 2976 11762 3004 12106
rect 4172 12084 4200 12718
rect 4724 12714 4752 13246
rect 4712 12708 4764 12714
rect 4712 12650 4764 12656
rect 4724 12306 4752 12650
rect 4712 12300 4764 12306
rect 4712 12242 4764 12248
rect 4804 12232 4856 12238
rect 4804 12174 4856 12180
rect 4080 12056 4200 12084
rect 4080 11898 4108 12056
rect 4220 11996 4516 12016
rect 4276 11994 4300 11996
rect 4356 11994 4380 11996
rect 4436 11994 4460 11996
rect 4298 11942 4300 11994
rect 4362 11942 4374 11994
rect 4436 11942 4438 11994
rect 4276 11940 4300 11942
rect 4356 11940 4380 11942
rect 4436 11940 4460 11942
rect 4220 11920 4516 11940
rect 4068 11892 4120 11898
rect 4068 11834 4120 11840
rect 4620 11892 4672 11898
rect 4620 11834 4672 11840
rect 2964 11756 3016 11762
rect 2964 11698 3016 11704
rect 4632 11218 4660 11834
rect 4816 11694 4844 12174
rect 4804 11688 4856 11694
rect 4804 11630 4856 11636
rect 4908 11558 4936 13262
rect 5000 12918 5028 13806
rect 4988 12912 5040 12918
rect 4988 12854 5040 12860
rect 4896 11552 4948 11558
rect 4896 11494 4948 11500
rect 5092 11354 5120 14282
rect 5368 14074 5396 15098
rect 5644 14958 5672 15506
rect 5816 15496 5868 15502
rect 5816 15438 5868 15444
rect 6276 15496 6328 15502
rect 6276 15438 6328 15444
rect 5632 14952 5684 14958
rect 5632 14894 5684 14900
rect 5448 14408 5500 14414
rect 5448 14350 5500 14356
rect 5356 14068 5408 14074
rect 5356 14010 5408 14016
rect 5460 13870 5488 14350
rect 5448 13864 5500 13870
rect 5448 13806 5500 13812
rect 5460 12782 5488 13806
rect 5448 12776 5500 12782
rect 5448 12718 5500 12724
rect 5264 12300 5316 12306
rect 5264 12242 5316 12248
rect 5276 11898 5304 12242
rect 5264 11892 5316 11898
rect 5264 11834 5316 11840
rect 5264 11688 5316 11694
rect 5264 11630 5316 11636
rect 5356 11688 5408 11694
rect 5356 11630 5408 11636
rect 5080 11348 5132 11354
rect 5080 11290 5132 11296
rect 2412 11212 2464 11218
rect 2412 11154 2464 11160
rect 4620 11212 4672 11218
rect 4620 11154 4672 11160
rect 2872 11144 2924 11150
rect 2872 11086 2924 11092
rect 2228 10600 2280 10606
rect 2228 10542 2280 10548
rect 2320 10464 2372 10470
rect 2320 10406 2372 10412
rect 2332 9518 2360 10406
rect 2778 9888 2834 9897
rect 2778 9823 2834 9832
rect 2792 9722 2820 9823
rect 2780 9716 2832 9722
rect 2780 9658 2832 9664
rect 2320 9512 2372 9518
rect 2320 9454 2372 9460
rect 2136 8968 2188 8974
rect 2136 8910 2188 8916
rect 2148 8498 2176 8910
rect 2136 8492 2188 8498
rect 2136 8434 2188 8440
rect 2332 8430 2360 9454
rect 2320 8424 2372 8430
rect 2320 8366 2372 8372
rect 2780 8356 2832 8362
rect 2780 8298 2832 8304
rect 2792 8090 2820 8298
rect 2780 8084 2832 8090
rect 2780 8026 2832 8032
rect 2596 7336 2648 7342
rect 2596 7278 2648 7284
rect 2608 6866 2636 7278
rect 2778 6896 2834 6905
rect 2596 6860 2648 6866
rect 2778 6831 2834 6840
rect 2596 6802 2648 6808
rect 2136 6792 2188 6798
rect 2136 6734 2188 6740
rect 2148 6390 2176 6734
rect 2136 6384 2188 6390
rect 2136 6326 2188 6332
rect 2792 5914 2820 6831
rect 2780 5908 2832 5914
rect 2780 5850 2832 5856
rect 2044 5160 2096 5166
rect 2044 5102 2096 5108
rect 2056 4826 2084 5102
rect 2044 4820 2096 4826
rect 2044 4762 2096 4768
rect 2596 3528 2648 3534
rect 2596 3470 2648 3476
rect 2608 2990 2636 3470
rect 2884 3058 2912 11086
rect 4620 11076 4672 11082
rect 4620 11018 4672 11024
rect 4220 10908 4516 10928
rect 4276 10906 4300 10908
rect 4356 10906 4380 10908
rect 4436 10906 4460 10908
rect 4298 10854 4300 10906
rect 4362 10854 4374 10906
rect 4436 10854 4438 10906
rect 4276 10852 4300 10854
rect 4356 10852 4380 10854
rect 4436 10852 4460 10854
rect 4220 10832 4516 10852
rect 4632 10674 4660 11018
rect 4620 10668 4672 10674
rect 4620 10610 4672 10616
rect 2964 10600 3016 10606
rect 2964 10542 3016 10548
rect 3148 10600 3200 10606
rect 4804 10600 4856 10606
rect 3148 10542 3200 10548
rect 3606 10568 3662 10577
rect 2976 10130 3004 10542
rect 3160 10266 3188 10542
rect 4804 10542 4856 10548
rect 3606 10503 3608 10512
rect 3660 10503 3662 10512
rect 3608 10474 3660 10480
rect 3148 10260 3200 10266
rect 3148 10202 3200 10208
rect 2964 10124 3016 10130
rect 2964 10066 3016 10072
rect 4620 10124 4672 10130
rect 4620 10066 4672 10072
rect 2976 8566 3004 10066
rect 3608 10056 3660 10062
rect 3608 9998 3660 10004
rect 3620 9382 3648 9998
rect 4220 9820 4516 9840
rect 4276 9818 4300 9820
rect 4356 9818 4380 9820
rect 4436 9818 4460 9820
rect 4298 9766 4300 9818
rect 4362 9766 4374 9818
rect 4436 9766 4438 9818
rect 4276 9764 4300 9766
rect 4356 9764 4380 9766
rect 4436 9764 4460 9766
rect 4220 9744 4516 9764
rect 3608 9376 3660 9382
rect 3608 9318 3660 9324
rect 4632 9110 4660 10066
rect 4620 9104 4672 9110
rect 4620 9046 4672 9052
rect 4712 8900 4764 8906
rect 4712 8842 4764 8848
rect 4220 8732 4516 8752
rect 4276 8730 4300 8732
rect 4356 8730 4380 8732
rect 4436 8730 4460 8732
rect 4298 8678 4300 8730
rect 4362 8678 4374 8730
rect 4436 8678 4438 8730
rect 4276 8676 4300 8678
rect 4356 8676 4380 8678
rect 4436 8676 4460 8678
rect 4220 8656 4516 8676
rect 2964 8560 3016 8566
rect 2964 8502 3016 8508
rect 2976 5030 3004 8502
rect 4724 8498 4752 8842
rect 4712 8492 4764 8498
rect 4712 8434 4764 8440
rect 4160 8424 4212 8430
rect 4160 8366 4212 8372
rect 4172 7954 4200 8366
rect 4528 8356 4580 8362
rect 4528 8298 4580 8304
rect 4540 8242 4568 8298
rect 4540 8214 4752 8242
rect 4160 7948 4212 7954
rect 4160 7890 4212 7896
rect 4620 7948 4672 7954
rect 4620 7890 4672 7896
rect 4220 7644 4516 7664
rect 4276 7642 4300 7644
rect 4356 7642 4380 7644
rect 4436 7642 4460 7644
rect 4298 7590 4300 7642
rect 4362 7590 4374 7642
rect 4436 7590 4438 7642
rect 4276 7588 4300 7590
rect 4356 7588 4380 7590
rect 4436 7588 4460 7590
rect 4220 7568 4516 7588
rect 4632 7546 4660 7890
rect 4620 7540 4672 7546
rect 4620 7482 4672 7488
rect 4160 7336 4212 7342
rect 4160 7278 4212 7284
rect 4172 6798 4200 7278
rect 4724 6866 4752 8214
rect 4816 7818 4844 10542
rect 5092 10130 5120 11290
rect 5276 10538 5304 11630
rect 5264 10532 5316 10538
rect 5264 10474 5316 10480
rect 5080 10124 5132 10130
rect 5080 10066 5132 10072
rect 4896 9512 4948 9518
rect 4896 9454 4948 9460
rect 4908 8634 4936 9454
rect 4896 8628 4948 8634
rect 4896 8570 4948 8576
rect 4988 7948 5040 7954
rect 4988 7890 5040 7896
rect 4804 7812 4856 7818
rect 4804 7754 4856 7760
rect 5000 7342 5028 7890
rect 5368 7410 5396 11630
rect 5540 9376 5592 9382
rect 5540 9318 5592 9324
rect 5552 9042 5580 9318
rect 5540 9036 5592 9042
rect 5540 8978 5592 8984
rect 5540 8424 5592 8430
rect 5540 8366 5592 8372
rect 5356 7404 5408 7410
rect 5356 7346 5408 7352
rect 4804 7336 4856 7342
rect 4804 7278 4856 7284
rect 4988 7336 5040 7342
rect 4988 7278 5040 7284
rect 4712 6860 4764 6866
rect 4712 6802 4764 6808
rect 4160 6792 4212 6798
rect 4160 6734 4212 6740
rect 4620 6792 4672 6798
rect 4620 6734 4672 6740
rect 3424 6656 3476 6662
rect 3424 6598 3476 6604
rect 3436 5778 3464 6598
rect 4220 6556 4516 6576
rect 4276 6554 4300 6556
rect 4356 6554 4380 6556
rect 4436 6554 4460 6556
rect 4298 6502 4300 6554
rect 4362 6502 4374 6554
rect 4436 6502 4438 6554
rect 4276 6500 4300 6502
rect 4356 6500 4380 6502
rect 4436 6500 4460 6502
rect 4220 6480 4516 6500
rect 4632 6254 4660 6734
rect 4068 6248 4120 6254
rect 4068 6190 4120 6196
rect 4620 6248 4672 6254
rect 4620 6190 4672 6196
rect 4080 5914 4108 6190
rect 4068 5908 4120 5914
rect 4068 5850 4120 5856
rect 3424 5772 3476 5778
rect 3424 5714 3476 5720
rect 4220 5468 4516 5488
rect 4276 5466 4300 5468
rect 4356 5466 4380 5468
rect 4436 5466 4460 5468
rect 4298 5414 4300 5466
rect 4362 5414 4374 5466
rect 4436 5414 4438 5466
rect 4276 5412 4300 5414
rect 4356 5412 4380 5414
rect 4436 5412 4460 5414
rect 4220 5392 4516 5412
rect 3240 5228 3292 5234
rect 3240 5170 3292 5176
rect 2964 5024 3016 5030
rect 2964 4966 3016 4972
rect 3252 4146 3280 5170
rect 4632 5166 4660 6190
rect 3792 5160 3844 5166
rect 3792 5102 3844 5108
rect 4620 5160 4672 5166
rect 4620 5102 4672 5108
rect 3424 5024 3476 5030
rect 3424 4966 3476 4972
rect 3240 4140 3292 4146
rect 3240 4082 3292 4088
rect 2964 4072 3016 4078
rect 2964 4014 3016 4020
rect 2976 3738 3004 4014
rect 2964 3732 3016 3738
rect 2964 3674 3016 3680
rect 3436 3534 3464 4966
rect 3804 4026 3832 5102
rect 4620 4480 4672 4486
rect 4620 4422 4672 4428
rect 4220 4380 4516 4400
rect 4276 4378 4300 4380
rect 4356 4378 4380 4380
rect 4436 4378 4460 4380
rect 4298 4326 4300 4378
rect 4362 4326 4374 4378
rect 4436 4326 4438 4378
rect 4276 4324 4300 4326
rect 4356 4324 4380 4326
rect 4436 4324 4460 4326
rect 4220 4304 4516 4324
rect 4632 4146 4660 4422
rect 4620 4140 4672 4146
rect 4620 4082 4672 4088
rect 3804 4010 4016 4026
rect 3804 4004 4028 4010
rect 3804 3998 3976 4004
rect 3424 3528 3476 3534
rect 3424 3470 3476 3476
rect 3804 3194 3832 3998
rect 3976 3946 4028 3952
rect 4816 3942 4844 7278
rect 5264 6724 5316 6730
rect 5264 6666 5316 6672
rect 4988 6656 5040 6662
rect 4988 6598 5040 6604
rect 5080 6656 5132 6662
rect 5080 6598 5132 6604
rect 5000 6322 5028 6598
rect 4988 6316 5040 6322
rect 4988 6258 5040 6264
rect 5092 5778 5120 6598
rect 5276 6186 5304 6666
rect 5552 6322 5580 8366
rect 5644 8362 5672 14894
rect 5828 14278 5856 15438
rect 5906 15192 5962 15201
rect 5906 15127 5962 15136
rect 5816 14272 5868 14278
rect 5816 14214 5868 14220
rect 5920 13870 5948 15127
rect 6288 15094 6316 15438
rect 6000 15088 6052 15094
rect 6000 15030 6052 15036
rect 6276 15088 6328 15094
rect 6276 15030 6328 15036
rect 5908 13864 5960 13870
rect 5908 13806 5960 13812
rect 6012 13394 6040 15030
rect 6184 14952 6236 14958
rect 6184 14894 6236 14900
rect 6000 13388 6052 13394
rect 6000 13330 6052 13336
rect 6000 13252 6052 13258
rect 6000 13194 6052 13200
rect 6012 12714 6040 13194
rect 6000 12708 6052 12714
rect 6000 12650 6052 12656
rect 5816 11824 5868 11830
rect 5816 11766 5868 11772
rect 5828 11218 5856 11766
rect 6196 11234 6224 14894
rect 6288 14890 6316 15030
rect 6276 14884 6328 14890
rect 6276 14826 6328 14832
rect 6368 13320 6420 13326
rect 6368 13262 6420 13268
rect 6380 12918 6408 13262
rect 6644 12980 6696 12986
rect 6644 12922 6696 12928
rect 6368 12912 6420 12918
rect 6368 12854 6420 12860
rect 6656 12782 6684 12922
rect 6644 12776 6696 12782
rect 6644 12718 6696 12724
rect 6460 12640 6512 12646
rect 6460 12582 6512 12588
rect 6644 12640 6696 12646
rect 6644 12582 6696 12588
rect 6276 11892 6328 11898
rect 6276 11834 6328 11840
rect 6288 11762 6316 11834
rect 6472 11762 6500 12582
rect 6552 12300 6604 12306
rect 6552 12242 6604 12248
rect 6276 11756 6328 11762
rect 6276 11698 6328 11704
rect 6460 11756 6512 11762
rect 6460 11698 6512 11704
rect 5816 11212 5868 11218
rect 5816 11154 5868 11160
rect 6104 11206 6224 11234
rect 6288 11218 6316 11698
rect 6472 11286 6500 11698
rect 6460 11280 6512 11286
rect 6460 11222 6512 11228
rect 6276 11212 6328 11218
rect 5816 10600 5868 10606
rect 5816 10542 5868 10548
rect 5828 10266 5856 10542
rect 5816 10260 5868 10266
rect 5816 10202 5868 10208
rect 5816 10056 5868 10062
rect 5816 9998 5868 10004
rect 5828 9382 5856 9998
rect 5816 9376 5868 9382
rect 5816 9318 5868 9324
rect 6000 8968 6052 8974
rect 6000 8910 6052 8916
rect 6012 8566 6040 8910
rect 6000 8560 6052 8566
rect 6000 8502 6052 8508
rect 5632 8356 5684 8362
rect 5632 8298 5684 8304
rect 5908 8356 5960 8362
rect 5908 8298 5960 8304
rect 5920 7018 5948 8298
rect 5828 6990 5948 7018
rect 5540 6316 5592 6322
rect 5540 6258 5592 6264
rect 5264 6180 5316 6186
rect 5264 6122 5316 6128
rect 5276 5778 5304 6122
rect 5080 5772 5132 5778
rect 5080 5714 5132 5720
rect 5264 5772 5316 5778
rect 5264 5714 5316 5720
rect 5276 5030 5304 5714
rect 5828 5166 5856 6990
rect 5908 6860 5960 6866
rect 5908 6802 5960 6808
rect 5920 6186 5948 6802
rect 6012 6254 6040 8502
rect 6104 7954 6132 11206
rect 6276 11154 6328 11160
rect 6184 11144 6236 11150
rect 6184 11086 6236 11092
rect 6196 10674 6224 11086
rect 6184 10668 6236 10674
rect 6184 10610 6236 10616
rect 6564 9586 6592 12242
rect 6656 10606 6684 12582
rect 6748 10674 6776 36110
rect 6840 34610 6868 36790
rect 6932 36582 6960 37266
rect 6920 36576 6972 36582
rect 6920 36518 6972 36524
rect 6932 35630 6960 36518
rect 7392 36378 7420 39200
rect 9416 37398 9444 39200
rect 9404 37392 9456 37398
rect 9404 37334 9456 37340
rect 7564 37324 7616 37330
rect 7564 37266 7616 37272
rect 7840 37324 7892 37330
rect 7840 37266 7892 37272
rect 7932 37324 7984 37330
rect 7932 37266 7984 37272
rect 9680 37324 9732 37330
rect 9864 37324 9916 37330
rect 9680 37266 9732 37272
rect 9784 37284 9864 37312
rect 7472 37188 7524 37194
rect 7472 37130 7524 37136
rect 7484 36922 7512 37130
rect 7472 36916 7524 36922
rect 7472 36858 7524 36864
rect 7576 36802 7604 37266
rect 7484 36774 7604 36802
rect 7484 36718 7512 36774
rect 7472 36712 7524 36718
rect 7472 36654 7524 36660
rect 7380 36372 7432 36378
rect 7380 36314 7432 36320
rect 7484 36224 7512 36654
rect 7392 36196 7512 36224
rect 6920 35624 6972 35630
rect 6920 35566 6972 35572
rect 7392 35154 7420 36196
rect 7748 35488 7800 35494
rect 7748 35430 7800 35436
rect 7380 35148 7432 35154
rect 7380 35090 7432 35096
rect 7012 35080 7064 35086
rect 7012 35022 7064 35028
rect 6920 34740 6972 34746
rect 6920 34682 6972 34688
rect 6828 34604 6880 34610
rect 6828 34546 6880 34552
rect 6932 33998 6960 34682
rect 7024 34474 7052 35022
rect 7288 34536 7340 34542
rect 7288 34478 7340 34484
rect 7012 34468 7064 34474
rect 7012 34410 7064 34416
rect 7024 34134 7052 34410
rect 7012 34128 7064 34134
rect 7012 34070 7064 34076
rect 6920 33992 6972 33998
rect 6920 33934 6972 33940
rect 7024 33658 7052 34070
rect 7300 34066 7328 34478
rect 7288 34060 7340 34066
rect 7288 34002 7340 34008
rect 7012 33652 7064 33658
rect 7012 33594 7064 33600
rect 6920 33448 6972 33454
rect 6920 33390 6972 33396
rect 6932 33130 6960 33390
rect 7300 33318 7328 34002
rect 7288 33312 7340 33318
rect 7288 33254 7340 33260
rect 6932 33102 7144 33130
rect 6828 32904 6880 32910
rect 6828 32846 6880 32852
rect 6840 31958 6868 32846
rect 7116 32026 7144 33102
rect 7300 32230 7328 33254
rect 7392 32774 7420 35090
rect 7760 35086 7788 35430
rect 7564 35080 7616 35086
rect 7564 35022 7616 35028
rect 7748 35080 7800 35086
rect 7748 35022 7800 35028
rect 7576 33590 7604 35022
rect 7656 34400 7708 34406
rect 7656 34342 7708 34348
rect 7564 33584 7616 33590
rect 7564 33526 7616 33532
rect 7668 33454 7696 34342
rect 7472 33448 7524 33454
rect 7470 33416 7472 33425
rect 7656 33448 7708 33454
rect 7524 33416 7526 33425
rect 7656 33390 7708 33396
rect 7470 33351 7526 33360
rect 7564 32836 7616 32842
rect 7564 32778 7616 32784
rect 7380 32768 7432 32774
rect 7380 32710 7432 32716
rect 7288 32224 7340 32230
rect 7288 32166 7340 32172
rect 7104 32020 7156 32026
rect 7104 31962 7156 31968
rect 6828 31952 6880 31958
rect 6828 31894 6880 31900
rect 6840 30802 6868 31894
rect 7116 31482 7144 31962
rect 7104 31476 7156 31482
rect 7104 31418 7156 31424
rect 7392 31346 7420 32710
rect 7380 31340 7432 31346
rect 7380 31282 7432 31288
rect 7012 31272 7064 31278
rect 7012 31214 7064 31220
rect 7024 30802 7052 31214
rect 6828 30796 6880 30802
rect 6828 30738 6880 30744
rect 7012 30796 7064 30802
rect 7012 30738 7064 30744
rect 7288 30252 7340 30258
rect 7288 30194 7340 30200
rect 7012 30184 7064 30190
rect 7012 30126 7064 30132
rect 7024 29646 7052 30126
rect 7196 30048 7248 30054
rect 7196 29990 7248 29996
rect 7012 29640 7064 29646
rect 7012 29582 7064 29588
rect 6828 29164 6880 29170
rect 6828 29106 6880 29112
rect 6840 27606 6868 29106
rect 7024 29102 7052 29582
rect 7012 29096 7064 29102
rect 7012 29038 7064 29044
rect 6920 29028 6972 29034
rect 6920 28970 6972 28976
rect 6932 28014 6960 28970
rect 6920 28008 6972 28014
rect 6920 27950 6972 27956
rect 6828 27600 6880 27606
rect 6828 27542 6880 27548
rect 7208 26926 7236 29990
rect 7300 27402 7328 30194
rect 7576 30190 7604 32778
rect 7656 32292 7708 32298
rect 7656 32234 7708 32240
rect 7668 31890 7696 32234
rect 7656 31884 7708 31890
rect 7656 31826 7708 31832
rect 7668 30802 7696 31826
rect 7656 30796 7708 30802
rect 7656 30738 7708 30744
rect 7380 30184 7432 30190
rect 7380 30126 7432 30132
rect 7564 30184 7616 30190
rect 7564 30126 7616 30132
rect 7392 29782 7420 30126
rect 7380 29776 7432 29782
rect 7380 29718 7432 29724
rect 7392 28762 7420 29718
rect 7576 29578 7604 30126
rect 7564 29572 7616 29578
rect 7564 29514 7616 29520
rect 7564 28960 7616 28966
rect 7564 28902 7616 28908
rect 7380 28756 7432 28762
rect 7380 28698 7432 28704
rect 7576 27878 7604 28902
rect 7564 27872 7616 27878
rect 7564 27814 7616 27820
rect 7288 27396 7340 27402
rect 7288 27338 7340 27344
rect 7380 26988 7432 26994
rect 7380 26930 7432 26936
rect 6920 26920 6972 26926
rect 6920 26862 6972 26868
rect 7196 26920 7248 26926
rect 7196 26862 7248 26868
rect 6828 25152 6880 25158
rect 6828 25094 6880 25100
rect 6840 24614 6868 25094
rect 6932 24750 6960 26862
rect 7208 26450 7236 26862
rect 7392 26790 7420 26930
rect 7380 26784 7432 26790
rect 7380 26726 7432 26732
rect 7472 26784 7524 26790
rect 7472 26726 7524 26732
rect 7196 26444 7248 26450
rect 7248 26404 7328 26432
rect 7196 26386 7248 26392
rect 7012 25832 7064 25838
rect 7012 25774 7064 25780
rect 7024 25498 7052 25774
rect 7012 25492 7064 25498
rect 7012 25434 7064 25440
rect 7012 25356 7064 25362
rect 7012 25298 7064 25304
rect 6920 24744 6972 24750
rect 6920 24686 6972 24692
rect 6828 24608 6880 24614
rect 6828 24550 6880 24556
rect 6840 23594 6868 24550
rect 7024 24342 7052 25298
rect 7196 25288 7248 25294
rect 7196 25230 7248 25236
rect 7208 24818 7236 25230
rect 7196 24812 7248 24818
rect 7196 24754 7248 24760
rect 7104 24676 7156 24682
rect 7104 24618 7156 24624
rect 7012 24336 7064 24342
rect 7012 24278 7064 24284
rect 7116 24274 7144 24618
rect 7104 24268 7156 24274
rect 7104 24210 7156 24216
rect 7300 23662 7328 26404
rect 7392 24018 7420 26726
rect 7484 24206 7512 26726
rect 7472 24200 7524 24206
rect 7472 24142 7524 24148
rect 7392 23990 7512 24018
rect 7288 23656 7340 23662
rect 7288 23598 7340 23604
rect 6828 23588 6880 23594
rect 6828 23530 6880 23536
rect 6840 23186 6868 23530
rect 7300 23254 7328 23598
rect 7288 23248 7340 23254
rect 7288 23190 7340 23196
rect 6828 23180 6880 23186
rect 6828 23122 6880 23128
rect 6840 22574 6868 23122
rect 7300 22710 7328 23190
rect 7380 23180 7432 23186
rect 7380 23122 7432 23128
rect 7392 23050 7420 23122
rect 7380 23044 7432 23050
rect 7380 22986 7432 22992
rect 7288 22704 7340 22710
rect 7288 22646 7340 22652
rect 7392 22642 7420 22986
rect 7380 22636 7432 22642
rect 7380 22578 7432 22584
rect 6828 22568 6880 22574
rect 6828 22510 6880 22516
rect 6840 22234 6868 22510
rect 7484 22234 7512 23990
rect 7576 23322 7604 27814
rect 7656 27532 7708 27538
rect 7656 27474 7708 27480
rect 7564 23316 7616 23322
rect 7564 23258 7616 23264
rect 6828 22228 6880 22234
rect 6828 22170 6880 22176
rect 7472 22228 7524 22234
rect 7472 22170 7524 22176
rect 7288 22024 7340 22030
rect 7288 21966 7340 21972
rect 7012 20936 7064 20942
rect 7012 20878 7064 20884
rect 7024 19310 7052 20878
rect 7104 20800 7156 20806
rect 7104 20742 7156 20748
rect 7116 20466 7144 20742
rect 7104 20460 7156 20466
rect 7104 20402 7156 20408
rect 7300 20398 7328 21966
rect 7668 21894 7696 27474
rect 7748 25968 7800 25974
rect 7748 25910 7800 25916
rect 7760 24818 7788 25910
rect 7748 24812 7800 24818
rect 7748 24754 7800 24760
rect 7748 24268 7800 24274
rect 7748 24210 7800 24216
rect 7760 22642 7788 24210
rect 7748 22636 7800 22642
rect 7748 22578 7800 22584
rect 7748 22500 7800 22506
rect 7748 22442 7800 22448
rect 7760 22166 7788 22442
rect 7748 22160 7800 22166
rect 7748 22102 7800 22108
rect 7656 21888 7708 21894
rect 7656 21830 7708 21836
rect 7380 21004 7432 21010
rect 7380 20946 7432 20952
rect 7288 20392 7340 20398
rect 7288 20334 7340 20340
rect 7300 19922 7328 20334
rect 7288 19916 7340 19922
rect 7288 19858 7340 19864
rect 7288 19780 7340 19786
rect 7288 19722 7340 19728
rect 7300 19310 7328 19722
rect 7392 19378 7420 20946
rect 7472 19848 7524 19854
rect 7472 19790 7524 19796
rect 7380 19372 7432 19378
rect 7380 19314 7432 19320
rect 7484 19310 7512 19790
rect 7012 19304 7064 19310
rect 7012 19246 7064 19252
rect 7288 19304 7340 19310
rect 7288 19246 7340 19252
rect 7472 19304 7524 19310
rect 7472 19246 7524 19252
rect 7024 18834 7052 19246
rect 7300 18834 7328 19246
rect 7484 18902 7512 19246
rect 7472 18896 7524 18902
rect 7472 18838 7524 18844
rect 7012 18828 7064 18834
rect 7012 18770 7064 18776
rect 7288 18828 7340 18834
rect 7288 18770 7340 18776
rect 6920 18080 6972 18086
rect 6920 18022 6972 18028
rect 6932 17134 6960 18022
rect 7024 17814 7052 18770
rect 7472 18624 7524 18630
rect 7472 18566 7524 18572
rect 7484 18222 7512 18566
rect 7472 18216 7524 18222
rect 7472 18158 7524 18164
rect 7012 17808 7064 17814
rect 7012 17750 7064 17756
rect 6920 17128 6972 17134
rect 6920 17070 6972 17076
rect 7196 16992 7248 16998
rect 7196 16934 7248 16940
rect 7564 16992 7616 16998
rect 7564 16934 7616 16940
rect 7104 16584 7156 16590
rect 7104 16526 7156 16532
rect 7116 16114 7144 16526
rect 7104 16108 7156 16114
rect 7104 16050 7156 16056
rect 7208 15570 7236 16934
rect 7576 16658 7604 16934
rect 7564 16652 7616 16658
rect 7564 16594 7616 16600
rect 7196 15564 7248 15570
rect 7196 15506 7248 15512
rect 6826 15056 6882 15065
rect 6826 14991 6882 15000
rect 7380 15020 7432 15026
rect 6840 14958 6868 14991
rect 7380 14962 7432 14968
rect 7564 15020 7616 15026
rect 7564 14962 7616 14968
rect 6828 14952 6880 14958
rect 6828 14894 6880 14900
rect 7104 14952 7156 14958
rect 7104 14894 7156 14900
rect 7012 14816 7064 14822
rect 7012 14758 7064 14764
rect 7024 14550 7052 14758
rect 7012 14544 7064 14550
rect 7012 14486 7064 14492
rect 6920 14476 6972 14482
rect 6920 14418 6972 14424
rect 6932 13870 6960 14418
rect 6920 13864 6972 13870
rect 6920 13806 6972 13812
rect 7024 13546 7052 14486
rect 7116 14414 7144 14894
rect 7104 14408 7156 14414
rect 7104 14350 7156 14356
rect 6840 13518 7052 13546
rect 6840 12646 6868 13518
rect 7012 13184 7064 13190
rect 7012 13126 7064 13132
rect 7024 12782 7052 13126
rect 7012 12776 7064 12782
rect 7012 12718 7064 12724
rect 6828 12640 6880 12646
rect 6828 12582 6880 12588
rect 6840 12306 6868 12582
rect 7024 12374 7052 12718
rect 7012 12368 7064 12374
rect 7012 12310 7064 12316
rect 6828 12300 6880 12306
rect 6828 12242 6880 12248
rect 6920 11212 6972 11218
rect 6920 11154 6972 11160
rect 6736 10668 6788 10674
rect 6736 10610 6788 10616
rect 6644 10600 6696 10606
rect 6644 10542 6696 10548
rect 6552 9580 6604 9586
rect 6552 9522 6604 9528
rect 6656 9518 6684 10542
rect 6736 9988 6788 9994
rect 6736 9930 6788 9936
rect 6644 9512 6696 9518
rect 6644 9454 6696 9460
rect 6460 9036 6512 9042
rect 6460 8978 6512 8984
rect 6092 7948 6144 7954
rect 6092 7890 6144 7896
rect 6104 7342 6132 7890
rect 6472 7818 6500 8978
rect 6748 8106 6776 9930
rect 6826 9072 6882 9081
rect 6826 9007 6828 9016
rect 6880 9007 6882 9016
rect 6828 8978 6880 8984
rect 6932 8634 6960 11154
rect 7024 9654 7052 12310
rect 7104 12164 7156 12170
rect 7104 12106 7156 12112
rect 7116 11694 7144 12106
rect 7392 11694 7420 14962
rect 7104 11688 7156 11694
rect 7104 11630 7156 11636
rect 7380 11688 7432 11694
rect 7380 11630 7432 11636
rect 7116 11354 7144 11630
rect 7104 11348 7156 11354
rect 7104 11290 7156 11296
rect 7576 11218 7604 14962
rect 7668 12986 7696 21830
rect 7760 21690 7788 22102
rect 7748 21684 7800 21690
rect 7748 21626 7800 21632
rect 7748 20528 7800 20534
rect 7748 20470 7800 20476
rect 7760 18222 7788 20470
rect 7748 18216 7800 18222
rect 7748 18158 7800 18164
rect 7760 17134 7788 18158
rect 7852 17542 7880 37266
rect 7944 36854 7972 37266
rect 9692 37194 9720 37266
rect 9680 37188 9732 37194
rect 9680 37130 9732 37136
rect 7932 36848 7984 36854
rect 7932 36790 7984 36796
rect 8208 36712 8260 36718
rect 8208 36654 8260 36660
rect 8220 36310 8248 36654
rect 8208 36304 8260 36310
rect 8208 36246 8260 36252
rect 8392 36236 8444 36242
rect 8392 36178 8444 36184
rect 8024 35488 8076 35494
rect 8024 35430 8076 35436
rect 7932 34604 7984 34610
rect 7932 34546 7984 34552
rect 7944 34066 7972 34546
rect 7932 34060 7984 34066
rect 7932 34002 7984 34008
rect 7932 33584 7984 33590
rect 7932 33526 7984 33532
rect 7944 33454 7972 33526
rect 7932 33448 7984 33454
rect 8036 33425 8064 35430
rect 8404 35290 8432 36178
rect 9784 36174 9812 37284
rect 9864 37266 9916 37272
rect 9864 37120 9916 37126
rect 9864 37062 9916 37068
rect 9876 36718 9904 37062
rect 9864 36712 9916 36718
rect 9864 36654 9916 36660
rect 11060 36712 11112 36718
rect 11060 36654 11112 36660
rect 11520 36712 11572 36718
rect 11520 36654 11572 36660
rect 10048 36576 10100 36582
rect 10048 36518 10100 36524
rect 9772 36168 9824 36174
rect 9772 36110 9824 36116
rect 10060 36106 10088 36518
rect 10140 36372 10192 36378
rect 10140 36314 10192 36320
rect 10152 36242 10180 36314
rect 10140 36236 10192 36242
rect 10416 36236 10468 36242
rect 10192 36196 10272 36224
rect 10140 36178 10192 36184
rect 10048 36100 10100 36106
rect 10048 36042 10100 36048
rect 8484 36032 8536 36038
rect 8484 35974 8536 35980
rect 9680 36032 9732 36038
rect 9680 35974 9732 35980
rect 8496 35698 8524 35974
rect 8484 35692 8536 35698
rect 8484 35634 8536 35640
rect 9692 35562 9720 35974
rect 10060 35630 10088 36042
rect 9956 35624 10008 35630
rect 9956 35566 10008 35572
rect 10048 35624 10100 35630
rect 10048 35566 10100 35572
rect 9680 35556 9732 35562
rect 9680 35498 9732 35504
rect 8392 35284 8444 35290
rect 8392 35226 8444 35232
rect 8300 34944 8352 34950
rect 8300 34886 8352 34892
rect 8312 33998 8340 34886
rect 8404 34066 8432 35226
rect 9680 35148 9732 35154
rect 9680 35090 9732 35096
rect 9692 35018 9720 35090
rect 9680 35012 9732 35018
rect 9680 34954 9732 34960
rect 8576 34672 8628 34678
rect 8576 34614 8628 34620
rect 8588 34202 8616 34614
rect 8576 34196 8628 34202
rect 8576 34138 8628 34144
rect 8392 34060 8444 34066
rect 8392 34002 8444 34008
rect 8300 33992 8352 33998
rect 8300 33934 8352 33940
rect 7932 33390 7984 33396
rect 8022 33416 8078 33425
rect 8022 33351 8078 33360
rect 8312 32960 8340 33934
rect 8484 33312 8536 33318
rect 8484 33254 8536 33260
rect 8496 33046 8524 33254
rect 8484 33040 8536 33046
rect 8484 32982 8536 32988
rect 8588 32978 8616 34138
rect 8760 34060 8812 34066
rect 8760 34002 8812 34008
rect 8772 33454 8800 34002
rect 9692 33658 9720 34954
rect 9968 34950 9996 35566
rect 10060 35222 10088 35566
rect 10244 35222 10272 36196
rect 10416 36178 10468 36184
rect 10428 35698 10456 36178
rect 10416 35692 10468 35698
rect 10416 35634 10468 35640
rect 11072 35630 11100 36654
rect 11428 36576 11480 36582
rect 11428 36518 11480 36524
rect 11152 36168 11204 36174
rect 11152 36110 11204 36116
rect 11164 35698 11192 36110
rect 11152 35692 11204 35698
rect 11152 35634 11204 35640
rect 10876 35624 10928 35630
rect 10876 35566 10928 35572
rect 11060 35624 11112 35630
rect 11060 35566 11112 35572
rect 10888 35222 10916 35566
rect 10048 35216 10100 35222
rect 10048 35158 10100 35164
rect 10232 35216 10284 35222
rect 10232 35158 10284 35164
rect 10876 35216 10928 35222
rect 10876 35158 10928 35164
rect 10324 35148 10376 35154
rect 10324 35090 10376 35096
rect 10784 35148 10836 35154
rect 10784 35090 10836 35096
rect 9864 34944 9916 34950
rect 9864 34886 9916 34892
rect 9956 34944 10008 34950
rect 9956 34886 10008 34892
rect 9876 34542 9904 34886
rect 10336 34610 10364 35090
rect 10796 34762 10824 35090
rect 10704 34734 10824 34762
rect 10324 34604 10376 34610
rect 10324 34546 10376 34552
rect 9864 34536 9916 34542
rect 9916 34496 10180 34524
rect 9864 34478 9916 34484
rect 10152 34134 10180 34496
rect 9772 34128 9824 34134
rect 9772 34070 9824 34076
rect 10140 34128 10192 34134
rect 10140 34070 10192 34076
rect 9680 33652 9732 33658
rect 9680 33594 9732 33600
rect 9784 33454 9812 34070
rect 8760 33448 8812 33454
rect 9128 33448 9180 33454
rect 8760 33390 8812 33396
rect 9126 33416 9128 33425
rect 9772 33448 9824 33454
rect 9180 33416 9182 33425
rect 8668 33380 8720 33386
rect 8668 33322 8720 33328
rect 8392 32972 8444 32978
rect 8312 32932 8392 32960
rect 7932 32564 7984 32570
rect 7932 32506 7984 32512
rect 7944 31822 7972 32506
rect 8024 32496 8076 32502
rect 8024 32438 8076 32444
rect 7932 31816 7984 31822
rect 7932 31758 7984 31764
rect 7932 30116 7984 30122
rect 7932 30058 7984 30064
rect 7944 29714 7972 30058
rect 7932 29708 7984 29714
rect 7932 29650 7984 29656
rect 7932 28620 7984 28626
rect 7932 28562 7984 28568
rect 7944 28150 7972 28562
rect 7932 28144 7984 28150
rect 7932 28086 7984 28092
rect 7944 27470 7972 28086
rect 7932 27464 7984 27470
rect 7932 27406 7984 27412
rect 7944 26926 7972 27406
rect 8036 26994 8064 32438
rect 8312 32366 8340 32932
rect 8392 32914 8444 32920
rect 8576 32972 8628 32978
rect 8576 32914 8628 32920
rect 8588 32434 8616 32914
rect 8576 32428 8628 32434
rect 8576 32370 8628 32376
rect 8208 32360 8260 32366
rect 8208 32302 8260 32308
rect 8300 32360 8352 32366
rect 8300 32302 8352 32308
rect 8220 32230 8248 32302
rect 8208 32224 8260 32230
rect 8208 32166 8260 32172
rect 8220 31890 8248 32166
rect 8116 31884 8168 31890
rect 8116 31826 8168 31832
rect 8208 31884 8260 31890
rect 8208 31826 8260 31832
rect 8128 31770 8156 31826
rect 8312 31770 8340 32302
rect 8392 32292 8444 32298
rect 8392 32234 8444 32240
rect 8128 31742 8340 31770
rect 8116 31272 8168 31278
rect 8116 31214 8168 31220
rect 8128 30870 8156 31214
rect 8116 30864 8168 30870
rect 8116 30806 8168 30812
rect 8404 30802 8432 32234
rect 8680 30802 8708 33322
rect 8772 33130 8800 33390
rect 9772 33390 9824 33396
rect 9126 33351 9182 33360
rect 8772 33102 8892 33130
rect 8864 32978 8892 33102
rect 8760 32972 8812 32978
rect 8760 32914 8812 32920
rect 8852 32972 8904 32978
rect 8852 32914 8904 32920
rect 8772 32366 8800 32914
rect 8864 32434 8892 32914
rect 9588 32904 9640 32910
rect 9588 32846 9640 32852
rect 9220 32768 9272 32774
rect 9220 32710 9272 32716
rect 8852 32428 8904 32434
rect 8852 32370 8904 32376
rect 8760 32360 8812 32366
rect 8760 32302 8812 32308
rect 8864 32026 8892 32370
rect 9232 32026 9260 32710
rect 8852 32020 8904 32026
rect 8852 31962 8904 31968
rect 9220 32020 9272 32026
rect 9220 31962 9272 31968
rect 9600 31890 9628 32846
rect 9784 32298 9812 33390
rect 9956 32904 10008 32910
rect 9956 32846 10008 32852
rect 9772 32292 9824 32298
rect 9772 32234 9824 32240
rect 8852 31884 8904 31890
rect 8852 31826 8904 31832
rect 9588 31884 9640 31890
rect 9588 31826 9640 31832
rect 8392 30796 8444 30802
rect 8392 30738 8444 30744
rect 8668 30796 8720 30802
rect 8668 30738 8720 30744
rect 8864 30326 8892 31826
rect 9784 31482 9812 32234
rect 9968 31686 9996 32846
rect 9956 31680 10008 31686
rect 9956 31622 10008 31628
rect 9772 31476 9824 31482
rect 9772 31418 9824 31424
rect 8944 30796 8996 30802
rect 8944 30738 8996 30744
rect 8852 30320 8904 30326
rect 8852 30262 8904 30268
rect 8392 30184 8444 30190
rect 8392 30126 8444 30132
rect 8404 29714 8432 30126
rect 8392 29708 8444 29714
rect 8392 29650 8444 29656
rect 8484 29504 8536 29510
rect 8484 29446 8536 29452
rect 8208 28416 8260 28422
rect 8208 28358 8260 28364
rect 8220 28218 8248 28358
rect 8208 28212 8260 28218
rect 8208 28154 8260 28160
rect 8116 27532 8168 27538
rect 8116 27474 8168 27480
rect 8128 27130 8156 27474
rect 8116 27124 8168 27130
rect 8116 27066 8168 27072
rect 8024 26988 8076 26994
rect 8024 26930 8076 26936
rect 7932 26920 7984 26926
rect 7932 26862 7984 26868
rect 7932 25832 7984 25838
rect 7932 25774 7984 25780
rect 7944 23866 7972 25774
rect 8024 24200 8076 24206
rect 8024 24142 8076 24148
rect 7932 23860 7984 23866
rect 7932 23802 7984 23808
rect 8036 22438 8064 24142
rect 8116 23656 8168 23662
rect 8116 23598 8168 23604
rect 8128 23186 8156 23598
rect 8116 23180 8168 23186
rect 8116 23122 8168 23128
rect 8128 22506 8156 23122
rect 8116 22500 8168 22506
rect 8116 22442 8168 22448
rect 8024 22432 8076 22438
rect 8024 22374 8076 22380
rect 8116 21344 8168 21350
rect 8116 21286 8168 21292
rect 8128 20398 8156 21286
rect 8220 21078 8248 28154
rect 8496 28014 8524 29446
rect 8668 29096 8720 29102
rect 8668 29038 8720 29044
rect 8680 28150 8708 29038
rect 8668 28144 8720 28150
rect 8668 28086 8720 28092
rect 8484 28008 8536 28014
rect 8484 27950 8536 27956
rect 8392 27532 8444 27538
rect 8392 27474 8444 27480
rect 8404 26314 8432 27474
rect 8392 26308 8444 26314
rect 8392 26250 8444 26256
rect 8392 25832 8444 25838
rect 8392 25774 8444 25780
rect 8404 25702 8432 25774
rect 8392 25696 8444 25702
rect 8392 25638 8444 25644
rect 8404 24818 8432 25638
rect 8392 24812 8444 24818
rect 8392 24754 8444 24760
rect 8404 24342 8432 24754
rect 8392 24336 8444 24342
rect 8392 24278 8444 24284
rect 8496 23322 8524 27950
rect 8680 26994 8708 28086
rect 8864 28014 8892 30262
rect 8852 28008 8904 28014
rect 8852 27950 8904 27956
rect 8956 27606 8984 30738
rect 9784 30734 9812 31418
rect 9956 31272 10008 31278
rect 9956 31214 10008 31220
rect 9772 30728 9824 30734
rect 9772 30670 9824 30676
rect 9220 30592 9272 30598
rect 9220 30534 9272 30540
rect 9128 30116 9180 30122
rect 9128 30058 9180 30064
rect 9036 29640 9088 29646
rect 9036 29582 9088 29588
rect 9048 29510 9076 29582
rect 9140 29510 9168 30058
rect 9036 29504 9088 29510
rect 9036 29446 9088 29452
rect 9128 29504 9180 29510
rect 9128 29446 9180 29452
rect 8944 27600 8996 27606
rect 8944 27542 8996 27548
rect 8852 27328 8904 27334
rect 8852 27270 8904 27276
rect 8668 26988 8720 26994
rect 8668 26930 8720 26936
rect 8864 26450 8892 27270
rect 9232 26994 9260 30534
rect 9404 30184 9456 30190
rect 9404 30126 9456 30132
rect 9416 29102 9444 30126
rect 9968 29306 9996 31214
rect 10048 31136 10100 31142
rect 10048 31078 10100 31084
rect 10060 30258 10088 31078
rect 10324 30796 10376 30802
rect 10324 30738 10376 30744
rect 10048 30252 10100 30258
rect 10048 30194 10100 30200
rect 9956 29300 10008 29306
rect 9956 29242 10008 29248
rect 9404 29096 9456 29102
rect 9404 29038 9456 29044
rect 9680 28960 9732 28966
rect 9680 28902 9732 28908
rect 9692 28150 9720 28902
rect 10336 28626 10364 30738
rect 10416 30592 10468 30598
rect 10416 30534 10468 30540
rect 10428 29170 10456 30534
rect 10598 30152 10654 30161
rect 10598 30087 10654 30096
rect 10612 29578 10640 30087
rect 10600 29572 10652 29578
rect 10600 29514 10652 29520
rect 10416 29164 10468 29170
rect 10416 29106 10468 29112
rect 10704 29102 10732 34734
rect 10784 34672 10836 34678
rect 10784 34614 10836 34620
rect 10796 34542 10824 34614
rect 10784 34536 10836 34542
rect 10784 34478 10836 34484
rect 10796 34218 10824 34478
rect 11072 34406 11100 35566
rect 11440 35154 11468 36518
rect 11532 35630 11560 36654
rect 11520 35624 11572 35630
rect 11520 35566 11572 35572
rect 11532 35154 11560 35566
rect 11428 35148 11480 35154
rect 11428 35090 11480 35096
rect 11520 35148 11572 35154
rect 11520 35090 11572 35096
rect 11520 34604 11572 34610
rect 11520 34546 11572 34552
rect 11152 34468 11204 34474
rect 11152 34410 11204 34416
rect 11060 34400 11112 34406
rect 11060 34342 11112 34348
rect 11164 34218 11192 34410
rect 10796 34190 11192 34218
rect 11244 34196 11296 34202
rect 10876 34128 10928 34134
rect 10876 34070 10928 34076
rect 10888 32366 10916 34070
rect 11072 34066 11100 34190
rect 11244 34138 11296 34144
rect 11060 34060 11112 34066
rect 11060 34002 11112 34008
rect 10876 32360 10928 32366
rect 10876 32302 10928 32308
rect 10888 31890 10916 32302
rect 11072 32298 11100 34002
rect 11256 33454 11284 34138
rect 11532 34066 11560 34546
rect 11520 34060 11572 34066
rect 11520 34002 11572 34008
rect 11244 33448 11296 33454
rect 11244 33390 11296 33396
rect 11244 33312 11296 33318
rect 11244 33254 11296 33260
rect 11256 33114 11284 33254
rect 11244 33108 11296 33114
rect 11244 33050 11296 33056
rect 11336 33040 11388 33046
rect 11336 32982 11388 32988
rect 11152 32972 11204 32978
rect 11152 32914 11204 32920
rect 11060 32292 11112 32298
rect 11060 32234 11112 32240
rect 10876 31884 10928 31890
rect 10876 31826 10928 31832
rect 10784 31680 10836 31686
rect 10784 31622 10836 31628
rect 10796 31346 10824 31622
rect 10784 31340 10836 31346
rect 10784 31282 10836 31288
rect 11164 30802 11192 32914
rect 11348 32366 11376 32982
rect 11336 32360 11388 32366
rect 11336 32302 11388 32308
rect 11244 31884 11296 31890
rect 11244 31826 11296 31832
rect 11256 31414 11284 31826
rect 11244 31408 11296 31414
rect 11244 31350 11296 31356
rect 11348 31278 11376 32302
rect 11428 31748 11480 31754
rect 11428 31690 11480 31696
rect 11336 31272 11388 31278
rect 11336 31214 11388 31220
rect 11152 30796 11204 30802
rect 11152 30738 11204 30744
rect 11440 30734 11468 31690
rect 11428 30728 11480 30734
rect 11428 30670 11480 30676
rect 11624 30190 11652 39200
rect 11704 37324 11756 37330
rect 11704 37266 11756 37272
rect 11716 35086 11744 37266
rect 12256 37120 12308 37126
rect 13648 37108 13676 39200
rect 15476 37256 15528 37262
rect 15476 37198 15528 37204
rect 13648 37080 13860 37108
rect 12256 37062 12308 37068
rect 11796 36576 11848 36582
rect 11796 36518 11848 36524
rect 11704 35080 11756 35086
rect 11704 35022 11756 35028
rect 11808 34066 11836 36518
rect 12268 36242 12296 37062
rect 13832 36854 13860 37080
rect 13820 36848 13872 36854
rect 13820 36790 13872 36796
rect 15488 36718 15516 37198
rect 12440 36712 12492 36718
rect 12440 36654 12492 36660
rect 12808 36712 12860 36718
rect 12808 36654 12860 36660
rect 15476 36712 15528 36718
rect 15476 36654 15528 36660
rect 12256 36236 12308 36242
rect 12256 36178 12308 36184
rect 12452 36174 12480 36654
rect 12440 36168 12492 36174
rect 12440 36110 12492 36116
rect 11888 35012 11940 35018
rect 11888 34954 11940 34960
rect 11900 34542 11928 34954
rect 11888 34536 11940 34542
rect 11888 34478 11940 34484
rect 11796 34060 11848 34066
rect 11796 34002 11848 34008
rect 12452 33930 12480 36110
rect 12532 35624 12584 35630
rect 12532 35566 12584 35572
rect 12544 34542 12572 35566
rect 12624 35148 12676 35154
rect 12624 35090 12676 35096
rect 12532 34536 12584 34542
rect 12532 34478 12584 34484
rect 12636 34202 12664 35090
rect 12624 34196 12676 34202
rect 12624 34138 12676 34144
rect 12440 33924 12492 33930
rect 12440 33866 12492 33872
rect 12348 32972 12400 32978
rect 12452 32960 12480 33866
rect 12636 33522 12664 34138
rect 12624 33516 12676 33522
rect 12624 33458 12676 33464
rect 12400 32932 12480 32960
rect 12348 32914 12400 32920
rect 12256 32904 12308 32910
rect 12256 32846 12308 32852
rect 12268 32502 12296 32846
rect 12256 32496 12308 32502
rect 12256 32438 12308 32444
rect 12072 31816 12124 31822
rect 12072 31758 12124 31764
rect 12716 31816 12768 31822
rect 12716 31758 12768 31764
rect 12084 31142 12112 31758
rect 12532 31680 12584 31686
rect 12532 31622 12584 31628
rect 12072 31136 12124 31142
rect 12072 31078 12124 31084
rect 12544 30190 12572 31622
rect 12728 30598 12756 31758
rect 12716 30592 12768 30598
rect 12716 30534 12768 30540
rect 12624 30320 12676 30326
rect 12624 30262 12676 30268
rect 11612 30184 11664 30190
rect 11612 30126 11664 30132
rect 12532 30184 12584 30190
rect 12532 30126 12584 30132
rect 11060 30116 11112 30122
rect 11060 30058 11112 30064
rect 10692 29096 10744 29102
rect 10692 29038 10744 29044
rect 9956 28620 10008 28626
rect 9956 28562 10008 28568
rect 10324 28620 10376 28626
rect 10324 28562 10376 28568
rect 10600 28620 10652 28626
rect 10600 28562 10652 28568
rect 9588 28144 9640 28150
rect 9588 28086 9640 28092
rect 9680 28144 9732 28150
rect 9680 28086 9732 28092
rect 9600 27996 9628 28086
rect 9692 27996 9720 28086
rect 9968 28082 9996 28562
rect 10612 28082 10640 28562
rect 9956 28076 10008 28082
rect 9956 28018 10008 28024
rect 10600 28076 10652 28082
rect 10600 28018 10652 28024
rect 9600 27968 9720 27996
rect 9772 28008 9824 28014
rect 9772 27950 9824 27956
rect 9784 27334 9812 27950
rect 11072 27878 11100 30058
rect 11612 30048 11664 30054
rect 11612 29990 11664 29996
rect 12348 30048 12400 30054
rect 12348 29990 12400 29996
rect 11336 29640 11388 29646
rect 11336 29582 11388 29588
rect 11348 28082 11376 29582
rect 11624 28762 11652 29990
rect 12360 29714 12388 29990
rect 12636 29850 12664 30262
rect 12624 29844 12676 29850
rect 12624 29786 12676 29792
rect 12348 29708 12400 29714
rect 12348 29650 12400 29656
rect 12728 29238 12756 30534
rect 12716 29232 12768 29238
rect 12716 29174 12768 29180
rect 12164 29164 12216 29170
rect 12164 29106 12216 29112
rect 11612 28756 11664 28762
rect 11612 28698 11664 28704
rect 11428 28688 11480 28694
rect 11428 28630 11480 28636
rect 11336 28076 11388 28082
rect 11336 28018 11388 28024
rect 11440 28014 11468 28630
rect 11624 28626 11652 28698
rect 11612 28620 11664 28626
rect 11612 28562 11664 28568
rect 12176 28490 12204 29106
rect 12716 29096 12768 29102
rect 12716 29038 12768 29044
rect 12728 28626 12756 29038
rect 12716 28620 12768 28626
rect 12716 28562 12768 28568
rect 12164 28484 12216 28490
rect 12164 28426 12216 28432
rect 12440 28144 12492 28150
rect 12440 28086 12492 28092
rect 11428 28008 11480 28014
rect 11428 27950 11480 27956
rect 12072 28008 12124 28014
rect 12072 27950 12124 27956
rect 11060 27872 11112 27878
rect 11060 27814 11112 27820
rect 11152 27668 11204 27674
rect 11152 27610 11204 27616
rect 10324 27532 10376 27538
rect 10324 27474 10376 27480
rect 9772 27328 9824 27334
rect 9772 27270 9824 27276
rect 9220 26988 9272 26994
rect 9220 26930 9272 26936
rect 9312 26988 9364 26994
rect 9312 26930 9364 26936
rect 8576 26444 8628 26450
rect 8576 26386 8628 26392
rect 8760 26444 8812 26450
rect 8760 26386 8812 26392
rect 8852 26444 8904 26450
rect 8852 26386 8904 26392
rect 8588 25906 8616 26386
rect 8576 25900 8628 25906
rect 8628 25860 8708 25888
rect 8576 25842 8628 25848
rect 8576 25152 8628 25158
rect 8576 25094 8628 25100
rect 8588 23662 8616 25094
rect 8680 24886 8708 25860
rect 8772 25770 8800 26386
rect 8864 25838 8892 26386
rect 8852 25832 8904 25838
rect 8852 25774 8904 25780
rect 8760 25764 8812 25770
rect 8760 25706 8812 25712
rect 8668 24880 8720 24886
rect 8668 24822 8720 24828
rect 8680 24274 8708 24822
rect 8772 24342 8800 25706
rect 8760 24336 8812 24342
rect 8760 24278 8812 24284
rect 8668 24268 8720 24274
rect 8668 24210 8720 24216
rect 8576 23656 8628 23662
rect 8576 23598 8628 23604
rect 8484 23316 8536 23322
rect 8484 23258 8536 23264
rect 8588 22574 8616 23598
rect 8680 23526 8708 24210
rect 8668 23520 8720 23526
rect 8668 23462 8720 23468
rect 8668 23316 8720 23322
rect 8668 23258 8720 23264
rect 8576 22568 8628 22574
rect 8576 22510 8628 22516
rect 8588 22098 8616 22510
rect 8576 22092 8628 22098
rect 8576 22034 8628 22040
rect 8576 21684 8628 21690
rect 8576 21626 8628 21632
rect 8588 21418 8616 21626
rect 8576 21412 8628 21418
rect 8576 21354 8628 21360
rect 8588 21146 8616 21354
rect 8576 21140 8628 21146
rect 8576 21082 8628 21088
rect 8208 21072 8260 21078
rect 8208 21014 8260 21020
rect 8116 20392 8168 20398
rect 8116 20334 8168 20340
rect 8208 20392 8260 20398
rect 8208 20334 8260 20340
rect 8220 19514 8248 20334
rect 8392 19984 8444 19990
rect 8392 19926 8444 19932
rect 8208 19508 8260 19514
rect 8208 19450 8260 19456
rect 8024 19440 8076 19446
rect 7930 19408 7986 19417
rect 7986 19388 8024 19394
rect 7986 19382 8076 19388
rect 7986 19366 8064 19382
rect 7930 19343 7986 19352
rect 7840 17536 7892 17542
rect 7840 17478 7892 17484
rect 7748 17128 7800 17134
rect 7748 17070 7800 17076
rect 7760 16046 7788 17070
rect 7748 16040 7800 16046
rect 7748 15982 7800 15988
rect 7656 12980 7708 12986
rect 7656 12922 7708 12928
rect 7944 12594 7972 19343
rect 8404 19310 8432 19926
rect 8392 19304 8444 19310
rect 8392 19246 8444 19252
rect 8404 18834 8432 19246
rect 8392 18828 8444 18834
rect 8392 18770 8444 18776
rect 8392 18216 8444 18222
rect 8392 18158 8444 18164
rect 8404 17882 8432 18158
rect 8392 17876 8444 17882
rect 8392 17818 8444 17824
rect 8392 17740 8444 17746
rect 8392 17682 8444 17688
rect 8024 17128 8076 17134
rect 8024 17070 8076 17076
rect 8036 16794 8064 17070
rect 8024 16788 8076 16794
rect 8024 16730 8076 16736
rect 8404 16250 8432 17682
rect 8680 17202 8708 23258
rect 8772 22642 8800 24278
rect 8864 24206 8892 25774
rect 9220 24744 9272 24750
rect 9220 24686 9272 24692
rect 9128 24268 9180 24274
rect 9128 24210 9180 24216
rect 8852 24200 8904 24206
rect 8852 24142 8904 24148
rect 9140 24070 9168 24210
rect 9128 24064 9180 24070
rect 9128 24006 9180 24012
rect 9232 23866 9260 24686
rect 9220 23860 9272 23866
rect 9220 23802 9272 23808
rect 8852 23180 8904 23186
rect 8852 23122 8904 23128
rect 8760 22636 8812 22642
rect 8760 22578 8812 22584
rect 8760 22228 8812 22234
rect 8760 22170 8812 22176
rect 8772 19310 8800 22170
rect 8864 22166 8892 23122
rect 8852 22160 8904 22166
rect 8852 22102 8904 22108
rect 8944 21004 8996 21010
rect 8944 20946 8996 20952
rect 8956 20602 8984 20946
rect 9036 20868 9088 20874
rect 9036 20810 9088 20816
rect 8944 20596 8996 20602
rect 8944 20538 8996 20544
rect 8956 19990 8984 20538
rect 9048 20466 9076 20810
rect 9036 20460 9088 20466
rect 9036 20402 9088 20408
rect 8944 19984 8996 19990
rect 8944 19926 8996 19932
rect 9036 19916 9088 19922
rect 9036 19858 9088 19864
rect 8760 19304 8812 19310
rect 8760 19246 8812 19252
rect 9048 18834 9076 19858
rect 9036 18828 9088 18834
rect 9036 18770 9088 18776
rect 9048 18426 9076 18770
rect 9036 18420 9088 18426
rect 9036 18362 9088 18368
rect 8944 17604 8996 17610
rect 8944 17546 8996 17552
rect 8668 17196 8720 17202
rect 8668 17138 8720 17144
rect 8956 16794 8984 17546
rect 8944 16788 8996 16794
rect 8944 16730 8996 16736
rect 8392 16244 8444 16250
rect 8392 16186 8444 16192
rect 8024 14952 8076 14958
rect 8024 14894 8076 14900
rect 9036 14952 9088 14958
rect 9036 14894 9088 14900
rect 8036 14006 8064 14894
rect 8944 14476 8996 14482
rect 8944 14418 8996 14424
rect 8760 14408 8812 14414
rect 8760 14350 8812 14356
rect 8484 14340 8536 14346
rect 8484 14282 8536 14288
rect 8024 14000 8076 14006
rect 8024 13942 8076 13948
rect 8024 12776 8076 12782
rect 8024 12718 8076 12724
rect 7760 12566 7972 12594
rect 7760 12322 7788 12566
rect 7668 12294 7788 12322
rect 7564 11212 7616 11218
rect 7564 11154 7616 11160
rect 7288 10532 7340 10538
rect 7288 10474 7340 10480
rect 7300 9722 7328 10474
rect 7288 9716 7340 9722
rect 7288 9658 7340 9664
rect 7012 9648 7064 9654
rect 7012 9590 7064 9596
rect 7104 9376 7156 9382
rect 7104 9318 7156 9324
rect 7012 9036 7064 9042
rect 7012 8978 7064 8984
rect 6920 8628 6972 8634
rect 6920 8570 6972 8576
rect 6564 8078 6776 8106
rect 6460 7812 6512 7818
rect 6460 7754 6512 7760
rect 6092 7336 6144 7342
rect 6092 7278 6144 7284
rect 6184 7200 6236 7206
rect 6184 7142 6236 7148
rect 6196 6798 6224 7142
rect 6184 6792 6236 6798
rect 6184 6734 6236 6740
rect 6460 6792 6512 6798
rect 6460 6734 6512 6740
rect 6000 6248 6052 6254
rect 6000 6190 6052 6196
rect 5908 6180 5960 6186
rect 5908 6122 5960 6128
rect 6000 6112 6052 6118
rect 6000 6054 6052 6060
rect 6012 5778 6040 6054
rect 6196 5846 6224 6734
rect 6472 6322 6500 6734
rect 6460 6316 6512 6322
rect 6460 6258 6512 6264
rect 6184 5840 6236 5846
rect 6184 5782 6236 5788
rect 6000 5772 6052 5778
rect 6000 5714 6052 5720
rect 5816 5160 5868 5166
rect 5816 5102 5868 5108
rect 5264 5024 5316 5030
rect 5264 4966 5316 4972
rect 5276 4690 5304 4966
rect 5264 4684 5316 4690
rect 5264 4626 5316 4632
rect 5448 4616 5500 4622
rect 5448 4558 5500 4564
rect 4804 3936 4856 3942
rect 4804 3878 4856 3884
rect 5172 3936 5224 3942
rect 5172 3878 5224 3884
rect 4068 3528 4120 3534
rect 4068 3470 4120 3476
rect 4712 3528 4764 3534
rect 4712 3470 4764 3476
rect 4080 3194 4108 3470
rect 4220 3292 4516 3312
rect 4276 3290 4300 3292
rect 4356 3290 4380 3292
rect 4436 3290 4460 3292
rect 4298 3238 4300 3290
rect 4362 3238 4374 3290
rect 4436 3238 4438 3290
rect 4276 3236 4300 3238
rect 4356 3236 4380 3238
rect 4436 3236 4460 3238
rect 4220 3216 4516 3236
rect 3792 3188 3844 3194
rect 3792 3130 3844 3136
rect 4068 3188 4120 3194
rect 4068 3130 4120 3136
rect 2872 3052 2924 3058
rect 2872 2994 2924 3000
rect 2596 2984 2648 2990
rect 2596 2926 2648 2932
rect 2608 2514 2636 2926
rect 4620 2916 4672 2922
rect 4620 2858 4672 2864
rect 1952 2508 2004 2514
rect 1952 2450 2004 2456
rect 2596 2508 2648 2514
rect 2596 2450 2648 2456
rect 2596 2304 2648 2310
rect 2596 2246 2648 2252
rect 2608 800 2636 2246
rect 4220 2204 4516 2224
rect 4276 2202 4300 2204
rect 4356 2202 4380 2204
rect 4436 2202 4460 2204
rect 4298 2150 4300 2202
rect 4362 2150 4374 2202
rect 4436 2150 4438 2202
rect 4276 2148 4300 2150
rect 4356 2148 4380 2150
rect 4436 2148 4460 2150
rect 4220 2128 4516 2148
rect 4632 800 4660 2858
rect 4724 2514 4752 3470
rect 4816 2854 4844 3878
rect 5184 3670 5212 3878
rect 5172 3664 5224 3670
rect 5172 3606 5224 3612
rect 5460 3602 5488 4558
rect 5828 3602 5856 5102
rect 6196 4690 6224 5782
rect 6368 4752 6420 4758
rect 6564 4706 6592 8078
rect 6644 7948 6696 7954
rect 6644 7890 6696 7896
rect 6656 5574 6684 7890
rect 6736 7880 6788 7886
rect 6736 7822 6788 7828
rect 6748 6866 6776 7822
rect 7024 7002 7052 8978
rect 7012 6996 7064 7002
rect 7012 6938 7064 6944
rect 6736 6860 6788 6866
rect 6736 6802 6788 6808
rect 7024 6254 7052 6938
rect 7012 6248 7064 6254
rect 7012 6190 7064 6196
rect 6828 6112 6880 6118
rect 6828 6054 6880 6060
rect 6840 5846 6868 6054
rect 6828 5840 6880 5846
rect 6828 5782 6880 5788
rect 6644 5568 6696 5574
rect 6644 5510 6696 5516
rect 6840 5030 6868 5782
rect 7012 5160 7064 5166
rect 7012 5102 7064 5108
rect 6828 5024 6880 5030
rect 6828 4966 6880 4972
rect 6420 4700 6592 4706
rect 6368 4694 6592 4700
rect 6184 4684 6236 4690
rect 6380 4678 6592 4694
rect 6840 4690 6868 4966
rect 6184 4626 6236 4632
rect 6564 3738 6592 4678
rect 6828 4684 6880 4690
rect 6828 4626 6880 4632
rect 7024 4282 7052 5102
rect 7012 4276 7064 4282
rect 7012 4218 7064 4224
rect 6920 4072 6972 4078
rect 6920 4014 6972 4020
rect 6552 3732 6604 3738
rect 6552 3674 6604 3680
rect 5448 3596 5500 3602
rect 5448 3538 5500 3544
rect 5816 3596 5868 3602
rect 5816 3538 5868 3544
rect 5724 2984 5776 2990
rect 5828 2972 5856 3538
rect 6932 3534 6960 4014
rect 6920 3528 6972 3534
rect 6920 3470 6972 3476
rect 6828 3460 6880 3466
rect 6828 3402 6880 3408
rect 6840 2990 6868 3402
rect 7116 2990 7144 9318
rect 7300 6202 7328 9658
rect 7380 8832 7432 8838
rect 7380 8774 7432 8780
rect 7392 8430 7420 8774
rect 7380 8424 7432 8430
rect 7380 8366 7432 8372
rect 7392 7886 7420 8366
rect 7380 7880 7432 7886
rect 7380 7822 7432 7828
rect 7392 7342 7420 7822
rect 7380 7336 7432 7342
rect 7380 7278 7432 7284
rect 7392 7018 7420 7278
rect 7392 6990 7512 7018
rect 7484 6934 7512 6990
rect 7472 6928 7524 6934
rect 7472 6870 7524 6876
rect 7472 6248 7524 6254
rect 7300 6174 7420 6202
rect 7472 6190 7524 6196
rect 7288 6112 7340 6118
rect 7288 6054 7340 6060
rect 7196 5704 7248 5710
rect 7196 5646 7248 5652
rect 7208 4146 7236 5646
rect 7300 5642 7328 6054
rect 7288 5636 7340 5642
rect 7288 5578 7340 5584
rect 7300 5302 7328 5578
rect 7288 5296 7340 5302
rect 7288 5238 7340 5244
rect 7392 5234 7420 6174
rect 7484 5574 7512 6190
rect 7472 5568 7524 5574
rect 7472 5510 7524 5516
rect 7380 5228 7432 5234
rect 7380 5170 7432 5176
rect 7196 4140 7248 4146
rect 7196 4082 7248 4088
rect 7392 3942 7420 5170
rect 7484 5166 7512 5510
rect 7472 5160 7524 5166
rect 7472 5102 7524 5108
rect 7484 4690 7512 5102
rect 7472 4684 7524 4690
rect 7472 4626 7524 4632
rect 7380 3936 7432 3942
rect 7380 3878 7432 3884
rect 7392 3534 7420 3878
rect 7472 3596 7524 3602
rect 7472 3538 7524 3544
rect 7380 3528 7432 3534
rect 7380 3470 7432 3476
rect 7484 3194 7512 3538
rect 7472 3188 7524 3194
rect 7472 3130 7524 3136
rect 7564 3052 7616 3058
rect 7564 2994 7616 3000
rect 5776 2944 5856 2972
rect 6644 2984 6696 2990
rect 5724 2926 5776 2932
rect 6644 2926 6696 2932
rect 6828 2984 6880 2990
rect 6828 2926 6880 2932
rect 7104 2984 7156 2990
rect 7104 2926 7156 2932
rect 7196 2984 7248 2990
rect 7196 2926 7248 2932
rect 4804 2848 4856 2854
rect 4804 2790 4856 2796
rect 6656 2650 6684 2926
rect 7208 2854 7236 2926
rect 7196 2848 7248 2854
rect 7196 2790 7248 2796
rect 7472 2848 7524 2854
rect 7472 2790 7524 2796
rect 6644 2644 6696 2650
rect 6644 2586 6696 2592
rect 4712 2508 4764 2514
rect 4712 2450 4764 2456
rect 6656 800 6684 2586
rect 7484 2582 7512 2790
rect 7472 2576 7524 2582
rect 7472 2518 7524 2524
rect 7576 2514 7604 2994
rect 6920 2508 6972 2514
rect 6920 2450 6972 2456
rect 7564 2508 7616 2514
rect 7564 2450 7616 2456
rect 6932 2038 6960 2450
rect 7668 2310 7696 12294
rect 8036 12238 8064 12718
rect 8300 12708 8352 12714
rect 8300 12650 8352 12656
rect 8024 12232 8076 12238
rect 8024 12174 8076 12180
rect 8036 11370 8064 12174
rect 8312 11898 8340 12650
rect 8392 12096 8444 12102
rect 8392 12038 8444 12044
rect 8300 11892 8352 11898
rect 8300 11834 8352 11840
rect 8404 11694 8432 12038
rect 8392 11688 8444 11694
rect 8392 11630 8444 11636
rect 8116 11552 8168 11558
rect 8116 11494 8168 11500
rect 7944 11354 8064 11370
rect 8128 11354 8156 11494
rect 7932 11348 8064 11354
rect 7984 11342 8064 11348
rect 8116 11348 8168 11354
rect 7932 11290 7984 11296
rect 8116 11290 8168 11296
rect 7944 9654 7972 11290
rect 8300 10600 8352 10606
rect 8300 10542 8352 10548
rect 8312 10266 8340 10542
rect 8392 10532 8444 10538
rect 8392 10474 8444 10480
rect 8300 10260 8352 10266
rect 8300 10202 8352 10208
rect 7932 9648 7984 9654
rect 7932 9590 7984 9596
rect 7840 9512 7892 9518
rect 7840 9454 7892 9460
rect 7852 8090 7880 9454
rect 7840 8084 7892 8090
rect 7840 8026 7892 8032
rect 7748 7948 7800 7954
rect 7748 7890 7800 7896
rect 7760 7478 7788 7890
rect 7748 7472 7800 7478
rect 7748 7414 7800 7420
rect 7852 7342 7880 8026
rect 7944 7954 7972 9590
rect 8300 9036 8352 9042
rect 8300 8978 8352 8984
rect 8312 8566 8340 8978
rect 8300 8560 8352 8566
rect 8300 8502 8352 8508
rect 7932 7948 7984 7954
rect 7932 7890 7984 7896
rect 7932 7404 7984 7410
rect 7932 7346 7984 7352
rect 7840 7336 7892 7342
rect 7840 7278 7892 7284
rect 7944 6322 7972 7346
rect 7932 6316 7984 6322
rect 7932 6258 7984 6264
rect 8312 5778 8340 8502
rect 8404 8090 8432 10474
rect 8392 8084 8444 8090
rect 8392 8026 8444 8032
rect 8392 7880 8444 7886
rect 8392 7822 8444 7828
rect 8404 7750 8432 7822
rect 8392 7744 8444 7750
rect 8392 7686 8444 7692
rect 8496 5778 8524 14282
rect 8668 13388 8720 13394
rect 8668 13330 8720 13336
rect 8576 11688 8628 11694
rect 8576 11630 8628 11636
rect 8588 10266 8616 11630
rect 8680 10810 8708 13330
rect 8772 12889 8800 14350
rect 8956 14074 8984 14418
rect 8944 14068 8996 14074
rect 8944 14010 8996 14016
rect 8758 12880 8814 12889
rect 8758 12815 8814 12824
rect 8772 12782 8800 12815
rect 8760 12776 8812 12782
rect 8760 12718 8812 12724
rect 9048 12306 9076 14894
rect 9232 14346 9260 23802
rect 9324 23186 9352 26930
rect 9680 26920 9732 26926
rect 9680 26862 9732 26868
rect 9692 25294 9720 26862
rect 10336 26858 10364 27474
rect 10324 26852 10376 26858
rect 10324 26794 10376 26800
rect 9864 26240 9916 26246
rect 9864 26182 9916 26188
rect 9876 25838 9904 26182
rect 9864 25832 9916 25838
rect 9864 25774 9916 25780
rect 9680 25288 9732 25294
rect 9732 25248 9812 25276
rect 9680 25230 9732 25236
rect 9784 24954 9812 25248
rect 9772 24948 9824 24954
rect 9772 24890 9824 24896
rect 9496 24676 9548 24682
rect 9496 24618 9548 24624
rect 9508 24274 9536 24618
rect 9496 24268 9548 24274
rect 9496 24210 9548 24216
rect 9588 24200 9640 24206
rect 9588 24142 9640 24148
rect 9404 23248 9456 23254
rect 9404 23190 9456 23196
rect 9312 23180 9364 23186
rect 9312 23122 9364 23128
rect 9416 22574 9444 23190
rect 9600 22574 9628 24142
rect 9680 22704 9732 22710
rect 9680 22646 9732 22652
rect 9404 22568 9456 22574
rect 9404 22510 9456 22516
rect 9588 22568 9640 22574
rect 9588 22510 9640 22516
rect 9416 21622 9444 22510
rect 9496 22092 9548 22098
rect 9496 22034 9548 22040
rect 9508 21865 9536 22034
rect 9494 21856 9550 21865
rect 9494 21791 9550 21800
rect 9404 21616 9456 21622
rect 9404 21558 9456 21564
rect 9692 21554 9720 22646
rect 9784 21962 9812 24890
rect 9876 23730 9904 25774
rect 9956 25288 10008 25294
rect 9956 25230 10008 25236
rect 9968 24274 9996 25230
rect 10048 24744 10100 24750
rect 10048 24686 10100 24692
rect 9956 24268 10008 24274
rect 9956 24210 10008 24216
rect 10060 24154 10088 24686
rect 9968 24126 10088 24154
rect 9864 23724 9916 23730
rect 9864 23666 9916 23672
rect 9968 23594 9996 24126
rect 10336 23730 10364 26794
rect 11164 26790 11192 27610
rect 11796 27532 11848 27538
rect 11796 27474 11848 27480
rect 11704 27396 11756 27402
rect 11704 27338 11756 27344
rect 11716 26926 11744 27338
rect 11808 27062 11836 27474
rect 11796 27056 11848 27062
rect 11796 26998 11848 27004
rect 11244 26920 11296 26926
rect 11244 26862 11296 26868
rect 11704 26920 11756 26926
rect 11704 26862 11756 26868
rect 11152 26784 11204 26790
rect 11152 26726 11204 26732
rect 11164 26518 11192 26726
rect 11152 26512 11204 26518
rect 11152 26454 11204 26460
rect 10784 26444 10836 26450
rect 10784 26386 10836 26392
rect 10796 24750 10824 26386
rect 11256 25770 11284 26862
rect 11888 26512 11940 26518
rect 11888 26454 11940 26460
rect 11704 26444 11756 26450
rect 11704 26386 11756 26392
rect 11244 25764 11296 25770
rect 11244 25706 11296 25712
rect 11612 25764 11664 25770
rect 11612 25706 11664 25712
rect 11060 25696 11112 25702
rect 11060 25638 11112 25644
rect 11152 25696 11204 25702
rect 11152 25638 11204 25644
rect 11072 25158 11100 25638
rect 11164 25498 11192 25638
rect 11152 25492 11204 25498
rect 11152 25434 11204 25440
rect 11060 25152 11112 25158
rect 11060 25094 11112 25100
rect 11164 24970 11192 25434
rect 11256 25430 11284 25706
rect 11244 25424 11296 25430
rect 11244 25366 11296 25372
rect 11624 25362 11652 25706
rect 11612 25356 11664 25362
rect 11612 25298 11664 25304
rect 11612 25152 11664 25158
rect 11612 25094 11664 25100
rect 10980 24942 11192 24970
rect 10784 24744 10836 24750
rect 10784 24686 10836 24692
rect 10692 24676 10744 24682
rect 10692 24618 10744 24624
rect 10508 24268 10560 24274
rect 10508 24210 10560 24216
rect 10520 24070 10548 24210
rect 10508 24064 10560 24070
rect 10508 24006 10560 24012
rect 10704 23730 10732 24618
rect 10324 23724 10376 23730
rect 10692 23724 10744 23730
rect 10376 23684 10456 23712
rect 10324 23666 10376 23672
rect 9956 23588 10008 23594
rect 9956 23530 10008 23536
rect 9968 23050 9996 23530
rect 10324 23112 10376 23118
rect 10324 23054 10376 23060
rect 9956 23044 10008 23050
rect 9956 22986 10008 22992
rect 10336 22574 10364 23054
rect 10048 22568 10100 22574
rect 10048 22510 10100 22516
rect 10324 22568 10376 22574
rect 10324 22510 10376 22516
rect 9864 22500 9916 22506
rect 9864 22442 9916 22448
rect 9772 21956 9824 21962
rect 9772 21898 9824 21904
rect 9680 21548 9732 21554
rect 9680 21490 9732 21496
rect 9784 21010 9812 21898
rect 9876 21486 9904 22442
rect 10060 22098 10088 22510
rect 10336 22166 10364 22510
rect 10428 22506 10456 23684
rect 10692 23666 10744 23672
rect 10980 23526 11008 24942
rect 11624 24750 11652 25094
rect 11612 24744 11664 24750
rect 11612 24686 11664 24692
rect 11716 24614 11744 26386
rect 11900 25702 11928 26454
rect 11888 25696 11940 25702
rect 11888 25638 11940 25644
rect 11980 25152 12032 25158
rect 11980 25094 12032 25100
rect 11992 24886 12020 25094
rect 11980 24880 12032 24886
rect 11980 24822 12032 24828
rect 12084 24750 12112 27950
rect 12452 27538 12480 28086
rect 12624 27600 12676 27606
rect 12624 27542 12676 27548
rect 12440 27532 12492 27538
rect 12492 27492 12572 27520
rect 12440 27474 12492 27480
rect 12544 26926 12572 27492
rect 12532 26920 12584 26926
rect 12532 26862 12584 26868
rect 12636 26586 12664 27542
rect 12728 27062 12756 28562
rect 12716 27056 12768 27062
rect 12716 26998 12768 27004
rect 12440 26580 12492 26586
rect 12440 26522 12492 26528
rect 12624 26580 12676 26586
rect 12624 26522 12676 26528
rect 12452 24818 12480 26522
rect 12532 26444 12584 26450
rect 12532 26386 12584 26392
rect 12544 25906 12572 26386
rect 12636 26042 12664 26522
rect 12624 26036 12676 26042
rect 12624 25978 12676 25984
rect 12532 25900 12584 25906
rect 12532 25842 12584 25848
rect 12624 25356 12676 25362
rect 12624 25298 12676 25304
rect 12636 24954 12664 25298
rect 12624 24948 12676 24954
rect 12624 24890 12676 24896
rect 12440 24812 12492 24818
rect 12440 24754 12492 24760
rect 12072 24744 12124 24750
rect 12072 24686 12124 24692
rect 11704 24608 11756 24614
rect 11704 24550 11756 24556
rect 11716 24342 11744 24550
rect 11060 24336 11112 24342
rect 11060 24278 11112 24284
rect 11704 24336 11756 24342
rect 11704 24278 11756 24284
rect 11072 23730 11100 24278
rect 12084 24206 12112 24686
rect 11704 24200 11756 24206
rect 11704 24142 11756 24148
rect 12072 24200 12124 24206
rect 12072 24142 12124 24148
rect 12164 24200 12216 24206
rect 12164 24142 12216 24148
rect 11060 23724 11112 23730
rect 11060 23666 11112 23672
rect 11716 23662 11744 24142
rect 11152 23656 11204 23662
rect 11152 23598 11204 23604
rect 11704 23656 11756 23662
rect 11704 23598 11756 23604
rect 10968 23520 11020 23526
rect 10968 23462 11020 23468
rect 11164 23118 11192 23598
rect 12176 23186 12204 24142
rect 12532 24132 12584 24138
rect 12532 24074 12584 24080
rect 12544 23662 12572 24074
rect 12624 23724 12676 23730
rect 12624 23666 12676 23672
rect 12532 23656 12584 23662
rect 12532 23598 12584 23604
rect 12532 23248 12584 23254
rect 12532 23190 12584 23196
rect 12164 23180 12216 23186
rect 12164 23122 12216 23128
rect 11152 23112 11204 23118
rect 11152 23054 11204 23060
rect 12176 22574 12204 23122
rect 12544 22574 12572 23190
rect 12636 23186 12664 23666
rect 12624 23180 12676 23186
rect 12624 23122 12676 23128
rect 12716 22976 12768 22982
rect 12716 22918 12768 22924
rect 11336 22568 11388 22574
rect 11336 22510 11388 22516
rect 12164 22568 12216 22574
rect 12532 22568 12584 22574
rect 12216 22528 12296 22556
rect 12164 22510 12216 22516
rect 10416 22500 10468 22506
rect 10416 22442 10468 22448
rect 10324 22160 10376 22166
rect 10324 22102 10376 22108
rect 10428 22098 10456 22442
rect 10048 22092 10100 22098
rect 10048 22034 10100 22040
rect 10416 22092 10468 22098
rect 10416 22034 10468 22040
rect 10600 22024 10652 22030
rect 10600 21966 10652 21972
rect 10612 21486 10640 21966
rect 11348 21486 11376 22510
rect 12268 22234 12296 22528
rect 12452 22528 12532 22556
rect 12452 22250 12480 22528
rect 12532 22510 12584 22516
rect 12532 22432 12584 22438
rect 12584 22380 12664 22386
rect 12532 22374 12664 22380
rect 12544 22358 12664 22374
rect 12256 22228 12308 22234
rect 12452 22222 12572 22250
rect 12256 22170 12308 22176
rect 12438 22128 12494 22137
rect 12438 22063 12494 22072
rect 9864 21480 9916 21486
rect 9864 21422 9916 21428
rect 10600 21480 10652 21486
rect 10600 21422 10652 21428
rect 11336 21480 11388 21486
rect 11336 21422 11388 21428
rect 11348 21146 11376 21422
rect 11336 21140 11388 21146
rect 11336 21082 11388 21088
rect 9772 21004 9824 21010
rect 9772 20946 9824 20952
rect 9496 20936 9548 20942
rect 9496 20878 9548 20884
rect 9508 20466 9536 20878
rect 12452 20534 12480 22063
rect 12544 21622 12572 22222
rect 12636 22098 12664 22358
rect 12624 22092 12676 22098
rect 12624 22034 12676 22040
rect 12728 22030 12756 22918
rect 12716 22024 12768 22030
rect 12716 21966 12768 21972
rect 12532 21616 12584 21622
rect 12532 21558 12584 21564
rect 12532 21344 12584 21350
rect 12532 21286 12584 21292
rect 12544 21010 12572 21286
rect 12532 21004 12584 21010
rect 12532 20946 12584 20952
rect 12440 20528 12492 20534
rect 12440 20470 12492 20476
rect 9496 20460 9548 20466
rect 9496 20402 9548 20408
rect 11428 20392 11480 20398
rect 11428 20334 11480 20340
rect 12532 20392 12584 20398
rect 12532 20334 12584 20340
rect 11440 20058 11468 20334
rect 12440 20256 12492 20262
rect 12440 20198 12492 20204
rect 11428 20052 11480 20058
rect 11428 19994 11480 20000
rect 11888 20052 11940 20058
rect 11888 19994 11940 20000
rect 11900 19922 11928 19994
rect 11888 19916 11940 19922
rect 11888 19858 11940 19864
rect 12348 19916 12400 19922
rect 12348 19858 12400 19864
rect 11060 19848 11112 19854
rect 11060 19790 11112 19796
rect 9680 19712 9732 19718
rect 9680 19654 9732 19660
rect 9692 18834 9720 19654
rect 11072 19514 11100 19790
rect 11060 19508 11112 19514
rect 11060 19450 11112 19456
rect 10600 19304 10652 19310
rect 10600 19246 10652 19252
rect 11612 19304 11664 19310
rect 11612 19246 11664 19252
rect 10232 19168 10284 19174
rect 10232 19110 10284 19116
rect 10244 18834 10272 19110
rect 9680 18828 9732 18834
rect 9680 18770 9732 18776
rect 10232 18828 10284 18834
rect 10232 18770 10284 18776
rect 10612 18766 10640 19246
rect 10600 18760 10652 18766
rect 10600 18702 10652 18708
rect 11244 18760 11296 18766
rect 11244 18702 11296 18708
rect 9772 18624 9824 18630
rect 9772 18566 9824 18572
rect 11152 18624 11204 18630
rect 11152 18566 11204 18572
rect 9784 17746 9812 18566
rect 11164 18290 11192 18566
rect 11152 18284 11204 18290
rect 11152 18226 11204 18232
rect 10140 18216 10192 18222
rect 10140 18158 10192 18164
rect 9772 17740 9824 17746
rect 9772 17682 9824 17688
rect 10152 17678 10180 18158
rect 11256 18154 11284 18702
rect 11336 18692 11388 18698
rect 11336 18634 11388 18640
rect 11348 18290 11376 18634
rect 11624 18426 11652 19246
rect 11900 18834 11928 19858
rect 11704 18828 11756 18834
rect 11704 18770 11756 18776
rect 11888 18828 11940 18834
rect 11888 18770 11940 18776
rect 11612 18420 11664 18426
rect 11612 18362 11664 18368
rect 11336 18284 11388 18290
rect 11336 18226 11388 18232
rect 11244 18148 11296 18154
rect 11244 18090 11296 18096
rect 9680 17672 9732 17678
rect 9680 17614 9732 17620
rect 10140 17672 10192 17678
rect 10140 17614 10192 17620
rect 9692 16590 9720 17614
rect 10692 17196 10744 17202
rect 10692 17138 10744 17144
rect 9864 17128 9916 17134
rect 9864 17070 9916 17076
rect 9772 16992 9824 16998
rect 9772 16934 9824 16940
rect 9784 16658 9812 16934
rect 9772 16652 9824 16658
rect 9772 16594 9824 16600
rect 9680 16584 9732 16590
rect 9680 16526 9732 16532
rect 9496 16040 9548 16046
rect 9496 15982 9548 15988
rect 9508 15570 9536 15982
rect 9876 15910 9904 17070
rect 10704 16114 10732 17138
rect 11060 17128 11112 17134
rect 11060 17070 11112 17076
rect 11072 16590 11100 17070
rect 11244 16720 11296 16726
rect 11244 16662 11296 16668
rect 11060 16584 11112 16590
rect 11060 16526 11112 16532
rect 11256 16250 11284 16662
rect 11428 16652 11480 16658
rect 11428 16594 11480 16600
rect 11244 16244 11296 16250
rect 11244 16186 11296 16192
rect 10692 16108 10744 16114
rect 10692 16050 10744 16056
rect 11256 16046 11284 16186
rect 10508 16040 10560 16046
rect 10428 16000 10508 16028
rect 9864 15904 9916 15910
rect 9864 15846 9916 15852
rect 9588 15700 9640 15706
rect 9588 15642 9640 15648
rect 9496 15564 9548 15570
rect 9496 15506 9548 15512
rect 9508 14822 9536 15506
rect 9600 14958 9628 15642
rect 9680 15496 9732 15502
rect 9680 15438 9732 15444
rect 9588 14952 9640 14958
rect 9588 14894 9640 14900
rect 9496 14816 9548 14822
rect 9496 14758 9548 14764
rect 9588 14816 9640 14822
rect 9588 14758 9640 14764
rect 9220 14340 9272 14346
rect 9220 14282 9272 14288
rect 9508 13682 9536 14758
rect 9600 13870 9628 14758
rect 9692 14346 9720 15438
rect 9876 15201 9904 15846
rect 10140 15700 10192 15706
rect 10140 15642 10192 15648
rect 9862 15192 9918 15201
rect 9862 15127 9918 15136
rect 10152 14958 10180 15642
rect 10232 15088 10284 15094
rect 10232 15030 10284 15036
rect 10140 14952 10192 14958
rect 10140 14894 10192 14900
rect 9772 14884 9824 14890
rect 9772 14826 9824 14832
rect 9680 14340 9732 14346
rect 9680 14282 9732 14288
rect 9784 13938 9812 14826
rect 10244 14482 10272 15030
rect 9956 14476 10008 14482
rect 9956 14418 10008 14424
rect 10232 14476 10284 14482
rect 10232 14418 10284 14424
rect 9864 14408 9916 14414
rect 9864 14350 9916 14356
rect 9772 13932 9824 13938
rect 9772 13874 9824 13880
rect 9588 13864 9640 13870
rect 9588 13806 9640 13812
rect 9508 13654 9720 13682
rect 9692 13394 9720 13654
rect 9680 13388 9732 13394
rect 9680 13330 9732 13336
rect 9404 13184 9456 13190
rect 9404 13126 9456 13132
rect 9416 12986 9444 13126
rect 9404 12980 9456 12986
rect 9404 12922 9456 12928
rect 9416 12782 9444 12922
rect 9404 12776 9456 12782
rect 9404 12718 9456 12724
rect 9416 12374 9444 12718
rect 9496 12708 9548 12714
rect 9496 12650 9548 12656
rect 9404 12368 9456 12374
rect 9404 12310 9456 12316
rect 9036 12300 9088 12306
rect 9036 12242 9088 12248
rect 8944 11756 8996 11762
rect 8944 11698 8996 11704
rect 8956 11218 8984 11698
rect 9128 11688 9180 11694
rect 9128 11630 9180 11636
rect 8944 11212 8996 11218
rect 8944 11154 8996 11160
rect 8668 10804 8720 10810
rect 8668 10746 8720 10752
rect 8576 10260 8628 10266
rect 8576 10202 8628 10208
rect 8588 10062 8616 10202
rect 8576 10056 8628 10062
rect 8576 9998 8628 10004
rect 8576 9172 8628 9178
rect 8576 9114 8628 9120
rect 8588 8430 8616 9114
rect 8680 8838 8708 10746
rect 8944 10124 8996 10130
rect 8944 10066 8996 10072
rect 8852 9512 8904 9518
rect 8852 9454 8904 9460
rect 8668 8832 8720 8838
rect 8668 8774 8720 8780
rect 8576 8424 8628 8430
rect 8576 8366 8628 8372
rect 8574 8120 8630 8129
rect 8574 8055 8630 8064
rect 8588 7954 8616 8055
rect 8576 7948 8628 7954
rect 8576 7890 8628 7896
rect 8760 7948 8812 7954
rect 8760 7890 8812 7896
rect 8772 7750 8800 7890
rect 8864 7818 8892 9454
rect 8852 7812 8904 7818
rect 8852 7754 8904 7760
rect 8760 7744 8812 7750
rect 8760 7686 8812 7692
rect 8864 7342 8892 7754
rect 8852 7336 8904 7342
rect 8852 7278 8904 7284
rect 8956 6730 8984 10066
rect 9036 9580 9088 9586
rect 9036 9522 9088 9528
rect 9048 8498 9076 9522
rect 9140 8974 9168 11630
rect 9508 10130 9536 12650
rect 9692 12306 9720 13330
rect 9784 12782 9812 13874
rect 9772 12776 9824 12782
rect 9772 12718 9824 12724
rect 9876 12442 9904 14350
rect 9968 13394 9996 14418
rect 10244 14226 10272 14418
rect 10244 14198 10364 14226
rect 9956 13388 10008 13394
rect 9956 13330 10008 13336
rect 10232 13388 10284 13394
rect 10232 13330 10284 13336
rect 9864 12436 9916 12442
rect 9864 12378 9916 12384
rect 9680 12300 9732 12306
rect 9680 12242 9732 12248
rect 9692 11914 9720 12242
rect 9692 11886 9812 11914
rect 9680 10600 9732 10606
rect 9680 10542 9732 10548
rect 9496 10124 9548 10130
rect 9496 10066 9548 10072
rect 9312 9920 9364 9926
rect 9312 9862 9364 9868
rect 9220 9036 9272 9042
rect 9220 8978 9272 8984
rect 9128 8968 9180 8974
rect 9128 8910 9180 8916
rect 9036 8492 9088 8498
rect 9036 8434 9088 8440
rect 9232 8294 9260 8978
rect 9220 8288 9272 8294
rect 9220 8230 9272 8236
rect 9232 7546 9260 8230
rect 9220 7540 9272 7546
rect 9220 7482 9272 7488
rect 8944 6724 8996 6730
rect 8944 6666 8996 6672
rect 8576 6452 8628 6458
rect 8576 6394 8628 6400
rect 8588 5914 8616 6394
rect 8576 5908 8628 5914
rect 8576 5850 8628 5856
rect 8300 5772 8352 5778
rect 8300 5714 8352 5720
rect 8484 5772 8536 5778
rect 8484 5714 8536 5720
rect 9036 5772 9088 5778
rect 9036 5714 9088 5720
rect 7840 4684 7892 4690
rect 7840 4626 7892 4632
rect 7852 4078 7880 4626
rect 7840 4072 7892 4078
rect 7840 4014 7892 4020
rect 7852 3126 7880 4014
rect 8668 3596 8720 3602
rect 8668 3538 8720 3544
rect 7932 3528 7984 3534
rect 7932 3470 7984 3476
rect 7840 3120 7892 3126
rect 7840 3062 7892 3068
rect 7656 2304 7708 2310
rect 7656 2246 7708 2252
rect 7944 2106 7972 3470
rect 8680 3194 8708 3538
rect 8668 3188 8720 3194
rect 8668 3130 8720 3136
rect 9048 2990 9076 5714
rect 9324 3534 9352 9862
rect 9496 9376 9548 9382
rect 9496 9318 9548 9324
rect 9508 9042 9536 9318
rect 9692 9110 9720 10542
rect 9784 9178 9812 11886
rect 9864 11756 9916 11762
rect 9864 11698 9916 11704
rect 9876 11014 9904 11698
rect 10244 11694 10272 13330
rect 10336 11694 10364 14198
rect 10428 12646 10456 16000
rect 10508 15982 10560 15988
rect 11244 16040 11296 16046
rect 11244 15982 11296 15988
rect 11440 15706 11468 16594
rect 11428 15700 11480 15706
rect 11428 15642 11480 15648
rect 11336 15360 11388 15366
rect 11336 15302 11388 15308
rect 10508 15020 10560 15026
rect 10508 14962 10560 14968
rect 10520 14482 10548 14962
rect 10876 14952 10928 14958
rect 10876 14894 10928 14900
rect 10888 14550 10916 14894
rect 10876 14544 10928 14550
rect 10876 14486 10928 14492
rect 10508 14476 10560 14482
rect 10508 14418 10560 14424
rect 10888 13938 10916 14486
rect 11348 14482 11376 15302
rect 11336 14476 11388 14482
rect 11336 14418 11388 14424
rect 11428 14340 11480 14346
rect 11428 14282 11480 14288
rect 11440 14006 11468 14282
rect 11428 14000 11480 14006
rect 11428 13942 11480 13948
rect 10876 13932 10928 13938
rect 10876 13874 10928 13880
rect 10692 13864 10744 13870
rect 10692 13806 10744 13812
rect 11060 13864 11112 13870
rect 11060 13806 11112 13812
rect 10704 13530 10732 13806
rect 10692 13524 10744 13530
rect 10692 13466 10744 13472
rect 10968 13524 11020 13530
rect 10968 13466 11020 13472
rect 10876 12844 10928 12850
rect 10876 12786 10928 12792
rect 10690 12744 10746 12753
rect 10690 12679 10746 12688
rect 10416 12640 10468 12646
rect 10416 12582 10468 12588
rect 9956 11688 10008 11694
rect 9956 11630 10008 11636
rect 10232 11688 10284 11694
rect 10232 11630 10284 11636
rect 10324 11688 10376 11694
rect 10324 11630 10376 11636
rect 9864 11008 9916 11014
rect 9864 10950 9916 10956
rect 9862 10432 9918 10441
rect 9862 10367 9918 10376
rect 9876 10130 9904 10367
rect 9864 10124 9916 10130
rect 9864 10066 9916 10072
rect 9968 9518 9996 11630
rect 10140 11552 10192 11558
rect 10140 11494 10192 11500
rect 10152 11286 10180 11494
rect 10140 11280 10192 11286
rect 10140 11222 10192 11228
rect 10152 10130 10180 11222
rect 10324 10736 10376 10742
rect 10324 10678 10376 10684
rect 10232 10532 10284 10538
rect 10232 10474 10284 10480
rect 10244 10130 10272 10474
rect 10336 10266 10364 10678
rect 10324 10260 10376 10266
rect 10324 10202 10376 10208
rect 10140 10124 10192 10130
rect 10140 10066 10192 10072
rect 10232 10124 10284 10130
rect 10232 10066 10284 10072
rect 9956 9512 10008 9518
rect 9956 9454 10008 9460
rect 9772 9172 9824 9178
rect 9772 9114 9824 9120
rect 9680 9104 9732 9110
rect 9680 9046 9732 9052
rect 9496 9036 9548 9042
rect 9496 8978 9548 8984
rect 9404 8016 9456 8022
rect 9404 7958 9456 7964
rect 9416 7410 9444 7958
rect 9404 7404 9456 7410
rect 9404 7346 9456 7352
rect 9508 6322 9536 8978
rect 10336 8974 10364 10202
rect 10428 9382 10456 12582
rect 10704 12442 10732 12679
rect 10888 12442 10916 12786
rect 10692 12436 10744 12442
rect 10692 12378 10744 12384
rect 10876 12436 10928 12442
rect 10876 12378 10928 12384
rect 10876 12232 10928 12238
rect 10876 12174 10928 12180
rect 10888 11830 10916 12174
rect 10692 11824 10744 11830
rect 10692 11766 10744 11772
rect 10876 11824 10928 11830
rect 10876 11766 10928 11772
rect 10600 11212 10652 11218
rect 10600 11154 10652 11160
rect 10508 11008 10560 11014
rect 10508 10950 10560 10956
rect 10520 10130 10548 10950
rect 10508 10124 10560 10130
rect 10508 10066 10560 10072
rect 10508 9580 10560 9586
rect 10508 9522 10560 9528
rect 10416 9376 10468 9382
rect 10416 9318 10468 9324
rect 10324 8968 10376 8974
rect 10324 8910 10376 8916
rect 9772 8900 9824 8906
rect 9772 8842 9824 8848
rect 9496 6316 9548 6322
rect 9496 6258 9548 6264
rect 9508 5846 9536 6258
rect 9680 6112 9732 6118
rect 9680 6054 9732 6060
rect 9496 5840 9548 5846
rect 9496 5782 9548 5788
rect 9508 5642 9536 5782
rect 9692 5778 9720 6054
rect 9680 5772 9732 5778
rect 9680 5714 9732 5720
rect 9496 5636 9548 5642
rect 9496 5578 9548 5584
rect 9784 4758 9812 8842
rect 10416 8424 10468 8430
rect 10416 8366 10468 8372
rect 10140 7948 10192 7954
rect 10140 7890 10192 7896
rect 10152 6866 10180 7890
rect 10428 7478 10456 8366
rect 10416 7472 10468 7478
rect 10416 7414 10468 7420
rect 10428 7274 10456 7414
rect 10520 7342 10548 9522
rect 10612 9466 10640 11154
rect 10704 11150 10732 11766
rect 10980 11218 11008 13466
rect 11072 12782 11100 13806
rect 11440 13258 11468 13942
rect 11428 13252 11480 13258
rect 11428 13194 11480 13200
rect 11244 12980 11296 12986
rect 11244 12922 11296 12928
rect 11336 12980 11388 12986
rect 11336 12922 11388 12928
rect 11152 12844 11204 12850
rect 11152 12786 11204 12792
rect 11060 12776 11112 12782
rect 11060 12718 11112 12724
rect 11060 12096 11112 12102
rect 11060 12038 11112 12044
rect 10968 11212 11020 11218
rect 10968 11154 11020 11160
rect 10692 11144 10744 11150
rect 10692 11086 10744 11092
rect 10704 10538 10732 11086
rect 11072 10849 11100 12038
rect 11164 11762 11192 12786
rect 11152 11756 11204 11762
rect 11152 11698 11204 11704
rect 11058 10840 11114 10849
rect 11058 10775 11114 10784
rect 10968 10600 11020 10606
rect 10968 10542 11020 10548
rect 10692 10532 10744 10538
rect 10692 10474 10744 10480
rect 10612 9438 10732 9466
rect 10600 9036 10652 9042
rect 10600 8978 10652 8984
rect 10508 7336 10560 7342
rect 10508 7278 10560 7284
rect 10416 7268 10468 7274
rect 10416 7210 10468 7216
rect 10140 6860 10192 6866
rect 10140 6802 10192 6808
rect 10232 6860 10284 6866
rect 10232 6802 10284 6808
rect 10152 6254 10180 6802
rect 10140 6248 10192 6254
rect 10140 6190 10192 6196
rect 10244 6118 10272 6802
rect 10508 6656 10560 6662
rect 10508 6598 10560 6604
rect 10232 6112 10284 6118
rect 10232 6054 10284 6060
rect 10244 5166 10272 6054
rect 10232 5160 10284 5166
rect 10232 5102 10284 5108
rect 10232 5024 10284 5030
rect 10232 4966 10284 4972
rect 9772 4752 9824 4758
rect 9692 4700 9772 4706
rect 9692 4694 9824 4700
rect 9692 4678 9812 4694
rect 10244 4690 10272 4966
rect 10232 4684 10284 4690
rect 9496 4616 9548 4622
rect 9496 4558 9548 4564
rect 9508 4214 9536 4558
rect 9496 4208 9548 4214
rect 9496 4150 9548 4156
rect 9312 3528 9364 3534
rect 9312 3470 9364 3476
rect 9036 2984 9088 2990
rect 9036 2926 9088 2932
rect 9324 2446 9352 3470
rect 9692 2514 9720 4678
rect 10232 4626 10284 4632
rect 10140 4548 10192 4554
rect 10140 4490 10192 4496
rect 9864 4072 9916 4078
rect 9864 4014 9916 4020
rect 9772 3664 9824 3670
rect 9876 3618 9904 4014
rect 9824 3612 9904 3618
rect 9772 3606 9904 3612
rect 9784 3590 9904 3606
rect 9876 2650 9904 3590
rect 10046 3088 10102 3097
rect 10046 3023 10048 3032
rect 10100 3023 10102 3032
rect 10048 2994 10100 3000
rect 10152 2990 10180 4490
rect 10244 4146 10272 4626
rect 10232 4140 10284 4146
rect 10232 4082 10284 4088
rect 10520 4078 10548 6598
rect 10612 6186 10640 8978
rect 10704 8514 10732 9438
rect 10784 9036 10836 9042
rect 10784 8978 10836 8984
rect 10796 8634 10824 8978
rect 10784 8628 10836 8634
rect 10784 8570 10836 8576
rect 10704 8486 10824 8514
rect 10796 7954 10824 8486
rect 10692 7948 10744 7954
rect 10692 7890 10744 7896
rect 10784 7948 10836 7954
rect 10784 7890 10836 7896
rect 10600 6180 10652 6186
rect 10600 6122 10652 6128
rect 10704 4690 10732 7890
rect 10980 6934 11008 10542
rect 11256 10452 11284 12922
rect 11348 12889 11376 12922
rect 11334 12880 11390 12889
rect 11334 12815 11390 12824
rect 11440 12782 11468 13194
rect 11428 12776 11480 12782
rect 11428 12718 11480 12724
rect 11336 12708 11388 12714
rect 11336 12650 11388 12656
rect 11348 12102 11376 12650
rect 11336 12096 11388 12102
rect 11336 12038 11388 12044
rect 11612 12096 11664 12102
rect 11612 12038 11664 12044
rect 11348 10606 11376 12038
rect 11520 11348 11572 11354
rect 11520 11290 11572 11296
rect 11532 10606 11560 11290
rect 11336 10600 11388 10606
rect 11336 10542 11388 10548
rect 11520 10600 11572 10606
rect 11520 10542 11572 10548
rect 11256 10424 11468 10452
rect 11336 10056 11388 10062
rect 11336 9998 11388 10004
rect 11152 9648 11204 9654
rect 11152 9590 11204 9596
rect 11164 8362 11192 9590
rect 11348 9518 11376 9998
rect 11336 9512 11388 9518
rect 11336 9454 11388 9460
rect 11336 8424 11388 8430
rect 11440 8412 11468 10424
rect 11520 9512 11572 9518
rect 11520 9454 11572 9460
rect 11388 8384 11468 8412
rect 11336 8366 11388 8372
rect 11152 8356 11204 8362
rect 11152 8298 11204 8304
rect 11348 7818 11376 8366
rect 11532 7970 11560 9454
rect 11624 8129 11652 12038
rect 11716 10033 11744 18770
rect 11900 17678 11928 18770
rect 12360 18426 12388 19858
rect 12452 19854 12480 20198
rect 12544 20058 12572 20334
rect 12532 20052 12584 20058
rect 12532 19994 12584 20000
rect 12440 19848 12492 19854
rect 12440 19790 12492 19796
rect 12452 19281 12480 19790
rect 12532 19712 12584 19718
rect 12532 19654 12584 19660
rect 12438 19272 12494 19281
rect 12438 19207 12494 19216
rect 12348 18420 12400 18426
rect 12348 18362 12400 18368
rect 12452 18222 12480 19207
rect 12544 18834 12572 19654
rect 12532 18828 12584 18834
rect 12532 18770 12584 18776
rect 12532 18420 12584 18426
rect 12532 18362 12584 18368
rect 12440 18216 12492 18222
rect 12440 18158 12492 18164
rect 12544 17746 12572 18362
rect 12624 18216 12676 18222
rect 12624 18158 12676 18164
rect 12636 17882 12664 18158
rect 12716 18080 12768 18086
rect 12716 18022 12768 18028
rect 12624 17876 12676 17882
rect 12624 17818 12676 17824
rect 12532 17740 12584 17746
rect 12532 17682 12584 17688
rect 11888 17672 11940 17678
rect 11888 17614 11940 17620
rect 12728 17542 12756 18022
rect 12716 17536 12768 17542
rect 12716 17478 12768 17484
rect 12728 17270 12756 17478
rect 12348 17264 12400 17270
rect 12348 17206 12400 17212
rect 12716 17264 12768 17270
rect 12716 17206 12768 17212
rect 11796 16516 11848 16522
rect 11796 16458 11848 16464
rect 11808 16250 11836 16458
rect 11796 16244 11848 16250
rect 11796 16186 11848 16192
rect 11808 10606 11836 16186
rect 12360 15910 12388 17206
rect 12624 17060 12676 17066
rect 12624 17002 12676 17008
rect 12440 16992 12492 16998
rect 12440 16934 12492 16940
rect 12452 16658 12480 16934
rect 12440 16652 12492 16658
rect 12440 16594 12492 16600
rect 12452 16046 12480 16594
rect 12636 16454 12664 17002
rect 12728 16658 12756 17206
rect 12820 16794 12848 36654
rect 13544 36236 13596 36242
rect 13544 36178 13596 36184
rect 15476 36236 15528 36242
rect 15476 36178 15528 36184
rect 15568 36236 15620 36242
rect 15568 36178 15620 36184
rect 13556 35630 13584 36178
rect 14188 36168 14240 36174
rect 14188 36110 14240 36116
rect 13912 36032 13964 36038
rect 13912 35974 13964 35980
rect 13544 35624 13596 35630
rect 13544 35566 13596 35572
rect 13360 35488 13412 35494
rect 13360 35430 13412 35436
rect 13372 35222 13400 35430
rect 13360 35216 13412 35222
rect 13360 35158 13412 35164
rect 13372 34542 13400 35158
rect 13556 35018 13584 35566
rect 13820 35556 13872 35562
rect 13820 35498 13872 35504
rect 13832 35154 13860 35498
rect 13820 35148 13872 35154
rect 13820 35090 13872 35096
rect 13924 35034 13952 35974
rect 14004 35624 14056 35630
rect 14004 35566 14056 35572
rect 13544 35012 13596 35018
rect 13544 34954 13596 34960
rect 13832 35006 13952 35034
rect 13832 34542 13860 35006
rect 14016 34542 14044 35566
rect 14200 35154 14228 36110
rect 14280 36032 14332 36038
rect 14280 35974 14332 35980
rect 14188 35148 14240 35154
rect 14188 35090 14240 35096
rect 14200 34542 14228 35090
rect 14292 34610 14320 35974
rect 14280 34604 14332 34610
rect 14280 34546 14332 34552
rect 15016 34604 15068 34610
rect 15016 34546 15068 34552
rect 13360 34536 13412 34542
rect 13360 34478 13412 34484
rect 13820 34536 13872 34542
rect 13820 34478 13872 34484
rect 14004 34536 14056 34542
rect 14004 34478 14056 34484
rect 14188 34536 14240 34542
rect 14188 34478 14240 34484
rect 14464 34536 14516 34542
rect 14464 34478 14516 34484
rect 13360 34060 13412 34066
rect 13360 34002 13412 34008
rect 13268 33992 13320 33998
rect 13268 33934 13320 33940
rect 13280 33658 13308 33934
rect 13268 33652 13320 33658
rect 13268 33594 13320 33600
rect 13372 33454 13400 34002
rect 14016 33454 14044 34478
rect 14200 33454 14228 34478
rect 14476 34202 14504 34478
rect 14464 34196 14516 34202
rect 14464 34138 14516 34144
rect 12992 33448 13044 33454
rect 12992 33390 13044 33396
rect 13360 33448 13412 33454
rect 13360 33390 13412 33396
rect 14004 33448 14056 33454
rect 14004 33390 14056 33396
rect 14188 33448 14240 33454
rect 14188 33390 14240 33396
rect 13004 33114 13032 33390
rect 12992 33108 13044 33114
rect 12992 33050 13044 33056
rect 14016 33046 14044 33390
rect 14004 33040 14056 33046
rect 14004 32982 14056 32988
rect 14280 32496 14332 32502
rect 14280 32438 14332 32444
rect 14292 31890 14320 32438
rect 14924 32360 14976 32366
rect 14924 32302 14976 32308
rect 14280 31884 14332 31890
rect 14280 31826 14332 31832
rect 14372 31884 14424 31890
rect 14372 31826 14424 31832
rect 13820 31816 13872 31822
rect 13820 31758 13872 31764
rect 13832 31346 13860 31758
rect 13820 31340 13872 31346
rect 13820 31282 13872 31288
rect 13084 31272 13136 31278
rect 13084 31214 13136 31220
rect 12900 31136 12952 31142
rect 12900 31078 12952 31084
rect 12912 30190 12940 31078
rect 12992 30252 13044 30258
rect 12992 30194 13044 30200
rect 12900 30184 12952 30190
rect 12900 30126 12952 30132
rect 12912 28558 12940 30126
rect 13004 29714 13032 30194
rect 12992 29708 13044 29714
rect 12992 29650 13044 29656
rect 12900 28552 12952 28558
rect 12900 28494 12952 28500
rect 13096 27538 13124 31214
rect 13728 30796 13780 30802
rect 13728 30738 13780 30744
rect 13740 29850 13768 30738
rect 13820 30660 13872 30666
rect 13820 30602 13872 30608
rect 13832 30394 13860 30602
rect 13820 30388 13872 30394
rect 13820 30330 13872 30336
rect 14384 30190 14412 31826
rect 14936 31822 14964 32302
rect 14924 31816 14976 31822
rect 14924 31758 14976 31764
rect 14648 31136 14700 31142
rect 14648 31078 14700 31084
rect 14660 30938 14688 31078
rect 14648 30932 14700 30938
rect 14648 30874 14700 30880
rect 14464 30728 14516 30734
rect 14464 30670 14516 30676
rect 14280 30184 14332 30190
rect 14280 30126 14332 30132
rect 14372 30184 14424 30190
rect 14372 30126 14424 30132
rect 13728 29844 13780 29850
rect 13728 29786 13780 29792
rect 14292 29238 14320 30126
rect 14476 29714 14504 30670
rect 14660 30258 14688 30874
rect 14740 30592 14792 30598
rect 14740 30534 14792 30540
rect 14648 30252 14700 30258
rect 14648 30194 14700 30200
rect 14556 30184 14608 30190
rect 14752 30138 14780 30534
rect 14556 30126 14608 30132
rect 14568 29850 14596 30126
rect 14660 30110 14780 30138
rect 14556 29844 14608 29850
rect 14556 29786 14608 29792
rect 14464 29708 14516 29714
rect 14464 29650 14516 29656
rect 14280 29232 14332 29238
rect 14280 29174 14332 29180
rect 13360 29028 13412 29034
rect 13360 28970 13412 28976
rect 13372 28762 13400 28970
rect 13268 28756 13320 28762
rect 13268 28698 13320 28704
rect 13360 28756 13412 28762
rect 13360 28698 13412 28704
rect 13280 28642 13308 28698
rect 13280 28626 13492 28642
rect 13280 28620 13504 28626
rect 13280 28614 13452 28620
rect 13452 28562 13504 28568
rect 13820 28008 13872 28014
rect 13820 27950 13872 27956
rect 13832 27538 13860 27950
rect 14292 27674 14320 29174
rect 14568 29170 14596 29786
rect 14556 29164 14608 29170
rect 14556 29106 14608 29112
rect 14372 29096 14424 29102
rect 14372 29038 14424 29044
rect 14384 28218 14412 29038
rect 14372 28212 14424 28218
rect 14372 28154 14424 28160
rect 14384 27946 14412 28154
rect 14372 27940 14424 27946
rect 14372 27882 14424 27888
rect 14464 27872 14516 27878
rect 14464 27814 14516 27820
rect 14280 27668 14332 27674
rect 14280 27610 14332 27616
rect 14476 27538 14504 27814
rect 13084 27532 13136 27538
rect 13084 27474 13136 27480
rect 13820 27532 13872 27538
rect 13820 27474 13872 27480
rect 14004 27532 14056 27538
rect 14004 27474 14056 27480
rect 14464 27532 14516 27538
rect 14464 27474 14516 27480
rect 14556 27532 14608 27538
rect 14556 27474 14608 27480
rect 13096 26926 13124 27474
rect 13820 27056 13872 27062
rect 13820 26998 13872 27004
rect 12992 26920 13044 26926
rect 12992 26862 13044 26868
rect 13084 26920 13136 26926
rect 13084 26862 13136 26868
rect 13004 26450 13032 26862
rect 13832 26450 13860 26998
rect 12992 26444 13044 26450
rect 12992 26386 13044 26392
rect 13820 26444 13872 26450
rect 13820 26386 13872 26392
rect 13084 26376 13136 26382
rect 13084 26318 13136 26324
rect 13096 26246 13124 26318
rect 13084 26240 13136 26246
rect 13084 26182 13136 26188
rect 12900 22976 12952 22982
rect 12900 22918 12952 22924
rect 12912 22137 12940 22918
rect 13096 22438 13124 26182
rect 13544 25900 13596 25906
rect 13544 25842 13596 25848
rect 13452 25764 13504 25770
rect 13452 25706 13504 25712
rect 13176 24268 13228 24274
rect 13176 24210 13228 24216
rect 13268 24268 13320 24274
rect 13268 24210 13320 24216
rect 13188 22642 13216 24210
rect 13280 23254 13308 24210
rect 13268 23248 13320 23254
rect 13268 23190 13320 23196
rect 13176 22636 13228 22642
rect 13176 22578 13228 22584
rect 13084 22432 13136 22438
rect 13084 22374 13136 22380
rect 12898 22128 12954 22137
rect 12898 22063 12954 22072
rect 13464 20058 13492 25706
rect 13556 25158 13584 25842
rect 13820 25832 13872 25838
rect 13820 25774 13872 25780
rect 13544 25152 13596 25158
rect 13544 25094 13596 25100
rect 13556 24818 13584 25094
rect 13544 24812 13596 24818
rect 13544 24754 13596 24760
rect 13832 24138 13860 25774
rect 13820 24132 13872 24138
rect 13820 24074 13872 24080
rect 13912 23180 13964 23186
rect 13912 23122 13964 23128
rect 13924 21894 13952 23122
rect 14016 23050 14044 27474
rect 14372 26784 14424 26790
rect 14372 26726 14424 26732
rect 14280 26376 14332 26382
rect 14280 26318 14332 26324
rect 14292 24750 14320 26318
rect 14384 25838 14412 26726
rect 14372 25832 14424 25838
rect 14372 25774 14424 25780
rect 14280 24744 14332 24750
rect 14280 24686 14332 24692
rect 14568 23798 14596 27474
rect 14660 25906 14688 30110
rect 14924 29096 14976 29102
rect 14924 29038 14976 29044
rect 14936 27946 14964 29038
rect 14924 27940 14976 27946
rect 14924 27882 14976 27888
rect 14740 27464 14792 27470
rect 14740 27406 14792 27412
rect 14752 27130 14780 27406
rect 14740 27124 14792 27130
rect 14740 27066 14792 27072
rect 14648 25900 14700 25906
rect 14648 25842 14700 25848
rect 15028 25242 15056 34546
rect 15292 33992 15344 33998
rect 15292 33934 15344 33940
rect 15304 33114 15332 33934
rect 15292 33108 15344 33114
rect 15292 33050 15344 33056
rect 15304 32910 15332 33050
rect 15292 32904 15344 32910
rect 15292 32846 15344 32852
rect 15304 31278 15332 32846
rect 15292 31272 15344 31278
rect 15292 31214 15344 31220
rect 15200 31204 15252 31210
rect 15200 31146 15252 31152
rect 15212 30802 15240 31146
rect 15200 30796 15252 30802
rect 15200 30738 15252 30744
rect 15212 30190 15240 30738
rect 15200 30184 15252 30190
rect 15200 30126 15252 30132
rect 15488 28744 15516 36178
rect 15580 35222 15608 36178
rect 15568 35216 15620 35222
rect 15568 35158 15620 35164
rect 15568 35080 15620 35086
rect 15568 35022 15620 35028
rect 15580 32978 15608 35022
rect 15568 32972 15620 32978
rect 15568 32914 15620 32920
rect 15568 32360 15620 32366
rect 15568 32302 15620 32308
rect 15580 31890 15608 32302
rect 15568 31884 15620 31890
rect 15568 31826 15620 31832
rect 15672 30274 15700 39200
rect 15752 37256 15804 37262
rect 15752 37198 15804 37204
rect 15764 36854 15792 37198
rect 16856 37120 16908 37126
rect 16856 37062 16908 37068
rect 15752 36848 15804 36854
rect 15752 36790 15804 36796
rect 16868 36786 16896 37062
rect 16856 36780 16908 36786
rect 16856 36722 16908 36728
rect 15752 36712 15804 36718
rect 15752 36654 15804 36660
rect 15764 36242 15792 36654
rect 17040 36576 17092 36582
rect 17040 36518 17092 36524
rect 15752 36236 15804 36242
rect 15804 36196 15884 36224
rect 15752 36178 15804 36184
rect 15752 36032 15804 36038
rect 15752 35974 15804 35980
rect 15764 35698 15792 35974
rect 15752 35692 15804 35698
rect 15752 35634 15804 35640
rect 15856 35630 15884 36196
rect 17052 36174 17080 36518
rect 17040 36168 17092 36174
rect 17040 36110 17092 36116
rect 15844 35624 15896 35630
rect 15844 35566 15896 35572
rect 16488 35624 16540 35630
rect 16488 35566 16540 35572
rect 16120 35556 16172 35562
rect 16120 35498 16172 35504
rect 15844 35080 15896 35086
rect 15844 35022 15896 35028
rect 15856 32026 15884 35022
rect 16132 34610 16160 35498
rect 16500 35290 16528 35566
rect 16488 35284 16540 35290
rect 16488 35226 16540 35232
rect 16488 35080 16540 35086
rect 16488 35022 16540 35028
rect 16120 34604 16172 34610
rect 16120 34546 16172 34552
rect 16500 34082 16528 35022
rect 16856 34672 16908 34678
rect 16856 34614 16908 34620
rect 16316 34054 16528 34082
rect 16868 34066 16896 34614
rect 16316 32774 16344 34054
rect 16396 33992 16448 33998
rect 16396 33934 16448 33940
rect 16408 33658 16436 33934
rect 16396 33652 16448 33658
rect 16500 33640 16528 34054
rect 16856 34060 16908 34066
rect 16856 34002 16908 34008
rect 16580 33652 16632 33658
rect 16500 33612 16580 33640
rect 16396 33594 16448 33600
rect 16580 33594 16632 33600
rect 16396 33516 16448 33522
rect 16448 33476 16620 33504
rect 16396 33458 16448 33464
rect 16304 32768 16356 32774
rect 16304 32710 16356 32716
rect 16316 32502 16344 32710
rect 16304 32496 16356 32502
rect 16224 32456 16304 32484
rect 15844 32020 15896 32026
rect 15844 31962 15896 31968
rect 16224 31822 16252 32456
rect 16304 32438 16356 32444
rect 16592 32434 16620 33476
rect 16948 32904 17000 32910
rect 16948 32846 17000 32852
rect 16856 32768 16908 32774
rect 16856 32710 16908 32716
rect 16580 32428 16632 32434
rect 16580 32370 16632 32376
rect 16304 32360 16356 32366
rect 16304 32302 16356 32308
rect 16672 32360 16724 32366
rect 16672 32302 16724 32308
rect 16212 31816 16264 31822
rect 16212 31758 16264 31764
rect 16316 31278 16344 32302
rect 16580 31884 16632 31890
rect 16580 31826 16632 31832
rect 16304 31272 16356 31278
rect 16304 31214 16356 31220
rect 16316 30938 16344 31214
rect 16304 30932 16356 30938
rect 16304 30874 16356 30880
rect 16396 30796 16448 30802
rect 16396 30738 16448 30744
rect 15672 30246 16344 30274
rect 15660 30048 15712 30054
rect 15660 29990 15712 29996
rect 15752 30048 15804 30054
rect 15752 29990 15804 29996
rect 16028 30048 16080 30054
rect 16028 29990 16080 29996
rect 15672 29850 15700 29990
rect 15660 29844 15712 29850
rect 15660 29786 15712 29792
rect 15764 29714 15792 29990
rect 16040 29714 16068 29990
rect 15752 29708 15804 29714
rect 15752 29650 15804 29656
rect 16028 29708 16080 29714
rect 16028 29650 16080 29656
rect 15844 29232 15896 29238
rect 15844 29174 15896 29180
rect 15304 28716 15516 28744
rect 15304 28150 15332 28716
rect 15384 28620 15436 28626
rect 15384 28562 15436 28568
rect 15752 28620 15804 28626
rect 15752 28562 15804 28568
rect 15292 28144 15344 28150
rect 15292 28086 15344 28092
rect 15304 27878 15332 28086
rect 15292 27872 15344 27878
rect 15292 27814 15344 27820
rect 15108 27668 15160 27674
rect 15108 27610 15160 27616
rect 15120 26926 15148 27610
rect 15108 26920 15160 26926
rect 15108 26862 15160 26868
rect 15108 26376 15160 26382
rect 15108 26318 15160 26324
rect 14844 25214 15056 25242
rect 14648 24744 14700 24750
rect 14648 24686 14700 24692
rect 14660 24274 14688 24686
rect 14648 24268 14700 24274
rect 14648 24210 14700 24216
rect 14556 23792 14608 23798
rect 14556 23734 14608 23740
rect 14660 23730 14688 24210
rect 14648 23724 14700 23730
rect 14648 23666 14700 23672
rect 14372 23316 14424 23322
rect 14372 23258 14424 23264
rect 14004 23044 14056 23050
rect 14004 22986 14056 22992
rect 14384 22574 14412 23258
rect 14464 23112 14516 23118
rect 14464 23054 14516 23060
rect 14372 22568 14424 22574
rect 14372 22510 14424 22516
rect 13912 21888 13964 21894
rect 13912 21830 13964 21836
rect 14370 21584 14426 21593
rect 14370 21519 14426 21528
rect 13820 21480 13872 21486
rect 13820 21422 13872 21428
rect 14004 21480 14056 21486
rect 14004 21422 14056 21428
rect 13728 21344 13780 21350
rect 13728 21286 13780 21292
rect 13544 20868 13596 20874
rect 13544 20810 13596 20816
rect 13452 20052 13504 20058
rect 13452 19994 13504 20000
rect 13556 19922 13584 20810
rect 13544 19916 13596 19922
rect 13544 19858 13596 19864
rect 13740 19378 13768 21286
rect 13832 20942 13860 21422
rect 13820 20936 13872 20942
rect 13820 20878 13872 20884
rect 14016 20602 14044 21422
rect 14096 21412 14148 21418
rect 14096 21354 14148 21360
rect 14004 20596 14056 20602
rect 14004 20538 14056 20544
rect 14108 19922 14136 21354
rect 14384 21350 14412 21519
rect 14372 21344 14424 21350
rect 14372 21286 14424 21292
rect 14188 20936 14240 20942
rect 14188 20878 14240 20884
rect 14004 19916 14056 19922
rect 14004 19858 14056 19864
rect 14096 19916 14148 19922
rect 14096 19858 14148 19864
rect 13820 19712 13872 19718
rect 13820 19654 13872 19660
rect 13728 19372 13780 19378
rect 13728 19314 13780 19320
rect 13544 19304 13596 19310
rect 13544 19246 13596 19252
rect 13556 18902 13584 19246
rect 13740 18902 13768 19314
rect 13544 18896 13596 18902
rect 13544 18838 13596 18844
rect 13728 18896 13780 18902
rect 13728 18838 13780 18844
rect 13636 17128 13688 17134
rect 13740 17116 13768 18838
rect 13832 18222 13860 19654
rect 13912 18692 13964 18698
rect 13912 18634 13964 18640
rect 13924 18222 13952 18634
rect 13820 18216 13872 18222
rect 13820 18158 13872 18164
rect 13912 18216 13964 18222
rect 13912 18158 13964 18164
rect 13820 17536 13872 17542
rect 13820 17478 13872 17484
rect 13832 17134 13860 17478
rect 13688 17088 13768 17116
rect 13820 17128 13872 17134
rect 13636 17070 13688 17076
rect 13820 17070 13872 17076
rect 12808 16788 12860 16794
rect 12808 16730 12860 16736
rect 12716 16652 12768 16658
rect 12768 16612 12848 16640
rect 12716 16594 12768 16600
rect 12624 16448 12676 16454
rect 12624 16390 12676 16396
rect 12820 16046 12848 16612
rect 14016 16130 14044 19858
rect 14200 19310 14228 20878
rect 14188 19304 14240 19310
rect 14188 19246 14240 19252
rect 14200 17134 14228 19246
rect 14280 19168 14332 19174
rect 14280 19110 14332 19116
rect 14292 18834 14320 19110
rect 14280 18828 14332 18834
rect 14280 18770 14332 18776
rect 14384 18714 14412 21286
rect 14476 21010 14504 23054
rect 14660 21146 14688 23666
rect 14648 21140 14700 21146
rect 14648 21082 14700 21088
rect 14464 21004 14516 21010
rect 14464 20946 14516 20952
rect 14844 20602 14872 25214
rect 14924 25152 14976 25158
rect 14924 25094 14976 25100
rect 14936 24750 14964 25094
rect 14924 24744 14976 24750
rect 14924 24686 14976 24692
rect 14924 24608 14976 24614
rect 14924 24550 14976 24556
rect 14936 24342 14964 24550
rect 14924 24336 14976 24342
rect 14924 24278 14976 24284
rect 14936 24070 14964 24278
rect 15120 24274 15148 26318
rect 15396 25974 15424 28562
rect 15568 26852 15620 26858
rect 15568 26794 15620 26800
rect 15384 25968 15436 25974
rect 15384 25910 15436 25916
rect 15200 25356 15252 25362
rect 15200 25298 15252 25304
rect 15108 24268 15160 24274
rect 15108 24210 15160 24216
rect 14924 24064 14976 24070
rect 14924 24006 14976 24012
rect 14936 23662 14964 24006
rect 14924 23656 14976 23662
rect 14924 23598 14976 23604
rect 14936 23118 14964 23598
rect 15120 23526 15148 24210
rect 15108 23520 15160 23526
rect 15108 23462 15160 23468
rect 15016 23316 15068 23322
rect 15016 23258 15068 23264
rect 14924 23112 14976 23118
rect 14924 23054 14976 23060
rect 15028 21962 15056 23258
rect 15108 23044 15160 23050
rect 15108 22986 15160 22992
rect 15120 22506 15148 22986
rect 15108 22500 15160 22506
rect 15108 22442 15160 22448
rect 15120 22166 15148 22442
rect 15108 22160 15160 22166
rect 15108 22102 15160 22108
rect 15016 21956 15068 21962
rect 15016 21898 15068 21904
rect 15212 21010 15240 25298
rect 15580 25158 15608 26794
rect 15660 25832 15712 25838
rect 15660 25774 15712 25780
rect 15672 25498 15700 25774
rect 15660 25492 15712 25498
rect 15660 25434 15712 25440
rect 15568 25152 15620 25158
rect 15568 25094 15620 25100
rect 15580 24614 15608 25094
rect 15660 24744 15712 24750
rect 15660 24686 15712 24692
rect 15568 24608 15620 24614
rect 15568 24550 15620 24556
rect 15672 24070 15700 24686
rect 15660 24064 15712 24070
rect 15660 24006 15712 24012
rect 15476 23656 15528 23662
rect 15476 23598 15528 23604
rect 15384 23588 15436 23594
rect 15384 23530 15436 23536
rect 15292 23180 15344 23186
rect 15292 23122 15344 23128
rect 15200 21004 15252 21010
rect 15200 20946 15252 20952
rect 14556 20596 14608 20602
rect 14556 20538 14608 20544
rect 14832 20596 14884 20602
rect 14832 20538 14884 20544
rect 14568 20398 14596 20538
rect 14556 20392 14608 20398
rect 14556 20334 14608 20340
rect 14740 20392 14792 20398
rect 14740 20334 14792 20340
rect 14832 20392 14884 20398
rect 14832 20334 14884 20340
rect 14292 18686 14412 18714
rect 14188 17128 14240 17134
rect 14188 17070 14240 17076
rect 14016 16102 14136 16130
rect 12440 16040 12492 16046
rect 12440 15982 12492 15988
rect 12808 16040 12860 16046
rect 12808 15982 12860 15988
rect 13912 16040 13964 16046
rect 13912 15982 13964 15988
rect 12348 15904 12400 15910
rect 12348 15846 12400 15852
rect 12256 14884 12308 14890
rect 12256 14826 12308 14832
rect 11888 14476 11940 14482
rect 11888 14418 11940 14424
rect 11900 12850 11928 14418
rect 11888 12844 11940 12850
rect 11888 12786 11940 12792
rect 11980 12300 12032 12306
rect 11980 12242 12032 12248
rect 11796 10600 11848 10606
rect 11796 10542 11848 10548
rect 11796 10464 11848 10470
rect 11796 10406 11848 10412
rect 11702 10024 11758 10033
rect 11702 9959 11758 9968
rect 11704 9920 11756 9926
rect 11704 9862 11756 9868
rect 11716 9518 11744 9862
rect 11704 9512 11756 9518
rect 11704 9454 11756 9460
rect 11610 8120 11666 8129
rect 11808 8090 11836 10406
rect 11888 10124 11940 10130
rect 11888 10066 11940 10072
rect 11900 8498 11928 10066
rect 11888 8492 11940 8498
rect 11888 8434 11940 8440
rect 11610 8055 11666 8064
rect 11796 8084 11848 8090
rect 11796 8026 11848 8032
rect 11992 7970 12020 12242
rect 12268 12102 12296 14826
rect 12360 14346 12388 15846
rect 12452 15094 12480 15982
rect 13268 15496 13320 15502
rect 13268 15438 13320 15444
rect 12532 15360 12584 15366
rect 12532 15302 12584 15308
rect 12440 15088 12492 15094
rect 12440 15030 12492 15036
rect 12452 14958 12480 15030
rect 12440 14952 12492 14958
rect 12440 14894 12492 14900
rect 12348 14340 12400 14346
rect 12348 14282 12400 14288
rect 12256 12096 12308 12102
rect 12256 12038 12308 12044
rect 12544 10130 12572 15302
rect 13280 15094 13308 15438
rect 13268 15088 13320 15094
rect 13268 15030 13320 15036
rect 12808 14952 12860 14958
rect 12808 14894 12860 14900
rect 13268 14952 13320 14958
rect 13268 14894 13320 14900
rect 12716 13932 12768 13938
rect 12716 13874 12768 13880
rect 12728 11121 12756 13874
rect 12820 13870 12848 14894
rect 13280 14550 13308 14894
rect 13268 14544 13320 14550
rect 13174 14512 13230 14521
rect 13268 14486 13320 14492
rect 13174 14447 13230 14456
rect 13188 14414 13216 14447
rect 13176 14408 13228 14414
rect 13176 14350 13228 14356
rect 12808 13864 12860 13870
rect 12808 13806 12860 13812
rect 13188 12918 13216 14350
rect 13924 14346 13952 15982
rect 14004 15496 14056 15502
rect 14004 15438 14056 15444
rect 14016 14482 14044 15438
rect 14004 14476 14056 14482
rect 14004 14418 14056 14424
rect 13912 14340 13964 14346
rect 13912 14282 13964 14288
rect 13268 14000 13320 14006
rect 13268 13942 13320 13948
rect 13280 13394 13308 13942
rect 13452 13864 13504 13870
rect 13452 13806 13504 13812
rect 13268 13388 13320 13394
rect 13268 13330 13320 13336
rect 13360 13184 13412 13190
rect 13360 13126 13412 13132
rect 13176 12912 13228 12918
rect 13176 12854 13228 12860
rect 13372 12782 13400 13126
rect 13464 12850 13492 13806
rect 13912 13184 13964 13190
rect 13912 13126 13964 13132
rect 13452 12844 13504 12850
rect 13452 12786 13504 12792
rect 13360 12776 13412 12782
rect 13360 12718 13412 12724
rect 13924 12714 13952 13126
rect 13912 12708 13964 12714
rect 13912 12650 13964 12656
rect 13176 12300 13228 12306
rect 13176 12242 13228 12248
rect 13188 12102 13216 12242
rect 13360 12232 13412 12238
rect 13360 12174 13412 12180
rect 13176 12096 13228 12102
rect 13176 12038 13228 12044
rect 12992 11688 13044 11694
rect 12992 11630 13044 11636
rect 12900 11620 12952 11626
rect 12900 11562 12952 11568
rect 12808 11212 12860 11218
rect 12808 11154 12860 11160
rect 12714 11112 12770 11121
rect 12714 11047 12770 11056
rect 12624 10192 12676 10198
rect 12624 10134 12676 10140
rect 12532 10124 12584 10130
rect 12532 10066 12584 10072
rect 12072 10056 12124 10062
rect 12072 9998 12124 10004
rect 12256 10056 12308 10062
rect 12256 9998 12308 10004
rect 12084 9602 12112 9998
rect 12084 9574 12204 9602
rect 12268 9586 12296 9998
rect 12176 9518 12204 9574
rect 12256 9580 12308 9586
rect 12256 9522 12308 9528
rect 12164 9512 12216 9518
rect 12164 9454 12216 9460
rect 12072 9444 12124 9450
rect 12072 9386 12124 9392
rect 12084 9042 12112 9386
rect 12072 9036 12124 9042
rect 12072 8978 12124 8984
rect 12176 8974 12204 9454
rect 12164 8968 12216 8974
rect 12164 8910 12216 8916
rect 11532 7942 11836 7970
rect 11992 7942 12112 7970
rect 12176 7954 12204 8910
rect 12268 8820 12296 9522
rect 12636 9382 12664 10134
rect 12728 9654 12756 11047
rect 12820 10588 12848 11154
rect 12912 11082 12940 11562
rect 13004 11286 13032 11630
rect 12992 11280 13044 11286
rect 12992 11222 13044 11228
rect 13084 11212 13136 11218
rect 13084 11154 13136 11160
rect 12900 11076 12952 11082
rect 12900 11018 12952 11024
rect 12992 10600 13044 10606
rect 12820 10560 12992 10588
rect 12992 10542 13044 10548
rect 12716 9648 12768 9654
rect 12716 9590 12768 9596
rect 12624 9376 12676 9382
rect 12624 9318 12676 9324
rect 12636 8838 12664 9318
rect 12624 8832 12676 8838
rect 12268 8792 12388 8820
rect 12256 8560 12308 8566
rect 12256 8502 12308 8508
rect 12360 8514 12388 8792
rect 12624 8774 12676 8780
rect 11152 7812 11204 7818
rect 11152 7754 11204 7760
rect 11336 7812 11388 7818
rect 11336 7754 11388 7760
rect 11164 7721 11192 7754
rect 11428 7744 11480 7750
rect 11150 7712 11206 7721
rect 11428 7686 11480 7692
rect 11150 7647 11206 7656
rect 11440 7449 11468 7686
rect 11426 7440 11482 7449
rect 11060 7404 11112 7410
rect 11808 7410 11836 7942
rect 11980 7880 12032 7886
rect 11980 7822 12032 7828
rect 11426 7375 11482 7384
rect 11796 7404 11848 7410
rect 11060 7346 11112 7352
rect 10968 6928 11020 6934
rect 10968 6870 11020 6876
rect 11072 5778 11100 7346
rect 11440 7342 11468 7375
rect 11796 7346 11848 7352
rect 11428 7336 11480 7342
rect 11428 7278 11480 7284
rect 11704 7336 11756 7342
rect 11704 7278 11756 7284
rect 11716 7002 11744 7278
rect 11992 7206 12020 7822
rect 11980 7200 12032 7206
rect 11980 7142 12032 7148
rect 11704 6996 11756 7002
rect 11704 6938 11756 6944
rect 11992 6254 12020 7142
rect 11244 6248 11296 6254
rect 11244 6190 11296 6196
rect 11980 6248 12032 6254
rect 11980 6190 12032 6196
rect 11256 5914 11284 6190
rect 11244 5908 11296 5914
rect 11244 5850 11296 5856
rect 11060 5772 11112 5778
rect 11060 5714 11112 5720
rect 11980 5772 12032 5778
rect 11980 5714 12032 5720
rect 10968 5704 11020 5710
rect 10968 5646 11020 5652
rect 10876 5228 10928 5234
rect 10876 5170 10928 5176
rect 10888 4690 10916 5170
rect 10980 5166 11008 5646
rect 11520 5568 11572 5574
rect 11520 5510 11572 5516
rect 11532 5166 11560 5510
rect 10968 5160 11020 5166
rect 10966 5128 10968 5137
rect 11520 5160 11572 5166
rect 11020 5128 11022 5137
rect 11520 5102 11572 5108
rect 10966 5063 11022 5072
rect 11532 4690 11560 5102
rect 11992 5030 12020 5714
rect 11980 5024 12032 5030
rect 11980 4966 12032 4972
rect 12084 4826 12112 7942
rect 12164 7948 12216 7954
rect 12164 7890 12216 7896
rect 12268 7750 12296 8502
rect 12360 8486 12940 8514
rect 12912 8430 12940 8486
rect 12624 8424 12676 8430
rect 12624 8366 12676 8372
rect 12900 8424 12952 8430
rect 12900 8366 12952 8372
rect 12256 7744 12308 7750
rect 12256 7686 12308 7692
rect 12164 7200 12216 7206
rect 12164 7142 12216 7148
rect 12176 6934 12204 7142
rect 12164 6928 12216 6934
rect 12164 6870 12216 6876
rect 12440 6860 12492 6866
rect 12268 6820 12440 6848
rect 12164 6792 12216 6798
rect 12268 6780 12296 6820
rect 12440 6802 12492 6808
rect 12216 6752 12296 6780
rect 12532 6792 12584 6798
rect 12164 6734 12216 6740
rect 12532 6734 12584 6740
rect 12544 6458 12572 6734
rect 12532 6452 12584 6458
rect 12532 6394 12584 6400
rect 12440 6248 12492 6254
rect 12440 6190 12492 6196
rect 12452 5302 12480 6190
rect 12532 5840 12584 5846
rect 12532 5782 12584 5788
rect 12440 5296 12492 5302
rect 12440 5238 12492 5244
rect 12072 4820 12124 4826
rect 12072 4762 12124 4768
rect 10692 4684 10744 4690
rect 10692 4626 10744 4632
rect 10876 4684 10928 4690
rect 10876 4626 10928 4632
rect 11244 4684 11296 4690
rect 11244 4626 11296 4632
rect 11520 4684 11572 4690
rect 11520 4626 11572 4632
rect 10704 4214 10732 4626
rect 10692 4208 10744 4214
rect 10692 4150 10744 4156
rect 10888 4146 10916 4626
rect 11256 4282 11284 4626
rect 11244 4276 11296 4282
rect 11244 4218 11296 4224
rect 11532 4146 11560 4626
rect 10876 4140 10928 4146
rect 10876 4082 10928 4088
rect 11520 4140 11572 4146
rect 11520 4082 11572 4088
rect 10508 4072 10560 4078
rect 10508 4014 10560 4020
rect 11428 4072 11480 4078
rect 11428 4014 11480 4020
rect 11440 3194 11468 4014
rect 12256 3596 12308 3602
rect 12256 3538 12308 3544
rect 11428 3188 11480 3194
rect 11428 3130 11480 3136
rect 12268 3126 12296 3538
rect 12440 3528 12492 3534
rect 12440 3470 12492 3476
rect 12348 3460 12400 3466
rect 12348 3402 12400 3408
rect 12256 3120 12308 3126
rect 12256 3062 12308 3068
rect 12360 3058 12388 3402
rect 12348 3052 12400 3058
rect 12348 2994 12400 3000
rect 10140 2984 10192 2990
rect 10140 2926 10192 2932
rect 10600 2848 10652 2854
rect 10652 2796 10732 2802
rect 10600 2790 10732 2796
rect 10612 2774 10732 2790
rect 9864 2644 9916 2650
rect 9864 2586 9916 2592
rect 9680 2508 9732 2514
rect 9680 2450 9732 2456
rect 9312 2440 9364 2446
rect 9312 2382 9364 2388
rect 7932 2100 7984 2106
rect 7932 2042 7984 2048
rect 6920 2032 6972 2038
rect 6920 1974 6972 1980
rect 8668 2032 8720 2038
rect 8668 1974 8720 1980
rect 8680 800 8708 1974
rect 10704 800 10732 2774
rect 12452 2514 12480 3470
rect 12544 2990 12572 5782
rect 12636 5778 12664 8366
rect 13004 7954 13032 10542
rect 12992 7948 13044 7954
rect 12992 7890 13044 7896
rect 13004 7449 13032 7890
rect 12990 7440 13046 7449
rect 12990 7375 13046 7384
rect 12716 7268 12768 7274
rect 12716 7210 12768 7216
rect 12728 6254 12756 7210
rect 13096 6730 13124 11154
rect 13188 10742 13216 12038
rect 13372 11694 13400 12174
rect 13360 11688 13412 11694
rect 13360 11630 13412 11636
rect 13820 11008 13872 11014
rect 13820 10950 13872 10956
rect 13176 10736 13228 10742
rect 13176 10678 13228 10684
rect 13268 10600 13320 10606
rect 13268 10542 13320 10548
rect 13280 9654 13308 10542
rect 13832 10130 13860 10950
rect 13820 10124 13872 10130
rect 13820 10066 13872 10072
rect 13268 9648 13320 9654
rect 13268 9590 13320 9596
rect 13924 9042 13952 12650
rect 14108 10674 14136 16102
rect 14188 15564 14240 15570
rect 14188 15506 14240 15512
rect 14200 14822 14228 15506
rect 14292 14890 14320 18686
rect 14568 18222 14596 20334
rect 14752 19718 14780 20334
rect 14740 19712 14792 19718
rect 14740 19654 14792 19660
rect 14844 19514 14872 20334
rect 15304 19802 15332 23122
rect 15396 21894 15424 23530
rect 15384 21888 15436 21894
rect 15384 21830 15436 21836
rect 15384 21480 15436 21486
rect 15384 21422 15436 21428
rect 15396 21146 15424 21422
rect 15384 21140 15436 21146
rect 15384 21082 15436 21088
rect 15488 20398 15516 23598
rect 15568 22568 15620 22574
rect 15568 22510 15620 22516
rect 15580 21622 15608 22510
rect 15568 21616 15620 21622
rect 15568 21558 15620 21564
rect 15568 21480 15620 21486
rect 15568 21422 15620 21428
rect 15476 20392 15528 20398
rect 15476 20334 15528 20340
rect 15476 19916 15528 19922
rect 15476 19858 15528 19864
rect 15304 19774 15424 19802
rect 14832 19508 14884 19514
rect 14832 19450 14884 19456
rect 15200 19304 15252 19310
rect 15200 19246 15252 19252
rect 15292 19304 15344 19310
rect 15292 19246 15344 19252
rect 14556 18216 14608 18222
rect 14556 18158 14608 18164
rect 14648 17672 14700 17678
rect 14648 17614 14700 17620
rect 14660 17202 14688 17614
rect 14648 17196 14700 17202
rect 14648 17138 14700 17144
rect 15108 17196 15160 17202
rect 15108 17138 15160 17144
rect 14372 16652 14424 16658
rect 14372 16594 14424 16600
rect 14280 14884 14332 14890
rect 14280 14826 14332 14832
rect 14188 14816 14240 14822
rect 14188 14758 14240 14764
rect 14200 14550 14228 14758
rect 14188 14544 14240 14550
rect 14188 14486 14240 14492
rect 14280 14340 14332 14346
rect 14280 14282 14332 14288
rect 14292 13938 14320 14282
rect 14280 13932 14332 13938
rect 14280 13874 14332 13880
rect 14188 13252 14240 13258
rect 14188 13194 14240 13200
rect 14096 10668 14148 10674
rect 14096 10610 14148 10616
rect 14004 10532 14056 10538
rect 14004 10474 14056 10480
rect 14016 10130 14044 10474
rect 14004 10124 14056 10130
rect 14004 10066 14056 10072
rect 14096 10056 14148 10062
rect 14096 9998 14148 10004
rect 14108 9722 14136 9998
rect 14096 9716 14148 9722
rect 14096 9658 14148 9664
rect 14096 9580 14148 9586
rect 14096 9522 14148 9528
rect 14004 9376 14056 9382
rect 14004 9318 14056 9324
rect 14016 9042 14044 9318
rect 13912 9036 13964 9042
rect 13912 8978 13964 8984
rect 14004 9036 14056 9042
rect 14004 8978 14056 8984
rect 13452 8968 13504 8974
rect 13452 8910 13504 8916
rect 13820 8968 13872 8974
rect 13820 8910 13872 8916
rect 13268 8832 13320 8838
rect 13268 8774 13320 8780
rect 13280 8430 13308 8774
rect 13464 8634 13492 8910
rect 13452 8628 13504 8634
rect 13452 8570 13504 8576
rect 13268 8424 13320 8430
rect 13268 8366 13320 8372
rect 13360 8424 13412 8430
rect 13360 8366 13412 8372
rect 13372 7886 13400 8366
rect 13832 8090 13860 8910
rect 13912 8424 13964 8430
rect 13912 8366 13964 8372
rect 13820 8084 13872 8090
rect 13820 8026 13872 8032
rect 13636 7948 13688 7954
rect 13636 7890 13688 7896
rect 13360 7880 13412 7886
rect 13360 7822 13412 7828
rect 13648 7478 13676 7890
rect 13636 7472 13688 7478
rect 13636 7414 13688 7420
rect 13924 7342 13952 8366
rect 14108 7342 14136 9522
rect 14200 7546 14228 13194
rect 14384 12306 14412 16594
rect 15120 16046 15148 17138
rect 15108 16040 15160 16046
rect 15108 15982 15160 15988
rect 14462 15192 14518 15201
rect 14462 15127 14464 15136
rect 14516 15127 14518 15136
rect 14464 15098 14516 15104
rect 15120 14890 15148 15982
rect 15108 14884 15160 14890
rect 15028 14844 15108 14872
rect 14464 14816 14516 14822
rect 14464 14758 14516 14764
rect 14476 13258 14504 14758
rect 15028 13870 15056 14844
rect 15108 14826 15160 14832
rect 15108 13932 15160 13938
rect 15108 13874 15160 13880
rect 15016 13864 15068 13870
rect 15016 13806 15068 13812
rect 14556 13388 14608 13394
rect 14556 13330 14608 13336
rect 14924 13388 14976 13394
rect 14924 13330 14976 13336
rect 14568 13258 14596 13330
rect 14464 13252 14516 13258
rect 14464 13194 14516 13200
rect 14556 13252 14608 13258
rect 14556 13194 14608 13200
rect 14648 12776 14700 12782
rect 14568 12724 14648 12730
rect 14568 12718 14700 12724
rect 14568 12702 14688 12718
rect 14372 12300 14424 12306
rect 14292 12260 14372 12288
rect 14292 8430 14320 12260
rect 14372 12242 14424 12248
rect 14464 11756 14516 11762
rect 14464 11698 14516 11704
rect 14372 11552 14424 11558
rect 14372 11494 14424 11500
rect 14384 11218 14412 11494
rect 14476 11218 14504 11698
rect 14372 11212 14424 11218
rect 14372 11154 14424 11160
rect 14464 11212 14516 11218
rect 14464 11154 14516 11160
rect 14464 9512 14516 9518
rect 14464 9454 14516 9460
rect 14476 9110 14504 9454
rect 14464 9104 14516 9110
rect 14464 9046 14516 9052
rect 14280 8424 14332 8430
rect 14280 8366 14332 8372
rect 14280 7948 14332 7954
rect 14280 7890 14332 7896
rect 14188 7540 14240 7546
rect 14188 7482 14240 7488
rect 13912 7336 13964 7342
rect 13912 7278 13964 7284
rect 14096 7336 14148 7342
rect 14096 7278 14148 7284
rect 13924 6866 13952 7278
rect 14108 6866 14136 7278
rect 13912 6860 13964 6866
rect 13912 6802 13964 6808
rect 14096 6860 14148 6866
rect 14096 6802 14148 6808
rect 13084 6724 13136 6730
rect 13084 6666 13136 6672
rect 13268 6384 13320 6390
rect 13268 6326 13320 6332
rect 12716 6248 12768 6254
rect 12716 6190 12768 6196
rect 12808 6180 12860 6186
rect 12808 6122 12860 6128
rect 12624 5772 12676 5778
rect 12624 5714 12676 5720
rect 12636 3942 12664 5714
rect 12716 5704 12768 5710
rect 12716 5646 12768 5652
rect 12728 4690 12756 5646
rect 12716 4684 12768 4690
rect 12716 4626 12768 4632
rect 12624 3936 12676 3942
rect 12624 3878 12676 3884
rect 12624 3732 12676 3738
rect 12624 3674 12676 3680
rect 12532 2984 12584 2990
rect 12532 2926 12584 2932
rect 12440 2508 12492 2514
rect 12440 2450 12492 2456
rect 12636 2446 12664 3674
rect 12820 3602 12848 6122
rect 13280 5914 13308 6326
rect 13912 6248 13964 6254
rect 13912 6190 13964 6196
rect 13268 5908 13320 5914
rect 13268 5850 13320 5856
rect 13728 5772 13780 5778
rect 13728 5714 13780 5720
rect 12992 5704 13044 5710
rect 12992 5646 13044 5652
rect 13004 5234 13032 5646
rect 13740 5574 13768 5714
rect 13728 5568 13780 5574
rect 13728 5510 13780 5516
rect 13924 5302 13952 6190
rect 13912 5296 13964 5302
rect 13912 5238 13964 5244
rect 12992 5228 13044 5234
rect 12992 5170 13044 5176
rect 13728 5228 13780 5234
rect 13728 5170 13780 5176
rect 13740 5137 13768 5170
rect 14292 5166 14320 7890
rect 14568 7410 14596 12702
rect 14740 12164 14792 12170
rect 14740 12106 14792 12112
rect 14648 12096 14700 12102
rect 14648 12038 14700 12044
rect 14660 11694 14688 12038
rect 14752 11898 14780 12106
rect 14740 11892 14792 11898
rect 14740 11834 14792 11840
rect 14648 11688 14700 11694
rect 14648 11630 14700 11636
rect 14738 11656 14794 11665
rect 14738 11591 14794 11600
rect 14648 11552 14700 11558
rect 14648 11494 14700 11500
rect 14660 11354 14688 11494
rect 14648 11348 14700 11354
rect 14648 11290 14700 11296
rect 14752 11286 14780 11591
rect 14740 11280 14792 11286
rect 14740 11222 14792 11228
rect 14936 7886 14964 13330
rect 15120 12782 15148 13874
rect 15108 12776 15160 12782
rect 15108 12718 15160 12724
rect 15016 10600 15068 10606
rect 15016 10542 15068 10548
rect 15028 10441 15056 10542
rect 15014 10432 15070 10441
rect 15014 10367 15070 10376
rect 15212 8566 15240 19246
rect 15304 18902 15332 19246
rect 15292 18896 15344 18902
rect 15292 18838 15344 18844
rect 15396 18850 15424 19774
rect 15488 18970 15516 19858
rect 15476 18964 15528 18970
rect 15476 18906 15528 18912
rect 15396 18822 15516 18850
rect 15292 17740 15344 17746
rect 15292 17682 15344 17688
rect 15304 16522 15332 17682
rect 15488 17610 15516 18822
rect 15580 18698 15608 21422
rect 15660 20936 15712 20942
rect 15660 20878 15712 20884
rect 15568 18692 15620 18698
rect 15568 18634 15620 18640
rect 15672 17898 15700 20878
rect 15764 20534 15792 28562
rect 15856 27538 15884 29174
rect 16040 29170 16068 29650
rect 16028 29164 16080 29170
rect 16028 29106 16080 29112
rect 15936 28008 15988 28014
rect 15936 27950 15988 27956
rect 15844 27532 15896 27538
rect 15844 27474 15896 27480
rect 15948 27334 15976 27950
rect 15936 27328 15988 27334
rect 15936 27270 15988 27276
rect 15844 26988 15896 26994
rect 15844 26930 15896 26936
rect 15856 26450 15884 26930
rect 15844 26444 15896 26450
rect 15844 26386 15896 26392
rect 15856 25702 15884 26386
rect 15844 25696 15896 25702
rect 15844 25638 15896 25644
rect 15856 25498 15884 25638
rect 15844 25492 15896 25498
rect 15844 25434 15896 25440
rect 16040 25430 16068 29106
rect 16212 28620 16264 28626
rect 16212 28562 16264 28568
rect 16120 28552 16172 28558
rect 16120 28494 16172 28500
rect 16132 28082 16160 28494
rect 16224 28150 16252 28562
rect 16212 28144 16264 28150
rect 16212 28086 16264 28092
rect 16120 28076 16172 28082
rect 16120 28018 16172 28024
rect 16120 26444 16172 26450
rect 16120 26386 16172 26392
rect 16132 25838 16160 26386
rect 16120 25832 16172 25838
rect 16120 25774 16172 25780
rect 16028 25424 16080 25430
rect 16028 25366 16080 25372
rect 15936 23724 15988 23730
rect 15936 23666 15988 23672
rect 15844 21412 15896 21418
rect 15844 21354 15896 21360
rect 15856 21010 15884 21354
rect 15844 21004 15896 21010
rect 15844 20946 15896 20952
rect 15752 20528 15804 20534
rect 15752 20470 15804 20476
rect 15948 19378 15976 23666
rect 16132 23644 16160 25774
rect 16212 24676 16264 24682
rect 16212 24618 16264 24624
rect 16224 24410 16252 24618
rect 16212 24404 16264 24410
rect 16212 24346 16264 24352
rect 16212 23656 16264 23662
rect 16132 23616 16212 23644
rect 16212 23598 16264 23604
rect 16224 22438 16252 23598
rect 16120 22432 16172 22438
rect 16120 22374 16172 22380
rect 16212 22432 16264 22438
rect 16212 22374 16264 22380
rect 16028 21616 16080 21622
rect 16028 21558 16080 21564
rect 16040 19922 16068 21558
rect 16132 21486 16160 22374
rect 16120 21480 16172 21486
rect 16120 21422 16172 21428
rect 16212 21344 16264 21350
rect 16212 21286 16264 21292
rect 16028 19916 16080 19922
rect 16028 19858 16080 19864
rect 15936 19372 15988 19378
rect 15936 19314 15988 19320
rect 16040 18834 16068 19858
rect 16028 18828 16080 18834
rect 16028 18770 16080 18776
rect 16120 18284 16172 18290
rect 16120 18226 16172 18232
rect 15580 17870 15700 17898
rect 15476 17604 15528 17610
rect 15476 17546 15528 17552
rect 15292 16516 15344 16522
rect 15292 16458 15344 16464
rect 15290 15056 15346 15065
rect 15290 14991 15292 15000
rect 15344 14991 15346 15000
rect 15292 14962 15344 14968
rect 15292 14000 15344 14006
rect 15292 13942 15344 13948
rect 15304 12850 15332 13942
rect 15476 13456 15528 13462
rect 15476 13398 15528 13404
rect 15384 13184 15436 13190
rect 15384 13126 15436 13132
rect 15292 12844 15344 12850
rect 15292 12786 15344 12792
rect 15292 12708 15344 12714
rect 15292 12650 15344 12656
rect 15304 11082 15332 12650
rect 15396 11830 15424 13126
rect 15384 11824 15436 11830
rect 15384 11766 15436 11772
rect 15488 11694 15516 13398
rect 15580 12442 15608 17870
rect 16132 17746 16160 18226
rect 15660 17740 15712 17746
rect 15660 17682 15712 17688
rect 16120 17740 16172 17746
rect 16120 17682 16172 17688
rect 15568 12436 15620 12442
rect 15568 12378 15620 12384
rect 15568 11824 15620 11830
rect 15568 11766 15620 11772
rect 15384 11688 15436 11694
rect 15384 11630 15436 11636
rect 15476 11688 15528 11694
rect 15476 11630 15528 11636
rect 15292 11076 15344 11082
rect 15292 11018 15344 11024
rect 15200 8560 15252 8566
rect 15200 8502 15252 8508
rect 15200 8084 15252 8090
rect 15200 8026 15252 8032
rect 14924 7880 14976 7886
rect 14924 7822 14976 7828
rect 14556 7404 14608 7410
rect 14556 7346 14608 7352
rect 14464 6792 14516 6798
rect 14464 6734 14516 6740
rect 14476 6322 14504 6734
rect 14740 6384 14792 6390
rect 14740 6326 14792 6332
rect 14464 6316 14516 6322
rect 14464 6258 14516 6264
rect 14556 6112 14608 6118
rect 14556 6054 14608 6060
rect 14752 6100 14780 6326
rect 14832 6112 14884 6118
rect 14752 6072 14832 6100
rect 14280 5160 14332 5166
rect 13726 5128 13782 5137
rect 14280 5102 14332 5108
rect 13726 5063 13782 5072
rect 14292 4826 14320 5102
rect 14280 4820 14332 4826
rect 14280 4762 14332 4768
rect 14568 4690 14596 6054
rect 14648 5568 14700 5574
rect 14648 5510 14700 5516
rect 14660 5166 14688 5510
rect 14648 5160 14700 5166
rect 14648 5102 14700 5108
rect 14556 4684 14608 4690
rect 14556 4626 14608 4632
rect 14752 4622 14780 6072
rect 14832 6054 14884 6060
rect 15016 5636 15068 5642
rect 15016 5578 15068 5584
rect 14740 4616 14792 4622
rect 14740 4558 14792 4564
rect 13452 4548 13504 4554
rect 13452 4490 13504 4496
rect 13464 3738 13492 4490
rect 13820 4480 13872 4486
rect 13820 4422 13872 4428
rect 13832 4214 13860 4422
rect 13820 4208 13872 4214
rect 13820 4150 13872 4156
rect 14752 4078 14780 4558
rect 15028 4146 15056 5578
rect 15212 5166 15240 8026
rect 15396 6730 15424 11630
rect 15580 11218 15608 11766
rect 15568 11212 15620 11218
rect 15488 11172 15568 11200
rect 15488 10470 15516 11172
rect 15568 11154 15620 11160
rect 15568 10600 15620 10606
rect 15568 10542 15620 10548
rect 15476 10464 15528 10470
rect 15476 10406 15528 10412
rect 15488 9042 15516 10406
rect 15580 9217 15608 10542
rect 15566 9208 15622 9217
rect 15672 9178 15700 17682
rect 16120 17264 16172 17270
rect 16120 17206 16172 17212
rect 16132 17134 16160 17206
rect 16120 17128 16172 17134
rect 16120 17070 16172 17076
rect 16120 16992 16172 16998
rect 16120 16934 16172 16940
rect 16132 16658 16160 16934
rect 16120 16652 16172 16658
rect 16120 16594 16172 16600
rect 16120 16244 16172 16250
rect 16120 16186 16172 16192
rect 16028 16040 16080 16046
rect 16028 15982 16080 15988
rect 16040 15706 16068 15982
rect 16028 15700 16080 15706
rect 16028 15642 16080 15648
rect 16132 15586 16160 16186
rect 16040 15558 16160 15586
rect 15752 14476 15804 14482
rect 15752 14418 15804 14424
rect 15764 12782 15792 14418
rect 15844 14408 15896 14414
rect 15844 14350 15896 14356
rect 15752 12776 15804 12782
rect 15752 12718 15804 12724
rect 15764 12646 15792 12718
rect 15752 12640 15804 12646
rect 15752 12582 15804 12588
rect 15856 11234 15884 14350
rect 16040 13394 16068 15558
rect 16120 14476 16172 14482
rect 16120 14418 16172 14424
rect 16028 13388 16080 13394
rect 16028 13330 16080 13336
rect 16132 12850 16160 14418
rect 16120 12844 16172 12850
rect 16120 12786 16172 12792
rect 16120 12232 16172 12238
rect 16120 12174 16172 12180
rect 15936 11688 15988 11694
rect 15936 11630 15988 11636
rect 15764 11206 15884 11234
rect 15764 10690 15792 11206
rect 15844 11144 15896 11150
rect 15844 11086 15896 11092
rect 15856 10849 15884 11086
rect 15842 10840 15898 10849
rect 15842 10775 15844 10784
rect 15896 10775 15898 10784
rect 15844 10746 15896 10752
rect 15764 10662 15884 10690
rect 15752 10124 15804 10130
rect 15752 10066 15804 10072
rect 15764 9722 15792 10066
rect 15752 9716 15804 9722
rect 15752 9658 15804 9664
rect 15856 9602 15884 10662
rect 15764 9574 15884 9602
rect 15566 9143 15622 9152
rect 15660 9172 15712 9178
rect 15660 9114 15712 9120
rect 15476 9036 15528 9042
rect 15476 8978 15528 8984
rect 15488 8498 15516 8978
rect 15476 8492 15528 8498
rect 15476 8434 15528 8440
rect 15764 8090 15792 9574
rect 15844 9036 15896 9042
rect 15844 8978 15896 8984
rect 15856 8634 15884 8978
rect 15948 8838 15976 11630
rect 16028 11212 16080 11218
rect 16028 11154 16080 11160
rect 16040 9994 16068 11154
rect 16028 9988 16080 9994
rect 16028 9930 16080 9936
rect 15936 8832 15988 8838
rect 15936 8774 15988 8780
rect 15844 8628 15896 8634
rect 15844 8570 15896 8576
rect 15844 8288 15896 8294
rect 15844 8230 15896 8236
rect 15752 8084 15804 8090
rect 15752 8026 15804 8032
rect 15660 7948 15712 7954
rect 15660 7890 15712 7896
rect 15568 7812 15620 7818
rect 15568 7754 15620 7760
rect 15580 7410 15608 7754
rect 15568 7404 15620 7410
rect 15568 7346 15620 7352
rect 15568 7200 15620 7206
rect 15568 7142 15620 7148
rect 15580 6934 15608 7142
rect 15568 6928 15620 6934
rect 15568 6870 15620 6876
rect 15476 6860 15528 6866
rect 15476 6802 15528 6808
rect 15384 6724 15436 6730
rect 15384 6666 15436 6672
rect 15292 6656 15344 6662
rect 15292 6598 15344 6604
rect 15304 6458 15332 6598
rect 15292 6452 15344 6458
rect 15292 6394 15344 6400
rect 15200 5160 15252 5166
rect 15200 5102 15252 5108
rect 15488 4146 15516 6802
rect 15568 6792 15620 6798
rect 15568 6734 15620 6740
rect 15580 6254 15608 6734
rect 15568 6248 15620 6254
rect 15568 6190 15620 6196
rect 15672 5896 15700 7890
rect 15764 7410 15792 8026
rect 15752 7404 15804 7410
rect 15752 7346 15804 7352
rect 15856 6866 15884 8230
rect 15948 7546 15976 8774
rect 16132 8634 16160 12174
rect 16224 11354 16252 21286
rect 16316 20754 16344 30246
rect 16408 30054 16436 30738
rect 16592 30716 16620 31826
rect 16684 31686 16712 32302
rect 16764 32292 16816 32298
rect 16764 32234 16816 32240
rect 16776 31958 16804 32234
rect 16764 31952 16816 31958
rect 16764 31894 16816 31900
rect 16868 31890 16896 32710
rect 16960 32366 16988 32846
rect 16948 32360 17000 32366
rect 16948 32302 17000 32308
rect 16856 31884 16908 31890
rect 16856 31826 16908 31832
rect 16672 31680 16724 31686
rect 16672 31622 16724 31628
rect 16868 31346 16896 31826
rect 16856 31340 16908 31346
rect 16856 31282 16908 31288
rect 16764 31136 16816 31142
rect 16764 31078 16816 31084
rect 16776 30870 16804 31078
rect 16764 30864 16816 30870
rect 16764 30806 16816 30812
rect 16764 30728 16816 30734
rect 16592 30688 16764 30716
rect 16764 30670 16816 30676
rect 16396 30048 16448 30054
rect 16396 29990 16448 29996
rect 16776 29646 16804 30670
rect 16948 30592 17000 30598
rect 16948 30534 17000 30540
rect 16764 29640 16816 29646
rect 16764 29582 16816 29588
rect 16396 26920 16448 26926
rect 16396 26862 16448 26868
rect 16580 26920 16632 26926
rect 16580 26862 16632 26868
rect 16408 21554 16436 26862
rect 16592 26586 16620 26862
rect 16580 26580 16632 26586
rect 16580 26522 16632 26528
rect 16776 26518 16804 29582
rect 16960 28626 16988 30534
rect 17052 30326 17080 36110
rect 17132 35148 17184 35154
rect 17132 35090 17184 35096
rect 17592 35148 17644 35154
rect 17592 35090 17644 35096
rect 17144 33454 17172 35090
rect 17604 34746 17632 35090
rect 17592 34740 17644 34746
rect 17592 34682 17644 34688
rect 17696 34610 17724 39200
rect 19720 37754 19748 39200
rect 21928 39166 21956 39200
rect 21916 39160 21968 39166
rect 21916 39102 21968 39108
rect 23756 39160 23808 39166
rect 23756 39102 23808 39108
rect 19720 37726 20300 37754
rect 19580 37564 19876 37584
rect 19636 37562 19660 37564
rect 19716 37562 19740 37564
rect 19796 37562 19820 37564
rect 19658 37510 19660 37562
rect 19722 37510 19734 37562
rect 19796 37510 19798 37562
rect 19636 37508 19660 37510
rect 19716 37508 19740 37510
rect 19796 37508 19820 37510
rect 19580 37488 19876 37508
rect 18328 36712 18380 36718
rect 18328 36654 18380 36660
rect 18052 36576 18104 36582
rect 18052 36518 18104 36524
rect 18064 36242 18092 36518
rect 18340 36310 18368 36654
rect 19432 36576 19484 36582
rect 19432 36518 19484 36524
rect 20076 36576 20128 36582
rect 20076 36518 20128 36524
rect 18328 36304 18380 36310
rect 18328 36246 18380 36252
rect 19444 36242 19472 36518
rect 19580 36476 19876 36496
rect 19636 36474 19660 36476
rect 19716 36474 19740 36476
rect 19796 36474 19820 36476
rect 19658 36422 19660 36474
rect 19722 36422 19734 36474
rect 19796 36422 19798 36474
rect 19636 36420 19660 36422
rect 19716 36420 19740 36422
rect 19796 36420 19820 36422
rect 19580 36400 19876 36420
rect 20088 36242 20116 36518
rect 18052 36236 18104 36242
rect 18052 36178 18104 36184
rect 19432 36236 19484 36242
rect 19432 36178 19484 36184
rect 20076 36236 20128 36242
rect 20076 36178 20128 36184
rect 19156 36168 19208 36174
rect 19156 36110 19208 36116
rect 19168 35630 19196 36110
rect 19444 35698 19472 36178
rect 19432 35692 19484 35698
rect 19432 35634 19484 35640
rect 17868 35624 17920 35630
rect 17868 35566 17920 35572
rect 19156 35624 19208 35630
rect 19156 35566 19208 35572
rect 17684 34604 17736 34610
rect 17684 34546 17736 34552
rect 17592 33856 17644 33862
rect 17592 33798 17644 33804
rect 17132 33448 17184 33454
rect 17132 33390 17184 33396
rect 17144 32502 17172 33390
rect 17224 33380 17276 33386
rect 17224 33322 17276 33328
rect 17236 32570 17264 33322
rect 17604 32892 17632 33798
rect 17684 32904 17736 32910
rect 17604 32864 17684 32892
rect 17684 32846 17736 32852
rect 17500 32836 17552 32842
rect 17500 32778 17552 32784
rect 17224 32564 17276 32570
rect 17224 32506 17276 32512
rect 17132 32496 17184 32502
rect 17132 32438 17184 32444
rect 17236 32230 17264 32506
rect 17224 32224 17276 32230
rect 17224 32166 17276 32172
rect 17316 30728 17368 30734
rect 17316 30670 17368 30676
rect 17040 30320 17092 30326
rect 17040 30262 17092 30268
rect 17328 30190 17356 30670
rect 17040 30184 17092 30190
rect 17038 30152 17040 30161
rect 17316 30184 17368 30190
rect 17092 30152 17094 30161
rect 17316 30126 17368 30132
rect 17038 30087 17094 30096
rect 17408 30116 17460 30122
rect 17512 30104 17540 32778
rect 17776 32360 17828 32366
rect 17776 32302 17828 32308
rect 17592 31884 17644 31890
rect 17592 31826 17644 31832
rect 17604 31686 17632 31826
rect 17592 31680 17644 31686
rect 17592 31622 17644 31628
rect 17604 30802 17632 31622
rect 17592 30796 17644 30802
rect 17592 30738 17644 30744
rect 17460 30076 17540 30104
rect 17408 30058 17460 30064
rect 17512 29714 17540 30076
rect 17500 29708 17552 29714
rect 17500 29650 17552 29656
rect 17132 29504 17184 29510
rect 17132 29446 17184 29452
rect 17040 29096 17092 29102
rect 17040 29038 17092 29044
rect 17052 28762 17080 29038
rect 17040 28756 17092 28762
rect 17040 28698 17092 28704
rect 16948 28620 17000 28626
rect 16948 28562 17000 28568
rect 17144 28218 17172 29446
rect 17132 28212 17184 28218
rect 17132 28154 17184 28160
rect 17500 28008 17552 28014
rect 17500 27950 17552 27956
rect 17408 27872 17460 27878
rect 17408 27814 17460 27820
rect 16856 27532 16908 27538
rect 16856 27474 16908 27480
rect 16764 26512 16816 26518
rect 16764 26454 16816 26460
rect 16488 26376 16540 26382
rect 16488 26318 16540 26324
rect 16500 24274 16528 26318
rect 16868 25702 16896 27474
rect 17224 27056 17276 27062
rect 17224 26998 17276 27004
rect 16948 26852 17000 26858
rect 16948 26794 17000 26800
rect 16960 25906 16988 26794
rect 16948 25900 17000 25906
rect 16948 25842 17000 25848
rect 16856 25696 16908 25702
rect 16856 25638 16908 25644
rect 16856 25356 16908 25362
rect 16856 25298 16908 25304
rect 16672 25220 16724 25226
rect 16672 25162 16724 25168
rect 16684 24750 16712 25162
rect 16868 25158 16896 25298
rect 16856 25152 16908 25158
rect 16856 25094 16908 25100
rect 16672 24744 16724 24750
rect 16672 24686 16724 24692
rect 17132 24744 17184 24750
rect 17132 24686 17184 24692
rect 16764 24336 16816 24342
rect 16764 24278 16816 24284
rect 16488 24268 16540 24274
rect 16488 24210 16540 24216
rect 16580 23656 16632 23662
rect 16580 23598 16632 23604
rect 16592 23050 16620 23598
rect 16672 23248 16724 23254
rect 16672 23190 16724 23196
rect 16580 23044 16632 23050
rect 16580 22986 16632 22992
rect 16684 22778 16712 23190
rect 16672 22772 16724 22778
rect 16672 22714 16724 22720
rect 16672 22568 16724 22574
rect 16672 22510 16724 22516
rect 16488 21616 16540 21622
rect 16488 21558 16540 21564
rect 16396 21548 16448 21554
rect 16396 21490 16448 21496
rect 16500 21350 16528 21558
rect 16488 21344 16540 21350
rect 16488 21286 16540 21292
rect 16316 20726 16528 20754
rect 16304 20392 16356 20398
rect 16304 20334 16356 20340
rect 16316 19990 16344 20334
rect 16304 19984 16356 19990
rect 16304 19926 16356 19932
rect 16500 19310 16528 20726
rect 16396 19304 16448 19310
rect 16396 19246 16448 19252
rect 16488 19304 16540 19310
rect 16488 19246 16540 19252
rect 16408 18426 16436 19246
rect 16396 18420 16448 18426
rect 16396 18362 16448 18368
rect 16396 16652 16448 16658
rect 16396 16594 16448 16600
rect 16488 16652 16540 16658
rect 16488 16594 16540 16600
rect 16304 15700 16356 15706
rect 16304 15642 16356 15648
rect 16316 15434 16344 15642
rect 16304 15428 16356 15434
rect 16304 15370 16356 15376
rect 16408 12782 16436 16594
rect 16500 15502 16528 16594
rect 16488 15496 16540 15502
rect 16488 15438 16540 15444
rect 16500 14074 16528 15438
rect 16580 15428 16632 15434
rect 16580 15370 16632 15376
rect 16592 15026 16620 15370
rect 16580 15020 16632 15026
rect 16580 14962 16632 14968
rect 16488 14068 16540 14074
rect 16488 14010 16540 14016
rect 16684 12918 16712 22510
rect 16776 21078 16804 24278
rect 16948 24268 17000 24274
rect 16948 24210 17000 24216
rect 16960 22710 16988 24210
rect 17144 23798 17172 24686
rect 17236 24206 17264 26998
rect 17420 26382 17448 27814
rect 17512 26432 17540 27950
rect 17604 26994 17632 30738
rect 17788 30161 17816 32302
rect 17774 30152 17830 30161
rect 17774 30087 17830 30096
rect 17684 28620 17736 28626
rect 17684 28562 17736 28568
rect 17696 28082 17724 28562
rect 17684 28076 17736 28082
rect 17684 28018 17736 28024
rect 17696 27062 17724 28018
rect 17684 27056 17736 27062
rect 17684 26998 17736 27004
rect 17592 26988 17644 26994
rect 17592 26930 17644 26936
rect 17776 26784 17828 26790
rect 17776 26726 17828 26732
rect 17592 26444 17644 26450
rect 17512 26404 17592 26432
rect 17592 26386 17644 26392
rect 17408 26376 17460 26382
rect 17408 26318 17460 26324
rect 17316 26308 17368 26314
rect 17316 26250 17368 26256
rect 17328 25362 17356 26250
rect 17420 25770 17448 26318
rect 17604 26246 17632 26386
rect 17592 26240 17644 26246
rect 17592 26182 17644 26188
rect 17408 25764 17460 25770
rect 17408 25706 17460 25712
rect 17316 25356 17368 25362
rect 17316 25298 17368 25304
rect 17604 25158 17632 26182
rect 17788 25974 17816 26726
rect 17776 25968 17828 25974
rect 17776 25910 17828 25916
rect 17592 25152 17644 25158
rect 17592 25094 17644 25100
rect 17224 24200 17276 24206
rect 17224 24142 17276 24148
rect 17132 23792 17184 23798
rect 17132 23734 17184 23740
rect 17132 23656 17184 23662
rect 17132 23598 17184 23604
rect 17144 23322 17172 23598
rect 17408 23588 17460 23594
rect 17408 23530 17460 23536
rect 17132 23316 17184 23322
rect 17132 23258 17184 23264
rect 17224 22772 17276 22778
rect 17224 22714 17276 22720
rect 16948 22704 17000 22710
rect 16948 22646 17000 22652
rect 17040 22092 17092 22098
rect 17040 22034 17092 22040
rect 17052 21690 17080 22034
rect 17236 22030 17264 22714
rect 17224 22024 17276 22030
rect 17224 21966 17276 21972
rect 17040 21684 17092 21690
rect 17040 21626 17092 21632
rect 17040 21480 17092 21486
rect 17040 21422 17092 21428
rect 17052 21078 17080 21422
rect 16764 21072 16816 21078
rect 16764 21014 16816 21020
rect 17040 21072 17092 21078
rect 17040 21014 17092 21020
rect 17052 20398 17080 21014
rect 17236 21010 17264 21966
rect 17224 21004 17276 21010
rect 17224 20946 17276 20952
rect 17236 20806 17264 20946
rect 17224 20800 17276 20806
rect 17224 20742 17276 20748
rect 17040 20392 17092 20398
rect 17040 20334 17092 20340
rect 17316 20256 17368 20262
rect 17316 20198 17368 20204
rect 16764 19712 16816 19718
rect 16764 19654 16816 19660
rect 16776 18902 16804 19654
rect 17328 19378 17356 20198
rect 17316 19372 17368 19378
rect 17316 19314 17368 19320
rect 16948 19236 17000 19242
rect 16948 19178 17000 19184
rect 17132 19236 17184 19242
rect 17132 19178 17184 19184
rect 16764 18896 16816 18902
rect 16764 18838 16816 18844
rect 16960 18222 16988 19178
rect 17144 18834 17172 19178
rect 17132 18828 17184 18834
rect 17132 18770 17184 18776
rect 16948 18216 17000 18222
rect 16948 18158 17000 18164
rect 17132 18216 17184 18222
rect 17132 18158 17184 18164
rect 17144 17134 17172 18158
rect 17328 17746 17356 19314
rect 17224 17740 17276 17746
rect 17224 17682 17276 17688
rect 17316 17740 17368 17746
rect 17316 17682 17368 17688
rect 17132 17128 17184 17134
rect 17132 17070 17184 17076
rect 16948 16448 17000 16454
rect 16948 16390 17000 16396
rect 16856 15904 16908 15910
rect 16856 15846 16908 15852
rect 16764 15428 16816 15434
rect 16764 15370 16816 15376
rect 16776 15162 16804 15370
rect 16764 15156 16816 15162
rect 16764 15098 16816 15104
rect 16764 15020 16816 15026
rect 16764 14962 16816 14968
rect 16776 14278 16804 14962
rect 16764 14272 16816 14278
rect 16764 14214 16816 14220
rect 16672 12912 16724 12918
rect 16672 12854 16724 12860
rect 16764 12912 16816 12918
rect 16764 12854 16816 12860
rect 16396 12776 16448 12782
rect 16776 12753 16804 12854
rect 16396 12718 16448 12724
rect 16762 12744 16818 12753
rect 16408 12374 16436 12718
rect 16762 12679 16818 12688
rect 16396 12368 16448 12374
rect 16396 12310 16448 12316
rect 16408 11694 16436 12310
rect 16396 11688 16448 11694
rect 16396 11630 16448 11636
rect 16212 11348 16264 11354
rect 16212 11290 16264 11296
rect 16672 11144 16724 11150
rect 16672 11086 16724 11092
rect 16580 10736 16632 10742
rect 16580 10678 16632 10684
rect 16210 10160 16266 10169
rect 16210 10095 16212 10104
rect 16264 10095 16266 10104
rect 16212 10066 16264 10072
rect 16592 9654 16620 10678
rect 16684 10198 16712 11086
rect 16868 10810 16896 15846
rect 16960 15570 16988 16390
rect 16948 15564 17000 15570
rect 17000 15524 17080 15552
rect 16948 15506 17000 15512
rect 16946 15192 17002 15201
rect 17052 15162 17080 15524
rect 17132 15496 17184 15502
rect 17132 15438 17184 15444
rect 16946 15127 17002 15136
rect 17040 15156 17092 15162
rect 16960 15094 16988 15127
rect 17040 15098 17092 15104
rect 16948 15088 17000 15094
rect 16948 15030 17000 15036
rect 16948 14272 17000 14278
rect 16948 14214 17000 14220
rect 16960 13190 16988 14214
rect 17144 14074 17172 15438
rect 17132 14068 17184 14074
rect 17132 14010 17184 14016
rect 17144 13394 17172 14010
rect 17132 13388 17184 13394
rect 17132 13330 17184 13336
rect 16948 13184 17000 13190
rect 16948 13126 17000 13132
rect 16856 10804 16908 10810
rect 16856 10746 16908 10752
rect 17236 10742 17264 17682
rect 17316 17128 17368 17134
rect 17316 17070 17368 17076
rect 17328 16046 17356 17070
rect 17316 16040 17368 16046
rect 17316 15982 17368 15988
rect 17316 13728 17368 13734
rect 17316 13670 17368 13676
rect 17328 13326 17356 13670
rect 17316 13320 17368 13326
rect 17316 13262 17368 13268
rect 17316 12096 17368 12102
rect 17316 12038 17368 12044
rect 17328 11762 17356 12038
rect 17420 11830 17448 23530
rect 17500 22568 17552 22574
rect 17500 22510 17552 22516
rect 17512 22234 17540 22510
rect 17880 22250 17908 35566
rect 18972 35556 19024 35562
rect 18972 35498 19024 35504
rect 18880 35284 18932 35290
rect 18880 35226 18932 35232
rect 18052 34536 18104 34542
rect 18052 34478 18104 34484
rect 18144 34536 18196 34542
rect 18144 34478 18196 34484
rect 18064 33658 18092 34478
rect 18052 33652 18104 33658
rect 18052 33594 18104 33600
rect 18156 32434 18184 34478
rect 18696 34468 18748 34474
rect 18696 34410 18748 34416
rect 18708 34066 18736 34410
rect 18696 34060 18748 34066
rect 18696 34002 18748 34008
rect 18420 33856 18472 33862
rect 18420 33798 18472 33804
rect 18432 33454 18460 33798
rect 18420 33448 18472 33454
rect 18420 33390 18472 33396
rect 18432 32570 18460 33390
rect 18512 32768 18564 32774
rect 18512 32710 18564 32716
rect 18788 32768 18840 32774
rect 18788 32710 18840 32716
rect 18420 32564 18472 32570
rect 18420 32506 18472 32512
rect 18144 32428 18196 32434
rect 18144 32370 18196 32376
rect 18236 32224 18288 32230
rect 18236 32166 18288 32172
rect 18248 31890 18276 32166
rect 18328 31952 18380 31958
rect 18328 31894 18380 31900
rect 18236 31884 18288 31890
rect 18236 31826 18288 31832
rect 18340 31822 18368 31894
rect 18328 31816 18380 31822
rect 18328 31758 18380 31764
rect 18432 31260 18460 32506
rect 18524 31958 18552 32710
rect 18800 32434 18828 32710
rect 18788 32428 18840 32434
rect 18788 32370 18840 32376
rect 18604 32360 18656 32366
rect 18604 32302 18656 32308
rect 18512 31952 18564 31958
rect 18512 31894 18564 31900
rect 18616 31822 18644 32302
rect 18604 31816 18656 31822
rect 18604 31758 18656 31764
rect 18800 31278 18828 32370
rect 18604 31272 18656 31278
rect 18432 31232 18604 31260
rect 18604 31214 18656 31220
rect 18788 31272 18840 31278
rect 18788 31214 18840 31220
rect 17960 30796 18012 30802
rect 17960 30738 18012 30744
rect 18512 30796 18564 30802
rect 18512 30738 18564 30744
rect 17972 29782 18000 30738
rect 18524 30258 18552 30738
rect 18512 30252 18564 30258
rect 18512 30194 18564 30200
rect 18052 30184 18104 30190
rect 18052 30126 18104 30132
rect 17960 29776 18012 29782
rect 17960 29718 18012 29724
rect 18064 29594 18092 30126
rect 17972 29578 18092 29594
rect 18236 29640 18288 29646
rect 18236 29582 18288 29588
rect 17960 29572 18092 29578
rect 18012 29566 18092 29572
rect 17960 29514 18012 29520
rect 18064 28014 18092 29566
rect 18248 29306 18276 29582
rect 18236 29300 18288 29306
rect 18236 29242 18288 29248
rect 18052 28008 18104 28014
rect 18052 27950 18104 27956
rect 18248 27538 18276 29242
rect 18328 28620 18380 28626
rect 18328 28562 18380 28568
rect 18340 28150 18368 28562
rect 18420 28552 18472 28558
rect 18420 28494 18472 28500
rect 18328 28144 18380 28150
rect 18328 28086 18380 28092
rect 18432 28014 18460 28494
rect 18420 28008 18472 28014
rect 18420 27950 18472 27956
rect 18236 27532 18288 27538
rect 18236 27474 18288 27480
rect 18328 26784 18380 26790
rect 18328 26726 18380 26732
rect 18052 26444 18104 26450
rect 18052 26386 18104 26392
rect 17960 25764 18012 25770
rect 17960 25706 18012 25712
rect 17972 25362 18000 25706
rect 18064 25498 18092 26386
rect 18236 26240 18288 26246
rect 18236 26182 18288 26188
rect 18248 25906 18276 26182
rect 18340 26042 18368 26726
rect 18432 26314 18460 27950
rect 18420 26308 18472 26314
rect 18420 26250 18472 26256
rect 18328 26036 18380 26042
rect 18328 25978 18380 25984
rect 18236 25900 18288 25906
rect 18236 25842 18288 25848
rect 18432 25838 18460 26250
rect 18616 25906 18644 31214
rect 18604 25900 18656 25906
rect 18604 25842 18656 25848
rect 18420 25832 18472 25838
rect 18420 25774 18472 25780
rect 18052 25492 18104 25498
rect 18052 25434 18104 25440
rect 17960 25356 18012 25362
rect 17960 25298 18012 25304
rect 18064 24886 18092 25434
rect 18052 24880 18104 24886
rect 18052 24822 18104 24828
rect 18800 24750 18828 31214
rect 18788 24744 18840 24750
rect 18788 24686 18840 24692
rect 18144 24676 18196 24682
rect 18144 24618 18196 24624
rect 18156 24274 18184 24618
rect 18892 24562 18920 35226
rect 18984 34066 19012 35498
rect 19168 35290 19196 35566
rect 19580 35388 19876 35408
rect 19636 35386 19660 35388
rect 19716 35386 19740 35388
rect 19796 35386 19820 35388
rect 19658 35334 19660 35386
rect 19722 35334 19734 35386
rect 19796 35334 19798 35386
rect 19636 35332 19660 35334
rect 19716 35332 19740 35334
rect 19796 35332 19820 35334
rect 19580 35312 19876 35332
rect 19156 35284 19208 35290
rect 19156 35226 19208 35232
rect 19064 34944 19116 34950
rect 19064 34886 19116 34892
rect 18972 34060 19024 34066
rect 18972 34002 19024 34008
rect 18972 30048 19024 30054
rect 18972 29990 19024 29996
rect 18984 29102 19012 29990
rect 18972 29096 19024 29102
rect 18972 29038 19024 29044
rect 18972 26920 19024 26926
rect 18972 26862 19024 26868
rect 18984 26450 19012 26862
rect 18972 26444 19024 26450
rect 18972 26386 19024 26392
rect 18972 24880 19024 24886
rect 18972 24822 19024 24828
rect 18984 24750 19012 24822
rect 18972 24744 19024 24750
rect 18972 24686 19024 24692
rect 18800 24534 18920 24562
rect 18144 24268 18196 24274
rect 18144 24210 18196 24216
rect 18512 23656 18564 23662
rect 18512 23598 18564 23604
rect 18524 23186 18552 23598
rect 18512 23180 18564 23186
rect 18512 23122 18564 23128
rect 17500 22228 17552 22234
rect 17880 22222 18000 22250
rect 17500 22170 17552 22176
rect 17776 21956 17828 21962
rect 17776 21898 17828 21904
rect 17592 21684 17644 21690
rect 17592 21626 17644 21632
rect 17604 19922 17632 21626
rect 17788 21010 17816 21898
rect 17972 21570 18000 22222
rect 18418 21992 18474 22001
rect 18418 21927 18474 21936
rect 17880 21542 18000 21570
rect 17776 21004 17828 21010
rect 17776 20946 17828 20952
rect 17880 20890 17908 21542
rect 17960 21480 18012 21486
rect 17960 21422 18012 21428
rect 17788 20862 17908 20890
rect 17684 20324 17736 20330
rect 17684 20266 17736 20272
rect 17592 19916 17644 19922
rect 17592 19858 17644 19864
rect 17696 17610 17724 20266
rect 17788 18680 17816 20862
rect 17868 20256 17920 20262
rect 17868 20198 17920 20204
rect 17880 20058 17908 20198
rect 17868 20052 17920 20058
rect 17868 19994 17920 20000
rect 17880 19310 17908 19994
rect 17868 19304 17920 19310
rect 17868 19246 17920 19252
rect 17972 18970 18000 21422
rect 18432 21010 18460 21927
rect 18524 21486 18552 23122
rect 18800 21962 18828 24534
rect 18880 23248 18932 23254
rect 18880 23190 18932 23196
rect 18892 22098 18920 23190
rect 18984 22982 19012 24686
rect 19076 23186 19104 34886
rect 19168 33114 19196 35226
rect 19248 34604 19300 34610
rect 19248 34546 19300 34552
rect 19260 34066 19288 34546
rect 19580 34300 19876 34320
rect 19636 34298 19660 34300
rect 19716 34298 19740 34300
rect 19796 34298 19820 34300
rect 19658 34246 19660 34298
rect 19722 34246 19734 34298
rect 19796 34246 19798 34298
rect 19636 34244 19660 34246
rect 19716 34244 19740 34246
rect 19796 34244 19820 34246
rect 19580 34224 19876 34244
rect 19248 34060 19300 34066
rect 19248 34002 19300 34008
rect 19340 33448 19392 33454
rect 19340 33390 19392 33396
rect 19432 33448 19484 33454
rect 19432 33390 19484 33396
rect 19156 33108 19208 33114
rect 19156 33050 19208 33056
rect 19352 32774 19380 33390
rect 19340 32768 19392 32774
rect 19340 32710 19392 32716
rect 19444 32008 19472 33390
rect 19984 33380 20036 33386
rect 19984 33322 20036 33328
rect 19580 33212 19876 33232
rect 19636 33210 19660 33212
rect 19716 33210 19740 33212
rect 19796 33210 19820 33212
rect 19658 33158 19660 33210
rect 19722 33158 19734 33210
rect 19796 33158 19798 33210
rect 19636 33156 19660 33158
rect 19716 33156 19740 33158
rect 19796 33156 19820 33158
rect 19580 33136 19876 33156
rect 19996 32978 20024 33322
rect 20076 33312 20128 33318
rect 20076 33254 20128 33260
rect 19984 32972 20036 32978
rect 19984 32914 20036 32920
rect 20088 32366 20116 33254
rect 19892 32360 19944 32366
rect 19892 32302 19944 32308
rect 20076 32360 20128 32366
rect 20076 32302 20128 32308
rect 19580 32124 19876 32144
rect 19636 32122 19660 32124
rect 19716 32122 19740 32124
rect 19796 32122 19820 32124
rect 19658 32070 19660 32122
rect 19722 32070 19734 32122
rect 19796 32070 19798 32122
rect 19636 32068 19660 32070
rect 19716 32068 19740 32070
rect 19796 32068 19820 32070
rect 19580 32048 19876 32068
rect 19444 31980 19564 32008
rect 19156 31748 19208 31754
rect 19156 31690 19208 31696
rect 19168 30870 19196 31690
rect 19536 31634 19564 31980
rect 19352 31606 19564 31634
rect 19156 30864 19208 30870
rect 19156 30806 19208 30812
rect 19168 29782 19196 30806
rect 19352 30274 19380 31606
rect 19580 31036 19876 31056
rect 19636 31034 19660 31036
rect 19716 31034 19740 31036
rect 19796 31034 19820 31036
rect 19658 30982 19660 31034
rect 19722 30982 19734 31034
rect 19796 30982 19798 31034
rect 19636 30980 19660 30982
rect 19716 30980 19740 30982
rect 19796 30980 19820 30982
rect 19580 30960 19876 30980
rect 19432 30796 19484 30802
rect 19432 30738 19484 30744
rect 19260 30246 19380 30274
rect 19156 29776 19208 29782
rect 19156 29718 19208 29724
rect 19156 29028 19208 29034
rect 19156 28970 19208 28976
rect 19168 28914 19196 28970
rect 19260 28914 19288 30246
rect 19444 30190 19472 30738
rect 19432 30184 19484 30190
rect 19432 30126 19484 30132
rect 19340 30116 19392 30122
rect 19340 30058 19392 30064
rect 19352 29170 19380 30058
rect 19444 29510 19472 30126
rect 19580 29948 19876 29968
rect 19636 29946 19660 29948
rect 19716 29946 19740 29948
rect 19796 29946 19820 29948
rect 19658 29894 19660 29946
rect 19722 29894 19734 29946
rect 19796 29894 19798 29946
rect 19636 29892 19660 29894
rect 19716 29892 19740 29894
rect 19796 29892 19820 29894
rect 19580 29872 19876 29892
rect 19706 29608 19762 29617
rect 19706 29543 19708 29552
rect 19760 29543 19762 29552
rect 19800 29572 19852 29578
rect 19708 29514 19760 29520
rect 19800 29514 19852 29520
rect 19432 29504 19484 29510
rect 19432 29446 19484 29452
rect 19444 29238 19472 29446
rect 19812 29306 19840 29514
rect 19800 29300 19852 29306
rect 19800 29242 19852 29248
rect 19432 29232 19484 29238
rect 19432 29174 19484 29180
rect 19340 29164 19392 29170
rect 19340 29106 19392 29112
rect 19812 29102 19840 29242
rect 19800 29096 19852 29102
rect 19800 29038 19852 29044
rect 19168 28886 19380 28914
rect 19352 27690 19380 28886
rect 19580 28860 19876 28880
rect 19636 28858 19660 28860
rect 19716 28858 19740 28860
rect 19796 28858 19820 28860
rect 19658 28806 19660 28858
rect 19722 28806 19734 28858
rect 19796 28806 19798 28858
rect 19636 28804 19660 28806
rect 19716 28804 19740 28806
rect 19796 28804 19820 28806
rect 19580 28784 19876 28804
rect 19904 28626 19932 32302
rect 20076 32020 20128 32026
rect 20076 31962 20128 31968
rect 20088 31890 20116 31962
rect 20076 31884 20128 31890
rect 20076 31826 20128 31832
rect 19984 31272 20036 31278
rect 19984 31214 20036 31220
rect 19996 30190 20024 31214
rect 19984 30184 20036 30190
rect 19984 30126 20036 30132
rect 20088 30054 20116 31826
rect 20272 31414 20300 37726
rect 21272 37324 21324 37330
rect 21272 37266 21324 37272
rect 21284 36718 21312 37266
rect 20812 36712 20864 36718
rect 20812 36654 20864 36660
rect 21272 36712 21324 36718
rect 21272 36654 21324 36660
rect 21548 36712 21600 36718
rect 21548 36654 21600 36660
rect 23020 36712 23072 36718
rect 23020 36654 23072 36660
rect 20824 36242 20852 36654
rect 20812 36236 20864 36242
rect 20812 36178 20864 36184
rect 20824 35834 20852 36178
rect 21284 35834 21312 36654
rect 21560 36378 21588 36654
rect 21548 36372 21600 36378
rect 21548 36314 21600 36320
rect 23032 36174 23060 36654
rect 23296 36644 23348 36650
rect 23296 36586 23348 36592
rect 23308 36242 23336 36586
rect 23296 36236 23348 36242
rect 23296 36178 23348 36184
rect 23020 36168 23072 36174
rect 23020 36110 23072 36116
rect 20812 35828 20864 35834
rect 20812 35770 20864 35776
rect 21272 35828 21324 35834
rect 21272 35770 21324 35776
rect 23032 35766 23060 36110
rect 23020 35760 23072 35766
rect 23020 35702 23072 35708
rect 21548 35624 21600 35630
rect 21548 35566 21600 35572
rect 20812 35556 20864 35562
rect 20812 35498 20864 35504
rect 20824 35086 20852 35498
rect 21560 35290 21588 35566
rect 22652 35556 22704 35562
rect 22652 35498 22704 35504
rect 21548 35284 21600 35290
rect 21548 35226 21600 35232
rect 22664 35154 22692 35498
rect 20996 35148 21048 35154
rect 20996 35090 21048 35096
rect 22652 35148 22704 35154
rect 22652 35090 22704 35096
rect 20812 35080 20864 35086
rect 20812 35022 20864 35028
rect 20352 33448 20404 33454
rect 20352 33390 20404 33396
rect 20364 32502 20392 33390
rect 20628 33312 20680 33318
rect 20628 33254 20680 33260
rect 20536 32972 20588 32978
rect 20536 32914 20588 32920
rect 20352 32496 20404 32502
rect 20352 32438 20404 32444
rect 20352 32360 20404 32366
rect 20352 32302 20404 32308
rect 20364 31958 20392 32302
rect 20352 31952 20404 31958
rect 20352 31894 20404 31900
rect 20352 31748 20404 31754
rect 20352 31690 20404 31696
rect 20260 31408 20312 31414
rect 20260 31350 20312 31356
rect 20168 31340 20220 31346
rect 20168 31282 20220 31288
rect 20076 30048 20128 30054
rect 20076 29990 20128 29996
rect 20180 29714 20208 31282
rect 20260 31204 20312 31210
rect 20260 31146 20312 31152
rect 20272 30938 20300 31146
rect 20260 30932 20312 30938
rect 20260 30874 20312 30880
rect 20168 29708 20220 29714
rect 20168 29650 20220 29656
rect 20076 29640 20128 29646
rect 20076 29582 20128 29588
rect 19984 29028 20036 29034
rect 19984 28970 20036 28976
rect 19892 28620 19944 28626
rect 19892 28562 19944 28568
rect 19432 28552 19484 28558
rect 19432 28494 19484 28500
rect 19260 27662 19380 27690
rect 19156 27328 19208 27334
rect 19156 27270 19208 27276
rect 19168 26790 19196 27270
rect 19260 27146 19288 27662
rect 19340 27532 19392 27538
rect 19340 27474 19392 27480
rect 19352 27334 19380 27474
rect 19444 27402 19472 28494
rect 19580 27772 19876 27792
rect 19636 27770 19660 27772
rect 19716 27770 19740 27772
rect 19796 27770 19820 27772
rect 19658 27718 19660 27770
rect 19722 27718 19734 27770
rect 19796 27718 19798 27770
rect 19636 27716 19660 27718
rect 19716 27716 19740 27718
rect 19796 27716 19820 27718
rect 19580 27696 19876 27716
rect 19996 27538 20024 28970
rect 20088 27606 20116 29582
rect 20168 29504 20220 29510
rect 20168 29446 20220 29452
rect 20180 28966 20208 29446
rect 20260 29096 20312 29102
rect 20260 29038 20312 29044
rect 20168 28960 20220 28966
rect 20168 28902 20220 28908
rect 20272 28558 20300 29038
rect 20260 28552 20312 28558
rect 20260 28494 20312 28500
rect 20272 27878 20300 28494
rect 20260 27872 20312 27878
rect 20260 27814 20312 27820
rect 20076 27600 20128 27606
rect 20076 27542 20128 27548
rect 19524 27532 19576 27538
rect 19524 27474 19576 27480
rect 19984 27532 20036 27538
rect 19984 27474 20036 27480
rect 19432 27396 19484 27402
rect 19432 27338 19484 27344
rect 19340 27328 19392 27334
rect 19340 27270 19392 27276
rect 19260 27118 19472 27146
rect 19340 26988 19392 26994
rect 19340 26930 19392 26936
rect 19156 26784 19208 26790
rect 19156 26726 19208 26732
rect 19352 26518 19380 26930
rect 19340 26512 19392 26518
rect 19340 26454 19392 26460
rect 19444 25294 19472 27118
rect 19536 26926 19564 27474
rect 19524 26920 19576 26926
rect 19524 26862 19576 26868
rect 19892 26920 19944 26926
rect 19892 26862 19944 26868
rect 19580 26684 19876 26704
rect 19636 26682 19660 26684
rect 19716 26682 19740 26684
rect 19796 26682 19820 26684
rect 19658 26630 19660 26682
rect 19722 26630 19734 26682
rect 19796 26630 19798 26682
rect 19636 26628 19660 26630
rect 19716 26628 19740 26630
rect 19796 26628 19820 26630
rect 19580 26608 19876 26628
rect 19708 26512 19760 26518
rect 19706 26480 19708 26489
rect 19760 26480 19762 26489
rect 19904 26450 19932 26862
rect 19984 26852 20036 26858
rect 19984 26794 20036 26800
rect 19996 26586 20024 26794
rect 20364 26738 20392 31690
rect 20444 31408 20496 31414
rect 20444 31350 20496 31356
rect 20456 29306 20484 31350
rect 20548 31142 20576 32914
rect 20640 32026 20668 33254
rect 20628 32020 20680 32026
rect 20628 31962 20680 31968
rect 20536 31136 20588 31142
rect 20536 31078 20588 31084
rect 20640 30802 20668 31962
rect 20824 31754 20852 35022
rect 21008 34134 21036 35090
rect 22376 35080 22428 35086
rect 22376 35022 22428 35028
rect 21180 34944 21232 34950
rect 21180 34886 21232 34892
rect 21192 34610 21220 34886
rect 22388 34610 22416 35022
rect 21180 34604 21232 34610
rect 21180 34546 21232 34552
rect 22376 34604 22428 34610
rect 22376 34546 22428 34552
rect 21364 34536 21416 34542
rect 21364 34478 21416 34484
rect 21732 34536 21784 34542
rect 21732 34478 21784 34484
rect 20996 34128 21048 34134
rect 20996 34070 21048 34076
rect 21088 32768 21140 32774
rect 21088 32710 21140 32716
rect 21100 32434 21128 32710
rect 21088 32428 21140 32434
rect 21088 32370 21140 32376
rect 20812 31748 20864 31754
rect 20812 31690 20864 31696
rect 20996 31272 21048 31278
rect 20996 31214 21048 31220
rect 20812 31204 20864 31210
rect 20812 31146 20864 31152
rect 20628 30796 20680 30802
rect 20628 30738 20680 30744
rect 20824 30734 20852 31146
rect 20812 30728 20864 30734
rect 20812 30670 20864 30676
rect 20824 30258 20852 30670
rect 20812 30252 20864 30258
rect 20812 30194 20864 30200
rect 21008 30190 21036 31214
rect 21088 30728 21140 30734
rect 21088 30670 21140 30676
rect 20628 30184 20680 30190
rect 20628 30126 20680 30132
rect 20996 30184 21048 30190
rect 20996 30126 21048 30132
rect 20536 29640 20588 29646
rect 20536 29582 20588 29588
rect 20444 29300 20496 29306
rect 20444 29242 20496 29248
rect 20444 29096 20496 29102
rect 20444 29038 20496 29044
rect 20456 28762 20484 29038
rect 20444 28756 20496 28762
rect 20444 28698 20496 28704
rect 20548 28694 20576 29582
rect 20640 28762 20668 30126
rect 20812 28960 20864 28966
rect 20812 28902 20864 28908
rect 20628 28756 20680 28762
rect 20628 28698 20680 28704
rect 20536 28688 20588 28694
rect 20536 28630 20588 28636
rect 20640 28082 20668 28698
rect 20824 28694 20852 28902
rect 20812 28688 20864 28694
rect 20812 28630 20864 28636
rect 20720 28620 20772 28626
rect 20720 28562 20772 28568
rect 20628 28076 20680 28082
rect 20628 28018 20680 28024
rect 20732 27606 20760 28562
rect 21008 27946 21036 30126
rect 21100 29578 21128 30670
rect 21180 29844 21232 29850
rect 21180 29786 21232 29792
rect 21088 29572 21140 29578
rect 21088 29514 21140 29520
rect 21192 29238 21220 29786
rect 21180 29232 21232 29238
rect 21180 29174 21232 29180
rect 21088 28960 21140 28966
rect 21088 28902 21140 28908
rect 21100 28626 21128 28902
rect 21088 28620 21140 28626
rect 21088 28562 21140 28568
rect 20996 27940 21048 27946
rect 20996 27882 21048 27888
rect 20720 27600 20772 27606
rect 20720 27542 20772 27548
rect 20444 27532 20496 27538
rect 20444 27474 20496 27480
rect 20456 26926 20484 27474
rect 21100 27402 21128 28562
rect 21180 28008 21232 28014
rect 21180 27950 21232 27956
rect 20812 27396 20864 27402
rect 20812 27338 20864 27344
rect 21088 27396 21140 27402
rect 21088 27338 21140 27344
rect 20628 27328 20680 27334
rect 20628 27270 20680 27276
rect 20640 26926 20668 27270
rect 20720 27056 20772 27062
rect 20720 26998 20772 27004
rect 20824 27010 20852 27338
rect 20444 26920 20496 26926
rect 20444 26862 20496 26868
rect 20628 26920 20680 26926
rect 20732 26897 20760 26998
rect 20824 26982 21128 27010
rect 21192 26994 21220 27950
rect 21100 26926 21128 26982
rect 21180 26988 21232 26994
rect 21180 26930 21232 26936
rect 20996 26920 21048 26926
rect 20628 26862 20680 26868
rect 20718 26888 20774 26897
rect 20180 26710 20392 26738
rect 19984 26580 20036 26586
rect 19984 26522 20036 26528
rect 20074 26480 20130 26489
rect 19706 26415 19762 26424
rect 19892 26444 19944 26450
rect 19892 26386 19944 26392
rect 19984 26444 20036 26450
rect 20074 26415 20130 26424
rect 19984 26386 20036 26392
rect 19996 25906 20024 26386
rect 19984 25900 20036 25906
rect 19984 25842 20036 25848
rect 19892 25832 19944 25838
rect 19892 25774 19944 25780
rect 19580 25596 19876 25616
rect 19636 25594 19660 25596
rect 19716 25594 19740 25596
rect 19796 25594 19820 25596
rect 19658 25542 19660 25594
rect 19722 25542 19734 25594
rect 19796 25542 19798 25594
rect 19636 25540 19660 25542
rect 19716 25540 19740 25542
rect 19796 25540 19820 25542
rect 19580 25520 19876 25540
rect 19904 25294 19932 25774
rect 19432 25288 19484 25294
rect 19432 25230 19484 25236
rect 19892 25288 19944 25294
rect 19892 25230 19944 25236
rect 19444 24954 19472 25230
rect 19432 24948 19484 24954
rect 19432 24890 19484 24896
rect 19904 24750 19932 25230
rect 20088 24886 20116 26415
rect 20076 24880 20128 24886
rect 20076 24822 20128 24828
rect 19892 24744 19944 24750
rect 19892 24686 19944 24692
rect 19340 24676 19392 24682
rect 19340 24618 19392 24624
rect 19352 24342 19380 24618
rect 19580 24508 19876 24528
rect 19636 24506 19660 24508
rect 19716 24506 19740 24508
rect 19796 24506 19820 24508
rect 19658 24454 19660 24506
rect 19722 24454 19734 24506
rect 19796 24454 19798 24506
rect 19636 24452 19660 24454
rect 19716 24452 19740 24454
rect 19796 24452 19820 24454
rect 19580 24432 19876 24452
rect 19340 24336 19392 24342
rect 19340 24278 19392 24284
rect 19984 24336 20036 24342
rect 19984 24278 20036 24284
rect 19352 24070 19380 24278
rect 19432 24268 19484 24274
rect 19432 24210 19484 24216
rect 19340 24064 19392 24070
rect 19340 24006 19392 24012
rect 19340 23724 19392 23730
rect 19340 23666 19392 23672
rect 19248 23656 19300 23662
rect 19248 23598 19300 23604
rect 19260 23254 19288 23598
rect 19248 23248 19300 23254
rect 19248 23190 19300 23196
rect 19064 23180 19116 23186
rect 19064 23122 19116 23128
rect 18972 22976 19024 22982
rect 18972 22918 19024 22924
rect 19352 22778 19380 23666
rect 19340 22772 19392 22778
rect 19340 22714 19392 22720
rect 19444 22658 19472 24210
rect 19580 23420 19876 23440
rect 19636 23418 19660 23420
rect 19716 23418 19740 23420
rect 19796 23418 19820 23420
rect 19658 23366 19660 23418
rect 19722 23366 19734 23418
rect 19796 23366 19798 23418
rect 19636 23364 19660 23366
rect 19716 23364 19740 23366
rect 19796 23364 19820 23366
rect 19580 23344 19876 23364
rect 19996 23322 20024 24278
rect 19984 23316 20036 23322
rect 19984 23258 20036 23264
rect 20076 23180 20128 23186
rect 20076 23122 20128 23128
rect 19352 22630 19472 22658
rect 18880 22092 18932 22098
rect 19064 22092 19116 22098
rect 18932 22052 19012 22080
rect 18880 22034 18932 22040
rect 18788 21956 18840 21962
rect 18788 21898 18840 21904
rect 18512 21480 18564 21486
rect 18512 21422 18564 21428
rect 18420 21004 18472 21010
rect 18420 20946 18472 20952
rect 18420 20392 18472 20398
rect 18420 20334 18472 20340
rect 18052 19304 18104 19310
rect 18050 19272 18052 19281
rect 18236 19304 18288 19310
rect 18104 19272 18106 19281
rect 18236 19246 18288 19252
rect 18050 19207 18106 19216
rect 17960 18964 18012 18970
rect 17960 18906 18012 18912
rect 17868 18692 17920 18698
rect 17788 18652 17868 18680
rect 17868 18634 17920 18640
rect 17776 18148 17828 18154
rect 17776 18090 17828 18096
rect 17788 17610 17816 18090
rect 17880 18086 17908 18634
rect 17868 18080 17920 18086
rect 17868 18022 17920 18028
rect 17684 17604 17736 17610
rect 17684 17546 17736 17552
rect 17776 17604 17828 17610
rect 17776 17546 17828 17552
rect 18064 17134 18092 19207
rect 18144 17604 18196 17610
rect 18144 17546 18196 17552
rect 18156 17134 18184 17546
rect 18052 17128 18104 17134
rect 18052 17070 18104 17076
rect 18144 17128 18196 17134
rect 18144 17070 18196 17076
rect 18144 16992 18196 16998
rect 18144 16934 18196 16940
rect 18052 16516 18104 16522
rect 18052 16458 18104 16464
rect 18064 16250 18092 16458
rect 18156 16454 18184 16934
rect 18144 16448 18196 16454
rect 18144 16390 18196 16396
rect 18052 16244 18104 16250
rect 18052 16186 18104 16192
rect 18144 15972 18196 15978
rect 18144 15914 18196 15920
rect 18156 15570 18184 15914
rect 17868 15564 17920 15570
rect 17868 15506 17920 15512
rect 18144 15564 18196 15570
rect 18144 15506 18196 15512
rect 17592 14884 17644 14890
rect 17592 14826 17644 14832
rect 17498 14376 17554 14385
rect 17498 14311 17500 14320
rect 17552 14311 17554 14320
rect 17500 14282 17552 14288
rect 17512 13462 17540 14282
rect 17500 13456 17552 13462
rect 17500 13398 17552 13404
rect 17500 12300 17552 12306
rect 17500 12242 17552 12248
rect 17408 11824 17460 11830
rect 17408 11766 17460 11772
rect 17316 11756 17368 11762
rect 17316 11698 17368 11704
rect 17224 10736 17276 10742
rect 17224 10678 17276 10684
rect 17408 10600 17460 10606
rect 17408 10542 17460 10548
rect 16672 10192 16724 10198
rect 16672 10134 16724 10140
rect 17420 10130 17448 10542
rect 17408 10124 17460 10130
rect 17408 10066 17460 10072
rect 16580 9648 16632 9654
rect 16580 9590 16632 9596
rect 16592 9042 16620 9590
rect 17512 9586 17540 12242
rect 17604 10130 17632 14826
rect 17776 14476 17828 14482
rect 17776 14418 17828 14424
rect 17684 14272 17736 14278
rect 17684 14214 17736 14220
rect 17696 13870 17724 14214
rect 17788 14074 17816 14418
rect 17776 14068 17828 14074
rect 17776 14010 17828 14016
rect 17684 13864 17736 13870
rect 17684 13806 17736 13812
rect 17880 13394 17908 15506
rect 17960 15496 18012 15502
rect 17960 15438 18012 15444
rect 17972 13462 18000 15438
rect 18052 14408 18104 14414
rect 18052 14350 18104 14356
rect 17960 13456 18012 13462
rect 17960 13398 18012 13404
rect 17868 13388 17920 13394
rect 17868 13330 17920 13336
rect 17880 13190 17908 13330
rect 17868 13184 17920 13190
rect 17868 13126 17920 13132
rect 17960 12776 18012 12782
rect 17960 12718 18012 12724
rect 17972 11286 18000 12718
rect 18064 12306 18092 14350
rect 18144 13796 18196 13802
rect 18144 13738 18196 13744
rect 18156 13394 18184 13738
rect 18144 13388 18196 13394
rect 18144 13330 18196 13336
rect 18248 13274 18276 19246
rect 18328 15496 18380 15502
rect 18328 15438 18380 15444
rect 18340 14550 18368 15438
rect 18432 14822 18460 20334
rect 18524 18170 18552 21422
rect 18800 20398 18828 21898
rect 18984 21486 19012 22052
rect 19064 22034 19116 22040
rect 18972 21480 19024 21486
rect 18972 21422 19024 21428
rect 18788 20392 18840 20398
rect 18788 20334 18840 20340
rect 18800 19854 18828 20334
rect 18984 20262 19012 21422
rect 18972 20256 19024 20262
rect 18972 20198 19024 20204
rect 18972 19916 19024 19922
rect 18972 19858 19024 19864
rect 18788 19848 18840 19854
rect 18788 19790 18840 19796
rect 18800 18766 18828 19790
rect 18984 19446 19012 19858
rect 18972 19440 19024 19446
rect 18972 19382 19024 19388
rect 18972 19168 19024 19174
rect 19076 19156 19104 22034
rect 19352 21706 19380 22630
rect 19432 22568 19484 22574
rect 19432 22510 19484 22516
rect 19984 22568 20036 22574
rect 19984 22510 20036 22516
rect 19260 21678 19380 21706
rect 19156 21616 19208 21622
rect 19156 21558 19208 21564
rect 19024 19128 19104 19156
rect 18972 19110 19024 19116
rect 18880 18828 18932 18834
rect 18880 18770 18932 18776
rect 18788 18760 18840 18766
rect 18788 18702 18840 18708
rect 18604 18624 18656 18630
rect 18604 18566 18656 18572
rect 18616 18290 18644 18566
rect 18800 18290 18828 18702
rect 18604 18284 18656 18290
rect 18604 18226 18656 18232
rect 18788 18284 18840 18290
rect 18788 18226 18840 18232
rect 18524 18142 18644 18170
rect 18616 17814 18644 18142
rect 18604 17808 18656 17814
rect 18604 17750 18656 17756
rect 18512 17060 18564 17066
rect 18512 17002 18564 17008
rect 18524 16658 18552 17002
rect 18512 16652 18564 16658
rect 18512 16594 18564 16600
rect 18420 14816 18472 14822
rect 18420 14758 18472 14764
rect 18328 14544 18380 14550
rect 18328 14486 18380 14492
rect 18512 13932 18564 13938
rect 18512 13874 18564 13880
rect 18328 13864 18380 13870
rect 18328 13806 18380 13812
rect 18340 13326 18368 13806
rect 18420 13388 18472 13394
rect 18420 13330 18472 13336
rect 18156 13246 18276 13274
rect 18328 13320 18380 13326
rect 18328 13262 18380 13268
rect 18052 12300 18104 12306
rect 18052 12242 18104 12248
rect 18052 11688 18104 11694
rect 18052 11630 18104 11636
rect 17960 11280 18012 11286
rect 17960 11222 18012 11228
rect 18064 11218 18092 11630
rect 18052 11212 18104 11218
rect 18052 11154 18104 11160
rect 17592 10124 17644 10130
rect 17592 10066 17644 10072
rect 17500 9580 17552 9586
rect 17500 9522 17552 9528
rect 17040 9376 17092 9382
rect 17040 9318 17092 9324
rect 17960 9376 18012 9382
rect 17960 9318 18012 9324
rect 17052 9178 17080 9318
rect 17040 9172 17092 9178
rect 17040 9114 17092 9120
rect 16762 9072 16818 9081
rect 16580 9036 16632 9042
rect 17052 9042 17080 9114
rect 16762 9007 16818 9016
rect 17040 9036 17092 9042
rect 16580 8978 16632 8984
rect 16120 8628 16172 8634
rect 16120 8570 16172 8576
rect 16212 8424 16264 8430
rect 16210 8392 16212 8401
rect 16580 8424 16632 8430
rect 16264 8392 16266 8401
rect 16210 8327 16266 8336
rect 16500 8384 16580 8412
rect 16500 8294 16528 8384
rect 16580 8366 16632 8372
rect 16488 8288 16540 8294
rect 16488 8230 16540 8236
rect 16028 8084 16080 8090
rect 16028 8026 16080 8032
rect 16040 7954 16068 8026
rect 16776 7954 16804 9007
rect 17040 8978 17092 8984
rect 17316 8424 17368 8430
rect 17314 8392 17316 8401
rect 17368 8392 17370 8401
rect 17314 8327 17370 8336
rect 16948 8288 17000 8294
rect 16854 8256 16910 8265
rect 16948 8230 17000 8236
rect 16854 8191 16910 8200
rect 16028 7948 16080 7954
rect 16028 7890 16080 7896
rect 16580 7948 16632 7954
rect 16580 7890 16632 7896
rect 16764 7948 16816 7954
rect 16764 7890 16816 7896
rect 15936 7540 15988 7546
rect 15936 7482 15988 7488
rect 15948 7002 15976 7482
rect 16488 7404 16540 7410
rect 16488 7346 16540 7352
rect 16500 7206 16528 7346
rect 16488 7200 16540 7206
rect 16488 7142 16540 7148
rect 15936 6996 15988 7002
rect 15936 6938 15988 6944
rect 15844 6860 15896 6866
rect 15844 6802 15896 6808
rect 16120 6724 16172 6730
rect 16120 6666 16172 6672
rect 16132 6322 16160 6666
rect 16120 6316 16172 6322
rect 16120 6258 16172 6264
rect 15672 5868 15976 5896
rect 15568 5840 15620 5846
rect 15568 5782 15620 5788
rect 15580 5574 15608 5782
rect 15672 5778 15700 5868
rect 15660 5772 15712 5778
rect 15660 5714 15712 5720
rect 15844 5772 15896 5778
rect 15844 5714 15896 5720
rect 15568 5568 15620 5574
rect 15568 5510 15620 5516
rect 15580 5166 15608 5510
rect 15568 5160 15620 5166
rect 15568 5102 15620 5108
rect 15752 4684 15804 4690
rect 15752 4626 15804 4632
rect 15016 4140 15068 4146
rect 15016 4082 15068 4088
rect 15476 4140 15528 4146
rect 15476 4082 15528 4088
rect 14004 4072 14056 4078
rect 14004 4014 14056 4020
rect 14740 4072 14792 4078
rect 14740 4014 14792 4020
rect 13452 3732 13504 3738
rect 13452 3674 13504 3680
rect 12808 3596 12860 3602
rect 12808 3538 12860 3544
rect 14016 3194 14044 4014
rect 14188 4004 14240 4010
rect 14188 3946 14240 3952
rect 14004 3188 14056 3194
rect 14004 3130 14056 3136
rect 12900 2576 12952 2582
rect 12900 2518 12952 2524
rect 12624 2440 12676 2446
rect 12624 2382 12676 2388
rect 12912 800 12940 2518
rect 14200 2446 14228 3946
rect 14752 3534 14780 4014
rect 14832 3732 14884 3738
rect 14832 3674 14884 3680
rect 14740 3528 14792 3534
rect 14740 3470 14792 3476
rect 14464 3392 14516 3398
rect 14464 3334 14516 3340
rect 14476 2514 14504 3334
rect 14844 3058 14872 3674
rect 15292 3596 15344 3602
rect 15292 3538 15344 3544
rect 14924 3392 14976 3398
rect 14924 3334 14976 3340
rect 14832 3052 14884 3058
rect 14832 2994 14884 3000
rect 14464 2508 14516 2514
rect 14464 2450 14516 2456
rect 14188 2440 14240 2446
rect 14188 2382 14240 2388
rect 14936 800 14964 3334
rect 15304 3058 15332 3538
rect 15292 3052 15344 3058
rect 15292 2994 15344 3000
rect 15488 2514 15516 4082
rect 15568 3596 15620 3602
rect 15568 3538 15620 3544
rect 15476 2508 15528 2514
rect 15476 2450 15528 2456
rect 15580 2378 15608 3538
rect 15764 3194 15792 4626
rect 15856 3602 15884 5714
rect 15948 5098 15976 5868
rect 16592 5710 16620 7890
rect 16868 7750 16896 8191
rect 16960 7886 16988 8230
rect 16948 7880 17000 7886
rect 16948 7822 17000 7828
rect 16856 7744 16908 7750
rect 16856 7686 16908 7692
rect 16868 6866 16896 7686
rect 16856 6860 16908 6866
rect 16856 6802 16908 6808
rect 16672 5908 16724 5914
rect 16672 5850 16724 5856
rect 16684 5778 16712 5850
rect 16672 5772 16724 5778
rect 16672 5714 16724 5720
rect 16580 5704 16632 5710
rect 16580 5646 16632 5652
rect 16684 5370 16712 5714
rect 16672 5364 16724 5370
rect 16672 5306 16724 5312
rect 16960 5166 16988 7822
rect 17328 7546 17356 8327
rect 17500 8288 17552 8294
rect 17500 8230 17552 8236
rect 17512 7954 17540 8230
rect 17500 7948 17552 7954
rect 17500 7890 17552 7896
rect 17684 7948 17736 7954
rect 17684 7890 17736 7896
rect 17498 7712 17554 7721
rect 17498 7647 17554 7656
rect 17316 7540 17368 7546
rect 17316 7482 17368 7488
rect 17512 6866 17540 7647
rect 17316 6860 17368 6866
rect 17316 6802 17368 6808
rect 17500 6860 17552 6866
rect 17500 6802 17552 6808
rect 17328 6118 17356 6802
rect 17316 6112 17368 6118
rect 17316 6054 17368 6060
rect 16488 5160 16540 5166
rect 16488 5102 16540 5108
rect 16948 5160 17000 5166
rect 16948 5102 17000 5108
rect 15936 5092 15988 5098
rect 15936 5034 15988 5040
rect 15948 4690 15976 5034
rect 15936 4684 15988 4690
rect 15936 4626 15988 4632
rect 15936 4480 15988 4486
rect 15936 4422 15988 4428
rect 15844 3596 15896 3602
rect 15844 3538 15896 3544
rect 15752 3188 15804 3194
rect 15752 3130 15804 3136
rect 15660 2916 15712 2922
rect 15660 2858 15712 2864
rect 15672 2514 15700 2858
rect 15948 2514 15976 4422
rect 16028 3936 16080 3942
rect 16028 3878 16080 3884
rect 16040 3738 16068 3878
rect 16028 3732 16080 3738
rect 16028 3674 16080 3680
rect 16500 3058 16528 5102
rect 16948 4684 17000 4690
rect 16948 4626 17000 4632
rect 16856 4548 16908 4554
rect 16856 4490 16908 4496
rect 16868 3602 16896 4490
rect 16960 4078 16988 4626
rect 16948 4072 17000 4078
rect 16948 4014 17000 4020
rect 17040 4072 17092 4078
rect 17040 4014 17092 4020
rect 16960 3602 16988 4014
rect 16856 3596 16908 3602
rect 16856 3538 16908 3544
rect 16948 3596 17000 3602
rect 16948 3538 17000 3544
rect 17052 3194 17080 4014
rect 17040 3188 17092 3194
rect 17040 3130 17092 3136
rect 16854 3088 16910 3097
rect 16488 3052 16540 3058
rect 16854 3023 16856 3032
rect 16488 2994 16540 3000
rect 16908 3023 16910 3032
rect 16856 2994 16908 3000
rect 17328 2990 17356 6054
rect 17696 5778 17724 7890
rect 17684 5772 17736 5778
rect 17684 5714 17736 5720
rect 17868 5704 17920 5710
rect 17868 5646 17920 5652
rect 17880 4690 17908 5646
rect 17972 5030 18000 9318
rect 17960 5024 18012 5030
rect 17960 4966 18012 4972
rect 17868 4684 17920 4690
rect 17868 4626 17920 4632
rect 17316 2984 17368 2990
rect 17316 2926 17368 2932
rect 15660 2508 15712 2514
rect 15660 2450 15712 2456
rect 15936 2508 15988 2514
rect 15936 2450 15988 2456
rect 15568 2372 15620 2378
rect 15568 2314 15620 2320
rect 17880 2310 17908 4626
rect 17972 3466 18000 4966
rect 18156 4554 18184 13246
rect 18432 12209 18460 13330
rect 18524 12782 18552 13874
rect 18512 12776 18564 12782
rect 18512 12718 18564 12724
rect 18616 12646 18644 17750
rect 18696 17740 18748 17746
rect 18696 17682 18748 17688
rect 18604 12640 18656 12646
rect 18604 12582 18656 12588
rect 18604 12300 18656 12306
rect 18524 12260 18604 12288
rect 18418 12200 18474 12209
rect 18418 12135 18474 12144
rect 18236 11348 18288 11354
rect 18236 11290 18288 11296
rect 18248 10198 18276 11290
rect 18420 11212 18472 11218
rect 18420 11154 18472 11160
rect 18328 11076 18380 11082
rect 18328 11018 18380 11024
rect 18340 10606 18368 11018
rect 18328 10600 18380 10606
rect 18328 10542 18380 10548
rect 18236 10192 18288 10198
rect 18236 10134 18288 10140
rect 18328 9376 18380 9382
rect 18328 9318 18380 9324
rect 18236 8356 18288 8362
rect 18236 8298 18288 8304
rect 18248 8022 18276 8298
rect 18236 8016 18288 8022
rect 18236 7958 18288 7964
rect 18340 7936 18368 9318
rect 18432 8974 18460 11154
rect 18420 8968 18472 8974
rect 18420 8910 18472 8916
rect 18420 7948 18472 7954
rect 18340 7908 18420 7936
rect 18420 7890 18472 7896
rect 18432 7818 18460 7890
rect 18420 7812 18472 7818
rect 18420 7754 18472 7760
rect 18432 7342 18460 7754
rect 18524 7698 18552 12260
rect 18604 12242 18656 12248
rect 18604 12164 18656 12170
rect 18604 12106 18656 12112
rect 18616 11898 18644 12106
rect 18604 11892 18656 11898
rect 18604 11834 18656 11840
rect 18616 11218 18644 11834
rect 18604 11212 18656 11218
rect 18604 11154 18656 11160
rect 18604 10600 18656 10606
rect 18604 10542 18656 10548
rect 18616 10198 18644 10542
rect 18604 10192 18656 10198
rect 18604 10134 18656 10140
rect 18604 9512 18656 9518
rect 18604 9454 18656 9460
rect 18616 8430 18644 9454
rect 18604 8424 18656 8430
rect 18604 8366 18656 8372
rect 18708 7834 18736 17682
rect 18788 16448 18840 16454
rect 18788 16390 18840 16396
rect 18800 11694 18828 16390
rect 18892 12306 18920 18770
rect 18984 18222 19012 19110
rect 19168 18748 19196 21558
rect 19260 20482 19288 21678
rect 19444 21593 19472 22510
rect 19580 22332 19876 22352
rect 19636 22330 19660 22332
rect 19716 22330 19740 22332
rect 19796 22330 19820 22332
rect 19658 22278 19660 22330
rect 19722 22278 19734 22330
rect 19796 22278 19798 22330
rect 19636 22276 19660 22278
rect 19716 22276 19740 22278
rect 19796 22276 19820 22278
rect 19580 22256 19876 22276
rect 19996 22166 20024 22510
rect 20088 22166 20116 23122
rect 19984 22160 20036 22166
rect 19984 22102 20036 22108
rect 20076 22160 20128 22166
rect 20076 22102 20128 22108
rect 19708 22092 19760 22098
rect 19760 22052 19840 22080
rect 19708 22034 19760 22040
rect 19430 21584 19486 21593
rect 19340 21548 19392 21554
rect 19430 21519 19486 21528
rect 19340 21490 19392 21496
rect 19352 20602 19380 21490
rect 19812 21486 19840 22052
rect 19892 21548 19944 21554
rect 19996 21536 20024 22102
rect 20074 21856 20130 21865
rect 20074 21791 20130 21800
rect 19944 21508 20024 21536
rect 19892 21490 19944 21496
rect 19800 21480 19852 21486
rect 19852 21428 19932 21434
rect 19800 21422 19932 21428
rect 19432 21412 19484 21418
rect 19812 21406 19932 21422
rect 19432 21354 19484 21360
rect 19444 20942 19472 21354
rect 19580 21244 19876 21264
rect 19636 21242 19660 21244
rect 19716 21242 19740 21244
rect 19796 21242 19820 21244
rect 19658 21190 19660 21242
rect 19722 21190 19734 21242
rect 19796 21190 19798 21242
rect 19636 21188 19660 21190
rect 19716 21188 19740 21190
rect 19796 21188 19820 21190
rect 19580 21168 19876 21188
rect 19904 21010 19932 21406
rect 19996 21078 20024 21508
rect 19984 21072 20036 21078
rect 19984 21014 20036 21020
rect 19892 21004 19944 21010
rect 19892 20946 19944 20952
rect 19432 20936 19484 20942
rect 19432 20878 19484 20884
rect 19340 20596 19392 20602
rect 19340 20538 19392 20544
rect 19260 20454 19472 20482
rect 19248 18760 19300 18766
rect 19168 18720 19248 18748
rect 19248 18702 19300 18708
rect 19064 18692 19116 18698
rect 19064 18634 19116 18640
rect 19076 18426 19104 18634
rect 19064 18420 19116 18426
rect 19064 18362 19116 18368
rect 18972 18216 19024 18222
rect 18972 18158 19024 18164
rect 19076 17678 19104 18362
rect 19064 17672 19116 17678
rect 19064 17614 19116 17620
rect 18972 17060 19024 17066
rect 19024 17020 19104 17048
rect 18972 17002 19024 17008
rect 19076 16522 19104 17020
rect 19064 16516 19116 16522
rect 19064 16458 19116 16464
rect 18972 16448 19024 16454
rect 18972 16390 19024 16396
rect 18984 15570 19012 16390
rect 19260 16250 19288 18702
rect 19340 17128 19392 17134
rect 19340 17070 19392 17076
rect 19248 16244 19300 16250
rect 19248 16186 19300 16192
rect 19064 16040 19116 16046
rect 19064 15982 19116 15988
rect 18972 15564 19024 15570
rect 18972 15506 19024 15512
rect 19076 15026 19104 15982
rect 19352 15706 19380 17070
rect 19444 16590 19472 20454
rect 19892 20392 19944 20398
rect 19892 20334 19944 20340
rect 19580 20156 19876 20176
rect 19636 20154 19660 20156
rect 19716 20154 19740 20156
rect 19796 20154 19820 20156
rect 19658 20102 19660 20154
rect 19722 20102 19734 20154
rect 19796 20102 19798 20154
rect 19636 20100 19660 20102
rect 19716 20100 19740 20102
rect 19796 20100 19820 20102
rect 19580 20080 19876 20100
rect 19580 19068 19876 19088
rect 19636 19066 19660 19068
rect 19716 19066 19740 19068
rect 19796 19066 19820 19068
rect 19658 19014 19660 19066
rect 19722 19014 19734 19066
rect 19796 19014 19798 19066
rect 19636 19012 19660 19014
rect 19716 19012 19740 19014
rect 19796 19012 19820 19014
rect 19580 18992 19876 19012
rect 19708 18828 19760 18834
rect 19708 18770 19760 18776
rect 19720 18426 19748 18770
rect 19904 18630 19932 20334
rect 20088 19786 20116 21791
rect 20180 21690 20208 26710
rect 20260 26580 20312 26586
rect 20260 26522 20312 26528
rect 20272 25838 20300 26522
rect 20260 25832 20312 25838
rect 20260 25774 20312 25780
rect 20456 25650 20484 26862
rect 20640 26450 20668 26862
rect 20996 26862 21048 26868
rect 21088 26920 21140 26926
rect 21088 26862 21140 26868
rect 20718 26823 20774 26832
rect 20628 26444 20680 26450
rect 20628 26386 20680 26392
rect 21008 26246 21036 26862
rect 21088 26444 21140 26450
rect 21088 26386 21140 26392
rect 21100 26314 21128 26386
rect 21088 26308 21140 26314
rect 21088 26250 21140 26256
rect 21272 26308 21324 26314
rect 21272 26250 21324 26256
rect 20996 26240 21048 26246
rect 20996 26182 21048 26188
rect 21284 25906 21312 26250
rect 21272 25900 21324 25906
rect 21272 25842 21324 25848
rect 20904 25832 20956 25838
rect 20904 25774 20956 25780
rect 20996 25832 21048 25838
rect 20996 25774 21048 25780
rect 20272 25622 20484 25650
rect 20272 24070 20300 25622
rect 20916 24274 20944 25774
rect 20904 24268 20956 24274
rect 20904 24210 20956 24216
rect 20260 24064 20312 24070
rect 20260 24006 20312 24012
rect 20168 21684 20220 21690
rect 20168 21626 20220 21632
rect 20272 21570 20300 24006
rect 20628 23656 20680 23662
rect 20628 23598 20680 23604
rect 20444 22500 20496 22506
rect 20444 22442 20496 22448
rect 20352 22432 20404 22438
rect 20352 22374 20404 22380
rect 20180 21542 20300 21570
rect 20076 19780 20128 19786
rect 20076 19722 20128 19728
rect 20076 19372 20128 19378
rect 20076 19314 20128 19320
rect 19984 18896 20036 18902
rect 19984 18838 20036 18844
rect 19892 18624 19944 18630
rect 19892 18566 19944 18572
rect 19708 18420 19760 18426
rect 19708 18362 19760 18368
rect 19996 18358 20024 18838
rect 19984 18352 20036 18358
rect 19984 18294 20036 18300
rect 19580 17980 19876 18000
rect 19636 17978 19660 17980
rect 19716 17978 19740 17980
rect 19796 17978 19820 17980
rect 19658 17926 19660 17978
rect 19722 17926 19734 17978
rect 19796 17926 19798 17978
rect 19636 17924 19660 17926
rect 19716 17924 19740 17926
rect 19796 17924 19820 17926
rect 19580 17904 19876 17924
rect 19996 17882 20024 18294
rect 19984 17876 20036 17882
rect 19984 17818 20036 17824
rect 19892 17536 19944 17542
rect 19892 17478 19944 17484
rect 19580 16892 19876 16912
rect 19636 16890 19660 16892
rect 19716 16890 19740 16892
rect 19796 16890 19820 16892
rect 19658 16838 19660 16890
rect 19722 16838 19734 16890
rect 19796 16838 19798 16890
rect 19636 16836 19660 16838
rect 19716 16836 19740 16838
rect 19796 16836 19820 16838
rect 19580 16816 19876 16836
rect 19432 16584 19484 16590
rect 19432 16526 19484 16532
rect 19580 15804 19876 15824
rect 19636 15802 19660 15804
rect 19716 15802 19740 15804
rect 19796 15802 19820 15804
rect 19658 15750 19660 15802
rect 19722 15750 19734 15802
rect 19796 15750 19798 15802
rect 19636 15748 19660 15750
rect 19716 15748 19740 15750
rect 19796 15748 19820 15750
rect 19580 15728 19876 15748
rect 19340 15700 19392 15706
rect 19340 15642 19392 15648
rect 19800 15632 19852 15638
rect 19904 15586 19932 17478
rect 19984 15904 20036 15910
rect 19984 15846 20036 15852
rect 19852 15580 19932 15586
rect 19800 15574 19932 15580
rect 19812 15558 19932 15574
rect 19064 15020 19116 15026
rect 19064 14962 19116 14968
rect 19064 14884 19116 14890
rect 19064 14826 19116 14832
rect 19248 14884 19300 14890
rect 19248 14826 19300 14832
rect 19076 14482 19104 14826
rect 19260 14618 19288 14826
rect 19432 14816 19484 14822
rect 19432 14758 19484 14764
rect 19248 14612 19300 14618
rect 19248 14554 19300 14560
rect 19340 14544 19392 14550
rect 19340 14486 19392 14492
rect 19064 14476 19116 14482
rect 19064 14418 19116 14424
rect 19156 14476 19208 14482
rect 19156 14418 19208 14424
rect 18972 14068 19024 14074
rect 18972 14010 19024 14016
rect 18984 13394 19012 14010
rect 19076 13530 19104 14418
rect 19168 13818 19196 14418
rect 19248 14408 19300 14414
rect 19248 14350 19300 14356
rect 19260 14006 19288 14350
rect 19248 14000 19300 14006
rect 19248 13942 19300 13948
rect 19168 13790 19288 13818
rect 19064 13524 19116 13530
rect 19064 13466 19116 13472
rect 19260 13462 19288 13790
rect 19248 13456 19300 13462
rect 19248 13398 19300 13404
rect 18972 13388 19024 13394
rect 18972 13330 19024 13336
rect 18984 13138 19012 13330
rect 18984 13110 19196 13138
rect 18972 12436 19024 12442
rect 18972 12378 19024 12384
rect 18880 12300 18932 12306
rect 18880 12242 18932 12248
rect 18788 11688 18840 11694
rect 18786 11656 18788 11665
rect 18840 11656 18842 11665
rect 18786 11591 18842 11600
rect 18984 11150 19012 12378
rect 19064 12232 19116 12238
rect 19064 12174 19116 12180
rect 19076 11898 19104 12174
rect 19064 11892 19116 11898
rect 19064 11834 19116 11840
rect 18972 11144 19024 11150
rect 18972 11086 19024 11092
rect 18984 9518 19012 11086
rect 19076 10198 19104 11834
rect 19168 11218 19196 13110
rect 19156 11212 19208 11218
rect 19156 11154 19208 11160
rect 19064 10192 19116 10198
rect 19064 10134 19116 10140
rect 19076 10062 19104 10134
rect 19156 10124 19208 10130
rect 19156 10066 19208 10072
rect 19064 10056 19116 10062
rect 19064 9998 19116 10004
rect 18972 9512 19024 9518
rect 18972 9454 19024 9460
rect 18880 9376 18932 9382
rect 18880 9318 18932 9324
rect 18892 7954 18920 9318
rect 18970 9208 19026 9217
rect 18970 9143 19026 9152
rect 18984 8566 19012 9143
rect 19064 9036 19116 9042
rect 19064 8978 19116 8984
rect 18972 8560 19024 8566
rect 18972 8502 19024 8508
rect 19076 8498 19104 8978
rect 19064 8492 19116 8498
rect 19064 8434 19116 8440
rect 18972 8424 19024 8430
rect 18972 8366 19024 8372
rect 18984 8265 19012 8366
rect 19064 8356 19116 8362
rect 19064 8298 19116 8304
rect 18970 8256 19026 8265
rect 18970 8191 19026 8200
rect 19076 7954 19104 8298
rect 18880 7948 18932 7954
rect 18880 7890 18932 7896
rect 19064 7948 19116 7954
rect 19064 7890 19116 7896
rect 18708 7806 19104 7834
rect 18524 7670 18736 7698
rect 18420 7336 18472 7342
rect 18420 7278 18472 7284
rect 18236 6792 18288 6798
rect 18236 6734 18288 6740
rect 18248 4690 18276 6734
rect 18512 5772 18564 5778
rect 18512 5714 18564 5720
rect 18328 5092 18380 5098
rect 18328 5034 18380 5040
rect 18236 4684 18288 4690
rect 18236 4626 18288 4632
rect 18144 4548 18196 4554
rect 18144 4490 18196 4496
rect 18052 4072 18104 4078
rect 18052 4014 18104 4020
rect 18064 3466 18092 4014
rect 17960 3460 18012 3466
rect 17960 3402 18012 3408
rect 18052 3460 18104 3466
rect 18052 3402 18104 3408
rect 18340 2990 18368 5034
rect 18524 4690 18552 5714
rect 18604 5160 18656 5166
rect 18604 5102 18656 5108
rect 18616 4826 18644 5102
rect 18604 4820 18656 4826
rect 18604 4762 18656 4768
rect 18512 4684 18564 4690
rect 18512 4626 18564 4632
rect 18616 4622 18644 4762
rect 18604 4616 18656 4622
rect 18604 4558 18656 4564
rect 18328 2984 18380 2990
rect 18328 2926 18380 2932
rect 17960 2916 18012 2922
rect 17960 2858 18012 2864
rect 17972 2582 18000 2858
rect 18708 2854 18736 7670
rect 18972 4548 19024 4554
rect 18972 4490 19024 4496
rect 18696 2848 18748 2854
rect 18696 2790 18748 2796
rect 17960 2576 18012 2582
rect 17960 2518 18012 2524
rect 18880 2440 18932 2446
rect 18880 2382 18932 2388
rect 16948 2304 17000 2310
rect 16948 2246 17000 2252
rect 17868 2304 17920 2310
rect 17868 2246 17920 2252
rect 16960 800 16988 2246
rect 18892 2038 18920 2382
rect 18880 2032 18932 2038
rect 18880 1974 18932 1980
rect 18984 800 19012 4490
rect 19076 4010 19104 7806
rect 19168 7410 19196 10066
rect 19260 10062 19288 13398
rect 19352 12782 19380 14486
rect 19444 13394 19472 14758
rect 19580 14716 19876 14736
rect 19636 14714 19660 14716
rect 19716 14714 19740 14716
rect 19796 14714 19820 14716
rect 19658 14662 19660 14714
rect 19722 14662 19734 14714
rect 19796 14662 19798 14714
rect 19636 14660 19660 14662
rect 19716 14660 19740 14662
rect 19796 14660 19820 14662
rect 19580 14640 19876 14660
rect 19890 14512 19946 14521
rect 19800 14476 19852 14482
rect 19890 14447 19892 14456
rect 19800 14418 19852 14424
rect 19944 14447 19946 14456
rect 19892 14418 19944 14424
rect 19812 13716 19840 14418
rect 19812 13688 19932 13716
rect 19580 13628 19876 13648
rect 19636 13626 19660 13628
rect 19716 13626 19740 13628
rect 19796 13626 19820 13628
rect 19658 13574 19660 13626
rect 19722 13574 19734 13626
rect 19796 13574 19798 13626
rect 19636 13572 19660 13574
rect 19716 13572 19740 13574
rect 19796 13572 19820 13574
rect 19580 13552 19876 13572
rect 19432 13388 19484 13394
rect 19432 13330 19484 13336
rect 19904 13190 19932 13688
rect 19996 13546 20024 15846
rect 20088 13734 20116 19314
rect 20180 17542 20208 21542
rect 20260 21480 20312 21486
rect 20260 21422 20312 21428
rect 20272 20058 20300 21422
rect 20364 21078 20392 22374
rect 20352 21072 20404 21078
rect 20352 21014 20404 21020
rect 20456 20874 20484 22442
rect 20536 21344 20588 21350
rect 20536 21286 20588 21292
rect 20548 20942 20576 21286
rect 20536 20936 20588 20942
rect 20536 20878 20588 20884
rect 20444 20868 20496 20874
rect 20444 20810 20496 20816
rect 20456 20398 20484 20810
rect 20548 20398 20576 20878
rect 20444 20392 20496 20398
rect 20444 20334 20496 20340
rect 20536 20392 20588 20398
rect 20536 20334 20588 20340
rect 20260 20052 20312 20058
rect 20260 19994 20312 20000
rect 20168 17536 20220 17542
rect 20168 17478 20220 17484
rect 20168 16992 20220 16998
rect 20168 16934 20220 16940
rect 20180 13870 20208 16934
rect 20168 13864 20220 13870
rect 20168 13806 20220 13812
rect 20272 13818 20300 19994
rect 20536 19304 20588 19310
rect 20536 19246 20588 19252
rect 20350 18728 20406 18737
rect 20350 18663 20352 18672
rect 20404 18663 20406 18672
rect 20352 18634 20404 18640
rect 20548 18086 20576 19246
rect 20536 18080 20588 18086
rect 20536 18022 20588 18028
rect 20444 17740 20496 17746
rect 20444 17682 20496 17688
rect 20352 17536 20404 17542
rect 20352 17478 20404 17484
rect 20364 14958 20392 17478
rect 20456 17270 20484 17682
rect 20444 17264 20496 17270
rect 20444 17206 20496 17212
rect 20548 16998 20576 18022
rect 20536 16992 20588 16998
rect 20536 16934 20588 16940
rect 20352 14952 20404 14958
rect 20352 14894 20404 14900
rect 20444 14408 20496 14414
rect 20444 14350 20496 14356
rect 20456 13938 20484 14350
rect 20444 13932 20496 13938
rect 20444 13874 20496 13880
rect 20076 13728 20128 13734
rect 20180 13716 20208 13806
rect 20272 13790 20484 13818
rect 20180 13688 20300 13716
rect 20076 13670 20128 13676
rect 19996 13518 20208 13546
rect 19984 13388 20036 13394
rect 19984 13330 20036 13336
rect 19892 13184 19944 13190
rect 19892 13126 19944 13132
rect 19892 12844 19944 12850
rect 19892 12786 19944 12792
rect 19340 12776 19392 12782
rect 19340 12718 19392 12724
rect 19432 12708 19484 12714
rect 19432 12650 19484 12656
rect 19444 12374 19472 12650
rect 19580 12540 19876 12560
rect 19636 12538 19660 12540
rect 19716 12538 19740 12540
rect 19796 12538 19820 12540
rect 19658 12486 19660 12538
rect 19722 12486 19734 12538
rect 19796 12486 19798 12538
rect 19636 12484 19660 12486
rect 19716 12484 19740 12486
rect 19796 12484 19820 12486
rect 19580 12464 19876 12484
rect 19432 12368 19484 12374
rect 19432 12310 19484 12316
rect 19340 12300 19392 12306
rect 19340 12242 19392 12248
rect 19708 12300 19760 12306
rect 19708 12242 19760 12248
rect 19352 10470 19380 12242
rect 19720 11898 19748 12242
rect 19708 11892 19760 11898
rect 19708 11834 19760 11840
rect 19904 11762 19932 12786
rect 19996 12782 20024 13330
rect 19984 12776 20036 12782
rect 19984 12718 20036 12724
rect 19892 11756 19944 11762
rect 19892 11698 19944 11704
rect 19432 11552 19484 11558
rect 19432 11494 19484 11500
rect 20076 11552 20128 11558
rect 20076 11494 20128 11500
rect 19444 11218 19472 11494
rect 19580 11452 19876 11472
rect 19636 11450 19660 11452
rect 19716 11450 19740 11452
rect 19796 11450 19820 11452
rect 19658 11398 19660 11450
rect 19722 11398 19734 11450
rect 19796 11398 19798 11450
rect 19636 11396 19660 11398
rect 19716 11396 19740 11398
rect 19796 11396 19820 11398
rect 19580 11376 19876 11396
rect 20088 11286 20116 11494
rect 20076 11280 20128 11286
rect 20076 11222 20128 11228
rect 19432 11212 19484 11218
rect 19432 11154 19484 11160
rect 19444 10606 19472 11154
rect 19432 10600 19484 10606
rect 19432 10542 19484 10548
rect 19340 10464 19392 10470
rect 19340 10406 19392 10412
rect 19444 10130 19472 10542
rect 19580 10364 19876 10384
rect 19636 10362 19660 10364
rect 19716 10362 19740 10364
rect 19796 10362 19820 10364
rect 19658 10310 19660 10362
rect 19722 10310 19734 10362
rect 19796 10310 19798 10362
rect 19636 10308 19660 10310
rect 19716 10308 19740 10310
rect 19796 10308 19820 10310
rect 19580 10288 19876 10308
rect 19340 10124 19392 10130
rect 19340 10066 19392 10072
rect 19432 10124 19484 10130
rect 19432 10066 19484 10072
rect 20076 10124 20128 10130
rect 20076 10066 20128 10072
rect 19248 10056 19300 10062
rect 19248 9998 19300 10004
rect 19248 9920 19300 9926
rect 19248 9862 19300 9868
rect 19260 8974 19288 9862
rect 19248 8968 19300 8974
rect 19248 8910 19300 8916
rect 19260 8362 19288 8910
rect 19248 8356 19300 8362
rect 19248 8298 19300 8304
rect 19156 7404 19208 7410
rect 19156 7346 19208 7352
rect 19352 7342 19380 10066
rect 19892 9580 19944 9586
rect 19892 9522 19944 9528
rect 19432 9444 19484 9450
rect 19432 9386 19484 9392
rect 19444 9081 19472 9386
rect 19580 9276 19876 9296
rect 19636 9274 19660 9276
rect 19716 9274 19740 9276
rect 19796 9274 19820 9276
rect 19658 9222 19660 9274
rect 19722 9222 19734 9274
rect 19796 9222 19798 9274
rect 19636 9220 19660 9222
rect 19716 9220 19740 9222
rect 19796 9220 19820 9222
rect 19580 9200 19876 9220
rect 19430 9072 19486 9081
rect 19430 9007 19486 9016
rect 19904 8906 19932 9522
rect 19984 9512 20036 9518
rect 19984 9454 20036 9460
rect 19996 9178 20024 9454
rect 19984 9172 20036 9178
rect 19984 9114 20036 9120
rect 19892 8900 19944 8906
rect 19892 8842 19944 8848
rect 19580 8188 19876 8208
rect 19636 8186 19660 8188
rect 19716 8186 19740 8188
rect 19796 8186 19820 8188
rect 19658 8134 19660 8186
rect 19722 8134 19734 8186
rect 19796 8134 19798 8186
rect 19636 8132 19660 8134
rect 19716 8132 19740 8134
rect 19796 8132 19820 8134
rect 19580 8112 19876 8132
rect 19432 7948 19484 7954
rect 19432 7890 19484 7896
rect 19892 7948 19944 7954
rect 19892 7890 19944 7896
rect 19340 7336 19392 7342
rect 19340 7278 19392 7284
rect 19156 6248 19208 6254
rect 19156 6190 19208 6196
rect 19168 5710 19196 6190
rect 19340 5772 19392 5778
rect 19340 5714 19392 5720
rect 19156 5704 19208 5710
rect 19156 5646 19208 5652
rect 19352 5234 19380 5714
rect 19340 5228 19392 5234
rect 19340 5170 19392 5176
rect 19444 5166 19472 7890
rect 19904 7818 19932 7890
rect 19892 7812 19944 7818
rect 19892 7754 19944 7760
rect 19892 7404 19944 7410
rect 19892 7346 19944 7352
rect 19580 7100 19876 7120
rect 19636 7098 19660 7100
rect 19716 7098 19740 7100
rect 19796 7098 19820 7100
rect 19658 7046 19660 7098
rect 19722 7046 19734 7098
rect 19796 7046 19798 7098
rect 19636 7044 19660 7046
rect 19716 7044 19740 7046
rect 19796 7044 19820 7046
rect 19580 7024 19876 7044
rect 19580 6012 19876 6032
rect 19636 6010 19660 6012
rect 19716 6010 19740 6012
rect 19796 6010 19820 6012
rect 19658 5958 19660 6010
rect 19722 5958 19734 6010
rect 19796 5958 19798 6010
rect 19636 5956 19660 5958
rect 19716 5956 19740 5958
rect 19796 5956 19820 5958
rect 19580 5936 19876 5956
rect 19904 5778 19932 7346
rect 19996 6934 20024 9114
rect 19984 6928 20036 6934
rect 19984 6870 20036 6876
rect 19984 5840 20036 5846
rect 19984 5782 20036 5788
rect 19892 5772 19944 5778
rect 19892 5714 19944 5720
rect 19892 5636 19944 5642
rect 19892 5578 19944 5584
rect 19432 5160 19484 5166
rect 19432 5102 19484 5108
rect 19340 4480 19392 4486
rect 19340 4422 19392 4428
rect 19352 4214 19380 4422
rect 19444 4282 19472 5102
rect 19580 4924 19876 4944
rect 19636 4922 19660 4924
rect 19716 4922 19740 4924
rect 19796 4922 19820 4924
rect 19658 4870 19660 4922
rect 19722 4870 19734 4922
rect 19796 4870 19798 4922
rect 19636 4868 19660 4870
rect 19716 4868 19740 4870
rect 19796 4868 19820 4870
rect 19580 4848 19876 4868
rect 19904 4554 19932 5578
rect 19996 4622 20024 5782
rect 20088 4672 20116 10066
rect 20180 9654 20208 13518
rect 20272 12714 20300 13688
rect 20352 12776 20404 12782
rect 20352 12718 20404 12724
rect 20260 12708 20312 12714
rect 20260 12650 20312 12656
rect 20272 11694 20300 12650
rect 20260 11688 20312 11694
rect 20260 11630 20312 11636
rect 20260 9988 20312 9994
rect 20260 9930 20312 9936
rect 20168 9648 20220 9654
rect 20168 9590 20220 9596
rect 20168 9512 20220 9518
rect 20168 9454 20220 9460
rect 20180 8838 20208 9454
rect 20272 8974 20300 9930
rect 20260 8968 20312 8974
rect 20260 8910 20312 8916
rect 20168 8832 20220 8838
rect 20168 8774 20220 8780
rect 20272 8616 20300 8910
rect 20364 8906 20392 12718
rect 20352 8900 20404 8906
rect 20352 8842 20404 8848
rect 20180 8588 20300 8616
rect 20180 8537 20208 8588
rect 20166 8528 20222 8537
rect 20166 8463 20222 8472
rect 20180 8090 20208 8463
rect 20260 8424 20312 8430
rect 20260 8366 20312 8372
rect 20168 8084 20220 8090
rect 20168 8026 20220 8032
rect 20180 7954 20208 8026
rect 20168 7948 20220 7954
rect 20168 7890 20220 7896
rect 20168 7268 20220 7274
rect 20168 7210 20220 7216
rect 20180 6390 20208 7210
rect 20272 7002 20300 8366
rect 20260 6996 20312 7002
rect 20260 6938 20312 6944
rect 20364 6848 20392 8842
rect 20272 6820 20392 6848
rect 20168 6384 20220 6390
rect 20168 6326 20220 6332
rect 20272 5642 20300 6820
rect 20456 6746 20484 13790
rect 20536 13184 20588 13190
rect 20536 13126 20588 13132
rect 20548 12782 20576 13126
rect 20536 12776 20588 12782
rect 20536 12718 20588 12724
rect 20640 10130 20668 23598
rect 20812 23248 20864 23254
rect 20812 23190 20864 23196
rect 20720 22500 20772 22506
rect 20720 22442 20772 22448
rect 20732 21010 20760 22442
rect 20720 21004 20772 21010
rect 20720 20946 20772 20952
rect 20824 20602 20852 23190
rect 21008 21865 21036 25774
rect 21272 25356 21324 25362
rect 21272 25298 21324 25304
rect 21088 24812 21140 24818
rect 21088 24754 21140 24760
rect 21100 24274 21128 24754
rect 21284 24750 21312 25298
rect 21272 24744 21324 24750
rect 21272 24686 21324 24692
rect 21088 24268 21140 24274
rect 21088 24210 21140 24216
rect 21376 23798 21404 34478
rect 21744 34134 21772 34478
rect 21732 34128 21784 34134
rect 21732 34070 21784 34076
rect 22388 33862 22416 34546
rect 21640 33856 21692 33862
rect 21640 33798 21692 33804
rect 22376 33856 22428 33862
rect 22376 33798 22428 33804
rect 21652 32978 21680 33798
rect 22376 33652 22428 33658
rect 22376 33594 22428 33600
rect 22388 32978 22416 33594
rect 23032 33522 23060 35702
rect 23388 35080 23440 35086
rect 23388 35022 23440 35028
rect 23400 34066 23428 35022
rect 23388 34060 23440 34066
rect 23388 34002 23440 34008
rect 23020 33516 23072 33522
rect 23020 33458 23072 33464
rect 23400 33454 23428 34002
rect 23768 33454 23796 39102
rect 23952 36802 23980 39200
rect 24952 37324 25004 37330
rect 24952 37266 25004 37272
rect 23860 36786 23980 36802
rect 23848 36780 23980 36786
rect 23900 36774 23980 36780
rect 23848 36722 23900 36728
rect 23940 36712 23992 36718
rect 23940 36654 23992 36660
rect 23952 36378 23980 36654
rect 23940 36372 23992 36378
rect 23940 36314 23992 36320
rect 24964 35834 24992 37266
rect 25044 36576 25096 36582
rect 25044 36518 25096 36524
rect 24952 35828 25004 35834
rect 24952 35770 25004 35776
rect 25056 35698 25084 36518
rect 25044 35692 25096 35698
rect 25044 35634 25096 35640
rect 24768 35148 24820 35154
rect 24768 35090 24820 35096
rect 24400 34944 24452 34950
rect 24400 34886 24452 34892
rect 24412 34610 24440 34886
rect 24400 34604 24452 34610
rect 24400 34546 24452 34552
rect 23848 34536 23900 34542
rect 23848 34478 23900 34484
rect 24216 34536 24268 34542
rect 24216 34478 24268 34484
rect 23860 33522 23888 34478
rect 24228 33998 24256 34478
rect 23940 33992 23992 33998
rect 23940 33934 23992 33940
rect 24216 33992 24268 33998
rect 24216 33934 24268 33940
rect 23952 33658 23980 33934
rect 24228 33862 24256 33934
rect 24216 33856 24268 33862
rect 24216 33798 24268 33804
rect 24676 33856 24728 33862
rect 24676 33798 24728 33804
rect 23940 33652 23992 33658
rect 23940 33594 23992 33600
rect 23848 33516 23900 33522
rect 23848 33458 23900 33464
rect 22652 33448 22704 33454
rect 22652 33390 22704 33396
rect 23388 33448 23440 33454
rect 23388 33390 23440 33396
rect 23756 33448 23808 33454
rect 23756 33390 23808 33396
rect 21640 32972 21692 32978
rect 21640 32914 21692 32920
rect 22376 32972 22428 32978
rect 22376 32914 22428 32920
rect 22192 32496 22244 32502
rect 22192 32438 22244 32444
rect 22008 32360 22060 32366
rect 22008 32302 22060 32308
rect 21824 32292 21876 32298
rect 21824 32234 21876 32240
rect 21836 31890 21864 32234
rect 22020 31958 22048 32302
rect 22008 31952 22060 31958
rect 22008 31894 22060 31900
rect 21824 31884 21876 31890
rect 21824 31826 21876 31832
rect 21836 31414 21864 31826
rect 21824 31408 21876 31414
rect 21824 31350 21876 31356
rect 21548 31272 21600 31278
rect 21548 31214 21600 31220
rect 21560 30326 21588 31214
rect 22008 30932 22060 30938
rect 22008 30874 22060 30880
rect 21548 30320 21600 30326
rect 21548 30262 21600 30268
rect 21560 28762 21588 30262
rect 21732 29300 21784 29306
rect 21732 29242 21784 29248
rect 21548 28756 21600 28762
rect 21548 28698 21600 28704
rect 21744 28694 21772 29242
rect 21732 28688 21784 28694
rect 21732 28630 21784 28636
rect 22020 28082 22048 30874
rect 22204 28626 22232 32438
rect 22376 32360 22428 32366
rect 22376 32302 22428 32308
rect 22388 31822 22416 32302
rect 22376 31816 22428 31822
rect 22376 31758 22428 31764
rect 22388 30938 22416 31758
rect 22664 31634 22692 33390
rect 23020 33380 23072 33386
rect 23020 33322 23072 33328
rect 22572 31606 22692 31634
rect 22376 30932 22428 30938
rect 22376 30874 22428 30880
rect 22284 30728 22336 30734
rect 22284 30670 22336 30676
rect 22296 28762 22324 30670
rect 22468 30184 22520 30190
rect 22468 30126 22520 30132
rect 22284 28756 22336 28762
rect 22284 28698 22336 28704
rect 22192 28620 22244 28626
rect 22192 28562 22244 28568
rect 22008 28076 22060 28082
rect 22008 28018 22060 28024
rect 21456 27940 21508 27946
rect 21456 27882 21508 27888
rect 21468 26450 21496 27882
rect 21548 27872 21600 27878
rect 21548 27814 21600 27820
rect 21560 26518 21588 27814
rect 22008 27532 22060 27538
rect 22008 27474 22060 27480
rect 22376 27532 22428 27538
rect 22376 27474 22428 27480
rect 22020 26790 22048 27474
rect 22284 27328 22336 27334
rect 22284 27270 22336 27276
rect 22100 26988 22152 26994
rect 22100 26930 22152 26936
rect 22112 26897 22140 26930
rect 22098 26888 22154 26897
rect 22098 26823 22154 26832
rect 22008 26784 22060 26790
rect 22008 26726 22060 26732
rect 21548 26512 21600 26518
rect 21548 26454 21600 26460
rect 21456 26444 21508 26450
rect 21456 26386 21508 26392
rect 21468 26042 21496 26386
rect 22020 26314 22048 26726
rect 22296 26450 22324 27270
rect 22388 26586 22416 27474
rect 22376 26580 22428 26586
rect 22376 26522 22428 26528
rect 22284 26444 22336 26450
rect 22284 26386 22336 26392
rect 22008 26308 22060 26314
rect 22008 26250 22060 26256
rect 22192 26240 22244 26246
rect 22192 26182 22244 26188
rect 21456 26036 21508 26042
rect 21456 25978 21508 25984
rect 22204 25906 22232 26182
rect 22192 25900 22244 25906
rect 22192 25842 22244 25848
rect 22296 25498 22324 26386
rect 22284 25492 22336 25498
rect 22284 25434 22336 25440
rect 22008 25356 22060 25362
rect 22008 25298 22060 25304
rect 21824 25220 21876 25226
rect 21824 25162 21876 25168
rect 21640 25152 21692 25158
rect 21640 25094 21692 25100
rect 21652 24750 21680 25094
rect 21836 24750 21864 25162
rect 22020 25158 22048 25298
rect 22008 25152 22060 25158
rect 22008 25094 22060 25100
rect 21640 24744 21692 24750
rect 21640 24686 21692 24692
rect 21824 24744 21876 24750
rect 21824 24686 21876 24692
rect 21732 24268 21784 24274
rect 21732 24210 21784 24216
rect 21364 23792 21416 23798
rect 21364 23734 21416 23740
rect 21744 23730 21772 24210
rect 21732 23724 21784 23730
rect 21732 23666 21784 23672
rect 21180 23656 21232 23662
rect 21180 23598 21232 23604
rect 21192 23186 21220 23598
rect 21548 23316 21600 23322
rect 21548 23258 21600 23264
rect 21180 23180 21232 23186
rect 21180 23122 21232 23128
rect 21560 22642 21588 23258
rect 21836 23118 21864 24686
rect 22020 24256 22048 25094
rect 22284 24948 22336 24954
rect 22284 24890 22336 24896
rect 22020 24228 22140 24256
rect 22008 23724 22060 23730
rect 22008 23666 22060 23672
rect 21916 23180 21968 23186
rect 21916 23122 21968 23128
rect 21640 23112 21692 23118
rect 21640 23054 21692 23060
rect 21824 23112 21876 23118
rect 21824 23054 21876 23060
rect 21548 22636 21600 22642
rect 21548 22578 21600 22584
rect 20994 21856 21050 21865
rect 20994 21791 21050 21800
rect 21652 21690 21680 23054
rect 21928 22710 21956 23122
rect 21916 22704 21968 22710
rect 21916 22646 21968 22652
rect 21916 22568 21968 22574
rect 21916 22510 21968 22516
rect 21732 22092 21784 22098
rect 21732 22034 21784 22040
rect 21824 22092 21876 22098
rect 21824 22034 21876 22040
rect 21744 21690 21772 22034
rect 21640 21684 21692 21690
rect 21640 21626 21692 21632
rect 21732 21684 21784 21690
rect 21732 21626 21784 21632
rect 21836 21486 21864 22034
rect 21180 21480 21232 21486
rect 21180 21422 21232 21428
rect 21824 21480 21876 21486
rect 21824 21422 21876 21428
rect 20812 20596 20864 20602
rect 20812 20538 20864 20544
rect 20904 20460 20956 20466
rect 20904 20402 20956 20408
rect 20720 19984 20772 19990
rect 20720 19926 20772 19932
rect 20732 18834 20760 19926
rect 20720 18828 20772 18834
rect 20720 18770 20772 18776
rect 20732 17882 20760 18770
rect 20812 18216 20864 18222
rect 20812 18158 20864 18164
rect 20720 17876 20772 17882
rect 20720 17818 20772 17824
rect 20720 16652 20772 16658
rect 20720 16594 20772 16600
rect 20732 16250 20760 16594
rect 20720 16244 20772 16250
rect 20720 16186 20772 16192
rect 20720 12640 20772 12646
rect 20720 12582 20772 12588
rect 20732 11082 20760 12582
rect 20720 11076 20772 11082
rect 20720 11018 20772 11024
rect 20824 10282 20852 18158
rect 20916 17542 20944 20402
rect 21192 19990 21220 21422
rect 21456 21140 21508 21146
rect 21456 21082 21508 21088
rect 21364 21072 21416 21078
rect 21364 21014 21416 21020
rect 21272 20528 21324 20534
rect 21272 20470 21324 20476
rect 21180 19984 21232 19990
rect 21180 19926 21232 19932
rect 21180 19712 21232 19718
rect 21180 19654 21232 19660
rect 21192 19378 21220 19654
rect 21180 19372 21232 19378
rect 21180 19314 21232 19320
rect 21284 19145 21312 20470
rect 21376 20466 21404 21014
rect 21364 20460 21416 20466
rect 21364 20402 21416 20408
rect 21468 20262 21496 21082
rect 21732 21004 21784 21010
rect 21732 20946 21784 20952
rect 21744 20534 21772 20946
rect 21548 20528 21600 20534
rect 21548 20470 21600 20476
rect 21732 20528 21784 20534
rect 21732 20470 21784 20476
rect 21456 20256 21508 20262
rect 21456 20198 21508 20204
rect 21468 19786 21496 20198
rect 21456 19780 21508 19786
rect 21456 19722 21508 19728
rect 21270 19136 21326 19145
rect 21270 19071 21326 19080
rect 20996 18896 21048 18902
rect 20996 18838 21048 18844
rect 21008 18290 21036 18838
rect 21560 18834 21588 20470
rect 21928 20074 21956 22510
rect 22020 20806 22048 23666
rect 22112 23662 22140 24228
rect 22100 23656 22152 23662
rect 22100 23598 22152 23604
rect 22100 22432 22152 22438
rect 22100 22374 22152 22380
rect 22008 20800 22060 20806
rect 22008 20742 22060 20748
rect 21744 20046 21956 20074
rect 21638 19680 21694 19689
rect 21638 19615 21694 19624
rect 21088 18828 21140 18834
rect 21088 18770 21140 18776
rect 21548 18828 21600 18834
rect 21548 18770 21600 18776
rect 20996 18284 21048 18290
rect 20996 18226 21048 18232
rect 21100 18086 21128 18770
rect 21088 18080 21140 18086
rect 21088 18022 21140 18028
rect 20904 17536 20956 17542
rect 20904 17478 20956 17484
rect 21100 17270 21128 18022
rect 21180 17604 21232 17610
rect 21180 17546 21232 17552
rect 21088 17264 21140 17270
rect 21088 17206 21140 17212
rect 21192 17134 21220 17546
rect 21272 17536 21324 17542
rect 21272 17478 21324 17484
rect 21180 17128 21232 17134
rect 21180 17070 21232 17076
rect 21192 16658 21220 17070
rect 21284 16794 21312 17478
rect 21272 16788 21324 16794
rect 21272 16730 21324 16736
rect 21088 16652 21140 16658
rect 21088 16594 21140 16600
rect 21180 16652 21232 16658
rect 21180 16594 21232 16600
rect 20904 16040 20956 16046
rect 20904 15982 20956 15988
rect 20916 15094 20944 15982
rect 20904 15088 20956 15094
rect 20904 15030 20956 15036
rect 20996 12776 21048 12782
rect 20996 12718 21048 12724
rect 20904 12232 20956 12238
rect 20904 12174 20956 12180
rect 20916 11694 20944 12174
rect 20904 11688 20956 11694
rect 20904 11630 20956 11636
rect 20732 10254 20852 10282
rect 20628 10124 20680 10130
rect 20628 10066 20680 10072
rect 20536 10056 20588 10062
rect 20536 9998 20588 10004
rect 20548 7342 20576 9998
rect 20628 9104 20680 9110
rect 20628 9046 20680 9052
rect 20640 7546 20668 9046
rect 20628 7540 20680 7546
rect 20628 7482 20680 7488
rect 20536 7336 20588 7342
rect 20536 7278 20588 7284
rect 20364 6718 20484 6746
rect 20260 5636 20312 5642
rect 20260 5578 20312 5584
rect 20272 5370 20300 5578
rect 20260 5364 20312 5370
rect 20260 5306 20312 5312
rect 20088 4644 20300 4672
rect 19984 4616 20036 4622
rect 19984 4558 20036 4564
rect 19892 4548 19944 4554
rect 19892 4490 19944 4496
rect 20076 4548 20128 4554
rect 20076 4490 20128 4496
rect 19432 4276 19484 4282
rect 19432 4218 19484 4224
rect 19340 4208 19392 4214
rect 19340 4150 19392 4156
rect 19064 4004 19116 4010
rect 19064 3946 19116 3952
rect 19248 3936 19300 3942
rect 19248 3878 19300 3884
rect 19260 2446 19288 3878
rect 19352 3670 19380 4150
rect 19432 3936 19484 3942
rect 19432 3878 19484 3884
rect 19340 3664 19392 3670
rect 19340 3606 19392 3612
rect 19444 3602 19472 3878
rect 19580 3836 19876 3856
rect 19636 3834 19660 3836
rect 19716 3834 19740 3836
rect 19796 3834 19820 3836
rect 19658 3782 19660 3834
rect 19722 3782 19734 3834
rect 19796 3782 19798 3834
rect 19636 3780 19660 3782
rect 19716 3780 19740 3782
rect 19796 3780 19820 3782
rect 19580 3760 19876 3780
rect 19432 3596 19484 3602
rect 19432 3538 19484 3544
rect 19904 3534 19932 4490
rect 20088 4146 20116 4490
rect 20076 4140 20128 4146
rect 20076 4082 20128 4088
rect 20168 4072 20220 4078
rect 20168 4014 20220 4020
rect 20076 4004 20128 4010
rect 20076 3946 20128 3952
rect 19892 3528 19944 3534
rect 19892 3470 19944 3476
rect 19580 2748 19876 2768
rect 19636 2746 19660 2748
rect 19716 2746 19740 2748
rect 19796 2746 19820 2748
rect 19658 2694 19660 2746
rect 19722 2694 19734 2746
rect 19796 2694 19798 2746
rect 19636 2692 19660 2694
rect 19716 2692 19740 2694
rect 19796 2692 19820 2694
rect 19580 2672 19876 2692
rect 19248 2440 19300 2446
rect 19248 2382 19300 2388
rect 20088 1970 20116 3946
rect 20180 3466 20208 4014
rect 20168 3460 20220 3466
rect 20168 3402 20220 3408
rect 20180 3194 20208 3402
rect 20272 3398 20300 4644
rect 20260 3392 20312 3398
rect 20260 3334 20312 3340
rect 20168 3188 20220 3194
rect 20168 3130 20220 3136
rect 20364 2310 20392 6718
rect 20548 6662 20576 7278
rect 20536 6656 20588 6662
rect 20536 6598 20588 6604
rect 20732 5846 20760 10254
rect 20812 10124 20864 10130
rect 20812 10066 20864 10072
rect 20824 9722 20852 10066
rect 20812 9716 20864 9722
rect 20812 9658 20864 9664
rect 20824 9042 20852 9658
rect 20904 9512 20956 9518
rect 20904 9454 20956 9460
rect 20812 9036 20864 9042
rect 20812 8978 20864 8984
rect 20916 8906 20944 9454
rect 20904 8900 20956 8906
rect 20904 8842 20956 8848
rect 20902 8528 20958 8537
rect 20902 8463 20904 8472
rect 20956 8463 20958 8472
rect 20904 8434 20956 8440
rect 20812 8424 20864 8430
rect 20812 8366 20864 8372
rect 20824 8022 20852 8366
rect 20904 8356 20956 8362
rect 20904 8298 20956 8304
rect 20916 8090 20944 8298
rect 20904 8084 20956 8090
rect 20904 8026 20956 8032
rect 20812 8016 20864 8022
rect 20812 7958 20864 7964
rect 20812 7268 20864 7274
rect 20812 7210 20864 7216
rect 20720 5840 20772 5846
rect 20720 5782 20772 5788
rect 20824 5234 20852 7210
rect 21008 5778 21036 12718
rect 21100 10146 21128 16594
rect 21192 15570 21220 16594
rect 21456 16040 21508 16046
rect 21454 16008 21456 16017
rect 21508 16008 21510 16017
rect 21454 15943 21510 15952
rect 21180 15564 21232 15570
rect 21180 15506 21232 15512
rect 21272 15088 21324 15094
rect 21272 15030 21324 15036
rect 21180 13320 21232 13326
rect 21180 13262 21232 13268
rect 21192 12306 21220 13262
rect 21180 12300 21232 12306
rect 21180 12242 21232 12248
rect 21284 11762 21312 15030
rect 21652 15026 21680 19615
rect 21744 19378 21772 20046
rect 21916 19916 21968 19922
rect 21916 19858 21968 19864
rect 21732 19372 21784 19378
rect 21732 19314 21784 19320
rect 21744 17610 21772 19314
rect 21928 18834 21956 19858
rect 22112 19689 22140 22374
rect 22192 22092 22244 22098
rect 22192 22034 22244 22040
rect 22204 21468 22232 22034
rect 22296 21622 22324 24890
rect 22480 24614 22508 30126
rect 22468 24608 22520 24614
rect 22468 24550 22520 24556
rect 22376 23792 22428 23798
rect 22376 23734 22428 23740
rect 22388 23254 22416 23734
rect 22376 23248 22428 23254
rect 22376 23190 22428 23196
rect 22376 22976 22428 22982
rect 22376 22918 22428 22924
rect 22388 22574 22416 22918
rect 22376 22568 22428 22574
rect 22376 22510 22428 22516
rect 22284 21616 22336 21622
rect 22284 21558 22336 21564
rect 22284 21480 22336 21486
rect 22204 21440 22284 21468
rect 22284 21422 22336 21428
rect 22296 20942 22324 21422
rect 22284 20936 22336 20942
rect 22284 20878 22336 20884
rect 22192 20324 22244 20330
rect 22192 20266 22244 20272
rect 22204 19922 22232 20266
rect 22296 20244 22324 20878
rect 22376 20256 22428 20262
rect 22296 20216 22376 20244
rect 22376 20198 22428 20204
rect 22192 19916 22244 19922
rect 22192 19858 22244 19864
rect 22098 19680 22154 19689
rect 22098 19615 22154 19624
rect 22204 19446 22232 19858
rect 22192 19440 22244 19446
rect 22192 19382 22244 19388
rect 22008 19304 22060 19310
rect 22060 19252 22140 19258
rect 22008 19246 22140 19252
rect 22020 19242 22140 19246
rect 22020 19236 22152 19242
rect 22020 19230 22100 19236
rect 22100 19178 22152 19184
rect 22006 19136 22062 19145
rect 22006 19071 22062 19080
rect 21916 18828 21968 18834
rect 21916 18770 21968 18776
rect 21732 17604 21784 17610
rect 21732 17546 21784 17552
rect 21824 17264 21876 17270
rect 21824 17206 21876 17212
rect 21836 16658 21864 17206
rect 22020 17134 22048 19071
rect 22204 18970 22232 19382
rect 22284 19168 22336 19174
rect 22284 19110 22336 19116
rect 22296 18970 22324 19110
rect 22192 18964 22244 18970
rect 22192 18906 22244 18912
rect 22284 18964 22336 18970
rect 22284 18906 22336 18912
rect 22100 18760 22152 18766
rect 22100 18702 22152 18708
rect 22112 18086 22140 18702
rect 22284 18216 22336 18222
rect 22284 18158 22336 18164
rect 22100 18080 22152 18086
rect 22100 18022 22152 18028
rect 22192 18080 22244 18086
rect 22192 18022 22244 18028
rect 22008 17128 22060 17134
rect 21928 17088 22008 17116
rect 21824 16652 21876 16658
rect 21744 16612 21824 16640
rect 21640 15020 21692 15026
rect 21640 14962 21692 14968
rect 21744 14958 21772 16612
rect 21824 16594 21876 16600
rect 21928 15570 21956 17088
rect 22008 17070 22060 17076
rect 22008 16720 22060 16726
rect 22008 16662 22060 16668
rect 21916 15564 21968 15570
rect 21916 15506 21968 15512
rect 21824 15496 21876 15502
rect 21824 15438 21876 15444
rect 21836 15094 21864 15438
rect 22020 15434 22048 16662
rect 22112 15978 22140 18022
rect 22204 17270 22232 18022
rect 22296 17746 22324 18158
rect 22284 17740 22336 17746
rect 22284 17682 22336 17688
rect 22192 17264 22244 17270
rect 22192 17206 22244 17212
rect 22192 16652 22244 16658
rect 22388 16640 22416 20198
rect 22468 18420 22520 18426
rect 22468 18362 22520 18368
rect 22480 18154 22508 18362
rect 22468 18148 22520 18154
rect 22468 18090 22520 18096
rect 22480 16658 22508 18090
rect 22244 16612 22416 16640
rect 22468 16652 22520 16658
rect 22192 16594 22244 16600
rect 22468 16594 22520 16600
rect 22204 16046 22232 16594
rect 22192 16040 22244 16046
rect 22192 15982 22244 15988
rect 22100 15972 22152 15978
rect 22100 15914 22152 15920
rect 22008 15428 22060 15434
rect 22008 15370 22060 15376
rect 21824 15088 21876 15094
rect 21824 15030 21876 15036
rect 21732 14952 21784 14958
rect 21732 14894 21784 14900
rect 21744 13734 21772 14894
rect 21836 14482 21864 15030
rect 21916 15020 21968 15026
rect 21916 14962 21968 14968
rect 21928 14550 21956 14962
rect 22112 14958 22140 15914
rect 22480 14958 22508 16594
rect 22100 14952 22152 14958
rect 22100 14894 22152 14900
rect 22468 14952 22520 14958
rect 22468 14894 22520 14900
rect 22008 14816 22060 14822
rect 22008 14758 22060 14764
rect 21916 14544 21968 14550
rect 21916 14486 21968 14492
rect 21824 14476 21876 14482
rect 21824 14418 21876 14424
rect 21824 14068 21876 14074
rect 21824 14010 21876 14016
rect 21732 13728 21784 13734
rect 21732 13670 21784 13676
rect 21744 13462 21772 13670
rect 21732 13456 21784 13462
rect 21732 13398 21784 13404
rect 21364 13320 21416 13326
rect 21364 13262 21416 13268
rect 21272 11756 21324 11762
rect 21272 11698 21324 11704
rect 21100 10118 21220 10146
rect 21088 9988 21140 9994
rect 21088 9930 21140 9936
rect 21100 9178 21128 9930
rect 21088 9172 21140 9178
rect 21088 9114 21140 9120
rect 21192 8430 21220 10118
rect 21272 10124 21324 10130
rect 21272 10066 21324 10072
rect 21284 9518 21312 10066
rect 21272 9512 21324 9518
rect 21272 9454 21324 9460
rect 21180 8424 21232 8430
rect 21180 8366 21232 8372
rect 21088 8288 21140 8294
rect 21088 8230 21140 8236
rect 21100 7750 21128 8230
rect 21088 7744 21140 7750
rect 21088 7686 21140 7692
rect 21284 7274 21312 9454
rect 21376 8566 21404 13262
rect 21456 11688 21508 11694
rect 21456 11630 21508 11636
rect 21468 11082 21496 11630
rect 21456 11076 21508 11082
rect 21456 11018 21508 11024
rect 21364 8560 21416 8566
rect 21364 8502 21416 8508
rect 21272 7268 21324 7274
rect 21272 7210 21324 7216
rect 21364 6248 21416 6254
rect 21364 6190 21416 6196
rect 20996 5772 21048 5778
rect 20996 5714 21048 5720
rect 21376 5642 21404 6190
rect 21364 5636 21416 5642
rect 21364 5578 21416 5584
rect 20812 5228 20864 5234
rect 20812 5170 20864 5176
rect 21272 5228 21324 5234
rect 21272 5170 21324 5176
rect 20628 5092 20680 5098
rect 20628 5034 20680 5040
rect 20720 5092 20772 5098
rect 20720 5034 20772 5040
rect 20444 4072 20496 4078
rect 20444 4014 20496 4020
rect 20456 3670 20484 4014
rect 20444 3664 20496 3670
rect 20444 3606 20496 3612
rect 20640 3074 20668 5034
rect 20732 4690 20760 5034
rect 20904 5024 20956 5030
rect 20904 4966 20956 4972
rect 20916 4690 20944 4966
rect 20720 4684 20772 4690
rect 20720 4626 20772 4632
rect 20904 4684 20956 4690
rect 20904 4626 20956 4632
rect 21284 3602 21312 5170
rect 21272 3596 21324 3602
rect 21272 3538 21324 3544
rect 20640 3046 20944 3074
rect 20916 2990 20944 3046
rect 20628 2984 20680 2990
rect 20628 2926 20680 2932
rect 20904 2984 20956 2990
rect 20904 2926 20956 2932
rect 20640 2446 20668 2926
rect 20628 2440 20680 2446
rect 20628 2382 20680 2388
rect 21364 2440 21416 2446
rect 21468 2428 21496 11018
rect 21836 10606 21864 14010
rect 21928 13394 21956 14486
rect 21916 13388 21968 13394
rect 21916 13330 21968 13336
rect 22020 12986 22048 14758
rect 22112 14482 22140 14894
rect 22192 14884 22244 14890
rect 22192 14826 22244 14832
rect 22204 14618 22232 14826
rect 22192 14612 22244 14618
rect 22192 14554 22244 14560
rect 22100 14476 22152 14482
rect 22100 14418 22152 14424
rect 22204 13394 22232 14554
rect 22284 14476 22336 14482
rect 22284 14418 22336 14424
rect 22192 13388 22244 13394
rect 22192 13330 22244 13336
rect 22296 12986 22324 14418
rect 22376 13932 22428 13938
rect 22376 13874 22428 13880
rect 22008 12980 22060 12986
rect 22008 12922 22060 12928
rect 22284 12980 22336 12986
rect 22284 12922 22336 12928
rect 22100 12096 22152 12102
rect 22100 12038 22152 12044
rect 22112 11694 22140 12038
rect 22100 11688 22152 11694
rect 22388 11642 22416 13874
rect 22572 13433 22600 31606
rect 23032 31482 23060 33322
rect 23400 33318 23428 33390
rect 23388 33312 23440 33318
rect 23388 33254 23440 33260
rect 23400 32434 23428 33254
rect 24228 32910 24256 33798
rect 24688 33454 24716 33798
rect 24676 33448 24728 33454
rect 24676 33390 24728 33396
rect 23848 32904 23900 32910
rect 23848 32846 23900 32852
rect 24216 32904 24268 32910
rect 24216 32846 24268 32852
rect 23756 32768 23808 32774
rect 23756 32710 23808 32716
rect 23388 32428 23440 32434
rect 23388 32370 23440 32376
rect 23400 32026 23428 32370
rect 23768 32366 23796 32710
rect 23756 32360 23808 32366
rect 23756 32302 23808 32308
rect 23388 32020 23440 32026
rect 23388 31962 23440 31968
rect 23860 31890 23888 32846
rect 24308 32768 24360 32774
rect 24308 32710 24360 32716
rect 24032 32292 24084 32298
rect 24032 32234 24084 32240
rect 24044 31890 24072 32234
rect 23204 31884 23256 31890
rect 23204 31826 23256 31832
rect 23848 31884 23900 31890
rect 23848 31826 23900 31832
rect 24032 31884 24084 31890
rect 24032 31826 24084 31832
rect 23020 31476 23072 31482
rect 23020 31418 23072 31424
rect 23216 31278 23244 31826
rect 24320 31278 24348 32710
rect 22836 31272 22888 31278
rect 22836 31214 22888 31220
rect 23204 31272 23256 31278
rect 23204 31214 23256 31220
rect 24308 31272 24360 31278
rect 24308 31214 24360 31220
rect 22652 30184 22704 30190
rect 22652 30126 22704 30132
rect 22664 29170 22692 30126
rect 22652 29164 22704 29170
rect 22652 29106 22704 29112
rect 22848 28098 22876 31214
rect 23572 30796 23624 30802
rect 23572 30738 23624 30744
rect 23480 30184 23532 30190
rect 23480 30126 23532 30132
rect 23204 29776 23256 29782
rect 23204 29718 23256 29724
rect 22928 29708 22980 29714
rect 22928 29650 22980 29656
rect 22940 29170 22968 29650
rect 22928 29164 22980 29170
rect 22928 29106 22980 29112
rect 23020 28620 23072 28626
rect 23020 28562 23072 28568
rect 23032 28218 23060 28562
rect 23020 28212 23072 28218
rect 23020 28154 23072 28160
rect 22848 28070 23060 28098
rect 22744 27940 22796 27946
rect 22744 27882 22796 27888
rect 22756 26790 22784 27882
rect 22836 27532 22888 27538
rect 22836 27474 22888 27480
rect 22744 26784 22796 26790
rect 22744 26726 22796 26732
rect 22756 26450 22784 26726
rect 22848 26518 22876 27474
rect 22928 27464 22980 27470
rect 22928 27406 22980 27412
rect 22940 27130 22968 27406
rect 22928 27124 22980 27130
rect 22928 27066 22980 27072
rect 22836 26512 22888 26518
rect 22834 26480 22836 26489
rect 22888 26480 22890 26489
rect 22744 26444 22796 26450
rect 22834 26415 22890 26424
rect 22744 26386 22796 26392
rect 22652 26308 22704 26314
rect 22652 26250 22704 26256
rect 22928 26308 22980 26314
rect 22928 26250 22980 26256
rect 22664 24750 22692 26250
rect 22744 25424 22796 25430
rect 22744 25366 22796 25372
rect 22756 24818 22784 25366
rect 22744 24812 22796 24818
rect 22744 24754 22796 24760
rect 22652 24744 22704 24750
rect 22652 24686 22704 24692
rect 22652 24268 22704 24274
rect 22652 24210 22704 24216
rect 22664 23594 22692 24210
rect 22744 23656 22796 23662
rect 22744 23598 22796 23604
rect 22652 23588 22704 23594
rect 22652 23530 22704 23536
rect 22664 22574 22692 23530
rect 22756 22778 22784 23598
rect 22744 22772 22796 22778
rect 22744 22714 22796 22720
rect 22652 22568 22704 22574
rect 22652 22510 22704 22516
rect 22744 22092 22796 22098
rect 22744 22034 22796 22040
rect 22756 21486 22784 22034
rect 22744 21480 22796 21486
rect 22744 21422 22796 21428
rect 22940 20602 22968 26250
rect 23032 25702 23060 28070
rect 23112 26580 23164 26586
rect 23112 26522 23164 26528
rect 23020 25696 23072 25702
rect 23020 25638 23072 25644
rect 23032 23866 23060 25638
rect 23124 25362 23152 26522
rect 23112 25356 23164 25362
rect 23112 25298 23164 25304
rect 23216 23866 23244 29718
rect 23296 29708 23348 29714
rect 23296 29650 23348 29656
rect 23308 29617 23336 29650
rect 23294 29608 23350 29617
rect 23294 29543 23350 29552
rect 23388 29028 23440 29034
rect 23388 28970 23440 28976
rect 23296 28008 23348 28014
rect 23296 27950 23348 27956
rect 23308 27146 23336 27950
rect 23400 27538 23428 28970
rect 23388 27532 23440 27538
rect 23388 27474 23440 27480
rect 23400 27334 23428 27474
rect 23492 27470 23520 30126
rect 23584 29714 23612 30738
rect 23848 30184 23900 30190
rect 23848 30126 23900 30132
rect 24216 30184 24268 30190
rect 24216 30126 24268 30132
rect 23572 29708 23624 29714
rect 23572 29650 23624 29656
rect 23860 29170 23888 30126
rect 24228 29782 24256 30126
rect 24216 29776 24268 29782
rect 24216 29718 24268 29724
rect 23848 29164 23900 29170
rect 23848 29106 23900 29112
rect 23664 28620 23716 28626
rect 23664 28562 23716 28568
rect 23572 28144 23624 28150
rect 23572 28086 23624 28092
rect 23480 27464 23532 27470
rect 23480 27406 23532 27412
rect 23388 27328 23440 27334
rect 23388 27270 23440 27276
rect 23308 27118 23428 27146
rect 23400 27062 23428 27118
rect 23388 27056 23440 27062
rect 23388 26998 23440 27004
rect 23400 26450 23428 26998
rect 23584 26926 23612 28086
rect 23572 26920 23624 26926
rect 23572 26862 23624 26868
rect 23584 26450 23612 26862
rect 23676 26858 23704 28562
rect 23848 27532 23900 27538
rect 23848 27474 23900 27480
rect 24124 27532 24176 27538
rect 24124 27474 24176 27480
rect 24216 27532 24268 27538
rect 24216 27474 24268 27480
rect 23860 26858 23888 27474
rect 24136 27062 24164 27474
rect 24124 27056 24176 27062
rect 24124 26998 24176 27004
rect 23664 26852 23716 26858
rect 23664 26794 23716 26800
rect 23848 26852 23900 26858
rect 23848 26794 23900 26800
rect 23388 26444 23440 26450
rect 23388 26386 23440 26392
rect 23572 26444 23624 26450
rect 23572 26386 23624 26392
rect 23020 23860 23072 23866
rect 23020 23802 23072 23808
rect 23204 23860 23256 23866
rect 23204 23802 23256 23808
rect 23400 22982 23428 26386
rect 23584 24614 23612 26386
rect 23664 26376 23716 26382
rect 23664 26318 23716 26324
rect 23676 25838 23704 26318
rect 23756 26036 23808 26042
rect 23756 25978 23808 25984
rect 23664 25832 23716 25838
rect 23664 25774 23716 25780
rect 23664 25288 23716 25294
rect 23664 25230 23716 25236
rect 23676 24886 23704 25230
rect 23664 24880 23716 24886
rect 23664 24822 23716 24828
rect 23676 24750 23704 24822
rect 23664 24744 23716 24750
rect 23664 24686 23716 24692
rect 23572 24608 23624 24614
rect 23572 24550 23624 24556
rect 23676 24274 23704 24686
rect 23664 24268 23716 24274
rect 23664 24210 23716 24216
rect 23388 22976 23440 22982
rect 23388 22918 23440 22924
rect 23400 22710 23428 22918
rect 23388 22704 23440 22710
rect 23388 22646 23440 22652
rect 23388 22568 23440 22574
rect 23388 22510 23440 22516
rect 23400 22234 23428 22510
rect 23112 22228 23164 22234
rect 23112 22170 23164 22176
rect 23388 22228 23440 22234
rect 23388 22170 23440 22176
rect 23020 20800 23072 20806
rect 23020 20742 23072 20748
rect 22928 20596 22980 20602
rect 22928 20538 22980 20544
rect 22744 20460 22796 20466
rect 22744 20402 22796 20408
rect 22756 18222 22784 20402
rect 22928 20256 22980 20262
rect 22928 20198 22980 20204
rect 22940 19786 22968 20198
rect 22928 19780 22980 19786
rect 22928 19722 22980 19728
rect 22836 19168 22888 19174
rect 22836 19110 22888 19116
rect 22744 18216 22796 18222
rect 22744 18158 22796 18164
rect 22652 18148 22704 18154
rect 22652 18090 22704 18096
rect 22664 17134 22692 18090
rect 22652 17128 22704 17134
rect 22652 17070 22704 17076
rect 22664 16114 22692 17070
rect 22652 16108 22704 16114
rect 22652 16050 22704 16056
rect 22848 15706 22876 19110
rect 23032 18222 23060 20742
rect 23124 19854 23152 22170
rect 23400 22098 23428 22170
rect 23388 22092 23440 22098
rect 23388 22034 23440 22040
rect 23572 21480 23624 21486
rect 23572 21422 23624 21428
rect 23480 20936 23532 20942
rect 23480 20878 23532 20884
rect 23112 19848 23164 19854
rect 23112 19790 23164 19796
rect 22928 18216 22980 18222
rect 22928 18158 22980 18164
rect 23020 18216 23072 18222
rect 23020 18158 23072 18164
rect 22940 17746 22968 18158
rect 23032 18086 23060 18158
rect 23020 18080 23072 18086
rect 23020 18022 23072 18028
rect 22928 17740 22980 17746
rect 22928 17682 22980 17688
rect 22940 15706 22968 17682
rect 23124 16266 23152 19790
rect 23296 19304 23348 19310
rect 23296 19246 23348 19252
rect 23308 18698 23336 19246
rect 23296 18692 23348 18698
rect 23296 18634 23348 18640
rect 23204 18624 23256 18630
rect 23204 18566 23256 18572
rect 23216 18426 23244 18566
rect 23204 18420 23256 18426
rect 23204 18362 23256 18368
rect 23204 18284 23256 18290
rect 23204 18226 23256 18232
rect 23216 17746 23244 18226
rect 23204 17740 23256 17746
rect 23204 17682 23256 17688
rect 23216 16658 23244 17682
rect 23308 17610 23336 18634
rect 23492 17814 23520 20878
rect 23584 20398 23612 21422
rect 23664 21344 23716 21350
rect 23664 21286 23716 21292
rect 23676 20942 23704 21286
rect 23664 20936 23716 20942
rect 23664 20878 23716 20884
rect 23676 20398 23704 20878
rect 23572 20392 23624 20398
rect 23572 20334 23624 20340
rect 23664 20392 23716 20398
rect 23664 20334 23716 20340
rect 23584 20058 23612 20334
rect 23572 20052 23624 20058
rect 23572 19994 23624 20000
rect 23664 18828 23716 18834
rect 23664 18770 23716 18776
rect 23572 18692 23624 18698
rect 23572 18634 23624 18640
rect 23480 17808 23532 17814
rect 23480 17750 23532 17756
rect 23388 17672 23440 17678
rect 23388 17614 23440 17620
rect 23296 17604 23348 17610
rect 23296 17546 23348 17552
rect 23204 16652 23256 16658
rect 23204 16594 23256 16600
rect 23204 16516 23256 16522
rect 23204 16458 23256 16464
rect 23032 16238 23152 16266
rect 22836 15700 22888 15706
rect 22836 15642 22888 15648
rect 22928 15700 22980 15706
rect 22928 15642 22980 15648
rect 22848 14498 22876 15642
rect 22756 14482 22876 14498
rect 22744 14476 22876 14482
rect 22796 14470 22876 14476
rect 22744 14418 22796 14424
rect 22836 14408 22888 14414
rect 22836 14350 22888 14356
rect 22558 13424 22614 13433
rect 22558 13359 22614 13368
rect 22652 12980 22704 12986
rect 22652 12922 22704 12928
rect 22100 11630 22152 11636
rect 22204 11614 22416 11642
rect 22468 11688 22520 11694
rect 22468 11630 22520 11636
rect 21914 11112 21970 11121
rect 21914 11047 21970 11056
rect 21928 11014 21956 11047
rect 21916 11008 21968 11014
rect 21916 10950 21968 10956
rect 22100 10736 22152 10742
rect 22100 10678 22152 10684
rect 21824 10600 21876 10606
rect 21824 10542 21876 10548
rect 22008 10600 22060 10606
rect 22008 10542 22060 10548
rect 21640 10464 21692 10470
rect 21640 10406 21692 10412
rect 21732 10464 21784 10470
rect 21732 10406 21784 10412
rect 21652 7018 21680 10406
rect 21744 10266 21772 10406
rect 21732 10260 21784 10266
rect 21732 10202 21784 10208
rect 21732 10056 21784 10062
rect 21732 9998 21784 10004
rect 21744 9042 21772 9998
rect 21836 9042 21864 10542
rect 22020 9994 22048 10542
rect 22008 9988 22060 9994
rect 22008 9930 22060 9936
rect 21916 9648 21968 9654
rect 21916 9590 21968 9596
rect 21928 9518 21956 9590
rect 22112 9586 22140 10678
rect 22204 10010 22232 11614
rect 22284 11552 22336 11558
rect 22284 11494 22336 11500
rect 22296 11218 22324 11494
rect 22376 11348 22428 11354
rect 22376 11290 22428 11296
rect 22284 11212 22336 11218
rect 22284 11154 22336 11160
rect 22296 10130 22324 11154
rect 22388 10606 22416 11290
rect 22480 11218 22508 11630
rect 22560 11620 22612 11626
rect 22560 11562 22612 11568
rect 22468 11212 22520 11218
rect 22468 11154 22520 11160
rect 22572 10810 22600 11562
rect 22560 10804 22612 10810
rect 22560 10746 22612 10752
rect 22376 10600 22428 10606
rect 22376 10542 22428 10548
rect 22468 10600 22520 10606
rect 22468 10542 22520 10548
rect 22284 10124 22336 10130
rect 22284 10066 22336 10072
rect 22204 9982 22324 10010
rect 22100 9580 22152 9586
rect 22100 9522 22152 9528
rect 21916 9512 21968 9518
rect 21916 9454 21968 9460
rect 22008 9512 22060 9518
rect 22008 9454 22060 9460
rect 21732 9036 21784 9042
rect 21732 8978 21784 8984
rect 21824 9036 21876 9042
rect 21824 8978 21876 8984
rect 21836 8430 21864 8978
rect 22020 8838 22048 9454
rect 22008 8832 22060 8838
rect 22008 8774 22060 8780
rect 21824 8424 21876 8430
rect 21824 8366 21876 8372
rect 21836 7954 21864 8366
rect 22112 8090 22140 9522
rect 22296 9110 22324 9982
rect 22388 9926 22416 10542
rect 22376 9920 22428 9926
rect 22376 9862 22428 9868
rect 22284 9104 22336 9110
rect 22284 9046 22336 9052
rect 22374 9072 22430 9081
rect 22374 9007 22430 9016
rect 22284 8968 22336 8974
rect 22284 8910 22336 8916
rect 22100 8084 22152 8090
rect 22100 8026 22152 8032
rect 21824 7948 21876 7954
rect 21824 7890 21876 7896
rect 22008 7880 22060 7886
rect 22008 7822 22060 7828
rect 21732 7472 21784 7478
rect 21730 7440 21732 7449
rect 21784 7440 21786 7449
rect 22020 7426 22048 7822
rect 21730 7375 21786 7384
rect 21928 7398 22048 7426
rect 22192 7404 22244 7410
rect 21928 7342 21956 7398
rect 22192 7346 22244 7352
rect 21916 7336 21968 7342
rect 22100 7336 22152 7342
rect 21916 7278 21968 7284
rect 22020 7296 22100 7324
rect 21824 7200 21876 7206
rect 21824 7142 21876 7148
rect 21548 6996 21600 7002
rect 21652 6990 21772 7018
rect 21548 6938 21600 6944
rect 21560 4282 21588 6938
rect 21640 6860 21692 6866
rect 21640 6802 21692 6808
rect 21652 5574 21680 6802
rect 21744 5846 21772 6990
rect 21836 6730 21864 7142
rect 21928 7002 21956 7278
rect 21916 6996 21968 7002
rect 21916 6938 21968 6944
rect 22020 6934 22048 7296
rect 22100 7278 22152 7284
rect 22008 6928 22060 6934
rect 22008 6870 22060 6876
rect 21824 6724 21876 6730
rect 21824 6666 21876 6672
rect 22020 6254 22048 6870
rect 22100 6792 22152 6798
rect 22100 6734 22152 6740
rect 22008 6248 22060 6254
rect 22008 6190 22060 6196
rect 21732 5840 21784 5846
rect 21732 5782 21784 5788
rect 22112 5681 22140 6734
rect 22204 5914 22232 7346
rect 22296 7274 22324 8910
rect 22388 8566 22416 9007
rect 22376 8560 22428 8566
rect 22376 8502 22428 8508
rect 22388 8430 22416 8502
rect 22480 8430 22508 10542
rect 22560 10124 22612 10130
rect 22560 10066 22612 10072
rect 22376 8424 22428 8430
rect 22376 8366 22428 8372
rect 22468 8424 22520 8430
rect 22468 8366 22520 8372
rect 22284 7268 22336 7274
rect 22284 7210 22336 7216
rect 22192 5908 22244 5914
rect 22192 5850 22244 5856
rect 22296 5710 22324 7210
rect 22480 6866 22508 8366
rect 22468 6860 22520 6866
rect 22468 6802 22520 6808
rect 22572 6746 22600 10066
rect 22664 6866 22692 12922
rect 22848 10742 22876 14350
rect 22928 14272 22980 14278
rect 22928 14214 22980 14220
rect 22940 12646 22968 14214
rect 23032 13938 23060 16238
rect 23112 16176 23164 16182
rect 23112 16118 23164 16124
rect 23020 13932 23072 13938
rect 23020 13874 23072 13880
rect 22928 12640 22980 12646
rect 22928 12582 22980 12588
rect 22836 10736 22888 10742
rect 22836 10678 22888 10684
rect 22836 10532 22888 10538
rect 22836 10474 22888 10480
rect 22744 9920 22796 9926
rect 22744 9862 22796 9868
rect 22652 6860 22704 6866
rect 22652 6802 22704 6808
rect 22480 6718 22600 6746
rect 22480 5778 22508 6718
rect 22560 6656 22612 6662
rect 22560 6598 22612 6604
rect 22468 5772 22520 5778
rect 22468 5714 22520 5720
rect 22284 5704 22336 5710
rect 22098 5672 22154 5681
rect 22284 5646 22336 5652
rect 22098 5607 22154 5616
rect 21640 5568 21692 5574
rect 21640 5510 21692 5516
rect 21652 5166 21680 5510
rect 21640 5160 21692 5166
rect 21640 5102 21692 5108
rect 21548 4276 21600 4282
rect 21548 4218 21600 4224
rect 21560 3670 21588 4218
rect 21548 3664 21600 3670
rect 21548 3606 21600 3612
rect 21652 3602 21680 5102
rect 22480 4554 22508 5714
rect 22468 4548 22520 4554
rect 22468 4490 22520 4496
rect 22572 4486 22600 6598
rect 22664 5778 22692 6802
rect 22652 5772 22704 5778
rect 22652 5714 22704 5720
rect 22664 5302 22692 5714
rect 22652 5296 22704 5302
rect 22652 5238 22704 5244
rect 22664 4758 22692 5238
rect 22756 4826 22784 9862
rect 22848 9178 22876 10474
rect 22940 9518 22968 12582
rect 22928 9512 22980 9518
rect 22928 9454 22980 9460
rect 22836 9172 22888 9178
rect 22836 9114 22888 9120
rect 23020 8628 23072 8634
rect 23020 8570 23072 8576
rect 22928 8424 22980 8430
rect 22928 8366 22980 8372
rect 22940 7954 22968 8366
rect 22928 7948 22980 7954
rect 22928 7890 22980 7896
rect 22836 7540 22888 7546
rect 22836 7482 22888 7488
rect 22848 7342 22876 7482
rect 22836 7336 22888 7342
rect 22836 7278 22888 7284
rect 22848 6254 22876 7278
rect 22836 6248 22888 6254
rect 22836 6190 22888 6196
rect 22926 5672 22982 5681
rect 22926 5607 22982 5616
rect 22940 5166 22968 5607
rect 22928 5160 22980 5166
rect 22928 5102 22980 5108
rect 22744 4820 22796 4826
rect 22744 4762 22796 4768
rect 22652 4752 22704 4758
rect 22652 4694 22704 4700
rect 22940 4690 22968 5102
rect 22928 4684 22980 4690
rect 22928 4626 22980 4632
rect 22744 4548 22796 4554
rect 22744 4490 22796 4496
rect 22560 4480 22612 4486
rect 22560 4422 22612 4428
rect 22100 4208 22152 4214
rect 22100 4150 22152 4156
rect 22112 4078 22140 4150
rect 22100 4072 22152 4078
rect 22020 4032 22100 4060
rect 22020 3942 22048 4032
rect 22100 4014 22152 4020
rect 22376 4072 22428 4078
rect 22376 4014 22428 4020
rect 22560 4072 22612 4078
rect 22560 4014 22612 4020
rect 22008 3936 22060 3942
rect 22008 3878 22060 3884
rect 21640 3596 21692 3602
rect 21640 3538 21692 3544
rect 22388 2650 22416 4014
rect 22572 3126 22600 4014
rect 22756 3602 22784 4490
rect 23032 3602 23060 8570
rect 23124 6866 23152 16118
rect 23216 15978 23244 16458
rect 23204 15972 23256 15978
rect 23204 15914 23256 15920
rect 23216 15570 23244 15914
rect 23204 15564 23256 15570
rect 23204 15506 23256 15512
rect 23216 15162 23244 15506
rect 23204 15156 23256 15162
rect 23204 15098 23256 15104
rect 23216 14414 23244 15098
rect 23296 14952 23348 14958
rect 23296 14894 23348 14900
rect 23204 14408 23256 14414
rect 23204 14350 23256 14356
rect 23216 13326 23244 14350
rect 23308 13870 23336 14894
rect 23400 14618 23428 17614
rect 23584 17542 23612 18634
rect 23676 18222 23704 18770
rect 23664 18216 23716 18222
rect 23664 18158 23716 18164
rect 23664 17740 23716 17746
rect 23664 17682 23716 17688
rect 23572 17536 23624 17542
rect 23572 17478 23624 17484
rect 23572 17332 23624 17338
rect 23572 17274 23624 17280
rect 23584 16726 23612 17274
rect 23572 16720 23624 16726
rect 23572 16662 23624 16668
rect 23676 16658 23704 17682
rect 23768 17134 23796 25978
rect 24032 25356 24084 25362
rect 24032 25298 24084 25304
rect 24044 24274 24072 25298
rect 24228 24750 24256 27474
rect 24320 25226 24348 31214
rect 24492 31136 24544 31142
rect 24492 31078 24544 31084
rect 24504 30433 24532 31078
rect 24780 30818 24808 35090
rect 25976 34950 26004 39200
rect 26240 37120 26292 37126
rect 26240 37062 26292 37068
rect 26252 36242 26280 37062
rect 26516 36712 26568 36718
rect 26516 36654 26568 36660
rect 27160 36712 27212 36718
rect 27160 36654 27212 36660
rect 26240 36236 26292 36242
rect 26240 36178 26292 36184
rect 26528 36174 26556 36654
rect 27172 36378 27200 36654
rect 27160 36372 27212 36378
rect 27160 36314 27212 36320
rect 26516 36168 26568 36174
rect 26516 36110 26568 36116
rect 26528 35698 26556 36110
rect 28000 35834 28028 39200
rect 30024 37346 30052 39200
rect 32048 37398 32076 39200
rect 29184 37324 29236 37330
rect 29184 37266 29236 37272
rect 29932 37318 30052 37346
rect 32036 37392 32088 37398
rect 32036 37334 32088 37340
rect 33140 37324 33192 37330
rect 29000 37256 29052 37262
rect 29000 37198 29052 37204
rect 28908 36644 28960 36650
rect 28908 36586 28960 36592
rect 28920 36242 28948 36586
rect 28908 36236 28960 36242
rect 28908 36178 28960 36184
rect 29012 36174 29040 37198
rect 29000 36168 29052 36174
rect 29000 36110 29052 36116
rect 29012 35834 29040 36110
rect 27988 35828 28040 35834
rect 27988 35770 28040 35776
rect 29000 35828 29052 35834
rect 29000 35770 29052 35776
rect 26516 35692 26568 35698
rect 26516 35634 26568 35640
rect 28908 35692 28960 35698
rect 28908 35634 28960 35640
rect 26332 35624 26384 35630
rect 26332 35566 26384 35572
rect 25964 34944 26016 34950
rect 25964 34886 26016 34892
rect 25504 34604 25556 34610
rect 25504 34546 25556 34552
rect 24952 33992 25004 33998
rect 24952 33934 25004 33940
rect 24964 33658 24992 33934
rect 24952 33652 25004 33658
rect 24952 33594 25004 33600
rect 25516 32502 25544 34546
rect 25872 33856 25924 33862
rect 25872 33798 25924 33804
rect 25964 33856 26016 33862
rect 25964 33798 26016 33804
rect 25780 33448 25832 33454
rect 25780 33390 25832 33396
rect 25792 32842 25820 33390
rect 25780 32836 25832 32842
rect 25780 32778 25832 32784
rect 25504 32496 25556 32502
rect 25504 32438 25556 32444
rect 25320 32360 25372 32366
rect 25320 32302 25372 32308
rect 25228 32224 25280 32230
rect 25228 32166 25280 32172
rect 24860 31884 24912 31890
rect 24860 31826 24912 31832
rect 24872 30938 24900 31826
rect 25240 31414 25268 32166
rect 25332 31822 25360 32302
rect 25320 31816 25372 31822
rect 25320 31758 25372 31764
rect 25228 31408 25280 31414
rect 25228 31350 25280 31356
rect 24860 30932 24912 30938
rect 24860 30874 24912 30880
rect 25136 30864 25188 30870
rect 24780 30790 24900 30818
rect 25136 30806 25188 30812
rect 24490 30424 24546 30433
rect 24490 30359 24546 30368
rect 24768 29708 24820 29714
rect 24768 29650 24820 29656
rect 24676 29164 24728 29170
rect 24676 29106 24728 29112
rect 24688 28014 24716 29106
rect 24780 29102 24808 29650
rect 24768 29096 24820 29102
rect 24768 29038 24820 29044
rect 24676 28008 24728 28014
rect 24676 27950 24728 27956
rect 24492 26852 24544 26858
rect 24492 26794 24544 26800
rect 24400 25832 24452 25838
rect 24400 25774 24452 25780
rect 24308 25220 24360 25226
rect 24308 25162 24360 25168
rect 24412 24993 24440 25774
rect 24504 25702 24532 26794
rect 24584 26444 24636 26450
rect 24584 26386 24636 26392
rect 24492 25696 24544 25702
rect 24492 25638 24544 25644
rect 24504 25362 24532 25638
rect 24492 25356 24544 25362
rect 24492 25298 24544 25304
rect 24492 25220 24544 25226
rect 24492 25162 24544 25168
rect 24398 24984 24454 24993
rect 24398 24919 24454 24928
rect 24216 24744 24268 24750
rect 24216 24686 24268 24692
rect 24400 24608 24452 24614
rect 24504 24596 24532 25162
rect 24452 24568 24532 24596
rect 24400 24550 24452 24556
rect 24032 24268 24084 24274
rect 24032 24210 24084 24216
rect 24032 23860 24084 23866
rect 24032 23802 24084 23808
rect 23940 23724 23992 23730
rect 23940 23666 23992 23672
rect 23848 23180 23900 23186
rect 23848 23122 23900 23128
rect 23860 20262 23888 23122
rect 23848 20256 23900 20262
rect 23848 20198 23900 20204
rect 23860 20058 23888 20198
rect 23848 20052 23900 20058
rect 23952 20040 23980 23666
rect 24044 23254 24072 23802
rect 24412 23508 24440 24550
rect 24596 24426 24624 26386
rect 24688 25838 24716 27950
rect 24780 26926 24808 29038
rect 24872 28778 24900 30790
rect 24952 30728 25004 30734
rect 24952 30670 25004 30676
rect 24964 30326 24992 30670
rect 24952 30320 25004 30326
rect 24952 30262 25004 30268
rect 25044 30116 25096 30122
rect 25044 30058 25096 30064
rect 25056 29714 25084 30058
rect 25044 29708 25096 29714
rect 25044 29650 25096 29656
rect 24872 28750 25084 28778
rect 24860 28620 24912 28626
rect 24860 28562 24912 28568
rect 24952 28620 25004 28626
rect 24952 28562 25004 28568
rect 24872 28150 24900 28562
rect 24860 28144 24912 28150
rect 24860 28086 24912 28092
rect 24964 27130 24992 28562
rect 24952 27124 25004 27130
rect 24952 27066 25004 27072
rect 24768 26920 24820 26926
rect 24768 26862 24820 26868
rect 24780 26382 24808 26862
rect 24768 26376 24820 26382
rect 24768 26318 24820 26324
rect 25056 26042 25084 28750
rect 25148 28014 25176 30806
rect 25332 29102 25360 31758
rect 25412 31272 25464 31278
rect 25412 31214 25464 31220
rect 25424 30666 25452 31214
rect 25412 30660 25464 30666
rect 25412 30602 25464 30608
rect 25516 29714 25544 32438
rect 25884 31346 25912 33798
rect 25976 32978 26004 33798
rect 25964 32972 26016 32978
rect 25964 32914 26016 32920
rect 25964 32836 26016 32842
rect 25964 32778 26016 32784
rect 25976 32366 26004 32778
rect 25964 32360 26016 32366
rect 25964 32302 26016 32308
rect 25976 31482 26004 32302
rect 25964 31476 26016 31482
rect 25964 31418 26016 31424
rect 25872 31340 25924 31346
rect 25872 31282 25924 31288
rect 25596 31272 25648 31278
rect 25596 31214 25648 31220
rect 25780 31272 25832 31278
rect 25780 31214 25832 31220
rect 25608 30258 25636 31214
rect 25596 30252 25648 30258
rect 25596 30194 25648 30200
rect 25792 29850 25820 31214
rect 25780 29844 25832 29850
rect 25780 29786 25832 29792
rect 25504 29708 25556 29714
rect 25504 29650 25556 29656
rect 25228 29096 25280 29102
rect 25228 29038 25280 29044
rect 25320 29096 25372 29102
rect 25320 29038 25372 29044
rect 25136 28008 25188 28014
rect 25136 27950 25188 27956
rect 25148 26518 25176 27950
rect 25136 26512 25188 26518
rect 25136 26454 25188 26460
rect 25044 26036 25096 26042
rect 25044 25978 25096 25984
rect 24676 25832 24728 25838
rect 24676 25774 24728 25780
rect 24768 25832 24820 25838
rect 24768 25774 24820 25780
rect 24688 24614 24716 25774
rect 24780 25430 24808 25774
rect 24768 25424 24820 25430
rect 24768 25366 24820 25372
rect 24676 24608 24728 24614
rect 24676 24550 24728 24556
rect 24504 24398 24716 24426
rect 24504 23662 24532 24398
rect 24688 24206 24716 24398
rect 24780 24274 24808 25366
rect 25044 24948 25096 24954
rect 25044 24890 25096 24896
rect 24952 24744 25004 24750
rect 24952 24686 25004 24692
rect 24964 24410 24992 24686
rect 24952 24404 25004 24410
rect 24952 24346 25004 24352
rect 25056 24274 25084 24890
rect 25240 24342 25268 29038
rect 25320 28620 25372 28626
rect 25320 28562 25372 28568
rect 25332 27062 25360 28562
rect 25320 27056 25372 27062
rect 25320 26998 25372 27004
rect 25884 26926 25912 31282
rect 26056 29708 26108 29714
rect 26056 29650 26108 29656
rect 26068 29102 26096 29650
rect 26056 29096 26108 29102
rect 26056 29038 26108 29044
rect 26068 28694 26096 29038
rect 26148 29028 26200 29034
rect 26148 28970 26200 28976
rect 26056 28688 26108 28694
rect 26056 28630 26108 28636
rect 26068 28014 26096 28630
rect 26056 28008 26108 28014
rect 26056 27950 26108 27956
rect 26068 26926 26096 27950
rect 25596 26920 25648 26926
rect 25596 26862 25648 26868
rect 25872 26920 25924 26926
rect 25872 26862 25924 26868
rect 26056 26920 26108 26926
rect 26056 26862 26108 26868
rect 25320 26512 25372 26518
rect 25320 26454 25372 26460
rect 25228 24336 25280 24342
rect 25228 24278 25280 24284
rect 24768 24268 24820 24274
rect 24768 24210 24820 24216
rect 25044 24268 25096 24274
rect 25044 24210 25096 24216
rect 24584 24200 24636 24206
rect 24584 24142 24636 24148
rect 24676 24200 24728 24206
rect 24676 24142 24728 24148
rect 24492 23656 24544 23662
rect 24492 23598 24544 23604
rect 24412 23480 24532 23508
rect 24032 23248 24084 23254
rect 24032 23190 24084 23196
rect 24216 23180 24268 23186
rect 24216 23122 24268 23128
rect 24124 22568 24176 22574
rect 24124 22510 24176 22516
rect 24136 21554 24164 22510
rect 24228 22506 24256 23122
rect 24400 23112 24452 23118
rect 24400 23054 24452 23060
rect 24412 22642 24440 23054
rect 24400 22636 24452 22642
rect 24400 22578 24452 22584
rect 24216 22500 24268 22506
rect 24216 22442 24268 22448
rect 24124 21548 24176 21554
rect 24124 21490 24176 21496
rect 24032 21480 24084 21486
rect 24032 21422 24084 21428
rect 24044 21010 24072 21422
rect 24136 21010 24164 21490
rect 24032 21004 24084 21010
rect 24032 20946 24084 20952
rect 24124 21004 24176 21010
rect 24124 20946 24176 20952
rect 24136 20602 24164 20946
rect 24124 20596 24176 20602
rect 24124 20538 24176 20544
rect 23952 20012 24072 20040
rect 23848 19994 23900 20000
rect 23940 19916 23992 19922
rect 23940 19858 23992 19864
rect 23848 18080 23900 18086
rect 23848 18022 23900 18028
rect 23860 17678 23888 18022
rect 23848 17672 23900 17678
rect 23848 17614 23900 17620
rect 23756 17128 23808 17134
rect 23756 17070 23808 17076
rect 23848 17128 23900 17134
rect 23848 17070 23900 17076
rect 23664 16652 23716 16658
rect 23664 16594 23716 16600
rect 23756 15360 23808 15366
rect 23756 15302 23808 15308
rect 23768 14958 23796 15302
rect 23756 14952 23808 14958
rect 23756 14894 23808 14900
rect 23388 14612 23440 14618
rect 23388 14554 23440 14560
rect 23400 14482 23428 14554
rect 23768 14482 23796 14894
rect 23860 14822 23888 17070
rect 23952 16998 23980 19858
rect 23940 16992 23992 16998
rect 23940 16934 23992 16940
rect 23848 14816 23900 14822
rect 23848 14758 23900 14764
rect 23388 14476 23440 14482
rect 23388 14418 23440 14424
rect 23756 14476 23808 14482
rect 23756 14418 23808 14424
rect 23664 14340 23716 14346
rect 23664 14282 23716 14288
rect 23296 13864 23348 13870
rect 23296 13806 23348 13812
rect 23308 13394 23336 13806
rect 23480 13796 23532 13802
rect 23480 13738 23532 13744
rect 23492 13530 23520 13738
rect 23572 13728 23624 13734
rect 23572 13670 23624 13676
rect 23480 13524 23532 13530
rect 23480 13466 23532 13472
rect 23296 13388 23348 13394
rect 23296 13330 23348 13336
rect 23204 13320 23256 13326
rect 23204 13262 23256 13268
rect 23492 12850 23520 13466
rect 23480 12844 23532 12850
rect 23480 12786 23532 12792
rect 23584 12782 23612 13670
rect 23572 12776 23624 12782
rect 23572 12718 23624 12724
rect 23296 10532 23348 10538
rect 23296 10474 23348 10480
rect 23308 10130 23336 10474
rect 23296 10124 23348 10130
rect 23296 10066 23348 10072
rect 23204 10056 23256 10062
rect 23204 9998 23256 10004
rect 23216 9586 23244 9998
rect 23296 9920 23348 9926
rect 23296 9862 23348 9868
rect 23204 9580 23256 9586
rect 23204 9522 23256 9528
rect 23216 8974 23244 9522
rect 23204 8968 23256 8974
rect 23204 8910 23256 8916
rect 23216 8430 23244 8910
rect 23204 8424 23256 8430
rect 23204 8366 23256 8372
rect 23204 8084 23256 8090
rect 23204 8026 23256 8032
rect 23216 7954 23244 8026
rect 23204 7948 23256 7954
rect 23204 7890 23256 7896
rect 23112 6860 23164 6866
rect 23112 6802 23164 6808
rect 23124 5778 23152 6802
rect 23112 5772 23164 5778
rect 23112 5714 23164 5720
rect 23124 5370 23152 5714
rect 23112 5364 23164 5370
rect 23112 5306 23164 5312
rect 23308 4690 23336 9862
rect 23480 8968 23532 8974
rect 23480 8910 23532 8916
rect 23388 8424 23440 8430
rect 23388 8366 23440 8372
rect 23400 6866 23428 8366
rect 23492 8090 23520 8910
rect 23480 8084 23532 8090
rect 23480 8026 23532 8032
rect 23388 6860 23440 6866
rect 23388 6802 23440 6808
rect 23584 6254 23612 12718
rect 23676 12102 23704 14282
rect 23768 13870 23796 14418
rect 23756 13864 23808 13870
rect 23756 13806 23808 13812
rect 23756 12776 23808 12782
rect 23756 12718 23808 12724
rect 23768 12238 23796 12718
rect 23756 12232 23808 12238
rect 23756 12174 23808 12180
rect 23664 12096 23716 12102
rect 23664 12038 23716 12044
rect 23676 10742 23704 12038
rect 23664 10736 23716 10742
rect 23664 10678 23716 10684
rect 23664 10600 23716 10606
rect 23664 10542 23716 10548
rect 23676 7002 23704 10542
rect 23860 8922 23888 14758
rect 24044 14464 24072 20012
rect 24124 17740 24176 17746
rect 24124 17682 24176 17688
rect 24136 16658 24164 17682
rect 24124 16652 24176 16658
rect 24124 16594 24176 16600
rect 23952 14436 24072 14464
rect 24124 14476 24176 14482
rect 23952 13734 23980 14436
rect 24124 14418 24176 14424
rect 24032 14340 24084 14346
rect 24032 14282 24084 14288
rect 23940 13728 23992 13734
rect 23940 13670 23992 13676
rect 23940 13252 23992 13258
rect 23940 13194 23992 13200
rect 23952 12850 23980 13194
rect 23940 12844 23992 12850
rect 23940 12786 23992 12792
rect 24044 12306 24072 14282
rect 24136 13394 24164 14418
rect 24124 13388 24176 13394
rect 24124 13330 24176 13336
rect 24228 12782 24256 22442
rect 24504 22166 24532 23480
rect 24596 22982 24624 24142
rect 24676 24064 24728 24070
rect 24676 24006 24728 24012
rect 24688 23730 24716 24006
rect 25056 23866 25084 24210
rect 25044 23860 25096 23866
rect 25044 23802 25096 23808
rect 24676 23724 24728 23730
rect 24676 23666 24728 23672
rect 24860 23656 24912 23662
rect 24860 23598 24912 23604
rect 24872 23118 24900 23598
rect 24860 23112 24912 23118
rect 24860 23054 24912 23060
rect 25332 23050 25360 26454
rect 25412 25152 25464 25158
rect 25412 25094 25464 25100
rect 25424 24750 25452 25094
rect 25608 24886 25636 26862
rect 26068 26586 26096 26862
rect 26056 26580 26108 26586
rect 26056 26522 26108 26528
rect 25688 26036 25740 26042
rect 25688 25978 25740 25984
rect 25596 24880 25648 24886
rect 25596 24822 25648 24828
rect 25412 24744 25464 24750
rect 25412 24686 25464 24692
rect 25700 24274 25728 25978
rect 26160 25362 26188 28970
rect 26240 27940 26292 27946
rect 26240 27882 26292 27888
rect 26252 27538 26280 27882
rect 26240 27532 26292 27538
rect 26240 27474 26292 27480
rect 26148 25356 26200 25362
rect 26148 25298 26200 25304
rect 26160 24750 26188 25298
rect 26148 24744 26200 24750
rect 26148 24686 26200 24692
rect 25688 24268 25740 24274
rect 25688 24210 25740 24216
rect 25700 23594 25728 24210
rect 25688 23588 25740 23594
rect 25688 23530 25740 23536
rect 26160 23526 26188 24686
rect 26148 23520 26200 23526
rect 26148 23462 26200 23468
rect 25320 23044 25372 23050
rect 25320 22986 25372 22992
rect 24584 22976 24636 22982
rect 24584 22918 24636 22924
rect 24952 22500 25004 22506
rect 24952 22442 25004 22448
rect 24492 22160 24544 22166
rect 24492 22102 24544 22108
rect 24964 22030 24992 22442
rect 25412 22092 25464 22098
rect 25412 22034 25464 22040
rect 24400 22024 24452 22030
rect 24400 21966 24452 21972
rect 24952 22024 25004 22030
rect 24952 21966 25004 21972
rect 24412 21350 24440 21966
rect 24400 21344 24452 21350
rect 24400 21286 24452 21292
rect 24308 21072 24360 21078
rect 24308 21014 24360 21020
rect 24320 13530 24348 21014
rect 24400 19304 24452 19310
rect 24400 19246 24452 19252
rect 24860 19304 24912 19310
rect 24860 19246 24912 19252
rect 24412 18834 24440 19246
rect 24768 19236 24820 19242
rect 24768 19178 24820 19184
rect 24584 18896 24636 18902
rect 24584 18838 24636 18844
rect 24400 18828 24452 18834
rect 24400 18770 24452 18776
rect 24412 17882 24440 18770
rect 24492 18080 24544 18086
rect 24492 18022 24544 18028
rect 24400 17876 24452 17882
rect 24400 17818 24452 17824
rect 24412 17338 24440 17818
rect 24400 17332 24452 17338
rect 24400 17274 24452 17280
rect 24504 17134 24532 18022
rect 24596 17746 24624 18838
rect 24780 18834 24808 19178
rect 24872 18902 24900 19246
rect 24860 18896 24912 18902
rect 24860 18838 24912 18844
rect 24768 18828 24820 18834
rect 24768 18770 24820 18776
rect 24584 17740 24636 17746
rect 24584 17682 24636 17688
rect 24860 17740 24912 17746
rect 24860 17682 24912 17688
rect 24676 17604 24728 17610
rect 24676 17546 24728 17552
rect 24492 17128 24544 17134
rect 24492 17070 24544 17076
rect 24400 17060 24452 17066
rect 24400 17002 24452 17008
rect 24412 15570 24440 17002
rect 24584 16992 24636 16998
rect 24584 16934 24636 16940
rect 24400 15564 24452 15570
rect 24400 15506 24452 15512
rect 24400 14952 24452 14958
rect 24400 14894 24452 14900
rect 24308 13524 24360 13530
rect 24308 13466 24360 13472
rect 24216 12776 24268 12782
rect 24216 12718 24268 12724
rect 24032 12300 24084 12306
rect 24032 12242 24084 12248
rect 24216 11892 24268 11898
rect 24216 11834 24268 11840
rect 24228 11354 24256 11834
rect 24216 11348 24268 11354
rect 24216 11290 24268 11296
rect 23940 10736 23992 10742
rect 23940 10678 23992 10684
rect 23952 9722 23980 10678
rect 23940 9716 23992 9722
rect 23940 9658 23992 9664
rect 24216 9512 24268 9518
rect 24216 9454 24268 9460
rect 24032 9376 24084 9382
rect 24032 9318 24084 9324
rect 23768 8894 23888 8922
rect 23768 8022 23796 8894
rect 23848 8832 23900 8838
rect 23848 8774 23900 8780
rect 23756 8016 23808 8022
rect 23756 7958 23808 7964
rect 23860 7342 23888 8774
rect 24044 8566 24072 9318
rect 24032 8560 24084 8566
rect 24032 8502 24084 8508
rect 24228 8430 24256 9454
rect 24216 8424 24268 8430
rect 24216 8366 24268 8372
rect 24320 8022 24348 13466
rect 24412 9330 24440 14894
rect 24596 13870 24624 16934
rect 24688 16658 24716 17546
rect 24872 17270 24900 17682
rect 24860 17264 24912 17270
rect 24860 17206 24912 17212
rect 24872 16658 24900 17206
rect 24964 17134 24992 21966
rect 25136 19984 25188 19990
rect 25136 19926 25188 19932
rect 25148 19310 25176 19926
rect 25228 19712 25280 19718
rect 25226 19680 25228 19689
rect 25280 19680 25282 19689
rect 25226 19615 25282 19624
rect 25044 19304 25096 19310
rect 25042 19272 25044 19281
rect 25136 19304 25188 19310
rect 25096 19272 25098 19281
rect 25136 19246 25188 19252
rect 25042 19207 25098 19216
rect 25148 18834 25176 19246
rect 25136 18828 25188 18834
rect 25136 18770 25188 18776
rect 25424 18154 25452 22034
rect 26056 20392 26108 20398
rect 26056 20334 26108 20340
rect 25872 20256 25924 20262
rect 25872 20198 25924 20204
rect 25884 19514 25912 20198
rect 26068 20058 26096 20334
rect 26056 20052 26108 20058
rect 26056 19994 26108 20000
rect 25872 19508 25924 19514
rect 25872 19450 25924 19456
rect 25884 18834 25912 19450
rect 26148 19304 26200 19310
rect 26148 19246 26200 19252
rect 25964 19168 26016 19174
rect 25964 19110 26016 19116
rect 25872 18828 25924 18834
rect 25872 18770 25924 18776
rect 25504 18216 25556 18222
rect 25504 18158 25556 18164
rect 25872 18216 25924 18222
rect 25872 18158 25924 18164
rect 25044 18148 25096 18154
rect 25044 18090 25096 18096
rect 25412 18148 25464 18154
rect 25412 18090 25464 18096
rect 24952 17128 25004 17134
rect 24952 17070 25004 17076
rect 24676 16652 24728 16658
rect 24676 16594 24728 16600
rect 24860 16652 24912 16658
rect 24860 16594 24912 16600
rect 24952 16652 25004 16658
rect 24952 16594 25004 16600
rect 24766 16144 24822 16153
rect 24766 16079 24768 16088
rect 24820 16079 24822 16088
rect 24768 16050 24820 16056
rect 24964 16046 24992 16594
rect 24952 16040 25004 16046
rect 24952 15982 25004 15988
rect 24952 15496 25004 15502
rect 24952 15438 25004 15444
rect 24964 14482 24992 15438
rect 24952 14476 25004 14482
rect 24952 14418 25004 14424
rect 24584 13864 24636 13870
rect 24584 13806 24636 13812
rect 24860 13728 24912 13734
rect 24860 13670 24912 13676
rect 24872 12782 24900 13670
rect 25056 13394 25084 18090
rect 25516 16522 25544 18158
rect 25688 17740 25740 17746
rect 25688 17682 25740 17688
rect 25700 16658 25728 17682
rect 25780 17672 25832 17678
rect 25780 17614 25832 17620
rect 25792 17134 25820 17614
rect 25884 17542 25912 18158
rect 25976 17882 26004 19110
rect 26056 18896 26108 18902
rect 26056 18838 26108 18844
rect 26068 18154 26096 18838
rect 26056 18148 26108 18154
rect 26056 18090 26108 18096
rect 25964 17876 26016 17882
rect 25964 17818 26016 17824
rect 25872 17536 25924 17542
rect 25872 17478 25924 17484
rect 25780 17128 25832 17134
rect 25780 17070 25832 17076
rect 25780 16788 25832 16794
rect 25780 16730 25832 16736
rect 25688 16652 25740 16658
rect 25688 16594 25740 16600
rect 25504 16516 25556 16522
rect 25504 16458 25556 16464
rect 25516 15570 25544 16458
rect 25792 15570 25820 16730
rect 25504 15564 25556 15570
rect 25504 15506 25556 15512
rect 25780 15564 25832 15570
rect 25780 15506 25832 15512
rect 25688 14952 25740 14958
rect 25688 14894 25740 14900
rect 25700 14618 25728 14894
rect 25688 14612 25740 14618
rect 25688 14554 25740 14560
rect 25320 13864 25372 13870
rect 25320 13806 25372 13812
rect 25044 13388 25096 13394
rect 25044 13330 25096 13336
rect 24676 12776 24728 12782
rect 24676 12718 24728 12724
rect 24860 12776 24912 12782
rect 24860 12718 24912 12724
rect 24688 11762 24716 12718
rect 24676 11756 24728 11762
rect 24676 11698 24728 11704
rect 24872 11354 24900 12718
rect 25332 11626 25360 13806
rect 25884 13802 25912 17478
rect 26160 16794 26188 19246
rect 26240 19168 26292 19174
rect 26240 19110 26292 19116
rect 26252 18358 26280 19110
rect 26240 18352 26292 18358
rect 26240 18294 26292 18300
rect 26240 17672 26292 17678
rect 26240 17614 26292 17620
rect 26148 16788 26200 16794
rect 26148 16730 26200 16736
rect 25964 15020 26016 15026
rect 25964 14962 26016 14968
rect 25976 14482 26004 14962
rect 26148 14612 26200 14618
rect 26148 14554 26200 14560
rect 25964 14476 26016 14482
rect 25964 14418 26016 14424
rect 25872 13796 25924 13802
rect 25872 13738 25924 13744
rect 25688 13728 25740 13734
rect 25688 13670 25740 13676
rect 25700 13394 25728 13670
rect 25688 13388 25740 13394
rect 25688 13330 25740 13336
rect 25504 12708 25556 12714
rect 25504 12650 25556 12656
rect 25516 12238 25544 12650
rect 25872 12640 25924 12646
rect 25872 12582 25924 12588
rect 25504 12232 25556 12238
rect 25504 12174 25556 12180
rect 25516 11830 25544 12174
rect 25596 12096 25648 12102
rect 25596 12038 25648 12044
rect 25504 11824 25556 11830
rect 25504 11766 25556 11772
rect 25320 11620 25372 11626
rect 25320 11562 25372 11568
rect 25516 11558 25544 11766
rect 25608 11626 25636 12038
rect 25596 11620 25648 11626
rect 25596 11562 25648 11568
rect 25412 11552 25464 11558
rect 25412 11494 25464 11500
rect 25504 11552 25556 11558
rect 25504 11494 25556 11500
rect 24860 11348 24912 11354
rect 24860 11290 24912 11296
rect 25424 10606 25452 11494
rect 25608 11218 25636 11562
rect 25596 11212 25648 11218
rect 25596 11154 25648 11160
rect 24952 10600 25004 10606
rect 24952 10542 25004 10548
rect 25412 10600 25464 10606
rect 25412 10542 25464 10548
rect 24964 9926 24992 10542
rect 25504 10124 25556 10130
rect 25504 10066 25556 10072
rect 25688 10124 25740 10130
rect 25688 10066 25740 10072
rect 24952 9920 25004 9926
rect 24952 9862 25004 9868
rect 25516 9722 25544 10066
rect 25504 9716 25556 9722
rect 25504 9658 25556 9664
rect 25700 9654 25728 10066
rect 25688 9648 25740 9654
rect 25688 9590 25740 9596
rect 25504 9512 25556 9518
rect 25504 9454 25556 9460
rect 24412 9302 24532 9330
rect 24400 8628 24452 8634
rect 24400 8570 24452 8576
rect 24412 8294 24440 8570
rect 24400 8288 24452 8294
rect 24400 8230 24452 8236
rect 24308 8016 24360 8022
rect 24308 7958 24360 7964
rect 24320 7478 24348 7958
rect 24412 7954 24440 8230
rect 24400 7948 24452 7954
rect 24400 7890 24452 7896
rect 24308 7472 24360 7478
rect 24308 7414 24360 7420
rect 23848 7336 23900 7342
rect 23848 7278 23900 7284
rect 24400 7336 24452 7342
rect 24400 7278 24452 7284
rect 23664 6996 23716 7002
rect 23664 6938 23716 6944
rect 23572 6248 23624 6254
rect 23572 6190 23624 6196
rect 23664 6112 23716 6118
rect 23664 6054 23716 6060
rect 23676 5166 23704 6054
rect 23860 5778 23888 7278
rect 24412 7206 24440 7278
rect 24400 7200 24452 7206
rect 24320 7160 24400 7188
rect 24320 5778 24348 7160
rect 24400 7142 24452 7148
rect 24504 6780 24532 9302
rect 25136 7948 25188 7954
rect 25136 7890 25188 7896
rect 25148 7478 25176 7890
rect 25136 7472 25188 7478
rect 24582 7440 24638 7449
rect 25136 7414 25188 7420
rect 24582 7375 24638 7384
rect 24596 7342 24624 7375
rect 24584 7336 24636 7342
rect 24584 7278 24636 7284
rect 24860 7200 24912 7206
rect 24860 7142 24912 7148
rect 24872 6866 24900 7142
rect 24860 6860 24912 6866
rect 24860 6802 24912 6808
rect 24584 6792 24636 6798
rect 24504 6752 24584 6780
rect 24584 6734 24636 6740
rect 23848 5772 23900 5778
rect 23848 5714 23900 5720
rect 24124 5772 24176 5778
rect 24124 5714 24176 5720
rect 24308 5772 24360 5778
rect 24308 5714 24360 5720
rect 23664 5160 23716 5166
rect 23664 5102 23716 5108
rect 23296 4684 23348 4690
rect 23296 4626 23348 4632
rect 23676 4486 23704 5102
rect 24136 4690 24164 5714
rect 24124 4684 24176 4690
rect 24124 4626 24176 4632
rect 23664 4480 23716 4486
rect 23664 4422 23716 4428
rect 24136 4162 24164 4626
rect 24044 4134 24164 4162
rect 24044 3670 24072 4134
rect 24596 4078 24624 6734
rect 25148 6458 25176 7414
rect 25516 6798 25544 9454
rect 25596 7336 25648 7342
rect 25596 7278 25648 7284
rect 25504 6792 25556 6798
rect 25504 6734 25556 6740
rect 25136 6452 25188 6458
rect 25136 6394 25188 6400
rect 25136 6248 25188 6254
rect 25136 6190 25188 6196
rect 25320 6248 25372 6254
rect 25320 6190 25372 6196
rect 24676 5772 24728 5778
rect 24676 5714 24728 5720
rect 24688 4690 24716 5714
rect 25148 5234 25176 6190
rect 25332 5846 25360 6190
rect 25320 5840 25372 5846
rect 25320 5782 25372 5788
rect 24860 5228 24912 5234
rect 24860 5170 24912 5176
rect 25136 5228 25188 5234
rect 25136 5170 25188 5176
rect 24676 4684 24728 4690
rect 24676 4626 24728 4632
rect 24584 4072 24636 4078
rect 24584 4014 24636 4020
rect 24124 4004 24176 4010
rect 24124 3946 24176 3952
rect 24032 3664 24084 3670
rect 24032 3606 24084 3612
rect 22744 3596 22796 3602
rect 22744 3538 22796 3544
rect 23020 3596 23072 3602
rect 23020 3538 23072 3544
rect 22836 3460 22888 3466
rect 22836 3402 22888 3408
rect 22560 3120 22612 3126
rect 22560 3062 22612 3068
rect 22848 3058 22876 3402
rect 23032 3126 23060 3538
rect 23940 3392 23992 3398
rect 23940 3334 23992 3340
rect 23020 3120 23072 3126
rect 23020 3062 23072 3068
rect 23952 3058 23980 3334
rect 22836 3052 22888 3058
rect 22836 2994 22888 3000
rect 23940 3052 23992 3058
rect 23940 2994 23992 3000
rect 23020 2848 23072 2854
rect 23020 2790 23072 2796
rect 22376 2644 22428 2650
rect 22376 2586 22428 2592
rect 21416 2400 21496 2428
rect 21364 2382 21416 2388
rect 20352 2304 20404 2310
rect 20352 2246 20404 2252
rect 20640 2038 20668 2382
rect 20996 2304 21048 2310
rect 20996 2246 21048 2252
rect 20628 2032 20680 2038
rect 20628 1974 20680 1980
rect 20076 1964 20128 1970
rect 20076 1906 20128 1912
rect 21008 800 21036 2246
rect 23032 800 23060 2790
rect 24136 2514 24164 3946
rect 24596 3534 24624 4014
rect 24688 3602 24716 4626
rect 24872 4146 24900 5170
rect 25228 5160 25280 5166
rect 25228 5102 25280 5108
rect 25240 4758 25268 5102
rect 25228 4752 25280 4758
rect 25228 4694 25280 4700
rect 25516 4690 25544 6734
rect 25608 4758 25636 7278
rect 25700 6866 25728 9590
rect 25688 6860 25740 6866
rect 25688 6802 25740 6808
rect 25596 4752 25648 4758
rect 25596 4694 25648 4700
rect 25504 4684 25556 4690
rect 25504 4626 25556 4632
rect 25700 4622 25728 6802
rect 25688 4616 25740 4622
rect 25688 4558 25740 4564
rect 24860 4140 24912 4146
rect 24860 4082 24912 4088
rect 24860 4004 24912 4010
rect 24860 3946 24912 3952
rect 24676 3596 24728 3602
rect 24676 3538 24728 3544
rect 24584 3528 24636 3534
rect 24584 3470 24636 3476
rect 24872 2514 24900 3946
rect 25596 3732 25648 3738
rect 25596 3674 25648 3680
rect 25608 3194 25636 3674
rect 25700 3398 25728 4558
rect 25780 4072 25832 4078
rect 25780 4014 25832 4020
rect 25792 3738 25820 4014
rect 25780 3732 25832 3738
rect 25780 3674 25832 3680
rect 25688 3392 25740 3398
rect 25688 3334 25740 3340
rect 25596 3188 25648 3194
rect 25596 3130 25648 3136
rect 25884 3058 25912 12582
rect 26160 11762 26188 14554
rect 26252 14074 26280 17614
rect 26240 14068 26292 14074
rect 26240 14010 26292 14016
rect 26252 13870 26280 14010
rect 26240 13864 26292 13870
rect 26240 13806 26292 13812
rect 26148 11756 26200 11762
rect 26148 11698 26200 11704
rect 25964 11620 26016 11626
rect 25964 11562 26016 11568
rect 25976 11286 26004 11562
rect 25964 11280 26016 11286
rect 25964 11222 26016 11228
rect 26148 11008 26200 11014
rect 26148 10950 26200 10956
rect 26160 10606 26188 10950
rect 26148 10600 26200 10606
rect 26148 10542 26200 10548
rect 26160 10130 26188 10542
rect 26240 10532 26292 10538
rect 26240 10474 26292 10480
rect 26148 10124 26200 10130
rect 26148 10066 26200 10072
rect 26252 9586 26280 10474
rect 26344 10470 26372 35566
rect 26516 35080 26568 35086
rect 26516 35022 26568 35028
rect 26528 34542 26556 35022
rect 27528 34944 27580 34950
rect 27528 34886 27580 34892
rect 27540 34610 27568 34886
rect 27528 34604 27580 34610
rect 27528 34546 27580 34552
rect 28920 34542 28948 35634
rect 29092 35624 29144 35630
rect 29092 35566 29144 35572
rect 29104 35290 29132 35566
rect 29092 35284 29144 35290
rect 29092 35226 29144 35232
rect 26516 34536 26568 34542
rect 26516 34478 26568 34484
rect 28908 34536 28960 34542
rect 28908 34478 28960 34484
rect 28448 34400 28500 34406
rect 28448 34342 28500 34348
rect 28460 34066 28488 34342
rect 28448 34060 28500 34066
rect 28448 34002 28500 34008
rect 28920 33998 28948 34478
rect 28908 33992 28960 33998
rect 28908 33934 28960 33940
rect 28920 33454 28948 33934
rect 29092 33856 29144 33862
rect 29092 33798 29144 33804
rect 28356 33448 28408 33454
rect 28356 33390 28408 33396
rect 28540 33448 28592 33454
rect 28540 33390 28592 33396
rect 28908 33448 28960 33454
rect 28908 33390 28960 33396
rect 27160 33312 27212 33318
rect 27160 33254 27212 33260
rect 27172 32978 27200 33254
rect 27160 32972 27212 32978
rect 27160 32914 27212 32920
rect 27804 32768 27856 32774
rect 27804 32710 27856 32716
rect 27988 32768 28040 32774
rect 27988 32710 28040 32716
rect 26608 31816 26660 31822
rect 26608 31758 26660 31764
rect 27712 31816 27764 31822
rect 27712 31758 27764 31764
rect 26620 30938 26648 31758
rect 27252 31748 27304 31754
rect 27252 31690 27304 31696
rect 27264 31346 27292 31690
rect 27724 31482 27752 31758
rect 27712 31476 27764 31482
rect 27712 31418 27764 31424
rect 27252 31340 27304 31346
rect 27252 31282 27304 31288
rect 26884 31272 26936 31278
rect 26884 31214 26936 31220
rect 26976 31272 27028 31278
rect 26976 31214 27028 31220
rect 26608 30932 26660 30938
rect 26608 30874 26660 30880
rect 26700 30796 26752 30802
rect 26700 30738 26752 30744
rect 26712 30394 26740 30738
rect 26700 30388 26752 30394
rect 26700 30330 26752 30336
rect 26424 30116 26476 30122
rect 26424 30058 26476 30064
rect 26436 29646 26464 30058
rect 26424 29640 26476 29646
rect 26424 29582 26476 29588
rect 26896 29306 26924 31214
rect 26988 30054 27016 31214
rect 27724 30802 27752 31418
rect 27160 30796 27212 30802
rect 27160 30738 27212 30744
rect 27712 30796 27764 30802
rect 27712 30738 27764 30744
rect 27172 30190 27200 30738
rect 27160 30184 27212 30190
rect 27160 30126 27212 30132
rect 26976 30048 27028 30054
rect 26976 29990 27028 29996
rect 26424 29300 26476 29306
rect 26424 29242 26476 29248
rect 26884 29300 26936 29306
rect 26884 29242 26936 29248
rect 26436 28014 26464 29242
rect 27172 29102 27200 30126
rect 27436 30048 27488 30054
rect 27436 29990 27488 29996
rect 27448 29578 27476 29990
rect 27620 29640 27672 29646
rect 27620 29582 27672 29588
rect 27436 29572 27488 29578
rect 27436 29514 27488 29520
rect 27160 29096 27212 29102
rect 27160 29038 27212 29044
rect 26516 28620 26568 28626
rect 26516 28562 26568 28568
rect 26424 28008 26476 28014
rect 26424 27950 26476 27956
rect 26528 27402 26556 28562
rect 26884 28552 26936 28558
rect 26884 28494 26936 28500
rect 26976 28552 27028 28558
rect 26976 28494 27028 28500
rect 26896 28082 26924 28494
rect 26884 28076 26936 28082
rect 26884 28018 26936 28024
rect 26792 27532 26844 27538
rect 26988 27520 27016 28494
rect 26844 27492 27016 27520
rect 26792 27474 26844 27480
rect 26516 27396 26568 27402
rect 26516 27338 26568 27344
rect 26804 26450 26832 27474
rect 27172 27470 27200 29038
rect 27344 27872 27396 27878
rect 27448 27826 27476 29514
rect 27632 29102 27660 29582
rect 27620 29096 27672 29102
rect 27620 29038 27672 29044
rect 27396 27820 27476 27826
rect 27344 27814 27476 27820
rect 27356 27798 27476 27814
rect 27160 27464 27212 27470
rect 27160 27406 27212 27412
rect 27448 27402 27476 27798
rect 27528 27464 27580 27470
rect 27528 27406 27580 27412
rect 27436 27396 27488 27402
rect 27436 27338 27488 27344
rect 26792 26444 26844 26450
rect 26792 26386 26844 26392
rect 26424 25968 26476 25974
rect 26424 25910 26476 25916
rect 26436 25430 26464 25910
rect 26516 25832 26568 25838
rect 26516 25774 26568 25780
rect 26424 25424 26476 25430
rect 26424 25366 26476 25372
rect 26528 25226 26556 25774
rect 26516 25220 26568 25226
rect 26516 25162 26568 25168
rect 26528 23118 26556 25162
rect 26804 24206 26832 26386
rect 27448 25226 27476 27338
rect 27540 26926 27568 27406
rect 27528 26920 27580 26926
rect 27528 26862 27580 26868
rect 27620 26444 27672 26450
rect 27620 26386 27672 26392
rect 27632 25294 27660 26386
rect 27620 25288 27672 25294
rect 27620 25230 27672 25236
rect 27436 25220 27488 25226
rect 27436 25162 27488 25168
rect 27816 24954 27844 32710
rect 28000 31890 28028 32710
rect 28368 31890 28396 33390
rect 27988 31884 28040 31890
rect 27988 31826 28040 31832
rect 28356 31884 28408 31890
rect 28356 31826 28408 31832
rect 27988 30728 28040 30734
rect 27988 30670 28040 30676
rect 27896 30592 27948 30598
rect 27896 30534 27948 30540
rect 27908 28558 27936 30534
rect 28000 30326 28028 30670
rect 27988 30320 28040 30326
rect 27988 30262 28040 30268
rect 28080 29640 28132 29646
rect 28080 29582 28132 29588
rect 28092 29238 28120 29582
rect 28080 29232 28132 29238
rect 28080 29174 28132 29180
rect 27896 28552 27948 28558
rect 27896 28494 27948 28500
rect 28552 28490 28580 33390
rect 29104 33046 29132 33798
rect 29092 33040 29144 33046
rect 29092 32982 29144 32988
rect 28632 32972 28684 32978
rect 28632 32914 28684 32920
rect 28644 31278 28672 32914
rect 28632 31272 28684 31278
rect 28632 31214 28684 31220
rect 29000 30184 29052 30190
rect 29000 30126 29052 30132
rect 29012 28490 29040 30126
rect 28540 28484 28592 28490
rect 28540 28426 28592 28432
rect 29000 28484 29052 28490
rect 29000 28426 29052 28432
rect 28264 27940 28316 27946
rect 28264 27882 28316 27888
rect 28276 27538 28304 27882
rect 28264 27532 28316 27538
rect 28264 27474 28316 27480
rect 28448 27464 28500 27470
rect 28448 27406 28500 27412
rect 28460 27062 28488 27406
rect 28448 27056 28500 27062
rect 28448 26998 28500 27004
rect 28448 26920 28500 26926
rect 28448 26862 28500 26868
rect 29092 26920 29144 26926
rect 29092 26862 29144 26868
rect 27988 26784 28040 26790
rect 27988 26726 28040 26732
rect 28000 25906 28028 26726
rect 28460 26314 28488 26862
rect 29000 26512 29052 26518
rect 29000 26454 29052 26460
rect 28172 26308 28224 26314
rect 28172 26250 28224 26256
rect 28448 26308 28500 26314
rect 28448 26250 28500 26256
rect 27988 25900 28040 25906
rect 27988 25842 28040 25848
rect 28184 25362 28212 26250
rect 28172 25356 28224 25362
rect 28172 25298 28224 25304
rect 27804 24948 27856 24954
rect 27804 24890 27856 24896
rect 28264 24812 28316 24818
rect 28264 24754 28316 24760
rect 27712 24744 27764 24750
rect 27712 24686 27764 24692
rect 28080 24744 28132 24750
rect 28080 24686 28132 24692
rect 27436 24268 27488 24274
rect 27436 24210 27488 24216
rect 26792 24200 26844 24206
rect 26792 24142 26844 24148
rect 26700 24064 26752 24070
rect 26700 24006 26752 24012
rect 26712 23730 26740 24006
rect 26700 23724 26752 23730
rect 26700 23666 26752 23672
rect 26608 23588 26660 23594
rect 26608 23530 26660 23536
rect 26620 23186 26648 23530
rect 26608 23180 26660 23186
rect 26608 23122 26660 23128
rect 26712 23118 26740 23666
rect 26792 23656 26844 23662
rect 26792 23598 26844 23604
rect 26976 23656 27028 23662
rect 26976 23598 27028 23604
rect 26516 23112 26568 23118
rect 26700 23112 26752 23118
rect 26516 23054 26568 23060
rect 26620 23060 26700 23066
rect 26620 23054 26752 23060
rect 26528 21486 26556 23054
rect 26620 23038 26740 23054
rect 26516 21480 26568 21486
rect 26516 21422 26568 21428
rect 26514 19408 26570 19417
rect 26514 19343 26516 19352
rect 26568 19343 26570 19352
rect 26516 19314 26568 19320
rect 26620 18737 26648 23038
rect 26712 22989 26740 23038
rect 26700 22636 26752 22642
rect 26700 22578 26752 22584
rect 26606 18728 26662 18737
rect 26606 18663 26662 18672
rect 26516 17740 26568 17746
rect 26516 17682 26568 17688
rect 26528 17270 26556 17682
rect 26516 17264 26568 17270
rect 26516 17206 26568 17212
rect 26424 17196 26476 17202
rect 26424 17138 26476 17144
rect 26436 13410 26464 17138
rect 26712 17134 26740 22578
rect 26804 22234 26832 23598
rect 26884 22772 26936 22778
rect 26884 22714 26936 22720
rect 26896 22574 26924 22714
rect 26988 22642 27016 23598
rect 26976 22636 27028 22642
rect 26976 22578 27028 22584
rect 26884 22568 26936 22574
rect 26884 22510 26936 22516
rect 26792 22228 26844 22234
rect 26792 22170 26844 22176
rect 26804 20398 26832 22170
rect 26896 22098 26924 22510
rect 27344 22500 27396 22506
rect 27344 22442 27396 22448
rect 27356 22098 27384 22442
rect 26884 22092 26936 22098
rect 26884 22034 26936 22040
rect 27344 22092 27396 22098
rect 27344 22034 27396 22040
rect 26792 20392 26844 20398
rect 26792 20334 26844 20340
rect 26896 19310 26924 22034
rect 26976 22024 27028 22030
rect 26976 21966 27028 21972
rect 26988 21554 27016 21966
rect 26976 21548 27028 21554
rect 26976 21490 27028 21496
rect 27068 21480 27120 21486
rect 27068 21422 27120 21428
rect 26976 19916 27028 19922
rect 26976 19858 27028 19864
rect 26884 19304 26936 19310
rect 26884 19246 26936 19252
rect 26988 19174 27016 19858
rect 26976 19168 27028 19174
rect 26976 19110 27028 19116
rect 26974 18864 27030 18873
rect 26974 18799 27030 18808
rect 26988 18766 27016 18799
rect 26976 18760 27028 18766
rect 26976 18702 27028 18708
rect 27080 17814 27108 21422
rect 27252 21412 27304 21418
rect 27252 21354 27304 21360
rect 27264 21146 27292 21354
rect 27252 21140 27304 21146
rect 27252 21082 27304 21088
rect 27160 20460 27212 20466
rect 27160 20402 27212 20408
rect 27172 19514 27200 20402
rect 27264 19922 27292 21082
rect 27448 20602 27476 24210
rect 27724 23526 27752 24686
rect 28092 24410 28120 24686
rect 28080 24404 28132 24410
rect 28080 24346 28132 24352
rect 28276 24274 28304 24754
rect 29012 24614 29040 26454
rect 29104 24886 29132 26862
rect 29092 24880 29144 24886
rect 29092 24822 29144 24828
rect 29000 24608 29052 24614
rect 29000 24550 29052 24556
rect 28724 24404 28776 24410
rect 28724 24346 28776 24352
rect 28264 24268 28316 24274
rect 28264 24210 28316 24216
rect 27896 24064 27948 24070
rect 27896 24006 27948 24012
rect 27908 23662 27936 24006
rect 27896 23656 27948 23662
rect 27896 23598 27948 23604
rect 27712 23520 27764 23526
rect 27712 23462 27764 23468
rect 27712 23316 27764 23322
rect 27712 23258 27764 23264
rect 27620 23180 27672 23186
rect 27620 23122 27672 23128
rect 27528 22092 27580 22098
rect 27528 22034 27580 22040
rect 27540 21418 27568 22034
rect 27528 21412 27580 21418
rect 27528 21354 27580 21360
rect 27540 21010 27568 21354
rect 27528 21004 27580 21010
rect 27528 20946 27580 20952
rect 27436 20596 27488 20602
rect 27436 20538 27488 20544
rect 27448 20262 27476 20538
rect 27436 20256 27488 20262
rect 27436 20198 27488 20204
rect 27540 19990 27568 20946
rect 27528 19984 27580 19990
rect 27528 19926 27580 19932
rect 27252 19916 27304 19922
rect 27252 19858 27304 19864
rect 27160 19508 27212 19514
rect 27160 19450 27212 19456
rect 27172 18766 27200 19450
rect 27342 19408 27398 19417
rect 27342 19343 27398 19352
rect 27250 19272 27306 19281
rect 27250 19207 27252 19216
rect 27304 19207 27306 19216
rect 27252 19178 27304 19184
rect 27160 18760 27212 18766
rect 27160 18702 27212 18708
rect 27356 18426 27384 19343
rect 27528 19304 27580 19310
rect 27448 19264 27528 19292
rect 27448 19174 27476 19264
rect 27528 19246 27580 19252
rect 27436 19168 27488 19174
rect 27436 19110 27488 19116
rect 27252 18420 27304 18426
rect 27252 18362 27304 18368
rect 27344 18420 27396 18426
rect 27344 18362 27396 18368
rect 27264 18306 27292 18362
rect 27264 18290 27384 18306
rect 27264 18284 27396 18290
rect 27264 18278 27344 18284
rect 27344 18226 27396 18232
rect 27160 18216 27212 18222
rect 27448 18170 27476 19110
rect 27632 18873 27660 23122
rect 27724 19174 27752 23258
rect 27908 22642 27936 23598
rect 28276 23254 28304 24210
rect 28632 23656 28684 23662
rect 28632 23598 28684 23604
rect 28264 23248 28316 23254
rect 28264 23190 28316 23196
rect 28644 22642 28672 23598
rect 27896 22636 27948 22642
rect 27896 22578 27948 22584
rect 28632 22636 28684 22642
rect 28632 22578 28684 22584
rect 28172 22228 28224 22234
rect 28172 22170 28224 22176
rect 27988 22024 28040 22030
rect 27988 21966 28040 21972
rect 27804 20528 27856 20534
rect 27804 20470 27856 20476
rect 27816 19922 27844 20470
rect 27804 19916 27856 19922
rect 27804 19858 27856 19864
rect 27896 19304 27948 19310
rect 27896 19246 27948 19252
rect 27712 19168 27764 19174
rect 27908 19145 27936 19246
rect 27712 19110 27764 19116
rect 27894 19136 27950 19145
rect 27894 19071 27950 19080
rect 27618 18864 27674 18873
rect 27618 18799 27674 18808
rect 27528 18624 27580 18630
rect 27528 18566 27580 18572
rect 27540 18222 27568 18566
rect 27160 18158 27212 18164
rect 27172 18086 27200 18158
rect 27356 18142 27476 18170
rect 27528 18216 27580 18222
rect 27528 18158 27580 18164
rect 27160 18080 27212 18086
rect 27160 18022 27212 18028
rect 27068 17808 27120 17814
rect 27068 17750 27120 17756
rect 26516 17128 26568 17134
rect 26514 17096 26516 17105
rect 26700 17128 26752 17134
rect 26568 17096 26570 17105
rect 26700 17070 26752 17076
rect 26514 17031 26570 17040
rect 26516 16652 26568 16658
rect 26516 16594 26568 16600
rect 26528 14890 26556 16594
rect 26608 16448 26660 16454
rect 26608 16390 26660 16396
rect 26620 15570 26648 16390
rect 27356 16182 27384 18142
rect 27436 16992 27488 16998
rect 27436 16934 27488 16940
rect 27448 16250 27476 16934
rect 27436 16244 27488 16250
rect 27436 16186 27488 16192
rect 27068 16176 27120 16182
rect 27068 16118 27120 16124
rect 27344 16176 27396 16182
rect 27344 16118 27396 16124
rect 26792 15904 26844 15910
rect 26792 15846 26844 15852
rect 26608 15564 26660 15570
rect 26608 15506 26660 15512
rect 26620 15450 26648 15506
rect 26804 15502 26832 15846
rect 27080 15570 27108 16118
rect 27344 16040 27396 16046
rect 27344 15982 27396 15988
rect 27252 15904 27304 15910
rect 27252 15846 27304 15852
rect 27068 15564 27120 15570
rect 27068 15506 27120 15512
rect 26792 15496 26844 15502
rect 26620 15434 26740 15450
rect 26792 15438 26844 15444
rect 26620 15428 26752 15434
rect 26620 15422 26700 15428
rect 26700 15370 26752 15376
rect 26608 15360 26660 15366
rect 26608 15302 26660 15308
rect 26620 14958 26648 15302
rect 26712 14958 26740 15370
rect 26608 14952 26660 14958
rect 26608 14894 26660 14900
rect 26700 14952 26752 14958
rect 26700 14894 26752 14900
rect 26516 14884 26568 14890
rect 26516 14826 26568 14832
rect 27080 14618 27108 15506
rect 27068 14612 27120 14618
rect 27068 14554 27120 14560
rect 26792 14408 26844 14414
rect 26792 14350 26844 14356
rect 26804 14006 26832 14350
rect 27160 14340 27212 14346
rect 27160 14282 27212 14288
rect 26792 14000 26844 14006
rect 26792 13942 26844 13948
rect 27068 13864 27120 13870
rect 27068 13806 27120 13812
rect 26436 13382 26740 13410
rect 26424 12776 26476 12782
rect 26424 12718 26476 12724
rect 26436 11694 26464 12718
rect 26424 11688 26476 11694
rect 26424 11630 26476 11636
rect 26516 11076 26568 11082
rect 26516 11018 26568 11024
rect 26528 10606 26556 11018
rect 26516 10600 26568 10606
rect 26516 10542 26568 10548
rect 26332 10464 26384 10470
rect 26332 10406 26384 10412
rect 26240 9580 26292 9586
rect 26240 9522 26292 9528
rect 25964 9512 26016 9518
rect 25964 9454 26016 9460
rect 25976 8838 26004 9454
rect 25964 8832 26016 8838
rect 25964 8774 26016 8780
rect 26332 8424 26384 8430
rect 26332 8366 26384 8372
rect 26344 7342 26372 8366
rect 26332 7336 26384 7342
rect 26332 7278 26384 7284
rect 26240 5636 26292 5642
rect 26240 5578 26292 5584
rect 26252 4282 26280 5578
rect 26712 5386 26740 13382
rect 27080 13190 27108 13806
rect 27068 13184 27120 13190
rect 27068 13126 27120 13132
rect 26976 11688 27028 11694
rect 26976 11630 27028 11636
rect 26988 10130 27016 11630
rect 27172 11218 27200 14282
rect 27264 12782 27292 15846
rect 27356 15026 27384 15982
rect 27448 15706 27476 16186
rect 27540 16046 27568 18158
rect 27804 18080 27856 18086
rect 27804 18022 27856 18028
rect 27620 17740 27672 17746
rect 27620 17682 27672 17688
rect 27632 16658 27660 17682
rect 27816 16697 27844 18022
rect 27896 17536 27948 17542
rect 27896 17478 27948 17484
rect 27908 17338 27936 17478
rect 27896 17332 27948 17338
rect 27896 17274 27948 17280
rect 27802 16688 27858 16697
rect 27620 16652 27672 16658
rect 27802 16623 27804 16632
rect 27620 16594 27672 16600
rect 27856 16623 27858 16632
rect 27804 16594 27856 16600
rect 27528 16040 27580 16046
rect 27528 15982 27580 15988
rect 27436 15700 27488 15706
rect 27436 15642 27488 15648
rect 27344 15020 27396 15026
rect 27344 14962 27396 14968
rect 27356 14482 27384 14962
rect 27448 14958 27476 15642
rect 27528 15564 27580 15570
rect 27816 15552 27844 16594
rect 28000 16046 28028 21966
rect 28080 20800 28132 20806
rect 28080 20742 28132 20748
rect 28092 19922 28120 20742
rect 28184 20398 28212 22170
rect 28644 21690 28672 22578
rect 28632 21684 28684 21690
rect 28632 21626 28684 21632
rect 28172 20392 28224 20398
rect 28172 20334 28224 20340
rect 28448 20392 28500 20398
rect 28448 20334 28500 20340
rect 28080 19916 28132 19922
rect 28080 19858 28132 19864
rect 28460 19514 28488 20334
rect 28448 19508 28500 19514
rect 28448 19450 28500 19456
rect 28356 18760 28408 18766
rect 28356 18702 28408 18708
rect 28172 18284 28224 18290
rect 28172 18226 28224 18232
rect 28184 17134 28212 18226
rect 28368 17338 28396 18702
rect 28540 18624 28592 18630
rect 28540 18566 28592 18572
rect 28356 17332 28408 17338
rect 28356 17274 28408 17280
rect 28172 17128 28224 17134
rect 28264 17128 28316 17134
rect 28172 17070 28224 17076
rect 28262 17096 28264 17105
rect 28316 17096 28318 17105
rect 28262 17031 28318 17040
rect 28356 17060 28408 17066
rect 28356 17002 28408 17008
rect 28172 16584 28224 16590
rect 28172 16526 28224 16532
rect 27988 16040 28040 16046
rect 27988 15982 28040 15988
rect 27580 15524 27844 15552
rect 27528 15506 27580 15512
rect 27436 14952 27488 14958
rect 27436 14894 27488 14900
rect 27448 14550 27476 14894
rect 27896 14884 27948 14890
rect 27896 14826 27948 14832
rect 27528 14816 27580 14822
rect 27528 14758 27580 14764
rect 27620 14816 27672 14822
rect 27620 14758 27672 14764
rect 27436 14544 27488 14550
rect 27436 14486 27488 14492
rect 27344 14476 27396 14482
rect 27344 14418 27396 14424
rect 27540 13394 27568 14758
rect 27632 13462 27660 14758
rect 27620 13456 27672 13462
rect 27620 13398 27672 13404
rect 27344 13388 27396 13394
rect 27344 13330 27396 13336
rect 27528 13388 27580 13394
rect 27528 13330 27580 13336
rect 27356 12850 27384 13330
rect 27344 12844 27396 12850
rect 27344 12786 27396 12792
rect 27252 12776 27304 12782
rect 27252 12718 27304 12724
rect 27264 12442 27292 12718
rect 27632 12442 27660 13398
rect 27712 13320 27764 13326
rect 27712 13262 27764 13268
rect 27724 12714 27752 13262
rect 27804 13252 27856 13258
rect 27804 13194 27856 13200
rect 27712 12708 27764 12714
rect 27712 12650 27764 12656
rect 27252 12436 27304 12442
rect 27252 12378 27304 12384
rect 27620 12436 27672 12442
rect 27620 12378 27672 12384
rect 27620 12300 27672 12306
rect 27620 12242 27672 12248
rect 27252 12096 27304 12102
rect 27252 12038 27304 12044
rect 27264 11694 27292 12038
rect 27632 11762 27660 12242
rect 27724 11898 27752 12650
rect 27816 12238 27844 13194
rect 27908 12782 27936 14826
rect 28000 14482 28028 15982
rect 28184 15638 28212 16526
rect 28172 15632 28224 15638
rect 28172 15574 28224 15580
rect 28184 14958 28212 15574
rect 28368 15162 28396 17002
rect 28552 15978 28580 18566
rect 28632 17740 28684 17746
rect 28632 17682 28684 17688
rect 28540 15972 28592 15978
rect 28540 15914 28592 15920
rect 28552 15570 28580 15914
rect 28540 15564 28592 15570
rect 28540 15506 28592 15512
rect 28356 15156 28408 15162
rect 28356 15098 28408 15104
rect 28172 14952 28224 14958
rect 28172 14894 28224 14900
rect 27988 14476 28040 14482
rect 27988 14418 28040 14424
rect 28368 13530 28396 15098
rect 28356 13524 28408 13530
rect 28356 13466 28408 13472
rect 28172 13388 28224 13394
rect 28172 13330 28224 13336
rect 28184 12986 28212 13330
rect 28172 12980 28224 12986
rect 28172 12922 28224 12928
rect 28552 12782 28580 15506
rect 28644 15094 28672 17682
rect 28736 17252 28764 24346
rect 29000 24268 29052 24274
rect 29000 24210 29052 24216
rect 29012 24154 29040 24210
rect 28920 24126 29040 24154
rect 28920 21010 28948 24126
rect 29000 23316 29052 23322
rect 29000 23258 29052 23264
rect 29012 22030 29040 23258
rect 29000 22024 29052 22030
rect 29000 21966 29052 21972
rect 28908 21004 28960 21010
rect 28908 20946 28960 20952
rect 29012 19990 29040 21966
rect 29196 21434 29224 37266
rect 29368 36576 29420 36582
rect 29368 36518 29420 36524
rect 29380 35154 29408 36518
rect 29932 35834 29960 37318
rect 33140 37266 33192 37272
rect 30012 37256 30064 37262
rect 30012 37198 30064 37204
rect 30024 36786 30052 37198
rect 31024 37120 31076 37126
rect 31024 37062 31076 37068
rect 30012 36780 30064 36786
rect 30012 36722 30064 36728
rect 30288 36780 30340 36786
rect 30288 36722 30340 36728
rect 30104 36644 30156 36650
rect 30104 36586 30156 36592
rect 30012 36032 30064 36038
rect 30012 35974 30064 35980
rect 29920 35828 29972 35834
rect 29920 35770 29972 35776
rect 30024 35698 30052 35974
rect 30012 35692 30064 35698
rect 30012 35634 30064 35640
rect 30116 35154 30144 36586
rect 30300 35630 30328 36722
rect 30840 36712 30892 36718
rect 30840 36654 30892 36660
rect 30380 36032 30432 36038
rect 30380 35974 30432 35980
rect 30288 35624 30340 35630
rect 30288 35566 30340 35572
rect 30392 35154 30420 35974
rect 30656 35488 30708 35494
rect 30656 35430 30708 35436
rect 30668 35222 30696 35430
rect 30656 35216 30708 35222
rect 30656 35158 30708 35164
rect 29368 35148 29420 35154
rect 29368 35090 29420 35096
rect 30104 35148 30156 35154
rect 30104 35090 30156 35096
rect 30380 35148 30432 35154
rect 30380 35090 30432 35096
rect 29552 34536 29604 34542
rect 29552 34478 29604 34484
rect 29564 34202 29592 34478
rect 29552 34196 29604 34202
rect 29552 34138 29604 34144
rect 29276 34060 29328 34066
rect 29276 34002 29328 34008
rect 29288 32026 29316 34002
rect 29368 33380 29420 33386
rect 29368 33322 29420 33328
rect 29276 32020 29328 32026
rect 29276 31962 29328 31968
rect 29276 30592 29328 30598
rect 29276 30534 29328 30540
rect 29288 29714 29316 30534
rect 29380 30326 29408 33322
rect 29828 32972 29880 32978
rect 29828 32914 29880 32920
rect 29736 32428 29788 32434
rect 29736 32370 29788 32376
rect 29460 32360 29512 32366
rect 29460 32302 29512 32308
rect 29472 32026 29500 32302
rect 29748 32026 29776 32370
rect 29460 32020 29512 32026
rect 29460 31962 29512 31968
rect 29736 32020 29788 32026
rect 29736 31962 29788 31968
rect 29368 30320 29420 30326
rect 29368 30262 29420 30268
rect 29472 30190 29500 31962
rect 29840 30190 29868 32914
rect 29460 30184 29512 30190
rect 29460 30126 29512 30132
rect 29644 30184 29696 30190
rect 29644 30126 29696 30132
rect 29828 30184 29880 30190
rect 29828 30126 29880 30132
rect 29276 29708 29328 29714
rect 29276 29650 29328 29656
rect 29288 28626 29316 29650
rect 29656 29646 29684 30126
rect 29920 29844 29972 29850
rect 29920 29786 29972 29792
rect 29644 29640 29696 29646
rect 29644 29582 29696 29588
rect 29460 29096 29512 29102
rect 29460 29038 29512 29044
rect 29368 28688 29420 28694
rect 29368 28630 29420 28636
rect 29276 28620 29328 28626
rect 29276 28562 29328 28568
rect 29380 28014 29408 28630
rect 29368 28008 29420 28014
rect 29368 27950 29420 27956
rect 29276 26376 29328 26382
rect 29276 26318 29328 26324
rect 29288 25838 29316 26318
rect 29276 25832 29328 25838
rect 29276 25774 29328 25780
rect 29288 24750 29316 25774
rect 29276 24744 29328 24750
rect 29276 24686 29328 24692
rect 29368 24200 29420 24206
rect 29368 24142 29420 24148
rect 29380 23866 29408 24142
rect 29368 23860 29420 23866
rect 29368 23802 29420 23808
rect 29368 22092 29420 22098
rect 29368 22034 29420 22040
rect 29380 21486 29408 22034
rect 29368 21480 29420 21486
rect 29196 21406 29316 21434
rect 29368 21422 29420 21428
rect 29184 21344 29236 21350
rect 29184 21286 29236 21292
rect 29288 21298 29316 21406
rect 29196 21010 29224 21286
rect 29288 21270 29408 21298
rect 29276 21140 29328 21146
rect 29276 21082 29328 21088
rect 29288 21010 29316 21082
rect 29184 21004 29236 21010
rect 29184 20946 29236 20952
rect 29276 21004 29328 21010
rect 29276 20946 29328 20952
rect 29276 20392 29328 20398
rect 29276 20334 29328 20340
rect 29184 20052 29236 20058
rect 29184 19994 29236 20000
rect 29000 19984 29052 19990
rect 29000 19926 29052 19932
rect 29196 19514 29224 19994
rect 29184 19508 29236 19514
rect 29184 19450 29236 19456
rect 29000 19440 29052 19446
rect 29000 19382 29052 19388
rect 28908 19304 28960 19310
rect 28908 19246 28960 19252
rect 28920 18630 28948 19246
rect 29012 18834 29040 19382
rect 29092 19372 29144 19378
rect 29092 19314 29144 19320
rect 29000 18828 29052 18834
rect 29000 18770 29052 18776
rect 28908 18624 28960 18630
rect 28908 18566 28960 18572
rect 28816 17876 28868 17882
rect 28816 17818 28868 17824
rect 28828 17746 28856 17818
rect 28816 17740 28868 17746
rect 28816 17682 28868 17688
rect 29000 17672 29052 17678
rect 29000 17614 29052 17620
rect 29012 17338 29040 17614
rect 29000 17332 29052 17338
rect 29000 17274 29052 17280
rect 28736 17224 28948 17252
rect 28632 15088 28684 15094
rect 28632 15030 28684 15036
rect 28632 14612 28684 14618
rect 28632 14554 28684 14560
rect 28644 14074 28672 14554
rect 28724 14272 28776 14278
rect 28724 14214 28776 14220
rect 28632 14068 28684 14074
rect 28632 14010 28684 14016
rect 28736 13954 28764 14214
rect 28644 13926 28764 13954
rect 28644 13870 28672 13926
rect 28632 13864 28684 13870
rect 28632 13806 28684 13812
rect 27896 12776 27948 12782
rect 27896 12718 27948 12724
rect 28540 12776 28592 12782
rect 28540 12718 28592 12724
rect 27908 12306 27936 12718
rect 27988 12436 28040 12442
rect 27988 12378 28040 12384
rect 27896 12300 27948 12306
rect 27896 12242 27948 12248
rect 27804 12232 27856 12238
rect 27804 12174 27856 12180
rect 27712 11892 27764 11898
rect 27712 11834 27764 11840
rect 27620 11756 27672 11762
rect 27620 11698 27672 11704
rect 27252 11688 27304 11694
rect 27252 11630 27304 11636
rect 27632 11354 27660 11698
rect 27724 11694 27752 11834
rect 27712 11688 27764 11694
rect 27712 11630 27764 11636
rect 27724 11354 27752 11630
rect 27620 11348 27672 11354
rect 27620 11290 27672 11296
rect 27712 11348 27764 11354
rect 27712 11290 27764 11296
rect 27160 11212 27212 11218
rect 27160 11154 27212 11160
rect 27528 11008 27580 11014
rect 27528 10950 27580 10956
rect 27540 10742 27568 10950
rect 27724 10742 27752 11290
rect 27528 10736 27580 10742
rect 27528 10678 27580 10684
rect 27712 10736 27764 10742
rect 27712 10678 27764 10684
rect 27816 10674 27844 12174
rect 28000 11898 28028 12378
rect 28552 12374 28580 12718
rect 28540 12368 28592 12374
rect 28540 12310 28592 12316
rect 28172 12096 28224 12102
rect 28172 12038 28224 12044
rect 27988 11892 28040 11898
rect 27988 11834 28040 11840
rect 28000 10674 28028 11834
rect 28080 11076 28132 11082
rect 28080 11018 28132 11024
rect 27804 10668 27856 10674
rect 27804 10610 27856 10616
rect 27988 10668 28040 10674
rect 27988 10610 28040 10616
rect 28092 10554 28120 11018
rect 28184 10606 28212 12038
rect 28644 11218 28672 13806
rect 28816 13388 28868 13394
rect 28816 13330 28868 13336
rect 28724 13184 28776 13190
rect 28724 13126 28776 13132
rect 28736 12170 28764 13126
rect 28828 12306 28856 13330
rect 28816 12300 28868 12306
rect 28816 12242 28868 12248
rect 28724 12164 28776 12170
rect 28724 12106 28776 12112
rect 28632 11212 28684 11218
rect 28632 11154 28684 11160
rect 28920 10742 28948 17224
rect 28998 16688 29054 16697
rect 28998 16623 29054 16632
rect 29012 16590 29040 16623
rect 29000 16584 29052 16590
rect 29000 16526 29052 16532
rect 29012 15570 29040 16526
rect 29000 15564 29052 15570
rect 29000 15506 29052 15512
rect 29000 14476 29052 14482
rect 29000 14418 29052 14424
rect 29012 11558 29040 14418
rect 29104 12424 29132 19314
rect 29184 18352 29236 18358
rect 29184 18294 29236 18300
rect 29196 15978 29224 18294
rect 29288 18034 29316 20334
rect 29380 19394 29408 21270
rect 29472 20058 29500 29038
rect 29656 28626 29684 29582
rect 29932 29170 29960 29786
rect 29920 29164 29972 29170
rect 29920 29106 29972 29112
rect 29644 28620 29696 28626
rect 29644 28562 29696 28568
rect 29656 26586 29684 28562
rect 30116 27674 30144 35090
rect 30748 35012 30800 35018
rect 30748 34954 30800 34960
rect 30656 34400 30708 34406
rect 30656 34342 30708 34348
rect 30472 33856 30524 33862
rect 30472 33798 30524 33804
rect 30484 32366 30512 33798
rect 30668 33522 30696 34342
rect 30656 33516 30708 33522
rect 30656 33458 30708 33464
rect 30760 33454 30788 34954
rect 30748 33448 30800 33454
rect 30748 33390 30800 33396
rect 30564 32972 30616 32978
rect 30564 32914 30616 32920
rect 30576 32502 30604 32914
rect 30748 32836 30800 32842
rect 30748 32778 30800 32784
rect 30564 32496 30616 32502
rect 30564 32438 30616 32444
rect 30760 32434 30788 32778
rect 30748 32428 30800 32434
rect 30748 32370 30800 32376
rect 30288 32360 30340 32366
rect 30288 32302 30340 32308
rect 30472 32360 30524 32366
rect 30472 32302 30524 32308
rect 30300 31278 30328 32302
rect 30484 31278 30512 32302
rect 30656 31884 30708 31890
rect 30656 31826 30708 31832
rect 30288 31272 30340 31278
rect 30288 31214 30340 31220
rect 30472 31272 30524 31278
rect 30472 31214 30524 31220
rect 30196 31136 30248 31142
rect 30196 31078 30248 31084
rect 30208 28014 30236 31078
rect 30300 30802 30328 31214
rect 30484 30802 30512 31214
rect 30564 31204 30616 31210
rect 30564 31146 30616 31152
rect 30576 30870 30604 31146
rect 30564 30864 30616 30870
rect 30564 30806 30616 30812
rect 30288 30796 30340 30802
rect 30288 30738 30340 30744
rect 30472 30796 30524 30802
rect 30472 30738 30524 30744
rect 30300 29714 30328 30738
rect 30484 29714 30512 30738
rect 30668 30666 30696 31826
rect 30748 31748 30800 31754
rect 30748 31690 30800 31696
rect 30760 31346 30788 31690
rect 30748 31340 30800 31346
rect 30748 31282 30800 31288
rect 30656 30660 30708 30666
rect 30656 30602 30708 30608
rect 30288 29708 30340 29714
rect 30288 29650 30340 29656
rect 30472 29708 30524 29714
rect 30472 29650 30524 29656
rect 30484 29102 30512 29650
rect 30380 29096 30432 29102
rect 30380 29038 30432 29044
rect 30472 29096 30524 29102
rect 30472 29038 30524 29044
rect 30196 28008 30248 28014
rect 30196 27950 30248 27956
rect 30288 28008 30340 28014
rect 30288 27950 30340 27956
rect 30104 27668 30156 27674
rect 30104 27610 30156 27616
rect 29920 27328 29972 27334
rect 29920 27270 29972 27276
rect 29932 26926 29960 27270
rect 30300 27062 30328 27950
rect 30392 27538 30420 29038
rect 30656 28620 30708 28626
rect 30656 28562 30708 28568
rect 30564 28484 30616 28490
rect 30564 28426 30616 28432
rect 30576 28014 30604 28426
rect 30564 28008 30616 28014
rect 30564 27950 30616 27956
rect 30380 27532 30432 27538
rect 30380 27474 30432 27480
rect 30288 27056 30340 27062
rect 30288 26998 30340 27004
rect 29920 26920 29972 26926
rect 29920 26862 29972 26868
rect 29644 26580 29696 26586
rect 29644 26522 29696 26528
rect 29656 26450 29684 26522
rect 29932 26518 29960 26862
rect 29920 26512 29972 26518
rect 29920 26454 29972 26460
rect 29644 26444 29696 26450
rect 29644 26386 29696 26392
rect 30300 25906 30328 26998
rect 30392 26926 30420 27474
rect 30668 27402 30696 28562
rect 30656 27396 30708 27402
rect 30656 27338 30708 27344
rect 30380 26920 30432 26926
rect 30380 26862 30432 26868
rect 30748 26376 30800 26382
rect 30748 26318 30800 26324
rect 30656 26308 30708 26314
rect 30656 26250 30708 26256
rect 30668 25906 30696 26250
rect 30288 25900 30340 25906
rect 30288 25842 30340 25848
rect 30656 25900 30708 25906
rect 30656 25842 30708 25848
rect 29920 25424 29972 25430
rect 29920 25366 29972 25372
rect 29828 25288 29880 25294
rect 29828 25230 29880 25236
rect 29840 24750 29868 25230
rect 29828 24744 29880 24750
rect 29828 24686 29880 24692
rect 29932 23594 29960 25366
rect 30760 25362 30788 26318
rect 30564 25356 30616 25362
rect 30564 25298 30616 25304
rect 30748 25356 30800 25362
rect 30748 25298 30800 25304
rect 30472 24744 30524 24750
rect 30472 24686 30524 24692
rect 30484 24070 30512 24686
rect 30472 24064 30524 24070
rect 30472 24006 30524 24012
rect 30576 23662 30604 25298
rect 30852 25242 30880 36654
rect 31036 35222 31064 37062
rect 32956 36712 33008 36718
rect 32956 36654 33008 36660
rect 32968 36310 32996 36654
rect 32956 36304 33008 36310
rect 32956 36246 33008 36252
rect 33152 36242 33180 37266
rect 33508 37256 33560 37262
rect 33508 37198 33560 37204
rect 32312 36236 32364 36242
rect 32312 36178 32364 36184
rect 33140 36236 33192 36242
rect 33140 36178 33192 36184
rect 31116 35488 31168 35494
rect 31116 35430 31168 35436
rect 31024 35216 31076 35222
rect 31024 35158 31076 35164
rect 31024 35080 31076 35086
rect 31024 35022 31076 35028
rect 31036 33998 31064 35022
rect 31024 33992 31076 33998
rect 31024 33934 31076 33940
rect 31036 32366 31064 33934
rect 31024 32360 31076 32366
rect 31024 32302 31076 32308
rect 30932 32292 30984 32298
rect 30932 32234 30984 32240
rect 30944 31278 30972 32234
rect 30932 31272 30984 31278
rect 30932 31214 30984 31220
rect 30944 30394 30972 31214
rect 31036 30734 31064 32302
rect 31024 30728 31076 30734
rect 31024 30670 31076 30676
rect 30932 30388 30984 30394
rect 30932 30330 30984 30336
rect 30932 30184 30984 30190
rect 30932 30126 30984 30132
rect 30944 29170 30972 30126
rect 31024 29708 31076 29714
rect 31024 29650 31076 29656
rect 31036 29306 31064 29650
rect 31024 29300 31076 29306
rect 31024 29242 31076 29248
rect 30932 29164 30984 29170
rect 30932 29106 30984 29112
rect 31128 26874 31156 35430
rect 31852 35080 31904 35086
rect 31852 35022 31904 35028
rect 32220 35080 32272 35086
rect 32220 35022 32272 35028
rect 31392 34536 31444 34542
rect 31392 34478 31444 34484
rect 31668 34536 31720 34542
rect 31668 34478 31720 34484
rect 31404 33454 31432 34478
rect 31680 34134 31708 34478
rect 31668 34128 31720 34134
rect 31668 34070 31720 34076
rect 31864 33522 31892 35022
rect 32232 34202 32260 35022
rect 32324 34746 32352 36178
rect 33152 34746 33180 36178
rect 33520 36174 33548 37198
rect 33508 36168 33560 36174
rect 33508 36110 33560 36116
rect 33416 36100 33468 36106
rect 33416 36042 33468 36048
rect 33428 35154 33456 36042
rect 33416 35148 33468 35154
rect 33416 35090 33468 35096
rect 32312 34740 32364 34746
rect 32312 34682 32364 34688
rect 33140 34740 33192 34746
rect 33140 34682 33192 34688
rect 33520 34542 33548 36110
rect 34256 35766 34284 39200
rect 35900 37324 35952 37330
rect 35900 37266 35952 37272
rect 35532 37256 35584 37262
rect 35532 37198 35584 37204
rect 34940 37020 35236 37040
rect 34996 37018 35020 37020
rect 35076 37018 35100 37020
rect 35156 37018 35180 37020
rect 35018 36966 35020 37018
rect 35082 36966 35094 37018
rect 35156 36966 35158 37018
rect 34996 36964 35020 36966
rect 35076 36964 35100 36966
rect 35156 36964 35180 36966
rect 34940 36944 35236 36964
rect 35544 36718 35572 37198
rect 35532 36712 35584 36718
rect 35532 36654 35584 36660
rect 35348 36644 35400 36650
rect 35348 36586 35400 36592
rect 35360 36242 35388 36586
rect 35544 36242 35572 36654
rect 35912 36582 35940 37266
rect 35992 36848 36044 36854
rect 36280 36802 36308 39200
rect 38106 37632 38162 37641
rect 38106 37567 38162 37576
rect 36452 37392 36504 37398
rect 36452 37334 36504 37340
rect 35992 36790 36044 36796
rect 36004 36718 36032 36790
rect 36188 36786 36308 36802
rect 36176 36780 36308 36786
rect 36228 36774 36308 36780
rect 36176 36722 36228 36728
rect 35992 36712 36044 36718
rect 35992 36654 36044 36660
rect 35900 36576 35952 36582
rect 35900 36518 35952 36524
rect 34704 36236 34756 36242
rect 34704 36178 34756 36184
rect 35348 36236 35400 36242
rect 35348 36178 35400 36184
rect 35532 36236 35584 36242
rect 35532 36178 35584 36184
rect 35624 36236 35676 36242
rect 35624 36178 35676 36184
rect 34520 36100 34572 36106
rect 34520 36042 34572 36048
rect 34244 35760 34296 35766
rect 34244 35702 34296 35708
rect 33784 35624 33836 35630
rect 33784 35566 33836 35572
rect 34152 35624 34204 35630
rect 34152 35566 34204 35572
rect 33796 35290 33824 35566
rect 33784 35284 33836 35290
rect 33784 35226 33836 35232
rect 34164 35222 34192 35566
rect 34152 35216 34204 35222
rect 34152 35158 34204 35164
rect 34532 34610 34560 36042
rect 34716 35766 34744 36178
rect 34940 35932 35236 35952
rect 34996 35930 35020 35932
rect 35076 35930 35100 35932
rect 35156 35930 35180 35932
rect 35018 35878 35020 35930
rect 35082 35878 35094 35930
rect 35156 35878 35158 35930
rect 34996 35876 35020 35878
rect 35076 35876 35100 35878
rect 35156 35876 35180 35878
rect 34940 35856 35236 35876
rect 34704 35760 34756 35766
rect 34704 35702 34756 35708
rect 35544 35222 35572 36178
rect 35636 35630 35664 36178
rect 35912 36174 35940 36518
rect 35900 36168 35952 36174
rect 35900 36110 35952 36116
rect 35624 35624 35676 35630
rect 35624 35566 35676 35572
rect 35808 35488 35860 35494
rect 35808 35430 35860 35436
rect 35820 35222 35848 35430
rect 35912 35290 35940 36110
rect 36004 35698 36032 36654
rect 36084 36644 36136 36650
rect 36084 36586 36136 36592
rect 35992 35692 36044 35698
rect 35992 35634 36044 35640
rect 35900 35284 35952 35290
rect 35900 35226 35952 35232
rect 35532 35216 35584 35222
rect 35532 35158 35584 35164
rect 35808 35216 35860 35222
rect 35808 35158 35860 35164
rect 35256 35012 35308 35018
rect 35256 34954 35308 34960
rect 34940 34844 35236 34864
rect 34996 34842 35020 34844
rect 35076 34842 35100 34844
rect 35156 34842 35180 34844
rect 35018 34790 35020 34842
rect 35082 34790 35094 34842
rect 35156 34790 35158 34842
rect 34996 34788 35020 34790
rect 35076 34788 35100 34790
rect 35156 34788 35180 34790
rect 34940 34768 35236 34788
rect 34520 34604 34572 34610
rect 34520 34546 34572 34552
rect 33508 34536 33560 34542
rect 33508 34478 33560 34484
rect 35268 34354 35296 34954
rect 35440 34944 35492 34950
rect 35440 34886 35492 34892
rect 35452 34542 35480 34886
rect 35820 34678 35848 35158
rect 36096 35154 36124 36586
rect 36464 36174 36492 37334
rect 37004 37324 37056 37330
rect 37004 37266 37056 37272
rect 37188 37324 37240 37330
rect 37188 37266 37240 37272
rect 37016 37210 37044 37266
rect 36728 37188 36780 37194
rect 36728 37130 36780 37136
rect 36924 37182 37044 37210
rect 37096 37188 37148 37194
rect 36740 36242 36768 37130
rect 36728 36236 36780 36242
rect 36728 36178 36780 36184
rect 36452 36168 36504 36174
rect 36452 36110 36504 36116
rect 36084 35148 36136 35154
rect 36084 35090 36136 35096
rect 36924 35086 36952 37182
rect 37096 37130 37148 37136
rect 37004 37120 37056 37126
rect 37004 37062 37056 37068
rect 37016 36786 37044 37062
rect 37108 36854 37136 37130
rect 37200 36922 37228 37266
rect 37188 36916 37240 36922
rect 37188 36858 37240 36864
rect 37096 36848 37148 36854
rect 37096 36790 37148 36796
rect 37004 36780 37056 36786
rect 37004 36722 37056 36728
rect 37096 36032 37148 36038
rect 37096 35974 37148 35980
rect 37108 35698 37136 35974
rect 37096 35692 37148 35698
rect 37096 35634 37148 35640
rect 36912 35080 36964 35086
rect 36912 35022 36964 35028
rect 36360 34740 36412 34746
rect 36360 34682 36412 34688
rect 35808 34672 35860 34678
rect 35808 34614 35860 34620
rect 35440 34536 35492 34542
rect 35440 34478 35492 34484
rect 35268 34326 35480 34354
rect 32220 34196 32272 34202
rect 32220 34138 32272 34144
rect 31944 34060 31996 34066
rect 31944 34002 31996 34008
rect 33048 34060 33100 34066
rect 33048 34002 33100 34008
rect 31852 33516 31904 33522
rect 31852 33458 31904 33464
rect 31392 33448 31444 33454
rect 31220 33408 31392 33436
rect 31220 32366 31248 33408
rect 31392 33390 31444 33396
rect 31760 32904 31812 32910
rect 31760 32846 31812 32852
rect 31208 32360 31260 32366
rect 31208 32302 31260 32308
rect 31772 31822 31800 32846
rect 31760 31816 31812 31822
rect 31760 31758 31812 31764
rect 31392 30388 31444 30394
rect 31392 30330 31444 30336
rect 31404 29170 31432 30330
rect 31852 30184 31904 30190
rect 31852 30126 31904 30132
rect 31668 30048 31720 30054
rect 31668 29990 31720 29996
rect 31680 29170 31708 29990
rect 31864 29782 31892 30126
rect 31852 29776 31904 29782
rect 31852 29718 31904 29724
rect 31760 29640 31812 29646
rect 31760 29582 31812 29588
rect 31392 29164 31444 29170
rect 31392 29106 31444 29112
rect 31668 29164 31720 29170
rect 31668 29106 31720 29112
rect 31484 28552 31536 28558
rect 31484 28494 31536 28500
rect 31208 27532 31260 27538
rect 31208 27474 31260 27480
rect 30760 25214 30880 25242
rect 30944 26846 31156 26874
rect 30656 24608 30708 24614
rect 30656 24550 30708 24556
rect 30564 23656 30616 23662
rect 30564 23598 30616 23604
rect 29552 23588 29604 23594
rect 29552 23530 29604 23536
rect 29920 23588 29972 23594
rect 29920 23530 29972 23536
rect 30380 23588 30432 23594
rect 30380 23530 30432 23536
rect 29564 22574 29592 23530
rect 29644 23520 29696 23526
rect 29644 23462 29696 23468
rect 29552 22568 29604 22574
rect 29552 22510 29604 22516
rect 29564 22166 29592 22510
rect 29552 22160 29604 22166
rect 29552 22102 29604 22108
rect 29564 21146 29592 22102
rect 29656 21486 29684 23462
rect 30288 23180 30340 23186
rect 30288 23122 30340 23128
rect 29828 23112 29880 23118
rect 29828 23054 29880 23060
rect 30012 23112 30064 23118
rect 30012 23054 30064 23060
rect 29840 22681 29868 23054
rect 30024 22710 30052 23054
rect 30012 22704 30064 22710
rect 29826 22672 29882 22681
rect 30012 22646 30064 22652
rect 29826 22607 29882 22616
rect 30300 22574 30328 23122
rect 30392 23118 30420 23530
rect 30472 23316 30524 23322
rect 30472 23258 30524 23264
rect 30380 23112 30432 23118
rect 30380 23054 30432 23060
rect 30288 22568 30340 22574
rect 30288 22510 30340 22516
rect 30392 22234 30420 23054
rect 30380 22228 30432 22234
rect 30380 22170 30432 22176
rect 30380 21616 30432 21622
rect 30380 21558 30432 21564
rect 29644 21480 29696 21486
rect 29644 21422 29696 21428
rect 29920 21480 29972 21486
rect 29920 21422 29972 21428
rect 29552 21140 29604 21146
rect 29552 21082 29604 21088
rect 29656 20602 29684 21422
rect 29644 20596 29696 20602
rect 29644 20538 29696 20544
rect 29460 20052 29512 20058
rect 29460 19994 29512 20000
rect 29644 19916 29696 19922
rect 29644 19858 29696 19864
rect 29380 19378 29500 19394
rect 29656 19378 29684 19858
rect 29380 19372 29512 19378
rect 29380 19366 29460 19372
rect 29460 19314 29512 19320
rect 29644 19372 29696 19378
rect 29644 19314 29696 19320
rect 29368 19304 29420 19310
rect 29368 19246 29420 19252
rect 29380 18902 29408 19246
rect 29736 19168 29788 19174
rect 29736 19110 29788 19116
rect 29368 18896 29420 18902
rect 29368 18838 29420 18844
rect 29552 18760 29604 18766
rect 29552 18702 29604 18708
rect 29644 18760 29696 18766
rect 29644 18702 29696 18708
rect 29564 18358 29592 18702
rect 29552 18352 29604 18358
rect 29552 18294 29604 18300
rect 29288 18006 29408 18034
rect 29276 17876 29328 17882
rect 29276 17818 29328 17824
rect 29288 16454 29316 17818
rect 29380 17746 29408 18006
rect 29368 17740 29420 17746
rect 29368 17682 29420 17688
rect 29656 17134 29684 18702
rect 29748 18154 29776 19110
rect 29828 18216 29880 18222
rect 29828 18158 29880 18164
rect 29736 18148 29788 18154
rect 29736 18090 29788 18096
rect 29644 17128 29696 17134
rect 29644 17070 29696 17076
rect 29748 17082 29776 18090
rect 29840 17202 29868 18158
rect 29828 17196 29880 17202
rect 29828 17138 29880 17144
rect 29656 16658 29684 17070
rect 29748 17054 29868 17082
rect 29460 16652 29512 16658
rect 29644 16652 29696 16658
rect 29460 16594 29512 16600
rect 29564 16612 29644 16640
rect 29276 16448 29328 16454
rect 29276 16390 29328 16396
rect 29184 15972 29236 15978
rect 29184 15914 29236 15920
rect 29184 15088 29236 15094
rect 29184 15030 29236 15036
rect 29196 12646 29224 15030
rect 29288 14090 29316 16390
rect 29368 15904 29420 15910
rect 29368 15846 29420 15852
rect 29380 15570 29408 15846
rect 29472 15570 29500 16594
rect 29368 15564 29420 15570
rect 29368 15506 29420 15512
rect 29460 15564 29512 15570
rect 29460 15506 29512 15512
rect 29380 14958 29408 15506
rect 29368 14952 29420 14958
rect 29368 14894 29420 14900
rect 29564 14278 29592 16612
rect 29644 16594 29696 16600
rect 29736 16040 29788 16046
rect 29736 15982 29788 15988
rect 29748 15706 29776 15982
rect 29736 15700 29788 15706
rect 29736 15642 29788 15648
rect 29840 14940 29868 17054
rect 29932 15094 29960 21422
rect 30196 21004 30248 21010
rect 30196 20946 30248 20952
rect 30208 20874 30236 20946
rect 30196 20868 30248 20874
rect 30196 20810 30248 20816
rect 30012 20392 30064 20398
rect 30012 20334 30064 20340
rect 30024 19446 30052 20334
rect 30104 20324 30156 20330
rect 30104 20266 30156 20272
rect 30116 19922 30144 20266
rect 30104 19916 30156 19922
rect 30104 19858 30156 19864
rect 30012 19440 30064 19446
rect 30012 19382 30064 19388
rect 30024 15994 30052 19382
rect 30208 19174 30236 20810
rect 30392 20262 30420 21558
rect 30484 21418 30512 23258
rect 30576 21690 30604 23598
rect 30668 22098 30696 24550
rect 30656 22092 30708 22098
rect 30656 22034 30708 22040
rect 30564 21684 30616 21690
rect 30564 21626 30616 21632
rect 30562 21584 30618 21593
rect 30562 21519 30618 21528
rect 30472 21412 30524 21418
rect 30472 21354 30524 21360
rect 30380 20256 30432 20262
rect 30380 20198 30432 20204
rect 30392 20058 30420 20198
rect 30380 20052 30432 20058
rect 30380 19994 30432 20000
rect 30472 19780 30524 19786
rect 30472 19722 30524 19728
rect 30380 19372 30432 19378
rect 30380 19314 30432 19320
rect 30288 19236 30340 19242
rect 30288 19178 30340 19184
rect 30196 19168 30248 19174
rect 30196 19110 30248 19116
rect 30196 18828 30248 18834
rect 30116 18788 30196 18816
rect 30116 17882 30144 18788
rect 30196 18770 30248 18776
rect 30300 18698 30328 19178
rect 30288 18692 30340 18698
rect 30288 18634 30340 18640
rect 30392 18358 30420 19314
rect 30380 18352 30432 18358
rect 30380 18294 30432 18300
rect 30196 18216 30248 18222
rect 30196 18158 30248 18164
rect 30104 17876 30156 17882
rect 30104 17818 30156 17824
rect 30104 17128 30156 17134
rect 30104 17070 30156 17076
rect 30116 16726 30144 17070
rect 30104 16720 30156 16726
rect 30104 16662 30156 16668
rect 30208 16182 30236 18158
rect 30484 17746 30512 19722
rect 30472 17740 30524 17746
rect 30472 17682 30524 17688
rect 30380 17536 30432 17542
rect 30380 17478 30432 17484
rect 30196 16176 30248 16182
rect 30196 16118 30248 16124
rect 30196 16040 30248 16046
rect 30024 15988 30196 15994
rect 30392 16017 30420 17478
rect 30484 17116 30512 17682
rect 30576 17542 30604 21519
rect 30668 20806 30696 22034
rect 30656 20800 30708 20806
rect 30656 20742 30708 20748
rect 30656 19712 30708 19718
rect 30656 19654 30708 19660
rect 30564 17536 30616 17542
rect 30564 17478 30616 17484
rect 30668 17270 30696 19654
rect 30760 18884 30788 25214
rect 30840 22568 30892 22574
rect 30840 22510 30892 22516
rect 30852 22098 30880 22510
rect 30840 22092 30892 22098
rect 30840 22034 30892 22040
rect 30852 21468 30880 22034
rect 30944 21593 30972 26846
rect 31116 26784 31168 26790
rect 31220 26772 31248 27474
rect 31168 26744 31248 26772
rect 31116 26726 31168 26732
rect 31024 26444 31076 26450
rect 31024 26386 31076 26392
rect 31036 23730 31064 26386
rect 31128 25702 31156 26726
rect 31496 26382 31524 28494
rect 31484 26376 31536 26382
rect 31536 26336 31616 26364
rect 31484 26318 31536 26324
rect 31116 25696 31168 25702
rect 31116 25638 31168 25644
rect 31024 23724 31076 23730
rect 31024 23666 31076 23672
rect 30930 21584 30986 21593
rect 30930 21519 30986 21528
rect 30932 21480 30984 21486
rect 30852 21440 30932 21468
rect 30932 21422 30984 21428
rect 30944 20602 30972 21422
rect 30932 20596 30984 20602
rect 30932 20538 30984 20544
rect 31036 20040 31064 23666
rect 31128 23118 31156 25638
rect 31208 25288 31260 25294
rect 31208 25230 31260 25236
rect 31220 24274 31248 25230
rect 31392 24744 31444 24750
rect 31392 24686 31444 24692
rect 31208 24268 31260 24274
rect 31208 24210 31260 24216
rect 31220 23662 31248 24210
rect 31208 23656 31260 23662
rect 31208 23598 31260 23604
rect 31220 23254 31248 23598
rect 31404 23322 31432 24686
rect 31484 24608 31536 24614
rect 31484 24550 31536 24556
rect 31496 23730 31524 24550
rect 31588 24138 31616 26336
rect 31772 25906 31800 29582
rect 31956 28218 31984 34002
rect 33060 33658 33088 34002
rect 33692 33992 33744 33998
rect 33692 33934 33744 33940
rect 33048 33652 33100 33658
rect 33048 33594 33100 33600
rect 33232 32972 33284 32978
rect 33232 32914 33284 32920
rect 33600 32972 33652 32978
rect 33600 32914 33652 32920
rect 32772 32904 32824 32910
rect 32772 32846 32824 32852
rect 32784 32570 32812 32846
rect 32772 32564 32824 32570
rect 32772 32506 32824 32512
rect 32784 31890 32812 32506
rect 32496 31884 32548 31890
rect 32496 31826 32548 31832
rect 32772 31884 32824 31890
rect 32772 31826 32824 31832
rect 32036 31816 32088 31822
rect 32036 31758 32088 31764
rect 32048 30666 32076 31758
rect 32508 31414 32536 31826
rect 32496 31408 32548 31414
rect 32496 31350 32548 31356
rect 33244 31278 33272 32914
rect 33612 32570 33640 32914
rect 33600 32564 33652 32570
rect 33600 32506 33652 32512
rect 33416 32292 33468 32298
rect 33416 32234 33468 32240
rect 33428 31958 33456 32234
rect 33416 31952 33468 31958
rect 33416 31894 33468 31900
rect 33232 31272 33284 31278
rect 33232 31214 33284 31220
rect 32772 31136 32824 31142
rect 32772 31078 32824 31084
rect 32784 30802 32812 31078
rect 32772 30796 32824 30802
rect 32772 30738 32824 30744
rect 33140 30728 33192 30734
rect 33140 30670 33192 30676
rect 32036 30660 32088 30666
rect 32036 30602 32088 30608
rect 32048 30190 32076 30602
rect 33152 30258 33180 30670
rect 33140 30252 33192 30258
rect 33140 30194 33192 30200
rect 33428 30190 33456 31894
rect 33600 31884 33652 31890
rect 33704 31872 33732 33934
rect 35348 33856 35400 33862
rect 35348 33798 35400 33804
rect 34940 33756 35236 33776
rect 34996 33754 35020 33756
rect 35076 33754 35100 33756
rect 35156 33754 35180 33756
rect 35018 33702 35020 33754
rect 35082 33702 35094 33754
rect 35156 33702 35158 33754
rect 34996 33700 35020 33702
rect 35076 33700 35100 33702
rect 35156 33700 35180 33702
rect 34940 33680 35236 33700
rect 35360 32978 35388 33798
rect 35452 33266 35480 34326
rect 35532 34060 35584 34066
rect 35532 34002 35584 34008
rect 35544 33454 35572 34002
rect 36176 33992 36228 33998
rect 36176 33934 36228 33940
rect 35532 33448 35584 33454
rect 35532 33390 35584 33396
rect 35452 33238 35572 33266
rect 35348 32972 35400 32978
rect 35348 32914 35400 32920
rect 34796 32904 34848 32910
rect 34796 32846 34848 32852
rect 34808 32434 34836 32846
rect 35440 32836 35492 32842
rect 35440 32778 35492 32784
rect 34940 32668 35236 32688
rect 34996 32666 35020 32668
rect 35076 32666 35100 32668
rect 35156 32666 35180 32668
rect 35018 32614 35020 32666
rect 35082 32614 35094 32666
rect 35156 32614 35158 32666
rect 34996 32612 35020 32614
rect 35076 32612 35100 32614
rect 35156 32612 35180 32614
rect 34940 32592 35236 32612
rect 34796 32428 34848 32434
rect 34796 32370 34848 32376
rect 34888 32360 34940 32366
rect 34888 32302 34940 32308
rect 35256 32360 35308 32366
rect 35256 32302 35308 32308
rect 34900 32026 34928 32302
rect 34888 32020 34940 32026
rect 34888 31962 34940 31968
rect 33652 31844 33732 31872
rect 33968 31884 34020 31890
rect 33600 31826 33652 31832
rect 33968 31826 34020 31832
rect 33612 30852 33640 31826
rect 33876 31816 33928 31822
rect 33876 31758 33928 31764
rect 33888 30938 33916 31758
rect 33980 31278 34008 31826
rect 34900 31770 34928 31962
rect 34808 31742 34928 31770
rect 34244 31340 34296 31346
rect 34244 31282 34296 31288
rect 33968 31272 34020 31278
rect 33968 31214 34020 31220
rect 33876 30932 33928 30938
rect 33876 30874 33928 30880
rect 33692 30864 33744 30870
rect 33612 30824 33692 30852
rect 33612 30394 33640 30824
rect 33692 30806 33744 30812
rect 34256 30802 34284 31282
rect 34808 31278 34836 31742
rect 34940 31580 35236 31600
rect 34996 31578 35020 31580
rect 35076 31578 35100 31580
rect 35156 31578 35180 31580
rect 35018 31526 35020 31578
rect 35082 31526 35094 31578
rect 35156 31526 35158 31578
rect 34996 31524 35020 31526
rect 35076 31524 35100 31526
rect 35156 31524 35180 31526
rect 34940 31504 35236 31524
rect 34796 31272 34848 31278
rect 34796 31214 34848 31220
rect 35268 30870 35296 32302
rect 35452 31362 35480 32778
rect 35544 31657 35572 33238
rect 35716 32904 35768 32910
rect 35716 32846 35768 32852
rect 35624 32768 35676 32774
rect 35624 32710 35676 32716
rect 35530 31648 35586 31657
rect 35530 31583 35586 31592
rect 35452 31334 35572 31362
rect 35348 31272 35400 31278
rect 35348 31214 35400 31220
rect 35256 30864 35308 30870
rect 35256 30806 35308 30812
rect 34244 30796 34296 30802
rect 34244 30738 34296 30744
rect 34940 30492 35236 30512
rect 34996 30490 35020 30492
rect 35076 30490 35100 30492
rect 35156 30490 35180 30492
rect 35018 30438 35020 30490
rect 35082 30438 35094 30490
rect 35156 30438 35158 30490
rect 34996 30436 35020 30438
rect 35076 30436 35100 30438
rect 35156 30436 35180 30438
rect 34940 30416 35236 30436
rect 33600 30388 33652 30394
rect 33600 30330 33652 30336
rect 32036 30184 32088 30190
rect 32036 30126 32088 30132
rect 32956 30184 33008 30190
rect 32956 30126 33008 30132
rect 33416 30184 33468 30190
rect 33416 30126 33468 30132
rect 32048 28490 32076 30126
rect 32772 30048 32824 30054
rect 32772 29990 32824 29996
rect 32784 29850 32812 29990
rect 32772 29844 32824 29850
rect 32772 29786 32824 29792
rect 32864 29708 32916 29714
rect 32864 29650 32916 29656
rect 32772 29572 32824 29578
rect 32772 29514 32824 29520
rect 32586 28792 32642 28801
rect 32312 28756 32364 28762
rect 32586 28727 32642 28736
rect 32312 28698 32364 28704
rect 32036 28484 32088 28490
rect 32036 28426 32088 28432
rect 31944 28212 31996 28218
rect 31944 28154 31996 28160
rect 32048 27130 32076 28426
rect 32324 28218 32352 28698
rect 32404 28620 32456 28626
rect 32404 28562 32456 28568
rect 32312 28212 32364 28218
rect 32312 28154 32364 28160
rect 32036 27124 32088 27130
rect 32036 27066 32088 27072
rect 32324 27010 32352 28154
rect 32416 28150 32444 28562
rect 32404 28144 32456 28150
rect 32404 28086 32456 28092
rect 32496 27464 32548 27470
rect 32496 27406 32548 27412
rect 32324 26982 32444 27010
rect 32312 26920 32364 26926
rect 32312 26862 32364 26868
rect 32220 26852 32272 26858
rect 32220 26794 32272 26800
rect 32232 26450 32260 26794
rect 32036 26444 32088 26450
rect 32036 26386 32088 26392
rect 32220 26444 32272 26450
rect 32220 26386 32272 26392
rect 32048 26042 32076 26386
rect 32036 26036 32088 26042
rect 32036 25978 32088 25984
rect 31760 25900 31812 25906
rect 31760 25842 31812 25848
rect 31944 25152 31996 25158
rect 31944 25094 31996 25100
rect 31956 24818 31984 25094
rect 31944 24812 31996 24818
rect 31944 24754 31996 24760
rect 31576 24132 31628 24138
rect 31576 24074 31628 24080
rect 31484 23724 31536 23730
rect 31484 23666 31536 23672
rect 31392 23316 31444 23322
rect 31392 23258 31444 23264
rect 31208 23248 31260 23254
rect 31208 23190 31260 23196
rect 31404 23202 31432 23258
rect 31116 23112 31168 23118
rect 31116 23054 31168 23060
rect 31220 22642 31248 23190
rect 31300 23180 31352 23186
rect 31404 23174 31524 23202
rect 31300 23122 31352 23128
rect 31208 22636 31260 22642
rect 31208 22578 31260 22584
rect 31208 22092 31260 22098
rect 31208 22034 31260 22040
rect 31220 21554 31248 22034
rect 31312 21622 31340 23122
rect 31392 23112 31444 23118
rect 31392 23054 31444 23060
rect 31300 21616 31352 21622
rect 31300 21558 31352 21564
rect 31208 21548 31260 21554
rect 31208 21490 31260 21496
rect 30944 20012 31064 20040
rect 30760 18856 30880 18884
rect 30748 17672 30800 17678
rect 30748 17614 30800 17620
rect 30656 17264 30708 17270
rect 30656 17206 30708 17212
rect 30564 17128 30616 17134
rect 30484 17088 30564 17116
rect 30564 17070 30616 17076
rect 30668 17066 30696 17206
rect 30656 17060 30708 17066
rect 30656 17002 30708 17008
rect 30760 16250 30788 17614
rect 30852 16794 30880 18856
rect 30840 16788 30892 16794
rect 30840 16730 30892 16736
rect 30748 16244 30800 16250
rect 30748 16186 30800 16192
rect 30024 15982 30248 15988
rect 30378 16008 30434 16017
rect 30024 15966 30236 15982
rect 30012 15496 30064 15502
rect 30012 15438 30064 15444
rect 29920 15088 29972 15094
rect 29920 15030 29972 15036
rect 29840 14912 29960 14940
rect 29644 14476 29696 14482
rect 29644 14418 29696 14424
rect 29552 14272 29604 14278
rect 29552 14214 29604 14220
rect 29288 14062 29592 14090
rect 29656 14074 29684 14418
rect 29460 12708 29512 12714
rect 29460 12650 29512 12656
rect 29184 12640 29236 12646
rect 29184 12582 29236 12588
rect 29368 12640 29420 12646
rect 29368 12582 29420 12588
rect 29104 12396 29316 12424
rect 29092 12300 29144 12306
rect 29092 12242 29144 12248
rect 29000 11552 29052 11558
rect 29000 11494 29052 11500
rect 29104 11150 29132 12242
rect 29184 11688 29236 11694
rect 29182 11656 29184 11665
rect 29236 11656 29238 11665
rect 29182 11591 29238 11600
rect 29182 11248 29238 11257
rect 29182 11183 29184 11192
rect 29236 11183 29238 11192
rect 29184 11154 29236 11160
rect 29092 11144 29144 11150
rect 29092 11086 29144 11092
rect 28540 10736 28592 10742
rect 28540 10678 28592 10684
rect 28908 10736 28960 10742
rect 28908 10678 28960 10684
rect 28000 10538 28120 10554
rect 28172 10600 28224 10606
rect 28172 10542 28224 10548
rect 27068 10532 27120 10538
rect 27068 10474 27120 10480
rect 27160 10532 27212 10538
rect 27160 10474 27212 10480
rect 27528 10532 27580 10538
rect 27528 10474 27580 10480
rect 27988 10532 28120 10538
rect 28040 10526 28120 10532
rect 27988 10474 28040 10480
rect 27080 10198 27108 10474
rect 27068 10192 27120 10198
rect 27068 10134 27120 10140
rect 26976 10124 27028 10130
rect 26976 10066 27028 10072
rect 26884 9444 26936 9450
rect 26884 9386 26936 9392
rect 26896 9042 26924 9386
rect 27080 9178 27108 10134
rect 27172 9926 27200 10474
rect 27344 10056 27396 10062
rect 27344 9998 27396 10004
rect 27160 9920 27212 9926
rect 27160 9862 27212 9868
rect 27356 9518 27384 9998
rect 27344 9512 27396 9518
rect 27344 9454 27396 9460
rect 27068 9172 27120 9178
rect 27068 9114 27120 9120
rect 27540 9042 27568 10474
rect 27620 10464 27672 10470
rect 27620 10406 27672 10412
rect 26884 9036 26936 9042
rect 26884 8978 26936 8984
rect 27528 9036 27580 9042
rect 27528 8978 27580 8984
rect 26976 8900 27028 8906
rect 26976 8842 27028 8848
rect 26792 8492 26844 8498
rect 26792 8434 26844 8440
rect 26804 5846 26832 8434
rect 26988 8022 27016 8842
rect 27068 8424 27120 8430
rect 27068 8366 27120 8372
rect 27252 8424 27304 8430
rect 27252 8366 27304 8372
rect 27344 8424 27396 8430
rect 27344 8366 27396 8372
rect 27080 8090 27108 8366
rect 27068 8084 27120 8090
rect 27068 8026 27120 8032
rect 26976 8016 27028 8022
rect 26976 7958 27028 7964
rect 26884 7404 26936 7410
rect 26884 7346 26936 7352
rect 26896 5846 26924 7346
rect 26988 7342 27016 7958
rect 27264 7954 27292 8366
rect 27252 7948 27304 7954
rect 27252 7890 27304 7896
rect 27160 7880 27212 7886
rect 27356 7834 27384 8366
rect 27436 7948 27488 7954
rect 27632 7936 27660 10406
rect 28000 10130 28028 10474
rect 27896 10124 27948 10130
rect 27896 10066 27948 10072
rect 27988 10124 28040 10130
rect 27988 10066 28040 10072
rect 27804 10056 27856 10062
rect 27804 9998 27856 10004
rect 27816 9042 27844 9998
rect 27804 9036 27856 9042
rect 27804 8978 27856 8984
rect 27908 8906 27936 10066
rect 27988 9988 28040 9994
rect 27988 9930 28040 9936
rect 28000 9450 28028 9930
rect 27988 9444 28040 9450
rect 27988 9386 28040 9392
rect 28184 9382 28212 10542
rect 28448 10464 28500 10470
rect 28448 10406 28500 10412
rect 28356 10124 28408 10130
rect 28356 10066 28408 10072
rect 28172 9376 28224 9382
rect 28172 9318 28224 9324
rect 28368 9178 28396 10066
rect 28460 9926 28488 10406
rect 28448 9920 28500 9926
rect 28448 9862 28500 9868
rect 28446 9616 28502 9625
rect 28446 9551 28502 9560
rect 28460 9518 28488 9551
rect 28448 9512 28500 9518
rect 28448 9454 28500 9460
rect 28356 9172 28408 9178
rect 28356 9114 28408 9120
rect 28172 8968 28224 8974
rect 28172 8910 28224 8916
rect 27896 8900 27948 8906
rect 27896 8842 27948 8848
rect 27896 8424 27948 8430
rect 27896 8366 27948 8372
rect 27488 7908 27660 7936
rect 27436 7890 27488 7896
rect 27160 7822 27212 7828
rect 26976 7336 27028 7342
rect 26976 7278 27028 7284
rect 27068 6792 27120 6798
rect 27068 6734 27120 6740
rect 27080 5914 27108 6734
rect 27068 5908 27120 5914
rect 27068 5850 27120 5856
rect 27172 5846 27200 7822
rect 27264 7818 27384 7834
rect 27252 7812 27384 7818
rect 27304 7806 27384 7812
rect 27252 7754 27304 7760
rect 27264 7342 27292 7754
rect 27344 7744 27396 7750
rect 27344 7686 27396 7692
rect 27356 7410 27384 7686
rect 27448 7546 27476 7890
rect 27436 7540 27488 7546
rect 27436 7482 27488 7488
rect 27344 7404 27396 7410
rect 27344 7346 27396 7352
rect 27252 7336 27304 7342
rect 27252 7278 27304 7284
rect 26792 5840 26844 5846
rect 26792 5782 26844 5788
rect 26884 5840 26936 5846
rect 26884 5782 26936 5788
rect 27160 5840 27212 5846
rect 27160 5782 27212 5788
rect 26712 5370 26924 5386
rect 26712 5364 26936 5370
rect 26712 5358 26884 5364
rect 26884 5306 26936 5312
rect 26792 5228 26844 5234
rect 26792 5170 26844 5176
rect 26804 4690 26832 5170
rect 26792 4684 26844 4690
rect 26792 4626 26844 4632
rect 26240 4276 26292 4282
rect 26240 4218 26292 4224
rect 26896 4078 26924 5306
rect 27160 5092 27212 5098
rect 27160 5034 27212 5040
rect 26884 4072 26936 4078
rect 26884 4014 26936 4020
rect 26516 4004 26568 4010
rect 26516 3946 26568 3952
rect 26528 3602 26556 3946
rect 27172 3602 27200 5034
rect 27264 3738 27292 7278
rect 27356 6866 27384 7346
rect 27908 7342 27936 8366
rect 27988 8356 28040 8362
rect 27988 8298 28040 8304
rect 28000 7954 28028 8298
rect 27988 7948 28040 7954
rect 27988 7890 28040 7896
rect 27896 7336 27948 7342
rect 27896 7278 27948 7284
rect 27528 7268 27580 7274
rect 27528 7210 27580 7216
rect 27344 6860 27396 6866
rect 27344 6802 27396 6808
rect 27436 6792 27488 6798
rect 27436 6734 27488 6740
rect 27448 6458 27476 6734
rect 27436 6452 27488 6458
rect 27436 6394 27488 6400
rect 27436 5772 27488 5778
rect 27540 5760 27568 7210
rect 27896 6860 27948 6866
rect 27896 6802 27948 6808
rect 27908 6254 27936 6802
rect 28184 6798 28212 8910
rect 28264 7336 28316 7342
rect 28264 7278 28316 7284
rect 28172 6792 28224 6798
rect 28172 6734 28224 6740
rect 27896 6248 27948 6254
rect 27896 6190 27948 6196
rect 27988 6248 28040 6254
rect 27988 6190 28040 6196
rect 27712 6180 27764 6186
rect 27712 6122 27764 6128
rect 27804 6180 27856 6186
rect 27804 6122 27856 6128
rect 27724 5914 27752 6122
rect 27712 5908 27764 5914
rect 27712 5850 27764 5856
rect 27816 5846 27844 6122
rect 27804 5840 27856 5846
rect 27804 5782 27856 5788
rect 27488 5732 27568 5760
rect 27436 5714 27488 5720
rect 27252 3732 27304 3738
rect 27252 3674 27304 3680
rect 26516 3596 26568 3602
rect 26516 3538 26568 3544
rect 27160 3596 27212 3602
rect 27160 3538 27212 3544
rect 25872 3052 25924 3058
rect 25872 2994 25924 3000
rect 26884 3052 26936 3058
rect 26884 2994 26936 3000
rect 26240 2984 26292 2990
rect 26240 2926 26292 2932
rect 26252 2650 26280 2926
rect 26240 2644 26292 2650
rect 26240 2586 26292 2592
rect 24124 2508 24176 2514
rect 24124 2450 24176 2456
rect 24860 2508 24912 2514
rect 24860 2450 24912 2456
rect 26896 2446 26924 2994
rect 27540 2922 27568 5732
rect 27908 2990 27936 6190
rect 28000 5846 28028 6190
rect 27988 5840 28040 5846
rect 27988 5782 28040 5788
rect 28172 5024 28224 5030
rect 28276 5012 28304 7278
rect 28552 6338 28580 10678
rect 28816 10532 28868 10538
rect 28816 10474 28868 10480
rect 28828 10198 28856 10474
rect 28816 10192 28868 10198
rect 28816 10134 28868 10140
rect 29196 10130 29224 11154
rect 29288 10577 29316 12396
rect 29274 10568 29330 10577
rect 29274 10503 29330 10512
rect 29000 10124 29052 10130
rect 29000 10066 29052 10072
rect 29184 10124 29236 10130
rect 29184 10066 29236 10072
rect 29012 9926 29040 10066
rect 29000 9920 29052 9926
rect 29000 9862 29052 9868
rect 28816 9172 28868 9178
rect 28816 9114 28868 9120
rect 28724 8968 28776 8974
rect 28724 8910 28776 8916
rect 28736 8566 28764 8910
rect 28724 8560 28776 8566
rect 28724 8502 28776 8508
rect 28552 6310 28672 6338
rect 28540 6248 28592 6254
rect 28540 6190 28592 6196
rect 28552 5846 28580 6190
rect 28540 5840 28592 5846
rect 28540 5782 28592 5788
rect 28644 5681 28672 6310
rect 28828 5778 28856 9114
rect 29012 9058 29040 9862
rect 29276 9648 29328 9654
rect 29276 9590 29328 9596
rect 29182 9072 29238 9081
rect 29012 9030 29182 9058
rect 29182 9007 29184 9016
rect 29236 9007 29238 9016
rect 29184 8978 29236 8984
rect 29184 7744 29236 7750
rect 29184 7686 29236 7692
rect 29000 7268 29052 7274
rect 29000 7210 29052 7216
rect 29012 6866 29040 7210
rect 29000 6860 29052 6866
rect 29000 6802 29052 6808
rect 28998 6760 29054 6769
rect 28998 6695 29054 6704
rect 28816 5772 28868 5778
rect 28816 5714 28868 5720
rect 28908 5772 28960 5778
rect 28908 5714 28960 5720
rect 28630 5672 28686 5681
rect 28630 5607 28686 5616
rect 28224 4984 28304 5012
rect 28172 4966 28224 4972
rect 28184 4622 28212 4966
rect 28920 4690 28948 5714
rect 29012 5574 29040 6695
rect 29196 6254 29224 7686
rect 29288 7478 29316 9590
rect 29380 7954 29408 12582
rect 29472 12374 29500 12650
rect 29460 12368 29512 12374
rect 29460 12310 29512 12316
rect 29460 11552 29512 11558
rect 29460 11494 29512 11500
rect 29472 10130 29500 11494
rect 29460 10124 29512 10130
rect 29460 10066 29512 10072
rect 29460 9920 29512 9926
rect 29460 9862 29512 9868
rect 29368 7948 29420 7954
rect 29368 7890 29420 7896
rect 29472 7750 29500 9862
rect 29460 7744 29512 7750
rect 29460 7686 29512 7692
rect 29472 7478 29500 7686
rect 29276 7472 29328 7478
rect 29276 7414 29328 7420
rect 29460 7472 29512 7478
rect 29460 7414 29512 7420
rect 29564 7342 29592 14062
rect 29644 14068 29696 14074
rect 29644 14010 29696 14016
rect 29828 13864 29880 13870
rect 29828 13806 29880 13812
rect 29840 13326 29868 13806
rect 29828 13320 29880 13326
rect 29828 13262 29880 13268
rect 29644 12776 29696 12782
rect 29644 12718 29696 12724
rect 29656 12646 29684 12718
rect 29932 12646 29960 14912
rect 29644 12640 29696 12646
rect 29644 12582 29696 12588
rect 29920 12640 29972 12646
rect 29920 12582 29972 12588
rect 30024 12442 30052 15438
rect 30116 15026 30144 15966
rect 30378 15943 30434 15952
rect 30944 15638 30972 20012
rect 31024 19916 31076 19922
rect 31024 19858 31076 19864
rect 31036 19446 31064 19858
rect 31024 19440 31076 19446
rect 31024 19382 31076 19388
rect 31036 17746 31064 19382
rect 31300 18828 31352 18834
rect 31300 18770 31352 18776
rect 31024 17740 31076 17746
rect 31024 17682 31076 17688
rect 31208 17740 31260 17746
rect 31208 17682 31260 17688
rect 31036 17134 31064 17682
rect 31116 17264 31168 17270
rect 31116 17206 31168 17212
rect 31024 17128 31076 17134
rect 31024 17070 31076 17076
rect 31128 16658 31156 17206
rect 31220 17202 31248 17682
rect 31312 17678 31340 18770
rect 31300 17672 31352 17678
rect 31300 17614 31352 17620
rect 31208 17196 31260 17202
rect 31208 17138 31260 17144
rect 31116 16652 31168 16658
rect 31116 16594 31168 16600
rect 31404 16130 31432 23054
rect 31496 21350 31524 23174
rect 31760 22636 31812 22642
rect 31760 22578 31812 22584
rect 31772 21418 31800 22578
rect 31852 22568 31904 22574
rect 31852 22510 31904 22516
rect 31864 22030 31892 22510
rect 31852 22024 31904 22030
rect 31852 21966 31904 21972
rect 31576 21412 31628 21418
rect 31576 21354 31628 21360
rect 31760 21412 31812 21418
rect 31760 21354 31812 21360
rect 31484 21344 31536 21350
rect 31484 21286 31536 21292
rect 31588 20890 31616 21354
rect 31956 21026 31984 24754
rect 32036 24744 32088 24750
rect 32036 24686 32088 24692
rect 32048 24138 32076 24686
rect 32324 24614 32352 26862
rect 32312 24608 32364 24614
rect 32312 24550 32364 24556
rect 32128 24268 32180 24274
rect 32128 24210 32180 24216
rect 32036 24132 32088 24138
rect 32036 24074 32088 24080
rect 32140 23866 32168 24210
rect 32128 23860 32180 23866
rect 32128 23802 32180 23808
rect 32416 23254 32444 26982
rect 32508 25838 32536 27406
rect 32496 25832 32548 25838
rect 32496 25774 32548 25780
rect 32600 24682 32628 28727
rect 32784 28626 32812 29514
rect 32772 28620 32824 28626
rect 32772 28562 32824 28568
rect 32876 28014 32904 29650
rect 32968 29646 32996 30126
rect 33140 29708 33192 29714
rect 33140 29650 33192 29656
rect 32956 29640 33008 29646
rect 32956 29582 33008 29588
rect 32968 29306 32996 29582
rect 32956 29300 33008 29306
rect 32956 29242 33008 29248
rect 33152 28694 33180 29650
rect 33140 28688 33192 28694
rect 33140 28630 33192 28636
rect 33428 28218 33456 30126
rect 33612 29714 33640 30330
rect 35268 30326 35296 30806
rect 35256 30320 35308 30326
rect 35256 30262 35308 30268
rect 34520 30184 34572 30190
rect 34520 30126 34572 30132
rect 34244 30116 34296 30122
rect 34244 30058 34296 30064
rect 33600 29708 33652 29714
rect 33600 29650 33652 29656
rect 34152 29640 34204 29646
rect 34152 29582 34204 29588
rect 33508 29028 33560 29034
rect 33508 28970 33560 28976
rect 33520 28762 33548 28970
rect 34164 28762 34192 29582
rect 33508 28756 33560 28762
rect 33508 28698 33560 28704
rect 34152 28756 34204 28762
rect 34152 28698 34204 28704
rect 33416 28212 33468 28218
rect 33416 28154 33468 28160
rect 32864 28008 32916 28014
rect 32864 27950 32916 27956
rect 33428 27606 33456 28154
rect 33520 28014 33548 28698
rect 34256 28626 34284 30058
rect 34428 29232 34480 29238
rect 34428 29174 34480 29180
rect 34244 28620 34296 28626
rect 34244 28562 34296 28568
rect 33784 28552 33836 28558
rect 33784 28494 33836 28500
rect 33508 28008 33560 28014
rect 33508 27950 33560 27956
rect 33416 27600 33468 27606
rect 33416 27542 33468 27548
rect 32956 27396 33008 27402
rect 32956 27338 33008 27344
rect 32772 26988 32824 26994
rect 32772 26930 32824 26936
rect 32680 26920 32732 26926
rect 32680 26862 32732 26868
rect 32692 26586 32720 26862
rect 32680 26580 32732 26586
rect 32680 26522 32732 26528
rect 32784 25362 32812 26930
rect 32968 26450 32996 27338
rect 33048 26512 33100 26518
rect 33048 26454 33100 26460
rect 32956 26444 33008 26450
rect 32956 26386 33008 26392
rect 32772 25356 32824 25362
rect 32772 25298 32824 25304
rect 32956 25288 33008 25294
rect 32956 25230 33008 25236
rect 32588 24676 32640 24682
rect 32588 24618 32640 24624
rect 32864 24608 32916 24614
rect 32864 24550 32916 24556
rect 32588 24064 32640 24070
rect 32588 24006 32640 24012
rect 32404 23248 32456 23254
rect 32404 23190 32456 23196
rect 32128 22092 32180 22098
rect 32128 22034 32180 22040
rect 32036 21412 32088 21418
rect 32036 21354 32088 21360
rect 31772 20998 31984 21026
rect 32048 21010 32076 21354
rect 32140 21078 32168 22034
rect 32600 21690 32628 24006
rect 32680 23180 32732 23186
rect 32680 23122 32732 23128
rect 32692 22642 32720 23122
rect 32680 22636 32732 22642
rect 32680 22578 32732 22584
rect 32680 22092 32732 22098
rect 32680 22034 32732 22040
rect 32692 21894 32720 22034
rect 32680 21888 32732 21894
rect 32680 21830 32732 21836
rect 32496 21684 32548 21690
rect 32496 21626 32548 21632
rect 32588 21684 32640 21690
rect 32588 21626 32640 21632
rect 32404 21616 32456 21622
rect 32404 21558 32456 21564
rect 32220 21412 32272 21418
rect 32220 21354 32272 21360
rect 32128 21072 32180 21078
rect 32128 21014 32180 21020
rect 32036 21004 32088 21010
rect 31772 20942 31800 20998
rect 32036 20946 32088 20952
rect 31496 20862 31616 20890
rect 31760 20936 31812 20942
rect 31760 20878 31812 20884
rect 31496 19310 31524 20862
rect 31668 20800 31720 20806
rect 31588 20760 31668 20788
rect 31588 20602 31616 20760
rect 31668 20742 31720 20748
rect 31576 20596 31628 20602
rect 31576 20538 31628 20544
rect 32048 20058 32076 20946
rect 32140 20330 32168 21014
rect 32128 20324 32180 20330
rect 32128 20266 32180 20272
rect 32036 20052 32088 20058
rect 32036 19994 32088 20000
rect 32128 19508 32180 19514
rect 32128 19450 32180 19456
rect 31484 19304 31536 19310
rect 31484 19246 31536 19252
rect 31760 19304 31812 19310
rect 31760 19246 31812 19252
rect 31496 18834 31524 19246
rect 31484 18828 31536 18834
rect 31484 18770 31536 18776
rect 31772 18154 31800 19246
rect 32036 18216 32088 18222
rect 32036 18158 32088 18164
rect 31760 18148 31812 18154
rect 31760 18090 31812 18096
rect 31772 17134 31800 18090
rect 32048 17882 32076 18158
rect 32036 17876 32088 17882
rect 32036 17818 32088 17824
rect 31760 17128 31812 17134
rect 31760 17070 31812 17076
rect 32036 16720 32088 16726
rect 32036 16662 32088 16668
rect 31668 16652 31720 16658
rect 31312 16102 31432 16130
rect 31588 16612 31668 16640
rect 31588 16114 31616 16612
rect 31668 16594 31720 16600
rect 31576 16108 31628 16114
rect 30932 15632 30984 15638
rect 30932 15574 30984 15580
rect 30748 15564 30800 15570
rect 30748 15506 30800 15512
rect 30104 15020 30156 15026
rect 30104 14962 30156 14968
rect 30116 14618 30144 14962
rect 30196 14952 30248 14958
rect 30196 14894 30248 14900
rect 30564 14952 30616 14958
rect 30564 14894 30616 14900
rect 30104 14612 30156 14618
rect 30104 14554 30156 14560
rect 30208 13394 30236 14894
rect 30576 14618 30604 14894
rect 30656 14816 30708 14822
rect 30656 14758 30708 14764
rect 30564 14612 30616 14618
rect 30564 14554 30616 14560
rect 30380 14476 30432 14482
rect 30380 14418 30432 14424
rect 30288 13796 30340 13802
rect 30288 13738 30340 13744
rect 30196 13388 30248 13394
rect 30196 13330 30248 13336
rect 30104 12776 30156 12782
rect 30104 12718 30156 12724
rect 29644 12436 29696 12442
rect 29644 12378 29696 12384
rect 30012 12436 30064 12442
rect 30012 12378 30064 12384
rect 29552 7336 29604 7342
rect 29552 7278 29604 7284
rect 29564 6866 29592 7278
rect 29552 6860 29604 6866
rect 29552 6802 29604 6808
rect 29276 6792 29328 6798
rect 29276 6734 29328 6740
rect 29288 6390 29316 6734
rect 29552 6656 29604 6662
rect 29552 6598 29604 6604
rect 29276 6384 29328 6390
rect 29276 6326 29328 6332
rect 29564 6322 29592 6598
rect 29552 6316 29604 6322
rect 29552 6258 29604 6264
rect 29184 6248 29236 6254
rect 29184 6190 29236 6196
rect 29092 6112 29144 6118
rect 29092 6054 29144 6060
rect 29000 5568 29052 5574
rect 29000 5510 29052 5516
rect 28908 4684 28960 4690
rect 28908 4626 28960 4632
rect 28172 4616 28224 4622
rect 28172 4558 28224 4564
rect 29104 4146 29132 6054
rect 29196 5234 29224 6190
rect 29656 6118 29684 12378
rect 30012 12096 30064 12102
rect 30012 12038 30064 12044
rect 29828 11892 29880 11898
rect 29828 11834 29880 11840
rect 29736 11620 29788 11626
rect 29736 11562 29788 11568
rect 29748 10674 29776 11562
rect 29840 11558 29868 11834
rect 29828 11552 29880 11558
rect 29828 11494 29880 11500
rect 29828 11212 29880 11218
rect 29828 11154 29880 11160
rect 29736 10668 29788 10674
rect 29736 10610 29788 10616
rect 29840 10606 29868 11154
rect 30024 10606 30052 12038
rect 30116 10742 30144 12718
rect 30208 11830 30236 13330
rect 30300 12306 30328 13738
rect 30392 13326 30420 14418
rect 30472 14340 30524 14346
rect 30472 14282 30524 14288
rect 30484 13870 30512 14282
rect 30472 13864 30524 13870
rect 30472 13806 30524 13812
rect 30668 13734 30696 14758
rect 30760 14482 30788 15506
rect 30748 14476 30800 14482
rect 30748 14418 30800 14424
rect 30932 14476 30984 14482
rect 30932 14418 30984 14424
rect 30944 13938 30972 14418
rect 30932 13932 30984 13938
rect 30932 13874 30984 13880
rect 30656 13728 30708 13734
rect 30656 13670 30708 13676
rect 30668 13394 30696 13670
rect 30656 13388 30708 13394
rect 30656 13330 30708 13336
rect 30380 13320 30432 13326
rect 30380 13262 30432 13268
rect 30288 12300 30340 12306
rect 30288 12242 30340 12248
rect 30300 12102 30328 12242
rect 30288 12096 30340 12102
rect 30288 12038 30340 12044
rect 30196 11824 30248 11830
rect 30196 11766 30248 11772
rect 30196 11688 30248 11694
rect 30196 11630 30248 11636
rect 30208 11257 30236 11630
rect 30194 11248 30250 11257
rect 30194 11183 30250 11192
rect 30104 10736 30156 10742
rect 30104 10678 30156 10684
rect 29828 10600 29880 10606
rect 29828 10542 29880 10548
rect 30012 10600 30064 10606
rect 30012 10542 30064 10548
rect 30196 10600 30248 10606
rect 30196 10542 30248 10548
rect 29736 9988 29788 9994
rect 29736 9930 29788 9936
rect 29748 9761 29776 9930
rect 29734 9752 29790 9761
rect 29734 9687 29790 9696
rect 29748 9518 29776 9687
rect 29736 9512 29788 9518
rect 29736 9454 29788 9460
rect 29736 9036 29788 9042
rect 29736 8978 29788 8984
rect 29748 8945 29776 8978
rect 29734 8936 29790 8945
rect 29840 8906 29868 10542
rect 30012 9988 30064 9994
rect 30012 9930 30064 9936
rect 30024 8974 30052 9930
rect 30012 8968 30064 8974
rect 30012 8910 30064 8916
rect 29734 8871 29790 8880
rect 29828 8900 29880 8906
rect 29828 8842 29880 8848
rect 30208 8430 30236 10542
rect 30392 10062 30420 13262
rect 30472 11688 30524 11694
rect 30472 11630 30524 11636
rect 30484 11354 30512 11630
rect 30472 11348 30524 11354
rect 30472 11290 30524 11296
rect 30564 11144 30616 11150
rect 30564 11086 30616 11092
rect 30576 10441 30604 11086
rect 30562 10432 30618 10441
rect 30562 10367 30618 10376
rect 30380 10056 30432 10062
rect 30380 9998 30432 10004
rect 30380 9920 30432 9926
rect 30380 9862 30432 9868
rect 30392 9654 30420 9862
rect 30380 9648 30432 9654
rect 30380 9590 30432 9596
rect 30288 9580 30340 9586
rect 30288 9522 30340 9528
rect 30196 8424 30248 8430
rect 30196 8366 30248 8372
rect 30104 8084 30156 8090
rect 30104 8026 30156 8032
rect 30116 7818 30144 8026
rect 30300 7954 30328 9522
rect 30562 8664 30618 8673
rect 30562 8599 30618 8608
rect 30472 8424 30524 8430
rect 30472 8366 30524 8372
rect 30288 7948 30340 7954
rect 30288 7890 30340 7896
rect 30104 7812 30156 7818
rect 30104 7754 30156 7760
rect 30300 7546 30328 7890
rect 30484 7886 30512 8366
rect 30472 7880 30524 7886
rect 30472 7822 30524 7828
rect 30484 7750 30512 7822
rect 30472 7744 30524 7750
rect 30472 7686 30524 7692
rect 30288 7540 30340 7546
rect 30288 7482 30340 7488
rect 29736 6928 29788 6934
rect 29736 6870 29788 6876
rect 29748 6662 29776 6870
rect 29736 6656 29788 6662
rect 29736 6598 29788 6604
rect 30196 6316 30248 6322
rect 30196 6258 30248 6264
rect 29644 6112 29696 6118
rect 29644 6054 29696 6060
rect 30208 5846 30236 6258
rect 30576 6254 30604 8599
rect 30668 8294 30696 13330
rect 31312 12306 31340 16102
rect 31576 16050 31628 16056
rect 31392 16040 31444 16046
rect 31392 15982 31444 15988
rect 31404 15502 31432 15982
rect 31392 15496 31444 15502
rect 31392 15438 31444 15444
rect 31392 14000 31444 14006
rect 31392 13942 31444 13948
rect 31404 13734 31432 13942
rect 31392 13728 31444 13734
rect 31392 13670 31444 13676
rect 31944 13728 31996 13734
rect 31944 13670 31996 13676
rect 31404 12918 31432 13670
rect 31852 13388 31904 13394
rect 31852 13330 31904 13336
rect 31576 13184 31628 13190
rect 31576 13126 31628 13132
rect 31392 12912 31444 12918
rect 31392 12854 31444 12860
rect 31300 12300 31352 12306
rect 31300 12242 31352 12248
rect 31208 12232 31260 12238
rect 31208 12174 31260 12180
rect 30748 12164 30800 12170
rect 30748 12106 30800 12112
rect 30760 11354 30788 12106
rect 31220 11694 31248 12174
rect 31312 12073 31340 12242
rect 31298 12064 31354 12073
rect 31298 11999 31354 12008
rect 31300 11892 31352 11898
rect 31300 11834 31352 11840
rect 31208 11688 31260 11694
rect 31208 11630 31260 11636
rect 30748 11348 30800 11354
rect 30748 11290 30800 11296
rect 30656 8288 30708 8294
rect 30656 8230 30708 8236
rect 30668 8022 30696 8230
rect 30656 8016 30708 8022
rect 30656 7958 30708 7964
rect 30760 7206 30788 11290
rect 31312 11218 31340 11834
rect 31588 11694 31616 13126
rect 31760 12232 31812 12238
rect 31760 12174 31812 12180
rect 31576 11688 31628 11694
rect 31576 11630 31628 11636
rect 31300 11212 31352 11218
rect 31300 11154 31352 11160
rect 31588 11064 31616 11630
rect 31668 11620 31720 11626
rect 31668 11562 31720 11568
rect 31312 11036 31616 11064
rect 31116 10532 31168 10538
rect 31036 10492 31116 10520
rect 30840 10056 30892 10062
rect 30840 9998 30892 10004
rect 30852 9518 30880 9998
rect 31036 9926 31064 10492
rect 31116 10474 31168 10480
rect 31208 10192 31260 10198
rect 31208 10134 31260 10140
rect 31116 10124 31168 10130
rect 31116 10066 31168 10072
rect 31024 9920 31076 9926
rect 31024 9862 31076 9868
rect 30840 9512 30892 9518
rect 30840 9454 30892 9460
rect 31036 8974 31064 9862
rect 31128 9654 31156 10066
rect 31116 9648 31168 9654
rect 31116 9590 31168 9596
rect 31024 8968 31076 8974
rect 31024 8910 31076 8916
rect 30932 8492 30984 8498
rect 30932 8434 30984 8440
rect 30944 8090 30972 8434
rect 31024 8424 31076 8430
rect 31024 8366 31076 8372
rect 30932 8084 30984 8090
rect 30932 8026 30984 8032
rect 30840 7336 30892 7342
rect 30840 7278 30892 7284
rect 30748 7200 30800 7206
rect 30748 7142 30800 7148
rect 30564 6248 30616 6254
rect 30564 6190 30616 6196
rect 30472 6112 30524 6118
rect 30472 6054 30524 6060
rect 30196 5840 30248 5846
rect 30196 5782 30248 5788
rect 30484 5710 30512 6054
rect 30012 5704 30064 5710
rect 30012 5646 30064 5652
rect 30472 5704 30524 5710
rect 30472 5646 30524 5652
rect 30024 5234 30052 5646
rect 29184 5228 29236 5234
rect 29184 5170 29236 5176
rect 30012 5228 30064 5234
rect 30012 5170 30064 5176
rect 29196 4146 29224 5170
rect 30656 5160 30708 5166
rect 30760 5148 30788 7142
rect 30852 6934 30880 7278
rect 30840 6928 30892 6934
rect 30840 6870 30892 6876
rect 30944 6458 30972 8026
rect 31036 6730 31064 8366
rect 31116 8288 31168 8294
rect 31116 8230 31168 8236
rect 31128 7410 31156 8230
rect 31116 7404 31168 7410
rect 31116 7346 31168 7352
rect 31024 6724 31076 6730
rect 31024 6666 31076 6672
rect 31220 6458 31248 10134
rect 31312 9518 31340 11036
rect 31680 10826 31708 11562
rect 31772 11218 31800 12174
rect 31760 11212 31812 11218
rect 31760 11154 31812 11160
rect 31864 11121 31892 13330
rect 31956 13326 31984 13670
rect 31944 13320 31996 13326
rect 31944 13262 31996 13268
rect 31956 11830 31984 13262
rect 31944 11824 31996 11830
rect 31944 11766 31996 11772
rect 31944 11688 31996 11694
rect 31942 11656 31944 11665
rect 31996 11656 31998 11665
rect 31942 11591 31998 11600
rect 31944 11280 31996 11286
rect 31944 11222 31996 11228
rect 31850 11112 31906 11121
rect 31760 11076 31812 11082
rect 31850 11047 31906 11056
rect 31760 11018 31812 11024
rect 31496 10798 31708 10826
rect 31392 9920 31444 9926
rect 31392 9862 31444 9868
rect 31300 9512 31352 9518
rect 31300 9454 31352 9460
rect 31312 9178 31340 9454
rect 31300 9172 31352 9178
rect 31300 9114 31352 9120
rect 31404 9042 31432 9862
rect 31496 9761 31524 10798
rect 31772 10690 31800 11018
rect 31680 10674 31800 10690
rect 31668 10668 31800 10674
rect 31720 10662 31800 10668
rect 31668 10610 31720 10616
rect 31956 10198 31984 11222
rect 31944 10192 31996 10198
rect 31944 10134 31996 10140
rect 31944 10056 31996 10062
rect 31944 9998 31996 10004
rect 31482 9752 31538 9761
rect 31482 9687 31538 9696
rect 31392 9036 31444 9042
rect 31392 8978 31444 8984
rect 31300 8968 31352 8974
rect 31300 8910 31352 8916
rect 31312 6798 31340 8910
rect 31496 7834 31524 9687
rect 31576 9376 31628 9382
rect 31576 9318 31628 9324
rect 31588 9110 31616 9318
rect 31668 9172 31720 9178
rect 31668 9114 31720 9120
rect 31576 9104 31628 9110
rect 31576 9046 31628 9052
rect 31496 7806 31616 7834
rect 31484 7744 31536 7750
rect 31484 7686 31536 7692
rect 31496 6866 31524 7686
rect 31484 6860 31536 6866
rect 31484 6802 31536 6808
rect 31588 6798 31616 7806
rect 31680 6866 31708 9114
rect 31758 9072 31814 9081
rect 31758 9007 31760 9016
rect 31812 9007 31814 9016
rect 31760 8978 31812 8984
rect 31956 8838 31984 9998
rect 31944 8832 31996 8838
rect 31944 8774 31996 8780
rect 31944 6996 31996 7002
rect 31944 6938 31996 6944
rect 31668 6860 31720 6866
rect 31668 6802 31720 6808
rect 31300 6792 31352 6798
rect 31300 6734 31352 6740
rect 31576 6792 31628 6798
rect 31576 6734 31628 6740
rect 30932 6452 30984 6458
rect 30932 6394 30984 6400
rect 31208 6452 31260 6458
rect 31208 6394 31260 6400
rect 31220 6322 31248 6394
rect 31956 6361 31984 6938
rect 31942 6352 31998 6361
rect 31208 6316 31260 6322
rect 31942 6287 31998 6296
rect 31208 6258 31260 6264
rect 31944 6248 31996 6254
rect 31944 6190 31996 6196
rect 31208 5704 31260 5710
rect 31208 5646 31260 5652
rect 30932 5568 30984 5574
rect 30932 5510 30984 5516
rect 30944 5370 30972 5510
rect 30932 5364 30984 5370
rect 30932 5306 30984 5312
rect 30708 5120 30788 5148
rect 30840 5160 30892 5166
rect 30656 5102 30708 5108
rect 30840 5102 30892 5108
rect 30380 4752 30432 4758
rect 30380 4694 30432 4700
rect 29828 4616 29880 4622
rect 29828 4558 29880 4564
rect 29092 4140 29144 4146
rect 29092 4082 29144 4088
rect 29184 4140 29236 4146
rect 29184 4082 29236 4088
rect 28448 4072 28500 4078
rect 28448 4014 28500 4020
rect 28080 4004 28132 4010
rect 28080 3946 28132 3952
rect 28092 3602 28120 3946
rect 28460 3738 28488 4014
rect 28448 3732 28500 3738
rect 28448 3674 28500 3680
rect 28080 3596 28132 3602
rect 28080 3538 28132 3544
rect 29104 2990 29132 4082
rect 29196 3534 29224 4082
rect 29368 4072 29420 4078
rect 29368 4014 29420 4020
rect 29552 4072 29604 4078
rect 29552 4014 29604 4020
rect 29380 3670 29408 4014
rect 29368 3664 29420 3670
rect 29368 3606 29420 3612
rect 29184 3528 29236 3534
rect 29184 3470 29236 3476
rect 29564 3058 29592 4014
rect 29840 3058 29868 4558
rect 30288 4140 30340 4146
rect 30288 4082 30340 4088
rect 30196 3936 30248 3942
rect 30196 3878 30248 3884
rect 30208 3738 30236 3878
rect 30196 3732 30248 3738
rect 30196 3674 30248 3680
rect 29552 3052 29604 3058
rect 29552 2994 29604 3000
rect 29828 3052 29880 3058
rect 29828 2994 29880 3000
rect 27896 2984 27948 2990
rect 27896 2926 27948 2932
rect 29092 2984 29144 2990
rect 29092 2926 29144 2932
rect 30300 2938 30328 4082
rect 30392 3602 30420 4694
rect 30852 4690 30880 5102
rect 30944 4826 30972 5306
rect 31116 5296 31168 5302
rect 31116 5238 31168 5244
rect 31128 5098 31156 5238
rect 31116 5092 31168 5098
rect 31116 5034 31168 5040
rect 31128 4826 31156 5034
rect 31220 4826 31248 5646
rect 31956 5642 31984 6190
rect 32048 5930 32076 16662
rect 32140 13870 32168 19450
rect 32232 18222 32260 21354
rect 32312 21140 32364 21146
rect 32312 21082 32364 21088
rect 32324 20398 32352 21082
rect 32416 21078 32444 21558
rect 32404 21072 32456 21078
rect 32404 21014 32456 21020
rect 32508 20942 32536 21626
rect 32496 20936 32548 20942
rect 32496 20878 32548 20884
rect 32312 20392 32364 20398
rect 32312 20334 32364 20340
rect 32324 18222 32352 20334
rect 32220 18216 32272 18222
rect 32220 18158 32272 18164
rect 32312 18216 32364 18222
rect 32312 18158 32364 18164
rect 32508 16590 32536 20878
rect 32600 19990 32628 21626
rect 32692 21418 32720 21830
rect 32772 21548 32824 21554
rect 32772 21490 32824 21496
rect 32680 21412 32732 21418
rect 32680 21354 32732 21360
rect 32588 19984 32640 19990
rect 32588 19926 32640 19932
rect 32784 19922 32812 21490
rect 32876 21010 32904 24550
rect 32968 23254 32996 25230
rect 33060 24750 33088 26454
rect 33428 25838 33456 27542
rect 33796 27334 33824 28494
rect 34336 27464 34388 27470
rect 34336 27406 34388 27412
rect 33784 27328 33836 27334
rect 33784 27270 33836 27276
rect 33796 27130 33824 27270
rect 33784 27124 33836 27130
rect 33784 27066 33836 27072
rect 34348 26994 34376 27406
rect 34336 26988 34388 26994
rect 34336 26930 34388 26936
rect 33968 26240 34020 26246
rect 33968 26182 34020 26188
rect 33980 25906 34008 26182
rect 33968 25900 34020 25906
rect 33968 25842 34020 25848
rect 33416 25832 33468 25838
rect 33416 25774 33468 25780
rect 33968 25356 34020 25362
rect 33968 25298 34020 25304
rect 33784 25152 33836 25158
rect 33784 25094 33836 25100
rect 33048 24744 33100 24750
rect 33048 24686 33100 24692
rect 33060 24070 33088 24686
rect 33600 24676 33652 24682
rect 33600 24618 33652 24624
rect 33416 24268 33468 24274
rect 33416 24210 33468 24216
rect 33324 24200 33376 24206
rect 33324 24142 33376 24148
rect 33048 24064 33100 24070
rect 33048 24006 33100 24012
rect 32956 23248 33008 23254
rect 32956 23190 33008 23196
rect 33140 22432 33192 22438
rect 33140 22374 33192 22380
rect 33152 21962 33180 22374
rect 33336 22098 33364 24142
rect 33324 22092 33376 22098
rect 33324 22034 33376 22040
rect 33140 21956 33192 21962
rect 33140 21898 33192 21904
rect 33232 21956 33284 21962
rect 33232 21898 33284 21904
rect 33244 21622 33272 21898
rect 33232 21616 33284 21622
rect 33232 21558 33284 21564
rect 33048 21548 33100 21554
rect 33048 21490 33100 21496
rect 33060 21146 33088 21490
rect 33244 21162 33272 21558
rect 33048 21140 33100 21146
rect 33048 21082 33100 21088
rect 33152 21134 33272 21162
rect 32864 21004 32916 21010
rect 32864 20946 32916 20952
rect 32956 20256 33008 20262
rect 32956 20198 33008 20204
rect 32968 19922 32996 20198
rect 32772 19916 32824 19922
rect 32772 19858 32824 19864
rect 32956 19916 33008 19922
rect 32956 19858 33008 19864
rect 32956 19304 33008 19310
rect 32956 19246 33008 19252
rect 32772 19168 32824 19174
rect 32772 19110 32824 19116
rect 32784 18222 32812 19110
rect 32968 18970 32996 19246
rect 33060 19242 33088 21082
rect 33152 19310 33180 21134
rect 33232 20392 33284 20398
rect 33232 20334 33284 20340
rect 33140 19304 33192 19310
rect 33140 19246 33192 19252
rect 33048 19236 33100 19242
rect 33048 19178 33100 19184
rect 32956 18964 33008 18970
rect 32956 18906 33008 18912
rect 32772 18216 32824 18222
rect 32772 18158 32824 18164
rect 33140 18216 33192 18222
rect 33140 18158 33192 18164
rect 32588 18080 32640 18086
rect 32588 18022 32640 18028
rect 32600 16794 32628 18022
rect 32784 17898 32812 18158
rect 32784 17870 32904 17898
rect 32772 17740 32824 17746
rect 32772 17682 32824 17688
rect 32588 16788 32640 16794
rect 32588 16730 32640 16736
rect 32496 16584 32548 16590
rect 32496 16526 32548 16532
rect 32508 15502 32536 16526
rect 32784 15706 32812 17682
rect 32772 15700 32824 15706
rect 32772 15642 32824 15648
rect 32496 15496 32548 15502
rect 32496 15438 32548 15444
rect 32784 14482 32812 15642
rect 32876 14618 32904 17870
rect 33048 17808 33100 17814
rect 33152 17796 33180 18158
rect 33100 17768 33180 17796
rect 33048 17750 33100 17756
rect 32956 17060 33008 17066
rect 32956 17002 33008 17008
rect 32864 14612 32916 14618
rect 32864 14554 32916 14560
rect 32772 14476 32824 14482
rect 32772 14418 32824 14424
rect 32220 14408 32272 14414
rect 32220 14350 32272 14356
rect 32128 13864 32180 13870
rect 32128 13806 32180 13812
rect 32232 12374 32260 14350
rect 32772 14272 32824 14278
rect 32772 14214 32824 14220
rect 32784 13870 32812 14214
rect 32772 13864 32824 13870
rect 32772 13806 32824 13812
rect 32876 13530 32904 14554
rect 32968 14482 32996 17002
rect 33060 16726 33088 17750
rect 33048 16720 33100 16726
rect 33048 16662 33100 16668
rect 33060 16250 33088 16662
rect 33048 16244 33100 16250
rect 33048 16186 33100 16192
rect 33048 15564 33100 15570
rect 33048 15506 33100 15512
rect 33060 14958 33088 15506
rect 33244 15484 33272 20334
rect 33428 19990 33456 24210
rect 33612 22624 33640 24618
rect 33692 24064 33744 24070
rect 33692 24006 33744 24012
rect 33704 23186 33732 24006
rect 33692 23180 33744 23186
rect 33692 23122 33744 23128
rect 33612 22596 33732 22624
rect 33600 22500 33652 22506
rect 33600 22442 33652 22448
rect 33508 22228 33560 22234
rect 33508 22170 33560 22176
rect 33416 19984 33468 19990
rect 33416 19926 33468 19932
rect 33324 19372 33376 19378
rect 33324 19314 33376 19320
rect 33336 18834 33364 19314
rect 33324 18828 33376 18834
rect 33324 18770 33376 18776
rect 33520 17354 33548 22170
rect 33612 19310 33640 22442
rect 33704 21894 33732 22596
rect 33796 22574 33824 25094
rect 33980 24818 34008 25298
rect 34348 25294 34376 26930
rect 34440 26042 34468 29174
rect 34532 28218 34560 30126
rect 34612 30048 34664 30054
rect 34612 29990 34664 29996
rect 34520 28212 34572 28218
rect 34520 28154 34572 28160
rect 34624 26926 34652 29990
rect 35256 29504 35308 29510
rect 35256 29446 35308 29452
rect 34940 29404 35236 29424
rect 34996 29402 35020 29404
rect 35076 29402 35100 29404
rect 35156 29402 35180 29404
rect 35018 29350 35020 29402
rect 35082 29350 35094 29402
rect 35156 29350 35158 29402
rect 34996 29348 35020 29350
rect 35076 29348 35100 29350
rect 35156 29348 35180 29350
rect 34940 29328 35236 29348
rect 35268 29102 35296 29446
rect 35360 29170 35388 31214
rect 35440 31204 35492 31210
rect 35440 31146 35492 31152
rect 35348 29164 35400 29170
rect 35348 29106 35400 29112
rect 35256 29096 35308 29102
rect 35256 29038 35308 29044
rect 34704 29028 34756 29034
rect 34704 28970 34756 28976
rect 34716 27538 34744 28970
rect 34940 28316 35236 28336
rect 34996 28314 35020 28316
rect 35076 28314 35100 28316
rect 35156 28314 35180 28316
rect 35018 28262 35020 28314
rect 35082 28262 35094 28314
rect 35156 28262 35158 28314
rect 34996 28260 35020 28262
rect 35076 28260 35100 28262
rect 35156 28260 35180 28262
rect 34940 28240 35236 28260
rect 35268 28014 35296 29038
rect 35452 29034 35480 31146
rect 35544 29594 35572 31334
rect 35636 30802 35664 32710
rect 35728 31822 35756 32846
rect 35808 32224 35860 32230
rect 35808 32166 35860 32172
rect 35820 31890 35848 32166
rect 35808 31884 35860 31890
rect 35808 31826 35860 31832
rect 35716 31816 35768 31822
rect 35716 31758 35768 31764
rect 35624 30796 35676 30802
rect 35624 30738 35676 30744
rect 35624 30184 35676 30190
rect 35624 30126 35676 30132
rect 35636 29714 35664 30126
rect 35900 30116 35952 30122
rect 35900 30058 35952 30064
rect 35624 29708 35676 29714
rect 35624 29650 35676 29656
rect 35544 29566 35664 29594
rect 35532 29096 35584 29102
rect 35532 29038 35584 29044
rect 35440 29028 35492 29034
rect 35440 28970 35492 28976
rect 35544 28626 35572 29038
rect 35532 28620 35584 28626
rect 35532 28562 35584 28568
rect 35544 28014 35572 28562
rect 35256 28008 35308 28014
rect 35256 27950 35308 27956
rect 35532 28008 35584 28014
rect 35532 27950 35584 27956
rect 34704 27532 34756 27538
rect 34704 27474 34756 27480
rect 35544 27334 35572 27950
rect 35532 27328 35584 27334
rect 35532 27270 35584 27276
rect 34940 27228 35236 27248
rect 34996 27226 35020 27228
rect 35076 27226 35100 27228
rect 35156 27226 35180 27228
rect 35018 27174 35020 27226
rect 35082 27174 35094 27226
rect 35156 27174 35158 27226
rect 34996 27172 35020 27174
rect 35076 27172 35100 27174
rect 35156 27172 35180 27174
rect 34940 27152 35236 27172
rect 34612 26920 34664 26926
rect 34612 26862 34664 26868
rect 34704 26444 34756 26450
rect 34704 26386 34756 26392
rect 35348 26444 35400 26450
rect 35348 26386 35400 26392
rect 34612 26240 34664 26246
rect 34612 26182 34664 26188
rect 34428 26036 34480 26042
rect 34428 25978 34480 25984
rect 34520 25900 34572 25906
rect 34520 25842 34572 25848
rect 34336 25288 34388 25294
rect 34336 25230 34388 25236
rect 33968 24812 34020 24818
rect 34020 24772 34100 24800
rect 33968 24754 34020 24760
rect 33966 24712 34022 24721
rect 33966 24647 33968 24656
rect 34020 24647 34022 24656
rect 33968 24618 34020 24624
rect 34072 22574 34100 24772
rect 34348 24682 34376 25230
rect 34532 24818 34560 25842
rect 34624 25838 34652 26182
rect 34612 25832 34664 25838
rect 34612 25774 34664 25780
rect 34520 24812 34572 24818
rect 34520 24754 34572 24760
rect 34612 24812 34664 24818
rect 34612 24754 34664 24760
rect 34336 24676 34388 24682
rect 34336 24618 34388 24624
rect 34520 24268 34572 24274
rect 34520 24210 34572 24216
rect 34244 24200 34296 24206
rect 34244 24142 34296 24148
rect 34256 23526 34284 24142
rect 34336 23588 34388 23594
rect 34336 23530 34388 23536
rect 34244 23520 34296 23526
rect 34244 23462 34296 23468
rect 33784 22568 33836 22574
rect 33784 22510 33836 22516
rect 34060 22568 34112 22574
rect 34060 22510 34112 22516
rect 34256 22166 34284 23462
rect 34244 22160 34296 22166
rect 34244 22102 34296 22108
rect 33692 21888 33744 21894
rect 33692 21830 33744 21836
rect 34244 21888 34296 21894
rect 34244 21830 34296 21836
rect 33968 21480 34020 21486
rect 33968 21422 34020 21428
rect 34256 21434 34284 21830
rect 34348 21554 34376 23530
rect 34532 23322 34560 24210
rect 34520 23316 34572 23322
rect 34520 23258 34572 23264
rect 34624 22642 34652 24754
rect 34716 24410 34744 26386
rect 34796 26376 34848 26382
rect 34796 26318 34848 26324
rect 34704 24404 34756 24410
rect 34704 24346 34756 24352
rect 34808 24342 34836 26318
rect 34940 26140 35236 26160
rect 34996 26138 35020 26140
rect 35076 26138 35100 26140
rect 35156 26138 35180 26140
rect 35018 26086 35020 26138
rect 35082 26086 35094 26138
rect 35156 26086 35158 26138
rect 34996 26084 35020 26086
rect 35076 26084 35100 26086
rect 35156 26084 35180 26086
rect 34940 26064 35236 26084
rect 35360 26042 35388 26386
rect 35348 26036 35400 26042
rect 35348 25978 35400 25984
rect 35544 25838 35572 27270
rect 35532 25832 35584 25838
rect 35532 25774 35584 25780
rect 35636 25650 35664 29566
rect 35912 27146 35940 30058
rect 35728 27118 35940 27146
rect 35728 26926 35756 27118
rect 35716 26920 35768 26926
rect 35716 26862 35768 26868
rect 35544 25622 35664 25650
rect 35440 25492 35492 25498
rect 35440 25434 35492 25440
rect 35452 25401 35480 25434
rect 35438 25392 35494 25401
rect 35438 25327 35494 25336
rect 35544 25276 35572 25622
rect 35624 25492 35676 25498
rect 35624 25434 35676 25440
rect 35452 25248 35572 25276
rect 34940 25052 35236 25072
rect 34996 25050 35020 25052
rect 35076 25050 35100 25052
rect 35156 25050 35180 25052
rect 35018 24998 35020 25050
rect 35082 24998 35094 25050
rect 35156 24998 35158 25050
rect 34996 24996 35020 24998
rect 35076 24996 35100 24998
rect 35156 24996 35180 24998
rect 34940 24976 35236 24996
rect 34796 24336 34848 24342
rect 34796 24278 34848 24284
rect 34704 24268 34756 24274
rect 34704 24210 34756 24216
rect 34716 22982 34744 24210
rect 34940 23964 35236 23984
rect 34996 23962 35020 23964
rect 35076 23962 35100 23964
rect 35156 23962 35180 23964
rect 35018 23910 35020 23962
rect 35082 23910 35094 23962
rect 35156 23910 35158 23962
rect 34996 23908 35020 23910
rect 35076 23908 35100 23910
rect 35156 23908 35180 23910
rect 34940 23888 35236 23908
rect 34796 23656 34848 23662
rect 34796 23598 34848 23604
rect 34704 22976 34756 22982
rect 34704 22918 34756 22924
rect 34612 22636 34664 22642
rect 34612 22578 34664 22584
rect 34808 22030 34836 23598
rect 35452 23474 35480 25248
rect 35532 25152 35584 25158
rect 35532 25094 35584 25100
rect 35544 23662 35572 25094
rect 35532 23656 35584 23662
rect 35532 23598 35584 23604
rect 35452 23446 35572 23474
rect 34940 22876 35236 22896
rect 34996 22874 35020 22876
rect 35076 22874 35100 22876
rect 35156 22874 35180 22876
rect 35018 22822 35020 22874
rect 35082 22822 35094 22874
rect 35156 22822 35158 22874
rect 34996 22820 35020 22822
rect 35076 22820 35100 22822
rect 35156 22820 35180 22822
rect 34940 22800 35236 22820
rect 35346 22672 35402 22681
rect 35346 22607 35402 22616
rect 35360 22574 35388 22607
rect 35348 22568 35400 22574
rect 35348 22510 35400 22516
rect 34796 22024 34848 22030
rect 34796 21966 34848 21972
rect 34428 21956 34480 21962
rect 34428 21898 34480 21904
rect 34440 21690 34468 21898
rect 34940 21788 35236 21808
rect 34996 21786 35020 21788
rect 35076 21786 35100 21788
rect 35156 21786 35180 21788
rect 35018 21734 35020 21786
rect 35082 21734 35094 21786
rect 35156 21734 35158 21786
rect 34996 21732 35020 21734
rect 35076 21732 35100 21734
rect 35156 21732 35180 21734
rect 34940 21712 35236 21732
rect 34428 21684 34480 21690
rect 34428 21626 34480 21632
rect 34336 21548 34388 21554
rect 34336 21490 34388 21496
rect 33876 21004 33928 21010
rect 33876 20946 33928 20952
rect 33600 19304 33652 19310
rect 33600 19246 33652 19252
rect 33784 18828 33836 18834
rect 33784 18770 33836 18776
rect 33796 17814 33824 18770
rect 33784 17808 33836 17814
rect 33784 17750 33836 17756
rect 33336 17326 33640 17354
rect 33336 17270 33364 17326
rect 33324 17264 33376 17270
rect 33324 17206 33376 17212
rect 33508 17196 33560 17202
rect 33508 17138 33560 17144
rect 33416 16652 33468 16658
rect 33416 16594 33468 16600
rect 33324 16584 33376 16590
rect 33324 16526 33376 16532
rect 33336 16046 33364 16526
rect 33428 16046 33456 16594
rect 33520 16522 33548 17138
rect 33508 16516 33560 16522
rect 33508 16458 33560 16464
rect 33324 16040 33376 16046
rect 33324 15982 33376 15988
rect 33416 16040 33468 16046
rect 33416 15982 33468 15988
rect 33428 15638 33456 15982
rect 33416 15632 33468 15638
rect 33416 15574 33468 15580
rect 33324 15496 33376 15502
rect 33244 15456 33324 15484
rect 33324 15438 33376 15444
rect 33048 14952 33100 14958
rect 33048 14894 33100 14900
rect 33508 14544 33560 14550
rect 33508 14486 33560 14492
rect 32956 14476 33008 14482
rect 32956 14418 33008 14424
rect 33520 14278 33548 14486
rect 33508 14272 33560 14278
rect 33508 14214 33560 14220
rect 33232 13932 33284 13938
rect 33232 13874 33284 13880
rect 32864 13524 32916 13530
rect 32864 13466 32916 13472
rect 33244 13394 33272 13874
rect 33324 13864 33376 13870
rect 33324 13806 33376 13812
rect 33232 13388 33284 13394
rect 33232 13330 33284 13336
rect 32772 13252 32824 13258
rect 32772 13194 32824 13200
rect 33140 13252 33192 13258
rect 33140 13194 33192 13200
rect 32784 12782 32812 13194
rect 32772 12776 32824 12782
rect 32772 12718 32824 12724
rect 32956 12708 33008 12714
rect 32956 12650 33008 12656
rect 32220 12368 32272 12374
rect 32220 12310 32272 12316
rect 32312 12368 32364 12374
rect 32312 12310 32364 12316
rect 32496 12368 32548 12374
rect 32496 12310 32548 12316
rect 32128 12232 32180 12238
rect 32128 12174 32180 12180
rect 32140 10470 32168 12174
rect 32220 11756 32272 11762
rect 32220 11698 32272 11704
rect 32232 10742 32260 11698
rect 32220 10736 32272 10742
rect 32220 10678 32272 10684
rect 32128 10464 32180 10470
rect 32128 10406 32180 10412
rect 32140 9518 32168 10406
rect 32324 10062 32352 12310
rect 32404 12300 32456 12306
rect 32404 12242 32456 12248
rect 32312 10056 32364 10062
rect 32312 9998 32364 10004
rect 32416 9722 32444 12242
rect 32508 11694 32536 12310
rect 32864 12232 32916 12238
rect 32864 12174 32916 12180
rect 32496 11688 32548 11694
rect 32496 11630 32548 11636
rect 32680 11620 32732 11626
rect 32680 11562 32732 11568
rect 32692 11218 32720 11562
rect 32680 11212 32732 11218
rect 32680 11154 32732 11160
rect 32876 10674 32904 12174
rect 32864 10668 32916 10674
rect 32864 10610 32916 10616
rect 32588 10600 32640 10606
rect 32586 10568 32588 10577
rect 32640 10568 32642 10577
rect 32586 10503 32642 10512
rect 32600 9926 32628 10503
rect 32968 10130 32996 12650
rect 33048 11552 33100 11558
rect 33048 11494 33100 11500
rect 33060 11218 33088 11494
rect 33152 11286 33180 13194
rect 33336 13190 33364 13806
rect 33324 13184 33376 13190
rect 33324 13126 33376 13132
rect 33336 11694 33364 13126
rect 33520 12238 33548 14214
rect 33508 12232 33560 12238
rect 33508 12174 33560 12180
rect 33414 12064 33470 12073
rect 33414 11999 33470 12008
rect 33324 11688 33376 11694
rect 33324 11630 33376 11636
rect 33140 11280 33192 11286
rect 33140 11222 33192 11228
rect 33048 11212 33100 11218
rect 33048 11154 33100 11160
rect 33048 10600 33100 10606
rect 33048 10542 33100 10548
rect 32956 10124 33008 10130
rect 32956 10066 33008 10072
rect 32864 9988 32916 9994
rect 32864 9930 32916 9936
rect 32588 9920 32640 9926
rect 32588 9862 32640 9868
rect 32404 9716 32456 9722
rect 32404 9658 32456 9664
rect 32128 9512 32180 9518
rect 32128 9454 32180 9460
rect 32312 9512 32364 9518
rect 32312 9454 32364 9460
rect 32140 8090 32168 9454
rect 32324 8090 32352 9454
rect 32416 9178 32444 9658
rect 32772 9444 32824 9450
rect 32772 9386 32824 9392
rect 32404 9172 32456 9178
rect 32404 9114 32456 9120
rect 32128 8084 32180 8090
rect 32128 8026 32180 8032
rect 32312 8084 32364 8090
rect 32312 8026 32364 8032
rect 32140 7002 32168 8026
rect 32220 7812 32272 7818
rect 32220 7754 32272 7760
rect 32128 6996 32180 7002
rect 32128 6938 32180 6944
rect 32232 6662 32260 7754
rect 32324 6866 32352 8026
rect 32416 7954 32444 9114
rect 32784 8430 32812 9386
rect 32876 8430 32904 9930
rect 32968 9518 32996 10066
rect 33060 10062 33088 10542
rect 33428 10130 33456 11999
rect 33520 10690 33548 12174
rect 33612 11150 33640 17326
rect 33888 15026 33916 20946
rect 33980 20398 34008 21422
rect 34256 21406 34376 21434
rect 34152 20936 34204 20942
rect 34152 20878 34204 20884
rect 33968 20392 34020 20398
rect 33968 20334 34020 20340
rect 33980 17882 34008 20334
rect 34164 19922 34192 20878
rect 34152 19916 34204 19922
rect 34152 19858 34204 19864
rect 34244 19304 34296 19310
rect 34244 19246 34296 19252
rect 34256 18902 34284 19246
rect 34244 18896 34296 18902
rect 34244 18838 34296 18844
rect 34152 18760 34204 18766
rect 34152 18702 34204 18708
rect 34164 18358 34192 18702
rect 34152 18352 34204 18358
rect 34152 18294 34204 18300
rect 33968 17876 34020 17882
rect 33968 17818 34020 17824
rect 33980 16522 34008 17818
rect 34348 17762 34376 21406
rect 34440 21010 34468 21626
rect 35256 21480 35308 21486
rect 35256 21422 35308 21428
rect 34428 21004 34480 21010
rect 34428 20946 34480 20952
rect 34704 21004 34756 21010
rect 34704 20946 34756 20952
rect 34428 20324 34480 20330
rect 34428 20266 34480 20272
rect 34256 17734 34376 17762
rect 34440 17746 34468 20266
rect 34716 20262 34744 20946
rect 34940 20700 35236 20720
rect 34996 20698 35020 20700
rect 35076 20698 35100 20700
rect 35156 20698 35180 20700
rect 35018 20646 35020 20698
rect 35082 20646 35094 20698
rect 35156 20646 35158 20698
rect 34996 20644 35020 20646
rect 35076 20644 35100 20646
rect 35156 20644 35180 20646
rect 34940 20624 35236 20644
rect 35268 20534 35296 21422
rect 35256 20528 35308 20534
rect 35256 20470 35308 20476
rect 34704 20256 34756 20262
rect 34704 20198 34756 20204
rect 34716 19242 34744 20198
rect 35268 19854 35296 20470
rect 35360 20262 35388 22510
rect 35544 22409 35572 23446
rect 35636 22506 35664 25434
rect 35716 25288 35768 25294
rect 35716 25230 35768 25236
rect 35728 23730 35756 25230
rect 35912 24342 35940 27118
rect 35992 26852 36044 26858
rect 35992 26794 36044 26800
rect 36004 26450 36032 26794
rect 35992 26444 36044 26450
rect 35992 26386 36044 26392
rect 36084 24744 36136 24750
rect 36084 24686 36136 24692
rect 35900 24336 35952 24342
rect 35900 24278 35952 24284
rect 35716 23724 35768 23730
rect 35716 23666 35768 23672
rect 35912 23118 35940 24278
rect 36096 23730 36124 24686
rect 36084 23724 36136 23730
rect 36084 23666 36136 23672
rect 35992 23180 36044 23186
rect 35992 23122 36044 23128
rect 35900 23112 35952 23118
rect 35900 23054 35952 23060
rect 35808 22976 35860 22982
rect 35808 22918 35860 22924
rect 35624 22500 35676 22506
rect 35624 22442 35676 22448
rect 35530 22400 35586 22409
rect 35636 22386 35664 22442
rect 35636 22358 35756 22386
rect 35530 22335 35586 22344
rect 35532 21956 35584 21962
rect 35532 21898 35584 21904
rect 35348 20256 35400 20262
rect 35348 20198 35400 20204
rect 35544 19990 35572 21898
rect 35728 21010 35756 22358
rect 35820 22098 35848 22918
rect 35808 22092 35860 22098
rect 35808 22034 35860 22040
rect 35716 21004 35768 21010
rect 35716 20946 35768 20952
rect 35716 20392 35768 20398
rect 35716 20334 35768 20340
rect 35728 20262 35756 20334
rect 35716 20256 35768 20262
rect 35716 20198 35768 20204
rect 35532 19984 35584 19990
rect 35532 19926 35584 19932
rect 35256 19848 35308 19854
rect 35256 19790 35308 19796
rect 34940 19612 35236 19632
rect 34996 19610 35020 19612
rect 35076 19610 35100 19612
rect 35156 19610 35180 19612
rect 35018 19558 35020 19610
rect 35082 19558 35094 19610
rect 35156 19558 35158 19610
rect 34996 19556 35020 19558
rect 35076 19556 35100 19558
rect 35156 19556 35180 19558
rect 34940 19536 35236 19556
rect 35544 19310 35572 19926
rect 34980 19304 35032 19310
rect 34980 19246 35032 19252
rect 35532 19304 35584 19310
rect 35532 19246 35584 19252
rect 34704 19236 34756 19242
rect 34704 19178 34756 19184
rect 34796 19168 34848 19174
rect 34796 19110 34848 19116
rect 34520 18760 34572 18766
rect 34520 18702 34572 18708
rect 34532 18290 34560 18702
rect 34704 18692 34756 18698
rect 34704 18634 34756 18640
rect 34520 18284 34572 18290
rect 34520 18226 34572 18232
rect 34716 18222 34744 18634
rect 34704 18216 34756 18222
rect 34704 18158 34756 18164
rect 34808 17746 34836 19110
rect 34992 18834 35020 19246
rect 34980 18828 35032 18834
rect 34980 18770 35032 18776
rect 35440 18828 35492 18834
rect 35440 18770 35492 18776
rect 34940 18524 35236 18544
rect 34996 18522 35020 18524
rect 35076 18522 35100 18524
rect 35156 18522 35180 18524
rect 35018 18470 35020 18522
rect 35082 18470 35094 18522
rect 35156 18470 35158 18522
rect 34996 18468 35020 18470
rect 35076 18468 35100 18470
rect 35156 18468 35180 18470
rect 34940 18448 35236 18468
rect 34980 18080 35032 18086
rect 34980 18022 35032 18028
rect 34992 17746 35020 18022
rect 34428 17740 34480 17746
rect 33968 16516 34020 16522
rect 33968 16458 34020 16464
rect 33980 15638 34008 16458
rect 33968 15632 34020 15638
rect 33968 15574 34020 15580
rect 33980 15094 34008 15574
rect 34060 15564 34112 15570
rect 34060 15506 34112 15512
rect 33968 15088 34020 15094
rect 33968 15030 34020 15036
rect 33876 15020 33928 15026
rect 33876 14962 33928 14968
rect 33968 14952 34020 14958
rect 33968 14894 34020 14900
rect 33980 14618 34008 14894
rect 33968 14612 34020 14618
rect 33968 14554 34020 14560
rect 33784 14000 33836 14006
rect 33784 13942 33836 13948
rect 33692 13728 33744 13734
rect 33692 13670 33744 13676
rect 33704 13190 33732 13670
rect 33692 13184 33744 13190
rect 33692 13126 33744 13132
rect 33704 11234 33732 13126
rect 33796 11762 33824 13942
rect 33980 13938 34008 14554
rect 33968 13932 34020 13938
rect 33968 13874 34020 13880
rect 34072 13818 34100 15506
rect 34256 15162 34284 17734
rect 34428 17682 34480 17688
rect 34796 17740 34848 17746
rect 34796 17682 34848 17688
rect 34980 17740 35032 17746
rect 34980 17682 35032 17688
rect 34336 17672 34388 17678
rect 34336 17614 34388 17620
rect 34348 17134 34376 17614
rect 34612 17604 34664 17610
rect 34612 17546 34664 17552
rect 34520 17536 34572 17542
rect 34520 17478 34572 17484
rect 34336 17128 34388 17134
rect 34336 17070 34388 17076
rect 34532 16658 34560 17478
rect 34520 16652 34572 16658
rect 34520 16594 34572 16600
rect 34244 15156 34296 15162
rect 34244 15098 34296 15104
rect 34152 14952 34204 14958
rect 34152 14894 34204 14900
rect 33888 13790 34100 13818
rect 33784 11756 33836 11762
rect 33784 11698 33836 11704
rect 33704 11206 33824 11234
rect 33600 11144 33652 11150
rect 33600 11086 33652 11092
rect 33520 10662 33732 10690
rect 33600 10600 33652 10606
rect 33600 10542 33652 10548
rect 33416 10124 33468 10130
rect 33416 10066 33468 10072
rect 33048 10056 33100 10062
rect 33048 9998 33100 10004
rect 33060 9926 33088 9998
rect 33048 9920 33100 9926
rect 33048 9862 33100 9868
rect 33428 9518 33456 10066
rect 32956 9512 33008 9518
rect 32956 9454 33008 9460
rect 33416 9512 33468 9518
rect 33416 9454 33468 9460
rect 33048 9036 33100 9042
rect 33048 8978 33100 8984
rect 33060 8566 33088 8978
rect 33048 8560 33100 8566
rect 33048 8502 33100 8508
rect 32496 8424 32548 8430
rect 32496 8366 32548 8372
rect 32772 8424 32824 8430
rect 32772 8366 32824 8372
rect 32864 8424 32916 8430
rect 32864 8366 32916 8372
rect 33416 8424 33468 8430
rect 33416 8366 33468 8372
rect 32508 8090 32536 8366
rect 32496 8084 32548 8090
rect 32496 8026 32548 8032
rect 32404 7948 32456 7954
rect 32404 7890 32456 7896
rect 33324 7948 33376 7954
rect 33324 7890 33376 7896
rect 33336 7410 33364 7890
rect 33428 7478 33456 8366
rect 33416 7472 33468 7478
rect 33416 7414 33468 7420
rect 33324 7404 33376 7410
rect 33324 7346 33376 7352
rect 33232 7336 33284 7342
rect 33152 7296 33232 7324
rect 33048 6928 33100 6934
rect 33048 6870 33100 6876
rect 32312 6860 32364 6866
rect 32312 6802 32364 6808
rect 32220 6656 32272 6662
rect 32220 6598 32272 6604
rect 32324 6390 32352 6802
rect 32496 6792 32548 6798
rect 32496 6734 32548 6740
rect 32508 6390 32536 6734
rect 32312 6384 32364 6390
rect 32312 6326 32364 6332
rect 32496 6384 32548 6390
rect 32496 6326 32548 6332
rect 33060 6322 33088 6870
rect 32220 6316 32272 6322
rect 32220 6258 32272 6264
rect 33048 6316 33100 6322
rect 33048 6258 33100 6264
rect 32232 6118 32260 6258
rect 32220 6112 32272 6118
rect 32220 6054 32272 6060
rect 32048 5902 32536 5930
rect 32048 5710 32076 5902
rect 32220 5840 32272 5846
rect 32220 5782 32272 5788
rect 32036 5704 32088 5710
rect 32036 5646 32088 5652
rect 32128 5704 32180 5710
rect 32128 5646 32180 5652
rect 31944 5636 31996 5642
rect 31944 5578 31996 5584
rect 31760 5160 31812 5166
rect 31760 5102 31812 5108
rect 31772 5030 31800 5102
rect 31760 5024 31812 5030
rect 31760 4966 31812 4972
rect 30932 4820 30984 4826
rect 30932 4762 30984 4768
rect 31116 4820 31168 4826
rect 31116 4762 31168 4768
rect 31208 4820 31260 4826
rect 31208 4762 31260 4768
rect 30930 4720 30986 4729
rect 30840 4684 30892 4690
rect 30930 4655 30932 4664
rect 30840 4626 30892 4632
rect 30984 4655 30986 4664
rect 30932 4626 30984 4632
rect 30656 4616 30708 4622
rect 30656 4558 30708 4564
rect 31024 4616 31076 4622
rect 31024 4558 31076 4564
rect 30668 4214 30696 4558
rect 31036 4282 31064 4558
rect 31024 4276 31076 4282
rect 31024 4218 31076 4224
rect 30656 4208 30708 4214
rect 30656 4150 30708 4156
rect 30380 3596 30432 3602
rect 30380 3538 30432 3544
rect 31772 3534 31800 4966
rect 32140 3534 32168 5646
rect 32232 4282 32260 5782
rect 32508 5710 32536 5902
rect 32772 5772 32824 5778
rect 32772 5714 32824 5720
rect 32404 5704 32456 5710
rect 32404 5646 32456 5652
rect 32496 5704 32548 5710
rect 32496 5646 32548 5652
rect 32416 4758 32444 5646
rect 32680 5092 32732 5098
rect 32680 5034 32732 5040
rect 32404 4752 32456 4758
rect 32404 4694 32456 4700
rect 32692 4690 32720 5034
rect 32784 4826 32812 5714
rect 33152 5556 33180 7296
rect 33232 7278 33284 7284
rect 33336 6882 33364 7346
rect 33336 6854 33548 6882
rect 33612 6866 33640 10542
rect 33232 6656 33284 6662
rect 33232 6598 33284 6604
rect 32876 5528 33180 5556
rect 32876 5370 32904 5528
rect 32864 5364 32916 5370
rect 32864 5306 32916 5312
rect 32876 5166 32904 5306
rect 33244 5166 33272 6598
rect 33324 6180 33376 6186
rect 33324 6122 33376 6128
rect 32864 5160 32916 5166
rect 32864 5102 32916 5108
rect 33232 5160 33284 5166
rect 33232 5102 33284 5108
rect 32956 5024 33008 5030
rect 32956 4966 33008 4972
rect 32968 4826 32996 4966
rect 32772 4820 32824 4826
rect 32772 4762 32824 4768
rect 32956 4820 33008 4826
rect 32956 4762 33008 4768
rect 32680 4684 32732 4690
rect 32680 4626 32732 4632
rect 32404 4548 32456 4554
rect 32404 4490 32456 4496
rect 32220 4276 32272 4282
rect 32220 4218 32272 4224
rect 31760 3528 31812 3534
rect 31760 3470 31812 3476
rect 32128 3528 32180 3534
rect 32128 3470 32180 3476
rect 32232 3126 32260 4218
rect 32416 4146 32444 4490
rect 32404 4140 32456 4146
rect 32404 4082 32456 4088
rect 32680 4140 32732 4146
rect 32680 4082 32732 4088
rect 32220 3120 32272 3126
rect 32220 3062 32272 3068
rect 30380 2984 30432 2990
rect 30300 2932 30380 2938
rect 30300 2926 30432 2932
rect 27528 2916 27580 2922
rect 27528 2858 27580 2864
rect 30300 2910 30420 2926
rect 32220 2916 32272 2922
rect 30300 2514 30328 2910
rect 32220 2858 32272 2864
rect 32128 2848 32180 2854
rect 32048 2796 32128 2802
rect 32048 2790 32180 2796
rect 32048 2774 32168 2790
rect 32048 2582 32076 2774
rect 32036 2576 32088 2582
rect 32036 2518 32088 2524
rect 32232 2514 32260 2858
rect 32692 2854 32720 4082
rect 33336 3602 33364 6122
rect 33520 5370 33548 6854
rect 33600 6860 33652 6866
rect 33600 6802 33652 6808
rect 33704 6662 33732 10662
rect 33796 10130 33824 11206
rect 33888 11014 33916 13790
rect 34060 13524 34112 13530
rect 34060 13466 34112 13472
rect 34072 13326 34100 13466
rect 34060 13320 34112 13326
rect 34060 13262 34112 13268
rect 33968 12300 34020 12306
rect 33968 12242 34020 12248
rect 33980 11830 34008 12242
rect 33968 11824 34020 11830
rect 33968 11766 34020 11772
rect 33876 11008 33928 11014
rect 33876 10950 33928 10956
rect 33980 10606 34008 11766
rect 34060 11688 34112 11694
rect 34060 11630 34112 11636
rect 34072 11218 34100 11630
rect 34164 11370 34192 14894
rect 34256 13938 34284 15098
rect 34520 15020 34572 15026
rect 34520 14962 34572 14968
rect 34532 14890 34560 14962
rect 34520 14884 34572 14890
rect 34520 14826 34572 14832
rect 34532 14550 34560 14826
rect 34520 14544 34572 14550
rect 34520 14486 34572 14492
rect 34520 14408 34572 14414
rect 34520 14350 34572 14356
rect 34336 14068 34388 14074
rect 34336 14010 34388 14016
rect 34244 13932 34296 13938
rect 34244 13874 34296 13880
rect 34348 13530 34376 14010
rect 34336 13524 34388 13530
rect 34336 13466 34388 13472
rect 34336 13320 34388 13326
rect 34336 13262 34388 13268
rect 34348 12918 34376 13262
rect 34336 12912 34388 12918
rect 34336 12854 34388 12860
rect 34244 12776 34296 12782
rect 34244 12718 34296 12724
rect 34256 12170 34284 12718
rect 34244 12164 34296 12170
rect 34244 12106 34296 12112
rect 34532 11880 34560 14350
rect 34624 14346 34652 17546
rect 34940 17436 35236 17456
rect 34996 17434 35020 17436
rect 35076 17434 35100 17436
rect 35156 17434 35180 17436
rect 35018 17382 35020 17434
rect 35082 17382 35094 17434
rect 35156 17382 35158 17434
rect 34996 17380 35020 17382
rect 35076 17380 35100 17382
rect 35156 17380 35180 17382
rect 34940 17360 35236 17380
rect 34796 16992 34848 16998
rect 34796 16934 34848 16940
rect 34808 16658 34836 16934
rect 35452 16658 35480 18770
rect 35820 18698 35848 22034
rect 35900 21344 35952 21350
rect 35900 21286 35952 21292
rect 35808 18692 35860 18698
rect 35808 18634 35860 18640
rect 35532 18624 35584 18630
rect 35532 18566 35584 18572
rect 34796 16652 34848 16658
rect 35440 16652 35492 16658
rect 34796 16594 34848 16600
rect 35268 16612 35440 16640
rect 34940 16348 35236 16368
rect 34996 16346 35020 16348
rect 35076 16346 35100 16348
rect 35156 16346 35180 16348
rect 35018 16294 35020 16346
rect 35082 16294 35094 16346
rect 35156 16294 35158 16346
rect 34996 16292 35020 16294
rect 35076 16292 35100 16294
rect 35156 16292 35180 16294
rect 34940 16272 35236 16292
rect 34978 16144 35034 16153
rect 34978 16079 34980 16088
rect 35032 16079 35034 16088
rect 34980 16050 35032 16056
rect 34940 15260 35236 15280
rect 34996 15258 35020 15260
rect 35076 15258 35100 15260
rect 35156 15258 35180 15260
rect 35018 15206 35020 15258
rect 35082 15206 35094 15258
rect 35156 15206 35158 15258
rect 34996 15204 35020 15206
rect 35076 15204 35100 15206
rect 35156 15204 35180 15206
rect 34940 15184 35236 15204
rect 35268 15026 35296 16612
rect 35440 16594 35492 16600
rect 35348 15496 35400 15502
rect 35348 15438 35400 15444
rect 35256 15020 35308 15026
rect 35256 14962 35308 14968
rect 34796 14544 34848 14550
rect 34796 14486 34848 14492
rect 34704 14476 34756 14482
rect 34704 14418 34756 14424
rect 34612 14340 34664 14346
rect 34612 14282 34664 14288
rect 34612 13524 34664 13530
rect 34612 13466 34664 13472
rect 34624 12306 34652 13466
rect 34612 12300 34664 12306
rect 34612 12242 34664 12248
rect 34532 11852 34652 11880
rect 34520 11756 34572 11762
rect 34520 11698 34572 11704
rect 34164 11342 34468 11370
rect 34060 11212 34112 11218
rect 34060 11154 34112 11160
rect 33968 10600 34020 10606
rect 33968 10542 34020 10548
rect 33784 10124 33836 10130
rect 33784 10066 33836 10072
rect 34072 8022 34100 11154
rect 34244 11144 34296 11150
rect 34244 11086 34296 11092
rect 34152 10600 34204 10606
rect 34152 10542 34204 10548
rect 34164 10198 34192 10542
rect 34152 10192 34204 10198
rect 34152 10134 34204 10140
rect 34256 9654 34284 11086
rect 34334 10432 34390 10441
rect 34334 10367 34390 10376
rect 34244 9648 34296 9654
rect 34244 9590 34296 9596
rect 34150 8936 34206 8945
rect 34150 8871 34206 8880
rect 34164 8430 34192 8871
rect 34152 8424 34204 8430
rect 34152 8366 34204 8372
rect 34060 8016 34112 8022
rect 34060 7958 34112 7964
rect 34256 7954 34284 9590
rect 34348 8566 34376 10367
rect 34336 8560 34388 8566
rect 34336 8502 34388 8508
rect 33876 7948 33928 7954
rect 33876 7890 33928 7896
rect 34244 7948 34296 7954
rect 34244 7890 34296 7896
rect 33692 6656 33744 6662
rect 33692 6598 33744 6604
rect 33508 5364 33560 5370
rect 33508 5306 33560 5312
rect 33600 5160 33652 5166
rect 33600 5102 33652 5108
rect 33612 4758 33640 5102
rect 33888 4758 33916 7890
rect 34256 7410 34284 7890
rect 34244 7404 34296 7410
rect 34244 7346 34296 7352
rect 34244 6860 34296 6866
rect 34244 6802 34296 6808
rect 33968 6792 34020 6798
rect 33966 6760 33968 6769
rect 34020 6760 34022 6769
rect 33966 6695 34022 6704
rect 33600 4752 33652 4758
rect 33600 4694 33652 4700
rect 33876 4752 33928 4758
rect 33876 4694 33928 4700
rect 33888 4622 33916 4694
rect 33876 4616 33928 4622
rect 33876 4558 33928 4564
rect 33980 4486 34008 6695
rect 34152 6248 34204 6254
rect 34152 6190 34204 6196
rect 33968 4480 34020 4486
rect 33968 4422 34020 4428
rect 33980 4214 34008 4422
rect 33968 4208 34020 4214
rect 33968 4150 34020 4156
rect 33876 3936 33928 3942
rect 33876 3878 33928 3884
rect 33324 3596 33376 3602
rect 33324 3538 33376 3544
rect 32772 3528 32824 3534
rect 32772 3470 32824 3476
rect 32784 2854 32812 3470
rect 33232 3052 33284 3058
rect 33284 3012 33364 3040
rect 33232 2994 33284 3000
rect 32680 2848 32732 2854
rect 32680 2790 32732 2796
rect 32772 2848 32824 2854
rect 32772 2790 32824 2796
rect 30288 2508 30340 2514
rect 30288 2450 30340 2456
rect 32220 2508 32272 2514
rect 32220 2450 32272 2456
rect 33140 2508 33192 2514
rect 33140 2450 33192 2456
rect 26884 2440 26936 2446
rect 26884 2382 26936 2388
rect 29276 2440 29328 2446
rect 29276 2382 29328 2388
rect 27252 2304 27304 2310
rect 27252 2246 27304 2252
rect 25228 1964 25280 1970
rect 25228 1906 25280 1912
rect 25240 800 25268 1906
rect 27264 800 27292 2246
rect 29288 800 29316 2382
rect 33152 2310 33180 2450
rect 31300 2304 31352 2310
rect 31300 2246 31352 2252
rect 33140 2304 33192 2310
rect 33140 2246 33192 2252
rect 31312 800 31340 2246
rect 33152 2106 33180 2246
rect 33140 2100 33192 2106
rect 33140 2042 33192 2048
rect 33336 800 33364 3012
rect 33888 2990 33916 3878
rect 34164 2990 34192 6190
rect 34256 4078 34284 6802
rect 34440 5302 34468 11342
rect 34532 9518 34560 11698
rect 34520 9512 34572 9518
rect 34520 9454 34572 9460
rect 34532 7886 34560 9454
rect 34624 8673 34652 11852
rect 34716 11642 34744 14418
rect 34808 11762 34836 14486
rect 35360 14482 35388 15438
rect 35440 15360 35492 15366
rect 35440 15302 35492 15308
rect 35452 14958 35480 15302
rect 35544 15094 35572 18566
rect 35716 17672 35768 17678
rect 35716 17614 35768 17620
rect 35728 16182 35756 17614
rect 35716 16176 35768 16182
rect 35716 16118 35768 16124
rect 35912 16046 35940 21286
rect 36004 20058 36032 23122
rect 36096 22574 36124 23666
rect 36084 22568 36136 22574
rect 36084 22510 36136 22516
rect 36084 21480 36136 21486
rect 36084 21422 36136 21428
rect 35992 20052 36044 20058
rect 35992 19994 36044 20000
rect 36096 19922 36124 21422
rect 36084 19916 36136 19922
rect 36084 19858 36136 19864
rect 35992 18624 36044 18630
rect 35992 18566 36044 18572
rect 36004 17134 36032 18566
rect 35992 17128 36044 17134
rect 35992 17070 36044 17076
rect 36096 16998 36124 19858
rect 36188 18358 36216 33934
rect 36268 33312 36320 33318
rect 36268 33254 36320 33260
rect 36280 29073 36308 33254
rect 36372 32978 36400 34682
rect 37002 34640 37058 34649
rect 37002 34575 37058 34584
rect 37280 34604 37332 34610
rect 36452 34196 36504 34202
rect 36452 34138 36504 34144
rect 36464 33454 36492 34138
rect 37016 34066 37044 34575
rect 37280 34546 37332 34552
rect 37188 34536 37240 34542
rect 37188 34478 37240 34484
rect 37004 34060 37056 34066
rect 37004 34002 37056 34008
rect 37200 33998 37228 34478
rect 36636 33992 36688 33998
rect 36636 33934 36688 33940
rect 37188 33992 37240 33998
rect 37188 33934 37240 33940
rect 36648 33522 36676 33934
rect 37200 33658 37228 33934
rect 37188 33652 37240 33658
rect 37188 33594 37240 33600
rect 36636 33516 36688 33522
rect 36636 33458 36688 33464
rect 36452 33448 36504 33454
rect 36452 33390 36504 33396
rect 36728 33448 36780 33454
rect 36728 33390 36780 33396
rect 36740 33114 36768 33390
rect 36728 33108 36780 33114
rect 36728 33050 36780 33056
rect 37292 32978 37320 34546
rect 36360 32972 36412 32978
rect 36360 32914 36412 32920
rect 37280 32972 37332 32978
rect 37280 32914 37332 32920
rect 36636 32564 36688 32570
rect 36636 32506 36688 32512
rect 36648 31346 36676 32506
rect 38120 32434 38148 37567
rect 38304 35834 38332 39200
rect 38292 35828 38344 35834
rect 38292 35770 38344 35776
rect 38108 32428 38160 32434
rect 38108 32370 38160 32376
rect 37924 32360 37976 32366
rect 37924 32302 37976 32308
rect 37556 32224 37608 32230
rect 37556 32166 37608 32172
rect 36728 31884 36780 31890
rect 36728 31826 36780 31832
rect 37464 31884 37516 31890
rect 37464 31826 37516 31832
rect 36636 31340 36688 31346
rect 36636 31282 36688 31288
rect 36452 31272 36504 31278
rect 36452 31214 36504 31220
rect 36464 30258 36492 31214
rect 36740 30938 36768 31826
rect 37280 31816 37332 31822
rect 37280 31758 37332 31764
rect 36912 31680 36964 31686
rect 36912 31622 36964 31628
rect 36728 30932 36780 30938
rect 36728 30874 36780 30880
rect 36820 30592 36872 30598
rect 36820 30534 36872 30540
rect 36452 30252 36504 30258
rect 36452 30194 36504 30200
rect 36464 29170 36492 30194
rect 36832 29714 36860 30534
rect 36820 29708 36872 29714
rect 36820 29650 36872 29656
rect 36728 29572 36780 29578
rect 36728 29514 36780 29520
rect 36740 29170 36768 29514
rect 36820 29504 36872 29510
rect 36820 29446 36872 29452
rect 36452 29164 36504 29170
rect 36452 29106 36504 29112
rect 36728 29164 36780 29170
rect 36728 29106 36780 29112
rect 36266 29064 36322 29073
rect 36832 29050 36860 29446
rect 36266 28999 36322 29008
rect 36740 29022 36860 29050
rect 36740 28966 36768 29022
rect 36728 28960 36780 28966
rect 36728 28902 36780 28908
rect 36360 28620 36412 28626
rect 36360 28562 36412 28568
rect 36452 28620 36504 28626
rect 36452 28562 36504 28568
rect 36372 28014 36400 28562
rect 36464 28082 36492 28562
rect 36544 28552 36596 28558
rect 36544 28494 36596 28500
rect 36452 28076 36504 28082
rect 36452 28018 36504 28024
rect 36360 28008 36412 28014
rect 36360 27950 36412 27956
rect 36556 27538 36584 28494
rect 36740 28014 36768 28902
rect 36728 28008 36780 28014
rect 36728 27950 36780 27956
rect 36636 27668 36688 27674
rect 36636 27610 36688 27616
rect 36544 27532 36596 27538
rect 36544 27474 36596 27480
rect 36360 26920 36412 26926
rect 36360 26862 36412 26868
rect 36372 25838 36400 26862
rect 36360 25832 36412 25838
rect 36360 25774 36412 25780
rect 36268 24948 36320 24954
rect 36268 24890 36320 24896
rect 36280 24274 36308 24890
rect 36372 24750 36400 25774
rect 36556 25702 36584 27474
rect 36544 25696 36596 25702
rect 36544 25638 36596 25644
rect 36544 25152 36596 25158
rect 36544 25094 36596 25100
rect 36360 24744 36412 24750
rect 36556 24721 36584 25094
rect 36360 24686 36412 24692
rect 36542 24712 36598 24721
rect 36542 24647 36598 24656
rect 36556 24274 36584 24647
rect 36268 24268 36320 24274
rect 36268 24210 36320 24216
rect 36544 24268 36596 24274
rect 36544 24210 36596 24216
rect 36360 24132 36412 24138
rect 36360 24074 36412 24080
rect 36268 20528 36320 20534
rect 36268 20470 36320 20476
rect 36280 20398 36308 20470
rect 36268 20392 36320 20398
rect 36268 20334 36320 20340
rect 36280 19378 36308 20334
rect 36268 19372 36320 19378
rect 36268 19314 36320 19320
rect 36268 18760 36320 18766
rect 36268 18702 36320 18708
rect 36176 18352 36228 18358
rect 36176 18294 36228 18300
rect 36280 18222 36308 18702
rect 36268 18216 36320 18222
rect 36268 18158 36320 18164
rect 36268 18080 36320 18086
rect 36268 18022 36320 18028
rect 36280 17542 36308 18022
rect 36268 17536 36320 17542
rect 36268 17478 36320 17484
rect 36372 17490 36400 24074
rect 36452 23180 36504 23186
rect 36452 23122 36504 23128
rect 36464 22030 36492 23122
rect 36452 22024 36504 22030
rect 36452 21966 36504 21972
rect 36648 21010 36676 27610
rect 36820 26784 36872 26790
rect 36820 26726 36872 26732
rect 36832 26450 36860 26726
rect 36820 26444 36872 26450
rect 36820 26386 36872 26392
rect 36924 25378 36952 31622
rect 37188 30048 37240 30054
rect 37188 29990 37240 29996
rect 37096 29640 37148 29646
rect 37096 29582 37148 29588
rect 37108 28082 37136 29582
rect 37200 28422 37228 29990
rect 37188 28416 37240 28422
rect 37188 28358 37240 28364
rect 37096 28076 37148 28082
rect 37096 28018 37148 28024
rect 37004 27940 37056 27946
rect 37004 27882 37056 27888
rect 37016 26926 37044 27882
rect 37004 26920 37056 26926
rect 37004 26862 37056 26868
rect 37016 26790 37044 26862
rect 37004 26784 37056 26790
rect 37004 26726 37056 26732
rect 37016 26450 37044 26726
rect 37004 26444 37056 26450
rect 37004 26386 37056 26392
rect 36832 25350 36952 25378
rect 36832 24614 36860 25350
rect 37200 24750 37228 28358
rect 37188 24744 37240 24750
rect 37188 24686 37240 24692
rect 36820 24608 36872 24614
rect 36820 24550 36872 24556
rect 36832 24274 36860 24550
rect 36820 24268 36872 24274
rect 36820 24210 36872 24216
rect 36832 23730 36860 24210
rect 36820 23724 36872 23730
rect 36820 23666 36872 23672
rect 36728 23656 36780 23662
rect 36728 23598 36780 23604
rect 36740 21894 36768 23598
rect 37292 22166 37320 31758
rect 37372 30184 37424 30190
rect 37372 30126 37424 30132
rect 37384 25362 37412 30126
rect 37372 25356 37424 25362
rect 37372 25298 37424 25304
rect 37476 22778 37504 31826
rect 37568 30190 37596 32166
rect 37740 30796 37792 30802
rect 37740 30738 37792 30744
rect 37556 30184 37608 30190
rect 37556 30126 37608 30132
rect 37556 30048 37608 30054
rect 37556 29990 37608 29996
rect 37464 22772 37516 22778
rect 37464 22714 37516 22720
rect 37568 22658 37596 29990
rect 37648 29708 37700 29714
rect 37648 29650 37700 29656
rect 37660 28762 37688 29650
rect 37752 29306 37780 30738
rect 37740 29300 37792 29306
rect 37740 29242 37792 29248
rect 37648 28756 37700 28762
rect 37648 28698 37700 28704
rect 37752 28642 37780 29242
rect 37936 29034 37964 32302
rect 37924 29028 37976 29034
rect 37924 28970 37976 28976
rect 38016 28960 38068 28966
rect 38016 28902 38068 28908
rect 37660 28626 37780 28642
rect 37648 28620 37780 28626
rect 37700 28614 37780 28620
rect 37648 28562 37700 28568
rect 37922 28384 37978 28393
rect 37922 28319 37978 28328
rect 37936 28218 37964 28319
rect 37924 28212 37976 28218
rect 37924 28154 37976 28160
rect 37740 27532 37792 27538
rect 37740 27474 37792 27480
rect 37752 26314 37780 27474
rect 37832 27328 37884 27334
rect 37832 27270 37884 27276
rect 37844 26994 37872 27270
rect 37832 26988 37884 26994
rect 37832 26930 37884 26936
rect 37740 26308 37792 26314
rect 37740 26250 37792 26256
rect 38028 24954 38056 28902
rect 38016 24948 38068 24954
rect 38016 24890 38068 24896
rect 37832 24744 37884 24750
rect 37832 24686 37884 24692
rect 37844 24410 37872 24686
rect 38016 24676 38068 24682
rect 38016 24618 38068 24624
rect 37832 24404 37884 24410
rect 37832 24346 37884 24352
rect 37832 23520 37884 23526
rect 37832 23462 37884 23468
rect 37844 23186 37872 23462
rect 37832 23180 37884 23186
rect 37832 23122 37884 23128
rect 37476 22630 37596 22658
rect 37280 22160 37332 22166
rect 37280 22102 37332 22108
rect 36728 21888 36780 21894
rect 36728 21830 36780 21836
rect 37004 21888 37056 21894
rect 37004 21830 37056 21836
rect 37016 21690 37044 21830
rect 37004 21684 37056 21690
rect 37004 21626 37056 21632
rect 37292 21554 37320 22102
rect 37280 21548 37332 21554
rect 37280 21490 37332 21496
rect 37372 21344 37424 21350
rect 37372 21286 37424 21292
rect 36636 21004 36688 21010
rect 36636 20946 36688 20952
rect 37004 21004 37056 21010
rect 37004 20946 37056 20952
rect 36820 20936 36872 20942
rect 36820 20878 36872 20884
rect 36832 19922 36860 20878
rect 36820 19916 36872 19922
rect 36820 19858 36872 19864
rect 36728 19780 36780 19786
rect 36728 19722 36780 19728
rect 36912 19780 36964 19786
rect 36912 19722 36964 19728
rect 36544 19304 36596 19310
rect 36544 19246 36596 19252
rect 36452 18828 36504 18834
rect 36452 18770 36504 18776
rect 36464 18426 36492 18770
rect 36452 18420 36504 18426
rect 36452 18362 36504 18368
rect 36556 18222 36584 19246
rect 36740 18290 36768 19722
rect 36728 18284 36780 18290
rect 36728 18226 36780 18232
rect 36544 18216 36596 18222
rect 36544 18158 36596 18164
rect 36280 17134 36308 17478
rect 36372 17462 36768 17490
rect 36268 17128 36320 17134
rect 36268 17070 36320 17076
rect 36084 16992 36136 16998
rect 36084 16934 36136 16940
rect 35992 16788 36044 16794
rect 35992 16730 36044 16736
rect 36004 16114 36032 16730
rect 35992 16108 36044 16114
rect 35992 16050 36044 16056
rect 35900 16040 35952 16046
rect 35900 15982 35952 15988
rect 35912 15706 35940 15982
rect 35900 15700 35952 15706
rect 35900 15642 35952 15648
rect 35716 15564 35768 15570
rect 35716 15506 35768 15512
rect 35532 15088 35584 15094
rect 35532 15030 35584 15036
rect 35440 14952 35492 14958
rect 35440 14894 35492 14900
rect 35532 14952 35584 14958
rect 35532 14894 35584 14900
rect 35452 14550 35480 14894
rect 35440 14544 35492 14550
rect 35440 14486 35492 14492
rect 35348 14476 35400 14482
rect 35348 14418 35400 14424
rect 34940 14172 35236 14192
rect 34996 14170 35020 14172
rect 35076 14170 35100 14172
rect 35156 14170 35180 14172
rect 35018 14118 35020 14170
rect 35082 14118 35094 14170
rect 35156 14118 35158 14170
rect 34996 14116 35020 14118
rect 35076 14116 35100 14118
rect 35156 14116 35180 14118
rect 34940 14096 35236 14116
rect 35360 13530 35388 14418
rect 35440 13932 35492 13938
rect 35440 13874 35492 13880
rect 35348 13524 35400 13530
rect 35348 13466 35400 13472
rect 35254 13424 35310 13433
rect 35254 13359 35310 13368
rect 34940 13084 35236 13104
rect 34996 13082 35020 13084
rect 35076 13082 35100 13084
rect 35156 13082 35180 13084
rect 35018 13030 35020 13082
rect 35082 13030 35094 13082
rect 35156 13030 35158 13082
rect 34996 13028 35020 13030
rect 35076 13028 35100 13030
rect 35156 13028 35180 13030
rect 34940 13008 35236 13028
rect 35268 12782 35296 13359
rect 35452 12850 35480 13874
rect 35544 13190 35572 14894
rect 35728 14414 35756 15506
rect 35992 15020 36044 15026
rect 35992 14962 36044 14968
rect 35716 14408 35768 14414
rect 35716 14350 35768 14356
rect 36004 13870 36032 14962
rect 36280 14958 36308 17070
rect 36544 17060 36596 17066
rect 36544 17002 36596 17008
rect 36556 16250 36584 17002
rect 36544 16244 36596 16250
rect 36544 16186 36596 16192
rect 36636 15564 36688 15570
rect 36636 15506 36688 15512
rect 36268 14952 36320 14958
rect 36268 14894 36320 14900
rect 36452 14952 36504 14958
rect 36452 14894 36504 14900
rect 36268 14476 36320 14482
rect 36268 14418 36320 14424
rect 36084 14068 36136 14074
rect 36084 14010 36136 14016
rect 35992 13864 36044 13870
rect 35992 13806 36044 13812
rect 35532 13184 35584 13190
rect 35532 13126 35584 13132
rect 35440 12844 35492 12850
rect 35440 12786 35492 12792
rect 35256 12776 35308 12782
rect 35256 12718 35308 12724
rect 35544 12628 35572 13126
rect 36096 12782 36124 14010
rect 36280 14006 36308 14418
rect 36464 14074 36492 14894
rect 36648 14482 36676 15506
rect 36636 14476 36688 14482
rect 36636 14418 36688 14424
rect 36452 14068 36504 14074
rect 36452 14010 36504 14016
rect 36268 14000 36320 14006
rect 36268 13942 36320 13948
rect 36464 13870 36492 14010
rect 36452 13864 36504 13870
rect 36452 13806 36504 13812
rect 36544 13864 36596 13870
rect 36544 13806 36596 13812
rect 36176 13320 36228 13326
rect 36176 13262 36228 13268
rect 36268 13320 36320 13326
rect 36268 13262 36320 13268
rect 36084 12776 36136 12782
rect 36084 12718 36136 12724
rect 35268 12600 35572 12628
rect 34940 11996 35236 12016
rect 34996 11994 35020 11996
rect 35076 11994 35100 11996
rect 35156 11994 35180 11996
rect 35018 11942 35020 11994
rect 35082 11942 35094 11994
rect 35156 11942 35158 11994
rect 34996 11940 35020 11942
rect 35076 11940 35100 11942
rect 35156 11940 35180 11942
rect 34940 11920 35236 11940
rect 34796 11756 34848 11762
rect 34796 11698 34848 11704
rect 34716 11614 34836 11642
rect 34704 10464 34756 10470
rect 34704 10406 34756 10412
rect 34716 10130 34744 10406
rect 34808 10146 34836 11614
rect 34940 10908 35236 10928
rect 34996 10906 35020 10908
rect 35076 10906 35100 10908
rect 35156 10906 35180 10908
rect 35018 10854 35020 10906
rect 35082 10854 35094 10906
rect 35156 10854 35158 10906
rect 34996 10852 35020 10854
rect 35076 10852 35100 10854
rect 35156 10852 35180 10854
rect 34940 10832 35236 10852
rect 34704 10124 34756 10130
rect 34808 10118 34928 10146
rect 34704 10066 34756 10072
rect 34796 10056 34848 10062
rect 34716 10004 34796 10010
rect 34716 9998 34848 10004
rect 34716 9982 34836 9998
rect 34716 8974 34744 9982
rect 34900 9908 34928 10118
rect 34808 9880 34928 9908
rect 34704 8968 34756 8974
rect 34704 8910 34756 8916
rect 34610 8664 34666 8673
rect 34610 8599 34666 8608
rect 34520 7880 34572 7886
rect 34520 7822 34572 7828
rect 34520 6792 34572 6798
rect 34520 6734 34572 6740
rect 34704 6792 34756 6798
rect 34704 6734 34756 6740
rect 34532 6390 34560 6734
rect 34520 6384 34572 6390
rect 34520 6326 34572 6332
rect 34520 6248 34572 6254
rect 34520 6190 34572 6196
rect 34428 5296 34480 5302
rect 34428 5238 34480 5244
rect 34532 5148 34560 6190
rect 34716 5778 34744 6734
rect 34808 6361 34836 9880
rect 34940 9820 35236 9840
rect 34996 9818 35020 9820
rect 35076 9818 35100 9820
rect 35156 9818 35180 9820
rect 35018 9766 35020 9818
rect 35082 9766 35094 9818
rect 35156 9766 35158 9818
rect 34996 9764 35020 9766
rect 35076 9764 35100 9766
rect 35156 9764 35180 9766
rect 34940 9744 35236 9764
rect 34940 8732 35236 8752
rect 34996 8730 35020 8732
rect 35076 8730 35100 8732
rect 35156 8730 35180 8732
rect 35018 8678 35020 8730
rect 35082 8678 35094 8730
rect 35156 8678 35158 8730
rect 34996 8676 35020 8678
rect 35076 8676 35100 8678
rect 35156 8676 35180 8678
rect 34940 8656 35236 8676
rect 35268 8362 35296 12600
rect 35440 12232 35492 12238
rect 35440 12174 35492 12180
rect 35348 12096 35400 12102
rect 35348 12038 35400 12044
rect 35360 11150 35388 12038
rect 35348 11144 35400 11150
rect 35348 11086 35400 11092
rect 35360 10062 35388 11086
rect 35348 10056 35400 10062
rect 35348 9998 35400 10004
rect 35348 9444 35400 9450
rect 35348 9386 35400 9392
rect 35256 8356 35308 8362
rect 35256 8298 35308 8304
rect 35268 7954 35296 8298
rect 35256 7948 35308 7954
rect 35256 7890 35308 7896
rect 34940 7644 35236 7664
rect 34996 7642 35020 7644
rect 35076 7642 35100 7644
rect 35156 7642 35180 7644
rect 35018 7590 35020 7642
rect 35082 7590 35094 7642
rect 35156 7590 35158 7642
rect 34996 7588 35020 7590
rect 35076 7588 35100 7590
rect 35156 7588 35180 7590
rect 34940 7568 35236 7588
rect 35360 7410 35388 9386
rect 35452 9110 35480 12174
rect 35808 11688 35860 11694
rect 35808 11630 35860 11636
rect 35716 11144 35768 11150
rect 35716 11086 35768 11092
rect 35532 9512 35584 9518
rect 35532 9454 35584 9460
rect 35624 9512 35676 9518
rect 35624 9454 35676 9460
rect 35440 9104 35492 9110
rect 35440 9046 35492 9052
rect 35440 8968 35492 8974
rect 35440 8910 35492 8916
rect 35452 8634 35480 8910
rect 35544 8838 35572 9454
rect 35532 8832 35584 8838
rect 35532 8774 35584 8780
rect 35440 8628 35492 8634
rect 35440 8570 35492 8576
rect 35544 8430 35572 8774
rect 35636 8430 35664 9454
rect 35532 8424 35584 8430
rect 35532 8366 35584 8372
rect 35624 8424 35676 8430
rect 35624 8366 35676 8372
rect 35440 7948 35492 7954
rect 35440 7890 35492 7896
rect 35452 7546 35480 7890
rect 35440 7540 35492 7546
rect 35440 7482 35492 7488
rect 35348 7404 35400 7410
rect 35348 7346 35400 7352
rect 35440 6792 35492 6798
rect 35440 6734 35492 6740
rect 34940 6556 35236 6576
rect 34996 6554 35020 6556
rect 35076 6554 35100 6556
rect 35156 6554 35180 6556
rect 35018 6502 35020 6554
rect 35082 6502 35094 6554
rect 35156 6502 35158 6554
rect 34996 6500 35020 6502
rect 35076 6500 35100 6502
rect 35156 6500 35180 6502
rect 34940 6480 35236 6500
rect 34794 6352 34850 6361
rect 35452 6322 35480 6734
rect 34794 6287 34850 6296
rect 35440 6316 35492 6322
rect 35440 6258 35492 6264
rect 35544 6254 35572 8366
rect 35636 7188 35664 8366
rect 35728 7342 35756 11086
rect 35820 10266 35848 11630
rect 35900 11008 35952 11014
rect 35900 10950 35952 10956
rect 35912 10674 35940 10950
rect 35900 10668 35952 10674
rect 35900 10610 35952 10616
rect 36084 10532 36136 10538
rect 36084 10474 36136 10480
rect 35808 10260 35860 10266
rect 35808 10202 35860 10208
rect 35820 10062 35848 10202
rect 35808 10056 35860 10062
rect 35808 9998 35860 10004
rect 35820 9518 35848 9998
rect 35808 9512 35860 9518
rect 35808 9454 35860 9460
rect 35992 9512 36044 9518
rect 35992 9454 36044 9460
rect 35900 8968 35952 8974
rect 35900 8910 35952 8916
rect 35912 8498 35940 8910
rect 36004 8634 36032 9454
rect 36096 8634 36124 10474
rect 35992 8628 36044 8634
rect 35992 8570 36044 8576
rect 36084 8628 36136 8634
rect 36084 8570 36136 8576
rect 35900 8492 35952 8498
rect 35900 8434 35952 8440
rect 36004 8430 36032 8570
rect 35992 8424 36044 8430
rect 35992 8366 36044 8372
rect 36096 7342 36124 8570
rect 36188 7478 36216 13262
rect 36280 9382 36308 13262
rect 36556 12850 36584 13806
rect 36544 12844 36596 12850
rect 36544 12786 36596 12792
rect 36452 11688 36504 11694
rect 36452 11630 36504 11636
rect 36464 10674 36492 11630
rect 36452 10668 36504 10674
rect 36452 10610 36504 10616
rect 36268 9376 36320 9382
rect 36268 9318 36320 9324
rect 36360 8968 36412 8974
rect 36360 8910 36412 8916
rect 36268 8424 36320 8430
rect 36268 8366 36320 8372
rect 36176 7472 36228 7478
rect 36176 7414 36228 7420
rect 35716 7336 35768 7342
rect 35716 7278 35768 7284
rect 36084 7336 36136 7342
rect 36084 7278 36136 7284
rect 36176 7336 36228 7342
rect 36280 7324 36308 8366
rect 36372 7410 36400 8910
rect 36360 7404 36412 7410
rect 36360 7346 36412 7352
rect 36228 7296 36308 7324
rect 36176 7278 36228 7284
rect 35636 7160 35940 7188
rect 35808 6860 35860 6866
rect 35808 6802 35860 6808
rect 35912 6848 35940 7160
rect 35992 6860 36044 6866
rect 35912 6820 35992 6848
rect 35716 6384 35768 6390
rect 35622 6352 35678 6361
rect 35716 6326 35768 6332
rect 35622 6287 35678 6296
rect 35636 6254 35664 6287
rect 35532 6248 35584 6254
rect 35532 6190 35584 6196
rect 35624 6248 35676 6254
rect 35624 6190 35676 6196
rect 35624 6112 35676 6118
rect 35624 6054 35676 6060
rect 34704 5772 34756 5778
rect 34704 5714 34756 5720
rect 34940 5468 35236 5488
rect 34996 5466 35020 5468
rect 35076 5466 35100 5468
rect 35156 5466 35180 5468
rect 35018 5414 35020 5466
rect 35082 5414 35094 5466
rect 35156 5414 35158 5466
rect 34996 5412 35020 5414
rect 35076 5412 35100 5414
rect 35156 5412 35180 5414
rect 34940 5392 35236 5412
rect 34440 5120 34560 5148
rect 34440 4554 34468 5120
rect 34612 4684 34664 4690
rect 34612 4626 34664 4632
rect 35440 4684 35492 4690
rect 35440 4626 35492 4632
rect 34520 4616 34572 4622
rect 34520 4558 34572 4564
rect 34428 4548 34480 4554
rect 34428 4490 34480 4496
rect 34336 4140 34388 4146
rect 34336 4082 34388 4088
rect 34244 4072 34296 4078
rect 34244 4014 34296 4020
rect 34348 3058 34376 4082
rect 34532 3670 34560 4558
rect 34624 3942 34652 4626
rect 35452 4486 35480 4626
rect 35532 4616 35584 4622
rect 35532 4558 35584 4564
rect 35440 4480 35492 4486
rect 35440 4422 35492 4428
rect 34940 4380 35236 4400
rect 34996 4378 35020 4380
rect 35076 4378 35100 4380
rect 35156 4378 35180 4380
rect 35018 4326 35020 4378
rect 35082 4326 35094 4378
rect 35156 4326 35158 4378
rect 34996 4324 35020 4326
rect 35076 4324 35100 4326
rect 35156 4324 35180 4326
rect 34940 4304 35236 4324
rect 34794 4176 34850 4185
rect 34794 4111 34850 4120
rect 34612 3936 34664 3942
rect 34612 3878 34664 3884
rect 34520 3664 34572 3670
rect 34520 3606 34572 3612
rect 34428 3528 34480 3534
rect 34428 3470 34480 3476
rect 34336 3052 34388 3058
rect 34336 2994 34388 3000
rect 33876 2984 33928 2990
rect 33876 2926 33928 2932
rect 34152 2984 34204 2990
rect 34152 2926 34204 2932
rect 34440 2582 34468 3470
rect 34532 2990 34560 3606
rect 34704 3528 34756 3534
rect 34704 3470 34756 3476
rect 34520 2984 34572 2990
rect 34520 2926 34572 2932
rect 34716 2854 34744 3470
rect 34808 3466 34836 4111
rect 35440 4004 35492 4010
rect 35440 3946 35492 3952
rect 34796 3460 34848 3466
rect 34796 3402 34848 3408
rect 34940 3292 35236 3312
rect 34996 3290 35020 3292
rect 35076 3290 35100 3292
rect 35156 3290 35180 3292
rect 35018 3238 35020 3290
rect 35082 3238 35094 3290
rect 35156 3238 35158 3290
rect 34996 3236 35020 3238
rect 35076 3236 35100 3238
rect 35156 3236 35180 3238
rect 34940 3216 35236 3236
rect 35452 3058 35480 3946
rect 35440 3052 35492 3058
rect 35440 2994 35492 3000
rect 34704 2848 34756 2854
rect 34704 2790 34756 2796
rect 34428 2576 34480 2582
rect 34428 2518 34480 2524
rect 35544 2514 35572 4558
rect 35636 4010 35664 6054
rect 35728 5166 35756 6326
rect 35820 5778 35848 6802
rect 35912 6322 35940 6820
rect 35992 6802 36044 6808
rect 35900 6316 35952 6322
rect 35900 6258 35952 6264
rect 35808 5772 35860 5778
rect 35808 5714 35860 5720
rect 35820 5234 35848 5714
rect 35808 5228 35860 5234
rect 35808 5170 35860 5176
rect 35716 5160 35768 5166
rect 35716 5102 35768 5108
rect 35728 4146 35756 5102
rect 35716 4140 35768 4146
rect 35716 4082 35768 4088
rect 35912 4078 35940 6258
rect 36084 6248 36136 6254
rect 36084 6190 36136 6196
rect 36096 5846 36124 6190
rect 36084 5840 36136 5846
rect 36084 5782 36136 5788
rect 36084 5568 36136 5574
rect 36188 5556 36216 7278
rect 36372 7002 36400 7346
rect 36360 6996 36412 7002
rect 36360 6938 36412 6944
rect 36136 5528 36216 5556
rect 36084 5510 36136 5516
rect 36096 5166 36124 5510
rect 36084 5160 36136 5166
rect 36084 5102 36136 5108
rect 36096 4078 36124 5102
rect 35900 4072 35952 4078
rect 35900 4014 35952 4020
rect 36084 4072 36136 4078
rect 36084 4014 36136 4020
rect 35624 4004 35676 4010
rect 35624 3946 35676 3952
rect 36096 3534 36124 4014
rect 36084 3528 36136 3534
rect 36084 3470 36136 3476
rect 36464 2990 36492 10610
rect 36648 10266 36676 14418
rect 36740 12782 36768 17462
rect 36924 15638 36952 19722
rect 37016 19718 37044 20946
rect 37280 19916 37332 19922
rect 37280 19858 37332 19864
rect 37004 19712 37056 19718
rect 37004 19654 37056 19660
rect 37016 18834 37044 19654
rect 37004 18828 37056 18834
rect 37004 18770 37056 18776
rect 37292 17814 37320 19858
rect 37384 19310 37412 21286
rect 37372 19304 37424 19310
rect 37372 19246 37424 19252
rect 37280 17808 37332 17814
rect 37280 17750 37332 17756
rect 37292 16114 37320 17750
rect 37280 16108 37332 16114
rect 37280 16050 37332 16056
rect 37188 16040 37240 16046
rect 37188 15982 37240 15988
rect 37004 15904 37056 15910
rect 37004 15846 37056 15852
rect 36912 15632 36964 15638
rect 36912 15574 36964 15580
rect 36820 12980 36872 12986
rect 36820 12922 36872 12928
rect 36728 12776 36780 12782
rect 36728 12718 36780 12724
rect 36728 11688 36780 11694
rect 36728 11630 36780 11636
rect 36740 10305 36768 11630
rect 36726 10296 36782 10305
rect 36636 10260 36688 10266
rect 36726 10231 36782 10240
rect 36636 10202 36688 10208
rect 36832 9042 36860 12922
rect 37016 11354 37044 15846
rect 37200 14346 37228 15982
rect 37292 15570 37320 16050
rect 37372 15972 37424 15978
rect 37372 15914 37424 15920
rect 37280 15564 37332 15570
rect 37280 15506 37332 15512
rect 37384 15502 37412 15914
rect 37372 15496 37424 15502
rect 37372 15438 37424 15444
rect 37384 15162 37412 15438
rect 37372 15156 37424 15162
rect 37372 15098 37424 15104
rect 37188 14340 37240 14346
rect 37188 14282 37240 14288
rect 37188 13320 37240 13326
rect 37188 13262 37240 13268
rect 37004 11348 37056 11354
rect 37004 11290 37056 11296
rect 37016 10130 37044 11290
rect 37200 10470 37228 13262
rect 37280 12232 37332 12238
rect 37278 12200 37280 12209
rect 37332 12200 37334 12209
rect 37278 12135 37334 12144
rect 37476 11898 37504 22630
rect 37648 22092 37700 22098
rect 37648 22034 37700 22040
rect 37660 21486 37688 22034
rect 37648 21480 37700 21486
rect 37648 21422 37700 21428
rect 37832 21480 37884 21486
rect 37832 21422 37884 21428
rect 37556 21072 37608 21078
rect 37556 21014 37608 21020
rect 37568 18358 37596 21014
rect 37660 20602 37688 21422
rect 37648 20596 37700 20602
rect 37648 20538 37700 20544
rect 37844 20398 37872 21422
rect 37832 20392 37884 20398
rect 37832 20334 37884 20340
rect 37922 19408 37978 19417
rect 37922 19343 37978 19352
rect 37740 18420 37792 18426
rect 37740 18362 37792 18368
rect 37556 18352 37608 18358
rect 37556 18294 37608 18300
rect 37752 17202 37780 18362
rect 37832 17536 37884 17542
rect 37832 17478 37884 17484
rect 37844 17338 37872 17478
rect 37832 17332 37884 17338
rect 37832 17274 37884 17280
rect 37740 17196 37792 17202
rect 37740 17138 37792 17144
rect 37936 16538 37964 19343
rect 37844 16510 37964 16538
rect 37740 13388 37792 13394
rect 37740 13330 37792 13336
rect 37556 12640 37608 12646
rect 37556 12582 37608 12588
rect 37464 11892 37516 11898
rect 37464 11834 37516 11840
rect 37568 10577 37596 12582
rect 37752 12306 37780 13330
rect 37740 12300 37792 12306
rect 37740 12242 37792 12248
rect 37844 11898 37872 16510
rect 37924 16448 37976 16454
rect 37922 16416 37924 16425
rect 37976 16416 37978 16425
rect 37922 16351 37978 16360
rect 37832 11892 37884 11898
rect 37832 11834 37884 11840
rect 37554 10568 37610 10577
rect 37554 10503 37610 10512
rect 37188 10464 37240 10470
rect 37188 10406 37240 10412
rect 37004 10124 37056 10130
rect 37004 10066 37056 10072
rect 36820 9036 36872 9042
rect 36820 8978 36872 8984
rect 37372 6792 37424 6798
rect 37372 6734 37424 6740
rect 37004 6248 37056 6254
rect 37004 6190 37056 6196
rect 37280 6248 37332 6254
rect 37280 6190 37332 6196
rect 36636 5908 36688 5914
rect 36636 5850 36688 5856
rect 36648 5234 36676 5850
rect 36728 5772 36780 5778
rect 36728 5714 36780 5720
rect 36636 5228 36688 5234
rect 36636 5170 36688 5176
rect 36542 4720 36598 4729
rect 36740 4706 36768 5714
rect 36598 4678 36768 4706
rect 36542 4655 36544 4664
rect 36596 4655 36598 4664
rect 36544 4626 36596 4632
rect 37016 4486 37044 6190
rect 37292 4758 37320 6190
rect 37384 5370 37412 6734
rect 37568 6254 37596 10503
rect 37740 10124 37792 10130
rect 37740 10066 37792 10072
rect 37752 9625 37780 10066
rect 37738 9616 37794 9625
rect 37738 9551 37794 9560
rect 38028 9518 38056 24618
rect 38120 16658 38148 32370
rect 38108 16652 38160 16658
rect 38108 16594 38160 16600
rect 38108 10532 38160 10538
rect 38108 10474 38160 10480
rect 38016 9512 38068 9518
rect 38016 9454 38068 9460
rect 37832 8900 37884 8906
rect 37832 8842 37884 8848
rect 37844 7546 37872 8842
rect 37832 7540 37884 7546
rect 37832 7482 37884 7488
rect 38120 7177 38148 10474
rect 38106 7168 38162 7177
rect 38106 7103 38162 7112
rect 37740 6452 37792 6458
rect 37740 6394 37792 6400
rect 37464 6248 37516 6254
rect 37464 6190 37516 6196
rect 37556 6248 37608 6254
rect 37556 6190 37608 6196
rect 37372 5364 37424 5370
rect 37372 5306 37424 5312
rect 37280 4752 37332 4758
rect 37280 4694 37332 4700
rect 37004 4480 37056 4486
rect 37004 4422 37056 4428
rect 37292 4282 37320 4694
rect 37280 4276 37332 4282
rect 37280 4218 37332 4224
rect 37292 3738 37320 4218
rect 37280 3732 37332 3738
rect 37280 3674 37332 3680
rect 37476 3670 37504 6190
rect 37464 3664 37516 3670
rect 37464 3606 37516 3612
rect 36452 2984 36504 2990
rect 36452 2926 36504 2932
rect 36268 2916 36320 2922
rect 36268 2858 36320 2864
rect 36280 2650 36308 2858
rect 36268 2644 36320 2650
rect 36268 2586 36320 2592
rect 35532 2508 35584 2514
rect 35532 2450 35584 2456
rect 36360 2440 36412 2446
rect 36464 2428 36492 2926
rect 37476 2514 37504 3606
rect 37568 3602 37596 6190
rect 37752 4690 37780 6394
rect 37922 5672 37978 5681
rect 37922 5607 37924 5616
rect 37976 5607 37978 5616
rect 37924 5578 37976 5584
rect 37740 4684 37792 4690
rect 37740 4626 37792 4632
rect 37924 4480 37976 4486
rect 37924 4422 37976 4428
rect 37556 3596 37608 3602
rect 37556 3538 37608 3544
rect 37936 2650 37964 4422
rect 38108 2916 38160 2922
rect 38108 2858 38160 2864
rect 37924 2644 37976 2650
rect 37924 2586 37976 2592
rect 37464 2508 37516 2514
rect 37464 2450 37516 2456
rect 36412 2400 36492 2428
rect 36360 2382 36412 2388
rect 35348 2304 35400 2310
rect 35348 2246 35400 2252
rect 37556 2304 37608 2310
rect 37556 2246 37608 2252
rect 34940 2204 35236 2224
rect 34996 2202 35020 2204
rect 35076 2202 35100 2204
rect 35156 2202 35180 2204
rect 35018 2150 35020 2202
rect 35082 2150 35094 2202
rect 35156 2150 35158 2202
rect 34996 2148 35020 2150
rect 35076 2148 35100 2150
rect 35156 2148 35180 2150
rect 34940 2128 35236 2148
rect 35360 800 35388 2246
rect 37568 800 37596 2246
rect 38120 1193 38148 2858
rect 38106 1184 38162 1193
rect 38106 1119 38162 1128
rect 570 0 626 800
rect 2594 0 2650 800
rect 4618 0 4674 800
rect 6642 0 6698 800
rect 8666 0 8722 800
rect 10690 0 10746 800
rect 12898 0 12954 800
rect 14922 0 14978 800
rect 16946 0 17002 800
rect 18970 0 19026 800
rect 20994 0 21050 800
rect 23018 0 23074 800
rect 25226 0 25282 800
rect 27250 0 27306 800
rect 29274 0 29330 800
rect 31298 0 31354 800
rect 33322 0 33378 800
rect 35346 0 35402 800
rect 37554 0 37610 800
<< via2 >>
rect 2778 37304 2834 37360
rect 4220 37018 4276 37020
rect 4300 37018 4356 37020
rect 4380 37018 4436 37020
rect 4460 37018 4516 37020
rect 4220 36966 4246 37018
rect 4246 36966 4276 37018
rect 4300 36966 4310 37018
rect 4310 36966 4356 37018
rect 4380 36966 4426 37018
rect 4426 36966 4436 37018
rect 4460 36966 4490 37018
rect 4490 36966 4516 37018
rect 4220 36964 4276 36966
rect 4300 36964 4356 36966
rect 4380 36964 4436 36966
rect 4460 36964 4516 36966
rect 4220 35930 4276 35932
rect 4300 35930 4356 35932
rect 4380 35930 4436 35932
rect 4460 35930 4516 35932
rect 4220 35878 4246 35930
rect 4246 35878 4276 35930
rect 4300 35878 4310 35930
rect 4310 35878 4356 35930
rect 4380 35878 4426 35930
rect 4426 35878 4436 35930
rect 4460 35878 4490 35930
rect 4490 35878 4516 35930
rect 4220 35876 4276 35878
rect 4300 35876 4356 35878
rect 4380 35876 4436 35878
rect 4460 35876 4516 35878
rect 3790 34040 3846 34096
rect 2134 31220 2136 31240
rect 2136 31220 2188 31240
rect 2188 31220 2190 31240
rect 2134 31184 2190 31220
rect 3146 31184 3202 31240
rect 1950 31048 2006 31104
rect 3054 28056 3110 28112
rect 570 3440 626 3496
rect 2778 22072 2834 22128
rect 3422 21972 3424 21992
rect 3424 21972 3476 21992
rect 3476 21972 3478 21992
rect 3422 21936 3478 21972
rect 4220 34842 4276 34844
rect 4300 34842 4356 34844
rect 4380 34842 4436 34844
rect 4460 34842 4516 34844
rect 4220 34790 4246 34842
rect 4246 34790 4276 34842
rect 4300 34790 4310 34842
rect 4310 34790 4356 34842
rect 4380 34790 4426 34842
rect 4426 34790 4436 34842
rect 4460 34790 4490 34842
rect 4490 34790 4516 34842
rect 4220 34788 4276 34790
rect 4300 34788 4356 34790
rect 4380 34788 4436 34790
rect 4460 34788 4516 34790
rect 4220 33754 4276 33756
rect 4300 33754 4356 33756
rect 4380 33754 4436 33756
rect 4460 33754 4516 33756
rect 4220 33702 4246 33754
rect 4246 33702 4276 33754
rect 4300 33702 4310 33754
rect 4310 33702 4356 33754
rect 4380 33702 4426 33754
rect 4426 33702 4436 33754
rect 4460 33702 4490 33754
rect 4490 33702 4516 33754
rect 4220 33700 4276 33702
rect 4300 33700 4356 33702
rect 4380 33700 4436 33702
rect 4460 33700 4516 33702
rect 4220 32666 4276 32668
rect 4300 32666 4356 32668
rect 4380 32666 4436 32668
rect 4460 32666 4516 32668
rect 4220 32614 4246 32666
rect 4246 32614 4276 32666
rect 4300 32614 4310 32666
rect 4310 32614 4356 32666
rect 4380 32614 4426 32666
rect 4426 32614 4436 32666
rect 4460 32614 4490 32666
rect 4490 32614 4516 32666
rect 4220 32612 4276 32614
rect 4300 32612 4356 32614
rect 4380 32612 4436 32614
rect 4460 32612 4516 32614
rect 4220 31578 4276 31580
rect 4300 31578 4356 31580
rect 4380 31578 4436 31580
rect 4460 31578 4516 31580
rect 4220 31526 4246 31578
rect 4246 31526 4276 31578
rect 4300 31526 4310 31578
rect 4310 31526 4356 31578
rect 4380 31526 4426 31578
rect 4426 31526 4436 31578
rect 4460 31526 4490 31578
rect 4490 31526 4516 31578
rect 4220 31524 4276 31526
rect 4300 31524 4356 31526
rect 4380 31524 4436 31526
rect 4460 31524 4516 31526
rect 4434 31220 4436 31240
rect 4436 31220 4488 31240
rect 4488 31220 4490 31240
rect 4434 31184 4490 31220
rect 4220 30490 4276 30492
rect 4300 30490 4356 30492
rect 4380 30490 4436 30492
rect 4460 30490 4516 30492
rect 4220 30438 4246 30490
rect 4246 30438 4276 30490
rect 4300 30438 4310 30490
rect 4310 30438 4356 30490
rect 4380 30438 4426 30490
rect 4426 30438 4436 30490
rect 4460 30438 4490 30490
rect 4490 30438 4516 30490
rect 4220 30436 4276 30438
rect 4300 30436 4356 30438
rect 4380 30436 4436 30438
rect 4460 30436 4516 30438
rect 4220 29402 4276 29404
rect 4300 29402 4356 29404
rect 4380 29402 4436 29404
rect 4460 29402 4516 29404
rect 4220 29350 4246 29402
rect 4246 29350 4276 29402
rect 4300 29350 4310 29402
rect 4310 29350 4356 29402
rect 4380 29350 4426 29402
rect 4426 29350 4436 29402
rect 4460 29350 4490 29402
rect 4490 29350 4516 29402
rect 4220 29348 4276 29350
rect 4300 29348 4356 29350
rect 4380 29348 4436 29350
rect 4460 29348 4516 29350
rect 4220 28314 4276 28316
rect 4300 28314 4356 28316
rect 4380 28314 4436 28316
rect 4460 28314 4516 28316
rect 4220 28262 4246 28314
rect 4246 28262 4276 28314
rect 4300 28262 4310 28314
rect 4310 28262 4356 28314
rect 4380 28262 4426 28314
rect 4426 28262 4436 28314
rect 4460 28262 4490 28314
rect 4490 28262 4516 28314
rect 4220 28260 4276 28262
rect 4300 28260 4356 28262
rect 4380 28260 4436 28262
rect 4460 28260 4516 28262
rect 4220 27226 4276 27228
rect 4300 27226 4356 27228
rect 4380 27226 4436 27228
rect 4460 27226 4516 27228
rect 4220 27174 4246 27226
rect 4246 27174 4276 27226
rect 4300 27174 4310 27226
rect 4310 27174 4356 27226
rect 4380 27174 4426 27226
rect 4426 27174 4436 27226
rect 4460 27174 4490 27226
rect 4490 27174 4516 27226
rect 4220 27172 4276 27174
rect 4300 27172 4356 27174
rect 4380 27172 4436 27174
rect 4460 27172 4516 27174
rect 4220 26138 4276 26140
rect 4300 26138 4356 26140
rect 4380 26138 4436 26140
rect 4460 26138 4516 26140
rect 4220 26086 4246 26138
rect 4246 26086 4276 26138
rect 4300 26086 4310 26138
rect 4310 26086 4356 26138
rect 4380 26086 4426 26138
rect 4426 26086 4436 26138
rect 4460 26086 4490 26138
rect 4490 26086 4516 26138
rect 4220 26084 4276 26086
rect 4300 26084 4356 26086
rect 4380 26084 4436 26086
rect 4460 26084 4516 26086
rect 3974 25064 4030 25120
rect 4220 25050 4276 25052
rect 4300 25050 4356 25052
rect 4380 25050 4436 25052
rect 4460 25050 4516 25052
rect 4220 24998 4246 25050
rect 4246 24998 4276 25050
rect 4300 24998 4310 25050
rect 4310 24998 4356 25050
rect 4380 24998 4426 25050
rect 4426 24998 4436 25050
rect 4460 24998 4490 25050
rect 4490 24998 4516 25050
rect 4220 24996 4276 24998
rect 4300 24996 4356 24998
rect 4380 24996 4436 24998
rect 4460 24996 4516 24998
rect 4220 23962 4276 23964
rect 4300 23962 4356 23964
rect 4380 23962 4436 23964
rect 4460 23962 4516 23964
rect 4220 23910 4246 23962
rect 4246 23910 4276 23962
rect 4300 23910 4310 23962
rect 4310 23910 4356 23962
rect 4380 23910 4426 23962
rect 4426 23910 4436 23962
rect 4460 23910 4490 23962
rect 4490 23910 4516 23962
rect 4220 23908 4276 23910
rect 4300 23908 4356 23910
rect 4380 23908 4436 23910
rect 4460 23908 4516 23910
rect 4220 22874 4276 22876
rect 4300 22874 4356 22876
rect 4380 22874 4436 22876
rect 4460 22874 4516 22876
rect 4220 22822 4246 22874
rect 4246 22822 4276 22874
rect 4300 22822 4310 22874
rect 4310 22822 4356 22874
rect 4380 22822 4426 22874
rect 4426 22822 4436 22874
rect 4460 22822 4490 22874
rect 4490 22822 4516 22874
rect 4220 22820 4276 22822
rect 4300 22820 4356 22822
rect 4380 22820 4436 22822
rect 4460 22820 4516 22822
rect 4220 21786 4276 21788
rect 4300 21786 4356 21788
rect 4380 21786 4436 21788
rect 4460 21786 4516 21788
rect 4220 21734 4246 21786
rect 4246 21734 4276 21786
rect 4300 21734 4310 21786
rect 4310 21734 4356 21786
rect 4380 21734 4426 21786
rect 4426 21734 4436 21786
rect 4460 21734 4490 21786
rect 4490 21734 4516 21786
rect 4220 21732 4276 21734
rect 4300 21732 4356 21734
rect 4380 21732 4436 21734
rect 4460 21732 4516 21734
rect 4220 20698 4276 20700
rect 4300 20698 4356 20700
rect 4380 20698 4436 20700
rect 4460 20698 4516 20700
rect 4220 20646 4246 20698
rect 4246 20646 4276 20698
rect 4300 20646 4310 20698
rect 4310 20646 4356 20698
rect 4380 20646 4426 20698
rect 4426 20646 4436 20698
rect 4460 20646 4490 20698
rect 4490 20646 4516 20698
rect 4220 20644 4276 20646
rect 4300 20644 4356 20646
rect 4380 20644 4436 20646
rect 4460 20644 4516 20646
rect 4220 19610 4276 19612
rect 4300 19610 4356 19612
rect 4380 19610 4436 19612
rect 4460 19610 4516 19612
rect 4220 19558 4246 19610
rect 4246 19558 4276 19610
rect 4300 19558 4310 19610
rect 4310 19558 4356 19610
rect 4380 19558 4426 19610
rect 4426 19558 4436 19610
rect 4460 19558 4490 19610
rect 4490 19558 4516 19610
rect 4220 19556 4276 19558
rect 4300 19556 4356 19558
rect 4380 19556 4436 19558
rect 4460 19556 4516 19558
rect 3974 19352 4030 19408
rect 4066 19080 4122 19136
rect 4220 18522 4276 18524
rect 4300 18522 4356 18524
rect 4380 18522 4436 18524
rect 4460 18522 4516 18524
rect 4220 18470 4246 18522
rect 4246 18470 4276 18522
rect 4300 18470 4310 18522
rect 4310 18470 4356 18522
rect 4380 18470 4426 18522
rect 4426 18470 4436 18522
rect 4460 18470 4490 18522
rect 4490 18470 4516 18522
rect 4220 18468 4276 18470
rect 4300 18468 4356 18470
rect 4380 18468 4436 18470
rect 4460 18468 4516 18470
rect 4220 17434 4276 17436
rect 4300 17434 4356 17436
rect 4380 17434 4436 17436
rect 4460 17434 4516 17436
rect 4220 17382 4246 17434
rect 4246 17382 4276 17434
rect 4300 17382 4310 17434
rect 4310 17382 4356 17434
rect 4380 17382 4426 17434
rect 4426 17382 4436 17434
rect 4460 17382 4490 17434
rect 4490 17382 4516 17434
rect 4220 17380 4276 17382
rect 4300 17380 4356 17382
rect 4380 17380 4436 17382
rect 4460 17380 4516 17382
rect 4220 16346 4276 16348
rect 4300 16346 4356 16348
rect 4380 16346 4436 16348
rect 4460 16346 4516 16348
rect 4220 16294 4246 16346
rect 4246 16294 4276 16346
rect 4300 16294 4310 16346
rect 4310 16294 4356 16346
rect 4380 16294 4426 16346
rect 4426 16294 4436 16346
rect 4460 16294 4490 16346
rect 4490 16294 4516 16346
rect 4220 16292 4276 16294
rect 4300 16292 4356 16294
rect 4380 16292 4436 16294
rect 4460 16292 4516 16294
rect 4066 15816 4122 15872
rect 4220 15258 4276 15260
rect 4300 15258 4356 15260
rect 4380 15258 4436 15260
rect 4460 15258 4516 15260
rect 4220 15206 4246 15258
rect 4246 15206 4276 15258
rect 4300 15206 4310 15258
rect 4310 15206 4356 15258
rect 4380 15206 4426 15258
rect 4426 15206 4436 15258
rect 4460 15206 4490 15258
rect 4490 15206 4516 15258
rect 4220 15204 4276 15206
rect 4300 15204 4356 15206
rect 4380 15204 4436 15206
rect 4460 15204 4516 15206
rect 3146 14320 3202 14376
rect 4220 14170 4276 14172
rect 4300 14170 4356 14172
rect 4380 14170 4436 14172
rect 4460 14170 4516 14172
rect 4220 14118 4246 14170
rect 4246 14118 4276 14170
rect 4300 14118 4310 14170
rect 4310 14118 4356 14170
rect 4380 14118 4426 14170
rect 4426 14118 4436 14170
rect 4460 14118 4490 14170
rect 4490 14118 4516 14170
rect 4220 14116 4276 14118
rect 4300 14116 4356 14118
rect 4380 14116 4436 14118
rect 4460 14116 4516 14118
rect 2870 13368 2926 13424
rect 2686 12824 2742 12880
rect 4220 13082 4276 13084
rect 4300 13082 4356 13084
rect 4380 13082 4436 13084
rect 4460 13082 4516 13084
rect 4220 13030 4246 13082
rect 4246 13030 4276 13082
rect 4300 13030 4310 13082
rect 4310 13030 4356 13082
rect 4380 13030 4426 13082
rect 4426 13030 4436 13082
rect 4460 13030 4490 13082
rect 4490 13030 4516 13082
rect 4220 13028 4276 13030
rect 4300 13028 4356 13030
rect 4380 13028 4436 13030
rect 4460 13028 4516 13030
rect 4220 11994 4276 11996
rect 4300 11994 4356 11996
rect 4380 11994 4436 11996
rect 4460 11994 4516 11996
rect 4220 11942 4246 11994
rect 4246 11942 4276 11994
rect 4300 11942 4310 11994
rect 4310 11942 4356 11994
rect 4380 11942 4426 11994
rect 4426 11942 4436 11994
rect 4460 11942 4490 11994
rect 4490 11942 4516 11994
rect 4220 11940 4276 11942
rect 4300 11940 4356 11942
rect 4380 11940 4436 11942
rect 4460 11940 4516 11942
rect 2778 9832 2834 9888
rect 2778 6840 2834 6896
rect 4220 10906 4276 10908
rect 4300 10906 4356 10908
rect 4380 10906 4436 10908
rect 4460 10906 4516 10908
rect 4220 10854 4246 10906
rect 4246 10854 4276 10906
rect 4300 10854 4310 10906
rect 4310 10854 4356 10906
rect 4380 10854 4426 10906
rect 4426 10854 4436 10906
rect 4460 10854 4490 10906
rect 4490 10854 4516 10906
rect 4220 10852 4276 10854
rect 4300 10852 4356 10854
rect 4380 10852 4436 10854
rect 4460 10852 4516 10854
rect 3606 10532 3662 10568
rect 3606 10512 3608 10532
rect 3608 10512 3660 10532
rect 3660 10512 3662 10532
rect 4220 9818 4276 9820
rect 4300 9818 4356 9820
rect 4380 9818 4436 9820
rect 4460 9818 4516 9820
rect 4220 9766 4246 9818
rect 4246 9766 4276 9818
rect 4300 9766 4310 9818
rect 4310 9766 4356 9818
rect 4380 9766 4426 9818
rect 4426 9766 4436 9818
rect 4460 9766 4490 9818
rect 4490 9766 4516 9818
rect 4220 9764 4276 9766
rect 4300 9764 4356 9766
rect 4380 9764 4436 9766
rect 4460 9764 4516 9766
rect 4220 8730 4276 8732
rect 4300 8730 4356 8732
rect 4380 8730 4436 8732
rect 4460 8730 4516 8732
rect 4220 8678 4246 8730
rect 4246 8678 4276 8730
rect 4300 8678 4310 8730
rect 4310 8678 4356 8730
rect 4380 8678 4426 8730
rect 4426 8678 4436 8730
rect 4460 8678 4490 8730
rect 4490 8678 4516 8730
rect 4220 8676 4276 8678
rect 4300 8676 4356 8678
rect 4380 8676 4436 8678
rect 4460 8676 4516 8678
rect 4220 7642 4276 7644
rect 4300 7642 4356 7644
rect 4380 7642 4436 7644
rect 4460 7642 4516 7644
rect 4220 7590 4246 7642
rect 4246 7590 4276 7642
rect 4300 7590 4310 7642
rect 4310 7590 4356 7642
rect 4380 7590 4426 7642
rect 4426 7590 4436 7642
rect 4460 7590 4490 7642
rect 4490 7590 4516 7642
rect 4220 7588 4276 7590
rect 4300 7588 4356 7590
rect 4380 7588 4436 7590
rect 4460 7588 4516 7590
rect 4220 6554 4276 6556
rect 4300 6554 4356 6556
rect 4380 6554 4436 6556
rect 4460 6554 4516 6556
rect 4220 6502 4246 6554
rect 4246 6502 4276 6554
rect 4300 6502 4310 6554
rect 4310 6502 4356 6554
rect 4380 6502 4426 6554
rect 4426 6502 4436 6554
rect 4460 6502 4490 6554
rect 4490 6502 4516 6554
rect 4220 6500 4276 6502
rect 4300 6500 4356 6502
rect 4380 6500 4436 6502
rect 4460 6500 4516 6502
rect 4220 5466 4276 5468
rect 4300 5466 4356 5468
rect 4380 5466 4436 5468
rect 4460 5466 4516 5468
rect 4220 5414 4246 5466
rect 4246 5414 4276 5466
rect 4300 5414 4310 5466
rect 4310 5414 4356 5466
rect 4380 5414 4426 5466
rect 4426 5414 4436 5466
rect 4460 5414 4490 5466
rect 4490 5414 4516 5466
rect 4220 5412 4276 5414
rect 4300 5412 4356 5414
rect 4380 5412 4436 5414
rect 4460 5412 4516 5414
rect 4220 4378 4276 4380
rect 4300 4378 4356 4380
rect 4380 4378 4436 4380
rect 4460 4378 4516 4380
rect 4220 4326 4246 4378
rect 4246 4326 4276 4378
rect 4300 4326 4310 4378
rect 4310 4326 4356 4378
rect 4380 4326 4426 4378
rect 4426 4326 4436 4378
rect 4460 4326 4490 4378
rect 4490 4326 4516 4378
rect 4220 4324 4276 4326
rect 4300 4324 4356 4326
rect 4380 4324 4436 4326
rect 4460 4324 4516 4326
rect 5906 15136 5962 15192
rect 7470 33396 7472 33416
rect 7472 33396 7524 33416
rect 7524 33396 7526 33416
rect 7470 33360 7526 33396
rect 6826 15000 6882 15056
rect 6826 9036 6882 9072
rect 6826 9016 6828 9036
rect 6828 9016 6880 9036
rect 6880 9016 6882 9036
rect 8022 33360 8078 33416
rect 9126 33396 9128 33416
rect 9128 33396 9180 33416
rect 9180 33396 9182 33416
rect 9126 33360 9182 33396
rect 10598 30096 10654 30152
rect 7930 19352 7986 19408
rect 4220 3290 4276 3292
rect 4300 3290 4356 3292
rect 4380 3290 4436 3292
rect 4460 3290 4516 3292
rect 4220 3238 4246 3290
rect 4246 3238 4276 3290
rect 4300 3238 4310 3290
rect 4310 3238 4356 3290
rect 4380 3238 4426 3290
rect 4426 3238 4436 3290
rect 4460 3238 4490 3290
rect 4490 3238 4516 3290
rect 4220 3236 4276 3238
rect 4300 3236 4356 3238
rect 4380 3236 4436 3238
rect 4460 3236 4516 3238
rect 4220 2202 4276 2204
rect 4300 2202 4356 2204
rect 4380 2202 4436 2204
rect 4460 2202 4516 2204
rect 4220 2150 4246 2202
rect 4246 2150 4276 2202
rect 4300 2150 4310 2202
rect 4310 2150 4356 2202
rect 4380 2150 4426 2202
rect 4426 2150 4436 2202
rect 4460 2150 4490 2202
rect 4490 2150 4516 2202
rect 4220 2148 4276 2150
rect 4300 2148 4356 2150
rect 4380 2148 4436 2150
rect 4460 2148 4516 2150
rect 8758 12824 8814 12880
rect 9494 21800 9550 21856
rect 12438 22072 12494 22128
rect 9862 15136 9918 15192
rect 8574 8064 8630 8120
rect 10690 12688 10746 12744
rect 9862 10376 9918 10432
rect 11058 10784 11114 10840
rect 10046 3052 10102 3088
rect 10046 3032 10048 3052
rect 10048 3032 10100 3052
rect 10100 3032 10102 3052
rect 11334 12824 11390 12880
rect 12438 19216 12494 19272
rect 12898 22072 12954 22128
rect 14370 21528 14426 21584
rect 11702 9968 11758 10024
rect 11610 8064 11666 8120
rect 13174 14456 13230 14512
rect 12714 11056 12770 11112
rect 11150 7656 11206 7712
rect 11426 7384 11482 7440
rect 10966 5108 10968 5128
rect 10968 5108 11020 5128
rect 11020 5108 11022 5128
rect 10966 5072 11022 5108
rect 12990 7384 13046 7440
rect 14462 15156 14518 15192
rect 14462 15136 14464 15156
rect 14464 15136 14516 15156
rect 14516 15136 14518 15156
rect 14738 11600 14794 11656
rect 15014 10376 15070 10432
rect 15290 15020 15346 15056
rect 15290 15000 15292 15020
rect 15292 15000 15344 15020
rect 15344 15000 15346 15020
rect 13726 5072 13782 5128
rect 15566 9152 15622 9208
rect 15842 10804 15898 10840
rect 15842 10784 15844 10804
rect 15844 10784 15896 10804
rect 15896 10784 15898 10804
rect 19580 37562 19636 37564
rect 19660 37562 19716 37564
rect 19740 37562 19796 37564
rect 19820 37562 19876 37564
rect 19580 37510 19606 37562
rect 19606 37510 19636 37562
rect 19660 37510 19670 37562
rect 19670 37510 19716 37562
rect 19740 37510 19786 37562
rect 19786 37510 19796 37562
rect 19820 37510 19850 37562
rect 19850 37510 19876 37562
rect 19580 37508 19636 37510
rect 19660 37508 19716 37510
rect 19740 37508 19796 37510
rect 19820 37508 19876 37510
rect 19580 36474 19636 36476
rect 19660 36474 19716 36476
rect 19740 36474 19796 36476
rect 19820 36474 19876 36476
rect 19580 36422 19606 36474
rect 19606 36422 19636 36474
rect 19660 36422 19670 36474
rect 19670 36422 19716 36474
rect 19740 36422 19786 36474
rect 19786 36422 19796 36474
rect 19820 36422 19850 36474
rect 19850 36422 19876 36474
rect 19580 36420 19636 36422
rect 19660 36420 19716 36422
rect 19740 36420 19796 36422
rect 19820 36420 19876 36422
rect 17038 30132 17040 30152
rect 17040 30132 17092 30152
rect 17092 30132 17094 30152
rect 17038 30096 17094 30132
rect 17774 30096 17830 30152
rect 16762 12688 16818 12744
rect 16210 10124 16266 10160
rect 16210 10104 16212 10124
rect 16212 10104 16264 10124
rect 16264 10104 16266 10124
rect 16946 15136 17002 15192
rect 19580 35386 19636 35388
rect 19660 35386 19716 35388
rect 19740 35386 19796 35388
rect 19820 35386 19876 35388
rect 19580 35334 19606 35386
rect 19606 35334 19636 35386
rect 19660 35334 19670 35386
rect 19670 35334 19716 35386
rect 19740 35334 19786 35386
rect 19786 35334 19796 35386
rect 19820 35334 19850 35386
rect 19850 35334 19876 35386
rect 19580 35332 19636 35334
rect 19660 35332 19716 35334
rect 19740 35332 19796 35334
rect 19820 35332 19876 35334
rect 18418 21936 18474 21992
rect 19580 34298 19636 34300
rect 19660 34298 19716 34300
rect 19740 34298 19796 34300
rect 19820 34298 19876 34300
rect 19580 34246 19606 34298
rect 19606 34246 19636 34298
rect 19660 34246 19670 34298
rect 19670 34246 19716 34298
rect 19740 34246 19786 34298
rect 19786 34246 19796 34298
rect 19820 34246 19850 34298
rect 19850 34246 19876 34298
rect 19580 34244 19636 34246
rect 19660 34244 19716 34246
rect 19740 34244 19796 34246
rect 19820 34244 19876 34246
rect 19580 33210 19636 33212
rect 19660 33210 19716 33212
rect 19740 33210 19796 33212
rect 19820 33210 19876 33212
rect 19580 33158 19606 33210
rect 19606 33158 19636 33210
rect 19660 33158 19670 33210
rect 19670 33158 19716 33210
rect 19740 33158 19786 33210
rect 19786 33158 19796 33210
rect 19820 33158 19850 33210
rect 19850 33158 19876 33210
rect 19580 33156 19636 33158
rect 19660 33156 19716 33158
rect 19740 33156 19796 33158
rect 19820 33156 19876 33158
rect 19580 32122 19636 32124
rect 19660 32122 19716 32124
rect 19740 32122 19796 32124
rect 19820 32122 19876 32124
rect 19580 32070 19606 32122
rect 19606 32070 19636 32122
rect 19660 32070 19670 32122
rect 19670 32070 19716 32122
rect 19740 32070 19786 32122
rect 19786 32070 19796 32122
rect 19820 32070 19850 32122
rect 19850 32070 19876 32122
rect 19580 32068 19636 32070
rect 19660 32068 19716 32070
rect 19740 32068 19796 32070
rect 19820 32068 19876 32070
rect 19580 31034 19636 31036
rect 19660 31034 19716 31036
rect 19740 31034 19796 31036
rect 19820 31034 19876 31036
rect 19580 30982 19606 31034
rect 19606 30982 19636 31034
rect 19660 30982 19670 31034
rect 19670 30982 19716 31034
rect 19740 30982 19786 31034
rect 19786 30982 19796 31034
rect 19820 30982 19850 31034
rect 19850 30982 19876 31034
rect 19580 30980 19636 30982
rect 19660 30980 19716 30982
rect 19740 30980 19796 30982
rect 19820 30980 19876 30982
rect 19580 29946 19636 29948
rect 19660 29946 19716 29948
rect 19740 29946 19796 29948
rect 19820 29946 19876 29948
rect 19580 29894 19606 29946
rect 19606 29894 19636 29946
rect 19660 29894 19670 29946
rect 19670 29894 19716 29946
rect 19740 29894 19786 29946
rect 19786 29894 19796 29946
rect 19820 29894 19850 29946
rect 19850 29894 19876 29946
rect 19580 29892 19636 29894
rect 19660 29892 19716 29894
rect 19740 29892 19796 29894
rect 19820 29892 19876 29894
rect 19706 29572 19762 29608
rect 19706 29552 19708 29572
rect 19708 29552 19760 29572
rect 19760 29552 19762 29572
rect 19580 28858 19636 28860
rect 19660 28858 19716 28860
rect 19740 28858 19796 28860
rect 19820 28858 19876 28860
rect 19580 28806 19606 28858
rect 19606 28806 19636 28858
rect 19660 28806 19670 28858
rect 19670 28806 19716 28858
rect 19740 28806 19786 28858
rect 19786 28806 19796 28858
rect 19820 28806 19850 28858
rect 19850 28806 19876 28858
rect 19580 28804 19636 28806
rect 19660 28804 19716 28806
rect 19740 28804 19796 28806
rect 19820 28804 19876 28806
rect 19580 27770 19636 27772
rect 19660 27770 19716 27772
rect 19740 27770 19796 27772
rect 19820 27770 19876 27772
rect 19580 27718 19606 27770
rect 19606 27718 19636 27770
rect 19660 27718 19670 27770
rect 19670 27718 19716 27770
rect 19740 27718 19786 27770
rect 19786 27718 19796 27770
rect 19820 27718 19850 27770
rect 19850 27718 19876 27770
rect 19580 27716 19636 27718
rect 19660 27716 19716 27718
rect 19740 27716 19796 27718
rect 19820 27716 19876 27718
rect 19580 26682 19636 26684
rect 19660 26682 19716 26684
rect 19740 26682 19796 26684
rect 19820 26682 19876 26684
rect 19580 26630 19606 26682
rect 19606 26630 19636 26682
rect 19660 26630 19670 26682
rect 19670 26630 19716 26682
rect 19740 26630 19786 26682
rect 19786 26630 19796 26682
rect 19820 26630 19850 26682
rect 19850 26630 19876 26682
rect 19580 26628 19636 26630
rect 19660 26628 19716 26630
rect 19740 26628 19796 26630
rect 19820 26628 19876 26630
rect 19706 26460 19708 26480
rect 19708 26460 19760 26480
rect 19760 26460 19762 26480
rect 19706 26424 19762 26460
rect 20074 26424 20130 26480
rect 19580 25594 19636 25596
rect 19660 25594 19716 25596
rect 19740 25594 19796 25596
rect 19820 25594 19876 25596
rect 19580 25542 19606 25594
rect 19606 25542 19636 25594
rect 19660 25542 19670 25594
rect 19670 25542 19716 25594
rect 19740 25542 19786 25594
rect 19786 25542 19796 25594
rect 19820 25542 19850 25594
rect 19850 25542 19876 25594
rect 19580 25540 19636 25542
rect 19660 25540 19716 25542
rect 19740 25540 19796 25542
rect 19820 25540 19876 25542
rect 19580 24506 19636 24508
rect 19660 24506 19716 24508
rect 19740 24506 19796 24508
rect 19820 24506 19876 24508
rect 19580 24454 19606 24506
rect 19606 24454 19636 24506
rect 19660 24454 19670 24506
rect 19670 24454 19716 24506
rect 19740 24454 19786 24506
rect 19786 24454 19796 24506
rect 19820 24454 19850 24506
rect 19850 24454 19876 24506
rect 19580 24452 19636 24454
rect 19660 24452 19716 24454
rect 19740 24452 19796 24454
rect 19820 24452 19876 24454
rect 19580 23418 19636 23420
rect 19660 23418 19716 23420
rect 19740 23418 19796 23420
rect 19820 23418 19876 23420
rect 19580 23366 19606 23418
rect 19606 23366 19636 23418
rect 19660 23366 19670 23418
rect 19670 23366 19716 23418
rect 19740 23366 19786 23418
rect 19786 23366 19796 23418
rect 19820 23366 19850 23418
rect 19850 23366 19876 23418
rect 19580 23364 19636 23366
rect 19660 23364 19716 23366
rect 19740 23364 19796 23366
rect 19820 23364 19876 23366
rect 18050 19252 18052 19272
rect 18052 19252 18104 19272
rect 18104 19252 18106 19272
rect 18050 19216 18106 19252
rect 17498 14340 17554 14376
rect 17498 14320 17500 14340
rect 17500 14320 17552 14340
rect 17552 14320 17554 14340
rect 16762 9016 16818 9072
rect 16210 8372 16212 8392
rect 16212 8372 16264 8392
rect 16264 8372 16266 8392
rect 16210 8336 16266 8372
rect 17314 8372 17316 8392
rect 17316 8372 17368 8392
rect 17368 8372 17370 8392
rect 17314 8336 17370 8372
rect 16854 8200 16910 8256
rect 17498 7656 17554 7712
rect 16854 3052 16910 3088
rect 16854 3032 16856 3052
rect 16856 3032 16908 3052
rect 16908 3032 16910 3052
rect 18418 12144 18474 12200
rect 19580 22330 19636 22332
rect 19660 22330 19716 22332
rect 19740 22330 19796 22332
rect 19820 22330 19876 22332
rect 19580 22278 19606 22330
rect 19606 22278 19636 22330
rect 19660 22278 19670 22330
rect 19670 22278 19716 22330
rect 19740 22278 19786 22330
rect 19786 22278 19796 22330
rect 19820 22278 19850 22330
rect 19850 22278 19876 22330
rect 19580 22276 19636 22278
rect 19660 22276 19716 22278
rect 19740 22276 19796 22278
rect 19820 22276 19876 22278
rect 19430 21528 19486 21584
rect 20074 21800 20130 21856
rect 19580 21242 19636 21244
rect 19660 21242 19716 21244
rect 19740 21242 19796 21244
rect 19820 21242 19876 21244
rect 19580 21190 19606 21242
rect 19606 21190 19636 21242
rect 19660 21190 19670 21242
rect 19670 21190 19716 21242
rect 19740 21190 19786 21242
rect 19786 21190 19796 21242
rect 19820 21190 19850 21242
rect 19850 21190 19876 21242
rect 19580 21188 19636 21190
rect 19660 21188 19716 21190
rect 19740 21188 19796 21190
rect 19820 21188 19876 21190
rect 19580 20154 19636 20156
rect 19660 20154 19716 20156
rect 19740 20154 19796 20156
rect 19820 20154 19876 20156
rect 19580 20102 19606 20154
rect 19606 20102 19636 20154
rect 19660 20102 19670 20154
rect 19670 20102 19716 20154
rect 19740 20102 19786 20154
rect 19786 20102 19796 20154
rect 19820 20102 19850 20154
rect 19850 20102 19876 20154
rect 19580 20100 19636 20102
rect 19660 20100 19716 20102
rect 19740 20100 19796 20102
rect 19820 20100 19876 20102
rect 19580 19066 19636 19068
rect 19660 19066 19716 19068
rect 19740 19066 19796 19068
rect 19820 19066 19876 19068
rect 19580 19014 19606 19066
rect 19606 19014 19636 19066
rect 19660 19014 19670 19066
rect 19670 19014 19716 19066
rect 19740 19014 19786 19066
rect 19786 19014 19796 19066
rect 19820 19014 19850 19066
rect 19850 19014 19876 19066
rect 19580 19012 19636 19014
rect 19660 19012 19716 19014
rect 19740 19012 19796 19014
rect 19820 19012 19876 19014
rect 20718 26832 20774 26888
rect 19580 17978 19636 17980
rect 19660 17978 19716 17980
rect 19740 17978 19796 17980
rect 19820 17978 19876 17980
rect 19580 17926 19606 17978
rect 19606 17926 19636 17978
rect 19660 17926 19670 17978
rect 19670 17926 19716 17978
rect 19740 17926 19786 17978
rect 19786 17926 19796 17978
rect 19820 17926 19850 17978
rect 19850 17926 19876 17978
rect 19580 17924 19636 17926
rect 19660 17924 19716 17926
rect 19740 17924 19796 17926
rect 19820 17924 19876 17926
rect 19580 16890 19636 16892
rect 19660 16890 19716 16892
rect 19740 16890 19796 16892
rect 19820 16890 19876 16892
rect 19580 16838 19606 16890
rect 19606 16838 19636 16890
rect 19660 16838 19670 16890
rect 19670 16838 19716 16890
rect 19740 16838 19786 16890
rect 19786 16838 19796 16890
rect 19820 16838 19850 16890
rect 19850 16838 19876 16890
rect 19580 16836 19636 16838
rect 19660 16836 19716 16838
rect 19740 16836 19796 16838
rect 19820 16836 19876 16838
rect 19580 15802 19636 15804
rect 19660 15802 19716 15804
rect 19740 15802 19796 15804
rect 19820 15802 19876 15804
rect 19580 15750 19606 15802
rect 19606 15750 19636 15802
rect 19660 15750 19670 15802
rect 19670 15750 19716 15802
rect 19740 15750 19786 15802
rect 19786 15750 19796 15802
rect 19820 15750 19850 15802
rect 19850 15750 19876 15802
rect 19580 15748 19636 15750
rect 19660 15748 19716 15750
rect 19740 15748 19796 15750
rect 19820 15748 19876 15750
rect 18786 11636 18788 11656
rect 18788 11636 18840 11656
rect 18840 11636 18842 11656
rect 18786 11600 18842 11636
rect 18970 9152 19026 9208
rect 18970 8200 19026 8256
rect 19580 14714 19636 14716
rect 19660 14714 19716 14716
rect 19740 14714 19796 14716
rect 19820 14714 19876 14716
rect 19580 14662 19606 14714
rect 19606 14662 19636 14714
rect 19660 14662 19670 14714
rect 19670 14662 19716 14714
rect 19740 14662 19786 14714
rect 19786 14662 19796 14714
rect 19820 14662 19850 14714
rect 19850 14662 19876 14714
rect 19580 14660 19636 14662
rect 19660 14660 19716 14662
rect 19740 14660 19796 14662
rect 19820 14660 19876 14662
rect 19890 14476 19946 14512
rect 19890 14456 19892 14476
rect 19892 14456 19944 14476
rect 19944 14456 19946 14476
rect 19580 13626 19636 13628
rect 19660 13626 19716 13628
rect 19740 13626 19796 13628
rect 19820 13626 19876 13628
rect 19580 13574 19606 13626
rect 19606 13574 19636 13626
rect 19660 13574 19670 13626
rect 19670 13574 19716 13626
rect 19740 13574 19786 13626
rect 19786 13574 19796 13626
rect 19820 13574 19850 13626
rect 19850 13574 19876 13626
rect 19580 13572 19636 13574
rect 19660 13572 19716 13574
rect 19740 13572 19796 13574
rect 19820 13572 19876 13574
rect 20350 18692 20406 18728
rect 20350 18672 20352 18692
rect 20352 18672 20404 18692
rect 20404 18672 20406 18692
rect 19580 12538 19636 12540
rect 19660 12538 19716 12540
rect 19740 12538 19796 12540
rect 19820 12538 19876 12540
rect 19580 12486 19606 12538
rect 19606 12486 19636 12538
rect 19660 12486 19670 12538
rect 19670 12486 19716 12538
rect 19740 12486 19786 12538
rect 19786 12486 19796 12538
rect 19820 12486 19850 12538
rect 19850 12486 19876 12538
rect 19580 12484 19636 12486
rect 19660 12484 19716 12486
rect 19740 12484 19796 12486
rect 19820 12484 19876 12486
rect 19580 11450 19636 11452
rect 19660 11450 19716 11452
rect 19740 11450 19796 11452
rect 19820 11450 19876 11452
rect 19580 11398 19606 11450
rect 19606 11398 19636 11450
rect 19660 11398 19670 11450
rect 19670 11398 19716 11450
rect 19740 11398 19786 11450
rect 19786 11398 19796 11450
rect 19820 11398 19850 11450
rect 19850 11398 19876 11450
rect 19580 11396 19636 11398
rect 19660 11396 19716 11398
rect 19740 11396 19796 11398
rect 19820 11396 19876 11398
rect 19580 10362 19636 10364
rect 19660 10362 19716 10364
rect 19740 10362 19796 10364
rect 19820 10362 19876 10364
rect 19580 10310 19606 10362
rect 19606 10310 19636 10362
rect 19660 10310 19670 10362
rect 19670 10310 19716 10362
rect 19740 10310 19786 10362
rect 19786 10310 19796 10362
rect 19820 10310 19850 10362
rect 19850 10310 19876 10362
rect 19580 10308 19636 10310
rect 19660 10308 19716 10310
rect 19740 10308 19796 10310
rect 19820 10308 19876 10310
rect 19580 9274 19636 9276
rect 19660 9274 19716 9276
rect 19740 9274 19796 9276
rect 19820 9274 19876 9276
rect 19580 9222 19606 9274
rect 19606 9222 19636 9274
rect 19660 9222 19670 9274
rect 19670 9222 19716 9274
rect 19740 9222 19786 9274
rect 19786 9222 19796 9274
rect 19820 9222 19850 9274
rect 19850 9222 19876 9274
rect 19580 9220 19636 9222
rect 19660 9220 19716 9222
rect 19740 9220 19796 9222
rect 19820 9220 19876 9222
rect 19430 9016 19486 9072
rect 19580 8186 19636 8188
rect 19660 8186 19716 8188
rect 19740 8186 19796 8188
rect 19820 8186 19876 8188
rect 19580 8134 19606 8186
rect 19606 8134 19636 8186
rect 19660 8134 19670 8186
rect 19670 8134 19716 8186
rect 19740 8134 19786 8186
rect 19786 8134 19796 8186
rect 19820 8134 19850 8186
rect 19850 8134 19876 8186
rect 19580 8132 19636 8134
rect 19660 8132 19716 8134
rect 19740 8132 19796 8134
rect 19820 8132 19876 8134
rect 19580 7098 19636 7100
rect 19660 7098 19716 7100
rect 19740 7098 19796 7100
rect 19820 7098 19876 7100
rect 19580 7046 19606 7098
rect 19606 7046 19636 7098
rect 19660 7046 19670 7098
rect 19670 7046 19716 7098
rect 19740 7046 19786 7098
rect 19786 7046 19796 7098
rect 19820 7046 19850 7098
rect 19850 7046 19876 7098
rect 19580 7044 19636 7046
rect 19660 7044 19716 7046
rect 19740 7044 19796 7046
rect 19820 7044 19876 7046
rect 19580 6010 19636 6012
rect 19660 6010 19716 6012
rect 19740 6010 19796 6012
rect 19820 6010 19876 6012
rect 19580 5958 19606 6010
rect 19606 5958 19636 6010
rect 19660 5958 19670 6010
rect 19670 5958 19716 6010
rect 19740 5958 19786 6010
rect 19786 5958 19796 6010
rect 19820 5958 19850 6010
rect 19850 5958 19876 6010
rect 19580 5956 19636 5958
rect 19660 5956 19716 5958
rect 19740 5956 19796 5958
rect 19820 5956 19876 5958
rect 19580 4922 19636 4924
rect 19660 4922 19716 4924
rect 19740 4922 19796 4924
rect 19820 4922 19876 4924
rect 19580 4870 19606 4922
rect 19606 4870 19636 4922
rect 19660 4870 19670 4922
rect 19670 4870 19716 4922
rect 19740 4870 19786 4922
rect 19786 4870 19796 4922
rect 19820 4870 19850 4922
rect 19850 4870 19876 4922
rect 19580 4868 19636 4870
rect 19660 4868 19716 4870
rect 19740 4868 19796 4870
rect 19820 4868 19876 4870
rect 20166 8472 20222 8528
rect 22098 26832 22154 26888
rect 20994 21800 21050 21856
rect 21270 19080 21326 19136
rect 21638 19624 21694 19680
rect 19580 3834 19636 3836
rect 19660 3834 19716 3836
rect 19740 3834 19796 3836
rect 19820 3834 19876 3836
rect 19580 3782 19606 3834
rect 19606 3782 19636 3834
rect 19660 3782 19670 3834
rect 19670 3782 19716 3834
rect 19740 3782 19786 3834
rect 19786 3782 19796 3834
rect 19820 3782 19850 3834
rect 19850 3782 19876 3834
rect 19580 3780 19636 3782
rect 19660 3780 19716 3782
rect 19740 3780 19796 3782
rect 19820 3780 19876 3782
rect 19580 2746 19636 2748
rect 19660 2746 19716 2748
rect 19740 2746 19796 2748
rect 19820 2746 19876 2748
rect 19580 2694 19606 2746
rect 19606 2694 19636 2746
rect 19660 2694 19670 2746
rect 19670 2694 19716 2746
rect 19740 2694 19786 2746
rect 19786 2694 19796 2746
rect 19820 2694 19850 2746
rect 19850 2694 19876 2746
rect 19580 2692 19636 2694
rect 19660 2692 19716 2694
rect 19740 2692 19796 2694
rect 19820 2692 19876 2694
rect 20902 8492 20958 8528
rect 20902 8472 20904 8492
rect 20904 8472 20956 8492
rect 20956 8472 20958 8492
rect 21454 15988 21456 16008
rect 21456 15988 21508 16008
rect 21508 15988 21510 16008
rect 21454 15952 21510 15988
rect 22098 19624 22154 19680
rect 22006 19080 22062 19136
rect 22834 26460 22836 26480
rect 22836 26460 22888 26480
rect 22888 26460 22890 26480
rect 22834 26424 22890 26460
rect 23294 29552 23350 29608
rect 22558 13368 22614 13424
rect 21914 11056 21970 11112
rect 22374 9016 22430 9072
rect 21730 7420 21732 7440
rect 21732 7420 21784 7440
rect 21784 7420 21786 7440
rect 21730 7384 21786 7420
rect 22098 5616 22154 5672
rect 22926 5616 22982 5672
rect 24490 30368 24546 30424
rect 24398 24928 24454 24984
rect 25226 19660 25228 19680
rect 25228 19660 25280 19680
rect 25280 19660 25282 19680
rect 25226 19624 25282 19660
rect 25042 19252 25044 19272
rect 25044 19252 25096 19272
rect 25096 19252 25098 19272
rect 25042 19216 25098 19252
rect 24766 16108 24822 16144
rect 24766 16088 24768 16108
rect 24768 16088 24820 16108
rect 24820 16088 24822 16108
rect 24582 7384 24638 7440
rect 26514 19372 26570 19408
rect 26514 19352 26516 19372
rect 26516 19352 26568 19372
rect 26568 19352 26570 19372
rect 26606 18672 26662 18728
rect 26974 18808 27030 18864
rect 27342 19352 27398 19408
rect 27250 19236 27306 19272
rect 27250 19216 27252 19236
rect 27252 19216 27304 19236
rect 27304 19216 27306 19236
rect 27894 19080 27950 19136
rect 27618 18808 27674 18864
rect 26514 17076 26516 17096
rect 26516 17076 26568 17096
rect 26568 17076 26570 17096
rect 26514 17040 26570 17076
rect 27802 16652 27858 16688
rect 27802 16632 27804 16652
rect 27804 16632 27856 16652
rect 27856 16632 27858 16652
rect 28262 17076 28264 17096
rect 28264 17076 28316 17096
rect 28316 17076 28318 17096
rect 28262 17040 28318 17076
rect 28998 16632 29054 16688
rect 34940 37018 34996 37020
rect 35020 37018 35076 37020
rect 35100 37018 35156 37020
rect 35180 37018 35236 37020
rect 34940 36966 34966 37018
rect 34966 36966 34996 37018
rect 35020 36966 35030 37018
rect 35030 36966 35076 37018
rect 35100 36966 35146 37018
rect 35146 36966 35156 37018
rect 35180 36966 35210 37018
rect 35210 36966 35236 37018
rect 34940 36964 34996 36966
rect 35020 36964 35076 36966
rect 35100 36964 35156 36966
rect 35180 36964 35236 36966
rect 38106 37576 38162 37632
rect 34940 35930 34996 35932
rect 35020 35930 35076 35932
rect 35100 35930 35156 35932
rect 35180 35930 35236 35932
rect 34940 35878 34966 35930
rect 34966 35878 34996 35930
rect 35020 35878 35030 35930
rect 35030 35878 35076 35930
rect 35100 35878 35146 35930
rect 35146 35878 35156 35930
rect 35180 35878 35210 35930
rect 35210 35878 35236 35930
rect 34940 35876 34996 35878
rect 35020 35876 35076 35878
rect 35100 35876 35156 35878
rect 35180 35876 35236 35878
rect 34940 34842 34996 34844
rect 35020 34842 35076 34844
rect 35100 34842 35156 34844
rect 35180 34842 35236 34844
rect 34940 34790 34966 34842
rect 34966 34790 34996 34842
rect 35020 34790 35030 34842
rect 35030 34790 35076 34842
rect 35100 34790 35146 34842
rect 35146 34790 35156 34842
rect 35180 34790 35210 34842
rect 35210 34790 35236 34842
rect 34940 34788 34996 34790
rect 35020 34788 35076 34790
rect 35100 34788 35156 34790
rect 35180 34788 35236 34790
rect 29826 22616 29882 22672
rect 30562 21528 30618 21584
rect 30930 21528 30986 21584
rect 34940 33754 34996 33756
rect 35020 33754 35076 33756
rect 35100 33754 35156 33756
rect 35180 33754 35236 33756
rect 34940 33702 34966 33754
rect 34966 33702 34996 33754
rect 35020 33702 35030 33754
rect 35030 33702 35076 33754
rect 35100 33702 35146 33754
rect 35146 33702 35156 33754
rect 35180 33702 35210 33754
rect 35210 33702 35236 33754
rect 34940 33700 34996 33702
rect 35020 33700 35076 33702
rect 35100 33700 35156 33702
rect 35180 33700 35236 33702
rect 34940 32666 34996 32668
rect 35020 32666 35076 32668
rect 35100 32666 35156 32668
rect 35180 32666 35236 32668
rect 34940 32614 34966 32666
rect 34966 32614 34996 32666
rect 35020 32614 35030 32666
rect 35030 32614 35076 32666
rect 35100 32614 35146 32666
rect 35146 32614 35156 32666
rect 35180 32614 35210 32666
rect 35210 32614 35236 32666
rect 34940 32612 34996 32614
rect 35020 32612 35076 32614
rect 35100 32612 35156 32614
rect 35180 32612 35236 32614
rect 34940 31578 34996 31580
rect 35020 31578 35076 31580
rect 35100 31578 35156 31580
rect 35180 31578 35236 31580
rect 34940 31526 34966 31578
rect 34966 31526 34996 31578
rect 35020 31526 35030 31578
rect 35030 31526 35076 31578
rect 35100 31526 35146 31578
rect 35146 31526 35156 31578
rect 35180 31526 35210 31578
rect 35210 31526 35236 31578
rect 34940 31524 34996 31526
rect 35020 31524 35076 31526
rect 35100 31524 35156 31526
rect 35180 31524 35236 31526
rect 35530 31592 35586 31648
rect 34940 30490 34996 30492
rect 35020 30490 35076 30492
rect 35100 30490 35156 30492
rect 35180 30490 35236 30492
rect 34940 30438 34966 30490
rect 34966 30438 34996 30490
rect 35020 30438 35030 30490
rect 35030 30438 35076 30490
rect 35100 30438 35146 30490
rect 35146 30438 35156 30490
rect 35180 30438 35210 30490
rect 35210 30438 35236 30490
rect 34940 30436 34996 30438
rect 35020 30436 35076 30438
rect 35100 30436 35156 30438
rect 35180 30436 35236 30438
rect 32586 28736 32642 28792
rect 29182 11636 29184 11656
rect 29184 11636 29236 11656
rect 29236 11636 29238 11656
rect 29182 11600 29238 11636
rect 29182 11212 29238 11248
rect 29182 11192 29184 11212
rect 29184 11192 29236 11212
rect 29236 11192 29238 11212
rect 28446 9560 28502 9616
rect 29274 10512 29330 10568
rect 29182 9036 29238 9072
rect 29182 9016 29184 9036
rect 29184 9016 29236 9036
rect 29236 9016 29238 9036
rect 28998 6704 29054 6760
rect 28630 5616 28686 5672
rect 30378 15952 30434 16008
rect 30194 11192 30250 11248
rect 29734 9696 29790 9752
rect 29734 8880 29790 8936
rect 30562 10376 30618 10432
rect 30562 8608 30618 8664
rect 31298 12008 31354 12064
rect 31942 11636 31944 11656
rect 31944 11636 31996 11656
rect 31996 11636 31998 11656
rect 31942 11600 31998 11636
rect 31850 11056 31906 11112
rect 31482 9696 31538 9752
rect 31758 9036 31814 9072
rect 31758 9016 31760 9036
rect 31760 9016 31812 9036
rect 31812 9016 31814 9036
rect 31942 6296 31998 6352
rect 34940 29402 34996 29404
rect 35020 29402 35076 29404
rect 35100 29402 35156 29404
rect 35180 29402 35236 29404
rect 34940 29350 34966 29402
rect 34966 29350 34996 29402
rect 35020 29350 35030 29402
rect 35030 29350 35076 29402
rect 35100 29350 35146 29402
rect 35146 29350 35156 29402
rect 35180 29350 35210 29402
rect 35210 29350 35236 29402
rect 34940 29348 34996 29350
rect 35020 29348 35076 29350
rect 35100 29348 35156 29350
rect 35180 29348 35236 29350
rect 34940 28314 34996 28316
rect 35020 28314 35076 28316
rect 35100 28314 35156 28316
rect 35180 28314 35236 28316
rect 34940 28262 34966 28314
rect 34966 28262 34996 28314
rect 35020 28262 35030 28314
rect 35030 28262 35076 28314
rect 35100 28262 35146 28314
rect 35146 28262 35156 28314
rect 35180 28262 35210 28314
rect 35210 28262 35236 28314
rect 34940 28260 34996 28262
rect 35020 28260 35076 28262
rect 35100 28260 35156 28262
rect 35180 28260 35236 28262
rect 34940 27226 34996 27228
rect 35020 27226 35076 27228
rect 35100 27226 35156 27228
rect 35180 27226 35236 27228
rect 34940 27174 34966 27226
rect 34966 27174 34996 27226
rect 35020 27174 35030 27226
rect 35030 27174 35076 27226
rect 35100 27174 35146 27226
rect 35146 27174 35156 27226
rect 35180 27174 35210 27226
rect 35210 27174 35236 27226
rect 34940 27172 34996 27174
rect 35020 27172 35076 27174
rect 35100 27172 35156 27174
rect 35180 27172 35236 27174
rect 33966 24676 34022 24712
rect 33966 24656 33968 24676
rect 33968 24656 34020 24676
rect 34020 24656 34022 24676
rect 34940 26138 34996 26140
rect 35020 26138 35076 26140
rect 35100 26138 35156 26140
rect 35180 26138 35236 26140
rect 34940 26086 34966 26138
rect 34966 26086 34996 26138
rect 35020 26086 35030 26138
rect 35030 26086 35076 26138
rect 35100 26086 35146 26138
rect 35146 26086 35156 26138
rect 35180 26086 35210 26138
rect 35210 26086 35236 26138
rect 34940 26084 34996 26086
rect 35020 26084 35076 26086
rect 35100 26084 35156 26086
rect 35180 26084 35236 26086
rect 35438 25336 35494 25392
rect 34940 25050 34996 25052
rect 35020 25050 35076 25052
rect 35100 25050 35156 25052
rect 35180 25050 35236 25052
rect 34940 24998 34966 25050
rect 34966 24998 34996 25050
rect 35020 24998 35030 25050
rect 35030 24998 35076 25050
rect 35100 24998 35146 25050
rect 35146 24998 35156 25050
rect 35180 24998 35210 25050
rect 35210 24998 35236 25050
rect 34940 24996 34996 24998
rect 35020 24996 35076 24998
rect 35100 24996 35156 24998
rect 35180 24996 35236 24998
rect 34940 23962 34996 23964
rect 35020 23962 35076 23964
rect 35100 23962 35156 23964
rect 35180 23962 35236 23964
rect 34940 23910 34966 23962
rect 34966 23910 34996 23962
rect 35020 23910 35030 23962
rect 35030 23910 35076 23962
rect 35100 23910 35146 23962
rect 35146 23910 35156 23962
rect 35180 23910 35210 23962
rect 35210 23910 35236 23962
rect 34940 23908 34996 23910
rect 35020 23908 35076 23910
rect 35100 23908 35156 23910
rect 35180 23908 35236 23910
rect 34940 22874 34996 22876
rect 35020 22874 35076 22876
rect 35100 22874 35156 22876
rect 35180 22874 35236 22876
rect 34940 22822 34966 22874
rect 34966 22822 34996 22874
rect 35020 22822 35030 22874
rect 35030 22822 35076 22874
rect 35100 22822 35146 22874
rect 35146 22822 35156 22874
rect 35180 22822 35210 22874
rect 35210 22822 35236 22874
rect 34940 22820 34996 22822
rect 35020 22820 35076 22822
rect 35100 22820 35156 22822
rect 35180 22820 35236 22822
rect 35346 22616 35402 22672
rect 34940 21786 34996 21788
rect 35020 21786 35076 21788
rect 35100 21786 35156 21788
rect 35180 21786 35236 21788
rect 34940 21734 34966 21786
rect 34966 21734 34996 21786
rect 35020 21734 35030 21786
rect 35030 21734 35076 21786
rect 35100 21734 35146 21786
rect 35146 21734 35156 21786
rect 35180 21734 35210 21786
rect 35210 21734 35236 21786
rect 34940 21732 34996 21734
rect 35020 21732 35076 21734
rect 35100 21732 35156 21734
rect 35180 21732 35236 21734
rect 32586 10548 32588 10568
rect 32588 10548 32640 10568
rect 32640 10548 32642 10568
rect 32586 10512 32642 10548
rect 33414 12008 33470 12064
rect 34940 20698 34996 20700
rect 35020 20698 35076 20700
rect 35100 20698 35156 20700
rect 35180 20698 35236 20700
rect 34940 20646 34966 20698
rect 34966 20646 34996 20698
rect 35020 20646 35030 20698
rect 35030 20646 35076 20698
rect 35100 20646 35146 20698
rect 35146 20646 35156 20698
rect 35180 20646 35210 20698
rect 35210 20646 35236 20698
rect 34940 20644 34996 20646
rect 35020 20644 35076 20646
rect 35100 20644 35156 20646
rect 35180 20644 35236 20646
rect 35530 22344 35586 22400
rect 34940 19610 34996 19612
rect 35020 19610 35076 19612
rect 35100 19610 35156 19612
rect 35180 19610 35236 19612
rect 34940 19558 34966 19610
rect 34966 19558 34996 19610
rect 35020 19558 35030 19610
rect 35030 19558 35076 19610
rect 35100 19558 35146 19610
rect 35146 19558 35156 19610
rect 35180 19558 35210 19610
rect 35210 19558 35236 19610
rect 34940 19556 34996 19558
rect 35020 19556 35076 19558
rect 35100 19556 35156 19558
rect 35180 19556 35236 19558
rect 34940 18522 34996 18524
rect 35020 18522 35076 18524
rect 35100 18522 35156 18524
rect 35180 18522 35236 18524
rect 34940 18470 34966 18522
rect 34966 18470 34996 18522
rect 35020 18470 35030 18522
rect 35030 18470 35076 18522
rect 35100 18470 35146 18522
rect 35146 18470 35156 18522
rect 35180 18470 35210 18522
rect 35210 18470 35236 18522
rect 34940 18468 34996 18470
rect 35020 18468 35076 18470
rect 35100 18468 35156 18470
rect 35180 18468 35236 18470
rect 30930 4684 30986 4720
rect 30930 4664 30932 4684
rect 30932 4664 30984 4684
rect 30984 4664 30986 4684
rect 34940 17434 34996 17436
rect 35020 17434 35076 17436
rect 35100 17434 35156 17436
rect 35180 17434 35236 17436
rect 34940 17382 34966 17434
rect 34966 17382 34996 17434
rect 35020 17382 35030 17434
rect 35030 17382 35076 17434
rect 35100 17382 35146 17434
rect 35146 17382 35156 17434
rect 35180 17382 35210 17434
rect 35210 17382 35236 17434
rect 34940 17380 34996 17382
rect 35020 17380 35076 17382
rect 35100 17380 35156 17382
rect 35180 17380 35236 17382
rect 34940 16346 34996 16348
rect 35020 16346 35076 16348
rect 35100 16346 35156 16348
rect 35180 16346 35236 16348
rect 34940 16294 34966 16346
rect 34966 16294 34996 16346
rect 35020 16294 35030 16346
rect 35030 16294 35076 16346
rect 35100 16294 35146 16346
rect 35146 16294 35156 16346
rect 35180 16294 35210 16346
rect 35210 16294 35236 16346
rect 34940 16292 34996 16294
rect 35020 16292 35076 16294
rect 35100 16292 35156 16294
rect 35180 16292 35236 16294
rect 34978 16108 35034 16144
rect 34978 16088 34980 16108
rect 34980 16088 35032 16108
rect 35032 16088 35034 16108
rect 34940 15258 34996 15260
rect 35020 15258 35076 15260
rect 35100 15258 35156 15260
rect 35180 15258 35236 15260
rect 34940 15206 34966 15258
rect 34966 15206 34996 15258
rect 35020 15206 35030 15258
rect 35030 15206 35076 15258
rect 35100 15206 35146 15258
rect 35146 15206 35156 15258
rect 35180 15206 35210 15258
rect 35210 15206 35236 15258
rect 34940 15204 34996 15206
rect 35020 15204 35076 15206
rect 35100 15204 35156 15206
rect 35180 15204 35236 15206
rect 34334 10376 34390 10432
rect 34150 8880 34206 8936
rect 33966 6740 33968 6760
rect 33968 6740 34020 6760
rect 34020 6740 34022 6760
rect 33966 6704 34022 6740
rect 37002 34584 37058 34640
rect 36266 29008 36322 29064
rect 36542 24656 36598 24712
rect 37922 28328 37978 28384
rect 34940 14170 34996 14172
rect 35020 14170 35076 14172
rect 35100 14170 35156 14172
rect 35180 14170 35236 14172
rect 34940 14118 34966 14170
rect 34966 14118 34996 14170
rect 35020 14118 35030 14170
rect 35030 14118 35076 14170
rect 35100 14118 35146 14170
rect 35146 14118 35156 14170
rect 35180 14118 35210 14170
rect 35210 14118 35236 14170
rect 34940 14116 34996 14118
rect 35020 14116 35076 14118
rect 35100 14116 35156 14118
rect 35180 14116 35236 14118
rect 35254 13368 35310 13424
rect 34940 13082 34996 13084
rect 35020 13082 35076 13084
rect 35100 13082 35156 13084
rect 35180 13082 35236 13084
rect 34940 13030 34966 13082
rect 34966 13030 34996 13082
rect 35020 13030 35030 13082
rect 35030 13030 35076 13082
rect 35100 13030 35146 13082
rect 35146 13030 35156 13082
rect 35180 13030 35210 13082
rect 35210 13030 35236 13082
rect 34940 13028 34996 13030
rect 35020 13028 35076 13030
rect 35100 13028 35156 13030
rect 35180 13028 35236 13030
rect 34940 11994 34996 11996
rect 35020 11994 35076 11996
rect 35100 11994 35156 11996
rect 35180 11994 35236 11996
rect 34940 11942 34966 11994
rect 34966 11942 34996 11994
rect 35020 11942 35030 11994
rect 35030 11942 35076 11994
rect 35100 11942 35146 11994
rect 35146 11942 35156 11994
rect 35180 11942 35210 11994
rect 35210 11942 35236 11994
rect 34940 11940 34996 11942
rect 35020 11940 35076 11942
rect 35100 11940 35156 11942
rect 35180 11940 35236 11942
rect 34940 10906 34996 10908
rect 35020 10906 35076 10908
rect 35100 10906 35156 10908
rect 35180 10906 35236 10908
rect 34940 10854 34966 10906
rect 34966 10854 34996 10906
rect 35020 10854 35030 10906
rect 35030 10854 35076 10906
rect 35100 10854 35146 10906
rect 35146 10854 35156 10906
rect 35180 10854 35210 10906
rect 35210 10854 35236 10906
rect 34940 10852 34996 10854
rect 35020 10852 35076 10854
rect 35100 10852 35156 10854
rect 35180 10852 35236 10854
rect 34610 8608 34666 8664
rect 34940 9818 34996 9820
rect 35020 9818 35076 9820
rect 35100 9818 35156 9820
rect 35180 9818 35236 9820
rect 34940 9766 34966 9818
rect 34966 9766 34996 9818
rect 35020 9766 35030 9818
rect 35030 9766 35076 9818
rect 35100 9766 35146 9818
rect 35146 9766 35156 9818
rect 35180 9766 35210 9818
rect 35210 9766 35236 9818
rect 34940 9764 34996 9766
rect 35020 9764 35076 9766
rect 35100 9764 35156 9766
rect 35180 9764 35236 9766
rect 34940 8730 34996 8732
rect 35020 8730 35076 8732
rect 35100 8730 35156 8732
rect 35180 8730 35236 8732
rect 34940 8678 34966 8730
rect 34966 8678 34996 8730
rect 35020 8678 35030 8730
rect 35030 8678 35076 8730
rect 35100 8678 35146 8730
rect 35146 8678 35156 8730
rect 35180 8678 35210 8730
rect 35210 8678 35236 8730
rect 34940 8676 34996 8678
rect 35020 8676 35076 8678
rect 35100 8676 35156 8678
rect 35180 8676 35236 8678
rect 34940 7642 34996 7644
rect 35020 7642 35076 7644
rect 35100 7642 35156 7644
rect 35180 7642 35236 7644
rect 34940 7590 34966 7642
rect 34966 7590 34996 7642
rect 35020 7590 35030 7642
rect 35030 7590 35076 7642
rect 35100 7590 35146 7642
rect 35146 7590 35156 7642
rect 35180 7590 35210 7642
rect 35210 7590 35236 7642
rect 34940 7588 34996 7590
rect 35020 7588 35076 7590
rect 35100 7588 35156 7590
rect 35180 7588 35236 7590
rect 34940 6554 34996 6556
rect 35020 6554 35076 6556
rect 35100 6554 35156 6556
rect 35180 6554 35236 6556
rect 34940 6502 34966 6554
rect 34966 6502 34996 6554
rect 35020 6502 35030 6554
rect 35030 6502 35076 6554
rect 35100 6502 35146 6554
rect 35146 6502 35156 6554
rect 35180 6502 35210 6554
rect 35210 6502 35236 6554
rect 34940 6500 34996 6502
rect 35020 6500 35076 6502
rect 35100 6500 35156 6502
rect 35180 6500 35236 6502
rect 34794 6296 34850 6352
rect 35622 6296 35678 6352
rect 34940 5466 34996 5468
rect 35020 5466 35076 5468
rect 35100 5466 35156 5468
rect 35180 5466 35236 5468
rect 34940 5414 34966 5466
rect 34966 5414 34996 5466
rect 35020 5414 35030 5466
rect 35030 5414 35076 5466
rect 35100 5414 35146 5466
rect 35146 5414 35156 5466
rect 35180 5414 35210 5466
rect 35210 5414 35236 5466
rect 34940 5412 34996 5414
rect 35020 5412 35076 5414
rect 35100 5412 35156 5414
rect 35180 5412 35236 5414
rect 34940 4378 34996 4380
rect 35020 4378 35076 4380
rect 35100 4378 35156 4380
rect 35180 4378 35236 4380
rect 34940 4326 34966 4378
rect 34966 4326 34996 4378
rect 35020 4326 35030 4378
rect 35030 4326 35076 4378
rect 35100 4326 35146 4378
rect 35146 4326 35156 4378
rect 35180 4326 35210 4378
rect 35210 4326 35236 4378
rect 34940 4324 34996 4326
rect 35020 4324 35076 4326
rect 35100 4324 35156 4326
rect 35180 4324 35236 4326
rect 34794 4120 34850 4176
rect 34940 3290 34996 3292
rect 35020 3290 35076 3292
rect 35100 3290 35156 3292
rect 35180 3290 35236 3292
rect 34940 3238 34966 3290
rect 34966 3238 34996 3290
rect 35020 3238 35030 3290
rect 35030 3238 35076 3290
rect 35100 3238 35146 3290
rect 35146 3238 35156 3290
rect 35180 3238 35210 3290
rect 35210 3238 35236 3290
rect 34940 3236 34996 3238
rect 35020 3236 35076 3238
rect 35100 3236 35156 3238
rect 35180 3236 35236 3238
rect 36726 10240 36782 10296
rect 37278 12180 37280 12200
rect 37280 12180 37332 12200
rect 37332 12180 37334 12200
rect 37278 12144 37334 12180
rect 37922 19352 37978 19408
rect 37922 16396 37924 16416
rect 37924 16396 37976 16416
rect 37976 16396 37978 16416
rect 37922 16360 37978 16396
rect 37554 10512 37610 10568
rect 36542 4684 36598 4720
rect 36542 4664 36544 4684
rect 36544 4664 36596 4684
rect 36596 4664 36598 4684
rect 37738 9560 37794 9616
rect 38106 7112 38162 7168
rect 37922 5636 37978 5672
rect 37922 5616 37924 5636
rect 37924 5616 37976 5636
rect 37976 5616 37978 5636
rect 34940 2202 34996 2204
rect 35020 2202 35076 2204
rect 35100 2202 35156 2204
rect 35180 2202 35236 2204
rect 34940 2150 34966 2202
rect 34966 2150 34996 2202
rect 35020 2150 35030 2202
rect 35030 2150 35076 2202
rect 35100 2150 35146 2202
rect 35146 2150 35156 2202
rect 35180 2150 35210 2202
rect 35210 2150 35236 2202
rect 34940 2148 34996 2150
rect 35020 2148 35076 2150
rect 35100 2148 35156 2150
rect 35180 2148 35236 2150
rect 38106 1128 38162 1184
<< metal3 >>
rect 38101 37634 38167 37637
rect 39200 37634 40000 37664
rect 38101 37632 40000 37634
rect 38101 37576 38106 37632
rect 38162 37576 40000 37632
rect 38101 37574 40000 37576
rect 38101 37571 38167 37574
rect 19568 37568 19888 37569
rect 19568 37504 19576 37568
rect 19640 37504 19656 37568
rect 19720 37504 19736 37568
rect 19800 37504 19816 37568
rect 19880 37504 19888 37568
rect 39200 37544 40000 37574
rect 19568 37503 19888 37504
rect 0 37362 800 37392
rect 2773 37362 2839 37365
rect 0 37360 2839 37362
rect 0 37304 2778 37360
rect 2834 37304 2839 37360
rect 0 37302 2839 37304
rect 0 37272 800 37302
rect 2773 37299 2839 37302
rect 4208 37024 4528 37025
rect 4208 36960 4216 37024
rect 4280 36960 4296 37024
rect 4360 36960 4376 37024
rect 4440 36960 4456 37024
rect 4520 36960 4528 37024
rect 4208 36959 4528 36960
rect 34928 37024 35248 37025
rect 34928 36960 34936 37024
rect 35000 36960 35016 37024
rect 35080 36960 35096 37024
rect 35160 36960 35176 37024
rect 35240 36960 35248 37024
rect 34928 36959 35248 36960
rect 19568 36480 19888 36481
rect 19568 36416 19576 36480
rect 19640 36416 19656 36480
rect 19720 36416 19736 36480
rect 19800 36416 19816 36480
rect 19880 36416 19888 36480
rect 19568 36415 19888 36416
rect 4208 35936 4528 35937
rect 4208 35872 4216 35936
rect 4280 35872 4296 35936
rect 4360 35872 4376 35936
rect 4440 35872 4456 35936
rect 4520 35872 4528 35936
rect 4208 35871 4528 35872
rect 34928 35936 35248 35937
rect 34928 35872 34936 35936
rect 35000 35872 35016 35936
rect 35080 35872 35096 35936
rect 35160 35872 35176 35936
rect 35240 35872 35248 35936
rect 34928 35871 35248 35872
rect 19568 35392 19888 35393
rect 19568 35328 19576 35392
rect 19640 35328 19656 35392
rect 19720 35328 19736 35392
rect 19800 35328 19816 35392
rect 19880 35328 19888 35392
rect 19568 35327 19888 35328
rect 4208 34848 4528 34849
rect 4208 34784 4216 34848
rect 4280 34784 4296 34848
rect 4360 34784 4376 34848
rect 4440 34784 4456 34848
rect 4520 34784 4528 34848
rect 4208 34783 4528 34784
rect 34928 34848 35248 34849
rect 34928 34784 34936 34848
rect 35000 34784 35016 34848
rect 35080 34784 35096 34848
rect 35160 34784 35176 34848
rect 35240 34784 35248 34848
rect 34928 34783 35248 34784
rect 36997 34642 37063 34645
rect 39200 34642 40000 34672
rect 36997 34640 40000 34642
rect 36997 34584 37002 34640
rect 37058 34584 40000 34640
rect 36997 34582 40000 34584
rect 36997 34579 37063 34582
rect 39200 34552 40000 34582
rect 19568 34304 19888 34305
rect 19568 34240 19576 34304
rect 19640 34240 19656 34304
rect 19720 34240 19736 34304
rect 19800 34240 19816 34304
rect 19880 34240 19888 34304
rect 19568 34239 19888 34240
rect 0 34098 800 34128
rect 3785 34098 3851 34101
rect 0 34096 3851 34098
rect 0 34040 3790 34096
rect 3846 34040 3851 34096
rect 0 34038 3851 34040
rect 0 34008 800 34038
rect 3785 34035 3851 34038
rect 4208 33760 4528 33761
rect 4208 33696 4216 33760
rect 4280 33696 4296 33760
rect 4360 33696 4376 33760
rect 4440 33696 4456 33760
rect 4520 33696 4528 33760
rect 4208 33695 4528 33696
rect 34928 33760 35248 33761
rect 34928 33696 34936 33760
rect 35000 33696 35016 33760
rect 35080 33696 35096 33760
rect 35160 33696 35176 33760
rect 35240 33696 35248 33760
rect 34928 33695 35248 33696
rect 7465 33418 7531 33421
rect 8017 33418 8083 33421
rect 9121 33418 9187 33421
rect 7465 33416 9187 33418
rect 7465 33360 7470 33416
rect 7526 33360 8022 33416
rect 8078 33360 9126 33416
rect 9182 33360 9187 33416
rect 7465 33358 9187 33360
rect 7465 33355 7531 33358
rect 8017 33355 8083 33358
rect 9121 33355 9187 33358
rect 19568 33216 19888 33217
rect 19568 33152 19576 33216
rect 19640 33152 19656 33216
rect 19720 33152 19736 33216
rect 19800 33152 19816 33216
rect 19880 33152 19888 33216
rect 19568 33151 19888 33152
rect 4208 32672 4528 32673
rect 4208 32608 4216 32672
rect 4280 32608 4296 32672
rect 4360 32608 4376 32672
rect 4440 32608 4456 32672
rect 4520 32608 4528 32672
rect 4208 32607 4528 32608
rect 34928 32672 35248 32673
rect 34928 32608 34936 32672
rect 35000 32608 35016 32672
rect 35080 32608 35096 32672
rect 35160 32608 35176 32672
rect 35240 32608 35248 32672
rect 34928 32607 35248 32608
rect 19568 32128 19888 32129
rect 19568 32064 19576 32128
rect 19640 32064 19656 32128
rect 19720 32064 19736 32128
rect 19800 32064 19816 32128
rect 19880 32064 19888 32128
rect 19568 32063 19888 32064
rect 35525 31650 35591 31653
rect 39200 31650 40000 31680
rect 35525 31648 40000 31650
rect 35525 31592 35530 31648
rect 35586 31592 40000 31648
rect 35525 31590 40000 31592
rect 35525 31587 35591 31590
rect 4208 31584 4528 31585
rect 4208 31520 4216 31584
rect 4280 31520 4296 31584
rect 4360 31520 4376 31584
rect 4440 31520 4456 31584
rect 4520 31520 4528 31584
rect 4208 31519 4528 31520
rect 34928 31584 35248 31585
rect 34928 31520 34936 31584
rect 35000 31520 35016 31584
rect 35080 31520 35096 31584
rect 35160 31520 35176 31584
rect 35240 31520 35248 31584
rect 39200 31560 40000 31590
rect 34928 31519 35248 31520
rect 2129 31242 2195 31245
rect 3141 31242 3207 31245
rect 4429 31242 4495 31245
rect 2129 31240 4495 31242
rect 2129 31184 2134 31240
rect 2190 31184 3146 31240
rect 3202 31184 4434 31240
rect 4490 31184 4495 31240
rect 2129 31182 4495 31184
rect 2129 31179 2195 31182
rect 3141 31179 3207 31182
rect 4429 31179 4495 31182
rect 0 31106 800 31136
rect 1945 31106 2011 31109
rect 0 31104 2011 31106
rect 0 31048 1950 31104
rect 2006 31048 2011 31104
rect 0 31046 2011 31048
rect 0 31016 800 31046
rect 1945 31043 2011 31046
rect 19568 31040 19888 31041
rect 19568 30976 19576 31040
rect 19640 30976 19656 31040
rect 19720 30976 19736 31040
rect 19800 30976 19816 31040
rect 19880 30976 19888 31040
rect 19568 30975 19888 30976
rect 4208 30496 4528 30497
rect 4208 30432 4216 30496
rect 4280 30432 4296 30496
rect 4360 30432 4376 30496
rect 4440 30432 4456 30496
rect 4520 30432 4528 30496
rect 4208 30431 4528 30432
rect 34928 30496 35248 30497
rect 34928 30432 34936 30496
rect 35000 30432 35016 30496
rect 35080 30432 35096 30496
rect 35160 30432 35176 30496
rect 35240 30432 35248 30496
rect 34928 30431 35248 30432
rect 24485 30428 24551 30429
rect 24485 30424 24532 30428
rect 24596 30426 24602 30428
rect 24485 30368 24490 30424
rect 24485 30364 24532 30368
rect 24596 30366 24642 30426
rect 24596 30364 24602 30366
rect 24485 30363 24551 30364
rect 10593 30154 10659 30157
rect 17033 30154 17099 30157
rect 17769 30154 17835 30157
rect 10593 30152 17835 30154
rect 10593 30096 10598 30152
rect 10654 30096 17038 30152
rect 17094 30096 17774 30152
rect 17830 30096 17835 30152
rect 10593 30094 17835 30096
rect 10593 30091 10659 30094
rect 17033 30091 17099 30094
rect 17769 30091 17835 30094
rect 19568 29952 19888 29953
rect 19568 29888 19576 29952
rect 19640 29888 19656 29952
rect 19720 29888 19736 29952
rect 19800 29888 19816 29952
rect 19880 29888 19888 29952
rect 19568 29887 19888 29888
rect 19701 29610 19767 29613
rect 23289 29610 23355 29613
rect 19701 29608 23355 29610
rect 19701 29552 19706 29608
rect 19762 29552 23294 29608
rect 23350 29552 23355 29608
rect 19701 29550 23355 29552
rect 19701 29547 19767 29550
rect 23289 29547 23355 29550
rect 4208 29408 4528 29409
rect 4208 29344 4216 29408
rect 4280 29344 4296 29408
rect 4360 29344 4376 29408
rect 4440 29344 4456 29408
rect 4520 29344 4528 29408
rect 4208 29343 4528 29344
rect 34928 29408 35248 29409
rect 34928 29344 34936 29408
rect 35000 29344 35016 29408
rect 35080 29344 35096 29408
rect 35160 29344 35176 29408
rect 35240 29344 35248 29408
rect 34928 29343 35248 29344
rect 36261 29066 36327 29069
rect 36126 29064 36327 29066
rect 36126 29008 36266 29064
rect 36322 29008 36327 29064
rect 36126 29006 36327 29008
rect 19568 28864 19888 28865
rect 19568 28800 19576 28864
rect 19640 28800 19656 28864
rect 19720 28800 19736 28864
rect 19800 28800 19816 28864
rect 19880 28800 19888 28864
rect 19568 28799 19888 28800
rect 32581 28794 32647 28797
rect 36126 28794 36186 29006
rect 36261 29003 36327 29006
rect 32581 28792 36186 28794
rect 32581 28736 32586 28792
rect 32642 28736 36186 28792
rect 32581 28734 36186 28736
rect 32581 28731 32647 28734
rect 37917 28386 37983 28389
rect 39200 28386 40000 28416
rect 37917 28384 40000 28386
rect 37917 28328 37922 28384
rect 37978 28328 40000 28384
rect 37917 28326 40000 28328
rect 37917 28323 37983 28326
rect 4208 28320 4528 28321
rect 4208 28256 4216 28320
rect 4280 28256 4296 28320
rect 4360 28256 4376 28320
rect 4440 28256 4456 28320
rect 4520 28256 4528 28320
rect 4208 28255 4528 28256
rect 34928 28320 35248 28321
rect 34928 28256 34936 28320
rect 35000 28256 35016 28320
rect 35080 28256 35096 28320
rect 35160 28256 35176 28320
rect 35240 28256 35248 28320
rect 39200 28296 40000 28326
rect 34928 28255 35248 28256
rect 0 28114 800 28144
rect 3049 28114 3115 28117
rect 0 28112 3115 28114
rect 0 28056 3054 28112
rect 3110 28056 3115 28112
rect 0 28054 3115 28056
rect 0 28024 800 28054
rect 3049 28051 3115 28054
rect 19568 27776 19888 27777
rect 19568 27712 19576 27776
rect 19640 27712 19656 27776
rect 19720 27712 19736 27776
rect 19800 27712 19816 27776
rect 19880 27712 19888 27776
rect 19568 27711 19888 27712
rect 4208 27232 4528 27233
rect 4208 27168 4216 27232
rect 4280 27168 4296 27232
rect 4360 27168 4376 27232
rect 4440 27168 4456 27232
rect 4520 27168 4528 27232
rect 4208 27167 4528 27168
rect 34928 27232 35248 27233
rect 34928 27168 34936 27232
rect 35000 27168 35016 27232
rect 35080 27168 35096 27232
rect 35160 27168 35176 27232
rect 35240 27168 35248 27232
rect 34928 27167 35248 27168
rect 20713 26890 20779 26893
rect 22093 26890 22159 26893
rect 20713 26888 22159 26890
rect 20713 26832 20718 26888
rect 20774 26832 22098 26888
rect 22154 26832 22159 26888
rect 20713 26830 22159 26832
rect 20713 26827 20779 26830
rect 22093 26827 22159 26830
rect 19568 26688 19888 26689
rect 19568 26624 19576 26688
rect 19640 26624 19656 26688
rect 19720 26624 19736 26688
rect 19800 26624 19816 26688
rect 19880 26624 19888 26688
rect 19568 26623 19888 26624
rect 19701 26482 19767 26485
rect 20069 26482 20135 26485
rect 22829 26482 22895 26485
rect 19701 26480 22895 26482
rect 19701 26424 19706 26480
rect 19762 26424 20074 26480
rect 20130 26424 22834 26480
rect 22890 26424 22895 26480
rect 19701 26422 22895 26424
rect 19701 26419 19767 26422
rect 20069 26419 20135 26422
rect 22829 26419 22895 26422
rect 4208 26144 4528 26145
rect 4208 26080 4216 26144
rect 4280 26080 4296 26144
rect 4360 26080 4376 26144
rect 4440 26080 4456 26144
rect 4520 26080 4528 26144
rect 4208 26079 4528 26080
rect 34928 26144 35248 26145
rect 34928 26080 34936 26144
rect 35000 26080 35016 26144
rect 35080 26080 35096 26144
rect 35160 26080 35176 26144
rect 35240 26080 35248 26144
rect 34928 26079 35248 26080
rect 19568 25600 19888 25601
rect 19568 25536 19576 25600
rect 19640 25536 19656 25600
rect 19720 25536 19736 25600
rect 19800 25536 19816 25600
rect 19880 25536 19888 25600
rect 19568 25535 19888 25536
rect 35433 25394 35499 25397
rect 39200 25394 40000 25424
rect 35433 25392 40000 25394
rect 35433 25336 35438 25392
rect 35494 25336 40000 25392
rect 35433 25334 40000 25336
rect 35433 25331 35499 25334
rect 39200 25304 40000 25334
rect 0 25122 800 25152
rect 3969 25122 4035 25125
rect 0 25120 4035 25122
rect 0 25064 3974 25120
rect 4030 25064 4035 25120
rect 0 25062 4035 25064
rect 0 25032 800 25062
rect 3969 25059 4035 25062
rect 4208 25056 4528 25057
rect 4208 24992 4216 25056
rect 4280 24992 4296 25056
rect 4360 24992 4376 25056
rect 4440 24992 4456 25056
rect 4520 24992 4528 25056
rect 4208 24991 4528 24992
rect 34928 25056 35248 25057
rect 34928 24992 34936 25056
rect 35000 24992 35016 25056
rect 35080 24992 35096 25056
rect 35160 24992 35176 25056
rect 35240 24992 35248 25056
rect 34928 24991 35248 24992
rect 24393 24988 24459 24989
rect 24342 24986 24348 24988
rect 24302 24926 24348 24986
rect 24412 24984 24459 24988
rect 24454 24928 24459 24984
rect 24342 24924 24348 24926
rect 24412 24924 24459 24928
rect 24393 24923 24459 24924
rect 33961 24714 34027 24717
rect 36537 24714 36603 24717
rect 33961 24712 36603 24714
rect 33961 24656 33966 24712
rect 34022 24656 36542 24712
rect 36598 24656 36603 24712
rect 33961 24654 36603 24656
rect 33961 24651 34027 24654
rect 36537 24651 36603 24654
rect 19568 24512 19888 24513
rect 19568 24448 19576 24512
rect 19640 24448 19656 24512
rect 19720 24448 19736 24512
rect 19800 24448 19816 24512
rect 19880 24448 19888 24512
rect 19568 24447 19888 24448
rect 4208 23968 4528 23969
rect 4208 23904 4216 23968
rect 4280 23904 4296 23968
rect 4360 23904 4376 23968
rect 4440 23904 4456 23968
rect 4520 23904 4528 23968
rect 4208 23903 4528 23904
rect 34928 23968 35248 23969
rect 34928 23904 34936 23968
rect 35000 23904 35016 23968
rect 35080 23904 35096 23968
rect 35160 23904 35176 23968
rect 35240 23904 35248 23968
rect 34928 23903 35248 23904
rect 19568 23424 19888 23425
rect 19568 23360 19576 23424
rect 19640 23360 19656 23424
rect 19720 23360 19736 23424
rect 19800 23360 19816 23424
rect 19880 23360 19888 23424
rect 19568 23359 19888 23360
rect 4208 22880 4528 22881
rect 4208 22816 4216 22880
rect 4280 22816 4296 22880
rect 4360 22816 4376 22880
rect 4440 22816 4456 22880
rect 4520 22816 4528 22880
rect 4208 22815 4528 22816
rect 34928 22880 35248 22881
rect 34928 22816 34936 22880
rect 35000 22816 35016 22880
rect 35080 22816 35096 22880
rect 35160 22816 35176 22880
rect 35240 22816 35248 22880
rect 34928 22815 35248 22816
rect 29821 22674 29887 22677
rect 35341 22674 35407 22677
rect 29821 22672 35407 22674
rect 29821 22616 29826 22672
rect 29882 22616 35346 22672
rect 35402 22616 35407 22672
rect 29821 22614 35407 22616
rect 29821 22611 29887 22614
rect 35341 22611 35407 22614
rect 35525 22402 35591 22405
rect 39200 22402 40000 22432
rect 35525 22400 40000 22402
rect 35525 22344 35530 22400
rect 35586 22344 40000 22400
rect 35525 22342 40000 22344
rect 35525 22339 35591 22342
rect 19568 22336 19888 22337
rect 19568 22272 19576 22336
rect 19640 22272 19656 22336
rect 19720 22272 19736 22336
rect 19800 22272 19816 22336
rect 19880 22272 19888 22336
rect 39200 22312 40000 22342
rect 19568 22271 19888 22272
rect 0 22130 800 22160
rect 2773 22130 2839 22133
rect 0 22128 2839 22130
rect 0 22072 2778 22128
rect 2834 22072 2839 22128
rect 0 22070 2839 22072
rect 0 22040 800 22070
rect 2773 22067 2839 22070
rect 12433 22130 12499 22133
rect 12893 22130 12959 22133
rect 12433 22128 12959 22130
rect 12433 22072 12438 22128
rect 12494 22072 12898 22128
rect 12954 22072 12959 22128
rect 12433 22070 12959 22072
rect 12433 22067 12499 22070
rect 12893 22067 12959 22070
rect 3417 21994 3483 21997
rect 18413 21994 18479 21997
rect 3417 21992 18479 21994
rect 3417 21936 3422 21992
rect 3478 21936 18418 21992
rect 18474 21936 18479 21992
rect 3417 21934 18479 21936
rect 3417 21931 3483 21934
rect 18413 21931 18479 21934
rect 9489 21858 9555 21861
rect 20069 21858 20135 21861
rect 20989 21858 21055 21861
rect 9489 21856 21055 21858
rect 9489 21800 9494 21856
rect 9550 21800 20074 21856
rect 20130 21800 20994 21856
rect 21050 21800 21055 21856
rect 9489 21798 21055 21800
rect 9489 21795 9555 21798
rect 20069 21795 20135 21798
rect 20989 21795 21055 21798
rect 4208 21792 4528 21793
rect 4208 21728 4216 21792
rect 4280 21728 4296 21792
rect 4360 21728 4376 21792
rect 4440 21728 4456 21792
rect 4520 21728 4528 21792
rect 4208 21727 4528 21728
rect 34928 21792 35248 21793
rect 34928 21728 34936 21792
rect 35000 21728 35016 21792
rect 35080 21728 35096 21792
rect 35160 21728 35176 21792
rect 35240 21728 35248 21792
rect 34928 21727 35248 21728
rect 14365 21586 14431 21589
rect 19425 21586 19491 21589
rect 14365 21584 19491 21586
rect 14365 21528 14370 21584
rect 14426 21528 19430 21584
rect 19486 21528 19491 21584
rect 14365 21526 19491 21528
rect 14365 21523 14431 21526
rect 19425 21523 19491 21526
rect 30557 21586 30623 21589
rect 30925 21586 30991 21589
rect 30557 21584 30991 21586
rect 30557 21528 30562 21584
rect 30618 21528 30930 21584
rect 30986 21528 30991 21584
rect 30557 21526 30991 21528
rect 30557 21523 30623 21526
rect 30925 21523 30991 21526
rect 19568 21248 19888 21249
rect 19568 21184 19576 21248
rect 19640 21184 19656 21248
rect 19720 21184 19736 21248
rect 19800 21184 19816 21248
rect 19880 21184 19888 21248
rect 19568 21183 19888 21184
rect 4208 20704 4528 20705
rect 4208 20640 4216 20704
rect 4280 20640 4296 20704
rect 4360 20640 4376 20704
rect 4440 20640 4456 20704
rect 4520 20640 4528 20704
rect 4208 20639 4528 20640
rect 34928 20704 35248 20705
rect 34928 20640 34936 20704
rect 35000 20640 35016 20704
rect 35080 20640 35096 20704
rect 35160 20640 35176 20704
rect 35240 20640 35248 20704
rect 34928 20639 35248 20640
rect 19568 20160 19888 20161
rect 19568 20096 19576 20160
rect 19640 20096 19656 20160
rect 19720 20096 19736 20160
rect 19800 20096 19816 20160
rect 19880 20096 19888 20160
rect 19568 20095 19888 20096
rect 21633 19682 21699 19685
rect 22093 19682 22159 19685
rect 25221 19682 25287 19685
rect 21633 19680 25287 19682
rect 21633 19624 21638 19680
rect 21694 19624 22098 19680
rect 22154 19624 25226 19680
rect 25282 19624 25287 19680
rect 21633 19622 25287 19624
rect 21633 19619 21699 19622
rect 22093 19619 22159 19622
rect 25221 19619 25287 19622
rect 4208 19616 4528 19617
rect 4208 19552 4216 19616
rect 4280 19552 4296 19616
rect 4360 19552 4376 19616
rect 4440 19552 4456 19616
rect 4520 19552 4528 19616
rect 4208 19551 4528 19552
rect 34928 19616 35248 19617
rect 34928 19552 34936 19616
rect 35000 19552 35016 19616
rect 35080 19552 35096 19616
rect 35160 19552 35176 19616
rect 35240 19552 35248 19616
rect 34928 19551 35248 19552
rect 3969 19410 4035 19413
rect 7925 19410 7991 19413
rect 3969 19408 7991 19410
rect 3969 19352 3974 19408
rect 4030 19352 7930 19408
rect 7986 19352 7991 19408
rect 3969 19350 7991 19352
rect 3969 19347 4035 19350
rect 7925 19347 7991 19350
rect 26509 19410 26575 19413
rect 27337 19410 27403 19413
rect 26509 19408 27403 19410
rect 26509 19352 26514 19408
rect 26570 19352 27342 19408
rect 27398 19352 27403 19408
rect 26509 19350 27403 19352
rect 26509 19347 26575 19350
rect 27337 19347 27403 19350
rect 37917 19410 37983 19413
rect 39200 19410 40000 19440
rect 37917 19408 40000 19410
rect 37917 19352 37922 19408
rect 37978 19352 40000 19408
rect 37917 19350 40000 19352
rect 37917 19347 37983 19350
rect 39200 19320 40000 19350
rect 12433 19274 12499 19277
rect 18045 19274 18111 19277
rect 12433 19272 18111 19274
rect 12433 19216 12438 19272
rect 12494 19216 18050 19272
rect 18106 19216 18111 19272
rect 12433 19214 18111 19216
rect 12433 19211 12499 19214
rect 18045 19211 18111 19214
rect 25037 19274 25103 19277
rect 27245 19274 27311 19277
rect 25037 19272 27311 19274
rect 25037 19216 25042 19272
rect 25098 19216 27250 19272
rect 27306 19216 27311 19272
rect 25037 19214 27311 19216
rect 25037 19211 25103 19214
rect 27245 19211 27311 19214
rect 0 19138 800 19168
rect 4061 19138 4127 19141
rect 0 19136 4127 19138
rect 0 19080 4066 19136
rect 4122 19080 4127 19136
rect 0 19078 4127 19080
rect 0 19048 800 19078
rect 4061 19075 4127 19078
rect 21265 19138 21331 19141
rect 22001 19138 22067 19141
rect 27889 19138 27955 19141
rect 21265 19136 27955 19138
rect 21265 19080 21270 19136
rect 21326 19080 22006 19136
rect 22062 19080 27894 19136
rect 27950 19080 27955 19136
rect 21265 19078 27955 19080
rect 21265 19075 21331 19078
rect 22001 19075 22067 19078
rect 27889 19075 27955 19078
rect 19568 19072 19888 19073
rect 19568 19008 19576 19072
rect 19640 19008 19656 19072
rect 19720 19008 19736 19072
rect 19800 19008 19816 19072
rect 19880 19008 19888 19072
rect 19568 19007 19888 19008
rect 26969 18866 27035 18869
rect 27613 18866 27679 18869
rect 26969 18864 27679 18866
rect 26969 18808 26974 18864
rect 27030 18808 27618 18864
rect 27674 18808 27679 18864
rect 26969 18806 27679 18808
rect 26969 18803 27035 18806
rect 27613 18803 27679 18806
rect 20345 18730 20411 18733
rect 26601 18730 26667 18733
rect 20345 18728 26667 18730
rect 20345 18672 20350 18728
rect 20406 18672 26606 18728
rect 26662 18672 26667 18728
rect 20345 18670 26667 18672
rect 20345 18667 20411 18670
rect 26601 18667 26667 18670
rect 4208 18528 4528 18529
rect 4208 18464 4216 18528
rect 4280 18464 4296 18528
rect 4360 18464 4376 18528
rect 4440 18464 4456 18528
rect 4520 18464 4528 18528
rect 4208 18463 4528 18464
rect 34928 18528 35248 18529
rect 34928 18464 34936 18528
rect 35000 18464 35016 18528
rect 35080 18464 35096 18528
rect 35160 18464 35176 18528
rect 35240 18464 35248 18528
rect 34928 18463 35248 18464
rect 19568 17984 19888 17985
rect 19568 17920 19576 17984
rect 19640 17920 19656 17984
rect 19720 17920 19736 17984
rect 19800 17920 19816 17984
rect 19880 17920 19888 17984
rect 19568 17919 19888 17920
rect 4208 17440 4528 17441
rect 4208 17376 4216 17440
rect 4280 17376 4296 17440
rect 4360 17376 4376 17440
rect 4440 17376 4456 17440
rect 4520 17376 4528 17440
rect 4208 17375 4528 17376
rect 34928 17440 35248 17441
rect 34928 17376 34936 17440
rect 35000 17376 35016 17440
rect 35080 17376 35096 17440
rect 35160 17376 35176 17440
rect 35240 17376 35248 17440
rect 34928 17375 35248 17376
rect 26509 17098 26575 17101
rect 28257 17098 28323 17101
rect 26509 17096 28323 17098
rect 26509 17040 26514 17096
rect 26570 17040 28262 17096
rect 28318 17040 28323 17096
rect 26509 17038 28323 17040
rect 26509 17035 26575 17038
rect 28257 17035 28323 17038
rect 19568 16896 19888 16897
rect 19568 16832 19576 16896
rect 19640 16832 19656 16896
rect 19720 16832 19736 16896
rect 19800 16832 19816 16896
rect 19880 16832 19888 16896
rect 19568 16831 19888 16832
rect 27797 16690 27863 16693
rect 28993 16690 29059 16693
rect 27797 16688 29059 16690
rect 27797 16632 27802 16688
rect 27858 16632 28998 16688
rect 29054 16632 29059 16688
rect 27797 16630 29059 16632
rect 27797 16627 27863 16630
rect 28993 16627 29059 16630
rect 37917 16418 37983 16421
rect 39200 16418 40000 16448
rect 37917 16416 40000 16418
rect 37917 16360 37922 16416
rect 37978 16360 40000 16416
rect 37917 16358 40000 16360
rect 37917 16355 37983 16358
rect 4208 16352 4528 16353
rect 4208 16288 4216 16352
rect 4280 16288 4296 16352
rect 4360 16288 4376 16352
rect 4440 16288 4456 16352
rect 4520 16288 4528 16352
rect 4208 16287 4528 16288
rect 34928 16352 35248 16353
rect 34928 16288 34936 16352
rect 35000 16288 35016 16352
rect 35080 16288 35096 16352
rect 35160 16288 35176 16352
rect 35240 16288 35248 16352
rect 39200 16328 40000 16358
rect 34928 16287 35248 16288
rect 24761 16146 24827 16149
rect 34973 16146 35039 16149
rect 24761 16144 35039 16146
rect 24761 16088 24766 16144
rect 24822 16088 34978 16144
rect 35034 16088 35039 16144
rect 24761 16086 35039 16088
rect 24761 16083 24827 16086
rect 34973 16083 35039 16086
rect 21449 16010 21515 16013
rect 30373 16010 30439 16013
rect 21449 16008 30439 16010
rect 21449 15952 21454 16008
rect 21510 15952 30378 16008
rect 30434 15952 30439 16008
rect 21449 15950 30439 15952
rect 21449 15947 21515 15950
rect 30373 15947 30439 15950
rect 0 15874 800 15904
rect 4061 15874 4127 15877
rect 0 15872 4127 15874
rect 0 15816 4066 15872
rect 4122 15816 4127 15872
rect 0 15814 4127 15816
rect 0 15784 800 15814
rect 4061 15811 4127 15814
rect 19568 15808 19888 15809
rect 19568 15744 19576 15808
rect 19640 15744 19656 15808
rect 19720 15744 19736 15808
rect 19800 15744 19816 15808
rect 19880 15744 19888 15808
rect 19568 15743 19888 15744
rect 4208 15264 4528 15265
rect 4208 15200 4216 15264
rect 4280 15200 4296 15264
rect 4360 15200 4376 15264
rect 4440 15200 4456 15264
rect 4520 15200 4528 15264
rect 4208 15199 4528 15200
rect 34928 15264 35248 15265
rect 34928 15200 34936 15264
rect 35000 15200 35016 15264
rect 35080 15200 35096 15264
rect 35160 15200 35176 15264
rect 35240 15200 35248 15264
rect 34928 15199 35248 15200
rect 5901 15194 5967 15197
rect 9857 15194 9923 15197
rect 5901 15192 9923 15194
rect 5901 15136 5906 15192
rect 5962 15136 9862 15192
rect 9918 15136 9923 15192
rect 5901 15134 9923 15136
rect 5901 15131 5967 15134
rect 9857 15131 9923 15134
rect 14457 15194 14523 15197
rect 16941 15194 17007 15197
rect 14457 15192 17007 15194
rect 14457 15136 14462 15192
rect 14518 15136 16946 15192
rect 17002 15136 17007 15192
rect 14457 15134 17007 15136
rect 14457 15131 14523 15134
rect 16941 15131 17007 15134
rect 6821 15058 6887 15061
rect 15285 15058 15351 15061
rect 6821 15056 15351 15058
rect 6821 15000 6826 15056
rect 6882 15000 15290 15056
rect 15346 15000 15351 15056
rect 6821 14998 15351 15000
rect 6821 14995 6887 14998
rect 15285 14995 15351 14998
rect 19568 14720 19888 14721
rect 19568 14656 19576 14720
rect 19640 14656 19656 14720
rect 19720 14656 19736 14720
rect 19800 14656 19816 14720
rect 19880 14656 19888 14720
rect 19568 14655 19888 14656
rect 13169 14514 13235 14517
rect 19885 14514 19951 14517
rect 13169 14512 19951 14514
rect 13169 14456 13174 14512
rect 13230 14456 19890 14512
rect 19946 14456 19951 14512
rect 13169 14454 19951 14456
rect 13169 14451 13235 14454
rect 19885 14451 19951 14454
rect 3141 14378 3207 14381
rect 17493 14378 17559 14381
rect 3141 14376 17559 14378
rect 3141 14320 3146 14376
rect 3202 14320 17498 14376
rect 17554 14320 17559 14376
rect 3141 14318 17559 14320
rect 3141 14315 3207 14318
rect 17493 14315 17559 14318
rect 4208 14176 4528 14177
rect 4208 14112 4216 14176
rect 4280 14112 4296 14176
rect 4360 14112 4376 14176
rect 4440 14112 4456 14176
rect 4520 14112 4528 14176
rect 4208 14111 4528 14112
rect 34928 14176 35248 14177
rect 34928 14112 34936 14176
rect 35000 14112 35016 14176
rect 35080 14112 35096 14176
rect 35160 14112 35176 14176
rect 35240 14112 35248 14176
rect 34928 14111 35248 14112
rect 19568 13632 19888 13633
rect 19568 13568 19576 13632
rect 19640 13568 19656 13632
rect 19720 13568 19736 13632
rect 19800 13568 19816 13632
rect 19880 13568 19888 13632
rect 19568 13567 19888 13568
rect 2865 13426 2931 13429
rect 22553 13426 22619 13429
rect 2865 13424 22619 13426
rect 2865 13368 2870 13424
rect 2926 13368 22558 13424
rect 22614 13368 22619 13424
rect 2865 13366 22619 13368
rect 2865 13363 2931 13366
rect 22553 13363 22619 13366
rect 35249 13426 35315 13429
rect 39200 13426 40000 13456
rect 35249 13424 40000 13426
rect 35249 13368 35254 13424
rect 35310 13368 40000 13424
rect 35249 13366 40000 13368
rect 35249 13363 35315 13366
rect 39200 13336 40000 13366
rect 4208 13088 4528 13089
rect 4208 13024 4216 13088
rect 4280 13024 4296 13088
rect 4360 13024 4376 13088
rect 4440 13024 4456 13088
rect 4520 13024 4528 13088
rect 4208 13023 4528 13024
rect 34928 13088 35248 13089
rect 34928 13024 34936 13088
rect 35000 13024 35016 13088
rect 35080 13024 35096 13088
rect 35160 13024 35176 13088
rect 35240 13024 35248 13088
rect 34928 13023 35248 13024
rect 0 12882 800 12912
rect 2681 12882 2747 12885
rect 0 12880 2747 12882
rect 0 12824 2686 12880
rect 2742 12824 2747 12880
rect 0 12822 2747 12824
rect 0 12792 800 12822
rect 2681 12819 2747 12822
rect 8753 12882 8819 12885
rect 11329 12882 11395 12885
rect 8753 12880 11395 12882
rect 8753 12824 8758 12880
rect 8814 12824 11334 12880
rect 11390 12824 11395 12880
rect 8753 12822 11395 12824
rect 8753 12819 8819 12822
rect 11329 12819 11395 12822
rect 10685 12746 10751 12749
rect 16757 12746 16823 12749
rect 10685 12744 16823 12746
rect 10685 12688 10690 12744
rect 10746 12688 16762 12744
rect 16818 12688 16823 12744
rect 10685 12686 16823 12688
rect 10685 12683 10751 12686
rect 16757 12683 16823 12686
rect 19568 12544 19888 12545
rect 19568 12480 19576 12544
rect 19640 12480 19656 12544
rect 19720 12480 19736 12544
rect 19800 12480 19816 12544
rect 19880 12480 19888 12544
rect 19568 12479 19888 12480
rect 18413 12202 18479 12205
rect 37273 12202 37339 12205
rect 18413 12200 37339 12202
rect 18413 12144 18418 12200
rect 18474 12144 37278 12200
rect 37334 12144 37339 12200
rect 18413 12142 37339 12144
rect 18413 12139 18479 12142
rect 37273 12139 37339 12142
rect 31293 12066 31359 12069
rect 33409 12066 33475 12069
rect 31293 12064 33475 12066
rect 31293 12008 31298 12064
rect 31354 12008 33414 12064
rect 33470 12008 33475 12064
rect 31293 12006 33475 12008
rect 31293 12003 31359 12006
rect 33409 12003 33475 12006
rect 4208 12000 4528 12001
rect 4208 11936 4216 12000
rect 4280 11936 4296 12000
rect 4360 11936 4376 12000
rect 4440 11936 4456 12000
rect 4520 11936 4528 12000
rect 4208 11935 4528 11936
rect 34928 12000 35248 12001
rect 34928 11936 34936 12000
rect 35000 11936 35016 12000
rect 35080 11936 35096 12000
rect 35160 11936 35176 12000
rect 35240 11936 35248 12000
rect 34928 11935 35248 11936
rect 14733 11658 14799 11661
rect 18781 11658 18847 11661
rect 14733 11656 18847 11658
rect 14733 11600 14738 11656
rect 14794 11600 18786 11656
rect 18842 11600 18847 11656
rect 14733 11598 18847 11600
rect 14733 11595 14799 11598
rect 18781 11595 18847 11598
rect 29177 11658 29243 11661
rect 31937 11658 32003 11661
rect 29177 11656 32003 11658
rect 29177 11600 29182 11656
rect 29238 11600 31942 11656
rect 31998 11600 32003 11656
rect 29177 11598 32003 11600
rect 29177 11595 29243 11598
rect 31937 11595 32003 11598
rect 19568 11456 19888 11457
rect 19568 11392 19576 11456
rect 19640 11392 19656 11456
rect 19720 11392 19736 11456
rect 19800 11392 19816 11456
rect 19880 11392 19888 11456
rect 19568 11391 19888 11392
rect 29177 11250 29243 11253
rect 30189 11250 30255 11253
rect 29177 11248 30255 11250
rect 29177 11192 29182 11248
rect 29238 11192 30194 11248
rect 30250 11192 30255 11248
rect 29177 11190 30255 11192
rect 29177 11187 29243 11190
rect 30189 11187 30255 11190
rect 12709 11114 12775 11117
rect 21909 11114 21975 11117
rect 31845 11114 31911 11117
rect 12709 11112 31911 11114
rect 12709 11056 12714 11112
rect 12770 11056 21914 11112
rect 21970 11056 31850 11112
rect 31906 11056 31911 11112
rect 12709 11054 31911 11056
rect 12709 11051 12775 11054
rect 21909 11051 21975 11054
rect 31845 11051 31911 11054
rect 4208 10912 4528 10913
rect 4208 10848 4216 10912
rect 4280 10848 4296 10912
rect 4360 10848 4376 10912
rect 4440 10848 4456 10912
rect 4520 10848 4528 10912
rect 4208 10847 4528 10848
rect 34928 10912 35248 10913
rect 34928 10848 34936 10912
rect 35000 10848 35016 10912
rect 35080 10848 35096 10912
rect 35160 10848 35176 10912
rect 35240 10848 35248 10912
rect 34928 10847 35248 10848
rect 11053 10842 11119 10845
rect 15837 10842 15903 10845
rect 11053 10840 15903 10842
rect 11053 10784 11058 10840
rect 11114 10784 15842 10840
rect 15898 10784 15903 10840
rect 11053 10782 15903 10784
rect 11053 10779 11119 10782
rect 15837 10779 15903 10782
rect 3601 10570 3667 10573
rect 29269 10570 29335 10573
rect 3601 10568 29335 10570
rect 3601 10512 3606 10568
rect 3662 10512 29274 10568
rect 29330 10512 29335 10568
rect 3601 10510 29335 10512
rect 3601 10507 3667 10510
rect 29269 10507 29335 10510
rect 32581 10570 32647 10573
rect 37549 10570 37615 10573
rect 32581 10568 37615 10570
rect 32581 10512 32586 10568
rect 32642 10512 37554 10568
rect 37610 10512 37615 10568
rect 32581 10510 37615 10512
rect 32581 10507 32647 10510
rect 37549 10507 37615 10510
rect 9857 10434 9923 10437
rect 15009 10434 15075 10437
rect 9857 10432 15075 10434
rect 9857 10376 9862 10432
rect 9918 10376 15014 10432
rect 15070 10376 15075 10432
rect 9857 10374 15075 10376
rect 9857 10371 9923 10374
rect 15009 10371 15075 10374
rect 30557 10434 30623 10437
rect 34329 10434 34395 10437
rect 30557 10432 34395 10434
rect 30557 10376 30562 10432
rect 30618 10376 34334 10432
rect 34390 10376 34395 10432
rect 30557 10374 34395 10376
rect 30557 10371 30623 10374
rect 34329 10371 34395 10374
rect 19568 10368 19888 10369
rect 19568 10304 19576 10368
rect 19640 10304 19656 10368
rect 19720 10304 19736 10368
rect 19800 10304 19816 10368
rect 19880 10304 19888 10368
rect 19568 10303 19888 10304
rect 36721 10298 36787 10301
rect 24166 10296 36787 10298
rect 24166 10240 36726 10296
rect 36782 10240 36787 10296
rect 24166 10238 36787 10240
rect 16205 10162 16271 10165
rect 24166 10162 24226 10238
rect 36721 10235 36787 10238
rect 39200 10162 40000 10192
rect 16205 10160 24226 10162
rect 16205 10104 16210 10160
rect 16266 10104 24226 10160
rect 16205 10102 24226 10104
rect 31894 10102 40000 10162
rect 16205 10099 16271 10102
rect 11697 10026 11763 10029
rect 31894 10026 31954 10102
rect 39200 10072 40000 10102
rect 11697 10024 31954 10026
rect 11697 9968 11702 10024
rect 11758 9968 31954 10024
rect 11697 9966 31954 9968
rect 11697 9963 11763 9966
rect 0 9890 800 9920
rect 2773 9890 2839 9893
rect 0 9888 2839 9890
rect 0 9832 2778 9888
rect 2834 9832 2839 9888
rect 0 9830 2839 9832
rect 0 9800 800 9830
rect 2773 9827 2839 9830
rect 4208 9824 4528 9825
rect 4208 9760 4216 9824
rect 4280 9760 4296 9824
rect 4360 9760 4376 9824
rect 4440 9760 4456 9824
rect 4520 9760 4528 9824
rect 4208 9759 4528 9760
rect 34928 9824 35248 9825
rect 34928 9760 34936 9824
rect 35000 9760 35016 9824
rect 35080 9760 35096 9824
rect 35160 9760 35176 9824
rect 35240 9760 35248 9824
rect 34928 9759 35248 9760
rect 29729 9754 29795 9757
rect 31477 9754 31543 9757
rect 29729 9752 31543 9754
rect 29729 9696 29734 9752
rect 29790 9696 31482 9752
rect 31538 9696 31543 9752
rect 29729 9694 31543 9696
rect 29729 9691 29795 9694
rect 31477 9691 31543 9694
rect 28441 9618 28507 9621
rect 37733 9618 37799 9621
rect 28441 9616 37799 9618
rect 28441 9560 28446 9616
rect 28502 9560 37738 9616
rect 37794 9560 37799 9616
rect 28441 9558 37799 9560
rect 28441 9555 28507 9558
rect 37733 9555 37799 9558
rect 19568 9280 19888 9281
rect 19568 9216 19576 9280
rect 19640 9216 19656 9280
rect 19720 9216 19736 9280
rect 19800 9216 19816 9280
rect 19880 9216 19888 9280
rect 19568 9215 19888 9216
rect 15561 9210 15627 9213
rect 18965 9210 19031 9213
rect 15561 9208 19031 9210
rect 15561 9152 15566 9208
rect 15622 9152 18970 9208
rect 19026 9152 19031 9208
rect 15561 9150 19031 9152
rect 15561 9147 15627 9150
rect 18965 9147 19031 9150
rect 6821 9074 6887 9077
rect 16757 9074 16823 9077
rect 6821 9072 16823 9074
rect 6821 9016 6826 9072
rect 6882 9016 16762 9072
rect 16818 9016 16823 9072
rect 6821 9014 16823 9016
rect 6821 9011 6887 9014
rect 16757 9011 16823 9014
rect 19425 9074 19491 9077
rect 22369 9074 22435 9077
rect 19425 9072 22435 9074
rect 19425 9016 19430 9072
rect 19486 9016 22374 9072
rect 22430 9016 22435 9072
rect 19425 9014 22435 9016
rect 19425 9011 19491 9014
rect 22369 9011 22435 9014
rect 29177 9074 29243 9077
rect 31753 9074 31819 9077
rect 29177 9072 31819 9074
rect 29177 9016 29182 9072
rect 29238 9016 31758 9072
rect 31814 9016 31819 9072
rect 29177 9014 31819 9016
rect 29177 9011 29243 9014
rect 31753 9011 31819 9014
rect 29729 8938 29795 8941
rect 34145 8938 34211 8941
rect 29729 8936 34211 8938
rect 29729 8880 29734 8936
rect 29790 8880 34150 8936
rect 34206 8880 34211 8936
rect 29729 8878 34211 8880
rect 29729 8875 29795 8878
rect 34145 8875 34211 8878
rect 4208 8736 4528 8737
rect 4208 8672 4216 8736
rect 4280 8672 4296 8736
rect 4360 8672 4376 8736
rect 4440 8672 4456 8736
rect 4520 8672 4528 8736
rect 4208 8671 4528 8672
rect 34928 8736 35248 8737
rect 34928 8672 34936 8736
rect 35000 8672 35016 8736
rect 35080 8672 35096 8736
rect 35160 8672 35176 8736
rect 35240 8672 35248 8736
rect 34928 8671 35248 8672
rect 30557 8666 30623 8669
rect 34605 8666 34671 8669
rect 30557 8664 34671 8666
rect 30557 8608 30562 8664
rect 30618 8608 34610 8664
rect 34666 8608 34671 8664
rect 30557 8606 34671 8608
rect 30557 8603 30623 8606
rect 34605 8603 34671 8606
rect 20161 8530 20227 8533
rect 20897 8530 20963 8533
rect 20161 8528 20963 8530
rect 20161 8472 20166 8528
rect 20222 8472 20902 8528
rect 20958 8472 20963 8528
rect 20161 8470 20963 8472
rect 20161 8467 20227 8470
rect 20897 8467 20963 8470
rect 16205 8394 16271 8397
rect 17309 8394 17375 8397
rect 16205 8392 17375 8394
rect 16205 8336 16210 8392
rect 16266 8336 17314 8392
rect 17370 8336 17375 8392
rect 16205 8334 17375 8336
rect 16205 8331 16271 8334
rect 17309 8331 17375 8334
rect 16849 8258 16915 8261
rect 18965 8258 19031 8261
rect 16849 8256 19031 8258
rect 16849 8200 16854 8256
rect 16910 8200 18970 8256
rect 19026 8200 19031 8256
rect 16849 8198 19031 8200
rect 16849 8195 16915 8198
rect 18965 8195 19031 8198
rect 19568 8192 19888 8193
rect 19568 8128 19576 8192
rect 19640 8128 19656 8192
rect 19720 8128 19736 8192
rect 19800 8128 19816 8192
rect 19880 8128 19888 8192
rect 19568 8127 19888 8128
rect 8569 8122 8635 8125
rect 11605 8122 11671 8125
rect 8569 8120 11671 8122
rect 8569 8064 8574 8120
rect 8630 8064 11610 8120
rect 11666 8064 11671 8120
rect 8569 8062 11671 8064
rect 8569 8059 8635 8062
rect 11605 8059 11671 8062
rect 11145 7714 11211 7717
rect 17493 7714 17559 7717
rect 11145 7712 17559 7714
rect 11145 7656 11150 7712
rect 11206 7656 17498 7712
rect 17554 7656 17559 7712
rect 11145 7654 17559 7656
rect 11145 7651 11211 7654
rect 17493 7651 17559 7654
rect 4208 7648 4528 7649
rect 4208 7584 4216 7648
rect 4280 7584 4296 7648
rect 4360 7584 4376 7648
rect 4440 7584 4456 7648
rect 4520 7584 4528 7648
rect 4208 7583 4528 7584
rect 34928 7648 35248 7649
rect 34928 7584 34936 7648
rect 35000 7584 35016 7648
rect 35080 7584 35096 7648
rect 35160 7584 35176 7648
rect 35240 7584 35248 7648
rect 34928 7583 35248 7584
rect 11421 7442 11487 7445
rect 12985 7442 13051 7445
rect 11421 7440 13051 7442
rect 11421 7384 11426 7440
rect 11482 7384 12990 7440
rect 13046 7384 13051 7440
rect 11421 7382 13051 7384
rect 11421 7379 11487 7382
rect 12985 7379 13051 7382
rect 21725 7442 21791 7445
rect 24577 7442 24643 7445
rect 21725 7440 24643 7442
rect 21725 7384 21730 7440
rect 21786 7384 24582 7440
rect 24638 7384 24643 7440
rect 21725 7382 24643 7384
rect 21725 7379 21791 7382
rect 24577 7379 24643 7382
rect 38101 7170 38167 7173
rect 39200 7170 40000 7200
rect 38101 7168 40000 7170
rect 38101 7112 38106 7168
rect 38162 7112 40000 7168
rect 38101 7110 40000 7112
rect 38101 7107 38167 7110
rect 19568 7104 19888 7105
rect 19568 7040 19576 7104
rect 19640 7040 19656 7104
rect 19720 7040 19736 7104
rect 19800 7040 19816 7104
rect 19880 7040 19888 7104
rect 39200 7080 40000 7110
rect 19568 7039 19888 7040
rect 0 6898 800 6928
rect 2773 6898 2839 6901
rect 0 6896 2839 6898
rect 0 6840 2778 6896
rect 2834 6840 2839 6896
rect 0 6838 2839 6840
rect 0 6808 800 6838
rect 2773 6835 2839 6838
rect 28993 6762 29059 6765
rect 33961 6762 34027 6765
rect 28993 6760 34027 6762
rect 28993 6704 28998 6760
rect 29054 6704 33966 6760
rect 34022 6704 34027 6760
rect 28993 6702 34027 6704
rect 28993 6699 29059 6702
rect 33961 6699 34027 6702
rect 4208 6560 4528 6561
rect 4208 6496 4216 6560
rect 4280 6496 4296 6560
rect 4360 6496 4376 6560
rect 4440 6496 4456 6560
rect 4520 6496 4528 6560
rect 4208 6495 4528 6496
rect 34928 6560 35248 6561
rect 34928 6496 34936 6560
rect 35000 6496 35016 6560
rect 35080 6496 35096 6560
rect 35160 6496 35176 6560
rect 35240 6496 35248 6560
rect 34928 6495 35248 6496
rect 31937 6354 32003 6357
rect 34789 6354 34855 6357
rect 35617 6354 35683 6357
rect 31937 6352 35683 6354
rect 31937 6296 31942 6352
rect 31998 6296 34794 6352
rect 34850 6296 35622 6352
rect 35678 6296 35683 6352
rect 31937 6294 35683 6296
rect 31937 6291 32003 6294
rect 34789 6291 34855 6294
rect 35617 6291 35683 6294
rect 19568 6016 19888 6017
rect 19568 5952 19576 6016
rect 19640 5952 19656 6016
rect 19720 5952 19736 6016
rect 19800 5952 19816 6016
rect 19880 5952 19888 6016
rect 19568 5951 19888 5952
rect 22093 5674 22159 5677
rect 22921 5674 22987 5677
rect 28625 5674 28691 5677
rect 37917 5674 37983 5677
rect 22093 5672 37983 5674
rect 22093 5616 22098 5672
rect 22154 5616 22926 5672
rect 22982 5616 28630 5672
rect 28686 5616 37922 5672
rect 37978 5616 37983 5672
rect 22093 5614 37983 5616
rect 22093 5611 22159 5614
rect 22921 5611 22987 5614
rect 28625 5611 28691 5614
rect 37917 5611 37983 5614
rect 4208 5472 4528 5473
rect 4208 5408 4216 5472
rect 4280 5408 4296 5472
rect 4360 5408 4376 5472
rect 4440 5408 4456 5472
rect 4520 5408 4528 5472
rect 4208 5407 4528 5408
rect 34928 5472 35248 5473
rect 34928 5408 34936 5472
rect 35000 5408 35016 5472
rect 35080 5408 35096 5472
rect 35160 5408 35176 5472
rect 35240 5408 35248 5472
rect 34928 5407 35248 5408
rect 10961 5130 11027 5133
rect 13721 5130 13787 5133
rect 10961 5128 13787 5130
rect 10961 5072 10966 5128
rect 11022 5072 13726 5128
rect 13782 5072 13787 5128
rect 10961 5070 13787 5072
rect 10961 5067 11027 5070
rect 13721 5067 13787 5070
rect 19568 4928 19888 4929
rect 19568 4864 19576 4928
rect 19640 4864 19656 4928
rect 19720 4864 19736 4928
rect 19800 4864 19816 4928
rect 19880 4864 19888 4928
rect 19568 4863 19888 4864
rect 30925 4722 30991 4725
rect 36537 4722 36603 4725
rect 30925 4720 36603 4722
rect 30925 4664 30930 4720
rect 30986 4664 36542 4720
rect 36598 4664 36603 4720
rect 30925 4662 36603 4664
rect 30925 4659 30991 4662
rect 36537 4659 36603 4662
rect 4208 4384 4528 4385
rect 4208 4320 4216 4384
rect 4280 4320 4296 4384
rect 4360 4320 4376 4384
rect 4440 4320 4456 4384
rect 4520 4320 4528 4384
rect 4208 4319 4528 4320
rect 34928 4384 35248 4385
rect 34928 4320 34936 4384
rect 35000 4320 35016 4384
rect 35080 4320 35096 4384
rect 35160 4320 35176 4384
rect 35240 4320 35248 4384
rect 34928 4319 35248 4320
rect 34789 4178 34855 4181
rect 39200 4178 40000 4208
rect 34789 4176 40000 4178
rect 34789 4120 34794 4176
rect 34850 4120 40000 4176
rect 34789 4118 40000 4120
rect 34789 4115 34855 4118
rect 39200 4088 40000 4118
rect 24526 4042 24532 4044
rect 2270 3982 24532 4042
rect 0 3906 800 3936
rect 2270 3906 2330 3982
rect 24526 3980 24532 3982
rect 24596 3980 24602 4044
rect 0 3846 2330 3906
rect 0 3816 800 3846
rect 19568 3840 19888 3841
rect 19568 3776 19576 3840
rect 19640 3776 19656 3840
rect 19720 3776 19736 3840
rect 19800 3776 19816 3840
rect 19880 3776 19888 3840
rect 19568 3775 19888 3776
rect 565 3498 631 3501
rect 24342 3498 24348 3500
rect 565 3496 24348 3498
rect 565 3440 570 3496
rect 626 3440 24348 3496
rect 565 3438 24348 3440
rect 565 3435 631 3438
rect 24342 3436 24348 3438
rect 24412 3436 24418 3500
rect 4208 3296 4528 3297
rect 4208 3232 4216 3296
rect 4280 3232 4296 3296
rect 4360 3232 4376 3296
rect 4440 3232 4456 3296
rect 4520 3232 4528 3296
rect 4208 3231 4528 3232
rect 34928 3296 35248 3297
rect 34928 3232 34936 3296
rect 35000 3232 35016 3296
rect 35080 3232 35096 3296
rect 35160 3232 35176 3296
rect 35240 3232 35248 3296
rect 34928 3231 35248 3232
rect 10041 3090 10107 3093
rect 16849 3090 16915 3093
rect 10041 3088 16915 3090
rect 10041 3032 10046 3088
rect 10102 3032 16854 3088
rect 16910 3032 16915 3088
rect 10041 3030 16915 3032
rect 10041 3027 10107 3030
rect 16849 3027 16915 3030
rect 19568 2752 19888 2753
rect 19568 2688 19576 2752
rect 19640 2688 19656 2752
rect 19720 2688 19736 2752
rect 19800 2688 19816 2752
rect 19880 2688 19888 2752
rect 19568 2687 19888 2688
rect 4208 2208 4528 2209
rect 4208 2144 4216 2208
rect 4280 2144 4296 2208
rect 4360 2144 4376 2208
rect 4440 2144 4456 2208
rect 4520 2144 4528 2208
rect 4208 2143 4528 2144
rect 34928 2208 35248 2209
rect 34928 2144 34936 2208
rect 35000 2144 35016 2208
rect 35080 2144 35096 2208
rect 35160 2144 35176 2208
rect 35240 2144 35248 2208
rect 34928 2143 35248 2144
rect 38101 1186 38167 1189
rect 39200 1186 40000 1216
rect 38101 1184 40000 1186
rect 38101 1128 38106 1184
rect 38162 1128 40000 1184
rect 38101 1126 40000 1128
rect 38101 1123 38167 1126
rect 39200 1096 40000 1126
<< via3 >>
rect 19576 37564 19640 37568
rect 19576 37508 19580 37564
rect 19580 37508 19636 37564
rect 19636 37508 19640 37564
rect 19576 37504 19640 37508
rect 19656 37564 19720 37568
rect 19656 37508 19660 37564
rect 19660 37508 19716 37564
rect 19716 37508 19720 37564
rect 19656 37504 19720 37508
rect 19736 37564 19800 37568
rect 19736 37508 19740 37564
rect 19740 37508 19796 37564
rect 19796 37508 19800 37564
rect 19736 37504 19800 37508
rect 19816 37564 19880 37568
rect 19816 37508 19820 37564
rect 19820 37508 19876 37564
rect 19876 37508 19880 37564
rect 19816 37504 19880 37508
rect 4216 37020 4280 37024
rect 4216 36964 4220 37020
rect 4220 36964 4276 37020
rect 4276 36964 4280 37020
rect 4216 36960 4280 36964
rect 4296 37020 4360 37024
rect 4296 36964 4300 37020
rect 4300 36964 4356 37020
rect 4356 36964 4360 37020
rect 4296 36960 4360 36964
rect 4376 37020 4440 37024
rect 4376 36964 4380 37020
rect 4380 36964 4436 37020
rect 4436 36964 4440 37020
rect 4376 36960 4440 36964
rect 4456 37020 4520 37024
rect 4456 36964 4460 37020
rect 4460 36964 4516 37020
rect 4516 36964 4520 37020
rect 4456 36960 4520 36964
rect 34936 37020 35000 37024
rect 34936 36964 34940 37020
rect 34940 36964 34996 37020
rect 34996 36964 35000 37020
rect 34936 36960 35000 36964
rect 35016 37020 35080 37024
rect 35016 36964 35020 37020
rect 35020 36964 35076 37020
rect 35076 36964 35080 37020
rect 35016 36960 35080 36964
rect 35096 37020 35160 37024
rect 35096 36964 35100 37020
rect 35100 36964 35156 37020
rect 35156 36964 35160 37020
rect 35096 36960 35160 36964
rect 35176 37020 35240 37024
rect 35176 36964 35180 37020
rect 35180 36964 35236 37020
rect 35236 36964 35240 37020
rect 35176 36960 35240 36964
rect 19576 36476 19640 36480
rect 19576 36420 19580 36476
rect 19580 36420 19636 36476
rect 19636 36420 19640 36476
rect 19576 36416 19640 36420
rect 19656 36476 19720 36480
rect 19656 36420 19660 36476
rect 19660 36420 19716 36476
rect 19716 36420 19720 36476
rect 19656 36416 19720 36420
rect 19736 36476 19800 36480
rect 19736 36420 19740 36476
rect 19740 36420 19796 36476
rect 19796 36420 19800 36476
rect 19736 36416 19800 36420
rect 19816 36476 19880 36480
rect 19816 36420 19820 36476
rect 19820 36420 19876 36476
rect 19876 36420 19880 36476
rect 19816 36416 19880 36420
rect 4216 35932 4280 35936
rect 4216 35876 4220 35932
rect 4220 35876 4276 35932
rect 4276 35876 4280 35932
rect 4216 35872 4280 35876
rect 4296 35932 4360 35936
rect 4296 35876 4300 35932
rect 4300 35876 4356 35932
rect 4356 35876 4360 35932
rect 4296 35872 4360 35876
rect 4376 35932 4440 35936
rect 4376 35876 4380 35932
rect 4380 35876 4436 35932
rect 4436 35876 4440 35932
rect 4376 35872 4440 35876
rect 4456 35932 4520 35936
rect 4456 35876 4460 35932
rect 4460 35876 4516 35932
rect 4516 35876 4520 35932
rect 4456 35872 4520 35876
rect 34936 35932 35000 35936
rect 34936 35876 34940 35932
rect 34940 35876 34996 35932
rect 34996 35876 35000 35932
rect 34936 35872 35000 35876
rect 35016 35932 35080 35936
rect 35016 35876 35020 35932
rect 35020 35876 35076 35932
rect 35076 35876 35080 35932
rect 35016 35872 35080 35876
rect 35096 35932 35160 35936
rect 35096 35876 35100 35932
rect 35100 35876 35156 35932
rect 35156 35876 35160 35932
rect 35096 35872 35160 35876
rect 35176 35932 35240 35936
rect 35176 35876 35180 35932
rect 35180 35876 35236 35932
rect 35236 35876 35240 35932
rect 35176 35872 35240 35876
rect 19576 35388 19640 35392
rect 19576 35332 19580 35388
rect 19580 35332 19636 35388
rect 19636 35332 19640 35388
rect 19576 35328 19640 35332
rect 19656 35388 19720 35392
rect 19656 35332 19660 35388
rect 19660 35332 19716 35388
rect 19716 35332 19720 35388
rect 19656 35328 19720 35332
rect 19736 35388 19800 35392
rect 19736 35332 19740 35388
rect 19740 35332 19796 35388
rect 19796 35332 19800 35388
rect 19736 35328 19800 35332
rect 19816 35388 19880 35392
rect 19816 35332 19820 35388
rect 19820 35332 19876 35388
rect 19876 35332 19880 35388
rect 19816 35328 19880 35332
rect 4216 34844 4280 34848
rect 4216 34788 4220 34844
rect 4220 34788 4276 34844
rect 4276 34788 4280 34844
rect 4216 34784 4280 34788
rect 4296 34844 4360 34848
rect 4296 34788 4300 34844
rect 4300 34788 4356 34844
rect 4356 34788 4360 34844
rect 4296 34784 4360 34788
rect 4376 34844 4440 34848
rect 4376 34788 4380 34844
rect 4380 34788 4436 34844
rect 4436 34788 4440 34844
rect 4376 34784 4440 34788
rect 4456 34844 4520 34848
rect 4456 34788 4460 34844
rect 4460 34788 4516 34844
rect 4516 34788 4520 34844
rect 4456 34784 4520 34788
rect 34936 34844 35000 34848
rect 34936 34788 34940 34844
rect 34940 34788 34996 34844
rect 34996 34788 35000 34844
rect 34936 34784 35000 34788
rect 35016 34844 35080 34848
rect 35016 34788 35020 34844
rect 35020 34788 35076 34844
rect 35076 34788 35080 34844
rect 35016 34784 35080 34788
rect 35096 34844 35160 34848
rect 35096 34788 35100 34844
rect 35100 34788 35156 34844
rect 35156 34788 35160 34844
rect 35096 34784 35160 34788
rect 35176 34844 35240 34848
rect 35176 34788 35180 34844
rect 35180 34788 35236 34844
rect 35236 34788 35240 34844
rect 35176 34784 35240 34788
rect 19576 34300 19640 34304
rect 19576 34244 19580 34300
rect 19580 34244 19636 34300
rect 19636 34244 19640 34300
rect 19576 34240 19640 34244
rect 19656 34300 19720 34304
rect 19656 34244 19660 34300
rect 19660 34244 19716 34300
rect 19716 34244 19720 34300
rect 19656 34240 19720 34244
rect 19736 34300 19800 34304
rect 19736 34244 19740 34300
rect 19740 34244 19796 34300
rect 19796 34244 19800 34300
rect 19736 34240 19800 34244
rect 19816 34300 19880 34304
rect 19816 34244 19820 34300
rect 19820 34244 19876 34300
rect 19876 34244 19880 34300
rect 19816 34240 19880 34244
rect 4216 33756 4280 33760
rect 4216 33700 4220 33756
rect 4220 33700 4276 33756
rect 4276 33700 4280 33756
rect 4216 33696 4280 33700
rect 4296 33756 4360 33760
rect 4296 33700 4300 33756
rect 4300 33700 4356 33756
rect 4356 33700 4360 33756
rect 4296 33696 4360 33700
rect 4376 33756 4440 33760
rect 4376 33700 4380 33756
rect 4380 33700 4436 33756
rect 4436 33700 4440 33756
rect 4376 33696 4440 33700
rect 4456 33756 4520 33760
rect 4456 33700 4460 33756
rect 4460 33700 4516 33756
rect 4516 33700 4520 33756
rect 4456 33696 4520 33700
rect 34936 33756 35000 33760
rect 34936 33700 34940 33756
rect 34940 33700 34996 33756
rect 34996 33700 35000 33756
rect 34936 33696 35000 33700
rect 35016 33756 35080 33760
rect 35016 33700 35020 33756
rect 35020 33700 35076 33756
rect 35076 33700 35080 33756
rect 35016 33696 35080 33700
rect 35096 33756 35160 33760
rect 35096 33700 35100 33756
rect 35100 33700 35156 33756
rect 35156 33700 35160 33756
rect 35096 33696 35160 33700
rect 35176 33756 35240 33760
rect 35176 33700 35180 33756
rect 35180 33700 35236 33756
rect 35236 33700 35240 33756
rect 35176 33696 35240 33700
rect 19576 33212 19640 33216
rect 19576 33156 19580 33212
rect 19580 33156 19636 33212
rect 19636 33156 19640 33212
rect 19576 33152 19640 33156
rect 19656 33212 19720 33216
rect 19656 33156 19660 33212
rect 19660 33156 19716 33212
rect 19716 33156 19720 33212
rect 19656 33152 19720 33156
rect 19736 33212 19800 33216
rect 19736 33156 19740 33212
rect 19740 33156 19796 33212
rect 19796 33156 19800 33212
rect 19736 33152 19800 33156
rect 19816 33212 19880 33216
rect 19816 33156 19820 33212
rect 19820 33156 19876 33212
rect 19876 33156 19880 33212
rect 19816 33152 19880 33156
rect 4216 32668 4280 32672
rect 4216 32612 4220 32668
rect 4220 32612 4276 32668
rect 4276 32612 4280 32668
rect 4216 32608 4280 32612
rect 4296 32668 4360 32672
rect 4296 32612 4300 32668
rect 4300 32612 4356 32668
rect 4356 32612 4360 32668
rect 4296 32608 4360 32612
rect 4376 32668 4440 32672
rect 4376 32612 4380 32668
rect 4380 32612 4436 32668
rect 4436 32612 4440 32668
rect 4376 32608 4440 32612
rect 4456 32668 4520 32672
rect 4456 32612 4460 32668
rect 4460 32612 4516 32668
rect 4516 32612 4520 32668
rect 4456 32608 4520 32612
rect 34936 32668 35000 32672
rect 34936 32612 34940 32668
rect 34940 32612 34996 32668
rect 34996 32612 35000 32668
rect 34936 32608 35000 32612
rect 35016 32668 35080 32672
rect 35016 32612 35020 32668
rect 35020 32612 35076 32668
rect 35076 32612 35080 32668
rect 35016 32608 35080 32612
rect 35096 32668 35160 32672
rect 35096 32612 35100 32668
rect 35100 32612 35156 32668
rect 35156 32612 35160 32668
rect 35096 32608 35160 32612
rect 35176 32668 35240 32672
rect 35176 32612 35180 32668
rect 35180 32612 35236 32668
rect 35236 32612 35240 32668
rect 35176 32608 35240 32612
rect 19576 32124 19640 32128
rect 19576 32068 19580 32124
rect 19580 32068 19636 32124
rect 19636 32068 19640 32124
rect 19576 32064 19640 32068
rect 19656 32124 19720 32128
rect 19656 32068 19660 32124
rect 19660 32068 19716 32124
rect 19716 32068 19720 32124
rect 19656 32064 19720 32068
rect 19736 32124 19800 32128
rect 19736 32068 19740 32124
rect 19740 32068 19796 32124
rect 19796 32068 19800 32124
rect 19736 32064 19800 32068
rect 19816 32124 19880 32128
rect 19816 32068 19820 32124
rect 19820 32068 19876 32124
rect 19876 32068 19880 32124
rect 19816 32064 19880 32068
rect 4216 31580 4280 31584
rect 4216 31524 4220 31580
rect 4220 31524 4276 31580
rect 4276 31524 4280 31580
rect 4216 31520 4280 31524
rect 4296 31580 4360 31584
rect 4296 31524 4300 31580
rect 4300 31524 4356 31580
rect 4356 31524 4360 31580
rect 4296 31520 4360 31524
rect 4376 31580 4440 31584
rect 4376 31524 4380 31580
rect 4380 31524 4436 31580
rect 4436 31524 4440 31580
rect 4376 31520 4440 31524
rect 4456 31580 4520 31584
rect 4456 31524 4460 31580
rect 4460 31524 4516 31580
rect 4516 31524 4520 31580
rect 4456 31520 4520 31524
rect 34936 31580 35000 31584
rect 34936 31524 34940 31580
rect 34940 31524 34996 31580
rect 34996 31524 35000 31580
rect 34936 31520 35000 31524
rect 35016 31580 35080 31584
rect 35016 31524 35020 31580
rect 35020 31524 35076 31580
rect 35076 31524 35080 31580
rect 35016 31520 35080 31524
rect 35096 31580 35160 31584
rect 35096 31524 35100 31580
rect 35100 31524 35156 31580
rect 35156 31524 35160 31580
rect 35096 31520 35160 31524
rect 35176 31580 35240 31584
rect 35176 31524 35180 31580
rect 35180 31524 35236 31580
rect 35236 31524 35240 31580
rect 35176 31520 35240 31524
rect 19576 31036 19640 31040
rect 19576 30980 19580 31036
rect 19580 30980 19636 31036
rect 19636 30980 19640 31036
rect 19576 30976 19640 30980
rect 19656 31036 19720 31040
rect 19656 30980 19660 31036
rect 19660 30980 19716 31036
rect 19716 30980 19720 31036
rect 19656 30976 19720 30980
rect 19736 31036 19800 31040
rect 19736 30980 19740 31036
rect 19740 30980 19796 31036
rect 19796 30980 19800 31036
rect 19736 30976 19800 30980
rect 19816 31036 19880 31040
rect 19816 30980 19820 31036
rect 19820 30980 19876 31036
rect 19876 30980 19880 31036
rect 19816 30976 19880 30980
rect 4216 30492 4280 30496
rect 4216 30436 4220 30492
rect 4220 30436 4276 30492
rect 4276 30436 4280 30492
rect 4216 30432 4280 30436
rect 4296 30492 4360 30496
rect 4296 30436 4300 30492
rect 4300 30436 4356 30492
rect 4356 30436 4360 30492
rect 4296 30432 4360 30436
rect 4376 30492 4440 30496
rect 4376 30436 4380 30492
rect 4380 30436 4436 30492
rect 4436 30436 4440 30492
rect 4376 30432 4440 30436
rect 4456 30492 4520 30496
rect 4456 30436 4460 30492
rect 4460 30436 4516 30492
rect 4516 30436 4520 30492
rect 4456 30432 4520 30436
rect 34936 30492 35000 30496
rect 34936 30436 34940 30492
rect 34940 30436 34996 30492
rect 34996 30436 35000 30492
rect 34936 30432 35000 30436
rect 35016 30492 35080 30496
rect 35016 30436 35020 30492
rect 35020 30436 35076 30492
rect 35076 30436 35080 30492
rect 35016 30432 35080 30436
rect 35096 30492 35160 30496
rect 35096 30436 35100 30492
rect 35100 30436 35156 30492
rect 35156 30436 35160 30492
rect 35096 30432 35160 30436
rect 35176 30492 35240 30496
rect 35176 30436 35180 30492
rect 35180 30436 35236 30492
rect 35236 30436 35240 30492
rect 35176 30432 35240 30436
rect 24532 30424 24596 30428
rect 24532 30368 24546 30424
rect 24546 30368 24596 30424
rect 24532 30364 24596 30368
rect 19576 29948 19640 29952
rect 19576 29892 19580 29948
rect 19580 29892 19636 29948
rect 19636 29892 19640 29948
rect 19576 29888 19640 29892
rect 19656 29948 19720 29952
rect 19656 29892 19660 29948
rect 19660 29892 19716 29948
rect 19716 29892 19720 29948
rect 19656 29888 19720 29892
rect 19736 29948 19800 29952
rect 19736 29892 19740 29948
rect 19740 29892 19796 29948
rect 19796 29892 19800 29948
rect 19736 29888 19800 29892
rect 19816 29948 19880 29952
rect 19816 29892 19820 29948
rect 19820 29892 19876 29948
rect 19876 29892 19880 29948
rect 19816 29888 19880 29892
rect 4216 29404 4280 29408
rect 4216 29348 4220 29404
rect 4220 29348 4276 29404
rect 4276 29348 4280 29404
rect 4216 29344 4280 29348
rect 4296 29404 4360 29408
rect 4296 29348 4300 29404
rect 4300 29348 4356 29404
rect 4356 29348 4360 29404
rect 4296 29344 4360 29348
rect 4376 29404 4440 29408
rect 4376 29348 4380 29404
rect 4380 29348 4436 29404
rect 4436 29348 4440 29404
rect 4376 29344 4440 29348
rect 4456 29404 4520 29408
rect 4456 29348 4460 29404
rect 4460 29348 4516 29404
rect 4516 29348 4520 29404
rect 4456 29344 4520 29348
rect 34936 29404 35000 29408
rect 34936 29348 34940 29404
rect 34940 29348 34996 29404
rect 34996 29348 35000 29404
rect 34936 29344 35000 29348
rect 35016 29404 35080 29408
rect 35016 29348 35020 29404
rect 35020 29348 35076 29404
rect 35076 29348 35080 29404
rect 35016 29344 35080 29348
rect 35096 29404 35160 29408
rect 35096 29348 35100 29404
rect 35100 29348 35156 29404
rect 35156 29348 35160 29404
rect 35096 29344 35160 29348
rect 35176 29404 35240 29408
rect 35176 29348 35180 29404
rect 35180 29348 35236 29404
rect 35236 29348 35240 29404
rect 35176 29344 35240 29348
rect 19576 28860 19640 28864
rect 19576 28804 19580 28860
rect 19580 28804 19636 28860
rect 19636 28804 19640 28860
rect 19576 28800 19640 28804
rect 19656 28860 19720 28864
rect 19656 28804 19660 28860
rect 19660 28804 19716 28860
rect 19716 28804 19720 28860
rect 19656 28800 19720 28804
rect 19736 28860 19800 28864
rect 19736 28804 19740 28860
rect 19740 28804 19796 28860
rect 19796 28804 19800 28860
rect 19736 28800 19800 28804
rect 19816 28860 19880 28864
rect 19816 28804 19820 28860
rect 19820 28804 19876 28860
rect 19876 28804 19880 28860
rect 19816 28800 19880 28804
rect 4216 28316 4280 28320
rect 4216 28260 4220 28316
rect 4220 28260 4276 28316
rect 4276 28260 4280 28316
rect 4216 28256 4280 28260
rect 4296 28316 4360 28320
rect 4296 28260 4300 28316
rect 4300 28260 4356 28316
rect 4356 28260 4360 28316
rect 4296 28256 4360 28260
rect 4376 28316 4440 28320
rect 4376 28260 4380 28316
rect 4380 28260 4436 28316
rect 4436 28260 4440 28316
rect 4376 28256 4440 28260
rect 4456 28316 4520 28320
rect 4456 28260 4460 28316
rect 4460 28260 4516 28316
rect 4516 28260 4520 28316
rect 4456 28256 4520 28260
rect 34936 28316 35000 28320
rect 34936 28260 34940 28316
rect 34940 28260 34996 28316
rect 34996 28260 35000 28316
rect 34936 28256 35000 28260
rect 35016 28316 35080 28320
rect 35016 28260 35020 28316
rect 35020 28260 35076 28316
rect 35076 28260 35080 28316
rect 35016 28256 35080 28260
rect 35096 28316 35160 28320
rect 35096 28260 35100 28316
rect 35100 28260 35156 28316
rect 35156 28260 35160 28316
rect 35096 28256 35160 28260
rect 35176 28316 35240 28320
rect 35176 28260 35180 28316
rect 35180 28260 35236 28316
rect 35236 28260 35240 28316
rect 35176 28256 35240 28260
rect 19576 27772 19640 27776
rect 19576 27716 19580 27772
rect 19580 27716 19636 27772
rect 19636 27716 19640 27772
rect 19576 27712 19640 27716
rect 19656 27772 19720 27776
rect 19656 27716 19660 27772
rect 19660 27716 19716 27772
rect 19716 27716 19720 27772
rect 19656 27712 19720 27716
rect 19736 27772 19800 27776
rect 19736 27716 19740 27772
rect 19740 27716 19796 27772
rect 19796 27716 19800 27772
rect 19736 27712 19800 27716
rect 19816 27772 19880 27776
rect 19816 27716 19820 27772
rect 19820 27716 19876 27772
rect 19876 27716 19880 27772
rect 19816 27712 19880 27716
rect 4216 27228 4280 27232
rect 4216 27172 4220 27228
rect 4220 27172 4276 27228
rect 4276 27172 4280 27228
rect 4216 27168 4280 27172
rect 4296 27228 4360 27232
rect 4296 27172 4300 27228
rect 4300 27172 4356 27228
rect 4356 27172 4360 27228
rect 4296 27168 4360 27172
rect 4376 27228 4440 27232
rect 4376 27172 4380 27228
rect 4380 27172 4436 27228
rect 4436 27172 4440 27228
rect 4376 27168 4440 27172
rect 4456 27228 4520 27232
rect 4456 27172 4460 27228
rect 4460 27172 4516 27228
rect 4516 27172 4520 27228
rect 4456 27168 4520 27172
rect 34936 27228 35000 27232
rect 34936 27172 34940 27228
rect 34940 27172 34996 27228
rect 34996 27172 35000 27228
rect 34936 27168 35000 27172
rect 35016 27228 35080 27232
rect 35016 27172 35020 27228
rect 35020 27172 35076 27228
rect 35076 27172 35080 27228
rect 35016 27168 35080 27172
rect 35096 27228 35160 27232
rect 35096 27172 35100 27228
rect 35100 27172 35156 27228
rect 35156 27172 35160 27228
rect 35096 27168 35160 27172
rect 35176 27228 35240 27232
rect 35176 27172 35180 27228
rect 35180 27172 35236 27228
rect 35236 27172 35240 27228
rect 35176 27168 35240 27172
rect 19576 26684 19640 26688
rect 19576 26628 19580 26684
rect 19580 26628 19636 26684
rect 19636 26628 19640 26684
rect 19576 26624 19640 26628
rect 19656 26684 19720 26688
rect 19656 26628 19660 26684
rect 19660 26628 19716 26684
rect 19716 26628 19720 26684
rect 19656 26624 19720 26628
rect 19736 26684 19800 26688
rect 19736 26628 19740 26684
rect 19740 26628 19796 26684
rect 19796 26628 19800 26684
rect 19736 26624 19800 26628
rect 19816 26684 19880 26688
rect 19816 26628 19820 26684
rect 19820 26628 19876 26684
rect 19876 26628 19880 26684
rect 19816 26624 19880 26628
rect 4216 26140 4280 26144
rect 4216 26084 4220 26140
rect 4220 26084 4276 26140
rect 4276 26084 4280 26140
rect 4216 26080 4280 26084
rect 4296 26140 4360 26144
rect 4296 26084 4300 26140
rect 4300 26084 4356 26140
rect 4356 26084 4360 26140
rect 4296 26080 4360 26084
rect 4376 26140 4440 26144
rect 4376 26084 4380 26140
rect 4380 26084 4436 26140
rect 4436 26084 4440 26140
rect 4376 26080 4440 26084
rect 4456 26140 4520 26144
rect 4456 26084 4460 26140
rect 4460 26084 4516 26140
rect 4516 26084 4520 26140
rect 4456 26080 4520 26084
rect 34936 26140 35000 26144
rect 34936 26084 34940 26140
rect 34940 26084 34996 26140
rect 34996 26084 35000 26140
rect 34936 26080 35000 26084
rect 35016 26140 35080 26144
rect 35016 26084 35020 26140
rect 35020 26084 35076 26140
rect 35076 26084 35080 26140
rect 35016 26080 35080 26084
rect 35096 26140 35160 26144
rect 35096 26084 35100 26140
rect 35100 26084 35156 26140
rect 35156 26084 35160 26140
rect 35096 26080 35160 26084
rect 35176 26140 35240 26144
rect 35176 26084 35180 26140
rect 35180 26084 35236 26140
rect 35236 26084 35240 26140
rect 35176 26080 35240 26084
rect 19576 25596 19640 25600
rect 19576 25540 19580 25596
rect 19580 25540 19636 25596
rect 19636 25540 19640 25596
rect 19576 25536 19640 25540
rect 19656 25596 19720 25600
rect 19656 25540 19660 25596
rect 19660 25540 19716 25596
rect 19716 25540 19720 25596
rect 19656 25536 19720 25540
rect 19736 25596 19800 25600
rect 19736 25540 19740 25596
rect 19740 25540 19796 25596
rect 19796 25540 19800 25596
rect 19736 25536 19800 25540
rect 19816 25596 19880 25600
rect 19816 25540 19820 25596
rect 19820 25540 19876 25596
rect 19876 25540 19880 25596
rect 19816 25536 19880 25540
rect 4216 25052 4280 25056
rect 4216 24996 4220 25052
rect 4220 24996 4276 25052
rect 4276 24996 4280 25052
rect 4216 24992 4280 24996
rect 4296 25052 4360 25056
rect 4296 24996 4300 25052
rect 4300 24996 4356 25052
rect 4356 24996 4360 25052
rect 4296 24992 4360 24996
rect 4376 25052 4440 25056
rect 4376 24996 4380 25052
rect 4380 24996 4436 25052
rect 4436 24996 4440 25052
rect 4376 24992 4440 24996
rect 4456 25052 4520 25056
rect 4456 24996 4460 25052
rect 4460 24996 4516 25052
rect 4516 24996 4520 25052
rect 4456 24992 4520 24996
rect 34936 25052 35000 25056
rect 34936 24996 34940 25052
rect 34940 24996 34996 25052
rect 34996 24996 35000 25052
rect 34936 24992 35000 24996
rect 35016 25052 35080 25056
rect 35016 24996 35020 25052
rect 35020 24996 35076 25052
rect 35076 24996 35080 25052
rect 35016 24992 35080 24996
rect 35096 25052 35160 25056
rect 35096 24996 35100 25052
rect 35100 24996 35156 25052
rect 35156 24996 35160 25052
rect 35096 24992 35160 24996
rect 35176 25052 35240 25056
rect 35176 24996 35180 25052
rect 35180 24996 35236 25052
rect 35236 24996 35240 25052
rect 35176 24992 35240 24996
rect 24348 24984 24412 24988
rect 24348 24928 24398 24984
rect 24398 24928 24412 24984
rect 24348 24924 24412 24928
rect 19576 24508 19640 24512
rect 19576 24452 19580 24508
rect 19580 24452 19636 24508
rect 19636 24452 19640 24508
rect 19576 24448 19640 24452
rect 19656 24508 19720 24512
rect 19656 24452 19660 24508
rect 19660 24452 19716 24508
rect 19716 24452 19720 24508
rect 19656 24448 19720 24452
rect 19736 24508 19800 24512
rect 19736 24452 19740 24508
rect 19740 24452 19796 24508
rect 19796 24452 19800 24508
rect 19736 24448 19800 24452
rect 19816 24508 19880 24512
rect 19816 24452 19820 24508
rect 19820 24452 19876 24508
rect 19876 24452 19880 24508
rect 19816 24448 19880 24452
rect 4216 23964 4280 23968
rect 4216 23908 4220 23964
rect 4220 23908 4276 23964
rect 4276 23908 4280 23964
rect 4216 23904 4280 23908
rect 4296 23964 4360 23968
rect 4296 23908 4300 23964
rect 4300 23908 4356 23964
rect 4356 23908 4360 23964
rect 4296 23904 4360 23908
rect 4376 23964 4440 23968
rect 4376 23908 4380 23964
rect 4380 23908 4436 23964
rect 4436 23908 4440 23964
rect 4376 23904 4440 23908
rect 4456 23964 4520 23968
rect 4456 23908 4460 23964
rect 4460 23908 4516 23964
rect 4516 23908 4520 23964
rect 4456 23904 4520 23908
rect 34936 23964 35000 23968
rect 34936 23908 34940 23964
rect 34940 23908 34996 23964
rect 34996 23908 35000 23964
rect 34936 23904 35000 23908
rect 35016 23964 35080 23968
rect 35016 23908 35020 23964
rect 35020 23908 35076 23964
rect 35076 23908 35080 23964
rect 35016 23904 35080 23908
rect 35096 23964 35160 23968
rect 35096 23908 35100 23964
rect 35100 23908 35156 23964
rect 35156 23908 35160 23964
rect 35096 23904 35160 23908
rect 35176 23964 35240 23968
rect 35176 23908 35180 23964
rect 35180 23908 35236 23964
rect 35236 23908 35240 23964
rect 35176 23904 35240 23908
rect 19576 23420 19640 23424
rect 19576 23364 19580 23420
rect 19580 23364 19636 23420
rect 19636 23364 19640 23420
rect 19576 23360 19640 23364
rect 19656 23420 19720 23424
rect 19656 23364 19660 23420
rect 19660 23364 19716 23420
rect 19716 23364 19720 23420
rect 19656 23360 19720 23364
rect 19736 23420 19800 23424
rect 19736 23364 19740 23420
rect 19740 23364 19796 23420
rect 19796 23364 19800 23420
rect 19736 23360 19800 23364
rect 19816 23420 19880 23424
rect 19816 23364 19820 23420
rect 19820 23364 19876 23420
rect 19876 23364 19880 23420
rect 19816 23360 19880 23364
rect 4216 22876 4280 22880
rect 4216 22820 4220 22876
rect 4220 22820 4276 22876
rect 4276 22820 4280 22876
rect 4216 22816 4280 22820
rect 4296 22876 4360 22880
rect 4296 22820 4300 22876
rect 4300 22820 4356 22876
rect 4356 22820 4360 22876
rect 4296 22816 4360 22820
rect 4376 22876 4440 22880
rect 4376 22820 4380 22876
rect 4380 22820 4436 22876
rect 4436 22820 4440 22876
rect 4376 22816 4440 22820
rect 4456 22876 4520 22880
rect 4456 22820 4460 22876
rect 4460 22820 4516 22876
rect 4516 22820 4520 22876
rect 4456 22816 4520 22820
rect 34936 22876 35000 22880
rect 34936 22820 34940 22876
rect 34940 22820 34996 22876
rect 34996 22820 35000 22876
rect 34936 22816 35000 22820
rect 35016 22876 35080 22880
rect 35016 22820 35020 22876
rect 35020 22820 35076 22876
rect 35076 22820 35080 22876
rect 35016 22816 35080 22820
rect 35096 22876 35160 22880
rect 35096 22820 35100 22876
rect 35100 22820 35156 22876
rect 35156 22820 35160 22876
rect 35096 22816 35160 22820
rect 35176 22876 35240 22880
rect 35176 22820 35180 22876
rect 35180 22820 35236 22876
rect 35236 22820 35240 22876
rect 35176 22816 35240 22820
rect 19576 22332 19640 22336
rect 19576 22276 19580 22332
rect 19580 22276 19636 22332
rect 19636 22276 19640 22332
rect 19576 22272 19640 22276
rect 19656 22332 19720 22336
rect 19656 22276 19660 22332
rect 19660 22276 19716 22332
rect 19716 22276 19720 22332
rect 19656 22272 19720 22276
rect 19736 22332 19800 22336
rect 19736 22276 19740 22332
rect 19740 22276 19796 22332
rect 19796 22276 19800 22332
rect 19736 22272 19800 22276
rect 19816 22332 19880 22336
rect 19816 22276 19820 22332
rect 19820 22276 19876 22332
rect 19876 22276 19880 22332
rect 19816 22272 19880 22276
rect 4216 21788 4280 21792
rect 4216 21732 4220 21788
rect 4220 21732 4276 21788
rect 4276 21732 4280 21788
rect 4216 21728 4280 21732
rect 4296 21788 4360 21792
rect 4296 21732 4300 21788
rect 4300 21732 4356 21788
rect 4356 21732 4360 21788
rect 4296 21728 4360 21732
rect 4376 21788 4440 21792
rect 4376 21732 4380 21788
rect 4380 21732 4436 21788
rect 4436 21732 4440 21788
rect 4376 21728 4440 21732
rect 4456 21788 4520 21792
rect 4456 21732 4460 21788
rect 4460 21732 4516 21788
rect 4516 21732 4520 21788
rect 4456 21728 4520 21732
rect 34936 21788 35000 21792
rect 34936 21732 34940 21788
rect 34940 21732 34996 21788
rect 34996 21732 35000 21788
rect 34936 21728 35000 21732
rect 35016 21788 35080 21792
rect 35016 21732 35020 21788
rect 35020 21732 35076 21788
rect 35076 21732 35080 21788
rect 35016 21728 35080 21732
rect 35096 21788 35160 21792
rect 35096 21732 35100 21788
rect 35100 21732 35156 21788
rect 35156 21732 35160 21788
rect 35096 21728 35160 21732
rect 35176 21788 35240 21792
rect 35176 21732 35180 21788
rect 35180 21732 35236 21788
rect 35236 21732 35240 21788
rect 35176 21728 35240 21732
rect 19576 21244 19640 21248
rect 19576 21188 19580 21244
rect 19580 21188 19636 21244
rect 19636 21188 19640 21244
rect 19576 21184 19640 21188
rect 19656 21244 19720 21248
rect 19656 21188 19660 21244
rect 19660 21188 19716 21244
rect 19716 21188 19720 21244
rect 19656 21184 19720 21188
rect 19736 21244 19800 21248
rect 19736 21188 19740 21244
rect 19740 21188 19796 21244
rect 19796 21188 19800 21244
rect 19736 21184 19800 21188
rect 19816 21244 19880 21248
rect 19816 21188 19820 21244
rect 19820 21188 19876 21244
rect 19876 21188 19880 21244
rect 19816 21184 19880 21188
rect 4216 20700 4280 20704
rect 4216 20644 4220 20700
rect 4220 20644 4276 20700
rect 4276 20644 4280 20700
rect 4216 20640 4280 20644
rect 4296 20700 4360 20704
rect 4296 20644 4300 20700
rect 4300 20644 4356 20700
rect 4356 20644 4360 20700
rect 4296 20640 4360 20644
rect 4376 20700 4440 20704
rect 4376 20644 4380 20700
rect 4380 20644 4436 20700
rect 4436 20644 4440 20700
rect 4376 20640 4440 20644
rect 4456 20700 4520 20704
rect 4456 20644 4460 20700
rect 4460 20644 4516 20700
rect 4516 20644 4520 20700
rect 4456 20640 4520 20644
rect 34936 20700 35000 20704
rect 34936 20644 34940 20700
rect 34940 20644 34996 20700
rect 34996 20644 35000 20700
rect 34936 20640 35000 20644
rect 35016 20700 35080 20704
rect 35016 20644 35020 20700
rect 35020 20644 35076 20700
rect 35076 20644 35080 20700
rect 35016 20640 35080 20644
rect 35096 20700 35160 20704
rect 35096 20644 35100 20700
rect 35100 20644 35156 20700
rect 35156 20644 35160 20700
rect 35096 20640 35160 20644
rect 35176 20700 35240 20704
rect 35176 20644 35180 20700
rect 35180 20644 35236 20700
rect 35236 20644 35240 20700
rect 35176 20640 35240 20644
rect 19576 20156 19640 20160
rect 19576 20100 19580 20156
rect 19580 20100 19636 20156
rect 19636 20100 19640 20156
rect 19576 20096 19640 20100
rect 19656 20156 19720 20160
rect 19656 20100 19660 20156
rect 19660 20100 19716 20156
rect 19716 20100 19720 20156
rect 19656 20096 19720 20100
rect 19736 20156 19800 20160
rect 19736 20100 19740 20156
rect 19740 20100 19796 20156
rect 19796 20100 19800 20156
rect 19736 20096 19800 20100
rect 19816 20156 19880 20160
rect 19816 20100 19820 20156
rect 19820 20100 19876 20156
rect 19876 20100 19880 20156
rect 19816 20096 19880 20100
rect 4216 19612 4280 19616
rect 4216 19556 4220 19612
rect 4220 19556 4276 19612
rect 4276 19556 4280 19612
rect 4216 19552 4280 19556
rect 4296 19612 4360 19616
rect 4296 19556 4300 19612
rect 4300 19556 4356 19612
rect 4356 19556 4360 19612
rect 4296 19552 4360 19556
rect 4376 19612 4440 19616
rect 4376 19556 4380 19612
rect 4380 19556 4436 19612
rect 4436 19556 4440 19612
rect 4376 19552 4440 19556
rect 4456 19612 4520 19616
rect 4456 19556 4460 19612
rect 4460 19556 4516 19612
rect 4516 19556 4520 19612
rect 4456 19552 4520 19556
rect 34936 19612 35000 19616
rect 34936 19556 34940 19612
rect 34940 19556 34996 19612
rect 34996 19556 35000 19612
rect 34936 19552 35000 19556
rect 35016 19612 35080 19616
rect 35016 19556 35020 19612
rect 35020 19556 35076 19612
rect 35076 19556 35080 19612
rect 35016 19552 35080 19556
rect 35096 19612 35160 19616
rect 35096 19556 35100 19612
rect 35100 19556 35156 19612
rect 35156 19556 35160 19612
rect 35096 19552 35160 19556
rect 35176 19612 35240 19616
rect 35176 19556 35180 19612
rect 35180 19556 35236 19612
rect 35236 19556 35240 19612
rect 35176 19552 35240 19556
rect 19576 19068 19640 19072
rect 19576 19012 19580 19068
rect 19580 19012 19636 19068
rect 19636 19012 19640 19068
rect 19576 19008 19640 19012
rect 19656 19068 19720 19072
rect 19656 19012 19660 19068
rect 19660 19012 19716 19068
rect 19716 19012 19720 19068
rect 19656 19008 19720 19012
rect 19736 19068 19800 19072
rect 19736 19012 19740 19068
rect 19740 19012 19796 19068
rect 19796 19012 19800 19068
rect 19736 19008 19800 19012
rect 19816 19068 19880 19072
rect 19816 19012 19820 19068
rect 19820 19012 19876 19068
rect 19876 19012 19880 19068
rect 19816 19008 19880 19012
rect 4216 18524 4280 18528
rect 4216 18468 4220 18524
rect 4220 18468 4276 18524
rect 4276 18468 4280 18524
rect 4216 18464 4280 18468
rect 4296 18524 4360 18528
rect 4296 18468 4300 18524
rect 4300 18468 4356 18524
rect 4356 18468 4360 18524
rect 4296 18464 4360 18468
rect 4376 18524 4440 18528
rect 4376 18468 4380 18524
rect 4380 18468 4436 18524
rect 4436 18468 4440 18524
rect 4376 18464 4440 18468
rect 4456 18524 4520 18528
rect 4456 18468 4460 18524
rect 4460 18468 4516 18524
rect 4516 18468 4520 18524
rect 4456 18464 4520 18468
rect 34936 18524 35000 18528
rect 34936 18468 34940 18524
rect 34940 18468 34996 18524
rect 34996 18468 35000 18524
rect 34936 18464 35000 18468
rect 35016 18524 35080 18528
rect 35016 18468 35020 18524
rect 35020 18468 35076 18524
rect 35076 18468 35080 18524
rect 35016 18464 35080 18468
rect 35096 18524 35160 18528
rect 35096 18468 35100 18524
rect 35100 18468 35156 18524
rect 35156 18468 35160 18524
rect 35096 18464 35160 18468
rect 35176 18524 35240 18528
rect 35176 18468 35180 18524
rect 35180 18468 35236 18524
rect 35236 18468 35240 18524
rect 35176 18464 35240 18468
rect 19576 17980 19640 17984
rect 19576 17924 19580 17980
rect 19580 17924 19636 17980
rect 19636 17924 19640 17980
rect 19576 17920 19640 17924
rect 19656 17980 19720 17984
rect 19656 17924 19660 17980
rect 19660 17924 19716 17980
rect 19716 17924 19720 17980
rect 19656 17920 19720 17924
rect 19736 17980 19800 17984
rect 19736 17924 19740 17980
rect 19740 17924 19796 17980
rect 19796 17924 19800 17980
rect 19736 17920 19800 17924
rect 19816 17980 19880 17984
rect 19816 17924 19820 17980
rect 19820 17924 19876 17980
rect 19876 17924 19880 17980
rect 19816 17920 19880 17924
rect 4216 17436 4280 17440
rect 4216 17380 4220 17436
rect 4220 17380 4276 17436
rect 4276 17380 4280 17436
rect 4216 17376 4280 17380
rect 4296 17436 4360 17440
rect 4296 17380 4300 17436
rect 4300 17380 4356 17436
rect 4356 17380 4360 17436
rect 4296 17376 4360 17380
rect 4376 17436 4440 17440
rect 4376 17380 4380 17436
rect 4380 17380 4436 17436
rect 4436 17380 4440 17436
rect 4376 17376 4440 17380
rect 4456 17436 4520 17440
rect 4456 17380 4460 17436
rect 4460 17380 4516 17436
rect 4516 17380 4520 17436
rect 4456 17376 4520 17380
rect 34936 17436 35000 17440
rect 34936 17380 34940 17436
rect 34940 17380 34996 17436
rect 34996 17380 35000 17436
rect 34936 17376 35000 17380
rect 35016 17436 35080 17440
rect 35016 17380 35020 17436
rect 35020 17380 35076 17436
rect 35076 17380 35080 17436
rect 35016 17376 35080 17380
rect 35096 17436 35160 17440
rect 35096 17380 35100 17436
rect 35100 17380 35156 17436
rect 35156 17380 35160 17436
rect 35096 17376 35160 17380
rect 35176 17436 35240 17440
rect 35176 17380 35180 17436
rect 35180 17380 35236 17436
rect 35236 17380 35240 17436
rect 35176 17376 35240 17380
rect 19576 16892 19640 16896
rect 19576 16836 19580 16892
rect 19580 16836 19636 16892
rect 19636 16836 19640 16892
rect 19576 16832 19640 16836
rect 19656 16892 19720 16896
rect 19656 16836 19660 16892
rect 19660 16836 19716 16892
rect 19716 16836 19720 16892
rect 19656 16832 19720 16836
rect 19736 16892 19800 16896
rect 19736 16836 19740 16892
rect 19740 16836 19796 16892
rect 19796 16836 19800 16892
rect 19736 16832 19800 16836
rect 19816 16892 19880 16896
rect 19816 16836 19820 16892
rect 19820 16836 19876 16892
rect 19876 16836 19880 16892
rect 19816 16832 19880 16836
rect 4216 16348 4280 16352
rect 4216 16292 4220 16348
rect 4220 16292 4276 16348
rect 4276 16292 4280 16348
rect 4216 16288 4280 16292
rect 4296 16348 4360 16352
rect 4296 16292 4300 16348
rect 4300 16292 4356 16348
rect 4356 16292 4360 16348
rect 4296 16288 4360 16292
rect 4376 16348 4440 16352
rect 4376 16292 4380 16348
rect 4380 16292 4436 16348
rect 4436 16292 4440 16348
rect 4376 16288 4440 16292
rect 4456 16348 4520 16352
rect 4456 16292 4460 16348
rect 4460 16292 4516 16348
rect 4516 16292 4520 16348
rect 4456 16288 4520 16292
rect 34936 16348 35000 16352
rect 34936 16292 34940 16348
rect 34940 16292 34996 16348
rect 34996 16292 35000 16348
rect 34936 16288 35000 16292
rect 35016 16348 35080 16352
rect 35016 16292 35020 16348
rect 35020 16292 35076 16348
rect 35076 16292 35080 16348
rect 35016 16288 35080 16292
rect 35096 16348 35160 16352
rect 35096 16292 35100 16348
rect 35100 16292 35156 16348
rect 35156 16292 35160 16348
rect 35096 16288 35160 16292
rect 35176 16348 35240 16352
rect 35176 16292 35180 16348
rect 35180 16292 35236 16348
rect 35236 16292 35240 16348
rect 35176 16288 35240 16292
rect 19576 15804 19640 15808
rect 19576 15748 19580 15804
rect 19580 15748 19636 15804
rect 19636 15748 19640 15804
rect 19576 15744 19640 15748
rect 19656 15804 19720 15808
rect 19656 15748 19660 15804
rect 19660 15748 19716 15804
rect 19716 15748 19720 15804
rect 19656 15744 19720 15748
rect 19736 15804 19800 15808
rect 19736 15748 19740 15804
rect 19740 15748 19796 15804
rect 19796 15748 19800 15804
rect 19736 15744 19800 15748
rect 19816 15804 19880 15808
rect 19816 15748 19820 15804
rect 19820 15748 19876 15804
rect 19876 15748 19880 15804
rect 19816 15744 19880 15748
rect 4216 15260 4280 15264
rect 4216 15204 4220 15260
rect 4220 15204 4276 15260
rect 4276 15204 4280 15260
rect 4216 15200 4280 15204
rect 4296 15260 4360 15264
rect 4296 15204 4300 15260
rect 4300 15204 4356 15260
rect 4356 15204 4360 15260
rect 4296 15200 4360 15204
rect 4376 15260 4440 15264
rect 4376 15204 4380 15260
rect 4380 15204 4436 15260
rect 4436 15204 4440 15260
rect 4376 15200 4440 15204
rect 4456 15260 4520 15264
rect 4456 15204 4460 15260
rect 4460 15204 4516 15260
rect 4516 15204 4520 15260
rect 4456 15200 4520 15204
rect 34936 15260 35000 15264
rect 34936 15204 34940 15260
rect 34940 15204 34996 15260
rect 34996 15204 35000 15260
rect 34936 15200 35000 15204
rect 35016 15260 35080 15264
rect 35016 15204 35020 15260
rect 35020 15204 35076 15260
rect 35076 15204 35080 15260
rect 35016 15200 35080 15204
rect 35096 15260 35160 15264
rect 35096 15204 35100 15260
rect 35100 15204 35156 15260
rect 35156 15204 35160 15260
rect 35096 15200 35160 15204
rect 35176 15260 35240 15264
rect 35176 15204 35180 15260
rect 35180 15204 35236 15260
rect 35236 15204 35240 15260
rect 35176 15200 35240 15204
rect 19576 14716 19640 14720
rect 19576 14660 19580 14716
rect 19580 14660 19636 14716
rect 19636 14660 19640 14716
rect 19576 14656 19640 14660
rect 19656 14716 19720 14720
rect 19656 14660 19660 14716
rect 19660 14660 19716 14716
rect 19716 14660 19720 14716
rect 19656 14656 19720 14660
rect 19736 14716 19800 14720
rect 19736 14660 19740 14716
rect 19740 14660 19796 14716
rect 19796 14660 19800 14716
rect 19736 14656 19800 14660
rect 19816 14716 19880 14720
rect 19816 14660 19820 14716
rect 19820 14660 19876 14716
rect 19876 14660 19880 14716
rect 19816 14656 19880 14660
rect 4216 14172 4280 14176
rect 4216 14116 4220 14172
rect 4220 14116 4276 14172
rect 4276 14116 4280 14172
rect 4216 14112 4280 14116
rect 4296 14172 4360 14176
rect 4296 14116 4300 14172
rect 4300 14116 4356 14172
rect 4356 14116 4360 14172
rect 4296 14112 4360 14116
rect 4376 14172 4440 14176
rect 4376 14116 4380 14172
rect 4380 14116 4436 14172
rect 4436 14116 4440 14172
rect 4376 14112 4440 14116
rect 4456 14172 4520 14176
rect 4456 14116 4460 14172
rect 4460 14116 4516 14172
rect 4516 14116 4520 14172
rect 4456 14112 4520 14116
rect 34936 14172 35000 14176
rect 34936 14116 34940 14172
rect 34940 14116 34996 14172
rect 34996 14116 35000 14172
rect 34936 14112 35000 14116
rect 35016 14172 35080 14176
rect 35016 14116 35020 14172
rect 35020 14116 35076 14172
rect 35076 14116 35080 14172
rect 35016 14112 35080 14116
rect 35096 14172 35160 14176
rect 35096 14116 35100 14172
rect 35100 14116 35156 14172
rect 35156 14116 35160 14172
rect 35096 14112 35160 14116
rect 35176 14172 35240 14176
rect 35176 14116 35180 14172
rect 35180 14116 35236 14172
rect 35236 14116 35240 14172
rect 35176 14112 35240 14116
rect 19576 13628 19640 13632
rect 19576 13572 19580 13628
rect 19580 13572 19636 13628
rect 19636 13572 19640 13628
rect 19576 13568 19640 13572
rect 19656 13628 19720 13632
rect 19656 13572 19660 13628
rect 19660 13572 19716 13628
rect 19716 13572 19720 13628
rect 19656 13568 19720 13572
rect 19736 13628 19800 13632
rect 19736 13572 19740 13628
rect 19740 13572 19796 13628
rect 19796 13572 19800 13628
rect 19736 13568 19800 13572
rect 19816 13628 19880 13632
rect 19816 13572 19820 13628
rect 19820 13572 19876 13628
rect 19876 13572 19880 13628
rect 19816 13568 19880 13572
rect 4216 13084 4280 13088
rect 4216 13028 4220 13084
rect 4220 13028 4276 13084
rect 4276 13028 4280 13084
rect 4216 13024 4280 13028
rect 4296 13084 4360 13088
rect 4296 13028 4300 13084
rect 4300 13028 4356 13084
rect 4356 13028 4360 13084
rect 4296 13024 4360 13028
rect 4376 13084 4440 13088
rect 4376 13028 4380 13084
rect 4380 13028 4436 13084
rect 4436 13028 4440 13084
rect 4376 13024 4440 13028
rect 4456 13084 4520 13088
rect 4456 13028 4460 13084
rect 4460 13028 4516 13084
rect 4516 13028 4520 13084
rect 4456 13024 4520 13028
rect 34936 13084 35000 13088
rect 34936 13028 34940 13084
rect 34940 13028 34996 13084
rect 34996 13028 35000 13084
rect 34936 13024 35000 13028
rect 35016 13084 35080 13088
rect 35016 13028 35020 13084
rect 35020 13028 35076 13084
rect 35076 13028 35080 13084
rect 35016 13024 35080 13028
rect 35096 13084 35160 13088
rect 35096 13028 35100 13084
rect 35100 13028 35156 13084
rect 35156 13028 35160 13084
rect 35096 13024 35160 13028
rect 35176 13084 35240 13088
rect 35176 13028 35180 13084
rect 35180 13028 35236 13084
rect 35236 13028 35240 13084
rect 35176 13024 35240 13028
rect 19576 12540 19640 12544
rect 19576 12484 19580 12540
rect 19580 12484 19636 12540
rect 19636 12484 19640 12540
rect 19576 12480 19640 12484
rect 19656 12540 19720 12544
rect 19656 12484 19660 12540
rect 19660 12484 19716 12540
rect 19716 12484 19720 12540
rect 19656 12480 19720 12484
rect 19736 12540 19800 12544
rect 19736 12484 19740 12540
rect 19740 12484 19796 12540
rect 19796 12484 19800 12540
rect 19736 12480 19800 12484
rect 19816 12540 19880 12544
rect 19816 12484 19820 12540
rect 19820 12484 19876 12540
rect 19876 12484 19880 12540
rect 19816 12480 19880 12484
rect 4216 11996 4280 12000
rect 4216 11940 4220 11996
rect 4220 11940 4276 11996
rect 4276 11940 4280 11996
rect 4216 11936 4280 11940
rect 4296 11996 4360 12000
rect 4296 11940 4300 11996
rect 4300 11940 4356 11996
rect 4356 11940 4360 11996
rect 4296 11936 4360 11940
rect 4376 11996 4440 12000
rect 4376 11940 4380 11996
rect 4380 11940 4436 11996
rect 4436 11940 4440 11996
rect 4376 11936 4440 11940
rect 4456 11996 4520 12000
rect 4456 11940 4460 11996
rect 4460 11940 4516 11996
rect 4516 11940 4520 11996
rect 4456 11936 4520 11940
rect 34936 11996 35000 12000
rect 34936 11940 34940 11996
rect 34940 11940 34996 11996
rect 34996 11940 35000 11996
rect 34936 11936 35000 11940
rect 35016 11996 35080 12000
rect 35016 11940 35020 11996
rect 35020 11940 35076 11996
rect 35076 11940 35080 11996
rect 35016 11936 35080 11940
rect 35096 11996 35160 12000
rect 35096 11940 35100 11996
rect 35100 11940 35156 11996
rect 35156 11940 35160 11996
rect 35096 11936 35160 11940
rect 35176 11996 35240 12000
rect 35176 11940 35180 11996
rect 35180 11940 35236 11996
rect 35236 11940 35240 11996
rect 35176 11936 35240 11940
rect 19576 11452 19640 11456
rect 19576 11396 19580 11452
rect 19580 11396 19636 11452
rect 19636 11396 19640 11452
rect 19576 11392 19640 11396
rect 19656 11452 19720 11456
rect 19656 11396 19660 11452
rect 19660 11396 19716 11452
rect 19716 11396 19720 11452
rect 19656 11392 19720 11396
rect 19736 11452 19800 11456
rect 19736 11396 19740 11452
rect 19740 11396 19796 11452
rect 19796 11396 19800 11452
rect 19736 11392 19800 11396
rect 19816 11452 19880 11456
rect 19816 11396 19820 11452
rect 19820 11396 19876 11452
rect 19876 11396 19880 11452
rect 19816 11392 19880 11396
rect 4216 10908 4280 10912
rect 4216 10852 4220 10908
rect 4220 10852 4276 10908
rect 4276 10852 4280 10908
rect 4216 10848 4280 10852
rect 4296 10908 4360 10912
rect 4296 10852 4300 10908
rect 4300 10852 4356 10908
rect 4356 10852 4360 10908
rect 4296 10848 4360 10852
rect 4376 10908 4440 10912
rect 4376 10852 4380 10908
rect 4380 10852 4436 10908
rect 4436 10852 4440 10908
rect 4376 10848 4440 10852
rect 4456 10908 4520 10912
rect 4456 10852 4460 10908
rect 4460 10852 4516 10908
rect 4516 10852 4520 10908
rect 4456 10848 4520 10852
rect 34936 10908 35000 10912
rect 34936 10852 34940 10908
rect 34940 10852 34996 10908
rect 34996 10852 35000 10908
rect 34936 10848 35000 10852
rect 35016 10908 35080 10912
rect 35016 10852 35020 10908
rect 35020 10852 35076 10908
rect 35076 10852 35080 10908
rect 35016 10848 35080 10852
rect 35096 10908 35160 10912
rect 35096 10852 35100 10908
rect 35100 10852 35156 10908
rect 35156 10852 35160 10908
rect 35096 10848 35160 10852
rect 35176 10908 35240 10912
rect 35176 10852 35180 10908
rect 35180 10852 35236 10908
rect 35236 10852 35240 10908
rect 35176 10848 35240 10852
rect 19576 10364 19640 10368
rect 19576 10308 19580 10364
rect 19580 10308 19636 10364
rect 19636 10308 19640 10364
rect 19576 10304 19640 10308
rect 19656 10364 19720 10368
rect 19656 10308 19660 10364
rect 19660 10308 19716 10364
rect 19716 10308 19720 10364
rect 19656 10304 19720 10308
rect 19736 10364 19800 10368
rect 19736 10308 19740 10364
rect 19740 10308 19796 10364
rect 19796 10308 19800 10364
rect 19736 10304 19800 10308
rect 19816 10364 19880 10368
rect 19816 10308 19820 10364
rect 19820 10308 19876 10364
rect 19876 10308 19880 10364
rect 19816 10304 19880 10308
rect 4216 9820 4280 9824
rect 4216 9764 4220 9820
rect 4220 9764 4276 9820
rect 4276 9764 4280 9820
rect 4216 9760 4280 9764
rect 4296 9820 4360 9824
rect 4296 9764 4300 9820
rect 4300 9764 4356 9820
rect 4356 9764 4360 9820
rect 4296 9760 4360 9764
rect 4376 9820 4440 9824
rect 4376 9764 4380 9820
rect 4380 9764 4436 9820
rect 4436 9764 4440 9820
rect 4376 9760 4440 9764
rect 4456 9820 4520 9824
rect 4456 9764 4460 9820
rect 4460 9764 4516 9820
rect 4516 9764 4520 9820
rect 4456 9760 4520 9764
rect 34936 9820 35000 9824
rect 34936 9764 34940 9820
rect 34940 9764 34996 9820
rect 34996 9764 35000 9820
rect 34936 9760 35000 9764
rect 35016 9820 35080 9824
rect 35016 9764 35020 9820
rect 35020 9764 35076 9820
rect 35076 9764 35080 9820
rect 35016 9760 35080 9764
rect 35096 9820 35160 9824
rect 35096 9764 35100 9820
rect 35100 9764 35156 9820
rect 35156 9764 35160 9820
rect 35096 9760 35160 9764
rect 35176 9820 35240 9824
rect 35176 9764 35180 9820
rect 35180 9764 35236 9820
rect 35236 9764 35240 9820
rect 35176 9760 35240 9764
rect 19576 9276 19640 9280
rect 19576 9220 19580 9276
rect 19580 9220 19636 9276
rect 19636 9220 19640 9276
rect 19576 9216 19640 9220
rect 19656 9276 19720 9280
rect 19656 9220 19660 9276
rect 19660 9220 19716 9276
rect 19716 9220 19720 9276
rect 19656 9216 19720 9220
rect 19736 9276 19800 9280
rect 19736 9220 19740 9276
rect 19740 9220 19796 9276
rect 19796 9220 19800 9276
rect 19736 9216 19800 9220
rect 19816 9276 19880 9280
rect 19816 9220 19820 9276
rect 19820 9220 19876 9276
rect 19876 9220 19880 9276
rect 19816 9216 19880 9220
rect 4216 8732 4280 8736
rect 4216 8676 4220 8732
rect 4220 8676 4276 8732
rect 4276 8676 4280 8732
rect 4216 8672 4280 8676
rect 4296 8732 4360 8736
rect 4296 8676 4300 8732
rect 4300 8676 4356 8732
rect 4356 8676 4360 8732
rect 4296 8672 4360 8676
rect 4376 8732 4440 8736
rect 4376 8676 4380 8732
rect 4380 8676 4436 8732
rect 4436 8676 4440 8732
rect 4376 8672 4440 8676
rect 4456 8732 4520 8736
rect 4456 8676 4460 8732
rect 4460 8676 4516 8732
rect 4516 8676 4520 8732
rect 4456 8672 4520 8676
rect 34936 8732 35000 8736
rect 34936 8676 34940 8732
rect 34940 8676 34996 8732
rect 34996 8676 35000 8732
rect 34936 8672 35000 8676
rect 35016 8732 35080 8736
rect 35016 8676 35020 8732
rect 35020 8676 35076 8732
rect 35076 8676 35080 8732
rect 35016 8672 35080 8676
rect 35096 8732 35160 8736
rect 35096 8676 35100 8732
rect 35100 8676 35156 8732
rect 35156 8676 35160 8732
rect 35096 8672 35160 8676
rect 35176 8732 35240 8736
rect 35176 8676 35180 8732
rect 35180 8676 35236 8732
rect 35236 8676 35240 8732
rect 35176 8672 35240 8676
rect 19576 8188 19640 8192
rect 19576 8132 19580 8188
rect 19580 8132 19636 8188
rect 19636 8132 19640 8188
rect 19576 8128 19640 8132
rect 19656 8188 19720 8192
rect 19656 8132 19660 8188
rect 19660 8132 19716 8188
rect 19716 8132 19720 8188
rect 19656 8128 19720 8132
rect 19736 8188 19800 8192
rect 19736 8132 19740 8188
rect 19740 8132 19796 8188
rect 19796 8132 19800 8188
rect 19736 8128 19800 8132
rect 19816 8188 19880 8192
rect 19816 8132 19820 8188
rect 19820 8132 19876 8188
rect 19876 8132 19880 8188
rect 19816 8128 19880 8132
rect 4216 7644 4280 7648
rect 4216 7588 4220 7644
rect 4220 7588 4276 7644
rect 4276 7588 4280 7644
rect 4216 7584 4280 7588
rect 4296 7644 4360 7648
rect 4296 7588 4300 7644
rect 4300 7588 4356 7644
rect 4356 7588 4360 7644
rect 4296 7584 4360 7588
rect 4376 7644 4440 7648
rect 4376 7588 4380 7644
rect 4380 7588 4436 7644
rect 4436 7588 4440 7644
rect 4376 7584 4440 7588
rect 4456 7644 4520 7648
rect 4456 7588 4460 7644
rect 4460 7588 4516 7644
rect 4516 7588 4520 7644
rect 4456 7584 4520 7588
rect 34936 7644 35000 7648
rect 34936 7588 34940 7644
rect 34940 7588 34996 7644
rect 34996 7588 35000 7644
rect 34936 7584 35000 7588
rect 35016 7644 35080 7648
rect 35016 7588 35020 7644
rect 35020 7588 35076 7644
rect 35076 7588 35080 7644
rect 35016 7584 35080 7588
rect 35096 7644 35160 7648
rect 35096 7588 35100 7644
rect 35100 7588 35156 7644
rect 35156 7588 35160 7644
rect 35096 7584 35160 7588
rect 35176 7644 35240 7648
rect 35176 7588 35180 7644
rect 35180 7588 35236 7644
rect 35236 7588 35240 7644
rect 35176 7584 35240 7588
rect 19576 7100 19640 7104
rect 19576 7044 19580 7100
rect 19580 7044 19636 7100
rect 19636 7044 19640 7100
rect 19576 7040 19640 7044
rect 19656 7100 19720 7104
rect 19656 7044 19660 7100
rect 19660 7044 19716 7100
rect 19716 7044 19720 7100
rect 19656 7040 19720 7044
rect 19736 7100 19800 7104
rect 19736 7044 19740 7100
rect 19740 7044 19796 7100
rect 19796 7044 19800 7100
rect 19736 7040 19800 7044
rect 19816 7100 19880 7104
rect 19816 7044 19820 7100
rect 19820 7044 19876 7100
rect 19876 7044 19880 7100
rect 19816 7040 19880 7044
rect 4216 6556 4280 6560
rect 4216 6500 4220 6556
rect 4220 6500 4276 6556
rect 4276 6500 4280 6556
rect 4216 6496 4280 6500
rect 4296 6556 4360 6560
rect 4296 6500 4300 6556
rect 4300 6500 4356 6556
rect 4356 6500 4360 6556
rect 4296 6496 4360 6500
rect 4376 6556 4440 6560
rect 4376 6500 4380 6556
rect 4380 6500 4436 6556
rect 4436 6500 4440 6556
rect 4376 6496 4440 6500
rect 4456 6556 4520 6560
rect 4456 6500 4460 6556
rect 4460 6500 4516 6556
rect 4516 6500 4520 6556
rect 4456 6496 4520 6500
rect 34936 6556 35000 6560
rect 34936 6500 34940 6556
rect 34940 6500 34996 6556
rect 34996 6500 35000 6556
rect 34936 6496 35000 6500
rect 35016 6556 35080 6560
rect 35016 6500 35020 6556
rect 35020 6500 35076 6556
rect 35076 6500 35080 6556
rect 35016 6496 35080 6500
rect 35096 6556 35160 6560
rect 35096 6500 35100 6556
rect 35100 6500 35156 6556
rect 35156 6500 35160 6556
rect 35096 6496 35160 6500
rect 35176 6556 35240 6560
rect 35176 6500 35180 6556
rect 35180 6500 35236 6556
rect 35236 6500 35240 6556
rect 35176 6496 35240 6500
rect 19576 6012 19640 6016
rect 19576 5956 19580 6012
rect 19580 5956 19636 6012
rect 19636 5956 19640 6012
rect 19576 5952 19640 5956
rect 19656 6012 19720 6016
rect 19656 5956 19660 6012
rect 19660 5956 19716 6012
rect 19716 5956 19720 6012
rect 19656 5952 19720 5956
rect 19736 6012 19800 6016
rect 19736 5956 19740 6012
rect 19740 5956 19796 6012
rect 19796 5956 19800 6012
rect 19736 5952 19800 5956
rect 19816 6012 19880 6016
rect 19816 5956 19820 6012
rect 19820 5956 19876 6012
rect 19876 5956 19880 6012
rect 19816 5952 19880 5956
rect 4216 5468 4280 5472
rect 4216 5412 4220 5468
rect 4220 5412 4276 5468
rect 4276 5412 4280 5468
rect 4216 5408 4280 5412
rect 4296 5468 4360 5472
rect 4296 5412 4300 5468
rect 4300 5412 4356 5468
rect 4356 5412 4360 5468
rect 4296 5408 4360 5412
rect 4376 5468 4440 5472
rect 4376 5412 4380 5468
rect 4380 5412 4436 5468
rect 4436 5412 4440 5468
rect 4376 5408 4440 5412
rect 4456 5468 4520 5472
rect 4456 5412 4460 5468
rect 4460 5412 4516 5468
rect 4516 5412 4520 5468
rect 4456 5408 4520 5412
rect 34936 5468 35000 5472
rect 34936 5412 34940 5468
rect 34940 5412 34996 5468
rect 34996 5412 35000 5468
rect 34936 5408 35000 5412
rect 35016 5468 35080 5472
rect 35016 5412 35020 5468
rect 35020 5412 35076 5468
rect 35076 5412 35080 5468
rect 35016 5408 35080 5412
rect 35096 5468 35160 5472
rect 35096 5412 35100 5468
rect 35100 5412 35156 5468
rect 35156 5412 35160 5468
rect 35096 5408 35160 5412
rect 35176 5468 35240 5472
rect 35176 5412 35180 5468
rect 35180 5412 35236 5468
rect 35236 5412 35240 5468
rect 35176 5408 35240 5412
rect 19576 4924 19640 4928
rect 19576 4868 19580 4924
rect 19580 4868 19636 4924
rect 19636 4868 19640 4924
rect 19576 4864 19640 4868
rect 19656 4924 19720 4928
rect 19656 4868 19660 4924
rect 19660 4868 19716 4924
rect 19716 4868 19720 4924
rect 19656 4864 19720 4868
rect 19736 4924 19800 4928
rect 19736 4868 19740 4924
rect 19740 4868 19796 4924
rect 19796 4868 19800 4924
rect 19736 4864 19800 4868
rect 19816 4924 19880 4928
rect 19816 4868 19820 4924
rect 19820 4868 19876 4924
rect 19876 4868 19880 4924
rect 19816 4864 19880 4868
rect 4216 4380 4280 4384
rect 4216 4324 4220 4380
rect 4220 4324 4276 4380
rect 4276 4324 4280 4380
rect 4216 4320 4280 4324
rect 4296 4380 4360 4384
rect 4296 4324 4300 4380
rect 4300 4324 4356 4380
rect 4356 4324 4360 4380
rect 4296 4320 4360 4324
rect 4376 4380 4440 4384
rect 4376 4324 4380 4380
rect 4380 4324 4436 4380
rect 4436 4324 4440 4380
rect 4376 4320 4440 4324
rect 4456 4380 4520 4384
rect 4456 4324 4460 4380
rect 4460 4324 4516 4380
rect 4516 4324 4520 4380
rect 4456 4320 4520 4324
rect 34936 4380 35000 4384
rect 34936 4324 34940 4380
rect 34940 4324 34996 4380
rect 34996 4324 35000 4380
rect 34936 4320 35000 4324
rect 35016 4380 35080 4384
rect 35016 4324 35020 4380
rect 35020 4324 35076 4380
rect 35076 4324 35080 4380
rect 35016 4320 35080 4324
rect 35096 4380 35160 4384
rect 35096 4324 35100 4380
rect 35100 4324 35156 4380
rect 35156 4324 35160 4380
rect 35096 4320 35160 4324
rect 35176 4380 35240 4384
rect 35176 4324 35180 4380
rect 35180 4324 35236 4380
rect 35236 4324 35240 4380
rect 35176 4320 35240 4324
rect 24532 3980 24596 4044
rect 19576 3836 19640 3840
rect 19576 3780 19580 3836
rect 19580 3780 19636 3836
rect 19636 3780 19640 3836
rect 19576 3776 19640 3780
rect 19656 3836 19720 3840
rect 19656 3780 19660 3836
rect 19660 3780 19716 3836
rect 19716 3780 19720 3836
rect 19656 3776 19720 3780
rect 19736 3836 19800 3840
rect 19736 3780 19740 3836
rect 19740 3780 19796 3836
rect 19796 3780 19800 3836
rect 19736 3776 19800 3780
rect 19816 3836 19880 3840
rect 19816 3780 19820 3836
rect 19820 3780 19876 3836
rect 19876 3780 19880 3836
rect 19816 3776 19880 3780
rect 24348 3436 24412 3500
rect 4216 3292 4280 3296
rect 4216 3236 4220 3292
rect 4220 3236 4276 3292
rect 4276 3236 4280 3292
rect 4216 3232 4280 3236
rect 4296 3292 4360 3296
rect 4296 3236 4300 3292
rect 4300 3236 4356 3292
rect 4356 3236 4360 3292
rect 4296 3232 4360 3236
rect 4376 3292 4440 3296
rect 4376 3236 4380 3292
rect 4380 3236 4436 3292
rect 4436 3236 4440 3292
rect 4376 3232 4440 3236
rect 4456 3292 4520 3296
rect 4456 3236 4460 3292
rect 4460 3236 4516 3292
rect 4516 3236 4520 3292
rect 4456 3232 4520 3236
rect 34936 3292 35000 3296
rect 34936 3236 34940 3292
rect 34940 3236 34996 3292
rect 34996 3236 35000 3292
rect 34936 3232 35000 3236
rect 35016 3292 35080 3296
rect 35016 3236 35020 3292
rect 35020 3236 35076 3292
rect 35076 3236 35080 3292
rect 35016 3232 35080 3236
rect 35096 3292 35160 3296
rect 35096 3236 35100 3292
rect 35100 3236 35156 3292
rect 35156 3236 35160 3292
rect 35096 3232 35160 3236
rect 35176 3292 35240 3296
rect 35176 3236 35180 3292
rect 35180 3236 35236 3292
rect 35236 3236 35240 3292
rect 35176 3232 35240 3236
rect 19576 2748 19640 2752
rect 19576 2692 19580 2748
rect 19580 2692 19636 2748
rect 19636 2692 19640 2748
rect 19576 2688 19640 2692
rect 19656 2748 19720 2752
rect 19656 2692 19660 2748
rect 19660 2692 19716 2748
rect 19716 2692 19720 2748
rect 19656 2688 19720 2692
rect 19736 2748 19800 2752
rect 19736 2692 19740 2748
rect 19740 2692 19796 2748
rect 19796 2692 19800 2748
rect 19736 2688 19800 2692
rect 19816 2748 19880 2752
rect 19816 2692 19820 2748
rect 19820 2692 19876 2748
rect 19876 2692 19880 2748
rect 19816 2688 19880 2692
rect 4216 2204 4280 2208
rect 4216 2148 4220 2204
rect 4220 2148 4276 2204
rect 4276 2148 4280 2204
rect 4216 2144 4280 2148
rect 4296 2204 4360 2208
rect 4296 2148 4300 2204
rect 4300 2148 4356 2204
rect 4356 2148 4360 2204
rect 4296 2144 4360 2148
rect 4376 2204 4440 2208
rect 4376 2148 4380 2204
rect 4380 2148 4436 2204
rect 4436 2148 4440 2204
rect 4376 2144 4440 2148
rect 4456 2204 4520 2208
rect 4456 2148 4460 2204
rect 4460 2148 4516 2204
rect 4516 2148 4520 2204
rect 4456 2144 4520 2148
rect 34936 2204 35000 2208
rect 34936 2148 34940 2204
rect 34940 2148 34996 2204
rect 34996 2148 35000 2204
rect 34936 2144 35000 2148
rect 35016 2204 35080 2208
rect 35016 2148 35020 2204
rect 35020 2148 35076 2204
rect 35076 2148 35080 2204
rect 35016 2144 35080 2148
rect 35096 2204 35160 2208
rect 35096 2148 35100 2204
rect 35100 2148 35156 2204
rect 35156 2148 35160 2204
rect 35096 2144 35160 2148
rect 35176 2204 35240 2208
rect 35176 2148 35180 2204
rect 35180 2148 35236 2204
rect 35236 2148 35240 2204
rect 35176 2144 35240 2148
<< metal4 >>
rect 4208 37024 4528 37584
rect 4208 36960 4216 37024
rect 4280 36960 4296 37024
rect 4360 36960 4376 37024
rect 4440 36960 4456 37024
rect 4520 36960 4528 37024
rect 4208 35936 4528 36960
rect 4208 35872 4216 35936
rect 4280 35872 4296 35936
rect 4360 35872 4376 35936
rect 4440 35872 4456 35936
rect 4520 35872 4528 35936
rect 4208 34848 4528 35872
rect 4208 34784 4216 34848
rect 4280 34784 4296 34848
rect 4360 34784 4376 34848
rect 4440 34784 4456 34848
rect 4520 34784 4528 34848
rect 4208 33760 4528 34784
rect 4208 33696 4216 33760
rect 4280 33696 4296 33760
rect 4360 33696 4376 33760
rect 4440 33696 4456 33760
rect 4520 33696 4528 33760
rect 4208 32672 4528 33696
rect 4208 32608 4216 32672
rect 4280 32608 4296 32672
rect 4360 32608 4376 32672
rect 4440 32608 4456 32672
rect 4520 32608 4528 32672
rect 4208 31584 4528 32608
rect 4208 31520 4216 31584
rect 4280 31520 4296 31584
rect 4360 31520 4376 31584
rect 4440 31520 4456 31584
rect 4520 31520 4528 31584
rect 4208 30496 4528 31520
rect 4208 30432 4216 30496
rect 4280 30432 4296 30496
rect 4360 30432 4376 30496
rect 4440 30432 4456 30496
rect 4520 30432 4528 30496
rect 4208 29408 4528 30432
rect 4208 29344 4216 29408
rect 4280 29344 4296 29408
rect 4360 29344 4376 29408
rect 4440 29344 4456 29408
rect 4520 29344 4528 29408
rect 4208 28320 4528 29344
rect 4208 28256 4216 28320
rect 4280 28256 4296 28320
rect 4360 28256 4376 28320
rect 4440 28256 4456 28320
rect 4520 28256 4528 28320
rect 4208 27232 4528 28256
rect 4208 27168 4216 27232
rect 4280 27168 4296 27232
rect 4360 27168 4376 27232
rect 4440 27168 4456 27232
rect 4520 27168 4528 27232
rect 4208 26144 4528 27168
rect 4208 26080 4216 26144
rect 4280 26080 4296 26144
rect 4360 26080 4376 26144
rect 4440 26080 4456 26144
rect 4520 26080 4528 26144
rect 4208 25056 4528 26080
rect 4208 24992 4216 25056
rect 4280 24992 4296 25056
rect 4360 24992 4376 25056
rect 4440 24992 4456 25056
rect 4520 24992 4528 25056
rect 4208 23968 4528 24992
rect 4208 23904 4216 23968
rect 4280 23904 4296 23968
rect 4360 23904 4376 23968
rect 4440 23904 4456 23968
rect 4520 23904 4528 23968
rect 4208 22880 4528 23904
rect 4208 22816 4216 22880
rect 4280 22816 4296 22880
rect 4360 22816 4376 22880
rect 4440 22816 4456 22880
rect 4520 22816 4528 22880
rect 4208 21792 4528 22816
rect 4208 21728 4216 21792
rect 4280 21728 4296 21792
rect 4360 21728 4376 21792
rect 4440 21728 4456 21792
rect 4520 21728 4528 21792
rect 4208 20704 4528 21728
rect 4208 20640 4216 20704
rect 4280 20640 4296 20704
rect 4360 20640 4376 20704
rect 4440 20640 4456 20704
rect 4520 20640 4528 20704
rect 4208 19616 4528 20640
rect 4208 19552 4216 19616
rect 4280 19552 4296 19616
rect 4360 19552 4376 19616
rect 4440 19552 4456 19616
rect 4520 19552 4528 19616
rect 4208 18528 4528 19552
rect 4208 18464 4216 18528
rect 4280 18464 4296 18528
rect 4360 18464 4376 18528
rect 4440 18464 4456 18528
rect 4520 18464 4528 18528
rect 4208 17440 4528 18464
rect 4208 17376 4216 17440
rect 4280 17376 4296 17440
rect 4360 17376 4376 17440
rect 4440 17376 4456 17440
rect 4520 17376 4528 17440
rect 4208 16352 4528 17376
rect 4208 16288 4216 16352
rect 4280 16288 4296 16352
rect 4360 16288 4376 16352
rect 4440 16288 4456 16352
rect 4520 16288 4528 16352
rect 4208 15264 4528 16288
rect 4208 15200 4216 15264
rect 4280 15200 4296 15264
rect 4360 15200 4376 15264
rect 4440 15200 4456 15264
rect 4520 15200 4528 15264
rect 4208 14176 4528 15200
rect 4208 14112 4216 14176
rect 4280 14112 4296 14176
rect 4360 14112 4376 14176
rect 4440 14112 4456 14176
rect 4520 14112 4528 14176
rect 4208 13088 4528 14112
rect 4208 13024 4216 13088
rect 4280 13024 4296 13088
rect 4360 13024 4376 13088
rect 4440 13024 4456 13088
rect 4520 13024 4528 13088
rect 4208 12000 4528 13024
rect 4208 11936 4216 12000
rect 4280 11936 4296 12000
rect 4360 11936 4376 12000
rect 4440 11936 4456 12000
rect 4520 11936 4528 12000
rect 4208 10912 4528 11936
rect 4208 10848 4216 10912
rect 4280 10848 4296 10912
rect 4360 10848 4376 10912
rect 4440 10848 4456 10912
rect 4520 10848 4528 10912
rect 4208 9824 4528 10848
rect 4208 9760 4216 9824
rect 4280 9760 4296 9824
rect 4360 9760 4376 9824
rect 4440 9760 4456 9824
rect 4520 9760 4528 9824
rect 4208 8736 4528 9760
rect 4208 8672 4216 8736
rect 4280 8672 4296 8736
rect 4360 8672 4376 8736
rect 4440 8672 4456 8736
rect 4520 8672 4528 8736
rect 4208 7648 4528 8672
rect 4208 7584 4216 7648
rect 4280 7584 4296 7648
rect 4360 7584 4376 7648
rect 4440 7584 4456 7648
rect 4520 7584 4528 7648
rect 4208 6560 4528 7584
rect 4208 6496 4216 6560
rect 4280 6496 4296 6560
rect 4360 6496 4376 6560
rect 4440 6496 4456 6560
rect 4520 6496 4528 6560
rect 4208 5472 4528 6496
rect 4208 5408 4216 5472
rect 4280 5408 4296 5472
rect 4360 5408 4376 5472
rect 4440 5408 4456 5472
rect 4520 5408 4528 5472
rect 4208 4384 4528 5408
rect 4208 4320 4216 4384
rect 4280 4320 4296 4384
rect 4360 4320 4376 4384
rect 4440 4320 4456 4384
rect 4520 4320 4528 4384
rect 4208 3296 4528 4320
rect 4208 3232 4216 3296
rect 4280 3232 4296 3296
rect 4360 3232 4376 3296
rect 4440 3232 4456 3296
rect 4520 3232 4528 3296
rect 4208 2208 4528 3232
rect 4208 2144 4216 2208
rect 4280 2144 4296 2208
rect 4360 2144 4376 2208
rect 4440 2144 4456 2208
rect 4520 2144 4528 2208
rect 4208 2128 4528 2144
rect 19568 37568 19888 37584
rect 19568 37504 19576 37568
rect 19640 37504 19656 37568
rect 19720 37504 19736 37568
rect 19800 37504 19816 37568
rect 19880 37504 19888 37568
rect 19568 36480 19888 37504
rect 19568 36416 19576 36480
rect 19640 36416 19656 36480
rect 19720 36416 19736 36480
rect 19800 36416 19816 36480
rect 19880 36416 19888 36480
rect 19568 35392 19888 36416
rect 19568 35328 19576 35392
rect 19640 35328 19656 35392
rect 19720 35328 19736 35392
rect 19800 35328 19816 35392
rect 19880 35328 19888 35392
rect 19568 34304 19888 35328
rect 19568 34240 19576 34304
rect 19640 34240 19656 34304
rect 19720 34240 19736 34304
rect 19800 34240 19816 34304
rect 19880 34240 19888 34304
rect 19568 33216 19888 34240
rect 19568 33152 19576 33216
rect 19640 33152 19656 33216
rect 19720 33152 19736 33216
rect 19800 33152 19816 33216
rect 19880 33152 19888 33216
rect 19568 32128 19888 33152
rect 19568 32064 19576 32128
rect 19640 32064 19656 32128
rect 19720 32064 19736 32128
rect 19800 32064 19816 32128
rect 19880 32064 19888 32128
rect 19568 31040 19888 32064
rect 19568 30976 19576 31040
rect 19640 30976 19656 31040
rect 19720 30976 19736 31040
rect 19800 30976 19816 31040
rect 19880 30976 19888 31040
rect 19568 29952 19888 30976
rect 34928 37024 35248 37584
rect 34928 36960 34936 37024
rect 35000 36960 35016 37024
rect 35080 36960 35096 37024
rect 35160 36960 35176 37024
rect 35240 36960 35248 37024
rect 34928 35936 35248 36960
rect 34928 35872 34936 35936
rect 35000 35872 35016 35936
rect 35080 35872 35096 35936
rect 35160 35872 35176 35936
rect 35240 35872 35248 35936
rect 34928 34848 35248 35872
rect 34928 34784 34936 34848
rect 35000 34784 35016 34848
rect 35080 34784 35096 34848
rect 35160 34784 35176 34848
rect 35240 34784 35248 34848
rect 34928 33760 35248 34784
rect 34928 33696 34936 33760
rect 35000 33696 35016 33760
rect 35080 33696 35096 33760
rect 35160 33696 35176 33760
rect 35240 33696 35248 33760
rect 34928 32672 35248 33696
rect 34928 32608 34936 32672
rect 35000 32608 35016 32672
rect 35080 32608 35096 32672
rect 35160 32608 35176 32672
rect 35240 32608 35248 32672
rect 34928 31584 35248 32608
rect 34928 31520 34936 31584
rect 35000 31520 35016 31584
rect 35080 31520 35096 31584
rect 35160 31520 35176 31584
rect 35240 31520 35248 31584
rect 34928 30496 35248 31520
rect 34928 30432 34936 30496
rect 35000 30432 35016 30496
rect 35080 30432 35096 30496
rect 35160 30432 35176 30496
rect 35240 30432 35248 30496
rect 24531 30428 24597 30429
rect 24531 30364 24532 30428
rect 24596 30364 24597 30428
rect 24531 30363 24597 30364
rect 19568 29888 19576 29952
rect 19640 29888 19656 29952
rect 19720 29888 19736 29952
rect 19800 29888 19816 29952
rect 19880 29888 19888 29952
rect 19568 28864 19888 29888
rect 19568 28800 19576 28864
rect 19640 28800 19656 28864
rect 19720 28800 19736 28864
rect 19800 28800 19816 28864
rect 19880 28800 19888 28864
rect 19568 27776 19888 28800
rect 19568 27712 19576 27776
rect 19640 27712 19656 27776
rect 19720 27712 19736 27776
rect 19800 27712 19816 27776
rect 19880 27712 19888 27776
rect 19568 26688 19888 27712
rect 19568 26624 19576 26688
rect 19640 26624 19656 26688
rect 19720 26624 19736 26688
rect 19800 26624 19816 26688
rect 19880 26624 19888 26688
rect 19568 25600 19888 26624
rect 19568 25536 19576 25600
rect 19640 25536 19656 25600
rect 19720 25536 19736 25600
rect 19800 25536 19816 25600
rect 19880 25536 19888 25600
rect 19568 24512 19888 25536
rect 24347 24988 24413 24989
rect 24347 24924 24348 24988
rect 24412 24924 24413 24988
rect 24347 24923 24413 24924
rect 19568 24448 19576 24512
rect 19640 24448 19656 24512
rect 19720 24448 19736 24512
rect 19800 24448 19816 24512
rect 19880 24448 19888 24512
rect 19568 23424 19888 24448
rect 19568 23360 19576 23424
rect 19640 23360 19656 23424
rect 19720 23360 19736 23424
rect 19800 23360 19816 23424
rect 19880 23360 19888 23424
rect 19568 22336 19888 23360
rect 19568 22272 19576 22336
rect 19640 22272 19656 22336
rect 19720 22272 19736 22336
rect 19800 22272 19816 22336
rect 19880 22272 19888 22336
rect 19568 21248 19888 22272
rect 19568 21184 19576 21248
rect 19640 21184 19656 21248
rect 19720 21184 19736 21248
rect 19800 21184 19816 21248
rect 19880 21184 19888 21248
rect 19568 20160 19888 21184
rect 19568 20096 19576 20160
rect 19640 20096 19656 20160
rect 19720 20096 19736 20160
rect 19800 20096 19816 20160
rect 19880 20096 19888 20160
rect 19568 19072 19888 20096
rect 19568 19008 19576 19072
rect 19640 19008 19656 19072
rect 19720 19008 19736 19072
rect 19800 19008 19816 19072
rect 19880 19008 19888 19072
rect 19568 17984 19888 19008
rect 19568 17920 19576 17984
rect 19640 17920 19656 17984
rect 19720 17920 19736 17984
rect 19800 17920 19816 17984
rect 19880 17920 19888 17984
rect 19568 16896 19888 17920
rect 19568 16832 19576 16896
rect 19640 16832 19656 16896
rect 19720 16832 19736 16896
rect 19800 16832 19816 16896
rect 19880 16832 19888 16896
rect 19568 15808 19888 16832
rect 19568 15744 19576 15808
rect 19640 15744 19656 15808
rect 19720 15744 19736 15808
rect 19800 15744 19816 15808
rect 19880 15744 19888 15808
rect 19568 14720 19888 15744
rect 19568 14656 19576 14720
rect 19640 14656 19656 14720
rect 19720 14656 19736 14720
rect 19800 14656 19816 14720
rect 19880 14656 19888 14720
rect 19568 13632 19888 14656
rect 19568 13568 19576 13632
rect 19640 13568 19656 13632
rect 19720 13568 19736 13632
rect 19800 13568 19816 13632
rect 19880 13568 19888 13632
rect 19568 12544 19888 13568
rect 19568 12480 19576 12544
rect 19640 12480 19656 12544
rect 19720 12480 19736 12544
rect 19800 12480 19816 12544
rect 19880 12480 19888 12544
rect 19568 11456 19888 12480
rect 19568 11392 19576 11456
rect 19640 11392 19656 11456
rect 19720 11392 19736 11456
rect 19800 11392 19816 11456
rect 19880 11392 19888 11456
rect 19568 10368 19888 11392
rect 19568 10304 19576 10368
rect 19640 10304 19656 10368
rect 19720 10304 19736 10368
rect 19800 10304 19816 10368
rect 19880 10304 19888 10368
rect 19568 9280 19888 10304
rect 19568 9216 19576 9280
rect 19640 9216 19656 9280
rect 19720 9216 19736 9280
rect 19800 9216 19816 9280
rect 19880 9216 19888 9280
rect 19568 8192 19888 9216
rect 19568 8128 19576 8192
rect 19640 8128 19656 8192
rect 19720 8128 19736 8192
rect 19800 8128 19816 8192
rect 19880 8128 19888 8192
rect 19568 7104 19888 8128
rect 19568 7040 19576 7104
rect 19640 7040 19656 7104
rect 19720 7040 19736 7104
rect 19800 7040 19816 7104
rect 19880 7040 19888 7104
rect 19568 6016 19888 7040
rect 19568 5952 19576 6016
rect 19640 5952 19656 6016
rect 19720 5952 19736 6016
rect 19800 5952 19816 6016
rect 19880 5952 19888 6016
rect 19568 4928 19888 5952
rect 19568 4864 19576 4928
rect 19640 4864 19656 4928
rect 19720 4864 19736 4928
rect 19800 4864 19816 4928
rect 19880 4864 19888 4928
rect 19568 3840 19888 4864
rect 19568 3776 19576 3840
rect 19640 3776 19656 3840
rect 19720 3776 19736 3840
rect 19800 3776 19816 3840
rect 19880 3776 19888 3840
rect 19568 2752 19888 3776
rect 24350 3501 24410 24923
rect 24534 4045 24594 30363
rect 34928 29408 35248 30432
rect 34928 29344 34936 29408
rect 35000 29344 35016 29408
rect 35080 29344 35096 29408
rect 35160 29344 35176 29408
rect 35240 29344 35248 29408
rect 34928 28320 35248 29344
rect 34928 28256 34936 28320
rect 35000 28256 35016 28320
rect 35080 28256 35096 28320
rect 35160 28256 35176 28320
rect 35240 28256 35248 28320
rect 34928 27232 35248 28256
rect 34928 27168 34936 27232
rect 35000 27168 35016 27232
rect 35080 27168 35096 27232
rect 35160 27168 35176 27232
rect 35240 27168 35248 27232
rect 34928 26144 35248 27168
rect 34928 26080 34936 26144
rect 35000 26080 35016 26144
rect 35080 26080 35096 26144
rect 35160 26080 35176 26144
rect 35240 26080 35248 26144
rect 34928 25056 35248 26080
rect 34928 24992 34936 25056
rect 35000 24992 35016 25056
rect 35080 24992 35096 25056
rect 35160 24992 35176 25056
rect 35240 24992 35248 25056
rect 34928 23968 35248 24992
rect 34928 23904 34936 23968
rect 35000 23904 35016 23968
rect 35080 23904 35096 23968
rect 35160 23904 35176 23968
rect 35240 23904 35248 23968
rect 34928 22880 35248 23904
rect 34928 22816 34936 22880
rect 35000 22816 35016 22880
rect 35080 22816 35096 22880
rect 35160 22816 35176 22880
rect 35240 22816 35248 22880
rect 34928 21792 35248 22816
rect 34928 21728 34936 21792
rect 35000 21728 35016 21792
rect 35080 21728 35096 21792
rect 35160 21728 35176 21792
rect 35240 21728 35248 21792
rect 34928 20704 35248 21728
rect 34928 20640 34936 20704
rect 35000 20640 35016 20704
rect 35080 20640 35096 20704
rect 35160 20640 35176 20704
rect 35240 20640 35248 20704
rect 34928 19616 35248 20640
rect 34928 19552 34936 19616
rect 35000 19552 35016 19616
rect 35080 19552 35096 19616
rect 35160 19552 35176 19616
rect 35240 19552 35248 19616
rect 34928 18528 35248 19552
rect 34928 18464 34936 18528
rect 35000 18464 35016 18528
rect 35080 18464 35096 18528
rect 35160 18464 35176 18528
rect 35240 18464 35248 18528
rect 34928 17440 35248 18464
rect 34928 17376 34936 17440
rect 35000 17376 35016 17440
rect 35080 17376 35096 17440
rect 35160 17376 35176 17440
rect 35240 17376 35248 17440
rect 34928 16352 35248 17376
rect 34928 16288 34936 16352
rect 35000 16288 35016 16352
rect 35080 16288 35096 16352
rect 35160 16288 35176 16352
rect 35240 16288 35248 16352
rect 34928 15264 35248 16288
rect 34928 15200 34936 15264
rect 35000 15200 35016 15264
rect 35080 15200 35096 15264
rect 35160 15200 35176 15264
rect 35240 15200 35248 15264
rect 34928 14176 35248 15200
rect 34928 14112 34936 14176
rect 35000 14112 35016 14176
rect 35080 14112 35096 14176
rect 35160 14112 35176 14176
rect 35240 14112 35248 14176
rect 34928 13088 35248 14112
rect 34928 13024 34936 13088
rect 35000 13024 35016 13088
rect 35080 13024 35096 13088
rect 35160 13024 35176 13088
rect 35240 13024 35248 13088
rect 34928 12000 35248 13024
rect 34928 11936 34936 12000
rect 35000 11936 35016 12000
rect 35080 11936 35096 12000
rect 35160 11936 35176 12000
rect 35240 11936 35248 12000
rect 34928 10912 35248 11936
rect 34928 10848 34936 10912
rect 35000 10848 35016 10912
rect 35080 10848 35096 10912
rect 35160 10848 35176 10912
rect 35240 10848 35248 10912
rect 34928 9824 35248 10848
rect 34928 9760 34936 9824
rect 35000 9760 35016 9824
rect 35080 9760 35096 9824
rect 35160 9760 35176 9824
rect 35240 9760 35248 9824
rect 34928 8736 35248 9760
rect 34928 8672 34936 8736
rect 35000 8672 35016 8736
rect 35080 8672 35096 8736
rect 35160 8672 35176 8736
rect 35240 8672 35248 8736
rect 34928 7648 35248 8672
rect 34928 7584 34936 7648
rect 35000 7584 35016 7648
rect 35080 7584 35096 7648
rect 35160 7584 35176 7648
rect 35240 7584 35248 7648
rect 34928 6560 35248 7584
rect 34928 6496 34936 6560
rect 35000 6496 35016 6560
rect 35080 6496 35096 6560
rect 35160 6496 35176 6560
rect 35240 6496 35248 6560
rect 34928 5472 35248 6496
rect 34928 5408 34936 5472
rect 35000 5408 35016 5472
rect 35080 5408 35096 5472
rect 35160 5408 35176 5472
rect 35240 5408 35248 5472
rect 34928 4384 35248 5408
rect 34928 4320 34936 4384
rect 35000 4320 35016 4384
rect 35080 4320 35096 4384
rect 35160 4320 35176 4384
rect 35240 4320 35248 4384
rect 24531 4044 24597 4045
rect 24531 3980 24532 4044
rect 24596 3980 24597 4044
rect 24531 3979 24597 3980
rect 24347 3500 24413 3501
rect 24347 3436 24348 3500
rect 24412 3436 24413 3500
rect 24347 3435 24413 3436
rect 19568 2688 19576 2752
rect 19640 2688 19656 2752
rect 19720 2688 19736 2752
rect 19800 2688 19816 2752
rect 19880 2688 19888 2752
rect 19568 2128 19888 2688
rect 34928 3296 35248 4320
rect 34928 3232 34936 3296
rect 35000 3232 35016 3296
rect 35080 3232 35096 3296
rect 35160 3232 35176 3296
rect 35240 3232 35248 3296
rect 34928 2208 35248 3232
rect 34928 2144 34936 2208
rect 35000 2144 35016 2208
rect 35080 2144 35096 2208
rect 35160 2144 35176 2208
rect 35240 2144 35248 2208
rect 34928 2128 35248 2144
use sky130_fd_sc_hd__decap_4  FILLER_1_12 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 2208 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 1380 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 3128 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1608254825
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _2509_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 2576 0 1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _2500_
timestamp 1608254825
transform 1 0 1380 0 -1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_2  _1908_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 1932 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_43
timestamp 1608254825
transform 1 0 5060 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_35
timestamp 1608254825
transform 1 0 4324 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32
timestamp 1608254825
transform 1 0 4048 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 3864 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2533_
timestamp 1608254825
transform 1 0 4600 0 -1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  _1915_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 4692 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_57
timestamp 1608254825
transform 1 0 6348 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_47
timestamp 1608254825
transform 1 0 5428 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57
timestamp 1608254825
transform 1 0 6348 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_4  _2343_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 5520 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_0_66
timestamp 1608254825
transform 1 0 7176 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61
timestamp 1608254825
transform 1 0 6716 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1608254825
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1608254825
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _2342_
timestamp 1608254825
transform 1 0 6900 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _2518_
timestamp 1608254825
transform 1 0 6808 0 1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_1_90
timestamp 1608254825
transform 1 0 9384 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_85
timestamp 1608254825
transform 1 0 8924 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_81
timestamp 1608254825
transform 1 0 8556 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_91 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 9476 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_83
timestamp 1608254825
transform 1 0 8740 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_4  _2344_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 7544 0 -1 2720
box -38 -48 1234 592
use sky130_fd_sc_hd__buf_2  _1912_
timestamp 1608254825
transform 1 0 9016 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_114
timestamp 1608254825
transform 1 0 11592 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_94
timestamp 1608254825
transform 1 0 9752 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_97
timestamp 1608254825
transform 1 0 10028 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1608254825
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2526_
timestamp 1608254825
transform 1 0 10396 0 -1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _2415_
timestamp 1608254825
transform 1 0 9844 0 1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_2  _1923_
timestamp 1608254825
transform 1 0 9752 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_136
timestamp 1608254825
transform 1 0 13616 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_132
timestamp 1608254825
transform 1 0 13248 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_120
timestamp 1608254825
transform 1 0 12144 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1608254825
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1608254825
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2520_
timestamp 1608254825
transform 1 0 12420 0 1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__and2_4  _1931_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 12604 0 -1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1925_
timestamp 1608254825
transform 1 0 13708 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_142
timestamp 1608254825
transform 1 0 14168 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_156
timestamp 1608254825
transform 1 0 15456 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_151
timestamp 1608254825
transform 1 0 14996 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_140
timestamp 1608254825
transform 1 0 13984 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1608254825
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2529_
timestamp 1608254825
transform 1 0 14536 0 1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _2525_
timestamp 1608254825
transform 1 0 15640 0 -1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__and2_4  _1951_
timestamp 1608254825
transform 1 0 14352 0 -1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_1_179
timestamp 1608254825
transform 1 0 17572 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_169
timestamp 1608254825
transform 1 0 16652 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_165
timestamp 1608254825
transform 1 0 16284 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_177
timestamp 1608254825
transform 1 0 17388 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_4  _1914_
timestamp 1608254825
transform 1 0 16744 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_1_203
timestamp 1608254825
transform 1 0 19780 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_190
timestamp 1608254825
transform 1 0 18584 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_185
timestamp 1608254825
transform 1 0 18124 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1608254825
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1608254825
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2528_
timestamp 1608254825
transform 1 0 18032 0 1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _2524_
timestamp 1608254825
transform 1 0 18952 0 -1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_2  _2277_
timestamp 1608254825
transform 1 0 18308 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_211
timestamp 1608254825
transform 1 0 20516 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_213
timestamp 1608254825
transform 1 0 20700 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1608254825
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2537_
timestamp 1608254825
transform 1 0 21160 0 -1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _2527_
timestamp 1608254825
transform 1 0 20608 0 1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_1_240
timestamp 1608254825
transform 1 0 23184 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_231
timestamp 1608254825
transform 1 0 22356 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_249
timestamp 1608254825
transform 1 0 24012 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_245
timestamp 1608254825
transform 1 0 23644 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_237
timestamp 1608254825
transform 1 0 22908 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1608254825
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1608254825
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2402_
timestamp 1608254825
transform 1 0 23644 0 1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_2  _1636_
timestamp 1608254825
transform 1 0 22908 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_1_264
timestamp 1608254825
transform 1 0 25392 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_274
timestamp 1608254825
transform 1 0 26312 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2523_
timestamp 1608254825
transform 1 0 24564 0 -1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _2514_
timestamp 1608254825
transform 1 0 25944 0 1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_1_296
timestamp 1608254825
transform 1 0 28336 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_289
timestamp 1608254825
transform 1 0 27692 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_278
timestamp 1608254825
transform 1 0 26680 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1608254825
transform 1 0 26772 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2531_
timestamp 1608254825
transform 1 0 26864 0 -1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_2  _1773_
timestamp 1608254825
transform 1 0 28060 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_304
timestamp 1608254825
transform 1 0 29072 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_307
timestamp 1608254825
transform 1 0 29348 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_299
timestamp 1608254825
transform 1 0 28612 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1608254825
transform 1 0 29164 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_318
timestamp 1608254825
transform 1 0 30360 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_314
timestamp 1608254825
transform 1 0 29992 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1608254825
transform 1 0 29624 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _2357_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 29716 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _2579_
timestamp 1608254825
transform 1 0 30360 0 -1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__o21a_4  _1792_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 29256 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_326
timestamp 1608254825
transform 1 0 31096 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_342
timestamp 1608254825
transform 1 0 32568 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_337
timestamp 1608254825
transform 1 0 32108 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1608254825
transform 1 0 32476 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2578_
timestamp 1608254825
transform 1 0 31188 0 1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_1_362
timestamp 1608254825
transform 1 0 34408 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_346
timestamp 1608254825
transform 1 0 32936 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_346
timestamp 1608254825
transform 1 0 32936 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_4 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 33028 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _2510_
timestamp 1608254825
transform 1 0 33212 0 -1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__o21a_4  _1812_
timestamp 1608254825
transform 1 0 33304 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_383
timestamp 1608254825
transform 1 0 36340 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_379
timestamp 1608254825
transform 1 0 35972 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_385
timestamp 1608254825
transform 1 0 36524 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_368
timestamp 1608254825
transform 1 0 34960 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1608254825
transform 1 0 34776 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1608254825
transform 1 0 35328 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2512_
timestamp 1608254825
transform 1 0 36432 0 1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__o21a_4  _1817_
timestamp 1608254825
transform 1 0 35420 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__o21a_4  _1815_
timestamp 1608254825
transform 1 0 34868 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_403
timestamp 1608254825
transform 1 0 38180 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_404
timestamp 1608254825
transform 1 0 38272 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_397
timestamp 1608254825
transform 1 0 37628 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_393
timestamp 1608254825
transform 1 0 37260 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1608254825
transform 1 0 38180 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1608254825
transform -1 0 38824 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1608254825
transform -1 0 38824 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2358_
timestamp 1608254825
transform 1 0 37352 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_7
timestamp 1608254825
transform 1 0 1748 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_3
timestamp 1608254825
transform 1 0 1380 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1608254825
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _2539_
timestamp 1608254825
transform 1 0 1840 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_2_40
timestamp 1608254825
transform 1 0 4784 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_32
timestamp 1608254825
transform 1 0 4048 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_27
timestamp 1608254825
transform 1 0 3588 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1608254825
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2431_
timestamp 1608254825
transform 1 0 5152 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__and2_4  _1919_
timestamp 1608254825
transform 1 0 4140 0 -1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_2_67
timestamp 1608254825
transform 1 0 7268 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_63
timestamp 1608254825
transform 1 0 6900 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__and2_4  _1955_
timestamp 1608254825
transform 1 0 7360 0 -1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_2_88
timestamp 1608254825
transform 1 0 9200 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_75
timestamp 1608254825
transform 1 0 8004 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_4  _1924_
timestamp 1608254825
transform 1 0 8372 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_2_112
timestamp 1608254825
transform 1 0 11408 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1608254825
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2530_
timestamp 1608254825
transform 1 0 9660 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_2_120
timestamp 1608254825
transform 1 0 12144 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2522_
timestamp 1608254825
transform 1 0 12512 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  _1921_
timestamp 1608254825
transform 1 0 11776 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_151
timestamp 1608254825
transform 1 0 14996 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_143
timestamp 1608254825
transform 1 0 14260 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1608254825
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _1926_
timestamp 1608254825
transform 1 0 15272 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_2_167
timestamp 1608254825
transform 1 0 16468 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_163
timestamp 1608254825
transform 1 0 16100 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2411_
timestamp 1608254825
transform 1 0 16560 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_2_195
timestamp 1608254825
transform 1 0 19044 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_187
timestamp 1608254825
transform 1 0 18308 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_4  _2135_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 19228 0 -1 3808
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_2_210
timestamp 1608254825
transform 1 0 20424 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1608254825
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__nand3_4  _2134_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 20884 0 -1 3808
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_2_251
timestamp 1608254825
transform 1 0 24196 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_229
timestamp 1608254825
transform 1 0 22172 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__a2bb2o_4  _2314_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 22724 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_2_271
timestamp 1608254825
transform 1 0 26036 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_4  _2317_
timestamp 1608254825
transform 1 0 24564 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_2_286
timestamp 1608254825
transform 1 0 27416 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_279
timestamp 1608254825
transform 1 0 26772 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1608254825
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2584_
timestamp 1608254825
transform 1 0 27784 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_2  _1765_
timestamp 1608254825
transform 1 0 27140 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1750_
timestamp 1608254825
transform 1 0 26496 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_309
timestamp 1608254825
transform 1 0 29532 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_4  _1797_
timestamp 1608254825
transform 1 0 29900 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_337
timestamp 1608254825
transform 1 0 32108 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_2_333
timestamp 1608254825
transform 1 0 31740 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_325
timestamp 1608254825
transform 1 0 31004 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1608254825
transform 1 0 32016 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_363
timestamp 1608254825
transform 1 0 34500 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_343
timestamp 1608254825
transform 1 0 32660 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2577_
timestamp 1608254825
transform 1 0 32752 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_2_386
timestamp 1608254825
transform 1 0 36616 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _2576_
timestamp 1608254825
transform 1 0 34868 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_2_406
timestamp 1608254825
transform 1 0 38456 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_402
timestamp 1608254825
transform 1 0 38088 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_2_394
timestamp 1608254825
transform 1 0 37352 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1608254825
transform 1 0 37628 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1608254825
transform -1 0 38824 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1810_
timestamp 1608254825
transform 1 0 37720 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_19
timestamp 1608254825
transform 1 0 2852 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_15
timestamp 1608254825
transform 1 0 2484 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_3_3
timestamp 1608254825
transform 1 0 1380 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1608254825
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _2429_
timestamp 1608254825
transform 1 0 2944 0 1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__nor2_4  _1905_
timestamp 1608254825
transform 1 0 1656 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_3_39
timestamp 1608254825
transform 1 0 4692 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_4  _1909_
timestamp 1608254825
transform 1 0 5060 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_3_60
timestamp 1608254825
transform 1 0 6624 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_52
timestamp 1608254825
transform 1 0 5888 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1608254825
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2433_
timestamp 1608254825
transform 1 0 6808 0 1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_3_89
timestamp 1608254825
transform 1 0 9292 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_81
timestamp 1608254825
transform 1 0 8556 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__o32ai_4  _2285_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 9384 0 1 3808
box -38 -48 2062 592
use sky130_fd_sc_hd__decap_8  FILLER_3_112
timestamp 1608254825
transform 1 0 11408 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_133
timestamp 1608254825
transform 1 0 13340 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_126
timestamp 1608254825
transform 1 0 12696 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_120
timestamp 1608254825
transform 1 0 12144 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1608254825
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _1953_
timestamp 1608254825
transform 1 0 13708 0 1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1844_
timestamp 1608254825
transform 1 0 13064 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1743_
timestamp 1608254825
transform 1 0 12420 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_144
timestamp 1608254825
transform 1 0 14352 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2413_
timestamp 1608254825
transform 1 0 14720 0 1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_3_179
timestamp 1608254825
transform 1 0 17572 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_171
timestamp 1608254825
transform 1 0 16836 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_167
timestamp 1608254825
transform 1 0 16468 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__and2_4  _1933_
timestamp 1608254825
transform 1 0 16928 0 1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_3_203
timestamp 1608254825
transform 1 0 19780 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1608254825
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2444_
timestamp 1608254825
transform 1 0 18032 0 1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_3_226
timestamp 1608254825
transform 1 0 21896 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2443_
timestamp 1608254825
transform 1 0 20148 0 1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_3_243
timestamp 1608254825
transform 1 0 23460 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_237
timestamp 1608254825
transform 1 0 22908 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1608254825
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _1934_
timestamp 1608254825
transform 1 0 23644 0 1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _1922_
timestamp 1608254825
transform 1 0 22264 0 1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_3_252
timestamp 1608254825
transform 1 0 24288 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  _2399_
timestamp 1608254825
transform 1 0 24840 0 1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_3_285
timestamp 1608254825
transform 1 0 27324 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_277
timestamp 1608254825
transform 1 0 26588 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_4  _1798_
timestamp 1608254825
transform 1 0 27692 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _1497_
timestamp 1608254825
transform 1 0 26956 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_301
timestamp 1608254825
transform 1 0 28796 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1608254825
transform 1 0 29164 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2587_
timestamp 1608254825
transform 1 0 29256 0 1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_3_331
timestamp 1608254825
transform 1 0 31556 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_325
timestamp 1608254825
transform 1 0 31004 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_4  _1811_
timestamp 1608254825
transform 1 0 31648 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_360
timestamp 1608254825
transform 1 0 34224 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_344
timestamp 1608254825
transform 1 0 32752 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_4  _1814_
timestamp 1608254825
transform 1 0 33120 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_372
timestamp 1608254825
transform 1 0 35328 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_367
timestamp 1608254825
transform 1 0 34868 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1608254825
transform 1 0 34776 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2575_
timestamp 1608254825
transform 1 0 36064 0 1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  _1788_
timestamp 1608254825
transform 1 0 34960 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_399
timestamp 1608254825
transform 1 0 37812 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1608254825
transform -1 0 38824 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_4_22
timestamp 1608254825
transform 1 0 3128 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1608254825
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _2541_
timestamp 1608254825
transform 1 0 1380 0 -1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_4_39
timestamp 1608254825
transform 1 0 4692 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_32
timestamp 1608254825
transform 1 0 4048 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_30
timestamp 1608254825
transform 1 0 3864 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1608254825
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__o32ai_4  _2252_
timestamp 1608254825
transform 1 0 5060 0 -1 4896
box -38 -48 2062 592
use sky130_fd_sc_hd__inv_2  _1904_
timestamp 1608254825
transform 1 0 4416 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_65
timestamp 1608254825
transform 1 0 7084 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_88
timestamp 1608254825
transform 1 0 9200 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2414_
timestamp 1608254825
transform 1 0 7452 0 -1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_4_93
timestamp 1608254825
transform 1 0 9660 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1608254825
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__o32ai_4  _2284_
timestamp 1608254825
transform 1 0 10028 0 -1 4896
box -38 -48 2062 592
use sky130_fd_sc_hd__decap_4  FILLER_4_119
timestamp 1608254825
transform 1 0 12052 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2416_
timestamp 1608254825
transform 1 0 12420 0 -1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_4_154
timestamp 1608254825
transform 1 0 15272 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_149
timestamp 1608254825
transform 1 0 14812 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_142
timestamp 1608254825
transform 1 0 14168 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1608254825
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _1932_
timestamp 1608254825
transform 1 0 15640 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1619_
timestamp 1608254825
transform 1 0 14536 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_4_165
timestamp 1608254825
transform 1 0 16284 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__o32ai_4  _2288_
timestamp 1608254825
transform 1 0 16836 0 -1 4896
box -38 -48 2062 592
use sky130_fd_sc_hd__decap_4  FILLER_4_193
timestamp 1608254825
transform 1 0 18860 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_4  _2132_
timestamp 1608254825
transform 1 0 19228 0 -1 4896
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_1  FILLER_4_222
timestamp 1608254825
transform 1 0 21528 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_218
timestamp 1608254825
transform 1 0 21160 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_210
timestamp 1608254825
transform 1 0 20424 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1608254825
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__nand3_4  _2130_
timestamp 1608254825
transform 1 0 21620 0 -1 4896
box -38 -48 1326 592
use sky130_fd_sc_hd__inv_2  _1929_
timestamp 1608254825
transform 1 0 20884 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_244
timestamp 1608254825
transform 1 0 23552 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_237
timestamp 1608254825
transform 1 0 22908 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_4  _2316_
timestamp 1608254825
transform 1 0 23920 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  _2223_
timestamp 1608254825
transform 1 0 23276 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_271
timestamp 1608254825
transform 1 0 26036 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_264
timestamp 1608254825
transform 1 0 25392 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1713_
timestamp 1608254825
transform 1 0 25760 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_276
timestamp 1608254825
transform 1 0 26496 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1608254825
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2586_
timestamp 1608254825
transform 1 0 26772 0 -1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_4_306
timestamp 1608254825
transform 1 0 29256 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_298
timestamp 1608254825
transform 1 0 28520 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_4  _1791_
timestamp 1608254825
transform 1 0 29440 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_328
timestamp 1608254825
transform 1 0 31280 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_320
timestamp 1608254825
transform 1 0 30544 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1608254825
transform 1 0 32016 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_4  _1796_
timestamp 1608254825
transform 1 0 32108 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _1790_
timestamp 1608254825
transform 1 0 30912 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_365
timestamp 1608254825
transform 1 0 34684 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_349
timestamp 1608254825
transform 1 0 33212 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_4  _1800_
timestamp 1608254825
transform 1 0 33580 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_381
timestamp 1608254825
transform 1 0 36156 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_4  _1816_
timestamp 1608254825
transform 1 0 35052 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _1813_
timestamp 1608254825
transform 1 0 36524 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_406
timestamp 1608254825
transform 1 0 38456 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_402
timestamp 1608254825
transform 1 0 38088 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_389
timestamp 1608254825
transform 1 0 36892 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1608254825
transform 1 0 37628 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1608254825
transform -1 0 38824 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1809_
timestamp 1608254825
transform 1 0 37720 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_16
timestamp 1608254825
transform 1 0 2576 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_5_3
timestamp 1608254825
transform 1 0 1380 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1608254825
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__and2_4  _1917_
timestamp 1608254825
transform 1 0 1932 0 1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__o32ai_4  _2256_
timestamp 1608254825
transform 1 0 3312 0 1 4896
box -38 -48 2062 592
use sky130_fd_sc_hd__decap_4  FILLER_5_65
timestamp 1608254825
transform 1 0 7084 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_57
timestamp 1608254825
transform 1 0 6348 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_52
timestamp 1608254825
transform 1 0 5888 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_46
timestamp 1608254825
transform 1 0 5336 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1608254825
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1950_
timestamp 1608254825
transform 1 0 5980 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1709_
timestamp 1608254825
transform 1 0 6808 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_88
timestamp 1608254825
transform 1 0 9200 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2417_
timestamp 1608254825
transform 1 0 7452 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_5_114
timestamp 1608254825
transform 1 0 11592 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__o32ai_4  _2282_
timestamp 1608254825
transform 1 0 9568 0 1 4896
box -38 -48 2062 592
use sky130_fd_sc_hd__decap_4  FILLER_5_132
timestamp 1608254825
transform 1 0 13248 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_127
timestamp 1608254825
transform 1 0 12788 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_123
timestamp 1608254825
transform 1 0 12420 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1608254825
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__o32ai_4  _2281_
timestamp 1608254825
transform 1 0 13616 0 1 4896
box -38 -48 2062 592
use sky130_fd_sc_hd__buf_2  _2280_
timestamp 1608254825
transform 1 0 12880 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_158
timestamp 1608254825
transform 1 0 15640 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_182
timestamp 1608254825
transform 1 0 17848 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_176
timestamp 1608254825
transform 1 0 17296 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_166
timestamp 1608254825
transform 1 0 16376 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _1928_
timestamp 1608254825
transform 1 0 16468 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_5_199
timestamp 1608254825
transform 1 0 19412 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_193
timestamp 1608254825
transform 1 0 18860 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1608254825
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__nand3_4  _2131_
timestamp 1608254825
transform 1 0 19504 0 1 4896
box -38 -48 1326 592
use sky130_fd_sc_hd__nor2_4  _1930_
timestamp 1608254825
transform 1 0 18032 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_5_222
timestamp 1608254825
transform 1 0 21528 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_214
timestamp 1608254825
transform 1 0 20792 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_4  _2127_
timestamp 1608254825
transform 1 0 21896 0 1 4896
box -38 -48 1326 592
use sky130_fd_sc_hd__buf_2  _2120_
timestamp 1608254825
transform 1 0 21160 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_249
timestamp 1608254825
transform 1 0 24012 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_5_240
timestamp 1608254825
transform 1 0 23184 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1608254825
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1873_
timestamp 1608254825
transform 1 0 23644 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_257
timestamp 1608254825
transform 1 0 24748 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _2400_
timestamp 1608254825
transform 1 0 24932 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_5_278
timestamp 1608254825
transform 1 0 26680 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2583_
timestamp 1608254825
transform 1 0 27048 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_5_306
timestamp 1608254825
transform 1 0 29256 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_301
timestamp 1608254825
transform 1 0 28796 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1608254825
transform 1 0 29164 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_4  _1793_
timestamp 1608254825
transform 1 0 29808 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_332
timestamp 1608254825
transform 1 0 31648 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_324
timestamp 1608254825
transform 1 0 30912 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_4  _1795_
timestamp 1608254825
transform 1 0 31924 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_363
timestamp 1608254825
transform 1 0 34500 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_355
timestamp 1608254825
transform 1 0 33764 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_5_347
timestamp 1608254825
transform 1 0 33028 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1462_
timestamp 1608254825
transform 1 0 33396 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_379
timestamp 1608254825
transform 1 0 35972 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1608254825
transform 1 0 34776 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2574_
timestamp 1608254825
transform 1 0 36340 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__o21a_4  _1801_
timestamp 1608254825
transform 1 0 34868 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_406
timestamp 1608254825
transform 1 0 38456 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_402
timestamp 1608254825
transform 1 0 38088 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1608254825
transform -1 0 38824 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_7_16
timestamp 1608254825
transform 1 0 2576 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_7_3
timestamp 1608254825
transform 1 0 1380 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_22
timestamp 1608254825
transform 1 0 3128 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1608254825
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1608254825
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _2535_
timestamp 1608254825
transform 1 0 1380 0 -1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__nor2_4  _1903_
timestamp 1608254825
transform 1 0 1748 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_7_24
timestamp 1608254825
transform 1 0 3312 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_42
timestamp 1608254825
transform 1 0 4968 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_36
timestamp 1608254825
transform 1 0 4416 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_32
timestamp 1608254825
transform 1 0 4048 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_30
timestamp 1608254825
transform 1 0 3864 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1608254825
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__o32ai_4  _2251_
timestamp 1608254825
transform 1 0 3404 0 1 5984
box -38 -48 2062 592
use sky130_fd_sc_hd__inv_2  _1902_
timestamp 1608254825
transform 1 0 4140 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1847_
timestamp 1608254825
transform 1 0 5060 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_66
timestamp 1608254825
transform 1 0 7176 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_55
timestamp 1608254825
transform 1 0 6164 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_47
timestamp 1608254825
transform 1 0 5428 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_46
timestamp 1608254825
transform 1 0 5336 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1608254825
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__o32ai_4  _2250_
timestamp 1608254825
transform 1 0 5704 0 -1 5984
box -38 -48 2062 592
use sky130_fd_sc_hd__buf_2  _2249_
timestamp 1608254825
transform 1 0 5796 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _2244_
timestamp 1608254825
transform 1 0 6808 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_89
timestamp 1608254825
transform 1 0 9292 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_91
timestamp 1608254825
transform 1 0 9476 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_83
timestamp 1608254825
transform 1 0 8740 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_72
timestamp 1608254825
transform 1 0 7728 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_0_0_addressalyzerBlock.SPI_CLK $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 8096 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _2426_
timestamp 1608254825
transform 1 0 7544 0 1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  _1935_
timestamp 1608254825
transform 1 0 8372 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_95
timestamp 1608254825
transform 1 0 9844 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_96
timestamp 1608254825
transform 1 0 9936 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1608254825
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _1710_
timestamp 1608254825
transform 1 0 9936 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1622_
timestamp 1608254825
transform 1 0 9660 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_105
timestamp 1608254825
transform 1 0 10764 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_102
timestamp 1608254825
transform 1 0 10488 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _1939_
timestamp 1608254825
transform 1 0 10580 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_4  _1936_
timestamp 1608254825
transform 1 0 11132 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_6_112
timestamp 1608254825
transform 1 0 11408 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_126
timestamp 1608254825
transform 1 0 12696 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_118
timestamp 1608254825
transform 1 0 11960 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_addressalyzerBlock.SPI_CLK
timestamp 1608254825
transform 1 0 13064 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1608254825
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2418_
timestamp 1608254825
transform 1 0 13340 0 1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__o32ai_4  _2283_
timestamp 1608254825
transform 1 0 11776 0 -1 5984
box -38 -48 2062 592
use sky130_fd_sc_hd__inv_2  _1705_
timestamp 1608254825
transform 1 0 12420 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_159
timestamp 1608254825
transform 1 0 15732 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_152
timestamp 1608254825
transform 1 0 15088 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_149
timestamp 1608254825
transform 1 0 14812 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_144
timestamp 1608254825
transform 1 0 14352 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_138
timestamp 1608254825
transform 1 0 13800 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_2_0_addressalyzerBlock.SPI_CLK
timestamp 1608254825
transform 1 0 15456 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1608254825
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__o32ai_4  _2286_
timestamp 1608254825
transform 1 0 15272 0 -1 5984
box -38 -48 2062 592
use sky130_fd_sc_hd__buf_2  _2278_
timestamp 1608254825
transform 1 0 14444 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_179
timestamp 1608254825
transform 1 0 17572 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_176
timestamp 1608254825
transform 1 0 17296 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2427_
timestamp 1608254825
transform 1 0 15824 0 1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  _2276_
timestamp 1608254825
transform 1 0 17664 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_191
timestamp 1608254825
transform 1 0 18676 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_187
timestamp 1608254825
transform 1 0 18308 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_192
timestamp 1608254825
transform 1 0 18768 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_184
timestamp 1608254825
transform 1 0 18032 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1608254825
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2445_
timestamp 1608254825
transform 1 0 18768 0 1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__o21ai_4  _2129_
timestamp 1608254825
transform 1 0 18952 0 -1 5984
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _1913_
timestamp 1608254825
transform 1 0 18032 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_7_211
timestamp 1608254825
transform 1 0 20516 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_213
timestamp 1608254825
transform 1 0 20700 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_207
timestamp 1608254825
transform 1 0 20148 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1608254825
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _2136_
timestamp 1608254825
transform 1 0 20884 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_219
timestamp 1608254825
transform 1 0 21252 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_225
timestamp 1608254825
transform 1 0 21804 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_218
timestamp 1608254825
transform 1 0 21160 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2119_
timestamp 1608254825
transform 1 0 21528 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_4  _2253_
timestamp 1608254825
transform 1 0 21344 0 1 5984
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_7_249
timestamp 1608254825
transform 1 0 24012 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_242
timestamp 1608254825
transform 1 0 23368 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_234
timestamp 1608254825
transform 1 0 22632 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_6_243
timestamp 1608254825
transform 1 0 23460 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1608254825
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _2318_
timestamp 1608254825
transform 1 0 24012 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__nand3_4  _2122_
timestamp 1608254825
transform 1 0 22172 0 -1 5984
box -38 -48 1326 592
use sky130_fd_sc_hd__buf_2  _1789_
timestamp 1608254825
transform 1 0 23644 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_258
timestamp 1608254825
transform 1 0 24840 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_253
timestamp 1608254825
transform 1 0 24380 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_273
timestamp 1608254825
transform 1 0 26220 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_265
timestamp 1608254825
transform 1 0 25484 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _2398_
timestamp 1608254825
transform 1 0 25208 0 1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  _1824_
timestamp 1608254825
transform 1 0 24472 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_281
timestamp 1608254825
transform 1 0 26956 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_288
timestamp 1608254825
transform 1 0 27600 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_6_276
timestamp 1608254825
transform 1 0 26496 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1608254825
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_4  _1823_
timestamp 1608254825
transform 1 0 27692 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__o21a_4  _1822_
timestamp 1608254825
transform 1 0 27968 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__and4_4  _1777_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 26772 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_7_301
timestamp 1608254825
transform 1 0 28796 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_304
timestamp 1608254825
transform 1 0 29072 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1608254825
transform 1 0 29164 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2608_
timestamp 1608254825
transform 1 0 29256 0 1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__o21a_4  _1794_
timestamp 1608254825
transform 1 0 29440 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_333
timestamp 1608254825
transform 1 0 31740 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_325
timestamp 1608254825
transform 1 0 31004 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_332
timestamp 1608254825
transform 1 0 31648 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_320
timestamp 1608254825
transform 1 0 30544 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1608254825
transform 1 0 32016 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2585_
timestamp 1608254825
transform 1 0 32108 0 -1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__o21a_4  _1821_
timestamp 1608254825
transform 1 0 31832 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _1477_
timestamp 1608254825
transform 1 0 31280 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_362
timestamp 1608254825
transform 1 0 34408 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_346
timestamp 1608254825
transform 1 0 32936 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_356
timestamp 1608254825
transform 1 0 33856 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  _2582_
timestamp 1608254825
transform 1 0 34408 0 -1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__o21a_4  _1819_
timestamp 1608254825
transform 1 0 33304 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_380
timestamp 1608254825
transform 1 0 36064 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_367
timestamp 1608254825
transform 1 0 34868 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_381
timestamp 1608254825
transform 1 0 36156 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1608254825
transform 1 0 34776 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_4  _1818_
timestamp 1608254825
transform 1 0 36432 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__o21a_4  _1802_
timestamp 1608254825
transform 1 0 34960 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _1787_
timestamp 1608254825
transform 1 0 36524 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_396
timestamp 1608254825
transform 1 0 37536 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_389
timestamp 1608254825
transform 1 0 36892 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1608254825
transform 1 0 37628 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_403
timestamp 1608254825
transform 1 0 38180 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_402
timestamp 1608254825
transform 1 0 38088 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1838_
timestamp 1608254825
transform 1 0 37720 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1808_
timestamp 1608254825
transform 1 0 37904 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_406
timestamp 1608254825
transform 1 0 38456 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1608254825
transform -1 0 38824 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1608254825
transform -1 0 38824 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_7
timestamp 1608254825
transform 1 0 1748 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_3
timestamp 1608254825
transform 1 0 1380 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1608254825
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _2432_
timestamp 1608254825
transform 1 0 1840 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_8_27
timestamp 1608254825
transform 1 0 3588 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_188
timestamp 1608254825
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__o32ai_4  _2254_
timestamp 1608254825
transform 1 0 4048 0 -1 7072
box -38 -48 2062 592
use sky130_fd_sc_hd__decap_4  FILLER_8_54
timestamp 1608254825
transform 1 0 6072 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2424_
timestamp 1608254825
transform 1 0 6440 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_8_91
timestamp 1608254825
transform 1 0 9476 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_85
timestamp 1608254825
transform 1 0 8924 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_77
timestamp 1608254825
transform 1 0 8188 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1625_
timestamp 1608254825
transform 1 0 8556 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_107
timestamp 1608254825
transform 1 0 10948 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_97
timestamp 1608254825
transform 1 0 10028 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_93
timestamp 1608254825
transform 1 0 9660 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_189
timestamp 1608254825
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _1706_
timestamp 1608254825
transform 1 0 10120 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_8_128
timestamp 1608254825
transform 1 0 12880 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_4  _2220_
timestamp 1608254825
transform 1 0 13432 0 -1 7072
box -38 -48 1234 592
use sky130_fd_sc_hd__a21oi_4  _1848_
timestamp 1608254825
transform 1 0 11684 0 -1 7072
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_6  FILLER_8_147
timestamp 1608254825
transform 1 0 14628 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_190
timestamp 1608254825
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_4  _2174_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 15272 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_8_163
timestamp 1608254825
transform 1 0 16100 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_3_0_addressalyzerBlock.SPI_CLK
timestamp 1608254825
transform 1 0 16468 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__o32ai_4  _2261_
timestamp 1608254825
transform 1 0 16744 0 -1 7072
box -38 -48 2062 592
use sky130_fd_sc_hd__decap_4  FILLER_8_192
timestamp 1608254825
transform 1 0 18768 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_4  _2260_
timestamp 1608254825
transform 1 0 19136 0 -1 7072
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_8_228
timestamp 1608254825
transform 1 0 22080 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_223
timestamp 1608254825
transform 1 0 21620 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_219
timestamp 1608254825
transform 1 0 21252 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_210
timestamp 1608254825
transform 1 0 20424 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_191
timestamp 1608254825
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _2311_
timestamp 1608254825
transform 1 0 21712 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _2123_
timestamp 1608254825
transform 1 0 20884 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_250
timestamp 1608254825
transform 1 0 24104 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_246
timestamp 1608254825
transform 1 0 23736 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2401_
timestamp 1608254825
transform 1 0 24196 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__nand3_4  _2133_
timestamp 1608254825
transform 1 0 22448 0 -1 7072
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_1  FILLER_8_274
timestamp 1608254825
transform 1 0 26312 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_270
timestamp 1608254825
transform 1 0 25944 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_294
timestamp 1608254825
transform 1 0 28152 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_276
timestamp 1608254825
transform 1 0 26496 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_192
timestamp 1608254825
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__a22oi_4  _1775_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 26588 0 -1 7072
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_8  FILLER_8_312
timestamp 1608254825
transform 1 0 29808 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_298
timestamp 1608254825
transform 1 0 28520 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_4  _1502_
timestamp 1608254825
transform 1 0 28612 0 -1 7072
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_8_332
timestamp 1608254825
transform 1 0 31648 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_193
timestamp 1608254825
transform 1 0 32016 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__a21o_4  _1516_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 30544 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__and4_4  _1457_
timestamp 1608254825
transform 1 0 32108 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_8_363
timestamp 1608254825
transform 1 0 34500 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_350
timestamp 1608254825
transform 1 0 33304 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_346
timestamp 1608254825
transform 1 0 32936 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_4  _1820_
timestamp 1608254825
transform 1 0 33396 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_386
timestamp 1608254825
transform 1 0 36616 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_8_379
timestamp 1608254825
transform 1 0 35972 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_4  _1803_
timestamp 1608254825
transform 1 0 34868 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1786_
timestamp 1608254825
transform 1 0 36340 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_406
timestamp 1608254825
transform 1 0 38456 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_398
timestamp 1608254825
transform 1 0 37720 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_394
timestamp 1608254825
transform 1 0 37352 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_194
timestamp 1608254825
transform 1 0 37628 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1608254825
transform -1 0 38824 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_15
timestamp 1608254825
transform 1 0 2484 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 1380 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1608254825
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _2430_
timestamp 1608254825
transform 1 0 2576 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_9_35
timestamp 1608254825
transform 1 0 4324 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_4  _2177_
timestamp 1608254825
transform 1 0 4692 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_9_62
timestamp 1608254825
transform 1 0 6808 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_57
timestamp 1608254825
transform 1 0 6348 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_52
timestamp 1608254825
transform 1 0 5888 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_48
timestamp 1608254825
transform 1 0 5520 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_195
timestamp 1608254825
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _2247_
timestamp 1608254825
transform 1 0 5980 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _2150_
timestamp 1608254825
transform 1 0 7084 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_69
timestamp 1608254825
transform 1 0 7452 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__o32ai_4  _2265_
timestamp 1608254825
transform 1 0 7820 0 1 7072
box -38 -48 2062 592
use sky130_fd_sc_hd__fill_1  FILLER_9_104
timestamp 1608254825
transform 1 0 10672 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_95
timestamp 1608254825
transform 1 0 9844 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_addressalyzerBlock.SPI_CLK
timestamp 1608254825
transform 1 0 10396 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_4  _1849_
timestamp 1608254825
transform 1 0 10764 0 1 7072
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_9_131
timestamp 1608254825
transform 1 0 13156 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_127
timestamp 1608254825
transform 1 0 12788 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_123
timestamp 1608254825
transform 1 0 12420 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_118
timestamp 1608254825
transform 1 0 11960 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_196
timestamp 1608254825
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _2243_
timestamp 1608254825
transform 1 0 12880 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_4  _1626_
timestamp 1608254825
transform 1 0 13524 0 1 7072
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_6  FILLER_9_148
timestamp 1608254825
transform 1 0 14720 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  _2412_
timestamp 1608254825
transform 1 0 15272 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_9_181
timestamp 1608254825
transform 1 0 17756 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_173
timestamp 1608254825
transform 1 0 17020 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_9_197
timestamp 1608254825
transform 1 0 19228 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_184
timestamp 1608254825
transform 1 0 18032 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_197
timestamp 1608254825
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__nand3_4  _2128_
timestamp 1608254825
transform 1 0 19596 0 1 7072
box -38 -48 1326 592
use sky130_fd_sc_hd__nor2_4  _1714_
timestamp 1608254825
transform 1 0 18400 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 1608254825
transform 1 0 21620 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_215
timestamp 1608254825
transform 1 0 20884 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__nand3_4  _2255_
timestamp 1608254825
transform 1 0 21712 0 1 7072
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_6  FILLER_9_238
timestamp 1608254825
transform 1 0 23000 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_198
timestamp 1608254825
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _2315_
timestamp 1608254825
transform 1 0 23644 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_9_271
timestamp 1608254825
transform 1 0 26036 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_261
timestamp 1608254825
transform 1 0 25116 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _1485_
timestamp 1608254825
transform 1 0 25668 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_292
timestamp 1608254825
transform 1 0 27968 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__a22oi_4  _1774_
timestamp 1608254825
transform 1 0 26404 0 1 7072
box -38 -48 1602 592
use sky130_fd_sc_hd__buf_2  _1459_
timestamp 1608254825
transform 1 0 28336 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_318
timestamp 1608254825
transform 1 0 30360 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_304
timestamp 1608254825
transform 1 0 29072 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_300
timestamp 1608254825
transform 1 0 28704 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_199
timestamp 1608254825
transform 1 0 29164 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__a21o_4  _1501_
timestamp 1608254825
transform 1 0 29256 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _2606_
timestamp 1608254825
transform 1 0 30912 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_9_365
timestamp 1608254825
transform 1 0 34684 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_361
timestamp 1608254825
transform 1 0 34316 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_347
timestamp 1608254825
transform 1 0 33028 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_343
timestamp 1608254825
transform 1 0 32660 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_4  _1478_
timestamp 1608254825
transform 1 0 33120 0 1 7072
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_9_380
timestamp 1608254825
transform 1 0 36064 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_367
timestamp 1608254825
transform 1 0 34868 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_200
timestamp 1608254825
transform 1 0 34776 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2573_
timestamp 1608254825
transform 1 0 36432 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__o21a_4  _1807_
timestamp 1608254825
transform 1 0 34960 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_403
timestamp 1608254825
transform 1 0 38180 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1608254825
transform -1 0 38824 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_10_22
timestamp 1608254825
transform 1 0 3128 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1608254825
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _2542_
timestamp 1608254825
transform 1 0 1380 0 -1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_10_43
timestamp 1608254825
transform 1 0 5060 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_10_32
timestamp 1608254825
transform 1 0 4048 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_30
timestamp 1608254825
transform 1 0 3864 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_201
timestamp 1608254825
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_4  _2154_
timestamp 1608254825
transform 1 0 4232 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_10_53
timestamp 1608254825
transform 1 0 5980 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__o32ai_4  _2269_
timestamp 1608254825
transform 1 0 6348 0 -1 8160
box -38 -48 2062 592
use sky130_fd_sc_hd__buf_2  _2258_
timestamp 1608254825
transform 1 0 5612 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_91
timestamp 1608254825
transform 1 0 9476 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_87
timestamp 1608254825
transform 1 0 9108 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_79
timestamp 1608254825
transform 1 0 8372 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1624_
timestamp 1608254825
transform 1 0 8740 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_112
timestamp 1608254825
transform 1 0 11408 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_108
timestamp 1608254825
transform 1 0 11040 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_93
timestamp 1608254825
transform 1 0 9660 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_202
timestamp 1608254825
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _1744_
timestamp 1608254825
transform 1 0 10212 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _1704_
timestamp 1608254825
transform 1 0 11500 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_136
timestamp 1608254825
transform 1 0 13616 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_117
timestamp 1608254825
transform 1 0 11868 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_4  _1627_
timestamp 1608254825
transform 1 0 12420 0 -1 8160
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_10_154
timestamp 1608254825
transform 1 0 15272 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_149
timestamp 1608254825
transform 1 0 14812 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_203
timestamp 1608254825
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__o32ai_4  _2287_
timestamp 1608254825
transform 1 0 15640 0 -1 8160
box -38 -48 2062 592
use sky130_fd_sc_hd__nor2_4  _1620_
timestamp 1608254825
transform 1 0 13984 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_10_180
timestamp 1608254825
transform 1 0 17664 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_10_200
timestamp 1608254825
transform 1 0 19504 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_4  _1852_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 18216 0 -1 8160
box -38 -48 1326 592
use sky130_fd_sc_hd__buf_2  _1631_
timestamp 1608254825
transform 1 0 19872 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_224
timestamp 1608254825
transform 1 0 21712 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_10_208
timestamp 1608254825
transform 1 0 20240 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_204
timestamp 1608254825
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _1751_
timestamp 1608254825
transform 1 0 20884 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_10_246
timestamp 1608254825
transform 1 0 23736 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_4  _2319_
timestamp 1608254825
transform 1 0 22264 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__nand3_4  _2257_
timestamp 1608254825
transform 1 0 24104 0 -1 8160
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_10_271
timestamp 1608254825
transform 1 0 26036 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_264
timestamp 1608254825
transform 1 0 25392 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1499_
timestamp 1608254825
transform 1 0 25760 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_296
timestamp 1608254825
transform 1 0 28336 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_10_276
timestamp 1608254825
transform 1 0 26496 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_205
timestamp 1608254825
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__a22oi_4  _1776_
timestamp 1608254825
transform 1 0 26772 0 -1 8160
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_10_319
timestamp 1608254825
transform 1 0 30452 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2607_
timestamp 1608254825
transform 1 0 28704 0 -1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_10_341
timestamp 1608254825
transform 1 0 32476 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_10_332
timestamp 1608254825
transform 1 0 31648 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_206
timestamp 1608254825
transform 1 0 32016 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1456_
timestamp 1608254825
transform 1 0 32108 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__and4_4  _1436_
timestamp 1608254825
transform 1 0 30820 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_10_362
timestamp 1608254825
transform 1 0 34408 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_4  _1498_
timestamp 1608254825
transform 1 0 33212 0 -1 8160
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_8  FILLER_10_386
timestamp 1608254825
transform 1 0 36616 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_10_379
timestamp 1608254825
transform 1 0 35972 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_4  _1515_
timestamp 1608254825
transform 1 0 34776 0 -1 8160
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _1512_
timestamp 1608254825
transform 1 0 36340 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_406
timestamp 1608254825
transform 1 0 38456 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_398
timestamp 1608254825
transform 1 0 37720 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_394
timestamp 1608254825
transform 1 0 37352 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_207
timestamp 1608254825
transform 1 0 37628 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1608254825
transform -1 0 38824 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_11
timestamp 1608254825
transform 1 0 2116 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_3
timestamp 1608254825
transform 1 0 1380 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1608254825
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__and2_4  _1916_
timestamp 1608254825
transform 1 0 1472 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_4  _1907_
timestamp 1608254825
transform 1 0 2484 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_11_32
timestamp 1608254825
transform 1 0 4048 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_28
timestamp 1608254825
transform 1 0 3680 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_24
timestamp 1608254825
transform 1 0 3312 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2428_
timestamp 1608254825
transform 1 0 4416 0 1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_2  _1906_
timestamp 1608254825
transform 1 0 3772 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_11_55
timestamp 1608254825
transform 1 0 6164 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_208
timestamp 1608254825
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_4  _2199_
timestamp 1608254825
transform 1 0 6808 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_11_77
timestamp 1608254825
transform 1 0 8188 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_71
timestamp 1608254825
transform 1 0 7636 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_addressalyzerBlock.SPI_CLK
timestamp 1608254825
transform 1 0 8280 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _2425_
timestamp 1608254825
transform 1 0 8556 0 1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_11_108
timestamp 1608254825
transform 1 0 11040 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_100
timestamp 1608254825
transform 1 0 10304 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_4  _1845_
timestamp 1608254825
transform 1 0 11132 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_11_135
timestamp 1608254825
transform 1 0 13524 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_118
timestamp 1608254825
transform 1 0 11960 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_209
timestamp 1608254825
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__a21o_4  _1629_
timestamp 1608254825
transform 1 0 12420 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_159
timestamp 1608254825
transform 1 0 15732 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_142
timestamp 1608254825
transform 1 0 14168 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_4  _1853_
timestamp 1608254825
transform 1 0 14536 0 1 8160
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _1617_
timestamp 1608254825
transform 1 0 13892 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_179
timestamp 1608254825
transform 1 0 17572 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_172
timestamp 1608254825
transform 1 0 16928 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_4  _2196_
timestamp 1608254825
transform 1 0 16100 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1927_
timestamp 1608254825
transform 1 0 17296 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_196
timestamp 1608254825
transform 1 0 19136 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_11_184
timestamp 1608254825
transform 1 0 18032 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_210
timestamp 1608254825
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__a211o_4  _1752_
timestamp 1608254825
transform 1 0 19504 0 1 8160
box -38 -48 1326 592
use sky130_fd_sc_hd__nor2_4  _1637_
timestamp 1608254825
transform 1 0 18308 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_11_222
timestamp 1608254825
transform 1 0 21528 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_214
timestamp 1608254825
transform 1 0 20792 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_4  _2320_
timestamp 1608254825
transform 1 0 21712 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_11_249
timestamp 1608254825
transform 1 0 24012 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_245
timestamp 1608254825
transform 1 0 23644 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_240
timestamp 1608254825
transform 1 0 23184 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_211
timestamp 1608254825
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2396_
timestamp 1608254825
transform 1 0 24104 0 1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_11_269
timestamp 1608254825
transform 1 0 25852 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_11_291
timestamp 1608254825
transform 1 0 27876 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_4  _1772_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 26588 0 1 8160
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_3  FILLER_11_306
timestamp 1608254825
transform 1 0 29256 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_301
timestamp 1608254825
transform 1 0 28796 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_212
timestamp 1608254825
transform 1 0 29164 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__a21o_4  _1513_
timestamp 1608254825
transform 1 0 29532 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _1481_
timestamp 1608254825
transform 1 0 28428 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_338
timestamp 1608254825
transform 1 0 32200 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_321
timestamp 1608254825
transform 1 0 30636 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_4  _1517_
timestamp 1608254825
transform 1 0 31004 0 1 8160
box -38 -48 1234 592
use sky130_fd_sc_hd__a21oi_4  _1480_
timestamp 1608254825
transform 1 0 32568 0 1 8160
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_11_362
timestamp 1608254825
transform 1 0 34408 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_355
timestamp 1608254825
transform 1 0 33764 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1511_
timestamp 1608254825
transform 1 0 34132 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_380
timestamp 1608254825
transform 1 0 36064 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_367
timestamp 1608254825
transform 1 0 34868 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_213
timestamp 1608254825
transform 1 0 34776 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2572_
timestamp 1608254825
transform 1 0 36432 0 1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__o21a_4  _1804_
timestamp 1608254825
transform 1 0 34960 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_403
timestamp 1608254825
transform 1 0 38180 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1608254825
transform -1 0 38824 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_12_7
timestamp 1608254825
transform 1 0 1748 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_3
timestamp 1608254825
transform 1 0 1380 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1608254825
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _2540_
timestamp 1608254825
transform 1 0 1840 0 -1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_12_43
timestamp 1608254825
transform 1 0 5060 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_32
timestamp 1608254825
transform 1 0 4048 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_12_27
timestamp 1608254825
transform 1 0 3588 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_214
timestamp 1608254825
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1623_
timestamp 1608254825
transform 1 0 4784 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__o32ai_4  _2259_
timestamp 1608254825
transform 1 0 5428 0 -1 9248
box -38 -48 2062 592
use sky130_fd_sc_hd__decap_4  FILLER_12_88
timestamp 1608254825
transform 1 0 9200 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_78
timestamp 1608254825
transform 1 0 8280 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_69
timestamp 1608254825
transform 1 0 7452 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_1_0_addressalyzerBlock.SPI_CLK
timestamp 1608254825
transform 1 0 8004 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_4  _2151_
timestamp 1608254825
transform 1 0 8372 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_12_110
timestamp 1608254825
transform 1 0 11224 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_12_93
timestamp 1608254825
transform 1 0 9660 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_215
timestamp 1608254825
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _1938_
timestamp 1608254825
transform 1 0 11592 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_4  _1711_
timestamp 1608254825
transform 1 0 9936 0 -1 9248
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_1  FILLER_12_127
timestamp 1608254825
transform 1 0 12788 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_123
timestamp 1608254825
transform 1 0 12420 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_4  _1621_
timestamp 1608254825
transform 1 0 12880 0 -1 9248
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_12_149
timestamp 1608254825
transform 1 0 14812 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_142
timestamp 1608254825
transform 1 0 14168 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_216
timestamp 1608254825
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1937_
timestamp 1608254825
transform 1 0 14536 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_4  _1639_
timestamp 1608254825
transform 1 0 15272 0 -1 9248
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_6  FILLER_12_175
timestamp 1608254825
transform 1 0 17204 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_167
timestamp 1608254825
transform 1 0 16468 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_4  _2181_
timestamp 1608254825
transform 1 0 17756 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _1616_
timestamp 1608254825
transform 1 0 16836 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_190
timestamp 1608254825
transform 1 0 18584 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_4  _1638_
timestamp 1608254825
transform 1 0 19136 0 -1 9248
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_12_228
timestamp 1608254825
transform 1 0 22080 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_210
timestamp 1608254825
transform 1 0 20424 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_217
timestamp 1608254825
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_4  _2126_
timestamp 1608254825
transform 1 0 20884 0 -1 9248
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_12_236
timestamp 1608254825
transform 1 0 22816 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2397_
timestamp 1608254825
transform 1 0 23184 0 -1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  _2313_
timestamp 1608254825
transform 1 0 22448 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_271
timestamp 1608254825
transform 1 0 26036 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_259
timestamp 1608254825
transform 1 0 24932 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1486_
timestamp 1608254825
transform 1 0 25668 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_295
timestamp 1608254825
transform 1 0 28244 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_276
timestamp 1608254825
transform 1 0 26496 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_218
timestamp 1608254825
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_4  _1496_
timestamp 1608254825
transform 1 0 27048 0 -1 9248
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_12_316
timestamp 1608254825
transform 1 0 30176 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__nand4_4  _1487_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 28612 0 -1 9248
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_12_340
timestamp 1608254825
transform 1 0 32384 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_332
timestamp 1608254825
transform 1 0 31648 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_219
timestamp 1608254825
transform 1 0 32016 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_4  _1825_
timestamp 1608254825
transform 1 0 30544 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1504_
timestamp 1608254825
transform 1 0 32108 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_363
timestamp 1608254825
transform 1 0 34500 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _2610_
timestamp 1608254825
transform 1 0 32752 0 -1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_12_384
timestamp 1608254825
transform 1 0 36432 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_371
timestamp 1608254825
transform 1 0 35236 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_4  _1805_
timestamp 1608254825
transform 1 0 35328 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _1799_
timestamp 1608254825
transform 1 0 36800 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_406
timestamp 1608254825
transform 1 0 38456 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_398
timestamp 1608254825
transform 1 0 37720 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_396
timestamp 1608254825
transform 1 0 37536 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_392
timestamp 1608254825
transform 1 0 37168 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_220
timestamp 1608254825
transform 1 0 37628 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1608254825
transform -1 0 38824 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_3
timestamp 1608254825
transform 1 0 1380 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_22
timestamp 1608254825
transform 1 0 3128 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1608254825
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1608254825
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _2538_
timestamp 1608254825
transform 1 0 1748 0 -1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _2536_
timestamp 1608254825
transform 1 0 1380 0 1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_14_32
timestamp 1608254825
transform 1 0 4048 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_30
timestamp 1608254825
transform 1 0 3864 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_26
timestamp 1608254825
transform 1 0 3496 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_227
timestamp 1608254825
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _1911_
timestamp 1608254825
transform 1 0 3496 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_14_41
timestamp 1608254825
transform 1 0 4876 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_35
timestamp 1608254825
transform 1 0 4324 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__and2_4  _1918_
timestamp 1608254825
transform 1 0 4232 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1910_
timestamp 1608254825
transform 1 0 4876 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_44
timestamp 1608254825
transform 1 0 5152 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_0_0_m1_clk_local
timestamp 1608254825
transform 1 0 5244 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_67
timestamp 1608254825
transform 1 0 7268 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_57
timestamp 1608254825
transform 1 0 6348 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_221
timestamp 1608254825
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2519_
timestamp 1608254825
transform 1 0 5520 0 -1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__nor2_4  _1942_
timestamp 1608254825
transform 1 0 6808 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_4  _1940_
timestamp 1608254825
transform 1 0 5520 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_14_85
timestamp 1608254825
transform 1 0 8924 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_71
timestamp 1608254825
transform 1 0 7636 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_71
timestamp 1608254825
transform 1 0 7636 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_2_0_m1_clk_local
timestamp 1608254825
transform 1 0 9292 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__o32ai_4  _2267_
timestamp 1608254825
transform 1 0 8004 0 1 9248
box -38 -48 2062 592
use sky130_fd_sc_hd__a21oi_4  _1747_
timestamp 1608254825
transform 1 0 7728 0 -1 10336
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_8  FILLER_14_105
timestamp 1608254825
transform 1 0 10764 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_105
timestamp 1608254825
transform 1 0 10764 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_97
timestamp 1608254825
transform 1 0 10028 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_228
timestamp 1608254825
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__a21o_4  _1850_
timestamp 1608254825
transform 1 0 10856 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__a211o_4  _1846_
timestamp 1608254825
transform 1 0 11500 0 -1 10336
box -38 -48 1326 592
use sky130_fd_sc_hd__a21o_4  _1749_
timestamp 1608254825
transform 1 0 9660 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_127
timestamp 1608254825
transform 1 0 12788 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_123
timestamp 1608254825
transform 1 0 12420 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_118
timestamp 1608254825
transform 1 0 11960 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_222
timestamp 1608254825
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__a21o_4  _2222_
timestamp 1608254825
transform 1 0 13156 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__a21oi_4  _2218_
timestamp 1608254825
transform 1 0 12788 0 1 9248
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_14_154
timestamp 1608254825
transform 1 0 15272 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_151
timestamp 1608254825
transform 1 0 14996 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_143
timestamp 1608254825
transform 1 0 14260 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_140
timestamp 1608254825
transform 1 0 13984 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_229
timestamp 1608254825
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2521_
timestamp 1608254825
transform 1 0 14352 0 1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__and2_4  _1952_
timestamp 1608254825
transform 1 0 15640 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_14_165
timestamp 1608254825
transform 1 0 16284 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_179
timestamp 1608254825
transform 1 0 17572 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_169
timestamp 1608254825
transform 1 0 16652 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_163
timestamp 1608254825
transform 1 0 16100 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_4  _2225_
timestamp 1608254825
transform 1 0 16652 0 -1 10336
box -38 -48 1326 592
use sky130_fd_sc_hd__nor2_4  _2203_
timestamp 1608254825
transform 1 0 16744 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_14_183
timestamp 1608254825
transform 1 0 17940 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_188
timestamp 1608254825
transform 1 0 18400 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_223
timestamp 1608254825
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _1851_
timestamp 1608254825
transform 1 0 18768 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _1630_
timestamp 1608254825
transform 1 0 18032 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_201
timestamp 1608254825
transform 1 0 19596 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_201
timestamp 1608254825
transform 1 0 19596 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2144_
timestamp 1608254825
transform 1 0 19964 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1633_
timestamp 1608254825
transform 1 0 19964 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_4  _1715_
timestamp 1608254825
transform 1 0 18308 0 -1 10336
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_1  FILLER_14_213
timestamp 1608254825
transform 1 0 20700 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_209
timestamp 1608254825
transform 1 0 20332 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_208
timestamp 1608254825
transform 1 0 20240 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_230
timestamp 1608254825
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2446_
timestamp 1608254825
transform 1 0 20608 0 1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__nand3_4  _2125_
timestamp 1608254825
transform 1 0 20884 0 -1 10336
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_1  FILLER_14_237
timestamp 1608254825
transform 1 0 22908 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_229
timestamp 1608254825
transform 1 0 22172 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_239
timestamp 1608254825
transform 1 0 23092 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_231
timestamp 1608254825
transform 1 0 22356 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _2124_
timestamp 1608254825
transform 1 0 22724 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_251
timestamp 1608254825
transform 1 0 24196 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_13_245
timestamp 1608254825
transform 1 0 23644 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_13_243
timestamp 1608254825
transform 1 0 23460 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_224
timestamp 1608254825
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1764_
timestamp 1608254825
transform 1 0 23920 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _2395_
timestamp 1608254825
transform 1 0 23000 0 -1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_14_271
timestamp 1608254825
transform 1 0 26036 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_261
timestamp 1608254825
transform 1 0 25116 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_257
timestamp 1608254825
transform 1 0 24748 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_4  _1768_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 24564 0 1 9248
box -38 -48 2062 592
use sky130_fd_sc_hd__nor2_4  _1766_
timestamp 1608254825
transform 1 0 25208 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_14_282
timestamp 1608254825
transform 1 0 27048 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_276
timestamp 1608254825
transform 1 0 26496 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_277
timestamp 1608254825
transform 1 0 26588 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_231
timestamp 1608254825
transform 1 0 26404 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__a2111o_4  _1769_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 26956 0 1 9248
box -38 -48 1602 592
use sky130_fd_sc_hd__a41oi_4  _1495_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 27416 0 -1 10336
box -38 -48 2062 592
use sky130_fd_sc_hd__buf_2  _1437_
timestamp 1608254825
transform 1 0 26680 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_308
timestamp 1608254825
transform 1 0 29440 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_306
timestamp 1608254825
transform 1 0 29256 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_304
timestamp 1608254825
transform 1 0 29072 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_298
timestamp 1608254825
transform 1 0 28520 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_225
timestamp 1608254825
transform 1 0 29164 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1470_
timestamp 1608254825
transform 1 0 29348 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_315
timestamp 1608254825
transform 1 0 30084 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_311
timestamp 1608254825
transform 1 0 29716 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_8_0_addressalyzerBlock.SPI_CLK
timestamp 1608254825
transform 1 0 29808 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_4  _1476_
timestamp 1608254825
transform 1 0 30268 0 -1 10336
box -38 -48 1234 592
use sky130_fd_sc_hd__a41oi_4  _1475_
timestamp 1608254825
transform 1 0 30084 0 1 9248
box -38 -48 2062 592
use sky130_fd_sc_hd__fill_1  FILLER_14_341
timestamp 1608254825
transform 1 0 32476 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_337
timestamp 1608254825
transform 1 0 32108 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_330
timestamp 1608254825
transform 1 0 31464 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_337
timestamp 1608254825
transform 1 0 32108 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_232
timestamp 1608254825
transform 1 0 32016 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_4  _1479_
timestamp 1608254825
transform 1 0 32476 0 1 9248
box -38 -48 1234 592
use sky130_fd_sc_hd__o21ai_4  _1464_
timestamp 1608254825
transform 1 0 32568 0 -1 10336
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_14_355
timestamp 1608254825
transform 1 0 33764 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_362
timestamp 1608254825
transform 1 0 34408 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_354
timestamp 1608254825
transform 1 0 33672 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_10_0_addressalyzerBlock.SPI_CLK
timestamp 1608254825
transform 1 0 34132 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _2611_
timestamp 1608254825
transform 1 0 34408 0 -1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  _1461_
timestamp 1608254825
transform 1 0 34040 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_381
timestamp 1608254825
transform 1 0 36156 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_380
timestamp 1608254825
transform 1 0 36064 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_367
timestamp 1608254825
transform 1 0 34868 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_226
timestamp 1608254825
transform 1 0 34776 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2591_
timestamp 1608254825
transform 1 0 36432 0 1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__o21a_4  _1806_
timestamp 1608254825
transform 1 0 34960 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _1520_
timestamp 1608254825
transform 1 0 36524 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_401
timestamp 1608254825
transform 1 0 37996 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_14_389
timestamp 1608254825
transform 1 0 36892 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_403
timestamp 1608254825
transform 1 0 38180 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_233
timestamp 1608254825
transform 1 0 37628 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1608254825
transform -1 0 38824 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1608254825
transform -1 0 38824 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1770_
timestamp 1608254825
transform 1 0 37720 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_15_15
timestamp 1608254825
transform 1 0 2484 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_15_3
timestamp 1608254825
transform 1 0 1380 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1608254825
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__and2_4  _1920_
timestamp 1608254825
transform 1 0 3036 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _1901_
timestamp 1608254825
transform 1 0 2116 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_28
timestamp 1608254825
transform 1 0 3680 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_4  _2156_
timestamp 1608254825
transform 1 0 4048 0 1 10336
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_1  FILLER_15_68
timestamp 1608254825
transform 1 0 7360 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_62
timestamp 1608254825
transform 1 0 6808 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_57
timestamp 1608254825
transform 1 0 6348 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_46
timestamp 1608254825
transform 1 0 5336 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_234
timestamp 1608254825
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _1954_
timestamp 1608254825
transform 1 0 5704 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_15_86
timestamp 1608254825
transform 1 0 9016 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_82
timestamp 1608254825
transform 1 0 8648 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_4  _1748_
timestamp 1608254825
transform 1 0 7452 0 1 10336
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_4  _1712_
timestamp 1608254825
transform 1 0 9108 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_15_114
timestamp 1608254825
transform 1 0 11592 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_15_96
timestamp 1608254825
transform 1 0 9936 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_4  _1707_
timestamp 1608254825
transform 1 0 10304 0 1 10336
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_6  FILLER_15_136
timestamp 1608254825
transform 1 0 13616 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_235
timestamp 1608254825
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_4  _2219_
timestamp 1608254825
transform 1 0 12420 0 1 10336
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_15_154
timestamp 1608254825
transform 1 0 15272 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_4  _1753_
timestamp 1608254825
transform 1 0 14168 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _1634_
timestamp 1608254825
transform 1 0 15640 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_179
timestamp 1608254825
transform 1 0 17572 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_162
timestamp 1608254825
transform 1 0 16008 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_4  _1717_
timestamp 1608254825
transform 1 0 16376 0 1 10336
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_6  FILLER_15_193
timestamp 1608254825
transform 1 0 18860 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_236
timestamp 1608254825
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _2158_
timestamp 1608254825
transform 1 0 19412 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  _1716_
timestamp 1608254825
transform 1 0 18032 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_15_220
timestamp 1608254825
transform 1 0 21344 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_216
timestamp 1608254825
transform 1 0 20976 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_208
timestamp 1608254825
transform 1 0 20240 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_4  _2321_
timestamp 1608254825
transform 1 0 21712 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  _1771_
timestamp 1608254825
transform 1 0 21068 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_248
timestamp 1608254825
transform 1 0 23920 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_240
timestamp 1608254825
transform 1 0 23184 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_237
timestamp 1608254825
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1503_
timestamp 1608254825
transform 1 0 23644 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_274
timestamp 1608254825
transform 1 0 26312 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_4  _1767_
timestamp 1608254825
transform 1 0 24288 0 1 10336
box -38 -48 2062 592
use sky130_fd_sc_hd__decap_4  FILLER_15_288
timestamp 1608254825
transform 1 0 27600 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_278
timestamp 1608254825
transform 1 0 26680 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__and4_4  _1494_
timestamp 1608254825
transform 1 0 26772 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__and4_4  _1473_
timestamp 1608254825
transform 1 0 27968 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_15_319
timestamp 1608254825
transform 1 0 30452 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_306
timestamp 1608254825
transform 1 0 29256 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_301
timestamp 1608254825
transform 1 0 28796 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_238
timestamp 1608254825
transform 1 0 29164 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__a21o_4  _1509_
timestamp 1608254825
transform 1 0 29348 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_329
timestamp 1608254825
transform 1 0 31372 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_4  _1827_
timestamp 1608254825
transform 1 0 31740 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _1439_
timestamp 1608254825
transform 1 0 31004 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_362
timestamp 1608254825
transform 1 0 34408 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_345
timestamp 1608254825
transform 1 0 32844 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_4  _1458_
timestamp 1608254825
transform 1 0 33212 0 1 10336
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_15_380
timestamp 1608254825
transform 1 0 36064 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_239
timestamp 1608254825
transform 1 0 34776 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2502_
timestamp 1608254825
transform 1 0 36432 0 1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__a21oi_4  _1465_
timestamp 1608254825
transform 1 0 34868 0 1 10336
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_15_403
timestamp 1608254825
transform 1 0 38180 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1608254825
transform -1 0 38824 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_20
timestamp 1608254825
transform 1 0 2944 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_11
timestamp 1608254825
transform 1 0 2116 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_3
timestamp 1608254825
transform 1 0 1380 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1608254825
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__and2_4  _1957_
timestamp 1608254825
transform 1 0 2300 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_16_41
timestamp 1608254825
transform 1 0 4876 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_16_28
timestamp 1608254825
transform 1 0 3680 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_m1_clk_local
timestamp 1608254825
transform 1 0 5244 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_240
timestamp 1608254825
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_4  _2155_
timestamp 1608254825
transform 1 0 4048 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_16_62
timestamp 1608254825
transform 1 0 6808 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _2262_
timestamp 1608254825
transform 1 0 7360 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_4  _2201_
timestamp 1608254825
transform 1 0 5520 0 -1 11424
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_16_88
timestamp 1608254825
transform 1 0 9200 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_72
timestamp 1608254825
transform 1 0 7728 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_4  _2157_
timestamp 1608254825
transform 1 0 8096 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_110
timestamp 1608254825
transform 1 0 11224 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_93
timestamp 1608254825
transform 1 0 9660 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_241
timestamp 1608254825
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__a211o_4  _1745_
timestamp 1608254825
transform 1 0 9936 0 -1 11424
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_16_133
timestamp 1608254825
transform 1 0 13340 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_118
timestamp 1608254825
transform 1 0 11960 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__o21ai_4  _2221_
timestamp 1608254825
transform 1 0 12144 0 -1 11424
box -38 -48 1234 592
use sky130_fd_sc_hd__a21o_4  _2180_
timestamp 1608254825
transform 1 0 13708 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_154
timestamp 1608254825
transform 1 0 15272 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_149
timestamp 1608254825
transform 1 0 14812 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_242
timestamp 1608254825
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_4  _2226_
timestamp 1608254825
transform 1 0 15364 0 -1 11424
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_16_177
timestamp 1608254825
transform 1 0 17388 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_172
timestamp 1608254825
transform 1 0 16928 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_168
timestamp 1608254825
transform 1 0 16560 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_4  _2182_
timestamp 1608254825
transform 1 0 17756 0 -1 11424
box -38 -48 1326 592
use sky130_fd_sc_hd__buf_2  _1635_
timestamp 1608254825
transform 1 0 17020 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_195
timestamp 1608254825
transform 1 0 19044 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_4  _2224_
timestamp 1608254825
transform 1 0 19412 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_16_228
timestamp 1608254825
transform 1 0 22080 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_221
timestamp 1608254825
transform 1 0 21436 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_16_215
timestamp 1608254825
transform 1 0 20884 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_16_208
timestamp 1608254825
transform 1 0 20240 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_243
timestamp 1608254825
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1533_
timestamp 1608254825
transform 1 0 21160 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1420_
timestamp 1608254825
transform 1 0 21804 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_246
timestamp 1608254825
transform 1 0 23736 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_236
timestamp 1608254825
transform 1 0 22816 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_11_0_m1_clk_local
timestamp 1608254825
transform 1 0 24104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1472_
timestamp 1608254825
transform 1 0 23368 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1471_
timestamp 1608254825
transform 1 0 22448 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_274
timestamp 1608254825
transform 1 0 26312 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_268
timestamp 1608254825
transform 1 0 25760 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_260
timestamp 1608254825
transform 1 0 25024 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_16_253
timestamp 1608254825
transform 1 0 24380 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1484_
timestamp 1608254825
transform 1 0 24656 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1431_
timestamp 1608254825
transform 1 0 25392 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_295
timestamp 1608254825
transform 1 0 28244 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_244
timestamp 1608254825
transform 1 0 26404 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2605_
timestamp 1608254825
transform 1 0 26496 0 -1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_16_316
timestamp 1608254825
transform 1 0 30176 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__nand4_4  _1505_
timestamp 1608254825
transform 1 0 28612 0 -1 11424
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_16_332
timestamp 1608254825
transform 1 0 31648 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_245
timestamp 1608254825
transform 1 0 32016 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_4  _1828_
timestamp 1608254825
transform 1 0 30544 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__a21oi_4  _1523_
timestamp 1608254825
transform 1 0 32108 0 -1 11424
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_6  FILLER_16_350
timestamp 1608254825
transform 1 0 33304 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_4  _1463_
timestamp 1608254825
transform 1 0 33856 0 -1 11424
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_16_369
timestamp 1608254825
transform 1 0 35052 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2580_
timestamp 1608254825
transform 1 0 35420 0 -1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_16_406
timestamp 1608254825
transform 1 0 38456 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_398
timestamp 1608254825
transform 1 0 37720 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_396
timestamp 1608254825
transform 1 0 37536 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_392
timestamp 1608254825
transform 1 0 37168 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_246
timestamp 1608254825
transform 1 0 37628 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1608254825
transform -1 0 38824 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_13
timestamp 1608254825
transform 1 0 2300 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_3
timestamp 1608254825
transform 1 0 1380 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1608254825
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _2422_
timestamp 1608254825
transform 1 0 2668 0 1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__nor2_4  _1945_
timestamp 1608254825
transform 1 0 1472 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_17_36
timestamp 1608254825
transform 1 0 4416 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_4  _2179_
timestamp 1608254825
transform 1 0 4784 0 1 11424
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_1  FILLER_17_60
timestamp 1608254825
transform 1 0 6624 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_54
timestamp 1608254825
transform 1 0 6072 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_247
timestamp 1608254825
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_4  _2200_
timestamp 1608254825
transform 1 0 6808 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_17_75
timestamp 1608254825
transform 1 0 8004 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_71
timestamp 1608254825
transform 1 0 7636 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_m1_clk_local
timestamp 1608254825
transform 1 0 8096 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_4  _2153_
timestamp 1608254825
transform 1 0 8372 0 1 11424
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_17_110
timestamp 1608254825
transform 1 0 11224 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_93
timestamp 1608254825
transform 1 0 9660 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_4  _2296_
timestamp 1608254825
transform 1 0 10028 0 1 11424
box -38 -48 1234 592
use sky130_fd_sc_hd__buf_2  _1628_
timestamp 1608254825
transform 1 0 11592 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_136
timestamp 1608254825
transform 1 0 13616 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_123
timestamp 1608254825
transform 1 0 12420 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_118
timestamp 1608254825
transform 1 0 11960 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_248
timestamp 1608254825
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__a21o_4  _2202_
timestamp 1608254825
transform 1 0 12512 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_156
timestamp 1608254825
transform 1 0 15456 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__nand3_4  _2176_
timestamp 1608254825
transform 1 0 14168 0 1 11424
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_1  FILLER_17_182
timestamp 1608254825
transform 1 0 17848 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_178
timestamp 1608254825
transform 1 0 17480 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_164
timestamp 1608254825
transform 1 0 16192 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_4  _2160_
timestamp 1608254825
transform 1 0 16284 0 1 11424
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_1  FILLER_17_199
timestamp 1608254825
transform 1 0 19412 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_195
timestamp 1608254825
transform 1 0 19044 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_188
timestamp 1608254825
transform 1 0 18400 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_249
timestamp 1608254825
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2442_
timestamp 1608254825
transform 1 0 19504 0 1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  _1703_
timestamp 1608254825
transform 1 0 18032 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1632_
timestamp 1608254825
transform 1 0 18768 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_17_219
timestamp 1608254825
transform 1 0 21252 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__and2_4  _1968_
timestamp 1608254825
transform 1 0 21988 0 1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_17_245
timestamp 1608254825
transform 1 0 23644 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_242
timestamp 1608254825
transform 1 0 23368 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_234
timestamp 1608254825
transform 1 0 22632 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_250
timestamp 1608254825
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _1607_
timestamp 1608254825
transform 1 0 23828 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_17_271
timestamp 1608254825
transform 1 0 26036 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_256
timestamp 1608254825
transform 1 0 24656 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__and4_4  _1483_
timestamp 1608254825
transform 1 0 25208 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__a41oi_4  _1518_
timestamp 1608254825
transform 1 0 26404 0 1 11424
box -38 -48 2062 592
use sky130_fd_sc_hd__fill_1  FILLER_17_301
timestamp 1608254825
transform 1 0 28796 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_297
timestamp 1608254825
transform 1 0 28428 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_addressalyzerBlock.SPI_CLK
timestamp 1608254825
transform 1 0 28888 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_251
timestamp 1608254825
transform 1 0 29164 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__a41o_4  _1508_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 29256 0 1 11424
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_17_340
timestamp 1608254825
transform 1 0 32384 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_323
timestamp 1608254825
transform 1 0 30820 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_4  _1519_
timestamp 1608254825
transform 1 0 31188 0 1 11424
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_8  FILLER_17_358
timestamp 1608254825
transform 1 0 34040 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_344
timestamp 1608254825
transform 1 0 32752 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_4  _1452_
timestamp 1608254825
transform 1 0 32844 0 1 11424
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_17_380
timestamp 1608254825
transform 1 0 36064 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_252
timestamp 1608254825
transform 1 0 34776 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2513_
timestamp 1608254825
transform 1 0 36432 0 1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__a21oi_4  _1521_
timestamp 1608254825
transform 1 0 34868 0 1 11424
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_17_403
timestamp 1608254825
transform 1 0 38180 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1608254825
transform -1 0 38824 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_18_22
timestamp 1608254825
transform 1 0 3128 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1608254825
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _2517_
timestamp 1608254825
transform 1 0 1380 0 -1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_18_41
timestamp 1608254825
transform 1 0 4876 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_30
timestamp 1608254825
transform 1 0 3864 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_253
timestamp 1608254825
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_4  _2178_
timestamp 1608254825
transform 1 0 4048 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1941_
timestamp 1608254825
transform 1 0 5244 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_48
timestamp 1608254825
transform 1 0 5520 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__o32ai_4  _2272_
timestamp 1608254825
transform 1 0 5888 0 -1 12512
box -38 -48 2062 592
use sky130_fd_sc_hd__fill_1  FILLER_18_91
timestamp 1608254825
transform 1 0 9476 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_87
timestamp 1608254825
transform 1 0 9108 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_74
timestamp 1608254825
transform 1 0 7912 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_4  _2152_
timestamp 1608254825
transform 1 0 8280 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_18_93
timestamp 1608254825
transform 1 0 9660 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_254
timestamp 1608254825
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2409_
timestamp 1608254825
transform 1 0 9936 0 -1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_18_122
timestamp 1608254825
transform 1 0 12328 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_115
timestamp 1608254825
transform 1 0 11684 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2268_
timestamp 1608254825
transform 1 0 12052 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_4  _2198_
timestamp 1608254825
transform 1 0 12696 0 -1 12512
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_2  FILLER_18_154
timestamp 1608254825
transform 1 0 15272 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_152
timestamp 1608254825
transform 1 0 15088 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_148
timestamp 1608254825
transform 1 0 14720 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_140
timestamp 1608254825
transform 1 0 13984 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_255
timestamp 1608254825
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_4  _2205_
timestamp 1608254825
transform 1 0 15456 0 -1 12512
box -38 -48 1234 592
use sky130_fd_sc_hd__buf_2  _1708_
timestamp 1608254825
transform 1 0 14352 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_169
timestamp 1608254825
transform 1 0 16652 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_4  _2204_
timestamp 1608254825
transform 1 0 17020 0 -1 12512
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_8  FILLER_18_205
timestamp 1608254825
transform 1 0 19964 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_18_187
timestamp 1608254825
transform 1 0 18308 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_4  _2159_
timestamp 1608254825
transform 1 0 18676 0 -1 12512
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_1  FILLER_18_213
timestamp 1608254825
transform 1 0 20700 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_256
timestamp 1608254825
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2506_
timestamp 1608254825
transform 1 0 20884 0 -1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_18_242
timestamp 1608254825
transform 1 0 23368 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_234
timestamp 1608254825
transform 1 0 22632 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2603_
timestamp 1608254825
transform 1 0 23736 0 -1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  _1430_
timestamp 1608254825
transform 1 0 23000 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_273
timestamp 1608254825
transform 1 0 26220 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_265
timestamp 1608254825
transform 1 0 25484 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_18_291
timestamp 1608254825
transform 1 0 27876 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_276
timestamp 1608254825
transform 1 0 26496 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_257
timestamp 1608254825
transform 1 0 26404 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_4  _1506_
timestamp 1608254825
transform 1 0 28244 0 -1 12512
box -38 -48 1234 592
use sky130_fd_sc_hd__and4_4  _1432_
timestamp 1608254825
transform 1 0 27048 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_18_315
timestamp 1608254825
transform 1 0 30084 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_308
timestamp 1608254825
transform 1 0 29440 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_4  _1522_
timestamp 1608254825
transform 1 0 30452 0 -1 12512
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _1447_
timestamp 1608254825
transform 1 0 29808 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_332
timestamp 1608254825
transform 1 0 31648 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_258
timestamp 1608254825
transform 1 0 32016 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__and4_4  _1438_
timestamp 1608254825
transform 1 0 32108 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_18_364
timestamp 1608254825
transform 1 0 34592 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_350
timestamp 1608254825
transform 1 0 33304 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_346
timestamp 1608254825
transform 1 0 32936 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_4  _1453_
timestamp 1608254825
transform 1 0 33396 0 -1 12512
box -38 -48 1234 592
use sky130_fd_sc_hd__dfxtp_4  _2581_
timestamp 1608254825
transform 1 0 35144 0 -1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_18_401
timestamp 1608254825
transform 1 0 37996 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_18_389
timestamp 1608254825
transform 1 0 36892 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_259
timestamp 1608254825
transform 1 0 37628 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1608254825
transform -1 0 38824 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2142_
timestamp 1608254825
transform 1 0 37720 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_22
timestamp 1608254825
transform 1 0 3128 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_14
timestamp 1608254825
transform 1 0 2392 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_3
timestamp 1608254825
transform 1 0 1380 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_3
timestamp 1608254825
transform 1 0 1380 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1608254825
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1608254825
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _2421_
timestamp 1608254825
transform 1 0 1656 0 1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__nor2_4  _1949_
timestamp 1608254825
transform 1 0 1564 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_20_42
timestamp 1608254825
transform 1 0 4968 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_35
timestamp 1608254825
transform 1 0 4324 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_27
timestamp 1608254825
transform 1 0 3588 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_25
timestamp 1608254825
transform 1 0 3404 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_266
timestamp 1608254825
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__o32ai_4  _2273_
timestamp 1608254825
transform 1 0 3772 0 1 12512
box -38 -48 2062 592
use sky130_fd_sc_hd__inv_2  _1948_
timestamp 1608254825
transform 1 0 3312 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1944_
timestamp 1608254825
transform 1 0 4048 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1746_
timestamp 1608254825
transform 1 0 4692 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_50
timestamp 1608254825
transform 1 0 5704 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_57
timestamp 1608254825
transform 1 0 6348 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_51
timestamp 1608254825
transform 1 0 5796 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_m1_clk_local
timestamp 1608254825
transform 1 0 6440 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_260
timestamp 1608254825
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2423_
timestamp 1608254825
transform 1 0 6072 0 -1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__o32ai_4  _2271_
timestamp 1608254825
transform 1 0 6808 0 1 12512
box -38 -48 2062 592
use sky130_fd_sc_hd__buf_2  _2264_
timestamp 1608254825
transform 1 0 5336 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_86
timestamp 1608254825
transform 1 0 9016 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_81
timestamp 1608254825
transform 1 0 8556 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_73
timestamp 1608254825
transform 1 0 7820 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_84
timestamp 1608254825
transform 1 0 8832 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_4  _2197_
timestamp 1608254825
transform 1 0 9200 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _1618_
timestamp 1608254825
transform 1 0 8648 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_112
timestamp 1608254825
transform 1 0 11408 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_97
timestamp 1608254825
transform 1 0 10028 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_3_0_m1_clk_local
timestamp 1608254825
transform 1 0 10396 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_267
timestamp 1608254825
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2407_
timestamp 1608254825
transform 1 0 9660 0 -1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__nand3_4  _2295_
timestamp 1608254825
transform 1 0 10672 0 1 12512
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_2  FILLER_19_123
timestamp 1608254825
transform 1 0 12420 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_118
timestamp 1608254825
transform 1 0 11960 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_261
timestamp 1608254825
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2410_
timestamp 1608254825
transform 1 0 12144 0 -1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__nand3_4  _2293_
timestamp 1608254825
transform 1 0 12604 0 1 12512
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_20_149
timestamp 1608254825
transform 1 0 14812 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_139
timestamp 1608254825
transform 1 0 13892 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_139
timestamp 1608254825
transform 1 0 13892 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_addressalyzerBlock.SPI_CLK
timestamp 1608254825
transform 1 0 14260 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_268
timestamp 1608254825
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _2266_
timestamp 1608254825
transform 1 0 14536 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_4  _2241_
timestamp 1608254825
transform 1 0 14628 0 1 12512
box -38 -48 1326 592
use sky130_fd_sc_hd__nand2_4  _2175_
timestamp 1608254825
transform 1 0 15272 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_20_167
timestamp 1608254825
transform 1 0 16468 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_163
timestamp 1608254825
transform 1 0 16100 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_179
timestamp 1608254825
transform 1 0 17572 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_165
timestamp 1608254825
transform 1 0 16284 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_161
timestamp 1608254825
transform 1 0 15916 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_4  _2183_
timestamp 1608254825
transform 1 0 16376 0 1 12512
box -38 -48 1234 592
use sky130_fd_sc_hd__o32ai_4  _2143_
timestamp 1608254825
transform 1 0 16560 0 -1 13600
box -38 -48 2062 592
use sky130_fd_sc_hd__decap_4  FILLER_20_190
timestamp 1608254825
transform 1 0 18584 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_194
timestamp 1608254825
transform 1 0 18952 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_187
timestamp 1608254825
transform 1 0 18308 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_262
timestamp 1608254825
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _2239_
timestamp 1608254825
transform 1 0 18032 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1962_
timestamp 1608254825
transform 1 0 18952 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1960_
timestamp 1608254825
transform 1 0 18676 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_197
timestamp 1608254825
transform 1 0 19228 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_4  _1961_
timestamp 1608254825
transform 1 0 19596 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__o32ai_4  _2140_
timestamp 1608254825
transform 1 0 19320 0 1 12512
box -38 -48 2062 592
use sky130_fd_sc_hd__fill_1  FILLER_20_219
timestamp 1608254825
transform 1 0 21252 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_215
timestamp 1608254825
transform 1 0 20884 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_210
timestamp 1608254825
transform 1 0 20424 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_220
timestamp 1608254825
transform 1 0 21344 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_269
timestamp 1608254825
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__a41o_4  _2248_
timestamp 1608254825
transform 1 0 21344 0 -1 13600
box -38 -48 1602 592
use sky130_fd_sc_hd__buf_2  _2121_
timestamp 1608254825
transform 1 0 22080 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_245
timestamp 1608254825
transform 1 0 23644 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_237
timestamp 1608254825
transform 1 0 22908 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_240
timestamp 1608254825
transform 1 0 23184 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_232
timestamp 1608254825
transform 1 0 22448 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_263
timestamp 1608254825
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2604_
timestamp 1608254825
transform 1 0 23644 0 1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  _1696_
timestamp 1608254825
transform 1 0 24012 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1695_
timestamp 1608254825
transform 1 0 23276 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1554_
timestamp 1608254825
transform 1 0 22816 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_271
timestamp 1608254825
transform 1 0 26036 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_257
timestamp 1608254825
transform 1 0 24748 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_253
timestamp 1608254825
transform 1 0 24380 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_272
timestamp 1608254825
transform 1 0 26128 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_268
timestamp 1608254825
transform 1 0 25760 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_264
timestamp 1608254825
transform 1 0 25392 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_10_0_m1_clk_local
timestamp 1608254825
transform 1 0 25852 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_4  _1536_
timestamp 1608254825
transform 1 0 24840 0 -1 13600
box -38 -48 1234 592
use sky130_fd_sc_hd__a41oi_4  _1524_
timestamp 1608254825
transform 1 0 26312 0 1 12512
box -38 -48 2062 592
use sky130_fd_sc_hd__fill_1  FILLER_20_293
timestamp 1608254825
transform 1 0 28060 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_289
timestamp 1608254825
transform 1 0 27692 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_296
timestamp 1608254825
transform 1 0 28336 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_270
timestamp 1608254825
transform 1 0 26404 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1555_
timestamp 1608254825
transform 1 0 28152 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_4  _1525_
timestamp 1608254825
transform 1 0 26496 0 -1 13600
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_20_298
timestamp 1608254825
transform 1 0 28520 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_319
timestamp 1608254825
transform 1 0 30452 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_304
timestamp 1608254825
transform 1 0 29072 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_264
timestamp 1608254825
transform 1 0 29164 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_4  _1510_
timestamp 1608254825
transform 1 0 29256 0 1 12512
box -38 -48 1234 592
use sky130_fd_sc_hd__o32ai_4  _1491_
timestamp 1608254825
transform 1 0 28888 0 -1 13600
box -38 -48 2062 592
use sky130_fd_sc_hd__fill_1  FILLER_20_337
timestamp 1608254825
transform 1 0 32108 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_332
timestamp 1608254825
transform 1 0 31648 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_324
timestamp 1608254825
transform 1 0 30912 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_332
timestamp 1608254825
transform 1 0 31648 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_271
timestamp 1608254825
transform 1 0 32016 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_4  _1507_
timestamp 1608254825
transform 1 0 30820 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  _1449_
timestamp 1608254825
transform 1 0 32016 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_4  _1441_
timestamp 1608254825
transform 1 0 32200 0 -1 13600
box -38 -48 1234 592
use sky130_fd_sc_hd__buf_2  _1433_
timestamp 1608254825
transform 1 0 31280 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_351
timestamp 1608254825
transform 1 0 33396 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_362
timestamp 1608254825
transform 1 0 34408 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_345
timestamp 1608254825
transform 1 0 32844 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_addressalyzerBlock.SPI_CLK
timestamp 1608254825
transform 1 0 33764 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _2612_
timestamp 1608254825
transform 1 0 34040 0 -1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__a21oi_4  _1455_
timestamp 1608254825
transform 1 0 33212 0 1 12512
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_20_377
timestamp 1608254825
transform 1 0 35788 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_377
timestamp 1608254825
transform 1 0 35788 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_19_367
timestamp 1608254825
transform 1 0 34868 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_265
timestamp 1608254825
transform 1 0 34776 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2461_
timestamp 1608254825
transform 1 0 36156 0 1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__and2_4  _2114_
timestamp 1608254825
transform 1 0 35144 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_4  _1826_
timestamp 1608254825
transform 1 0 36156 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_406
timestamp 1608254825
transform 1 0 38456 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_402
timestamp 1608254825
transform 1 0 38088 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_393
timestamp 1608254825
transform 1 0 37260 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_406
timestamp 1608254825
transform 1 0 38456 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_400
timestamp 1608254825
transform 1 0 37904 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_272
timestamp 1608254825
transform 1 0 37628 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1608254825
transform -1 0 38824 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1608254825
transform -1 0 38824 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1514_
timestamp 1608254825
transform 1 0 37720 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_7
timestamp 1608254825
transform 1 0 1748 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_3
timestamp 1608254825
transform 1 0 1380 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1608254825
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _2419_
timestamp 1608254825
transform 1 0 1840 0 1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_21_27
timestamp 1608254825
transform 1 0 3588 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__o32ai_4  _2275_
timestamp 1608254825
transform 1 0 3956 0 1 13600
box -38 -48 2062 592
use sky130_fd_sc_hd__decap_4  FILLER_21_62
timestamp 1608254825
transform 1 0 6808 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_53
timestamp 1608254825
transform 1 0 5980 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_273
timestamp 1608254825
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_4  _2307_
timestamp 1608254825
transform 1 0 7176 0 1 13600
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_21_79
timestamp 1608254825
transform 1 0 8372 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_4  _2306_
timestamp 1608254825
transform 1 0 8740 0 1 13600
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_21_97
timestamp 1608254825
transform 1 0 10028 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_4  _2300_
timestamp 1608254825
transform 1 0 10396 0 1 13600
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_21_136
timestamp 1608254825
transform 1 0 13616 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_121
timestamp 1608254825
transform 1 0 12236 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_115
timestamp 1608254825
transform 1 0 11684 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_274
timestamp 1608254825
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_4  _2294_
timestamp 1608254825
transform 1 0 12420 0 1 13600
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_21_159
timestamp 1608254825
transform 1 0 15732 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2434_
timestamp 1608254825
transform 1 0 13984 0 1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_21_175
timestamp 1608254825
transform 1 0 17204 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_21_167
timestamp 1608254825
transform 1 0 16468 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _2240_
timestamp 1608254825
transform 1 0 16836 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1601_
timestamp 1608254825
transform 1 0 16100 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_203
timestamp 1608254825
transform 1 0 19780 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_275
timestamp 1608254825
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2440_
timestamp 1608254825
transform 1 0 18032 0 1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_21_226
timestamp 1608254825
transform 1 0 21896 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2441_
timestamp 1608254825
transform 1 0 20148 0 1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_21_240
timestamp 1608254825
transform 1 0 23184 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_230
timestamp 1608254825
transform 1 0 22264 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_276
timestamp 1608254825
transform 1 0 23552 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__and4_4  _2312_
timestamp 1608254825
transform 1 0 23644 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__and4_4  _2238_
timestamp 1608254825
transform 1 0 22356 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_21_274
timestamp 1608254825
transform 1 0 26312 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_254
timestamp 1608254825
transform 1 0 24472 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_m1_clk_local
timestamp 1608254825
transform 1 0 24840 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_4  _1532_
timestamp 1608254825
transform 1 0 25116 0 1 13600
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_6  FILLER_21_291
timestamp 1608254825
transform 1 0 27876 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_4  _1540_
timestamp 1608254825
transform 1 0 26680 0 1 13600
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_21_301
timestamp 1608254825
transform 1 0 28796 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_277
timestamp 1608254825
transform 1 0 29164 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__a22oi_4  _1492_
timestamp 1608254825
transform 1 0 29256 0 1 13600
box -38 -48 1602 592
use sky130_fd_sc_hd__buf_2  _1488_
timestamp 1608254825
transform 1 0 28428 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_338
timestamp 1608254825
transform 1 0 32200 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_331
timestamp 1608254825
transform 1 0 31556 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_323
timestamp 1608254825
transform 1 0 30820 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_addressalyzerBlock.SPI_CLK
timestamp 1608254825
transform 1 0 31924 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1448_
timestamp 1608254825
transform 1 0 31188 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__nand4_4  _1440_
timestamp 1608254825
transform 1 0 32384 0 1 13600
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_2  FILLER_21_364
timestamp 1608254825
transform 1 0 34592 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_357
timestamp 1608254825
transform 1 0 33948 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_11_0_addressalyzerBlock.SPI_CLK
timestamp 1608254825
transform 1 0 34316 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_380
timestamp 1608254825
transform 1 0 36064 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_367
timestamp 1608254825
transform 1 0 34868 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_278
timestamp 1608254825
transform 1 0 34776 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2450_
timestamp 1608254825
transform 1 0 36432 0 1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__and2_4  _2113_
timestamp 1608254825
transform 1 0 35420 0 1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_21_403
timestamp 1608254825
transform 1 0 38180 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1608254825
transform -1 0 38824 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_22_22
timestamp 1608254825
transform 1 0 3128 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1608254825
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _2515_
timestamp 1608254825
transform 1 0 1380 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  FILLER_22_32
timestamp 1608254825
transform 1 0 4048 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_1_0_m1_clk_local
timestamp 1608254825
transform 1 0 3680 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_279
timestamp 1608254825
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__o32ai_4  _2274_
timestamp 1608254825
transform 1 0 4324 0 -1 14688
box -38 -48 2062 592
use sky130_fd_sc_hd__fill_2  FILLER_22_65
timestamp 1608254825
transform 1 0 7084 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_57
timestamp 1608254825
transform 1 0 6348 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1943_
timestamp 1608254825
transform 1 0 7268 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_88
timestamp 1608254825
transform 1 0 9200 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_71
timestamp 1608254825
transform 1 0 7636 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_4  _2301_
timestamp 1608254825
transform 1 0 8004 0 -1 14688
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_22_106
timestamp 1608254825
transform 1 0 10856 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_280
timestamp 1608254825
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_4  _2303_
timestamp 1608254825
transform 1 0 9660 0 -1 14688
box -38 -48 1234 592
use sky130_fd_sc_hd__nand3_4  _2298_
timestamp 1608254825
transform 1 0 11224 0 -1 14688
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_6  FILLER_22_124
timestamp 1608254825
transform 1 0 12512 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_4  _2305_
timestamp 1608254825
transform 1 0 13064 0 -1 14688
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_2  FILLER_22_151
timestamp 1608254825
transform 1 0 14996 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_143
timestamp 1608254825
transform 1 0 14260 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_281
timestamp 1608254825
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_4  _2242_
timestamp 1608254825
transform 1 0 15272 0 -1 14688
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_6  FILLER_22_181
timestamp 1608254825
transform 1 0 17756 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_174
timestamp 1608254825
transform 1 0 17112 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_167
timestamp 1608254825
transform 1 0 16468 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2138_
timestamp 1608254825
transform 1 0 16836 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1964_
timestamp 1608254825
transform 1 0 17480 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_22_187
timestamp 1608254825
transform 1 0 18308 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__o32ai_4  _2141_
timestamp 1608254825
transform 1 0 18400 0 -1 14688
box -38 -48 2062 592
use sky130_fd_sc_hd__decap_4  FILLER_22_210
timestamp 1608254825
transform 1 0 20424 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_282
timestamp 1608254825
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__a41o_4  _2139_
timestamp 1608254825
transform 1 0 20884 0 -1 14688
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_22_232
timestamp 1608254825
transform 1 0 22448 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__a41o_4  _2310_
timestamp 1608254825
transform 1 0 22816 0 -1 14688
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_1  FILLER_22_274
timestamp 1608254825
transform 1 0 26312 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_270
timestamp 1608254825
transform 1 0 25944 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_253
timestamp 1608254825
transform 1 0 24380 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_4  _1543_
timestamp 1608254825
transform 1 0 24748 0 -1 14688
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_6  FILLER_22_293
timestamp 1608254825
transform 1 0 28060 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_276
timestamp 1608254825
transform 1 0 26496 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_283
timestamp 1608254825
transform 1 0 26404 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__nor3_4  _1482_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 26864 0 -1 14688
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_22_315
timestamp 1608254825
transform 1 0 30084 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_299
timestamp 1608254825
transform 1 0 28612 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_9_0_addressalyzerBlock.SPI_CLK
timestamp 1608254825
transform 1 0 28704 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_4  _1493_
timestamp 1608254825
transform 1 0 30452 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_4  _1489_
timestamp 1608254825
transform 1 0 28980 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_337
timestamp 1608254825
transform 1 0 32108 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_22_328
timestamp 1608254825
transform 1 0 31280 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_284
timestamp 1608254825
transform 1 0 32016 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_359
timestamp 1608254825
transform 1 0 34132 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_355
timestamp 1608254825
transform 1 0 33764 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_347
timestamp 1608254825
transform 1 0 33028 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_4  _1578_
timestamp 1608254825
transform 1 0 34224 0 -1 14688
box -38 -48 1234 592
use sky130_fd_sc_hd__buf_2  _1450_
timestamp 1608254825
transform 1 0 33396 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1422_
timestamp 1608254825
transform 1 0 32660 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_373
timestamp 1608254825
transform 1 0 35420 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_4  _1778_
timestamp 1608254825
transform 1 0 35788 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_401
timestamp 1608254825
transform 1 0 37996 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_22_389
timestamp 1608254825
transform 1 0 36892 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_285
timestamp 1608254825
transform 1 0 37628 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1608254825
transform -1 0 38824 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1423_
timestamp 1608254825
transform 1 0 37720 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_23_22
timestamp 1608254825
transform 1 0 3128 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_18
timestamp 1608254825
transform 1 0 2760 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_3
timestamp 1608254825
transform 1 0 1380 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1608254825
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__and2_4  _1959_
timestamp 1608254825
transform 1 0 2116 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_23_26
timestamp 1608254825
transform 1 0 3496 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2420_
timestamp 1608254825
transform 1 0 3864 0 1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_2  _1946_
timestamp 1608254825
transform 1 0 3220 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_23_66
timestamp 1608254825
transform 1 0 7176 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_57
timestamp 1608254825
transform 1 0 6348 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_49
timestamp 1608254825
transform 1 0 5612 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_286
timestamp 1608254825
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _2270_
timestamp 1608254825
transform 1 0 6808 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1956_
timestamp 1608254825
transform 1 0 5980 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_91
timestamp 1608254825
transform 1 0 9476 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2404_
timestamp 1608254825
transform 1 0 7728 0 1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_23_113
timestamp 1608254825
transform 1 0 11500 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_109
timestamp 1608254825
transform 1 0 11132 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_4  _2302_
timestamp 1608254825
transform 1 0 9844 0 1 14688
box -38 -48 1326 592
use sky130_fd_sc_hd__buf_2  _2291_
timestamp 1608254825
transform 1 0 11592 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_136
timestamp 1608254825
transform 1 0 13616 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_118
timestamp 1608254825
transform 1 0 11960 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_287
timestamp 1608254825
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_4  _2299_
timestamp 1608254825
transform 1 0 12420 0 1 14688
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_23_156
timestamp 1608254825
transform 1 0 15456 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_152
timestamp 1608254825
transform 1 0 15088 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_144
timestamp 1608254825
transform 1 0 14352 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _2297_
timestamp 1608254825
transform 1 0 13984 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2246_
timestamp 1608254825
transform 1 0 15180 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_179
timestamp 1608254825
transform 1 0 17572 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2439_
timestamp 1608254825
transform 1 0 15824 0 1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_23_200
timestamp 1608254825
transform 1 0 19504 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_23_187
timestamp 1608254825
transform 1 0 18308 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_288
timestamp 1608254825
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1966_
timestamp 1608254825
transform 1 0 18032 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_4  _1963_
timestamp 1608254825
transform 1 0 18676 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_23_213
timestamp 1608254825
transform 1 0 20700 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_208
timestamp 1608254825
transform 1 0 20240 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__a41o_4  _2263_
timestamp 1608254825
transform 1 0 21068 0 1 14688
box -38 -48 1602 592
use sky130_fd_sc_hd__buf_2  _1597_
timestamp 1608254825
transform 1 0 20332 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_249
timestamp 1608254825
transform 1 0 24012 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_242
timestamp 1608254825
transform 1 0 23368 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_234
timestamp 1608254825
transform 1 0 22632 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_289
timestamp 1608254825
transform 1 0 23552 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1581_
timestamp 1608254825
transform 1 0 23644 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_274
timestamp 1608254825
transform 1 0 26312 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_257
timestamp 1608254825
transform 1 0 24748 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_253
timestamp 1608254825
transform 1 0 24380 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_4  _1539_
timestamp 1608254825
transform 1 0 25116 0 1 14688
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _1490_
timestamp 1608254825
transform 1 0 24472 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_23_280
timestamp 1608254825
transform 1 0 26864 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__nor4_4  _1469_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 26956 0 1 14688
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_23_313
timestamp 1608254825
transform 1 0 29900 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_23_306
timestamp 1608254825
transform 1 0 29256 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_23_304
timestamp 1608254825
transform 1 0 29072 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_298
timestamp 1608254825
transform 1 0 28520 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_290
timestamp 1608254825
transform 1 0 29164 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2609_
timestamp 1608254825
transform 1 0 30268 0 1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  _1474_
timestamp 1608254825
transform 1 0 29532 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_336
timestamp 1608254825
transform 1 0 32016 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_23_362
timestamp 1608254825
transform 1 0 34408 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_344
timestamp 1608254825
transform 1 0 32752 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__nand4_4  _2326_
timestamp 1608254825
transform 1 0 32844 0 1 14688
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_23_380
timestamp 1608254825
transform 1 0 36064 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_291
timestamp 1608254825
transform 1 0 34776 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2451_
timestamp 1608254825
transform 1 0 36432 0 1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__o21ai_4  _1588_
timestamp 1608254825
transform 1 0 34868 0 1 14688
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_23_403
timestamp 1608254825
transform 1 0 38180 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1608254825
transform -1 0 38824 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_24_15
timestamp 1608254825
transform 1 0 2484 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_3
timestamp 1608254825
transform 1 0 1380 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1608254825
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_4  _1965_
timestamp 1608254825
transform 1 0 2576 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_24_42
timestamp 1608254825
transform 1 0 4968 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_32
timestamp 1608254825
transform 1 0 4048 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_25
timestamp 1608254825
transform 1 0 3404 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_292
timestamp 1608254825
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _1947_
timestamp 1608254825
transform 1 0 4140 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_24_50
timestamp 1608254825
transform 1 0 5704 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  _2406_
timestamp 1608254825
transform 1 0 6256 0 -1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  _1255_
timestamp 1608254825
transform 1 0 5336 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_91
timestamp 1608254825
transform 1 0 9476 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_87
timestamp 1608254825
transform 1 0 9108 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_75
timestamp 1608254825
transform 1 0 8004 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_105
timestamp 1608254825
transform 1 0 10764 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_93
timestamp 1608254825
transform 1 0 9660 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_293
timestamp 1608254825
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2408_
timestamp 1608254825
transform 1 0 11132 0 -1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_24_132
timestamp 1608254825
transform 1 0 13248 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_128
timestamp 1608254825
transform 1 0 12880 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_4  _2304_
timestamp 1608254825
transform 1 0 13340 0 -1 15776
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_6  FILLER_24_154
timestamp 1608254825
transform 1 0 15272 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_24_147
timestamp 1608254825
transform 1 0 14628 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_294
timestamp 1608254825
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_163
timestamp 1608254825
transform 1 0 16100 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__o32ai_4  _2145_
timestamp 1608254825
transform 1 0 16468 0 -1 15776
box -38 -48 2062 592
use sky130_fd_sc_hd__inv_2  _2117_
timestamp 1608254825
transform 1 0 15824 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_197
timestamp 1608254825
transform 1 0 19228 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_193
timestamp 1608254825
transform 1 0 18860 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_189
timestamp 1608254825
transform 1 0 18492 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_4  _2137_
timestamp 1608254825
transform 1 0 19596 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1603_
timestamp 1608254825
transform 1 0 18952 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_24_228
timestamp 1608254825
transform 1 0 22080 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_24_210
timestamp 1608254825
transform 1 0 20424 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_295
timestamp 1608254825
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__nor3_4  _2245_
timestamp 1608254825
transform 1 0 20884 0 -1 15776
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_24_246
timestamp 1608254825
transform 1 0 23736 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_236
timestamp 1608254825
transform 1 0 22816 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_4  _1600_
timestamp 1608254825
transform 1 0 22908 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _1580_
timestamp 1608254825
transform 1 0 24104 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_271
timestamp 1608254825
transform 1 0 26036 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_258
timestamp 1608254825
transform 1 0 24840 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_254
timestamp 1608254825
transform 1 0 24472 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_4  _1542_
timestamp 1608254825
transform 1 0 24932 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_293
timestamp 1608254825
transform 1 0 28060 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_296
timestamp 1608254825
transform 1 0 26404 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__o41a_4  _1538_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 26496 0 -1 15776
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_8  FILLER_24_315
timestamp 1608254825
transform 1 0 30084 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_297
timestamp 1608254825
transform 1 0 28428 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__nor4_4  _1548_
timestamp 1608254825
transform 1 0 28520 0 -1 15776
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_24_340
timestamp 1608254825
transform 1 0 32384 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_332
timestamp 1608254825
transform 1 0 31648 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_297
timestamp 1608254825
transform 1 0 32016 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _1983_
timestamp 1608254825
transform 1 0 30820 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1421_
timestamp 1608254825
transform 1 0 32108 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_361
timestamp 1608254825
transform 1 0 34316 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__nand4_4  _2335_
timestamp 1608254825
transform 1 0 32752 0 -1 15776
box -38 -48 1602 592
use sky130_fd_sc_hd__buf_2  _1217_
timestamp 1608254825
transform 1 0 34684 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_375
timestamp 1608254825
transform 1 0 35604 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_369
timestamp 1608254825
transform 1 0 35052 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__nand4_4  _1783_
timestamp 1608254825
transform 1 0 35696 0 -1 15776
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_1  FILLER_24_406
timestamp 1608254825
transform 1 0 38456 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_402
timestamp 1608254825
transform 1 0 38088 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_393
timestamp 1608254825
transform 1 0 37260 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_298
timestamp 1608254825
transform 1 0 37628 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1608254825
transform -1 0 38824 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1460_
timestamp 1608254825
transform 1 0 37720 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_3
timestamp 1608254825
transform 1 0 1380 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1608254825
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _2504_
timestamp 1608254825
transform 1 0 1932 0 1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_25_28
timestamp 1608254825
transform 1 0 3680 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  _2516_
timestamp 1608254825
transform 1 0 4232 0 1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_25_53
timestamp 1608254825
transform 1 0 5980 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_299
timestamp 1608254825
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2503_
timestamp 1608254825
transform 1 0 6808 0 1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  FILLER_25_89
timestamp 1608254825
transform 1 0 9292 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_25_81
timestamp 1608254825
transform 1 0 8556 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_25_111
timestamp 1608254825
transform 1 0 11316 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2403_
timestamp 1608254825
transform 1 0 9568 0 1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_25_130
timestamp 1608254825
transform 1 0 13064 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_25_123
timestamp 1608254825
transform 1 0 12420 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_118
timestamp 1608254825
transform 1 0 11960 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_300
timestamp 1608254825
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2405_
timestamp 1608254825
transform 1 0 13616 0 1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  _2292_
timestamp 1608254825
transform 1 0 12696 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2089_
timestamp 1608254825
transform 1 0 11684 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_155
timestamp 1608254825
transform 1 0 15364 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2447_
timestamp 1608254825
transform 1 0 15732 0 1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_25_182
timestamp 1608254825
transform 1 0 17848 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_178
timestamp 1608254825
transform 1 0 17480 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_188
timestamp 1608254825
transform 1 0 18400 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_301
timestamp 1608254825
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2505_
timestamp 1608254825
transform 1 0 18768 0 1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  _1886_
timestamp 1608254825
transform 1 0 18032 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_222
timestamp 1608254825
transform 1 0 21528 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_211
timestamp 1608254825
transform 1 0 20516 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__and2_4  _1969_
timestamp 1608254825
transform 1 0 20884 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_4  _1561_
timestamp 1608254825
transform 1 0 21896 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_25_245
timestamp 1608254825
transform 1 0 23644 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_243
timestamp 1608254825
transform 1 0 23460 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_235
timestamp 1608254825
transform 1 0 22724 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_302
timestamp 1608254825
transform 1 0 23552 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__a211o_4  _1599_
timestamp 1608254825
transform 1 0 24012 0 1 15776
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_25_271
timestamp 1608254825
transform 1 0 26036 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_267
timestamp 1608254825
transform 1 0 25668 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_263
timestamp 1608254825
transform 1 0 25300 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1467_
timestamp 1608254825
transform 1 0 25760 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_25_296
timestamp 1608254825
transform 1 0 28336 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_292
timestamp 1608254825
transform 1 0 27968 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_279
timestamp 1608254825
transform 1 0 26772 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1468_
timestamp 1608254825
transform 1 0 26404 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_4  _1429_
timestamp 1608254825
transform 1 0 27140 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_25_319
timestamp 1608254825
transform 1 0 30452 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_301
timestamp 1608254825
transform 1 0 28796 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_303
timestamp 1608254825
transform 1 0 29164 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_4  _1550_
timestamp 1608254825
transform 1 0 29256 0 1 15776
box -38 -48 1234 592
use sky130_fd_sc_hd__buf_2  _1451_
timestamp 1608254825
transform 1 0 28428 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_325
timestamp 1608254825
transform 1 0 31004 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2494_
timestamp 1608254825
transform 1 0 31096 0 1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_25_358
timestamp 1608254825
transform 1 0 34040 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_25_345
timestamp 1608254825
transform 1 0 32844 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_4  _1526_
timestamp 1608254825
transform 1 0 33212 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_25_380
timestamp 1608254825
transform 1 0 36064 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_367
timestamp 1608254825
transform 1 0 34868 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_304
timestamp 1608254825
transform 1 0 34776 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__nand3_4  _1779_
timestamp 1608254825
transform 1 0 36432 0 1 15776
box -38 -48 1326 592
use sky130_fd_sc_hd__o21a_4  _1598_
timestamp 1608254825
transform 1 0 34960 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_406
timestamp 1608254825
transform 1 0 38456 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_398
timestamp 1608254825
transform 1 0 37720 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1608254825
transform -1 0 38824 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_13
timestamp 1608254825
transform 1 0 2300 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_9
timestamp 1608254825
transform 1 0 1932 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_3
timestamp 1608254825
transform 1 0 1380 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_26_22
timestamp 1608254825
transform 1 0 3128 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1608254825
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1608254825
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _2507_
timestamp 1608254825
transform 1 0 1380 0 -1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_2  _1264_
timestamp 1608254825
transform 1 0 2024 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_4  _1263_
timestamp 1608254825
transform 1 0 2668 0 1 16864
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_8  FILLER_27_31
timestamp 1608254825
transform 1 0 3956 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_26_39
timestamp 1608254825
transform 1 0 4692 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_30
timestamp 1608254825
transform 1 0 3864 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_305
timestamp 1608254825
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _1970_
timestamp 1608254825
transform 1 0 4048 0 -1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__nand3_4  _1289_
timestamp 1608254825
transform 1 0 4692 0 1 16864
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_27_68
timestamp 1608254825
transform 1 0 7360 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_62
timestamp 1608254825
transform 1 0 6808 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_53
timestamp 1608254825
transform 1 0 5980 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_67
timestamp 1608254825
transform 1 0 7268 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_54
timestamp 1608254825
transform 1 0 6072 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_312
timestamp 1608254825
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _1967_
timestamp 1608254825
transform 1 0 6440 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__and2_4  _1958_
timestamp 1608254825
transform 1 0 5428 0 -1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _1254_
timestamp 1608254825
transform 1 0 6992 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_91
timestamp 1608254825
transform 1 0 9476 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_91
timestamp 1608254825
transform 1 0 9476 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_87
timestamp 1608254825
transform 1 0 9108 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_80
timestamp 1608254825
transform 1 0 8464 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2469_
timestamp 1608254825
transform 1 0 7728 0 1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__nor2_4  _2090_
timestamp 1608254825
transform 1 0 7636 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1290_
timestamp 1608254825
transform 1 0 8832 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_27_108
timestamp 1608254825
transform 1 0 11040 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_104
timestamp 1608254825
transform 1 0 10672 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_100
timestamp 1608254825
transform 1 0 10304 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_306
timestamp 1608254825
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_4  _2309_
timestamp 1608254825
transform 1 0 9844 0 1 16864
box -38 -48 1234 592
use sky130_fd_sc_hd__nand3_4  _2308_
timestamp 1608254825
transform 1 0 10764 0 -1 16864
box -38 -48 1326 592
use sky130_fd_sc_hd__and2_4  _2088_
timestamp 1608254825
transform 1 0 9660 0 -1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_27_130
timestamp 1608254825
transform 1 0 13064 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_123
timestamp 1608254825
transform 1 0 12420 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_120
timestamp 1608254825
transform 1 0 12144 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_125
timestamp 1608254825
transform 1 0 12604 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_119
timestamp 1608254825
transform 1 0 12052 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_313
timestamp 1608254825
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2448_
timestamp 1608254825
transform 1 0 12696 0 -1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_2  _2290_
timestamp 1608254825
transform 1 0 12788 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_4  _1615_
timestamp 1608254825
transform 1 0 13432 0 1 16864
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_1  FILLER_27_151
timestamp 1608254825
transform 1 0 14996 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_147
timestamp 1608254825
transform 1 0 14628 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_154
timestamp 1608254825
transform 1 0 15272 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_26_145
timestamp 1608254825
transform 1 0 14444 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_307
timestamp 1608254825
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2557_
timestamp 1608254825
transform 1 0 15088 0 1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_27_179
timestamp 1608254825
transform 1 0 17572 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_171
timestamp 1608254825
transform 1 0 16836 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_169
timestamp 1608254825
transform 1 0 16652 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2449_
timestamp 1608254825
transform 1 0 17020 0 -1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  _1880_
timestamp 1608254825
transform 1 0 17204 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_4  _1701_
timestamp 1608254825
transform 1 0 15824 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_27_191
timestamp 1608254825
transform 1 0 18676 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_192
timestamp 1608254825
transform 1 0 18768 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_314
timestamp 1608254825
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2597_
timestamp 1608254825
transform 1 0 19044 0 1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__and2_4  _1883_
timestamp 1608254825
transform 1 0 18032 0 1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__nand3_4  _1602_
timestamp 1608254825
transform 1 0 19136 0 -1 16864
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_27_214
timestamp 1608254825
transform 1 0 20792 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_215
timestamp 1608254825
transform 1 0 20884 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_210
timestamp 1608254825
transform 1 0 20424 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_308
timestamp 1608254825
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__nor4_4  _2289_
timestamp 1608254825
transform 1 0 21160 0 1 16864
box -38 -48 1602 592
use sky130_fd_sc_hd__a41o_4  _2279_
timestamp 1608254825
transform 1 0 21068 0 -1 16864
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_3  FILLER_27_245
timestamp 1608254825
transform 1 0 23644 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_27_235
timestamp 1608254825
transform 1 0 22724 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_26_234
timestamp 1608254825
transform 1 0 22632 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_m1_clk_local
timestamp 1608254825
transform 1 0 23276 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_315
timestamp 1608254825
transform 1 0 23552 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__a41oi_4  _2115_
timestamp 1608254825
transform 1 0 23184 0 -1 16864
box -38 -48 2062 592
use sky130_fd_sc_hd__o21ai_4  _1582_
timestamp 1608254825
transform 1 0 23920 0 1 16864
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_27_261
timestamp 1608254825
transform 1 0 25116 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_274
timestamp 1608254825
transform 1 0 26312 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_270
timestamp 1608254825
transform 1 0 25944 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_262
timestamp 1608254825
transform 1 0 25208 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__a32oi_4  _1563_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 25484 0 1 16864
box -38 -48 2062 592
use sky130_fd_sc_hd__buf_2  _1541_
timestamp 1608254825
transform 1 0 25576 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_287
timestamp 1608254825
transform 1 0 27508 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_296
timestamp 1608254825
transform 1 0 28336 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_279
timestamp 1608254825
transform 1 0 26772 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_309
timestamp 1608254825
transform 1 0 26404 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__and3_4  _1557_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 27876 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_4  _1552_
timestamp 1608254825
transform 1 0 27140 0 -1 16864
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _1466_
timestamp 1608254825
transform 1 0 26496 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_306
timestamp 1608254825
transform 1 0 29256 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_304
timestamp 1608254825
transform 1 0 29072 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_300
timestamp 1608254825
transform 1 0 28704 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_313
timestamp 1608254825
transform 1 0 29900 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_316
timestamp 1608254825
transform 1 0 29164 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__a41o_4  _1546_
timestamp 1608254825
transform 1 0 29440 0 1 16864
box -38 -48 1602 592
use sky130_fd_sc_hd__o21ai_4  _1544_
timestamp 1608254825
transform 1 0 28704 0 -1 16864
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_27_325
timestamp 1608254825
transform 1 0 31004 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_337
timestamp 1608254825
transform 1 0 32108 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_332
timestamp 1608254825
transform 1 0 31648 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_321
timestamp 1608254825
transform 1 0 30636 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_310
timestamp 1608254825
transform 1 0 32016 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_4  _2333_
timestamp 1608254825
transform 1 0 30820 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_4  _1547_
timestamp 1608254825
transform 1 0 32292 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__nand3_4  _1446_
timestamp 1608254825
transform 1 0 31372 0 1 16864
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_27_362
timestamp 1608254825
transform 1 0 34408 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_343
timestamp 1608254825
transform 1 0 32660 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_359
timestamp 1608254825
transform 1 0 34132 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_351
timestamp 1608254825
transform 1 0 33396 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2389_
timestamp 1608254825
transform 1 0 34500 0 -1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__a21oi_4  _2334_
timestamp 1608254825
transform 1 0 33212 0 1 16864
box -38 -48 1234 592
use sky130_fd_sc_hd__buf_2  _1184_
timestamp 1608254825
transform 1 0 33764 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_380
timestamp 1608254825
transform 1 0 36064 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_382
timestamp 1608254825
transform 1 0 36248 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_317
timestamp 1608254825
transform 1 0 34776 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2589_
timestamp 1608254825
transform 1 0 36432 0 1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__a21oi_4  _1782_
timestamp 1608254825
transform 1 0 34868 0 1 16864
box -38 -48 1234 592
use sky130_fd_sc_hd__buf_2  _1577_
timestamp 1608254825
transform 1 0 36616 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_403
timestamp 1608254825
transform 1 0 38180 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_406
timestamp 1608254825
transform 1 0 38456 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_402
timestamp 1608254825
transform 1 0 38088 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_396
timestamp 1608254825
transform 1 0 37536 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_390
timestamp 1608254825
transform 1 0 36984 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_311
timestamp 1608254825
transform 1 0 37628 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1608254825
transform -1 0 38824 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1608254825
transform -1 0 38824 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _2360_
timestamp 1608254825
transform 1 0 37720 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_7
timestamp 1608254825
transform 1 0 1748 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_3
timestamp 1608254825
transform 1 0 1380 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1608254825
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _2644_
timestamp 1608254825
transform 1 0 1840 0 -1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_28_45
timestamp 1608254825
transform 1 0 5244 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_41
timestamp 1608254825
transform 1 0 4876 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_27
timestamp 1608254825
transform 1 0 3588 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_318
timestamp 1608254825
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_4  _1252_
timestamp 1608254825
transform 1 0 4048 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_28_65
timestamp 1608254825
transform 1 0 7084 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2639_
timestamp 1608254825
transform 1 0 5336 0 -1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_28_91
timestamp 1608254825
transform 1 0 9476 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_85
timestamp 1608254825
transform 1 0 8924 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_81
timestamp 1608254825
transform 1 0 8556 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_77
timestamp 1608254825
transform 1 0 8188 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_69
timestamp 1608254825
transform 1 0 7452 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _1971_
timestamp 1608254825
transform 1 0 7544 0 -1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1279_
timestamp 1608254825
transform 1 0 8648 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_28_97
timestamp 1608254825
transform 1 0 10028 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_93
timestamp 1608254825
transform 1 0 9660 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_319
timestamp 1608254825
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2566_
timestamp 1608254825
transform 1 0 10120 0 -1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_28_117
timestamp 1608254825
transform 1 0 11868 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2558_
timestamp 1608254825
transform 1 0 12236 0 -1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_28_149
timestamp 1608254825
transform 1 0 14812 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_140
timestamp 1608254825
transform 1 0 13984 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_320
timestamp 1608254825
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1702_
timestamp 1608254825
transform 1 0 14536 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_4  _1642_
timestamp 1608254825
transform 1 0 15272 0 -1 17952
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_28_167
timestamp 1608254825
transform 1 0 16468 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_4  _1718_
timestamp 1608254825
transform 1 0 16836 0 -1 17952
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_28_203
timestamp 1608254825
transform 1 0 19780 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_195
timestamp 1608254825
transform 1 0 19044 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_184
timestamp 1608254825
transform 1 0 18032 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__and2_4  _1871_
timestamp 1608254825
transform 1 0 18400 0 -1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _1534_
timestamp 1608254825
transform 1 0 19412 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_220
timestamp 1608254825
transform 1 0 21344 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_215
timestamp 1608254825
transform 1 0 20884 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_210
timestamp 1608254825
transform 1 0 20424 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_321
timestamp 1608254825
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__a21o_4  _1595_
timestamp 1608254825
transform 1 0 21712 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1591_
timestamp 1608254825
transform 1 0 20148 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1427_
timestamp 1608254825
transform 1 0 20976 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_236
timestamp 1608254825
transform 1 0 22816 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__a41oi_4  _1587_
timestamp 1608254825
transform 1 0 23184 0 -1 17952
box -38 -48 2062 592
use sky130_fd_sc_hd__decap_4  FILLER_28_271
timestamp 1608254825
transform 1 0 26036 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_266
timestamp 1608254825
transform 1 0 25576 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_262
timestamp 1608254825
transform 1 0 25208 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1531_
timestamp 1608254825
transform 1 0 25668 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_287
timestamp 1608254825
transform 1 0 27508 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_283
timestamp 1608254825
transform 1 0 27140 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_322
timestamp 1608254825
transform 1 0 26404 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _1564_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 26496 0 -1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_4  _1553_
timestamp 1608254825
transform 1 0 27600 0 -1 17952
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_28_314
timestamp 1608254825
transform 1 0 29992 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_302
timestamp 1608254825
transform 1 0 28888 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__nand3_4  _1530_
timestamp 1608254825
transform 1 0 30360 0 -1 17952
box -38 -48 1326 592
use sky130_fd_sc_hd__buf_2  _1500_
timestamp 1608254825
transform 1 0 29624 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_332
timestamp 1608254825
transform 1 0 31648 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_323
timestamp 1608254825
transform 1 0 32016 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__a21o_4  _1442_
timestamp 1608254825
transform 1 0 32108 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_349
timestamp 1608254825
transform 1 0 33212 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_4  _1681_
timestamp 1608254825
transform 1 0 33764 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_373
timestamp 1608254825
transform 1 0 35420 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_367
timestamp 1608254825
transform 1 0 34868 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  _2595_
timestamp 1608254825
transform 1 0 35512 0 -1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_28_401
timestamp 1608254825
transform 1 0 37996 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_393
timestamp 1608254825
transform 1 0 37260 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_324
timestamp 1608254825
transform 1 0 37628 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1608254825
transform -1 0 38824 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1527_
timestamp 1608254825
transform 1 0 37720 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_29_22
timestamp 1608254825
transform 1 0 3128 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1608254825
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _2643_
timestamp 1608254825
transform 1 0 1380 0 1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_29_30
timestamp 1608254825
transform 1 0 3864 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__nand4_4  _1250_
timestamp 1608254825
transform 1 0 4048 0 1 17952
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_29_65
timestamp 1608254825
transform 1 0 7084 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_60
timestamp 1608254825
transform 1 0 6624 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_56
timestamp 1608254825
transform 1 0 6256 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_49
timestamp 1608254825
transform 1 0 5612 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_325
timestamp 1608254825
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1287_
timestamp 1608254825
transform 1 0 6808 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1267_
timestamp 1608254825
transform 1 0 5980 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_72
timestamp 1608254825
transform 1 0 7728 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2642_
timestamp 1608254825
transform 1 0 8096 0 1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_2  _1249_
timestamp 1608254825
transform 1 0 7452 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_95
timestamp 1608254825
transform 1 0 9844 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2564_
timestamp 1608254825
transform 1 0 10212 0 1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_29_130
timestamp 1608254825
transform 1 0 13064 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_118
timestamp 1608254825
transform 1 0 11960 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_4_0_addressalyzerBlock.SPI_CLK
timestamp 1608254825
transform 1 0 13616 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_326
timestamp 1608254825
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _1882_
timestamp 1608254825
transform 1 0 12420 0 1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_29_146
timestamp 1608254825
transform 1 0 14536 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2565_
timestamp 1608254825
transform 1 0 14904 0 1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__or2_4  _1641_
timestamp 1608254825
transform 1 0 13892 0 1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_29_179
timestamp 1608254825
transform 1 0 17572 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_169
timestamp 1608254825
transform 1 0 16652 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _1874_
timestamp 1608254825
transform 1 0 17204 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_29_184
timestamp 1608254825
transform 1 0 18032 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_327
timestamp 1608254825
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2560_
timestamp 1608254825
transform 1 0 18308 0 1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_29_224
timestamp 1608254825
transform 1 0 21712 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_213
timestamp 1608254825
transform 1 0 20700 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_206
timestamp 1608254825
transform 1 0 20056 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_6_0_addressalyzerBlock.SPI_CLK
timestamp 1608254825
transform 1 0 20424 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__and4_4  _2118_
timestamp 1608254825
transform 1 0 20884 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_4  _1586_
timestamp 1608254825
transform 1 0 22080 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_249
timestamp 1608254825
transform 1 0 24012 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_240
timestamp 1608254825
transform 1 0 23184 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_328
timestamp 1608254825
transform 1 0 23552 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1594_
timestamp 1608254825
transform 1 0 23644 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_272
timestamp 1608254825
transform 1 0 26128 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_29_256
timestamp 1608254825
transform 1 0 24656 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1562_
timestamp 1608254825
transform 1 0 24380 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_4  _1535_
timestamp 1608254825
transform 1 0 25024 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_289
timestamp 1608254825
transform 1 0 27692 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_4  _1556_
timestamp 1608254825
transform 1 0 26864 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _1537_
timestamp 1608254825
transform 1 0 28060 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_319
timestamp 1608254825
transform 1 0 30452 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_297
timestamp 1608254825
transform 1 0 28428 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_329
timestamp 1608254825
transform 1 0 29164 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_4  _1551_
timestamp 1608254825
transform 1 0 29256 0 1 17952
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_29_326
timestamp 1608254825
transform 1 0 31096 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__a41o_4  _1576_
timestamp 1608254825
transform 1 0 31464 0 1 17952
box -38 -48 1602 592
use sky130_fd_sc_hd__inv_2  _1443_
timestamp 1608254825
transform 1 0 30820 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_29_360
timestamp 1608254825
transform 1 0 34224 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_347
timestamp 1608254825
transform 1 0 33028 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_4  _1528_
timestamp 1608254825
transform 1 0 33396 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_29_380
timestamp 1608254825
transform 1 0 36064 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_330
timestamp 1608254825
transform 1 0 34776 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2588_
timestamp 1608254825
transform 1 0 36432 0 1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__a21oi_4  _1686_
timestamp 1608254825
transform 1 0 34868 0 1 17952
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_29_403
timestamp 1608254825
transform 1 0 38180 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1608254825
transform -1 0 38824 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_30_9
timestamp 1608254825
transform 1 0 1932 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_3
timestamp 1608254825
transform 1 0 1380 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1608254825
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__nand4_4  _1262_
timestamp 1608254825
transform 1 0 2024 0 -1 19040
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_6  FILLER_30_35
timestamp 1608254825
transform 1 0 4324 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_27
timestamp 1608254825
transform 1 0 3588 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_331
timestamp 1608254825
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_4  _1268_
timestamp 1608254825
transform 1 0 4876 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1251_
timestamp 1608254825
transform 1 0 4048 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_50
timestamp 1608254825
transform 1 0 5704 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__nand4_4  _1266_
timestamp 1608254825
transform 1 0 6072 0 -1 19040
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_6  FILLER_30_86
timestamp 1608254825
transform 1 0 9016 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_30_71
timestamp 1608254825
transform 1 0 7636 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_4  _1248_
timestamp 1608254825
transform 1 0 8188 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_30_113
timestamp 1608254825
transform 1 0 11500 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_102
timestamp 1608254825
transform 1 0 10488 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_1
timestamp 1608254825
transform 1 0 10672 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_332
timestamp 1608254825
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _1875_
timestamp 1608254825
transform 1 0 10856 0 -1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_4  _1278_
timestamp 1608254825
transform 1 0 9660 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_30_136
timestamp 1608254825
transform 1 0 13616 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2556_
timestamp 1608254825
transform 1 0 11868 0 -1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_30_152
timestamp 1608254825
transform 1 0 15088 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_148
timestamp 1608254825
transform 1 0 14720 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_140
timestamp 1608254825
transform 1 0 13984 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_333
timestamp 1608254825
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_4  _2217_
timestamp 1608254825
transform 1 0 15272 0 -1 19040
box -38 -48 1234 592
use sky130_fd_sc_hd__or2_4  _1854_
timestamp 1608254825
transform 1 0 14076 0 -1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_30_167
timestamp 1608254825
transform 1 0 16468 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2559_
timestamp 1608254825
transform 1 0 16836 0 -1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_30_190
timestamp 1608254825
transform 1 0 18584 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__and2_4  _1889_
timestamp 1608254825
transform 1 0 19596 0 -1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _1879_
timestamp 1608254825
transform 1 0 18952 0 -1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_30_218
timestamp 1608254825
transform 1 0 21160 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_212
timestamp 1608254825
transform 1 0 20608 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_334
timestamp 1608254825
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__nor3_4  _1669_
timestamp 1608254825
transform 1 0 21528 0 -1 19040
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _1589_
timestamp 1608254825
transform 1 0 20884 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1560_
timestamp 1608254825
transform 1 0 20240 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_235
timestamp 1608254825
transform 1 0 22724 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__a41oi_4  _2116_
timestamp 1608254825
transform 1 0 23276 0 -1 19040
box -38 -48 2062 592
use sky130_fd_sc_hd__decap_4  FILLER_30_271
timestamp 1608254825
transform 1 0 26036 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_263
timestamp 1608254825
transform 1 0 25300 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1694_
timestamp 1608254825
transform 1 0 25668 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_279
timestamp 1608254825
transform 1 0 26772 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_335
timestamp 1608254825
transform 1 0 26404 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2601_
timestamp 1608254825
transform 1 0 27140 0 -1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_2  _1424_
timestamp 1608254825
transform 1 0 26496 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_302
timestamp 1608254825
transform 1 0 28888 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2602_
timestamp 1608254825
transform 1 0 29256 0 -1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  FILLER_30_337
timestamp 1608254825
transform 1 0 32108 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_332
timestamp 1608254825
transform 1 0 31648 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_325
timestamp 1608254825
transform 1 0 31004 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_336
timestamp 1608254825
transform 1 0 32016 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__a21o_4  _1685_
timestamp 1608254825
transform 1 0 32384 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1435_
timestamp 1608254825
transform 1 0 31372 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_352
timestamp 1608254825
transform 1 0 33488 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__o41ai_4  _1682_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 33856 0 -1 19040
box -38 -48 2062 592
use sky130_fd_sc_hd__decap_6  FILLER_30_378
timestamp 1608254825
transform 1 0 35880 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_4  _1780_
timestamp 1608254825
transform 1 0 36432 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_30_401
timestamp 1608254825
transform 1 0 37996 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_393
timestamp 1608254825
transform 1 0 37260 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_337
timestamp 1608254825
transform 1 0 37628 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1608254825
transform -1 0 38824 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1444_
timestamp 1608254825
transform 1 0 37720 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_31_11
timestamp 1608254825
transform 1 0 2116 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_31_3
timestamp 1608254825
transform 1 0 1380 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1608254825
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _2640_
timestamp 1608254825
transform 1 0 2392 0 1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_31_40
timestamp 1608254825
transform 1 0 4784 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_33
timestamp 1608254825
transform 1 0 4140 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__and3_4  _1271_
timestamp 1608254825
transform 1 0 5152 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1256_
timestamp 1608254825
transform 1 0 4508 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_31_53
timestamp 1608254825
transform 1 0 5980 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_338
timestamp 1608254825
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__nand4_4  _1272_
timestamp 1608254825
transform 1 0 6808 0 1 19040
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_1  FILLER_31_85
timestamp 1608254825
transform 1 0 8924 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_79
timestamp 1608254825
transform 1 0 8372 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_4  _1276_
timestamp 1608254825
transform 1 0 9016 0 1 19040
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_31_110
timestamp 1608254825
transform 1 0 11224 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_99
timestamp 1608254825
transform 1 0 10212 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__and2_4  _1876_
timestamp 1608254825
transform 1 0 10580 0 1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1273_
timestamp 1608254825
transform 1 0 11592 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_31_131
timestamp 1608254825
transform 1 0 13156 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_123
timestamp 1608254825
transform 1 0 12420 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_121
timestamp 1608254825
transform 1 0 12236 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_117
timestamp 1608254825
transform 1 0 11868 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_339
timestamp 1608254825
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_4  _1843_
timestamp 1608254825
transform 1 0 13248 0 1 19040
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_31_145
timestamp 1608254825
transform 1 0 14444 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_4  _1855_
timestamp 1608254825
transform 1 0 14812 0 1 19040
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_1  FILLER_31_179
timestamp 1608254825
transform 1 0 17572 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_173
timestamp 1608254825
transform 1 0 17020 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_162
timestamp 1608254825
transform 1 0 16008 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_addressalyzerBlock.SPI_CLK
timestamp 1608254825
transform 1 0 17664 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__and2_4  _1872_
timestamp 1608254825
transform 1 0 16376 0 1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_31_195
timestamp 1608254825
transform 1 0 19044 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_191
timestamp 1608254825
transform 1 0 18676 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_addressalyzerBlock.SPI_CLK $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 19136 0 1 19040
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_340
timestamp 1608254825
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _1881_
timestamp 1608254825
transform 1 0 18032 0 1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_4  _2598_
timestamp 1608254825
transform 1 0 20976 0 1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_31_243
timestamp 1608254825
transform 1 0 23460 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_239
timestamp 1608254825
transform 1 0 23092 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_341
timestamp 1608254825
transform 1 0 23552 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__a41oi_4  _1596_
timestamp 1608254825
transform 1 0 23644 0 1 19040
box -38 -48 2062 592
use sky130_fd_sc_hd__buf_2  _1220_
timestamp 1608254825
transform 1 0 22724 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_271
timestamp 1608254825
transform 1 0 26036 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_267
timestamp 1608254825
transform 1 0 25668 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1549_
timestamp 1608254825
transform 1 0 26128 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_31_295
timestamp 1608254825
transform 1 0 28244 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_31_275
timestamp 1608254825
transform 1 0 26404 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_4  _1692_
timestamp 1608254825
transform 1 0 26772 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_31_315
timestamp 1608254825
transform 1 0 30084 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_31_303
timestamp 1608254825
transform 1 0 28980 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_342
timestamp 1608254825
transform 1 0 29164 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _1608_
timestamp 1608254825
transform 1 0 29256 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_31_339
timestamp 1608254825
transform 1 0 32292 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_321
timestamp 1608254825
transform 1 0 30636 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__nand4_4  _1445_
timestamp 1608254825
transform 1 0 30728 0 1 19040
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_1  FILLER_31_365
timestamp 1608254825
transform 1 0 34684 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_357
timestamp 1608254825
transform 1 0 33948 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__nand3_4  _1684_
timestamp 1608254825
transform 1 0 32660 0 1 19040
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_8  FILLER_31_376
timestamp 1608254825
transform 1 0 35696 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_343
timestamp 1608254825
transform 1 0 34776 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2462_
timestamp 1608254825
transform 1 0 36432 0 1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__nor2_4  _1679_
timestamp 1608254825
transform 1 0 34868 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_31_403
timestamp 1608254825
transform 1 0 38180 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1608254825
transform -1 0 38824 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_32_11
timestamp 1608254825
transform 1 0 2116 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_32_3
timestamp 1608254825
transform 1 0 1380 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1608254825
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_4  _1286_
timestamp 1608254825
transform 1 0 2392 0 -1 20128
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_1  FILLER_32_32
timestamp 1608254825
transform 1 0 4048 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_27
timestamp 1608254825
transform 1 0 3588 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_344
timestamp 1608254825
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__nor4_4  _1261_
timestamp 1608254825
transform 1 0 4140 0 -1 20128
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_32_66
timestamp 1608254825
transform 1 0 7176 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_56
timestamp 1608254825
transform 1 0 6256 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_50
timestamp 1608254825
transform 1 0 5704 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_4  _1265_
timestamp 1608254825
transform 1 0 6348 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_32_91
timestamp 1608254825
transform 1 0 9476 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_87
timestamp 1608254825
transform 1 0 9108 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__nand4_4  _1277_
timestamp 1608254825
transform 1 0 7544 0 -1 20128
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_1  FILLER_32_97
timestamp 1608254825
transform 1 0 10028 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_93
timestamp 1608254825
transform 1 0 9660 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_345
timestamp 1608254825
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2563_
timestamp 1608254825
transform 1 0 10120 0 -1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_32_132
timestamp 1608254825
transform 1 0 13248 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_128
timestamp 1608254825
transform 1 0 12880 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_117
timestamp 1608254825
transform 1 0 11868 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__and2_4  _1884_
timestamp 1608254825
transform 1 0 12236 0 -1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_4  _1756_
timestamp 1608254825
transform 1 0 13340 0 -1 20128
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_32_146
timestamp 1608254825
transform 1 0 14536 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_addressalyzerBlock.SPI_CLK
timestamp 1608254825
transform 1 0 14904 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_346
timestamp 1608254825
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _1719_
timestamp 1608254825
transform 1 0 15272 0 -1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_32_161
timestamp 1608254825
transform 1 0 15916 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2551_
timestamp 1608254825
transform 1 0 16284 0 -1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_32_192
timestamp 1608254825
transform 1 0 18768 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_184
timestamp 1608254825
transform 1 0 18032 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_m1_clk_local
timestamp 1608254825
transform 1 0 18952 0 -1 20128
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_1  FILLER_32_219
timestamp 1608254825
transform 1 0 21252 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_215
timestamp 1608254825
transform 1 0 20884 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_347
timestamp 1608254825
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _1590_
timestamp 1608254825
transform 1 0 21344 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_32_242
timestamp 1608254825
transform 1 0 23368 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_229
timestamp 1608254825
transform 1 0 22172 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_m1_clk_local
timestamp 1608254825
transform 1 0 23736 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_4  _1606_
timestamp 1608254825
transform 1 0 22540 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_4  _1593_
timestamp 1608254825
transform 1 0 24012 0 -1 20128
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_32_271
timestamp 1608254825
transform 1 0 26036 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_262
timestamp 1608254825
transform 1 0 25208 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1687_
timestamp 1608254825
transform 1 0 25760 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_295
timestamp 1608254825
transform 1 0 28244 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_276
timestamp 1608254825
transform 1 0 26496 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_348
timestamp 1608254825
transform 1 0 26404 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_4  _1699_
timestamp 1608254825
transform 1 0 27048 0 -1 20128
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_32_315
timestamp 1608254825
transform 1 0 30084 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_307
timestamp 1608254825
transform 1 0 29348 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_302
timestamp 1608254825
transform 1 0 28888 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_addressalyzerBlock.SPI_CLK
timestamp 1608254825
transform 1 0 28612 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1585_
timestamp 1608254825
transform 1 0 29716 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1529_
timestamp 1608254825
transform 1 0 29072 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1221_
timestamp 1608254825
transform 1 0 30452 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_337
timestamp 1608254825
transform 1 0 32108 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_335
timestamp 1608254825
transform 1 0 31924 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_331
timestamp 1608254825
transform 1 0 31556 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_323
timestamp 1608254825
transform 1 0 30820 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_349
timestamp 1608254825
transform 1 0 32016 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1545_
timestamp 1608254825
transform 1 0 31188 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_352
timestamp 1608254825
transform 1 0 33488 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2387_
timestamp 1608254825
transform 1 0 33856 0 -1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__and3_4  _2338_
timestamp 1608254825
transform 1 0 32660 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_32_379
timestamp 1608254825
transform 1 0 35972 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_375
timestamp 1608254825
transform 1 0 35604 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_4  _1785_
timestamp 1608254825
transform 1 0 36064 0 -1 20128
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_6  FILLER_32_401
timestamp 1608254825
transform 1 0 37996 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_393
timestamp 1608254825
transform 1 0 37260 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_350
timestamp 1608254825
transform 1 0 37628 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1608254825
transform -1 0 38824 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1678_
timestamp 1608254825
transform 1 0 37720 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_14
timestamp 1608254825
transform 1 0 2392 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_3
timestamp 1608254825
transform 1 0 1380 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_22
timestamp 1608254825
transform 1 0 3128 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1608254825
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1608254825
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _2638_
timestamp 1608254825
transform 1 0 1380 0 1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__nand2_4  _1296_
timestamp 1608254825
transform 1 0 1564 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  _1227_
timestamp 1608254825
transform 1 0 2760 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_34_36
timestamp 1608254825
transform 1 0 4416 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_32
timestamp 1608254825
transform 1 0 4048 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_27
timestamp 1608254825
transform 1 0 3588 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_29
timestamp 1608254825
transform 1 0 3772 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_357
timestamp 1608254825
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1293_
timestamp 1608254825
transform 1 0 3496 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_4  _1288_
timestamp 1608254825
transform 1 0 4324 0 1 20128
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _1259_
timestamp 1608254825
transform 1 0 4140 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__nor4_4  _1247_
timestamp 1608254825
transform 1 0 4784 0 -1 21216
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_8  FILLER_34_57
timestamp 1608254825
transform 1 0 6348 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_60
timestamp 1608254825
transform 1 0 6624 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_56
timestamp 1608254825
transform 1 0 6256 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_48
timestamp 1608254825
transform 1 0 5520 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_351
timestamp 1608254825
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__and3_4  _1282_
timestamp 1608254825
transform 1 0 7084 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__o41ai_4  _1281_
timestamp 1608254825
transform 1 0 6808 0 1 20128
box -38 -48 2062 592
use sky130_fd_sc_hd__buf_2  _1257_
timestamp 1608254825
transform 1 0 5888 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_88
timestamp 1608254825
transform 1 0 9200 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_81
timestamp 1608254825
transform 1 0 8556 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_74
timestamp 1608254825
transform 1 0 7912 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_84
timestamp 1608254825
transform 1 0 8832 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2641_
timestamp 1608254825
transform 1 0 9200 0 1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_2  _1280_
timestamp 1608254825
transform 1 0 8924 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1224_
timestamp 1608254825
transform 1 0 8280 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_34_113
timestamp 1608254825
transform 1 0 11500 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_93
timestamp 1608254825
transform 1 0 9660 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_107
timestamp 1608254825
transform 1 0 10948 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_358
timestamp 1608254825
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2633_
timestamp 1608254825
transform 1 0 9752 0 -1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__and2_4  _1885_
timestamp 1608254825
transform 1 0 11316 0 1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_34_125
timestamp 1608254825
transform 1 0 12604 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_118
timestamp 1608254825
transform 1 0 11960 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_352
timestamp 1608254825
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2555_
timestamp 1608254825
transform 1 0 12420 0 1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__o21ai_4  _1755_
timestamp 1608254825
transform 1 0 12788 0 -1 21216
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_6  FILLER_34_140
timestamp 1608254825
transform 1 0 13984 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_142
timestamp 1608254825
transform 1 0 14168 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_5_0_addressalyzerBlock.SPI_CLK
timestamp 1608254825
transform 1 0 14536 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1741_
timestamp 1608254825
transform 1 0 14536 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_154
timestamp 1608254825
transform 1 0 15272 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_149
timestamp 1608254825
transform 1 0 14812 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_152
timestamp 1608254825
transform 1 0 15088 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_359
timestamp 1608254825
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1691_
timestamp 1608254825
transform 1 0 14812 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_4  _2207_
timestamp 1608254825
transform 1 0 15640 0 -1 21216
box -38 -48 1234 592
use sky130_fd_sc_hd__a21oi_4  _1720_
timestamp 1608254825
transform 1 0 15456 0 1 20128
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_34_171
timestamp 1608254825
transform 1 0 16836 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_177
timestamp 1608254825
transform 1 0 17388 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_169
timestamp 1608254825
transform 1 0 16652 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2oi_4  _2206_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 17204 0 -1 21216
box -38 -48 1970 592
use sky130_fd_sc_hd__buf_2  _1614_
timestamp 1608254825
transform 1 0 17020 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_200
timestamp 1608254825
transform 1 0 19504 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_196
timestamp 1608254825
transform 1 0 19136 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_184
timestamp 1608254825
transform 1 0 18032 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_addressalyzerBlock.SPI_CLK
timestamp 1608254825
transform 1 0 18400 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_353
timestamp 1608254825
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2552_
timestamp 1608254825
transform 1 0 18676 0 1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__and4_4  _1643_
timestamp 1608254825
transform 1 0 19596 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_34_219
timestamp 1608254825
transform 1 0 21252 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_215
timestamp 1608254825
transform 1 0 20884 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_210
timestamp 1608254825
transform 1 0 20424 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_218
timestamp 1608254825
transform 1 0 21160 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_360
timestamp 1608254825
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _2148_
timestamp 1608254825
transform 1 0 20792 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_4  _1664_
timestamp 1608254825
transform 1 0 21344 0 -1 21216
box -38 -48 1326 592
use sky130_fd_sc_hd__buf_2  _1650_
timestamp 1608254825
transform 1 0 20424 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_4  _1592_
timestamp 1608254825
transform 1 0 21344 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_34_234
timestamp 1608254825
transform 1 0 22632 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_249
timestamp 1608254825
transform 1 0 24012 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_237
timestamp 1608254825
transform 1 0 22908 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_229
timestamp 1608254825
transform 1 0 22172 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_8_0_m1_clk_local
timestamp 1608254825
transform 1 0 23276 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_354
timestamp 1608254825
transform 1 0 23552 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2599_
timestamp 1608254825
transform 1 0 23000 0 -1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  _1579_
timestamp 1608254825
transform 1 0 23644 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1426_
timestamp 1608254825
transform 1 0 22540 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_273
timestamp 1608254825
transform 1 0 26220 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_34_265
timestamp 1608254825
transform 1 0 25484 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_34_257
timestamp 1608254825
transform 1 0 24748 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_264
timestamp 1608254825
transform 1 0 25392 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_256
timestamp 1608254825
transform 1 0 24656 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _2594_
timestamp 1608254825
transform 1 0 25484 0 1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  _1583_
timestamp 1608254825
transform 1 0 25116 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1558_
timestamp 1608254825
transform 1 0 24380 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_34_280
timestamp 1608254825
transform 1 0 26864 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_276
timestamp 1608254825
transform 1 0 26496 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_284
timestamp 1608254825
transform 1 0 27232 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_361
timestamp 1608254825
transform 1 0 26404 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__nand4_4  _1698_
timestamp 1608254825
transform 1 0 26956 0 -1 21216
box -38 -48 1602 592
use sky130_fd_sc_hd__o21ai_4  _1693_
timestamp 1608254825
transform 1 0 27600 0 1 20128
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_34_298
timestamp 1608254825
transform 1 0 28520 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_310
timestamp 1608254825
transform 1 0 29624 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_301
timestamp 1608254825
transform 1 0 28796 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_355
timestamp 1608254825
transform 1 0 29164 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2393_
timestamp 1608254825
transform 1 0 28888 0 -1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _2388_
timestamp 1608254825
transform 1 0 29992 0 1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  _2101_
timestamp 1608254825
transform 1 0 29256 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_332
timestamp 1608254825
transform 1 0 31648 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_327
timestamp 1608254825
transform 1 0 31188 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_34_321
timestamp 1608254825
transform 1 0 30636 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_333
timestamp 1608254825
transform 1 0 31740 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_362
timestamp 1608254825
transform 1 0 32016 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_4  _2336_
timestamp 1608254825
transform 1 0 32108 0 1 20128
box -38 -48 1234 592
use sky130_fd_sc_hd__a21o_4  _2328_
timestamp 1608254825
transform 1 0 32108 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _1454_
timestamp 1608254825
transform 1 0 31280 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_349
timestamp 1608254825
transform 1 0 33212 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_362
timestamp 1608254825
transform 1 0 34408 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_354
timestamp 1608254825
transform 1 0 33672 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_350
timestamp 1608254825
transform 1 0 33304 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__o41ai_4  _2327_
timestamp 1608254825
transform 1 0 33580 0 -1 21216
box -38 -48 2062 592
use sky130_fd_sc_hd__or2_4  _1680_
timestamp 1608254825
transform 1 0 33764 0 1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_34_383
timestamp 1608254825
transform 1 0 36340 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_375
timestamp 1608254825
transform 1 0 35604 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_33_378
timestamp 1608254825
transform 1 0 35880 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_367
timestamp 1608254825
transform 1 0 34868 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_356
timestamp 1608254825
transform 1 0 34776 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2453_
timestamp 1608254825
transform 1 0 36248 0 1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__nand2_4  _2111_
timestamp 1608254825
transform 1 0 35052 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  _1784_
timestamp 1608254825
transform 1 0 36432 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_34_401
timestamp 1608254825
transform 1 0 37996 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_393
timestamp 1608254825
transform 1 0 37260 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_401
timestamp 1608254825
transform 1 0 37996 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_363
timestamp 1608254825
transform 1 0 37628 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1608254825
transform -1 0 38824 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1608254825
transform -1 0 38824 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1575_
timestamp 1608254825
transform 1 0 37720 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_7
timestamp 1608254825
transform 1 0 1748 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_3
timestamp 1608254825
transform 1 0 1380 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1608254825
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1297_
timestamp 1608254825
transform 1 0 1472 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__nand4_4  _1295_
timestamp 1608254825
transform 1 0 2116 0 1 21216
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_1  FILLER_35_34
timestamp 1608254825
transform 1 0 4232 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_28
timestamp 1608254825
transform 1 0 3680 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__o41a_4  _1285_
timestamp 1608254825
transform 1 0 4324 0 1 21216
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_6  FILLER_35_62
timestamp 1608254825
transform 1 0 6808 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_60
timestamp 1608254825
transform 1 0 6624 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_52
timestamp 1608254825
transform 1 0 5888 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_364
timestamp 1608254825
transform 1 0 6716 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1225_
timestamp 1608254825
transform 1 0 7360 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_82
timestamp 1608254825
transform 1 0 8648 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_78
timestamp 1608254825
transform 1 0 8280 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_72
timestamp 1608254825
transform 1 0 7728 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_4  _1326_
timestamp 1608254825
transform 1 0 9016 0 1 21216
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _1245_
timestamp 1608254825
transform 1 0 8372 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_35_110
timestamp 1608254825
transform 1 0 11224 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_106
timestamp 1608254825
transform 1 0 10856 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_99
timestamp 1608254825
transform 1 0 10212 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1323_
timestamp 1608254825
transform 1 0 10580 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1315_
timestamp 1608254825
transform 1 0 11316 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_130
timestamp 1608254825
transform 1 0 13064 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_126
timestamp 1608254825
transform 1 0 12696 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_121
timestamp 1608254825
transform 1 0 12236 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_115
timestamp 1608254825
transform 1 0 11684 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_365
timestamp 1608254825
transform 1 0 12328 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_4  _1754_
timestamp 1608254825
transform 1 0 13156 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1327_
timestamp 1608254825
transform 1 0 12420 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_150
timestamp 1608254825
transform 1 0 14904 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_143
timestamp 1608254825
transform 1 0 14260 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_4  _2228_
timestamp 1608254825
transform 1 0 15272 0 1 21216
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _1648_
timestamp 1608254825
transform 1 0 14628 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_35_175
timestamp 1608254825
transform 1 0 17204 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_167
timestamp 1608254825
transform 1 0 16468 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__and2_4  _1890_
timestamp 1608254825
transform 1 0 17296 0 1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _1640_
timestamp 1608254825
transform 1 0 16836 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_366
timestamp 1608254825
transform 1 0 17940 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_4  _2195_
timestamp 1608254825
transform 1 0 18032 0 1 21216
box -38 -48 1234 592
use sky130_fd_sc_hd__nand4_4  _1613_
timestamp 1608254825
transform 1 0 19228 0 1 21216
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_8  FILLER_35_214
timestamp 1608254825
transform 1 0 20792 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__nand3_4  _1567_
timestamp 1608254825
transform 1 0 21528 0 1 21216
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_1  FILLER_35_243
timestamp 1608254825
transform 1 0 23460 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_236
timestamp 1608254825
transform 1 0 22816 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_9_0_m1_clk_local
timestamp 1608254825
transform 1 0 23184 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_367
timestamp 1608254825
transform 1 0 23552 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _1604_
timestamp 1608254825
transform 1 0 23644 0 1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_35_252
timestamp 1608254825
transform 1 0 24288 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2600_
timestamp 1608254825
transform 1 0 24656 0 1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_35_296
timestamp 1608254825
transform 1 0 28336 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_292
timestamp 1608254825
transform 1 0 27968 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_275
timestamp 1608254825
transform 1 0 26404 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_4  _1573_
timestamp 1608254825
transform 1 0 26772 0 1 21216
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_35_319
timestamp 1608254825
transform 1 0 30452 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_301
timestamp 1608254825
transform 1 0 28796 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_368
timestamp 1608254825
transform 1 0 29164 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__nor3_4  _2340_
timestamp 1608254825
transform 1 0 29256 0 1 21216
box -38 -48 1234 592
use sky130_fd_sc_hd__buf_2  _1565_
timestamp 1608254825
transform 1 0 28428 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_332
timestamp 1608254825
transform 1 0 31648 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_4  _2337_
timestamp 1608254825
transform 1 0 32200 0 1 21216
box -38 -48 1326 592
use sky130_fd_sc_hd__nor2_4  _1434_
timestamp 1608254825
transform 1 0 30820 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_35_365
timestamp 1608254825
transform 1 0 34684 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_359
timestamp 1608254825
transform 1 0 34132 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_352
timestamp 1608254825
transform 1 0 33488 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1185_
timestamp 1608254825
transform 1 0 33856 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_386
timestamp 1608254825
transform 1 0 36616 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_369
timestamp 1608254825
transform 1 0 34776 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2390_
timestamp 1608254825
transform 1 0 34868 0 1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_35_403
timestamp 1608254825
transform 1 0 38180 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1608254825
transform -1 0 38824 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_4  _2100_
timestamp 1608254825
transform 1 0 36984 0 1 21216
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_36_10
timestamp 1608254825
transform 1 0 2024 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_3
timestamp 1608254825
transform 1 0 1380 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1608254825
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_4  _1294_
timestamp 1608254825
transform 1 0 2392 0 -1 22304
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _1291_
timestamp 1608254825
transform 1 0 1748 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_36_41
timestamp 1608254825
transform 1 0 4876 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_36_27
timestamp 1608254825
transform 1 0 3588 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_370
timestamp 1608254825
transform 1 0 3956 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_4  _1300_
timestamp 1608254825
transform 1 0 4048 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_36_52
timestamp 1608254825
transform 1 0 5888 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_47
timestamp 1608254825
transform 1 0 5428 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1304_
timestamp 1608254825
transform 1 0 5520 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__nand4_4  _1260_
timestamp 1608254825
transform 1 0 6624 0 -1 22304
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_36_85
timestamp 1608254825
transform 1 0 8924 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_77
timestamp 1608254825
transform 1 0 8188 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_m1_clk_local
timestamp 1608254825
transform 1 0 9292 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1311_
timestamp 1608254825
transform 1 0 8556 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_107
timestamp 1608254825
transform 1 0 10948 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_371
timestamp 1608254825
transform 1 0 9568 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__nand3_4  _1322_
timestamp 1608254825
transform 1 0 9660 0 -1 22304
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_36_134
timestamp 1608254825
transform 1 0 13432 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2634_
timestamp 1608254825
transform 1 0 11684 0 -1 22304
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_36_147
timestamp 1608254825
transform 1 0 14628 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_372
timestamp 1608254825
transform 1 0 15180 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__and3_4  _1856_
timestamp 1608254825
transform 1 0 15272 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__and3_4  _1652_
timestamp 1608254825
transform 1 0 13800 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_36_167
timestamp 1608254825
transform 1 0 16468 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_163
timestamp 1608254825
transform 1 0 16100 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2oi_4  _2184_
timestamp 1608254825
transform 1 0 16560 0 -1 22304
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_3  FILLER_36_196
timestamp 1608254825
transform 1 0 19136 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_189
timestamp 1608254825
transform 1 0 18492 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_7_0_addressalyzerBlock.SPI_CLK
timestamp 1608254825
transform 1 0 18860 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__and4_4  _1609_
timestamp 1608254825
transform 1 0 19412 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_36_219
timestamp 1608254825
transform 1 0 21252 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_36_208
timestamp 1608254825
transform 1 0 20240 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_373
timestamp 1608254825
transform 1 0 20792 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1605_
timestamp 1608254825
transform 1 0 20884 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__nand4_4  _1428_
timestamp 1608254825
transform 1 0 21988 0 -1 22304
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_36_244
timestamp 1608254825
transform 1 0 23552 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1425_
timestamp 1608254825
transform 1 0 23920 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_271
timestamp 1608254825
transform 1 0 26036 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_252
timestamp 1608254825
transform 1 0 24288 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_4  _1572_
timestamp 1608254825
transform 1 0 24840 0 -1 22304
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_36_291
timestamp 1608254825
transform 1 0 27876 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_276
timestamp 1608254825
transform 1 0 26496 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_374
timestamp 1608254825
transform 1 0 26404 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__nor3_4  _1690_
timestamp 1608254825
transform 1 0 28244 0 -1 22304
box -38 -48 1234 592
use sky130_fd_sc_hd__nor3_4  _1688_
timestamp 1608254825
transform 1 0 26680 0 -1 22304
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_36_308
timestamp 1608254825
transform 1 0 29440 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_4  _1729_
timestamp 1608254825
transform 1 0 29808 0 -1 22304
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_36_332
timestamp 1608254825
transform 1 0 31648 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_325
timestamp 1608254825
transform 1 0 31004 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_375
timestamp 1608254825
transform 1 0 32016 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__o32ai_4  _2329_
timestamp 1608254825
transform 1 0 32108 0 -1 22304
box -38 -48 2062 592
use sky130_fd_sc_hd__inv_2  _1574_
timestamp 1608254825
transform 1 0 31372 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_359
timestamp 1608254825
transform 1 0 34132 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__a22oi_4  _2330_
timestamp 1608254825
transform 1 0 34500 0 -1 22304
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_36_380
timestamp 1608254825
transform 1 0 36064 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__and3_4  _2099_
timestamp 1608254825
transform 1 0 36432 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_36_401
timestamp 1608254825
transform 1 0 37996 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_36_393
timestamp 1608254825
transform 1 0 37260 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_376
timestamp 1608254825
transform 1 0 37628 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1608254825
transform -1 0 38824 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1683_
timestamp 1608254825
transform 1 0 37720 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_22
timestamp 1608254825
transform 1 0 3128 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1608254825
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _2637_
timestamp 1608254825
transform 1 0 1380 0 1 22304
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_37_40
timestamp 1608254825
transform 1 0 4784 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_4  _1292_
timestamp 1608254825
transform 1 0 3496 0 1 22304
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_6  FILLER_37_62
timestamp 1608254825
transform 1 0 6808 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_37_55
timestamp 1608254825
transform 1 0 6164 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_377
timestamp 1608254825
transform 1 0 6716 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__and4_4  _1305_
timestamp 1608254825
transform 1 0 7360 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  _1226_
timestamp 1608254825
transform 1 0 5336 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_37_81
timestamp 1608254825
transform 1 0 8556 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_77
timestamp 1608254825
transform 1 0 8188 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__a41oi_4  _1325_
timestamp 1608254825
transform 1 0 8648 0 1 22304
box -38 -48 2062 592
use sky130_fd_sc_hd__fill_1  FILLER_37_108
timestamp 1608254825
transform 1 0 11040 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_104
timestamp 1608254825
transform 1 0 10672 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_4  _1244_
timestamp 1608254825
transform 1 0 11132 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_37_132
timestamp 1608254825
transform 1 0 13248 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_37_118
timestamp 1608254825
transform 1 0 11960 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_378
timestamp 1608254825
transform 1 0 12328 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__and4_4  _1316_
timestamp 1608254825
transform 1 0 12420 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_37_159
timestamp 1608254825
transform 1 0 15732 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__a2bb2oi_4  _2227_
timestamp 1608254825
transform 1 0 13800 0 1 22304
box -38 -48 1970 592
use sky130_fd_sc_hd__fill_1  FILLER_37_182
timestamp 1608254825
transform 1 0 17848 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_178
timestamp 1608254825
transform 1 0 17480 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_4  _2185_
timestamp 1608254825
transform 1 0 16284 0 1 22304
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_37_203
timestamp 1608254825
transform 1 0 19780 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_188
timestamp 1608254825
transform 1 0 18400 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_379
timestamp 1608254825
transform 1 0 17940 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _1649_
timestamp 1608254825
transform 1 0 18952 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _1644_
timestamp 1608254825
transform 1 0 18032 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_224
timestamp 1608254825
transform 1 0 21712 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_216
timestamp 1608254825
transform 1 0 20976 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_4  _1647_
timestamp 1608254825
transform 1 0 20148 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _1584_
timestamp 1608254825
transform 1 0 21804 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_243
timestamp 1608254825
transform 1 0 23460 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_37_237
timestamp 1608254825
transform 1 0 22908 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_37_229
timestamp 1608254825
transform 1 0 22172 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_380
timestamp 1608254825
transform 1 0 23552 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1659_
timestamp 1608254825
transform 1 0 22540 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_4  _1559_
timestamp 1608254825
transform 1 0 23644 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_37_262
timestamp 1608254825
transform 1 0 25208 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_254
timestamp 1608254825
transform 1 0 24472 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_4  _1569_
timestamp 1608254825
transform 1 0 25300 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_283
timestamp 1608254825
transform 1 0 27140 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_275
timestamp 1608254825
transform 1 0 26404 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_4  _2324_
timestamp 1608254825
transform 1 0 27324 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_319
timestamp 1608254825
transform 1 0 30452 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_297
timestamp 1608254825
transform 1 0 28428 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_381
timestamp 1608254825
transform 1 0 29164 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__nor3_4  _1728_
timestamp 1608254825
transform 1 0 29256 0 1 22304
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_37_327
timestamp 1608254825
transform 1 0 31188 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2386_
timestamp 1608254825
transform 1 0 31556 0 1 22304
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  _1566_
timestamp 1608254825
transform 1 0 30820 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_362
timestamp 1608254825
transform 1 0 34408 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_354
timestamp 1608254825
transform 1 0 33672 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_350
timestamp 1608254825
transform 1 0 33304 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__or2_4  _2105_
timestamp 1608254825
transform 1 0 33764 0 1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_37_376
timestamp 1608254825
transform 1 0 35696 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_382
timestamp 1608254825
transform 1 0 34776 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2452_
timestamp 1608254825
transform 1 0 36064 0 1 22304
box -38 -48 1786 592
use sky130_fd_sc_hd__nand2_4  _2112_
timestamp 1608254825
transform 1 0 34868 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_37_399
timestamp 1608254825
transform 1 0 37812 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1608254825
transform -1 0 38824 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_9
timestamp 1608254825
transform 1 0 1932 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_38_3
timestamp 1608254825
transform 1 0 1380 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1608254825
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1302_
timestamp 1608254825
transform 1 0 1656 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_4  _1301_
timestamp 1608254825
transform 1 0 2300 0 -1 23392
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_2  FILLER_38_32
timestamp 1608254825
transform 1 0 4048 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_27
timestamp 1608254825
transform 1 0 3588 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_383
timestamp 1608254825
transform 1 0 3956 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2635_
timestamp 1608254825
transform 1 0 4232 0 -1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_38_57
timestamp 1608254825
transform 1 0 6348 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_53
timestamp 1608254825
transform 1 0 5980 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__a41oi_4  _1312_
timestamp 1608254825
transform 1 0 6440 0 -1 23392
box -38 -48 2062 592
use sky130_fd_sc_hd__decap_4  FILLER_38_88
timestamp 1608254825
transform 1 0 9200 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_80
timestamp 1608254825
transform 1 0 8464 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1303_
timestamp 1608254825
transform 1 0 8832 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_38_101
timestamp 1608254825
transform 1 0 10396 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_38_93
timestamp 1608254825
transform 1 0 9660 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_384
timestamp 1608254825
transform 1 0 9568 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__nand4_4  _1318_
timestamp 1608254825
transform 1 0 10672 0 -1 23392
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_8  FILLER_38_128
timestamp 1608254825
transform 1 0 12880 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_38_121
timestamp 1608254825
transform 1 0 12236 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_4  _1653_
timestamp 1608254825
transform 1 0 13616 0 -1 23392
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _1320_
timestamp 1608254825
transform 1 0 12604 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_38_154
timestamp 1608254825
transform 1 0 15272 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_149
timestamp 1608254825
transform 1 0 14812 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_385
timestamp 1608254825
transform 1 0 15180 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1651_
timestamp 1608254825
transform 1 0 15456 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_160
timestamp 1608254825
transform 1 0 15824 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2oi_4  _2161_
timestamp 1608254825
transform 1 0 16192 0 -1 23392
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_4  FILLER_38_202
timestamp 1608254825
transform 1 0 19688 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_185
timestamp 1608254825
transform 1 0 18124 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_4  _2149_
timestamp 1608254825
transform 1 0 18492 0 -1 23392
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_38_228
timestamp 1608254825
transform 1 0 22080 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_210
timestamp 1608254825
transform 1 0 20424 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_386
timestamp 1608254825
transform 1 0 20792 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__nor3_4  _1654_
timestamp 1608254825
transform 1 0 20884 0 -1 23392
box -38 -48 1234 592
use sky130_fd_sc_hd__buf_2  _1610_
timestamp 1608254825
transform 1 0 20056 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_244
timestamp 1608254825
transform 1 0 23552 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_236
timestamp 1608254825
transform 1 0 22816 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__and4_4  _1667_
timestamp 1608254825
transform 1 0 23920 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _1568_
timestamp 1608254825
transform 1 0 23184 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1219_
timestamp 1608254825
transform 1 0 22448 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_273
timestamp 1608254825
transform 1 0 26220 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_265
timestamp 1608254825
transform 1 0 25484 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_38_257
timestamp 1608254825
transform 1 0 24748 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1668_
timestamp 1608254825
transform 1 0 25116 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_295
timestamp 1608254825
transform 1 0 28244 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_387
timestamp 1608254825
transform 1 0 26404 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2394_
timestamp 1608254825
transform 1 0 26496 0 -1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_38_302
timestamp 1608254825
transform 1 0 28888 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_4  _1730_
timestamp 1608254825
transform 1 0 29256 0 -1 23392
box -38 -48 1326 592
use sky130_fd_sc_hd__inv_2  _1670_
timestamp 1608254825
transform 1 0 28612 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_38_337
timestamp 1608254825
transform 1 0 32108 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_332
timestamp 1608254825
transform 1 0 31648 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_320
timestamp 1608254825
transform 1 0 30544 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_388
timestamp 1608254825
transform 1 0 32016 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _2106_
timestamp 1608254825
transform 1 0 32384 0 -1 23392
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _1781_
timestamp 1608254825
transform 1 0 31280 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_347
timestamp 1608254825
transform 1 0 33028 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2385_
timestamp 1608254825
transform 1 0 33396 0 -1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_38_388
timestamp 1608254825
transform 1 0 36800 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_378
timestamp 1608254825
transform 1 0 35880 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_370
timestamp 1608254825
transform 1 0 35144 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_4  _1736_
timestamp 1608254825
transform 1 0 35972 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_38_401
timestamp 1608254825
transform 1 0 37996 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_396
timestamp 1608254825
transform 1 0 37536 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_389
timestamp 1608254825
transform 1 0 37628 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1608254825
transform -1 0 38824 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1839_
timestamp 1608254825
transform 1 0 37720 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_9
timestamp 1608254825
transform 1 0 1932 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_40_3
timestamp 1608254825
transform 1 0 1380 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_39_7
timestamp 1608254825
transform 1 0 1748 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_3
timestamp 1608254825
transform 1 0 1380 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1608254825
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1608254825
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2345_
timestamp 1608254825
transform 1 0 1656 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_20
timestamp 1608254825
transform 1 0 2944 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_4  _2086_
timestamp 1608254825
transform 1 0 1840 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__a21oi_4  _2085_
timestamp 1608254825
transform 1 0 2300 0 -1 24480
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_8  FILLER_40_32
timestamp 1608254825
transform 1 0 4048 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_30
timestamp 1608254825
transform 1 0 3864 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_26
timestamp 1608254825
transform 1 0 3496 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_27
timestamp 1608254825
transform 1 0 3588 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_396
timestamp 1608254825
transform 1 0 3956 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1299_
timestamp 1608254825
transform 1 0 3312 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_38
timestamp 1608254825
transform 1 0 4600 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1314_
timestamp 1608254825
transform 1 0 4324 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _2636_
timestamp 1608254825
transform 1 0 4784 0 -1 24480
box -38 -48 1786 592
use sky130_fd_sc_hd__o21ai_4  _1313_
timestamp 1608254825
transform 1 0 4968 0 1 23392
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_40_59
timestamp 1608254825
transform 1 0 6532 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_62
timestamp 1608254825
transform 1 0 6808 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_55
timestamp 1608254825
transform 1 0 6164 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_390
timestamp 1608254825
transform 1 0 6716 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1339_
timestamp 1608254825
transform 1 0 7176 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_4  _1307_
timestamp 1608254825
transform 1 0 6900 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_88
timestamp 1608254825
transform 1 0 9200 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_75
timestamp 1608254825
transform 1 0 8004 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_91
timestamp 1608254825
transform 1 0 9476 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_70
timestamp 1608254825
transform 1 0 7544 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__and4_4  _1338_
timestamp 1608254825
transform 1 0 8372 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__nand4_4  _1246_
timestamp 1608254825
transform 1 0 7912 0 1 23392
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_8  FILLER_40_105
timestamp 1608254825
transform 1 0 10764 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_39_105
timestamp 1608254825
transform 1 0 10764 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_95
timestamp 1608254825
transform 1 0 9844 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_397
timestamp 1608254825
transform 1 0 9568 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_4  _1341_
timestamp 1608254825
transform 1 0 9660 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__and4_4  _1330_
timestamp 1608254825
transform 1 0 9936 0 1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  _1319_
timestamp 1608254825
transform 1 0 11132 0 1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_4  _1317_
timestamp 1608254825
transform 1 0 11500 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_131
timestamp 1608254825
transform 1 0 13156 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_40_125
timestamp 1608254825
transform 1 0 12604 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_136
timestamp 1608254825
transform 1 0 13616 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_123
timestamp 1608254825
transform 1 0 12420 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_118
timestamp 1608254825
transform 1 0 11960 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_391
timestamp 1608254825
transform 1 0 12328 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_4  _2186_
timestamp 1608254825
transform 1 0 12512 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__o21ai_4  _1742_
timestamp 1608254825
transform 1 0 13248 0 -1 24480
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_6  FILLER_40_158
timestamp 1608254825
transform 1 0 15640 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_40_145
timestamp 1608254825
transform 1 0 14444 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_39_153
timestamp 1608254825
transform 1 0 15180 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_398
timestamp 1608254825
transform 1 0 15180 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_4  _1857_
timestamp 1608254825
transform 1 0 13984 0 1 23392
box -38 -48 1234 592
use sky130_fd_sc_hd__buf_2  _1646_
timestamp 1608254825
transform 1 0 15272 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1645_
timestamp 1608254825
transform 1 0 15548 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_40_177
timestamp 1608254825
transform 1 0 17388 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_39_177
timestamp 1608254825
transform 1 0 17388 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_160
timestamp 1608254825
transform 1 0 15824 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_4  _2188_
timestamp 1608254825
transform 1 0 16192 0 -1 24480
box -38 -48 1234 592
use sky130_fd_sc_hd__o21ai_4  _2162_
timestamp 1608254825
transform 1 0 16192 0 1 23392
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_1  FILLER_40_205
timestamp 1608254825
transform 1 0 19964 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_197
timestamp 1608254825
transform 1 0 19228 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_183
timestamp 1608254825
transform 1 0 17940 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_39_205
timestamp 1608254825
transform 1 0 19964 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_201
timestamp 1608254825
transform 1 0 19596 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_184
timestamp 1608254825
transform 1 0 18032 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_392
timestamp 1608254825
transform 1 0 17940 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_4  _2210_
timestamp 1608254825
transform 1 0 18032 0 -1 24480
box -38 -48 1234 592
use sky130_fd_sc_hd__o21ai_4  _2173_
timestamp 1608254825
transform 1 0 18400 0 1 23392
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_6  FILLER_40_228
timestamp 1608254825
transform 1 0 22080 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_40_210
timestamp 1608254825
transform 1 0 20424 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_215
timestamp 1608254825
transform 1 0 20884 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_399
timestamp 1608254825
transform 1 0 20792 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_4  _2190_
timestamp 1608254825
transform 1 0 20884 0 -1 24480
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_4  _2189_
timestamp 1608254825
transform 1 0 20056 0 1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__nor3_4  _1665_
timestamp 1608254825
transform 1 0 21252 0 1 23392
box -38 -48 1234 592
use sky130_fd_sc_hd__buf_2  _1405_
timestamp 1608254825
transform 1 0 20056 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_239
timestamp 1608254825
transform 1 0 23092 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_234
timestamp 1608254825
transform 1 0 22632 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_232
timestamp 1608254825
transform 1 0 22448 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1570_
timestamp 1608254825
transform 1 0 22724 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1190_
timestamp 1608254825
transform 1 0 22816 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_245
timestamp 1608254825
transform 1 0 23644 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_240
timestamp 1608254825
transform 1 0 23184 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_393
timestamp 1608254825
transform 1 0 23552 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__a211o_4  _1724_
timestamp 1608254825
transform 1 0 23828 0 1 23392
box -38 -48 1326 592
use sky130_fd_sc_hd__nor3_4  _1671_
timestamp 1608254825
transform 1 0 23460 0 -1 24480
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_40_271
timestamp 1608254825
transform 1 0 26036 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_263
timestamp 1608254825
transform 1 0 25300 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_256
timestamp 1608254825
transform 1 0 24656 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_269
timestamp 1608254825
transform 1 0 25852 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_261
timestamp 1608254825
transform 1 0 25116 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_4  _2325_
timestamp 1608254825
transform 1 0 25944 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _1663_
timestamp 1608254825
transform 1 0 25668 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1189_
timestamp 1608254825
transform 1 0 25024 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_40_286
timestamp 1608254825
transform 1 0 27416 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_40_280
timestamp 1608254825
transform 1 0 26864 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_282
timestamp 1608254825
transform 1 0 27048 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_400
timestamp 1608254825
transform 1 0 26404 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1870_
timestamp 1608254825
transform 1 0 26496 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_4  _1732_
timestamp 1608254825
transform 1 0 27508 0 -1 24480
box -38 -48 1234 592
use sky130_fd_sc_hd__nor3_4  _1731_
timestamp 1608254825
transform 1 0 27416 0 1 23392
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_40_300
timestamp 1608254825
transform 1 0 28704 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_39_306
timestamp 1608254825
transform 1 0 29256 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_39_299
timestamp 1608254825
transform 1 0 28612 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_394
timestamp 1608254825
transform 1 0 29164 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2391_
timestamp 1608254825
transform 1 0 29072 0 -1 24480
box -38 -48 1786 592
use sky130_fd_sc_hd__a211o_4  _2332_
timestamp 1608254825
transform 1 0 29532 0 1 23392
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_40_332
timestamp 1608254825
transform 1 0 31648 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_327
timestamp 1608254825
transform 1 0 31188 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_323
timestamp 1608254825
transform 1 0 30820 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_323
timestamp 1608254825
transform 1 0 30820 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_401
timestamp 1608254825
transform 1 0 32016 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2392_
timestamp 1608254825
transform 1 0 31188 0 1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__nand2_4  _2322_
timestamp 1608254825
transform 1 0 32108 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _1212_
timestamp 1608254825
transform 1 0 31280 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_346
timestamp 1608254825
transform 1 0 32936 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_362
timestamp 1608254825
transform 1 0 34408 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_352
timestamp 1608254825
transform 1 0 33488 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_346
timestamp 1608254825
transform 1 0 32936 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_4  _2339_
timestamp 1608254825
transform 1 0 33488 0 -1 24480
box -38 -48 1326 592
use sky130_fd_sc_hd__nor2_4  _2331_
timestamp 1608254825
transform 1 0 33580 0 1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_40_366
timestamp 1608254825
transform 1 0 34776 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_383
timestamp 1608254825
transform 1 0 36340 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_379
timestamp 1608254825
transform 1 0 35972 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_39_367
timestamp 1608254825
transform 1 0 34868 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_395
timestamp 1608254825
transform 1 0 34776 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2463_
timestamp 1608254825
transform 1 0 36432 0 1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__nor4_4  _2102_
timestamp 1608254825
transform 1 0 35512 0 -1 24480
box -38 -48 1602 592
use sky130_fd_sc_hd__nor2_4  _2092_
timestamp 1608254825
transform 1 0 35144 0 1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_40_401
timestamp 1608254825
transform 1 0 37996 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_40_391
timestamp 1608254825
transform 1 0 37076 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_403
timestamp 1608254825
transform 1 0 38180 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_402
timestamp 1608254825
transform 1 0 37628 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1608254825
transform -1 0 38824 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1608254825
transform -1 0 38824 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1737_
timestamp 1608254825
transform 1 0 37720 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_41_14
timestamp 1608254825
transform 1 0 2392 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_3
timestamp 1608254825
transform 1 0 1380 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1608254825
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _2471_
timestamp 1608254825
transform 1 0 2760 0 1 24480
box -38 -48 1786 592
use sky130_fd_sc_hd__nor2_4  _2087_
timestamp 1608254825
transform 1 0 1564 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_41_41
timestamp 1608254825
transform 1 0 4876 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_37
timestamp 1608254825
transform 1 0 4508 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_4  _1308_
timestamp 1608254825
transform 1 0 4968 0 1 24480
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_41_62
timestamp 1608254825
transform 1 0 6808 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_60
timestamp 1608254825
transform 1 0 6624 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_56
timestamp 1608254825
transform 1 0 6256 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_403
timestamp 1608254825
transform 1 0 6716 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_4  _1343_
timestamp 1608254825
transform 1 0 7176 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_86
timestamp 1608254825
transform 1 0 9016 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_41_78
timestamp 1608254825
transform 1 0 8280 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__a41oi_4  _1340_
timestamp 1608254825
transform 1 0 9200 0 1 24480
box -38 -48 2062 592
use sky130_fd_sc_hd__decap_4  FILLER_41_110
timestamp 1608254825
transform 1 0 11224 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1328_
timestamp 1608254825
transform 1 0 11592 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_135
timestamp 1608254825
transform 1 0 13524 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_118
timestamp 1608254825
transform 1 0 11960 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_404
timestamp 1608254825
transform 1 0 12328 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_4  _1331_
timestamp 1608254825
transform 1 0 12420 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_41_157
timestamp 1608254825
transform 1 0 15548 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_41_151
timestamp 1608254825
transform 1 0 14996 0 1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_4  _2163_
timestamp 1608254825
transform 1 0 13892 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _1655_
timestamp 1608254825
transform 1 0 15640 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_179
timestamp 1608254825
transform 1 0 17572 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_162
timestamp 1608254825
transform 1 0 16008 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_4  _2165_
timestamp 1608254825
transform 1 0 16376 0 1 24480
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_1  FILLER_41_203
timestamp 1608254825
transform 1 0 19780 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_41_197
timestamp 1608254825
transform 1 0 19228 0 1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_184
timestamp 1608254825
transform 1 0 18032 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_405
timestamp 1608254825
transform 1 0 17940 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__a21o_4  _2209_
timestamp 1608254825
transform 1 0 18124 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _1406_
timestamp 1608254825
transform 1 0 19872 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_208
timestamp 1608254825
transform 1 0 20240 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__o41ai_4  _2172_
timestamp 1608254825
transform 1 0 20976 0 1 24480
box -38 -48 2062 592
use sky130_fd_sc_hd__decap_6  FILLER_41_249
timestamp 1608254825
transform 1 0 24012 0 1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_41_238
timestamp 1608254825
transform 1 0 23000 0 1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_406
timestamp 1608254825
transform 1 0 23552 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1571_
timestamp 1608254825
transform 1 0 23644 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_268
timestamp 1608254825
transform 1 0 25760 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_4  _2212_
timestamp 1608254825
transform 1 0 24564 0 1 24480
box -38 -48 1234 592
use sky130_fd_sc_hd__buf_2  _1666_
timestamp 1608254825
transform 1 0 26128 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_276
timestamp 1608254825
transform 1 0 26496 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_4  _1733_
timestamp 1608254825
transform 1 0 27232 0 1 24480
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_41_315
timestamp 1608254825
transform 1 0 30084 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_297
timestamp 1608254825
transform 1 0 28428 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_407
timestamp 1608254825
transform 1 0 29164 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _2236_
timestamp 1608254825
transform 1 0 29256 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1689_
timestamp 1608254825
transform 1 0 30452 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_41_341
timestamp 1608254825
transform 1 0 32476 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_322
timestamp 1608254825
transform 1 0 30728 0 1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_4  _2323_
timestamp 1608254825
transform 1 0 31280 0 1 24480
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_41_362
timestamp 1608254825
transform 1 0 34408 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_349
timestamp 1608254825
transform 1 0 33212 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__and4_4  _2104_
timestamp 1608254825
transform 1 0 33580 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _1186_
timestamp 1608254825
transform 1 0 32844 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_386
timestamp 1608254825
transform 1 0 36616 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_408
timestamp 1608254825
transform 1 0 34776 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2459_
timestamp 1608254825
transform 1 0 34868 0 1 24480
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_41_399
timestamp 1608254825
transform 1 0 37812 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1608254825
transform -1 0 38824 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_4  _1738_
timestamp 1608254825
transform 1 0 36984 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_42_22
timestamp 1608254825
transform 1 0 3128 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1608254825
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _2472_
timestamp 1608254825
transform 1 0 1380 0 -1 25568
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_42_44
timestamp 1608254825
transform 1 0 5152 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_36
timestamp 1608254825
transform 1 0 4416 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_30
timestamp 1608254825
transform 1 0 3864 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_409
timestamp 1608254825
transform 1 0 3956 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _2078_
timestamp 1608254825
transform 1 0 4048 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_4  _1309_
timestamp 1608254825
transform 1 0 5244 0 -1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_42_54
timestamp 1608254825
transform 1 0 6072 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2630_
timestamp 1608254825
transform 1 0 6440 0 -1 25568
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_42_91
timestamp 1608254825
transform 1 0 9476 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_85
timestamp 1608254825
transform 1 0 8924 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_77
timestamp 1608254825
transform 1 0 8188 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1243_
timestamp 1608254825
transform 1 0 8556 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_112
timestamp 1608254825
transform 1 0 11408 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_410
timestamp 1608254825
transform 1 0 9568 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2631_
timestamp 1608254825
transform 1 0 9660 0 -1 25568
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_42_124
timestamp 1608254825
transform 1 0 12512 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_120
timestamp 1608254825
transform 1 0 12144 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2632_
timestamp 1608254825
transform 1 0 12604 0 -1 25568
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  _1329_
timestamp 1608254825
transform 1 0 11776 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_154
timestamp 1608254825
transform 1 0 15272 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_152
timestamp 1608254825
transform 1 0 15088 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_144
timestamp 1608254825
transform 1 0 14352 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_411
timestamp 1608254825
transform 1 0 15180 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1611_
timestamp 1608254825
transform 1 0 15640 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_178
timestamp 1608254825
transform 1 0 17480 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_162
timestamp 1608254825
transform 1 0 16008 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_4  _2164_
timestamp 1608254825
transform 1 0 16376 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1337_
timestamp 1608254825
transform 1 0 17848 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_185
timestamp 1608254825
transform 1 0 18124 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2613_
timestamp 1608254825
transform 1 0 18492 0 -1 25568
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_42_215
timestamp 1608254825
transform 1 0 20884 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_42_208
timestamp 1608254825
transform 1 0 20240 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_412
timestamp 1608254825
transform 1 0 20792 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__o41ai_4  _2194_
timestamp 1608254825
transform 1 0 21436 0 -1 25568
box -38 -48 2062 592
use sky130_fd_sc_hd__decap_6  FILLER_42_243
timestamp 1608254825
transform 1 0 23460 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__or4_4  _2234_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 24012 0 -1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_42_271
timestamp 1608254825
transform 1 0 26036 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_258
timestamp 1608254825
transform 1 0 24840 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_4  _2211_
timestamp 1608254825
transform 1 0 25208 0 -1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_42_285
timestamp 1608254825
transform 1 0 27324 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_413
timestamp 1608254825
transform 1 0 26404 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2435_
timestamp 1608254825
transform 1 0 27876 0 -1 25568
box -38 -48 1786 592
use sky130_fd_sc_hd__nand2_4  _2235_
timestamp 1608254825
transform 1 0 26496 0 -1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_42_310
timestamp 1608254825
transform 1 0 29624 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_4  _1218_
timestamp 1608254825
transform 1 0 30360 0 -1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_42_340
timestamp 1608254825
transform 1 0 32384 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_335
timestamp 1608254825
transform 1 0 31924 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_327
timestamp 1608254825
transform 1 0 31188 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_414
timestamp 1608254825
transform 1 0 32016 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1697_
timestamp 1608254825
transform 1 0 32108 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_42_363
timestamp 1608254825
transform 1 0 34500 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _2458_
timestamp 1608254825
transform 1 0 32752 0 -1 25568
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_42_371
timestamp 1608254825
transform 1 0 35236 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2468_
timestamp 1608254825
transform 1 0 35328 0 -1 25568
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_42_406
timestamp 1608254825
transform 1 0 38456 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_402
timestamp 1608254825
transform 1 0 38088 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_391
timestamp 1608254825
transform 1 0 37076 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_415
timestamp 1608254825
transform 1 0 37628 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1608254825
transform -1 0 38824 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1222_
timestamp 1608254825
transform 1 0 37720 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_11
timestamp 1608254825
transform 1 0 2116 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_7
timestamp 1608254825
transform 1 0 1748 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_3
timestamp 1608254825
transform 1 0 1380 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1608254825
transform 1 0 1104 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2080_
timestamp 1608254825
transform 1 0 1840 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_4  _2079_
timestamp 1608254825
transform 1 0 2484 0 1 25568
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_43_40
timestamp 1608254825
transform 1 0 4784 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_29
timestamp 1608254825
transform 1 0 3772 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__or2_4  _2081_
timestamp 1608254825
transform 1 0 4140 0 1 25568
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _1284_
timestamp 1608254825
transform 1 0 5152 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_67
timestamp 1608254825
transform 1 0 7268 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_62
timestamp 1608254825
transform 1 0 6808 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_43_55
timestamp 1608254825
transform 1 0 6164 0 1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_48
timestamp 1608254825
transform 1 0 5520 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_416
timestamp 1608254825
transform 1 0 6716 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1334_
timestamp 1608254825
transform 1 0 6900 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1310_
timestamp 1608254825
transform 1 0 5888 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__a41oi_4  _1342_
timestamp 1608254825
transform 1 0 7636 0 1 25568
box -38 -48 2062 592
use sky130_fd_sc_hd__fill_1  FILLER_43_105
timestamp 1608254825
transform 1 0 10764 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_101
timestamp 1608254825
transform 1 0 10396 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_93
timestamp 1608254825
transform 1 0 9660 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1321_
timestamp 1608254825
transform 1 0 10028 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__and4_4  _1242_
timestamp 1608254825
transform 1 0 10856 0 1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_43_134
timestamp 1608254825
transform 1 0 13432 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_126
timestamp 1608254825
transform 1 0 12696 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_121
timestamp 1608254825
transform 1 0 12236 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_43_115
timestamp 1608254825
transform 1 0 11684 0 1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_417
timestamp 1608254825
transform 1 0 12328 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_4  _1758_
timestamp 1608254825
transform 1 0 13524 0 1 25568
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _1332_
timestamp 1608254825
transform 1 0 12420 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_148
timestamp 1608254825
transform 1 0 14720 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_4  _1700_
timestamp 1608254825
transform 1 0 15088 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_179
timestamp 1608254825
transform 1 0 17572 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_164
timestamp 1608254825
transform 1 0 16192 0 1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__and3_4  _1419_
timestamp 1608254825
transform 1 0 16744 0 1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_43_200
timestamp 1608254825
transform 1 0 19504 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_196
timestamp 1608254825
transform 1 0 19136 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_418
timestamp 1608254825
transform 1 0 17940 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__a21o_4  _2230_
timestamp 1608254825
transform 1 0 18032 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__nand4_4  _1232_
timestamp 1608254825
transform 1 0 19596 0 1 25568
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_6  FILLER_43_218
timestamp 1608254825
transform 1 0 21160 0 1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_m1_clk_local
timestamp 1608254825
transform 1 0 21712 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_4  _2233_
timestamp 1608254825
transform 1 0 21988 0 1 25568
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_43_240
timestamp 1608254825
transform 1 0 23184 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_419
timestamp 1608254825
transform 1 0 23552 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__a21boi_4  _2232_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 23644 0 1 25568
box -38 -48 1418 592
use sky130_fd_sc_hd__fill_1  FILLER_43_274
timestamp 1608254825
transform 1 0 26312 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_43_268
timestamp 1608254825
transform 1 0 25760 0 1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_260
timestamp 1608254825
transform 1 0 25024 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1660_
timestamp 1608254825
transform 1 0 25392 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_294
timestamp 1608254825
transform 1 0 28152 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2592_
timestamp 1608254825
transform 1 0 26404 0 1 25568
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_43_314
timestamp 1608254825
transform 1 0 29992 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_306
timestamp 1608254825
transform 1 0 29256 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_301
timestamp 1608254825
transform 1 0 28796 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_420
timestamp 1608254825
transform 1 0 29164 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2645_
timestamp 1608254825
transform 1 0 30360 0 1 25568
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_2  _1662_
timestamp 1608254825
transform 1 0 28520 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1213_
timestamp 1608254825
transform 1 0 29624 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_337
timestamp 1608254825
transform 1 0 32108 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_4  _1216_
timestamp 1608254825
transform 1 0 32476 0 1 25568
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_43_362
timestamp 1608254825
transform 1 0 34408 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_355
timestamp 1608254825
transform 1 0 33764 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1841_
timestamp 1608254825
transform 1 0 34132 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_380
timestamp 1608254825
transform 1 0 36064 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_367
timestamp 1608254825
transform 1 0 34868 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_421
timestamp 1608254825
transform 1 0 34776 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2460_
timestamp 1608254825
transform 1 0 36432 0 1 25568
box -38 -48 1786 592
use sky130_fd_sc_hd__nand2_4  _1833_
timestamp 1608254825
transform 1 0 35236 0 1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_43_403
timestamp 1608254825
transform 1 0 38180 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1608254825
transform -1 0 38824 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_44_22
timestamp 1608254825
transform 1 0 3128 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1608254825
transform 1 0 1104 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _2473_
timestamp 1608254825
transform 1 0 1380 0 -1 26656
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_44_36
timestamp 1608254825
transform 1 0 4416 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_32
timestamp 1608254825
transform 1 0 4048 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_30
timestamp 1608254825
transform 1 0 3864 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_422
timestamp 1608254825
transform 1 0 3956 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2474_
timestamp 1608254825
transform 1 0 4508 0 -1 26656
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_44_64
timestamp 1608254825
transform 1 0 6992 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_44_56
timestamp 1608254825
transform 1 0 6256 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1391_
timestamp 1608254825
transform 1 0 7176 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_88
timestamp 1608254825
transform 1 0 9200 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_44_70
timestamp 1608254825
transform 1 0 7544 0 -1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_4  _1344_
timestamp 1608254825
transform 1 0 8096 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_104
timestamp 1608254825
transform 1 0 10672 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_93
timestamp 1608254825
transform 1 0 9660 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_423
timestamp 1608254825
transform 1 0 9568 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_4  _1336_
timestamp 1608254825
transform 1 0 9844 0 -1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__nand4_4  _1335_
timestamp 1608254825
transform 1 0 11040 0 -1 26656
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_1  FILLER_44_136
timestamp 1608254825
transform 1 0 13616 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_132
timestamp 1608254825
transform 1 0 13248 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_125
timestamp 1608254825
transform 1 0 12604 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_4  _2208_
timestamp 1608254825
transform 1 0 13708 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1241_
timestamp 1608254825
transform 1 0 12972 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_44_154
timestamp 1608254825
transform 1 0 15272 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_44_149
timestamp 1608254825
transform 1 0 14812 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_424
timestamp 1608254825
transform 1 0 15180 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_4  _2229_
timestamp 1608254825
transform 1 0 15548 0 -1 26656
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_44_170
timestamp 1608254825
transform 1 0 16744 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_4  _2187_
timestamp 1608254825
transform 1 0 17112 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_199
timestamp 1608254825
transform 1 0 19412 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_186
timestamp 1608254825
transform 1 0 18216 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_4  _1414_
timestamp 1608254825
transform 1 0 18584 0 -1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__or2_4  _1411_
timestamp 1608254825
transform 1 0 19780 0 -1 26656
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_44_224
timestamp 1608254825
transform 1 0 21712 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_210
timestamp 1608254825
transform 1 0 20424 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_425
timestamp 1608254825
transform 1 0 20792 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__o41ai_4  _2216_
timestamp 1608254825
transform 1 0 22080 0 -1 26656
box -38 -48 2062 592
use sky130_fd_sc_hd__and3_4  _1412_
timestamp 1608254825
transform 1 0 20884 0 -1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_44_250
timestamp 1608254825
transform 1 0 24104 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_271
timestamp 1608254825
transform 1 0 26036 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_263
timestamp 1608254825
transform 1 0 25300 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_4  _2168_
timestamp 1608254825
transform 1 0 24472 0 -1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _1672_
timestamp 1608254825
transform 1 0 25668 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_283
timestamp 1608254825
transform 1 0 27140 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_44_276
timestamp 1608254825
transform 1 0 26496 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_426
timestamp 1608254825
transform 1 0 26404 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_4  _2237_
timestamp 1608254825
transform 1 0 27508 0 -1 26656
box -38 -48 1234 592
use sky130_fd_sc_hd__buf_2  _1761_
timestamp 1608254825
transform 1 0 26772 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_317
timestamp 1608254825
transform 1 0 30268 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_313
timestamp 1608254825
transform 1 0 29900 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_300
timestamp 1608254825
transform 1 0 28704 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_4  _2214_
timestamp 1608254825
transform 1 0 29072 0 -1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_4  _1223_
timestamp 1608254825
transform 1 0 30360 0 -1 26656
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_1  FILLER_44_337
timestamp 1608254825
transform 1 0 32108 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_44_335
timestamp 1608254825
transform 1 0 31924 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_331
timestamp 1608254825
transform 1 0 31556 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_427
timestamp 1608254825
transform 1 0 32016 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_4  _1215_
timestamp 1608254825
transform 1 0 32200 0 -1 26656
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_44_359
timestamp 1608254825
transform 1 0 34132 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_351
timestamp 1608254825
transform 1 0 33396 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_4  _1840_
timestamp 1608254825
transform 1 0 34500 0 -1 26656
box -38 -48 1326 592
use sky130_fd_sc_hd__buf_2  _1188_
timestamp 1608254825
transform 1 0 33764 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_377
timestamp 1608254825
transform 1 0 35788 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_4  _1836_
timestamp 1608254825
transform 1 0 36156 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_401
timestamp 1608254825
transform 1 0 37996 0 -1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_44_393
timestamp 1608254825
transform 1 0 37260 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_428
timestamp 1608254825
transform 1 0 37628 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1608254825
transform -1 0 38824 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1834_
timestamp 1608254825
transform 1 0 37720 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_45_13
timestamp 1608254825
transform 1 0 2300 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_3
timestamp 1608254825
transform 1 0 1380 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1608254825
transform 1 0 1104 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__and3_4  _2084_
timestamp 1608254825
transform 1 0 1472 0 1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__nand4_4  _1991_
timestamp 1608254825
transform 1 0 2668 0 1 26656
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_45_34
timestamp 1608254825
transform 1 0 4232 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__and3_4  _2082_
timestamp 1608254825
transform 1 0 4600 0 1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_45_62
timestamp 1608254825
transform 1 0 6808 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_57
timestamp 1608254825
transform 1 0 6348 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_53
timestamp 1608254825
transform 1 0 5980 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_45_47
timestamp 1608254825
transform 1 0 5428 0 1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_429
timestamp 1608254825
transform 1 0 6716 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1345_
timestamp 1608254825
transform 1 0 6072 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1275_
timestamp 1608254825
transform 1 0 7176 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_84
timestamp 1608254825
transform 1 0 8832 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_45_78
timestamp 1608254825
transform 1 0 8280 0 1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_45_70
timestamp 1608254825
transform 1 0 7544 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2629_
timestamp 1608254825
transform 1 0 8924 0 1 26656
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  _1306_
timestamp 1608254825
transform 1 0 7912 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_108
timestamp 1608254825
transform 1 0 11040 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_104
timestamp 1608254825
transform 1 0 10672 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_4  _1239_
timestamp 1608254825
transform 1 0 11132 0 1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_45_136
timestamp 1608254825
transform 1 0 13616 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_118
timestamp 1608254825
transform 1 0 11960 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_430
timestamp 1608254825
transform 1 0 12328 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__nor3_4  _1258_
timestamp 1608254825
transform 1 0 12420 0 1 26656
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_6  FILLER_45_153
timestamp 1608254825
transform 1 0 15180 0 1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_4  _2231_
timestamp 1608254825
transform 1 0 15732 0 1 26656
box -38 -48 1234 592
use sky130_fd_sc_hd__a21oi_4  _1757_
timestamp 1608254825
transform 1 0 13984 0 1 26656
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_45_179
timestamp 1608254825
transform 1 0 17572 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_172
timestamp 1608254825
transform 1 0 16928 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1413_
timestamp 1608254825
transform 1 0 17296 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_45_191
timestamp 1608254825
transform 1 0 18676 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_431
timestamp 1608254825
transform 1 0 17940 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _1418_
timestamp 1608254825
transform 1 0 18032 0 1 26656
box -38 -48 682 592
use sky130_fd_sc_hd__nand3_4  _1409_
timestamp 1608254825
transform 1 0 19044 0 1 26656
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_45_209
timestamp 1608254825
transform 1 0 20332 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2615_
timestamp 1608254825
transform 1 0 20700 0 1 26656
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_45_245
timestamp 1608254825
transform 1 0 23644 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_45_243
timestamp 1608254825
transform 1 0 23460 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_239
timestamp 1608254825
transform 1 0 23092 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_232
timestamp 1608254825
transform 1 0 22448 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_432
timestamp 1608254825
transform 1 0 23552 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__or4_4  _1661_
timestamp 1608254825
transform 1 0 23828 0 1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1417_
timestamp 1608254825
transform 1 0 22816 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_45_256
timestamp 1608254825
transform 1 0 24656 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__a22oi_4  _2213_
timestamp 1608254825
transform 1 0 25024 0 1 26656
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_2  FILLER_45_285
timestamp 1608254825
transform 1 0 27324 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_45_277
timestamp 1608254825
transform 1 0 26588 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_4  _2215_
timestamp 1608254825
transform 1 0 27508 0 1 26656
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_45_309
timestamp 1608254825
transform 1 0 29532 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_304
timestamp 1608254825
transform 1 0 29072 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_300
timestamp 1608254825
transform 1 0 28704 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_433
timestamp 1608254825
transform 1 0 29164 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1734_
timestamp 1608254825
transform 1 0 29256 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_4  _1214_
timestamp 1608254825
transform 1 0 29900 0 1 26656
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_45_336
timestamp 1608254825
transform 1 0 32016 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_326
timestamp 1608254825
transform 1 0 31096 0 1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  _2646_
timestamp 1608254825
transform 1 0 32384 0 1 26656
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  _1187_
timestamp 1608254825
transform 1 0 31648 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_359
timestamp 1608254825
transform 1 0 34132 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_14_0_addressalyzerBlock.SPI_CLK
timestamp 1608254825
transform 1 0 34500 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_45_380
timestamp 1608254825
transform 1 0 36064 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_434
timestamp 1608254825
transform 1 0 34776 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2570_
timestamp 1608254825
transform 1 0 36432 0 1 26656
box -38 -48 1786 592
use sky130_fd_sc_hd__o21ai_4  _1835_
timestamp 1608254825
transform 1 0 34868 0 1 26656
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_45_403
timestamp 1608254825
transform 1 0 38180 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1608254825
transform -1 0 38824 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_47_10
timestamp 1608254825
transform 1 0 2024 0 1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_47_3
timestamp 1608254825
transform 1 0 1380 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_11
timestamp 1608254825
transform 1 0 2116 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_3
timestamp 1608254825
transform 1 0 1380 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1608254825
transform 1 0 1104 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1608254825
transform 1 0 1104 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_4  _2083_
timestamp 1608254825
transform 1 0 2208 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _2070_
timestamp 1608254825
transform 1 0 1748 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_4  _2053_
timestamp 1608254825
transform 1 0 2576 0 1 27744
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_47_29
timestamp 1608254825
transform 1 0 3772 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_30
timestamp 1608254825
transform 1 0 3864 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_46_24
timestamp 1608254825
transform 1 0 3312 0 -1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_435
timestamp 1608254825
transform 1 0 3956 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _2059_
timestamp 1608254825
transform 1 0 4048 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _2058_
timestamp 1608254825
transform 1 0 4140 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_41
timestamp 1608254825
transform 1 0 4876 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_37
timestamp 1608254825
transform 1 0 4508 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_43
timestamp 1608254825
transform 1 0 5060 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_36
timestamp 1608254825
transform 1 0 4416 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_4_0_m1_clk_local
timestamp 1608254825
transform 1 0 4784 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _2475_
timestamp 1608254825
transform 1 0 5152 0 -1 27744
box -38 -48 1786 592
use sky130_fd_sc_hd__o21ai_4  _2076_
timestamp 1608254825
transform 1 0 4968 0 1 27744
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_47_68
timestamp 1608254825
transform 1 0 7360 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_62
timestamp 1608254825
transform 1 0 6808 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_47_55
timestamp 1608254825
transform 1 0 6164 0 1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_46_63
timestamp 1608254825
transform 1 0 6900 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_m1_clk_local
timestamp 1608254825
transform 1 0 7268 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_442
timestamp 1608254825
transform 1 0 6716 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1298_
timestamp 1608254825
transform 1 0 6992 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_76
timestamp 1608254825
transform 1 0 8096 0 1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_46_86
timestamp 1608254825
transform 1 0 9016 0 -1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_46_70
timestamp 1608254825
transform 1 0 7544 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_6_0_m1_clk_local
timestamp 1608254825
transform 1 0 8648 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_4  _1353_
timestamp 1608254825
transform 1 0 8924 0 1 27744
box -38 -48 1326 592
use sky130_fd_sc_hd__nand3_4  _1347_
timestamp 1608254825
transform 1 0 7728 0 -1 27744
box -38 -48 1326 592
use sky130_fd_sc_hd__buf_2  _1269_
timestamp 1608254825
transform 1 0 7728 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_99
timestamp 1608254825
transform 1 0 10212 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_105
timestamp 1608254825
transform 1 0 10764 0 -1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_46_97
timestamp 1608254825
transform 1 0 10028 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_436
timestamp 1608254825
transform 1 0 9568 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_4  _1352_
timestamp 1608254825
transform 1 0 10580 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _1346_
timestamp 1608254825
transform 1 0 10396 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__nor4_4  _1333_
timestamp 1608254825
transform 1 0 11316 0 -1 27744
box -38 -48 1602 592
use sky130_fd_sc_hd__buf_2  _1324_
timestamp 1608254825
transform 1 0 9660 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_136
timestamp 1608254825
transform 1 0 13616 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_132
timestamp 1608254825
transform 1 0 13248 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_121
timestamp 1608254825
transform 1 0 12236 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_47_115
timestamp 1608254825
transform 1 0 11684 0 1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_46_128
timestamp 1608254825
transform 1 0 12880 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_443
timestamp 1608254825
transform 1 0 12328 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_4  _1658_
timestamp 1608254825
transform 1 0 13616 0 -1 27744
box -38 -48 1234 592
use sky130_fd_sc_hd__a21oi_4  _1657_
timestamp 1608254825
transform 1 0 13708 0 1 27744
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_4  _1240_
timestamp 1608254825
transform 1 0 12420 0 1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_47_150
timestamp 1608254825
transform 1 0 14904 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_149
timestamp 1608254825
transform 1 0 14812 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_437
timestamp 1608254825
transform 1 0 15180 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_4  _1859_
timestamp 1608254825
transform 1 0 15272 0 -1 27744
box -38 -48 1234 592
use sky130_fd_sc_hd__a21oi_4  _1721_
timestamp 1608254825
transform 1 0 15272 0 1 27744
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_8  FILLER_47_175
timestamp 1608254825
transform 1 0 17204 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_47_167
timestamp 1608254825
transform 1 0 16468 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_181
timestamp 1608254825
transform 1 0 17756 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_46_175
timestamp 1608254825
transform 1 0 17204 0 -1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_46_167
timestamp 1608254825
transform 1 0 16468 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2614_
timestamp 1608254825
transform 1 0 17848 0 -1 27744
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  _1656_
timestamp 1608254825
transform 1 0 16836 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1612_
timestamp 1608254825
transform 1 0 16836 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_197
timestamp 1608254825
transform 1 0 19228 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_46_201
timestamp 1608254825
transform 1 0 19596 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_444
timestamp 1608254825
transform 1 0 17940 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_4  _1415_
timestamp 1608254825
transform 1 0 18032 0 1 27744
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _1404_
timestamp 1608254825
transform 1 0 19964 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_4  _1401_
timestamp 1608254825
transform 1 0 19964 0 1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_47_221
timestamp 1608254825
transform 1 0 21436 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_47_214
timestamp 1608254825
transform 1 0 20792 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_208
timestamp 1608254825
transform 1 0 20240 0 -1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_438
timestamp 1608254825
transform 1 0 20792 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1410_
timestamp 1608254825
transform 1 0 21160 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__a41oi_4  _1407_
timestamp 1608254825
transform 1 0 20884 0 -1 27744
box -38 -48 2062 592
use sky130_fd_sc_hd__fill_1  FILLER_47_249
timestamp 1608254825
transform 1 0 24012 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_245
timestamp 1608254825
transform 1 0 23644 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_240
timestamp 1608254825
transform 1 0 23184 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_229
timestamp 1608254825
transform 1 0 22172 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_237
timestamp 1608254825
transform 1 0 22908 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_445
timestamp 1608254825
transform 1 0 23552 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__o41ai_4  _2147_
timestamp 1608254825
transform 1 0 23276 0 -1 27744
box -38 -48 2062 592
use sky130_fd_sc_hd__or4_4  _1860_
timestamp 1608254825
transform 1 0 22356 0 1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__nor4_4  _1673_
timestamp 1608254825
transform 1 0 24104 0 1 27744
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_1  FILLER_47_273
timestamp 1608254825
transform 1 0 26220 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_47_267
timestamp 1608254825
transform 1 0 25668 0 1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_46_271
timestamp 1608254825
transform 1 0 26036 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_263
timestamp 1608254825
transform 1 0 25300 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_12_0_addressalyzerBlock.SPI_CLK
timestamp 1608254825
transform 1 0 26312 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1675_
timestamp 1608254825
transform 1 0 25668 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_296
timestamp 1608254825
transform 1 0 28336 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_46_290
timestamp 1608254825
transform 1 0 27784 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_280
timestamp 1608254825
transform 1 0 26864 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_276
timestamp 1608254825
transform 1 0 26496 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_439
timestamp 1608254825
transform 1 0 26404 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2596_
timestamp 1608254825
transform 1 0 26588 0 1 27744
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _2436_
timestamp 1608254825
transform 1 0 28152 0 -1 27744
box -38 -48 1786 592
use sky130_fd_sc_hd__nand2_4  _1676_
timestamp 1608254825
transform 1 0 26956 0 -1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_47_313
timestamp 1608254825
transform 1 0 29900 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_304
timestamp 1608254825
transform 1 0 29072 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_313
timestamp 1608254825
transform 1 0 29900 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_446
timestamp 1608254825
transform 1 0 29164 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2652_
timestamp 1608254825
transform 1 0 30268 0 1 27744
box -38 -48 1786 592
use sky130_fd_sc_hd__o21ai_4  _2355_
timestamp 1608254825
transform 1 0 30268 0 -1 27744
box -38 -48 1234 592
use sky130_fd_sc_hd__or2_4  _2353_
timestamp 1608254825
transform 1 0 29256 0 1 27744
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_47_336
timestamp 1608254825
transform 1 0 32016 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_46_337
timestamp 1608254825
transform 1 0 32108 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_46_330
timestamp 1608254825
transform 1 0 31464 0 -1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_440
timestamp 1608254825
transform 1 0 32016 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_4  _2354_
timestamp 1608254825
transform 1 0 32384 0 1 27744
box -38 -48 1234 592
use sky130_fd_sc_hd__o21ai_4  _1211_
timestamp 1608254825
transform 1 0 32384 0 -1 27744
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_1  FILLER_47_365
timestamp 1608254825
transform 1 0 34684 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_361
timestamp 1608254825
transform 1 0 34316 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_353
timestamp 1608254825
transform 1 0 33580 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_361
timestamp 1608254825
transform 1 0 34316 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_353
timestamp 1608254825
transform 1 0 33580 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _2569_
timestamp 1608254825
transform 1 0 34408 0 -1 27744
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  _1181_
timestamp 1608254825
transform 1 0 33948 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_378
timestamp 1608254825
transform 1 0 35880 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_374
timestamp 1608254825
transform 1 0 35512 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_381
timestamp 1608254825
transform 1 0 36156 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_447
timestamp 1608254825
transform 1 0 34776 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__nand3_4  _1830_
timestamp 1608254825
transform 1 0 35972 0 1 27744
box -38 -48 1326 592
use sky130_fd_sc_hd__or2_4  _1210_
timestamp 1608254825
transform 1 0 36524 0 -1 27744
box -38 -48 682 592
use sky130_fd_sc_hd__or2_4  _1202_
timestamp 1608254825
transform 1 0 34868 0 1 27744
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_47_393
timestamp 1608254825
transform 1 0 37260 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_392
timestamp 1608254825
transform 1 0 37168 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_397
timestamp 1608254825
transform 1 0 37628 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_46_401
timestamp 1608254825
transform 1 0 37996 0 -1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_396
timestamp 1608254825
transform 1 0 37536 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_441
timestamp 1608254825
transform 1 0 37628 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _2362_
timestamp 1608254825
transform 1 0 37720 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1837_
timestamp 1608254825
transform 1 0 37720 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_47_406
timestamp 1608254825
transform 1 0 38456 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_402
timestamp 1608254825
transform 1 0 38088 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1608254825
transform -1 0 38824 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1608254825
transform -1 0 38824 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_48_22
timestamp 1608254825
transform 1 0 3128 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1608254825
transform 1 0 1104 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _2477_
timestamp 1608254825
transform 1 0 1380 0 -1 28832
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_48_45
timestamp 1608254825
transform 1 0 5244 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_30
timestamp 1608254825
transform 1 0 3864 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_448
timestamp 1608254825
transform 1 0 3956 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_4  _2069_
timestamp 1608254825
transform 1 0 4048 0 -1 28832
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_48_62
timestamp 1608254825
transform 1 0 6808 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_4  _2077_
timestamp 1608254825
transform 1 0 5612 0 -1 28832
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_4  _2072_
timestamp 1608254825
transform 1 0 7176 0 -1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_48_91
timestamp 1608254825
transform 1 0 9476 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_83
timestamp 1608254825
transform 1 0 8740 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_48_75
timestamp 1608254825
transform 1 0 8004 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1270_
timestamp 1608254825
transform 1 0 8372 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_102
timestamp 1608254825
transform 1 0 10488 0 -1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_449
timestamp 1608254825
transform 1 0 9568 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_4  _1354_
timestamp 1608254825
transform 1 0 9660 0 -1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__nor3_4  _1351_
timestamp 1608254825
transform 1 0 11040 0 -1 28832
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_48_121
timestamp 1608254825
transform 1 0 12236 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_4  _1357_
timestamp 1608254825
transform 1 0 12604 0 -1 28832
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_1  FILLER_48_154
timestamp 1608254825
transform 1 0 15272 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_145
timestamp 1608254825
transform 1 0 14444 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_48_138
timestamp 1608254825
transform 1 0 13800 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_450
timestamp 1608254825
transform 1 0 15180 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_4  _1722_
timestamp 1608254825
transform 1 0 15364 0 -1 28832
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _1356_
timestamp 1608254825
transform 1 0 14168 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_48_179
timestamp 1608254825
transform 1 0 17572 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_175
timestamp 1608254825
transform 1 0 17204 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_168
timestamp 1608254825
transform 1 0 16560 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_4  _1416_
timestamp 1608254825
transform 1 0 17664 0 -1 28832
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _1378_
timestamp 1608254825
transform 1 0 16928 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_48_193
timestamp 1608254825
transform 1 0 18860 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_4  _1408_
timestamp 1608254825
transform 1 0 19228 0 -1 28832
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_48_225
timestamp 1608254825
transform 1 0 21804 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_218
timestamp 1608254825
transform 1 0 21160 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_210
timestamp 1608254825
transform 1 0 20424 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_451
timestamp 1608254825
transform 1 0 20792 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1396_
timestamp 1608254825
transform 1 0 21528 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1230_
timestamp 1608254825
transform 1 0 20884 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_48_251
timestamp 1608254825
transform 1 0 24196 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_236
timestamp 1608254825
transform 1 0 22816 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_232
timestamp 1608254825
transform 1 0 22448 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_4  _1861_
timestamp 1608254825
transform 1 0 22908 0 -1 28832
box -38 -48 1326 592
use sky130_fd_sc_hd__inv_2  _1400_
timestamp 1608254825
transform 1 0 22172 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_48_269
timestamp 1608254825
transform 1 0 25852 0 -1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_4  _1674_
timestamp 1608254825
transform 1 0 24564 0 -1 28832
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_48_285
timestamp 1608254825
transform 1 0 27324 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_452
timestamp 1608254825
transform 1 0 26404 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _1739_
timestamp 1608254825
transform 1 0 27692 0 -1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  _1677_
timestamp 1608254825
transform 1 0 26496 0 -1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_48_311
timestamp 1608254825
transform 1 0 29716 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_48_298
timestamp 1608254825
transform 1 0 28520 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_4  _2356_
timestamp 1608254825
transform 1 0 30452 0 -1 28832
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_4  _2170_
timestamp 1608254825
transform 1 0 28888 0 -1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_48_337
timestamp 1608254825
transform 1 0 32108 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_332
timestamp 1608254825
transform 1 0 31648 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_453
timestamp 1608254825
transform 1 0 32016 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _1206_
timestamp 1608254825
transform 1 0 32476 0 -1 28832
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_48_365
timestamp 1608254825
transform 1 0 34684 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_348
timestamp 1608254825
transform 1 0 33120 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_4  _1205_
timestamp 1608254825
transform 1 0 33488 0 -1 28832
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_48_372
timestamp 1608254825
transform 1 0 35328 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__nand4_4  _1735_
timestamp 1608254825
transform 1 0 35696 0 -1 28832
box -38 -48 1602 592
use sky130_fd_sc_hd__inv_2  _1180_
timestamp 1608254825
transform 1 0 35052 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_48_406
timestamp 1608254825
transform 1 0 38456 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_402
timestamp 1608254825
transform 1 0 38088 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_393
timestamp 1608254825
transform 1 0 37260 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_454
timestamp 1608254825
transform 1 0 37628 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1608254825
transform -1 0 38824 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1178_
timestamp 1608254825
transform 1 0 37720 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_11
timestamp 1608254825
transform 1 0 2116 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_7
timestamp 1608254825
transform 1 0 1748 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_3
timestamp 1608254825
transform 1 0 1380 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1608254825
transform 1 0 1104 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__nor4_4  _1992_
timestamp 1608254825
transform 1 0 2484 0 1 28832
box -38 -48 1602 592
use sky130_fd_sc_hd__inv_2  _1988_
timestamp 1608254825
transform 1 0 1840 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_49_32
timestamp 1608254825
transform 1 0 4048 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_4  _2068_
timestamp 1608254825
transform 1 0 4416 0 1 28832
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_49_57
timestamp 1608254825
transform 1 0 6348 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_49
timestamp 1608254825
transform 1 0 5612 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_455
timestamp 1608254825
transform 1 0 6716 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _2027_
timestamp 1608254825
transform 1 0 5980 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_4  _1990_
timestamp 1608254825
transform 1 0 6808 0 1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_49_75
timestamp 1608254825
transform 1 0 8004 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_71
timestamp 1608254825
transform 1 0 7636 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2628_
timestamp 1608254825
transform 1 0 8096 0 1 28832
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_49_113
timestamp 1608254825
transform 1 0 11500 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_49_95
timestamp 1608254825
transform 1 0 9844 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_4  _1358_
timestamp 1608254825
transform 1 0 10212 0 1 28832
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_8  FILLER_49_132
timestamp 1608254825
transform 1 0 13248 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_121
timestamp 1608254825
transform 1 0 12236 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_456
timestamp 1608254825
transform 1 0 12328 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_4  _1228_
timestamp 1608254825
transform 1 0 12420 0 1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_49_159
timestamp 1608254825
transform 1 0 15732 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_155
timestamp 1608254825
transform 1 0 15364 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_140
timestamp 1608254825
transform 1 0 13984 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__a21oi_4  _1858_
timestamp 1608254825
transform 1 0 14168 0 1 28832
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_49_179
timestamp 1608254825
transform 1 0 17572 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2624_
timestamp 1608254825
transform 1 0 15824 0 1 28832
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_49_198
timestamp 1608254825
transform 1 0 19320 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_184
timestamp 1608254825
transform 1 0 18032 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_457
timestamp 1608254825
transform 1 0 17940 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_4  _1403_
timestamp 1608254825
transform 1 0 18124 0 1 28832
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_49_226
timestamp 1608254825
transform 1 0 21896 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_206
timestamp 1608254825
transform 1 0 20056 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2616_
timestamp 1608254825
transform 1 0 20148 0 1 28832
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_49_248
timestamp 1608254825
transform 1 0 23920 0 1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_243
timestamp 1608254825
transform 1 0 23460 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_239
timestamp 1608254825
transform 1 0 23092 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_458
timestamp 1608254825
transform 1 0 23552 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_4  _2166_
timestamp 1608254825
transform 1 0 22264 0 1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _2146_
timestamp 1608254825
transform 1 0 23644 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_49_272
timestamp 1608254825
transform 1 0 26128 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_254
timestamp 1608254825
transform 1 0 24472 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__a22oi_4  _2191_
timestamp 1608254825
transform 1 0 24564 0 1 28832
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_6  FILLER_49_296
timestamp 1608254825
transform 1 0 28336 0 1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_addressalyzerBlock.SPI_CLK
timestamp 1608254825
transform 1 0 26864 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_4  _2193_
timestamp 1608254825
transform 1 0 27140 0 1 28832
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_6  FILLER_49_306
timestamp 1608254825
transform 1 0 29256 0 1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_addressalyzerBlock.SPI_CLK
timestamp 1608254825
transform 1 0 28888 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_459
timestamp 1608254825
transform 1 0 29164 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_4  _1208_
timestamp 1608254825
transform 1 0 29808 0 1 28832
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_49_325
timestamp 1608254825
transform 1 0 31004 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2647_
timestamp 1608254825
transform 1 0 31372 0 1 28832
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_49_362
timestamp 1608254825
transform 1 0 34408 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_354
timestamp 1608254825
transform 1 0 33672 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_49_348
timestamp 1608254825
transform 1 0 33120 0 1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__or2_4  _1198_
timestamp 1608254825
transform 1 0 33764 0 1 28832
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_49_383
timestamp 1608254825
transform 1 0 36340 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_379
timestamp 1608254825
transform 1 0 35972 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_460
timestamp 1608254825
transform 1 0 34776 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2571_
timestamp 1608254825
transform 1 0 36432 0 1 28832
box -38 -48 1786 592
use sky130_fd_sc_hd__o21a_4  _1842_
timestamp 1608254825
transform 1 0 34868 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_403
timestamp 1608254825
transform 1 0 38180 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1608254825
transform -1 0 38824 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_50_15
timestamp 1608254825
transform 1 0 2484 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_11
timestamp 1608254825
transform 1 0 2116 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_3
timestamp 1608254825
transform 1 0 1380 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1608254825
transform 1 0 1104 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _2054_
timestamp 1608254825
transform 1 0 2852 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1989_
timestamp 1608254825
transform 1 0 2208 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_50_45
timestamp 1608254825
transform 1 0 5244 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_41
timestamp 1608254825
transform 1 0 4876 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_50_23
timestamp 1608254825
transform 1 0 3220 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_461
timestamp 1608254825
transform 1 0 3956 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _2060_
timestamp 1608254825
transform 1 0 4048 0 -1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_50_65
timestamp 1608254825
transform 1 0 7084 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2476_
timestamp 1608254825
transform 1 0 5336 0 -1 29920
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_50_88
timestamp 1608254825
transform 1 0 9200 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_81
timestamp 1608254825
transform 1 0 8556 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_4  _2074_
timestamp 1608254825
transform 1 0 7452 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1253_
timestamp 1608254825
transform 1 0 8924 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_50_105
timestamp 1608254825
transform 1 0 10764 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_50_97
timestamp 1608254825
transform 1 0 10028 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_462
timestamp 1608254825
transform 1 0 9568 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1374_
timestamp 1608254825
transform 1 0 10396 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_4  _1362_
timestamp 1608254825
transform 1 0 11500 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _1283_
timestamp 1608254825
transform 1 0 9660 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_125
timestamp 1608254825
transform 1 0 12604 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2626_
timestamp 1608254825
transform 1 0 12972 0 -1 29920
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_50_157
timestamp 1608254825
transform 1 0 15548 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_152
timestamp 1608254825
transform 1 0 15088 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_148
timestamp 1608254825
transform 1 0 14720 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_463
timestamp 1608254825
transform 1 0 15180 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1369_
timestamp 1608254825
transform 1 0 15272 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_50_175
timestamp 1608254825
transform 1 0 17204 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__nand3_4  _1376_
timestamp 1608254825
transform 1 0 15916 0 -1 29920
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_50_203
timestamp 1608254825
transform 1 0 19780 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_183
timestamp 1608254825
transform 1 0 17940 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2617_
timestamp 1608254825
transform 1 0 18032 0 -1 29920
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_50_215
timestamp 1608254825
transform 1 0 20884 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_210
timestamp 1608254825
transform 1 0 20424 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_464
timestamp 1608254825
transform 1 0 20792 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__a21o_4  _1725_
timestamp 1608254825
transform 1 0 21252 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1235_
timestamp 1608254825
transform 1 0 20148 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_50_248
timestamp 1608254825
transform 1 0 23920 0 -1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_50_231
timestamp 1608254825
transform 1 0 22356 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_4  _1723_
timestamp 1608254825
transform 1 0 22724 0 -1 29920
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_50_271
timestamp 1608254825
transform 1 0 26036 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__a22oi_4  _2169_
timestamp 1608254825
transform 1 0 24472 0 -1 29920
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_50_286
timestamp 1608254825
transform 1 0 27416 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_276
timestamp 1608254825
transform 1 0 26496 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_465
timestamp 1608254825
transform 1 0 26404 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2437_
timestamp 1608254825
transform 1 0 27784 0 -1 29920
box -38 -48 1786 592
use sky130_fd_sc_hd__nand2_4  _2192_
timestamp 1608254825
transform 1 0 26588 0 -1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_50_309
timestamp 1608254825
transform 1 0 29532 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_4  _1204_
timestamp 1608254825
transform 1 0 29900 0 -1 29920
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_2  FILLER_50_337
timestamp 1608254825
transform 1 0 32108 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_50_333
timestamp 1608254825
transform 1 0 31740 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_50_326
timestamp 1608254825
transform 1 0 31096 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_addressalyzerBlock.SPI_CLK
timestamp 1608254825
transform 1 0 31464 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_466
timestamp 1608254825
transform 1 0 32016 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_4  _1207_
timestamp 1608254825
transform 1 0 32292 0 -1 29920
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_50_352
timestamp 1608254825
transform 1 0 33488 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2648_
timestamp 1608254825
transform 1 0 33856 0 -1 29920
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_50_379
timestamp 1608254825
transform 1 0 35972 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_375
timestamp 1608254825
transform 1 0 35604 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_4  _1832_
timestamp 1608254825
transform 1 0 36064 0 -1 29920
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_1  FILLER_50_406
timestamp 1608254825
transform 1 0 38456 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_402
timestamp 1608254825
transform 1 0 38088 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_393
timestamp 1608254825
transform 1 0 37260 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_467
timestamp 1608254825
transform 1 0 37628 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1608254825
transform -1 0 38824 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1179_
timestamp 1608254825
transform 1 0 37720 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_22
timestamp 1608254825
transform 1 0 3128 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1608254825
transform 1 0 1104 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _2478_
timestamp 1608254825
transform 1 0 1380 0 1 29920
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_51_39
timestamp 1608254825
transform 1 0 4692 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_m1_clk_local
timestamp 1608254825
transform 1 0 5060 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_4  _2066_
timestamp 1608254825
transform 1 0 3496 0 1 29920
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_51_57
timestamp 1608254825
transform 1 0 6348 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_49
timestamp 1608254825
transform 1 0 5612 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_468
timestamp 1608254825
transform 1 0 6716 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_4  _2073_
timestamp 1608254825
transform 1 0 6808 0 1 29920
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _2071_
timestamp 1608254825
transform 1 0 5336 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1388_
timestamp 1608254825
transform 1 0 5980 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_83
timestamp 1608254825
transform 1 0 8740 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_75
timestamp 1608254825
transform 1 0 8004 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_m1_clk_local
timestamp 1608254825
transform 1 0 9108 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _2627_
timestamp 1608254825
transform 1 0 9384 0 1 29920
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  _1274_
timestamp 1608254825
transform 1 0 8372 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_109
timestamp 1608254825
transform 1 0 11132 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1349_
timestamp 1608254825
transform 1 0 11500 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_51_132
timestamp 1608254825
transform 1 0 13248 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_51_116
timestamp 1608254825
transform 1 0 11776 0 1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_469
timestamp 1608254825
transform 1 0 12328 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__nand4_4  _1367_
timestamp 1608254825
transform 1 0 13616 0 1 29920
box -38 -48 1602 592
use sky130_fd_sc_hd__nor2_4  _1361_
timestamp 1608254825
transform 1 0 12420 0 1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_51_153
timestamp 1608254825
transform 1 0 15180 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1372_
timestamp 1608254825
transform 1 0 15548 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_179
timestamp 1608254825
transform 1 0 17572 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_51_161
timestamp 1608254825
transform 1 0 15916 0 1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_4  _1375_
timestamp 1608254825
transform 1 0 16468 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_51_203
timestamp 1608254825
transform 1 0 19780 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_199
timestamp 1608254825
transform 1 0 19412 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_51_184
timestamp 1608254825
transform 1 0 18032 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_470
timestamp 1608254825
transform 1 0 17940 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_4  _1402_
timestamp 1608254825
transform 1 0 18216 0 1 29920
box -38 -48 1234 592
use sky130_fd_sc_hd__nor3_4  _1363_
timestamp 1608254825
transform 1 0 19872 0 1 29920
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_8  FILLER_51_217
timestamp 1608254825
transform 1 0 21068 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_4  _2167_
timestamp 1608254825
transform 1 0 21804 0 1 29920
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_6  FILLER_51_238
timestamp 1608254825
transform 1 0 23000 0 1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_471
timestamp 1608254825
transform 1 0 23552 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_4  _1759_
timestamp 1608254825
transform 1 0 23644 0 1 29920
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_1  FILLER_51_262
timestamp 1608254825
transform 1 0 25208 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_258
timestamp 1608254825
transform 1 0 24840 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2593_
timestamp 1608254825
transform 1 0 25300 0 1 29920
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_51_282
timestamp 1608254825
transform 1 0 27048 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_4  _2171_
timestamp 1608254825
transform 1 0 27416 0 1 29920
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_8  FILLER_51_315
timestamp 1608254825
transform 1 0 30084 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_51_299
timestamp 1608254825
transform 1 0 28612 0 1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_472
timestamp 1608254825
transform 1 0 29164 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_4  _1862_
timestamp 1608254825
transform 1 0 29256 0 1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_51_339
timestamp 1608254825
transform 1 0 32292 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_51_323
timestamp 1608254825
transform 1 0 30820 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_4  _1209_
timestamp 1608254825
transform 1 0 31096 0 1 29920
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_51_362
timestamp 1608254825
transform 1 0 34408 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_51_346
timestamp 1608254825
transform 1 0 32936 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_15_0_addressalyzerBlock.SPI_CLK
timestamp 1608254825
transform 1 0 32660 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_4  _1203_
timestamp 1608254825
transform 1 0 33212 0 1 29920
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_51_380
timestamp 1608254825
transform 1 0 36064 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_367
timestamp 1608254825
transform 1 0 34868 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_473
timestamp 1608254825
transform 1 0 34776 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2455_
timestamp 1608254825
transform 1 0 36432 0 1 29920
box -38 -48 1786 592
use sky130_fd_sc_hd__nand2_4  _1831_
timestamp 1608254825
transform 1 0 35236 0 1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_51_403
timestamp 1608254825
transform 1 0 38180 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1608254825
transform -1 0 38824 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_53_14
timestamp 1608254825
transform 1 0 2392 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_53_3
timestamp 1608254825
transform 1 0 1380 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_11
timestamp 1608254825
transform 1 0 2116 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_52_3
timestamp 1608254825
transform 1 0 1380 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1608254825
transform 1 0 1104 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1608254825
transform 1 0 1104 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_4  _2067_
timestamp 1608254825
transform 1 0 2300 0 -1 31008
box -38 -48 1234 592
use sky130_fd_sc_hd__and4_4  _2062_
timestamp 1608254825
transform 1 0 1564 0 1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__a41oi_4  _2061_
timestamp 1608254825
transform 1 0 2760 0 1 31008
box -38 -48 2062 592
use sky130_fd_sc_hd__decap_8  FILLER_53_40
timestamp 1608254825
transform 1 0 4784 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_52_45
timestamp 1608254825
transform 1 0 5244 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_52_40
timestamp 1608254825
transform 1 0 4784 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_52_32
timestamp 1608254825
transform 1 0 4048 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_30
timestamp 1608254825
transform 1 0 3864 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_26
timestamp 1608254825
transform 1 0 3496 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_474
timestamp 1608254825
transform 1 0 3956 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _2075_
timestamp 1608254825
transform 1 0 4968 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_53_62
timestamp 1608254825
transform 1 0 6808 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_57
timestamp 1608254825
transform 1 0 6348 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_52_52
timestamp 1608254825
transform 1 0 5888 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_481
timestamp 1608254825
transform 1 0 6716 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _2039_
timestamp 1608254825
transform 1 0 5612 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_4  _2038_
timestamp 1608254825
transform 1 0 5520 0 1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1996_
timestamp 1608254825
transform 1 0 7176 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_4  _1995_
timestamp 1608254825
transform 1 0 6624 0 -1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_53_69
timestamp 1608254825
transform 1 0 7452 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_91
timestamp 1608254825
transform 1 0 9476 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_52_85
timestamp 1608254825
transform 1 0 8924 0 -1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_52_69
timestamp 1608254825
transform 1 0 7452 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2487_
timestamp 1608254825
transform 1 0 7820 0 1 31008
box -38 -48 1786 592
use sky130_fd_sc_hd__o21a_4  _2034_
timestamp 1608254825
transform 1 0 7820 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_99
timestamp 1608254825
transform 1 0 10212 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_92
timestamp 1608254825
transform 1 0 9568 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_96
timestamp 1608254825
transform 1 0 9936 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_475
timestamp 1608254825
transform 1 0 9568 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1359_
timestamp 1608254825
transform 1 0 9936 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1355_
timestamp 1608254825
transform 1 0 10304 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1348_
timestamp 1608254825
transform 1 0 9660 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_52_103
timestamp 1608254825
transform 1 0 10580 0 -1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  _2625_
timestamp 1608254825
transform 1 0 11132 0 -1 31008
box -38 -48 1786 592
use sky130_fd_sc_hd__o21ai_4  _1370_
timestamp 1608254825
transform 1 0 10580 0 1 31008
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_8  FILLER_53_127
timestamp 1608254825
transform 1 0 12788 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_53_116
timestamp 1608254825
transform 1 0 11776 0 1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_52_128
timestamp 1608254825
transform 1 0 12880 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_482
timestamp 1608254825
transform 1 0 12328 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2623_
timestamp 1608254825
transform 1 0 13524 0 1 31008
box -38 -48 1786 592
use sky130_fd_sc_hd__nand2_4  _1368_
timestamp 1608254825
transform 1 0 13248 0 -1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _1350_
timestamp 1608254825
transform 1 0 12420 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_154
timestamp 1608254825
transform 1 0 15272 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_154
timestamp 1608254825
transform 1 0 15272 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_149
timestamp 1608254825
transform 1 0 14812 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_145
timestamp 1608254825
transform 1 0 14444 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_141
timestamp 1608254825
transform 1 0 14076 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_476
timestamp 1608254825
transform 1 0 15180 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__nand4_4  _1238_
timestamp 1608254825
transform 1 0 15640 0 1 31008
box -38 -48 1602 592
use sky130_fd_sc_hd__inv_2  _1237_
timestamp 1608254825
transform 1 0 14536 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_4  _1236_
timestamp 1608254825
transform 1 0 15364 0 -1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_53_175
timestamp 1608254825
transform 1 0 17204 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_52_179
timestamp 1608254825
transform 1 0 17572 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_52_164
timestamp 1608254825
transform 1 0 16192 0 -1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__and4_4  _1373_
timestamp 1608254825
transform 1 0 16744 0 -1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_53_197
timestamp 1608254825
transform 1 0 19228 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_193
timestamp 1608254825
transform 1 0 18860 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_200
timestamp 1608254825
transform 1 0 19504 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_192
timestamp 1608254825
transform 1 0 18768 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_483
timestamp 1608254825
transform 1 0 17940 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_4  _1377_
timestamp 1608254825
transform 1 0 17940 0 -1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  _1234_
timestamp 1608254825
transform 1 0 18032 0 1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__nor4_4  _1233_
timestamp 1608254825
transform 1 0 19320 0 1 31008
box -38 -48 1602 592
use sky130_fd_sc_hd__nand2_4  _1231_
timestamp 1608254825
transform 1 0 19596 0 -1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_53_215
timestamp 1608254825
transform 1 0 20884 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_226
timestamp 1608254825
transform 1 0 21896 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_218
timestamp 1608254825
transform 1 0 21160 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_52_210
timestamp 1608254825
transform 1 0 20424 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_477
timestamp 1608254825
transform 1 0 20792 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2618_
timestamp 1608254825
transform 1 0 21988 0 -1 31008
box -38 -48 1786 592
use sky130_fd_sc_hd__nor3_4  _1397_
timestamp 1608254825
transform 1 0 21252 0 1 31008
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _1229_
timestamp 1608254825
transform 1 0 20884 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_53_245
timestamp 1608254825
transform 1 0 23644 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_240
timestamp 1608254825
transform 1 0 23184 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_232
timestamp 1608254825
transform 1 0 22448 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_246
timestamp 1608254825
transform 1 0 23736 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_484
timestamp 1608254825
transform 1 0 23552 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__or3_4  _2352_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 24012 0 1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _1898_
timestamp 1608254825
transform 1 0 22816 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_4  _1760_
timestamp 1608254825
transform 1 0 24104 0 -1 31008
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_53_271
timestamp 1608254825
transform 1 0 26036 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_258
timestamp 1608254825
transform 1 0 24840 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_271
timestamp 1608254825
transform 1 0 26036 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_267
timestamp 1608254825
transform 1 0 25668 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_263
timestamp 1608254825
transform 1 0 25300 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1740_
timestamp 1608254825
transform 1 0 25760 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_4  _1727_
timestamp 1608254825
transform 1 0 25208 0 1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_53_278
timestamp 1608254825
transform 1 0 26680 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_52_285
timestamp 1608254825
transform 1 0 27324 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_13_0_addressalyzerBlock.SPI_CLK
timestamp 1608254825
transform 1 0 26404 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_478
timestamp 1608254825
transform 1 0 26404 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2590_
timestamp 1608254825
transform 1 0 26956 0 1 31008
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _2438_
timestamp 1608254825
transform 1 0 27692 0 -1 31008
box -38 -48 1786 592
use sky130_fd_sc_hd__nand2_4  _1726_
timestamp 1608254825
transform 1 0 26496 0 -1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_53_306
timestamp 1608254825
transform 1 0 29256 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_53_304
timestamp 1608254825
transform 1 0 29072 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_300
timestamp 1608254825
transform 1 0 28704 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_308
timestamp 1608254825
transform 1 0 29440 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_485
timestamp 1608254825
transform 1 0 29164 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_4  _1200_
timestamp 1608254825
transform 1 0 29440 0 1 31008
box -38 -48 1234 592
use sky130_fd_sc_hd__o21ai_4  _1192_
timestamp 1608254825
transform 1 0 29808 0 -1 31008
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_53_321
timestamp 1608254825
transform 1 0 30636 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_337
timestamp 1608254825
transform 1 0 32108 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_52_333
timestamp 1608254825
transform 1 0 31740 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_52_325
timestamp 1608254825
transform 1 0 31004 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_479
timestamp 1608254825
transform 1 0 32016 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2651_
timestamp 1608254825
transform 1 0 31004 0 1 31008
box -38 -48 1786 592
use sky130_fd_sc_hd__and2_4  _2109_
timestamp 1608254825
transform 1 0 32476 0 -1 31008
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_53_365
timestamp 1608254825
transform 1 0 34684 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_361
timestamp 1608254825
transform 1 0 34316 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_344
timestamp 1608254825
transform 1 0 32752 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_52_365
timestamp 1608254825
transform 1 0 34684 0 -1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_52_348
timestamp 1608254825
transform 1 0 33120 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_4  _1201_
timestamp 1608254825
transform 1 0 33488 0 -1 31008
box -38 -48 1234 592
use sky130_fd_sc_hd__o21ai_4  _1183_
timestamp 1608254825
transform 1 0 33120 0 1 31008
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_53_380
timestamp 1608254825
transform 1 0 36064 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_371
timestamp 1608254825
transform 1 0 35236 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_486
timestamp 1608254825
transform 1 0 34776 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2467_
timestamp 1608254825
transform 1 0 35328 0 -1 31008
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _2454_
timestamp 1608254825
transform 1 0 36432 0 1 31008
box -38 -48 1786 592
use sky130_fd_sc_hd__o21ai_4  _1199_
timestamp 1608254825
transform 1 0 34868 0 1 31008
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_53_403
timestamp 1608254825
transform 1 0 38180 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_52_401
timestamp 1608254825
transform 1 0 37996 0 -1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_52_391
timestamp 1608254825
transform 1 0 37076 0 -1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_480
timestamp 1608254825
transform 1 0 37628 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1608254825
transform -1 0 38824 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1608254825
transform -1 0 38824 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1829_
timestamp 1608254825
transform 1 0 37720 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_54_22
timestamp 1608254825
transform 1 0 3128 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1608254825
transform 1 0 1104 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _2480_
timestamp 1608254825
transform 1 0 1380 0 -1 32096
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_54_43
timestamp 1608254825
transform 1 0 5060 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_39
timestamp 1608254825
transform 1 0 4692 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_32
timestamp 1608254825
transform 1 0 4048 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_30
timestamp 1608254825
transform 1 0 3864 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_5_0_m1_clk_local
timestamp 1608254825
transform 1 0 4416 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_487
timestamp 1608254825
transform 1 0 3956 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2486_
timestamp 1608254825
transform 1 0 5152 0 -1 32096
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_54_63
timestamp 1608254825
transform 1 0 6900 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__nand4_4  _2037_
timestamp 1608254825
transform 1 0 7268 0 -1 32096
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_1  FILLER_54_91
timestamp 1608254825
transform 1 0 9476 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_84
timestamp 1608254825
transform 1 0 8832 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_7_0_m1_clk_local
timestamp 1608254825
transform 1 0 9200 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_54_102
timestamp 1608254825
transform 1 0 10488 0 -1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_488
timestamp 1608254825
transform 1 0 9568 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__and3_4  _2028_
timestamp 1608254825
transform 1 0 9660 0 -1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_4  _1371_
timestamp 1608254825
transform 1 0 11040 0 -1 32096
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_1  FILLER_54_136
timestamp 1608254825
transform 1 0 13616 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_128
timestamp 1608254825
transform 1 0 12880 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_54_121
timestamp 1608254825
transform 1 0 12236 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_4  _1382_
timestamp 1608254825
transform 1 0 13708 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1360_
timestamp 1608254825
transform 1 0 12604 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_54_149
timestamp 1608254825
transform 1 0 14812 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_489
timestamp 1608254825
transform 1 0 15180 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_4  _1392_
timestamp 1608254825
transform 1 0 15272 0 -1 32096
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_8  FILLER_54_175
timestamp 1608254825
transform 1 0 17204 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_54_167
timestamp 1608254825
transform 1 0 16468 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1364_
timestamp 1608254825
transform 1 0 16836 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_200
timestamp 1608254825
transform 1 0 19504 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_192
timestamp 1608254825
transform 1 0 18768 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_4  _1394_
timestamp 1608254825
transform 1 0 19596 0 -1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__and4_4  _1365_
timestamp 1608254825
transform 1 0 17940 0 -1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_54_215
timestamp 1608254825
transform 1 0 20884 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_210
timestamp 1608254825
transform 1 0 20424 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_490
timestamp 1608254825
transform 1 0 20792 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_4  _1398_
timestamp 1608254825
transform 1 0 21252 0 -1 32096
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_54_242
timestamp 1608254825
transform 1 0 23368 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_54_232
timestamp 1608254825
transform 1 0 22448 0 -1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  _2545_
timestamp 1608254825
transform 1 0 23736 0 -1 32096
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  _1892_
timestamp 1608254825
transform 1 0 23000 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_54_273
timestamp 1608254825
transform 1 0 26220 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_54_265
timestamp 1608254825
transform 1 0 25484 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_54_289
timestamp 1608254825
transform 1 0 27692 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_491
timestamp 1608254825
transform 1 0 26404 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2568_
timestamp 1608254825
transform 1 0 28060 0 -1 32096
box -38 -48 1786 592
use sky130_fd_sc_hd__o21ai_4  _1763_
timestamp 1608254825
transform 1 0 26496 0 -1 32096
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_1  FILLER_54_318
timestamp 1608254825
transform 1 0 30360 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_54_312
timestamp 1608254825
transform 1 0 29808 0 -1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_4  _1193_
timestamp 1608254825
transform 1 0 30452 0 -1 32096
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_1  FILLER_54_341
timestamp 1608254825
transform 1 0 32476 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_337
timestamp 1608254825
transform 1 0 32108 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_332
timestamp 1608254825
transform 1 0 31648 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_492
timestamp 1608254825
transform 1 0 32016 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _1182_
timestamp 1608254825
transform 1 0 32568 0 -1 32096
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_54_349
timestamp 1608254825
transform 1 0 33212 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2649_
timestamp 1608254825
transform 1 0 33580 0 -1 32096
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_54_383
timestamp 1608254825
transform 1 0 36340 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_372
timestamp 1608254825
transform 1 0 35328 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__and2_4  _2094_
timestamp 1608254825
transform 1 0 35696 0 -1 32096
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _2091_
timestamp 1608254825
transform 1 0 36708 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_54_401
timestamp 1608254825
transform 1 0 37996 0 -1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_396
timestamp 1608254825
transform 1 0 37536 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_54_390
timestamp 1608254825
transform 1 0 36984 0 -1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_493
timestamp 1608254825
transform 1 0 37628 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1608254825
transform -1 0 38824 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2098_
timestamp 1608254825
transform 1 0 37720 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_55_16
timestamp 1608254825
transform 1 0 2576 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1608254825
transform 1 0 1104 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__a41oi_4  _2064_
timestamp 1608254825
transform 1 0 2944 0 1 32096
box -38 -48 2062 592
use sky130_fd_sc_hd__nor3_4  _2063_
timestamp 1608254825
transform 1 0 1380 0 1 32096
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_6  FILLER_55_42
timestamp 1608254825
transform 1 0 4968 0 1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_55_68
timestamp 1608254825
transform 1 0 7360 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_55_62
timestamp 1608254825
transform 1 0 6808 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_57
timestamp 1608254825
transform 1 0 6348 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_494
timestamp 1608254825
transform 1 0 6716 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__and4_4  _2035_
timestamp 1608254825
transform 1 0 5520 0 1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _2031_
timestamp 1608254825
transform 1 0 6992 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__a41oi_4  _2033_
timestamp 1608254825
transform 1 0 7728 0 1 32096
box -38 -48 2062 592
use sky130_fd_sc_hd__decap_8  FILLER_55_94
timestamp 1608254825
transform 1 0 9752 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_4  _2024_
timestamp 1608254825
transform 1 0 10488 0 1 32096
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_6  FILLER_55_136
timestamp 1608254825
transform 1 0 13616 0 1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_121
timestamp 1608254825
transform 1 0 12236 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_55_115
timestamp 1608254825
transform 1 0 11684 0 1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_495
timestamp 1608254825
transform 1 0 12328 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_4  _2025_
timestamp 1608254825
transform 1 0 12420 0 1 32096
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_1  FILLER_55_142
timestamp 1608254825
transform 1 0 14168 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__a41oi_4  _1381_
timestamp 1608254825
transform 1 0 14260 0 1 32096
box -38 -48 2062 592
use sky130_fd_sc_hd__decap_4  FILLER_55_179
timestamp 1608254825
transform 1 0 17572 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_169
timestamp 1608254825
transform 1 0 16652 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_165
timestamp 1608254825
transform 1 0 16284 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__and4_4  _1383_
timestamp 1608254825
transform 1 0 16744 0 1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_55_196
timestamp 1608254825
transform 1 0 19136 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_496
timestamp 1608254825
transform 1 0 17940 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__nor3_4  _1395_
timestamp 1608254825
transform 1 0 19504 0 1 32096
box -38 -48 1234 592
use sky130_fd_sc_hd__o21a_4  _1384_
timestamp 1608254825
transform 1 0 18032 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_55_221
timestamp 1608254825
transform 1 0 21436 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_213
timestamp 1608254825
transform 1 0 20700 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_4  _1399_
timestamp 1608254825
transform 1 0 21528 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_55_242
timestamp 1608254825
transform 1 0 23368 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_55_234
timestamp 1608254825
transform 1 0 22632 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_497
timestamp 1608254825
transform 1 0 23552 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _1897_
timestamp 1608254825
transform 1 0 23644 0 1 32096
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_55_266
timestamp 1608254825
transform 1 0 25576 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_256
timestamp 1608254825
transform 1 0 24656 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_252
timestamp 1608254825
transform 1 0 24288 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2466_
timestamp 1608254825
transform 1 0 25944 0 1 32096
box -38 -48 1786 592
use sky130_fd_sc_hd__or3_4  _2351_
timestamp 1608254825
transform 1 0 24748 0 1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_55_293
timestamp 1608254825
transform 1 0 28060 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_289
timestamp 1608254825
transform 1 0 27692 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__and2_4  _2110_
timestamp 1608254825
transform 1 0 28152 0 1 32096
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_55_306
timestamp 1608254825
transform 1 0 29256 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_301
timestamp 1608254825
transform 1 0 28796 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_498
timestamp 1608254825
transform 1 0 29164 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_4  _1196_
timestamp 1608254825
transform 1 0 29624 0 1 32096
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_55_323
timestamp 1608254825
transform 1 0 30820 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2650_
timestamp 1608254825
transform 1 0 31188 0 1 32096
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_55_362
timestamp 1608254825
transform 1 0 34408 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_354
timestamp 1608254825
transform 1 0 33672 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_346
timestamp 1608254825
transform 1 0 32936 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__or2_4  _1194_
timestamp 1608254825
transform 1 0 33764 0 1 32096
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_55_373
timestamp 1608254825
transform 1 0 35420 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_55_367
timestamp 1608254825
transform 1 0 34868 0 1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_499
timestamp 1608254825
transform 1 0 34776 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2465_
timestamp 1608254825
transform 1 0 35512 0 1 32096
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_55_406
timestamp 1608254825
transform 1 0 38456 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_55_400
timestamp 1608254825
transform 1 0 37904 0 1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_55_393
timestamp 1608254825
transform 1 0 37260 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1608254825
transform -1 0 38824 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2103_
timestamp 1608254825
transform 1 0 37628 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_56_9
timestamp 1608254825
transform 1 0 1932 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_56_3
timestamp 1608254825
transform 1 0 1380 0 -1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1608254825
transform 1 0 1104 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__a41o_4  _2056_
timestamp 1608254825
transform 1 0 2024 0 -1 33184
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_56_44
timestamp 1608254825
transform 1 0 5152 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_27
timestamp 1608254825
transform 1 0 3588 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_500
timestamp 1608254825
transform 1 0 3956 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_4  _2065_
timestamp 1608254825
transform 1 0 4048 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_67
timestamp 1608254825
transform 1 0 7268 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_51
timestamp 1608254825
transform 1 0 5796 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2041_
timestamp 1608254825
transform 1 0 5520 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_4  _2036_
timestamp 1608254825
transform 1 0 6164 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_88
timestamp 1608254825
transform 1 0 9200 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__a41o_4  _2026_
timestamp 1608254825
transform 1 0 7636 0 -1 33184
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_6  FILLER_56_112
timestamp 1608254825
transform 1 0 11408 0 -1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_501
timestamp 1608254825
transform 1 0 9568 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2488_
timestamp 1608254825
transform 1 0 9660 0 -1 33184
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_56_137
timestamp 1608254825
transform 1 0 13708 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _2489_
timestamp 1608254825
transform 1 0 11960 0 -1 33184
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_56_149
timestamp 1608254825
transform 1 0 14812 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_502
timestamp 1608254825
transform 1 0 15180 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2620_
timestamp 1608254825
transform 1 0 15272 0 -1 33184
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  _1380_
timestamp 1608254825
transform 1 0 14444 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_181
timestamp 1608254825
transform 1 0 17756 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_173
timestamp 1608254825
transform 1 0 17020 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1366_
timestamp 1608254825
transform 1 0 17388 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_56_204
timestamp 1608254825
transform 1 0 19872 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _2622_
timestamp 1608254825
transform 1 0 18124 0 -1 33184
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_56_219
timestamp 1608254825
transform 1 0 21252 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_56_212
timestamp 1608254825
transform 1 0 20608 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_503
timestamp 1608254825
transform 1 0 20792 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2549_
timestamp 1608254825
transform 1 0 21620 0 -1 33184
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  _1379_
timestamp 1608254825
transform 1 0 20884 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_248
timestamp 1608254825
transform 1 0 23920 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_56_242
timestamp 1608254825
transform 1 0 23368 0 -1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  _2543_
timestamp 1608254825
transform 1 0 24012 0 -1 33184
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_56_274
timestamp 1608254825
transform 1 0 26312 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_56_268
timestamp 1608254825
transform 1 0 25760 0 -1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_56_295
timestamp 1608254825
transform 1 0 28244 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_504
timestamp 1608254825
transform 1 0 26404 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2384_
timestamp 1608254825
transform 1 0 26496 0 -1 33184
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  FILLER_56_316
timestamp 1608254825
transform 1 0 30176 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_56_308
timestamp 1608254825
transform 1 0 29440 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_4  _1762_
timestamp 1608254825
transform 1 0 28612 0 -1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_4  _1197_
timestamp 1608254825
transform 1 0 30452 0 -1 33184
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_6  FILLER_56_337
timestamp 1608254825
transform 1 0 32108 0 -1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_56_332
timestamp 1608254825
transform 1 0 31648 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_505
timestamp 1608254825
transform 1 0 32016 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_356
timestamp 1608254825
transform 1 0 33856 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__and2_4  _2095_
timestamp 1608254825
transform 1 0 34224 0 -1 33184
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_4  _1195_
timestamp 1608254825
transform 1 0 32660 0 -1 33184
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_1  FILLER_56_382
timestamp 1608254825
transform 1 0 36248 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_378
timestamp 1608254825
transform 1 0 35880 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_367
timestamp 1608254825
transform 1 0 34868 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__and2_4  _2093_
timestamp 1608254825
transform 1 0 35236 0 -1 33184
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_4  _1869_
timestamp 1608254825
transform 1 0 36340 0 -1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_56_406
timestamp 1608254825
transform 1 0 38456 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_398
timestamp 1608254825
transform 1 0 37720 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_396
timestamp 1608254825
transform 1 0 37536 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_392
timestamp 1608254825
transform 1 0 37168 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_506
timestamp 1608254825
transform 1 0 37628 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1608254825
transform -1 0 38824 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_57_12
timestamp 1608254825
transform 1 0 2208 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1608254825
transform 1 0 1104 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _2479_
timestamp 1608254825
transform 1 0 2576 0 1 33184
box -38 -48 1786 592
use sky130_fd_sc_hd__and3_4  _2057_
timestamp 1608254825
transform 1 0 1380 0 1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_57_43
timestamp 1608254825
transform 1 0 5060 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_35
timestamp 1608254825
transform 1 0 4324 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _2055_
timestamp 1608254825
transform 1 0 4692 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_57
timestamp 1608254825
transform 1 0 6348 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_47
timestamp 1608254825
transform 1 0 5428 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_507
timestamp 1608254825
transform 1 0 6716 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__nor3_4  _2046_
timestamp 1608254825
transform 1 0 6808 0 1 33184
box -38 -48 1234 592
use sky130_fd_sc_hd__and4_4  _2032_
timestamp 1608254825
transform 1 0 5520 0 1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_57_75
timestamp 1608254825
transform 1 0 8004 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__nand4_4  _1997_
timestamp 1608254825
transform 1 0 8372 0 1 33184
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_1  FILLER_57_104
timestamp 1608254825
transform 1 0 10672 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_96
timestamp 1608254825
transform 1 0 9936 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__nor3_4  _2019_
timestamp 1608254825
transform 1 0 10764 0 1 33184
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_57_118
timestamp 1608254825
transform 1 0 11960 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_508
timestamp 1608254825
transform 1 0 12328 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__a41oi_4  _2018_
timestamp 1608254825
transform 1 0 12420 0 1 33184
box -38 -48 2062 592
use sky130_fd_sc_hd__decap_4  FILLER_57_145
timestamp 1608254825
transform 1 0 14444 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_4  _1390_
timestamp 1608254825
transform 1 0 14812 0 1 33184
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_57_179
timestamp 1608254825
transform 1 0 17572 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_162
timestamp 1608254825
transform 1 0 16008 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_4  _1389_
timestamp 1608254825
transform 1 0 16376 0 1 33184
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_1  FILLER_57_205
timestamp 1608254825
transform 1 0 19964 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_201
timestamp 1608254825
transform 1 0 19596 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_509
timestamp 1608254825
transform 1 0 17940 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__nand4_4  _1385_
timestamp 1608254825
transform 1 0 18032 0 1 33184
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_2  FILLER_57_225
timestamp 1608254825
transform 1 0 21804 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_0
timestamp 1608254825
transform 1 0 21988 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _2619_
timestamp 1608254825
transform 1 0 20056 0 1 33184
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_57_236
timestamp 1608254825
transform 1 0 22816 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_510
timestamp 1608254825
transform 1 0 23552 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _1895_
timestamp 1608254825
transform 1 0 23644 0 1 33184
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _1893_
timestamp 1608254825
transform 1 0 22172 0 1 33184
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_57_267
timestamp 1608254825
transform 1 0 25668 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_263
timestamp 1608254825
transform 1 0 25300 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_252
timestamp 1608254825
transform 1 0 24288 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2383_
timestamp 1608254825
transform 1 0 25760 0 1 33184
box -38 -48 1786 592
use sky130_fd_sc_hd__and2_4  _1899_
timestamp 1608254825
transform 1 0 24656 0 1 33184
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_57_291
timestamp 1608254825
transform 1 0 27876 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_287
timestamp 1608254825
transform 1 0 27508 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_4  _1863_
timestamp 1608254825
transform 1 0 27968 0 1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_57_306
timestamp 1608254825
transform 1 0 29256 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_57_301
timestamp 1608254825
transform 1 0 28796 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_511
timestamp 1608254825
transform 1 0 29164 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2381_
timestamp 1608254825
transform 1 0 29532 0 1 33184
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_57_336
timestamp 1608254825
transform 1 0 32016 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_328
timestamp 1608254825
transform 1 0 31280 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _2456_
timestamp 1608254825
transform 1 0 32108 0 1 33184
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_57_364
timestamp 1608254825
transform 1 0 34592 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_57_356
timestamp 1608254825
transform 1 0 33856 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_57_380
timestamp 1608254825
transform 1 0 36064 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_367
timestamp 1608254825
transform 1 0 34868 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_512
timestamp 1608254825
transform 1 0 34776 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2567_
timestamp 1608254825
transform 1 0 36432 0 1 33184
box -38 -48 1786 592
use sky130_fd_sc_hd__nand2_4  _2346_
timestamp 1608254825
transform 1 0 35236 0 1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_57_403
timestamp 1608254825
transform 1 0 38180 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1608254825
transform -1 0 38824 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_58_22
timestamp 1608254825
transform 1 0 3128 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1608254825
transform 1 0 1104 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _2481_
timestamp 1608254825
transform 1 0 1380 0 -1 34272
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_58_32
timestamp 1608254825
transform 1 0 4048 0 -1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_30
timestamp 1608254825
transform 1 0 3864 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_513
timestamp 1608254825
transform 1 0 3956 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2485_
timestamp 1608254825
transform 1 0 4600 0 -1 34272
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_58_57
timestamp 1608254825
transform 1 0 6348 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__nand4_4  _2043_
timestamp 1608254825
transform 1 0 6716 0 -1 34272
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_6  FILLER_58_86
timestamp 1608254825
transform 1 0 9016 0 -1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_58_78
timestamp 1608254825
transform 1 0 8280 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _2016_
timestamp 1608254825
transform 1 0 8648 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_102
timestamp 1608254825
transform 1 0 10488 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_514
timestamp 1608254825
transform 1 0 9568 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__and4_4  _2017_
timestamp 1608254825
transform 1 0 9660 0 -1 34272
box -38 -48 866 592
use sky130_fd_sc_hd__nor4_4  _2013_
timestamp 1608254825
transform 1 0 10856 0 -1 34272
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_6  FILLER_58_123
timestamp 1608254825
transform 1 0 12420 0 -1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  _2491_
timestamp 1608254825
transform 1 0 12972 0 -1 34272
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  FILLER_58_154
timestamp 1608254825
transform 1 0 15272 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_58_152
timestamp 1608254825
transform 1 0 15088 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_148
timestamp 1608254825
transform 1 0 14720 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_515
timestamp 1608254825
transform 1 0 15180 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1387_
timestamp 1608254825
transform 1 0 15548 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_58_160
timestamp 1608254825
transform 1 0 15824 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2621_
timestamp 1608254825
transform 1 0 16192 0 -1 34272
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_58_183
timestamp 1608254825
transform 1 0 17940 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _2561_
timestamp 1608254825
transform 1 0 18676 0 -1 34272
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_58_225
timestamp 1608254825
transform 1 0 21804 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_58_215
timestamp 1608254825
transform 1 0 20884 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_58_210
timestamp 1608254825
transform 1 0 20424 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_516
timestamp 1608254825
transform 1 0 20792 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _1894_
timestamp 1608254825
transform 1 0 21160 0 -1 34272
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_58_248
timestamp 1608254825
transform 1 0 23920 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2547_
timestamp 1608254825
transform 1 0 22172 0 -1 34272
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_58_271
timestamp 1608254825
transform 1 0 26036 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2544_
timestamp 1608254825
transform 1 0 24288 0 -1 34272
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  FILLER_58_291
timestamp 1608254825
transform 1 0 27876 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_58_283
timestamp 1608254825
transform 1 0 27140 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_517
timestamp 1608254825
transform 1 0 26404 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2379_
timestamp 1608254825
transform 1 0 28152 0 -1 34272
box -38 -48 1786 592
use sky130_fd_sc_hd__and2_4  _1900_
timestamp 1608254825
transform 1 0 26496 0 -1 34272
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_58_313
timestamp 1608254825
transform 1 0 29900 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1191_
timestamp 1608254825
transform 1 0 30268 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_341
timestamp 1608254825
transform 1 0 32476 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_332
timestamp 1608254825
transform 1 0 31648 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_321
timestamp 1608254825
transform 1 0 30636 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_518
timestamp 1608254825
transform 1 0 32016 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _2097_
timestamp 1608254825
transform 1 0 31004 0 -1 34272
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _2096_
timestamp 1608254825
transform 1 0 32108 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_352
timestamp 1608254825
transform 1 0 33488 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2457_
timestamp 1608254825
transform 1 0 33856 0 -1 34272
box -38 -48 1786 592
use sky130_fd_sc_hd__and2_4  _2107_
timestamp 1608254825
transform 1 0 32844 0 -1 34272
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_58_375
timestamp 1608254825
transform 1 0 35604 0 -1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_4  _2347_
timestamp 1608254825
transform 1 0 36156 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_406
timestamp 1608254825
transform 1 0 38456 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_398
timestamp 1608254825
transform 1 0 37720 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_58_393
timestamp 1608254825
transform 1 0 37260 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_519
timestamp 1608254825
transform 1 0 37628 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1608254825
transform -1 0 38824 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_60_7
timestamp 1608254825
transform 1 0 1748 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_12
timestamp 1608254825
transform 1 0 2208 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1608254825
transform 1 0 1104 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1608254825
transform 1 0 1104 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_4  _2052_
timestamp 1608254825
transform 1 0 2116 0 -1 35360
box -38 -48 1234 592
use sky130_fd_sc_hd__and3_4  _2044_
timestamp 1608254825
transform 1 0 1380 0 1 34272
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _2040_
timestamp 1608254825
transform 1 0 1380 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__nand4_4  _1993_
timestamp 1608254825
transform 1 0 2576 0 1 34272
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_6  FILLER_60_45
timestamp 1608254825
transform 1 0 5244 0 -1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_30
timestamp 1608254825
transform 1 0 3864 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_60_24
timestamp 1608254825
transform 1 0 3312 0 -1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_59_33
timestamp 1608254825
transform 1 0 4140 0 1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_526
timestamp 1608254825
transform 1 0 3956 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_4  _2048_
timestamp 1608254825
transform 1 0 4048 0 -1 35360
box -38 -48 1234 592
use sky130_fd_sc_hd__a41o_4  _2042_
timestamp 1608254825
transform 1 0 4692 0 1 34272
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_6  FILLER_60_61
timestamp 1608254825
transform 1 0 6716 0 -1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_51
timestamp 1608254825
transform 1 0 5796 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_59_62
timestamp 1608254825
transform 1 0 6808 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_59_60
timestamp 1608254825
transform 1 0 6624 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_56
timestamp 1608254825
transform 1 0 6256 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_520
timestamp 1608254825
transform 1 0 6716 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2484_
timestamp 1608254825
transform 1 0 7268 0 -1 35360
box -38 -48 1786 592
use sky130_fd_sc_hd__a21oi_4  _2045_
timestamp 1608254825
transform 1 0 7084 0 1 34272
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_4  _2029_
timestamp 1608254825
transform 1 0 5888 0 -1 35360
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_60_86
timestamp 1608254825
transform 1 0 9016 0 -1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_59_86
timestamp 1608254825
transform 1 0 9016 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_59_78
timestamp 1608254825
transform 1 0 8280 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_4  _2021_
timestamp 1608254825
transform 1 0 9200 0 1 34272
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_1  FILLER_60_103
timestamp 1608254825
transform 1 0 10580 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_60_97
timestamp 1608254825
transform 1 0 10028 0 -1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_59_101
timestamp 1608254825
transform 1 0 10396 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_527
timestamp 1608254825
transform 1 0 9568 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__nand3_4  _2022_
timestamp 1608254825
transform 1 0 10672 0 -1 35360
box -38 -48 1326 592
use sky130_fd_sc_hd__buf_2  _2012_
timestamp 1608254825
transform 1 0 9660 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_4  _2004_
timestamp 1608254825
transform 1 0 10764 0 1 34272
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_2  FILLER_60_126
timestamp 1608254825
transform 1 0 12696 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_60_118
timestamp 1608254825
transform 1 0 11960 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_59_127
timestamp 1608254825
transform 1 0 12788 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_118
timestamp 1608254825
transform 1 0 11960 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_521
timestamp 1608254825
transform 1 0 12328 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__a41o_4  _2009_
timestamp 1608254825
transform 1 0 13156 0 1 34272
box -38 -48 1602 592
use sky130_fd_sc_hd__buf_2  _2002_
timestamp 1608254825
transform 1 0 12420 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__nand4_4  _1999_
timestamp 1608254825
transform 1 0 12880 0 -1 35360
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_8  FILLER_60_145
timestamp 1608254825
transform 1 0 14444 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_59_159
timestamp 1608254825
transform 1 0 15732 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_155
timestamp 1608254825
transform 1 0 15364 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_148
timestamp 1608254825
transform 1 0 14720 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_528
timestamp 1608254825
transform 1 0 15180 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _2003_
timestamp 1608254825
transform 1 0 15088 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_4  _1393_
timestamp 1608254825
transform 1 0 15272 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_174
timestamp 1608254825
transform 1 0 17112 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_60_166
timestamp 1608254825
transform 1 0 16376 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_59_179
timestamp 1608254825
transform 1 0 17572 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2562_
timestamp 1608254825
transform 1 0 15824 0 1 34272
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _2554_
timestamp 1608254825
transform 1 0 17204 0 -1 35360
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_60_205
timestamp 1608254825
transform 1 0 19964 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_194
timestamp 1608254825
transform 1 0 18952 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_197
timestamp 1608254825
transform 1 0 19228 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_193
timestamp 1608254825
transform 1 0 18860 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_522
timestamp 1608254825
transform 1 0 17940 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2553_
timestamp 1608254825
transform 1 0 19320 0 1 34272
box -38 -48 1786 592
use sky130_fd_sc_hd__and2_4  _1887_
timestamp 1608254825
transform 1 0 19320 0 -1 35360
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_4  _1386_
timestamp 1608254825
transform 1 0 18032 0 1 34272
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_60_222
timestamp 1608254825
transform 1 0 21528 0 -1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_60_212
timestamp 1608254825
transform 1 0 20608 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_217
timestamp 1608254825
transform 1 0 21068 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_12_0_m1_clk_local
timestamp 1608254825
transform 1 0 20332 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_m1_clk_local
timestamp 1608254825
transform 1 0 22080 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_529
timestamp 1608254825
transform 1 0 20792 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2548_
timestamp 1608254825
transform 1 0 21436 0 1 34272
box -38 -48 1786 592
use sky130_fd_sc_hd__and2_4  _1888_
timestamp 1608254825
transform 1 0 20884 0 -1 35360
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_60_250
timestamp 1608254825
transform 1 0 24104 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_249
timestamp 1608254825
transform 1 0 24012 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_245
timestamp 1608254825
transform 1 0 23644 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_240
timestamp 1608254825
transform 1 0 23184 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_523
timestamp 1608254825
transform 1 0 23552 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2550_
timestamp 1608254825
transform 1 0 22356 0 -1 35360
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _2546_
timestamp 1608254825
transform 1 0 24104 0 1 34272
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_60_274
timestamp 1608254825
transform 1 0 26312 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_60_268
timestamp 1608254825
transform 1 0 25760 0 -1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_60_261
timestamp 1608254825
transform 1 0 25116 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_59_269
timestamp 1608254825
transform 1 0 25852 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_m1_clk_local
timestamp 1608254825
transform 1 0 25484 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__and2_4  _1896_
timestamp 1608254825
transform 1 0 24472 0 -1 35360
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_60_295
timestamp 1608254825
transform 1 0 28244 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_281
timestamp 1608254825
transform 1 0 26956 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_530
timestamp 1608254825
transform 1 0 26404 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2378_
timestamp 1608254825
transform 1 0 27048 0 1 34272
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _2377_
timestamp 1608254825
transform 1 0 26496 0 -1 35360
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_60_318
timestamp 1608254825
transform 1 0 30360 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_60_302
timestamp 1608254825
transform 1 0 28888 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_59_301
timestamp 1608254825
transform 1 0 28796 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_m1_clk_local
timestamp 1608254825
transform 1 0 28612 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_524
timestamp 1608254825
transform 1 0 29164 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2380_
timestamp 1608254825
transform 1 0 29256 0 1 34272
box -38 -48 1786 592
use sky130_fd_sc_hd__a21oi_4  _2350_
timestamp 1608254825
transform 1 0 29164 0 -1 35360
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_1  FILLER_60_337
timestamp 1608254825
transform 1 0 32108 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_332
timestamp 1608254825
transform 1 0 31648 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_325
timestamp 1608254825
transform 1 0 31004 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_14_0_m1_clk_local
timestamp 1608254825
transform 1 0 30728 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_531
timestamp 1608254825
transform 1 0 32016 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2498_
timestamp 1608254825
transform 1 0 32200 0 -1 35360
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _2464_
timestamp 1608254825
transform 1 0 31372 0 1 34272
box -38 -48 1786 592
use sky130_fd_sc_hd__and2_4  _2108_
timestamp 1608254825
transform 1 0 31004 0 -1 35360
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_60_357
timestamp 1608254825
transform 1 0 33948 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_362
timestamp 1608254825
transform 1 0 34408 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_352
timestamp 1608254825
transform 1 0 33488 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_348
timestamp 1608254825
transform 1 0 33120 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__or3_4  _1981_
timestamp 1608254825
transform 1 0 33580 0 1 34272
box -38 -48 866 592
use sky130_fd_sc_hd__nor3_4  _1867_
timestamp 1608254825
transform 1 0 34316 0 -1 35360
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_8  FILLER_60_387
timestamp 1608254825
transform 1 0 36708 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_60_374
timestamp 1608254825
transform 1 0 35512 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_373
timestamp 1608254825
transform 1 0 35420 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_59_367
timestamp 1608254825
transform 1 0 34868 0 1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_525
timestamp 1608254825
transform 1 0 34776 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__xnor2_4  _1868_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 35512 0 1 34272
box -38 -48 2062 592
use sky130_fd_sc_hd__nand2_4  _1866_
timestamp 1608254825
transform 1 0 35880 0 -1 35360
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_60_406
timestamp 1608254825
transform 1 0 38456 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_60_398
timestamp 1608254825
transform 1 0 37720 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_395
timestamp 1608254825
transform 1 0 37444 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_59_404
timestamp 1608254825
transform 1 0 38272 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_59_396
timestamp 1608254825
transform 1 0 37536 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_532
timestamp 1608254825
transform 1 0 37628 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1608254825
transform -1 0 38824 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1608254825
transform -1 0 38824 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_61_3
timestamp 1608254825
transform 1 0 1380 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1608254825
transform 1 0 1104 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _2482_
timestamp 1608254825
transform 1 0 2116 0 1 35360
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_61_38
timestamp 1608254825
transform 1 0 4600 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_61_30
timestamp 1608254825
transform 1 0 3864 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__nor3_4  _2015_
timestamp 1608254825
transform 1 0 4784 0 1 35360
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_8  FILLER_61_53
timestamp 1608254825
transform 1 0 5980 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_533
timestamp 1608254825
transform 1 0 6716 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__nor4_4  _1994_
timestamp 1608254825
transform 1 0 6808 0 1 35360
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_1  FILLER_61_85
timestamp 1608254825
transform 1 0 8924 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_61_79
timestamp 1608254825
transform 1 0 8372 0 1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_4  _2001_
timestamp 1608254825
transform 1 0 9016 0 1 35360
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_61_95
timestamp 1608254825
transform 1 0 9844 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__nand4_4  _2005_
timestamp 1608254825
transform 1 0 10212 0 1 35360
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_61_126
timestamp 1608254825
transform 1 0 12696 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_61_116
timestamp 1608254825
transform 1 0 11776 0 1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_534
timestamp 1608254825
transform 1 0 12328 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _1998_
timestamp 1608254825
transform 1 0 13064 0 1 35360
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1984_
timestamp 1608254825
transform 1 0 12420 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_61_139
timestamp 1608254825
transform 1 0 13892 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2492_
timestamp 1608254825
transform 1 0 14260 0 1 35360
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_61_181
timestamp 1608254825
transform 1 0 17756 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_61_173
timestamp 1608254825
transform 1 0 17020 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_61_162
timestamp 1608254825
transform 1 0 16008 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__and2_4  _1877_
timestamp 1608254825
transform 1 0 16376 0 1 35360
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_61_193
timestamp 1608254825
transform 1 0 18860 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_61_184
timestamp 1608254825
transform 1 0 18032 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_535
timestamp 1608254825
transform 1 0 17940 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2366_
timestamp 1608254825
transform 1 0 19228 0 1 35360
box -38 -48 1786 592
use sky130_fd_sc_hd__and2_4  _1878_
timestamp 1608254825
transform 1 0 18216 0 1 35360
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_61_227
timestamp 1608254825
transform 1 0 21988 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_223
timestamp 1608254825
transform 1 0 21620 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_216
timestamp 1608254825
transform 1 0 20976 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_13_0_m1_clk_local
timestamp 1608254825
transform 1 0 21344 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__and2_4  _1891_
timestamp 1608254825
transform 1 0 22080 0 1 35360
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  FILLER_61_245
timestamp 1608254825
transform 1 0 23644 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_61_243
timestamp 1608254825
transform 1 0 23460 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_235
timestamp 1608254825
transform 1 0 22724 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_536
timestamp 1608254825
transform 1 0 23552 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2371_
timestamp 1608254825
transform 1 0 23920 0 1 35360
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_61_267
timestamp 1608254825
transform 1 0 25668 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2534_
timestamp 1608254825
transform 1 0 26036 0 1 35360
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_61_290
timestamp 1608254825
transform 1 0 27784 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_15_0_m1_clk_local
timestamp 1608254825
transform 1 0 28888 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_537
timestamp 1608254825
transform 1 0 29164 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2376_
timestamp 1608254825
transform 1 0 29256 0 1 35360
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_61_325
timestamp 1608254825
transform 1 0 31004 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_3
timestamp 1608254825
transform 1 0 31188 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _2501_
timestamp 1608254825
transform 1 0 31372 0 1 35360
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_61_362
timestamp 1608254825
transform 1 0 34408 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_352
timestamp 1608254825
transform 1 0 33488 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_348
timestamp 1608254825
transform 1 0 33120 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_4  _1973_
timestamp 1608254825
transform 1 0 33580 0 1 35360
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_61_380
timestamp 1608254825
transform 1 0 36064 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_538
timestamp 1608254825
transform 1 0 34776 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2495_
timestamp 1608254825
transform 1 0 36432 0 1 35360
box -38 -48 1786 592
use sky130_fd_sc_hd__a21oi_4  _1974_
timestamp 1608254825
transform 1 0 34868 0 1 35360
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_61_403
timestamp 1608254825
transform 1 0 38180 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1608254825
transform -1 0 38824 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_62_11
timestamp 1608254825
transform 1 0 2116 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_3
timestamp 1608254825
transform 1 0 1380 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1608254825
transform 1 0 1104 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_4  _2051_
timestamp 1608254825
transform 1 0 2208 0 -1 36448
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_6  FILLER_62_25
timestamp 1608254825
transform 1 0 3404 0 -1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_539
timestamp 1608254825
transform 1 0 3956 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__nand3_4  _2049_
timestamp 1608254825
transform 1 0 4048 0 -1 36448
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_2  FILLER_62_54
timestamp 1608254825
transform 1 0 6072 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_62_46
timestamp 1608254825
transform 1 0 5336 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _2511_
timestamp 1608254825
transform 1 0 6256 0 -1 36448
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_62_90
timestamp 1608254825
transform 1 0 9384 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_62_82
timestamp 1608254825
transform 1 0 8648 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_62_75
timestamp 1608254825
transform 1 0 8004 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1987_
timestamp 1608254825
transform 1 0 8372 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_62_114
timestamp 1608254825
transform 1 0 11592 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_107
timestamp 1608254825
transform 1 0 10948 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_540
timestamp 1608254825
transform 1 0 9568 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__nand3_4  _2006_
timestamp 1608254825
transform 1 0 9660 0 -1 36448
box -38 -48 1326 592
use sky130_fd_sc_hd__inv_2  _2000_
timestamp 1608254825
transform 1 0 11316 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_62_137
timestamp 1608254825
transform 1 0 13708 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2490_
timestamp 1608254825
transform 1 0 11960 0 -1 36448
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_62_152
timestamp 1608254825
transform 1 0 15088 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_144
timestamp 1608254825
transform 1 0 14352 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_541
timestamp 1608254825
transform 1 0 15180 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__and3_4  _2010_
timestamp 1608254825
transform 1 0 15272 0 -1 36448
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _2008_
timestamp 1608254825
transform 1 0 14076 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_62_163
timestamp 1608254825
transform 1 0 16100 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _2364_
timestamp 1608254825
transform 1 0 16836 0 -1 36448
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_62_196
timestamp 1608254825
transform 1 0 19136 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_62_190
timestamp 1608254825
transform 1 0 18584 0 -1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_4  _1865_
timestamp 1608254825
transform 1 0 19228 0 -1 36448
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_62_210
timestamp 1608254825
transform 1 0 20424 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_542
timestamp 1608254825
transform 1 0 20792 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2367_
timestamp 1608254825
transform 1 0 20884 0 -1 36448
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_62_234
timestamp 1608254825
transform 1 0 22632 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2369_
timestamp 1608254825
transform 1 0 23000 0 -1 36448
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_62_269
timestamp 1608254825
transform 1 0 25852 0 -1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_62_257
timestamp 1608254825
transform 1 0 24748 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_295
timestamp 1608254825
transform 1 0 28244 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_543
timestamp 1608254825
transform 1 0 26404 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2373_
timestamp 1608254825
transform 1 0 26496 0 -1 36448
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_62_318
timestamp 1608254825
transform 1 0 30360 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _2375_
timestamp 1608254825
transform 1 0 28612 0 -1 36448
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_62_341
timestamp 1608254825
transform 1 0 32476 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_337
timestamp 1608254825
transform 1 0 32108 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_335
timestamp 1608254825
transform 1 0 31924 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_62_329
timestamp 1608254825
transform 1 0 31372 0 -1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_544
timestamp 1608254825
transform 1 0 32016 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _2348_
timestamp 1608254825
transform 1 0 31096 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_4  _1975_
timestamp 1608254825
transform 1 0 32568 0 -1 36448
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_3  FILLER_62_363
timestamp 1608254825
transform 1 0 34500 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_62_355
timestamp 1608254825
transform 1 0 33764 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_62_380
timestamp 1608254825
transform 1 0 36064 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__and3_4  _1978_
timestamp 1608254825
transform 1 0 36432 0 -1 36448
box -38 -48 866 592
use sky130_fd_sc_hd__nand3_4  _1972_
timestamp 1608254825
transform 1 0 34776 0 -1 36448
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_6  FILLER_62_401
timestamp 1608254825
transform 1 0 37996 0 -1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_62_393
timestamp 1608254825
transform 1 0 37260 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_545
timestamp 1608254825
transform 1 0 37628 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1608254825
transform -1 0 38824 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1982_
timestamp 1608254825
transform 1 0 37720 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_63_19
timestamp 1608254825
transform 1 0 2852 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_11
timestamp 1608254825
transform 1 0 2116 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_3
timestamp 1608254825
transform 1 0 1380 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_2
timestamp 1608254825
transform 1 0 2300 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1608254825
transform 1 0 1104 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _2361_
timestamp 1608254825
transform 1 0 2484 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _2359_
timestamp 1608254825
transform 1 0 1748 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_27
timestamp 1608254825
transform 1 0 3588 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_23
timestamp 1608254825
transform 1 0 3220 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2483_
timestamp 1608254825
transform 1 0 3956 0 1 36448
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_2  _2050_
timestamp 1608254825
transform 1 0 3312 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_63_66
timestamp 1608254825
transform 1 0 7176 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_57
timestamp 1608254825
transform 1 0 6348 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_50
timestamp 1608254825
transform 1 0 5704 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_546
timestamp 1608254825
transform 1 0 6716 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _2030_
timestamp 1608254825
transform 1 0 6808 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1985_
timestamp 1608254825
transform 1 0 6072 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_63_78
timestamp 1608254825
transform 1 0 8280 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2493_
timestamp 1608254825
transform 1 0 8648 0 1 36448
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_63_111
timestamp 1608254825
transform 1 0 11316 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_107
timestamp 1608254825
transform 1 0 10948 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_63_101
timestamp 1608254825
transform 1 0 10396 0 1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _2020_
timestamp 1608254825
transform 1 0 11040 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_63_118
timestamp 1608254825
transform 1 0 11960 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_547
timestamp 1608254825
transform 1 0 12328 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2470_
timestamp 1608254825
transform 1 0 12420 0 1 36448
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_2  _2011_
timestamp 1608254825
transform 1 0 11684 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_63_153
timestamp 1608254825
transform 1 0 15180 0 1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_63_142
timestamp 1608254825
transform 1 0 14168 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _2363_
timestamp 1608254825
transform 1 0 15732 0 1 36448
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_2  _2341_
timestamp 1608254825
transform 1 0 14904 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_63_182
timestamp 1608254825
transform 1 0 17848 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_178
timestamp 1608254825
transform 1 0 17480 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_63_203
timestamp 1608254825
transform 1 0 19780 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_548
timestamp 1608254825
transform 1 0 17940 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2365_
timestamp 1608254825
transform 1 0 18032 0 1 36448
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_63_218
timestamp 1608254825
transform 1 0 21160 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_214
timestamp 1608254825
transform 1 0 20792 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2368_
timestamp 1608254825
transform 1 0 21252 0 1 36448
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_2  _1864_
timestamp 1608254825
transform 1 0 20516 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_63_238
timestamp 1608254825
transform 1 0 23000 0 1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_549
timestamp 1608254825
transform 1 0 23552 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2370_
timestamp 1608254825
transform 1 0 23644 0 1 36448
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_63_264
timestamp 1608254825
transform 1 0 25392 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_276
timestamp 1608254825
transform 1 0 26496 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2374_
timestamp 1608254825
transform 1 0 26864 0 1 36448
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_63_319
timestamp 1608254825
transform 1 0 30452 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_315
timestamp 1608254825
transform 1 0 30084 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_63_299
timestamp 1608254825
transform 1 0 28612 0 1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_550
timestamp 1608254825
transform 1 0 29164 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _2349_
timestamp 1608254825
transform 1 0 29256 0 1 36448
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_63_339
timestamp 1608254825
transform 1 0 32292 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2508_
timestamp 1608254825
transform 1 0 30544 0 1 36448
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_63_362
timestamp 1608254825
transform 1 0 34408 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2497_
timestamp 1608254825
transform 1 0 32660 0 1 36448
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_63_375
timestamp 1608254825
transform 1 0 35604 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_367
timestamp 1608254825
transform 1 0 34868 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_551
timestamp 1608254825
transform 1 0 34776 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2496_
timestamp 1608254825
transform 1 0 35972 0 1 36448
box -38 -48 1786 592
use sky130_fd_sc_hd__or2_4  _1979_
timestamp 1608254825
transform 1 0 34960 0 1 36448
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_63_406
timestamp 1608254825
transform 1 0 38456 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_398
timestamp 1608254825
transform 1 0 37720 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1608254825
transform -1 0 38824 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_15
timestamp 1608254825
transform 1 0 2484 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_3
timestamp 1608254825
transform 1 0 1380 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1608254825
transform 1 0 1104 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_64_44
timestamp 1608254825
transform 1 0 5152 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_37
timestamp 1608254825
transform 1 0 4508 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_32
timestamp 1608254825
transform 1 0 4048 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_27
timestamp 1608254825
transform 1 0 3588 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_552
timestamp 1608254825
transform 1 0 3956 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _2047_
timestamp 1608254825
transform 1 0 4232 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1986_
timestamp 1608254825
transform 1 0 4876 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_64_63
timestamp 1608254825
transform 1 0 6900 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_64_60
timestamp 1608254825
transform 1 0 6624 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_52
timestamp 1608254825
transform 1 0 5888 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_553
timestamp 1608254825
transform 1 0 6808 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _2014_
timestamp 1608254825
transform 1 0 5520 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_89
timestamp 1608254825
transform 1 0 9292 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_69
timestamp 1608254825
transform 1 0 7452 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2499_
timestamp 1608254825
transform 1 0 7544 0 -1 37536
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_64_109
timestamp 1608254825
transform 1 0 11132 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_64_97
timestamp 1608254825
transform 1 0 10028 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_554
timestamp 1608254825
transform 1 0 9660 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _2007_
timestamp 1608254825
transform 1 0 9752 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_137
timestamp 1608254825
transform 1 0 13708 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_125
timestamp 1608254825
transform 1 0 12604 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_118
timestamp 1608254825
transform 1 0 11960 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_555
timestamp 1608254825
transform 1 0 12512 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _2023_
timestamp 1608254825
transform 1 0 11684 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_64_149
timestamp 1608254825
transform 1 0 14812 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_556
timestamp 1608254825
transform 1 0 15364 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2382_
timestamp 1608254825
transform 1 0 15456 0 -1 37536
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_64_175
timestamp 1608254825
transform 1 0 17204 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_64_199
timestamp 1608254825
transform 1 0 19412 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_187
timestamp 1608254825
transform 1 0 18308 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_183
timestamp 1608254825
transform 1 0 17940 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_557
timestamp 1608254825
transform 1 0 18216 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_218
timestamp 1608254825
transform 1 0 21160 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_211
timestamp 1608254825
transform 1 0 20516 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_558
timestamp 1608254825
transform 1 0 21068 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_64_249
timestamp 1608254825
transform 1 0 24012 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_64_242
timestamp 1608254825
transform 1 0 23368 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_64_230
timestamp 1608254825
transform 1 0 22264 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_559
timestamp 1608254825
transform 1 0 23920 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_64_255
timestamp 1608254825
transform 1 0 24564 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2372_
timestamp 1608254825
transform 1 0 24656 0 -1 37536
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_64_292
timestamp 1608254825
transform 1 0 27968 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_280
timestamp 1608254825
transform 1 0 26864 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_275
timestamp 1608254825
transform 1 0 26404 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_560
timestamp 1608254825
transform 1 0 26772 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_64_311
timestamp 1608254825
transform 1 0 29716 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_64_304
timestamp 1608254825
transform 1 0 29072 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_5
timestamp 1608254825
transform 1 0 29808 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_561
timestamp 1608254825
transform 1 0 29624 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2532_
timestamp 1608254825
transform 1 0 29992 0 -1 37536
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_64_342
timestamp 1608254825
transform 1 0 32568 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_333
timestamp 1608254825
transform 1 0 31740 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_562
timestamp 1608254825
transform 1 0 32476 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_363
timestamp 1608254825
transform 1 0 34500 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_4  _1976_
timestamp 1608254825
transform 1 0 33672 0 -1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_64_385
timestamp 1608254825
transform 1 0 36524 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_371
timestamp 1608254825
transform 1 0 35236 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_563
timestamp 1608254825
transform 1 0 35328 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__a21o_4  _1977_
timestamp 1608254825
transform 1 0 35420 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_404
timestamp 1608254825
transform 1 0 38272 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_64_402
timestamp 1608254825
transform 1 0 38088 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_398
timestamp 1608254825
transform 1 0 37720 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_564
timestamp 1608254825
transform 1 0 38180 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1608254825
transform -1 0 38824 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__and3_4  _1980_
timestamp 1608254825
transform 1 0 36892 0 -1 37536
box -38 -48 866 592
<< labels >>
rlabel metal2 s 3330 39200 3386 40000 6 CLK_LED
port 0 nsew signal tristate
rlabel metal2 s 21914 39200 21970 40000 6 DATA_AVAILABLE[0]
port 1 nsew signal input
rlabel metal2 s 17682 39200 17738 40000 6 DATA_AVAILABLE[1]
port 2 nsew signal input
rlabel metal3 s 0 12792 800 12912 6 DATA_AVAILABLE[2]
port 3 nsew signal input
rlabel metal2 s 34242 39200 34298 40000 6 DATA_AVAILABLE[3]
port 4 nsew signal input
rlabel metal2 s 18970 0 19026 800 6 DATA_FROM_HASH[0]
port 5 nsew signal input
rlabel metal2 s 23018 0 23074 800 6 DATA_FROM_HASH[1]
port 6 nsew signal input
rlabel metal2 s 30010 39200 30066 40000 6 DATA_FROM_HASH[2]
port 7 nsew signal input
rlabel metal2 s 5354 39200 5410 40000 6 DATA_FROM_HASH[3]
port 8 nsew signal input
rlabel metal3 s 0 19048 800 19168 6 DATA_FROM_HASH[4]
port 9 nsew signal input
rlabel metal3 s 39200 10072 40000 10192 6 DATA_FROM_HASH[5]
port 10 nsew signal input
rlabel metal2 s 15658 39200 15714 40000 6 DATA_FROM_HASH[6]
port 11 nsew signal input
rlabel metal2 s 25226 0 25282 800 6 DATA_FROM_HASH[7]
port 12 nsew signal input
rlabel metal3 s 0 28024 800 28144 6 DATA_TO_HASH[0]
port 13 nsew signal tristate
rlabel metal2 s 36266 39200 36322 40000 6 DATA_TO_HASH[1]
port 14 nsew signal tristate
rlabel metal2 s 4618 0 4674 800 6 DATA_TO_HASH[2]
port 15 nsew signal tristate
rlabel metal2 s 35346 0 35402 800 6 DATA_TO_HASH[3]
port 16 nsew signal tristate
rlabel metal2 s 7378 39200 7434 40000 6 DATA_TO_HASH[4]
port 17 nsew signal tristate
rlabel metal3 s 39200 1096 40000 1216 6 DATA_TO_HASH[5]
port 18 nsew signal tristate
rlabel metal3 s 39200 19320 40000 19440 6 DATA_TO_HASH[6]
port 19 nsew signal tristate
rlabel metal2 s 33322 0 33378 800 6 DATA_TO_HASH[7]
port 20 nsew signal tristate
rlabel metal2 s 23938 39200 23994 40000 6 EXT_RESET_N_fromHost
port 21 nsew signal input
rlabel metal3 s 0 31016 800 31136 6 EXT_RESET_N_toClient
port 22 nsew signal tristate
rlabel metal2 s 31298 0 31354 800 6 HASH_ADDR[0]
port 23 nsew signal tristate
rlabel metal2 s 32034 39200 32090 40000 6 HASH_ADDR[1]
port 24 nsew signal tristate
rlabel metal2 s 10690 0 10746 800 6 HASH_ADDR[2]
port 25 nsew signal tristate
rlabel metal2 s 27986 39200 28042 40000 6 HASH_ADDR[3]
port 26 nsew signal tristate
rlabel metal3 s 0 6808 800 6928 6 HASH_ADDR[4]
port 27 nsew signal tristate
rlabel metal3 s 0 9800 800 9920 6 HASH_ADDR[5]
port 28 nsew signal tristate
rlabel metal2 s 13634 39200 13690 40000 6 HASH_EN
port 29 nsew signal tristate
rlabel metal3 s 0 15784 800 15904 6 HASH_LED
port 30 nsew signal tristate
rlabel metal3 s 39200 13336 40000 13456 6 ID_fromClient
port 31 nsew signal input
rlabel metal3 s 0 34008 800 34128 6 ID_toHost
port 32 nsew signal tristate
rlabel metal3 s 39200 22312 40000 22432 6 IRQ_OUT_fromClient
port 33 nsew signal input
rlabel metal3 s 0 3816 800 3936 6 IRQ_OUT_toHost
port 34 nsew signal tristate
rlabel metal2 s 8666 0 8722 800 6 M1_CLK_IN
port 35 nsew signal input
rlabel metal2 s 6642 0 6698 800 6 M1_CLK_SELECT
port 36 nsew signal input
rlabel metal2 s 27250 0 27306 800 6 MACRO_RD_SELECT[0]
port 37 nsew signal tristate
rlabel metal2 s 20994 0 21050 800 6 MACRO_RD_SELECT[1]
port 38 nsew signal tristate
rlabel metal2 s 16946 0 17002 800 6 MACRO_RD_SELECT[2]
port 39 nsew signal tristate
rlabel metal2 s 12898 0 12954 800 6 MACRO_RD_SELECT[3]
port 40 nsew signal tristate
rlabel metal2 s 9402 39200 9458 40000 6 MACRO_WR_SELECT[0]
port 41 nsew signal tristate
rlabel metal2 s 2594 0 2650 800 6 MACRO_WR_SELECT[1]
port 42 nsew signal tristate
rlabel metal2 s 38290 39200 38346 40000 6 MACRO_WR_SELECT[2]
port 43 nsew signal tristate
rlabel metal3 s 39200 7080 40000 7200 6 MACRO_WR_SELECT[3]
port 44 nsew signal tristate
rlabel metal2 s 1306 39200 1362 40000 6 MISO_fromClient
port 45 nsew signal input
rlabel metal2 s 25962 39200 26018 40000 6 MISO_toHost
port 46 nsew signal tristate
rlabel metal3 s 39200 37544 40000 37664 6 MOSI_fromHost
port 47 nsew signal input
rlabel metal3 s 39200 16328 40000 16448 6 MOSI_toClient
port 48 nsew signal tristate
rlabel metal3 s 39200 4088 40000 4208 6 PLL_INPUT
port 49 nsew signal input
rlabel metal3 s 0 22040 800 22160 6 S1_CLK_IN
port 50 nsew signal input
rlabel metal3 s 39200 34552 40000 34672 6 S1_CLK_SELECT
port 51 nsew signal input
rlabel metal3 s 39200 31560 40000 31680 6 SCLK_fromHost
port 52 nsew signal input
rlabel metal3 s 0 37272 800 37392 6 SCLK_toClient
port 53 nsew signal tristate
rlabel metal2 s 19706 39200 19762 40000 6 SCSN_fromHost
port 54 nsew signal input
rlabel metal3 s 39200 28296 40000 28416 6 SCSN_toClient
port 55 nsew signal tristate
rlabel metal2 s 570 0 626 800 6 THREAD_COUNT[0]
port 56 nsew signal input
rlabel metal3 s 39200 25304 40000 25424 6 THREAD_COUNT[1]
port 57 nsew signal input
rlabel metal2 s 14922 0 14978 800 6 THREAD_COUNT[2]
port 58 nsew signal input
rlabel metal2 s 11610 39200 11666 40000 6 THREAD_COUNT[3]
port 59 nsew signal input
rlabel metal3 s 0 25032 800 25152 6 m1_clk_local
port 60 nsew signal tristate
rlabel metal2 s 29274 0 29330 800 6 one
port 61 nsew signal tristate
rlabel metal2 s 37554 0 37610 800 6 zero
port 62 nsew signal tristate
rlabel metal4 s 34928 2128 35248 37584 6 VPWR
port 63 nsew power bidirectional
rlabel metal4 s 4208 2128 4528 37584 6 VPWR
port 64 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 37584 6 VGND
port 65 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 40000 40000
<< end >>

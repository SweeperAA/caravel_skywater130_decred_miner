* NGSPICE file created from decred_controller.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_4 abstract view
.subckt sky130_fd_sc_hd__a41o_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_4 abstract view
.subckt sky130_fd_sc_hd__and4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_4 abstract view
.subckt sky130_fd_sc_hd__nand4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41oi_4 abstract view
.subckt sky130_fd_sc_hd__a41oi_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41ai_4 abstract view
.subckt sky130_fd_sc_hd__o41ai_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_4 abstract view
.subckt sky130_fd_sc_hd__a211o_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_4 abstract view
.subckt sky130_fd_sc_hd__o32a_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_4 abstract view
.subckt sky130_fd_sc_hd__o41a_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_4 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_4 abstract view
.subckt sky130_fd_sc_hd__a21boi_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_4 abstract view
.subckt sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_4 abstract view
.subckt sky130_fd_sc_hd__a2111o_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_4 abstract view
.subckt sky130_fd_sc_hd__nor4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2oi_4 abstract view
.subckt sky130_fd_sc_hd__a2bb2oi_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_4 abstract view
.subckt sky130_fd_sc_hd__o32ai_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_4 abstract view
.subckt sky130_fd_sc_hd__a2111oi_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

.subckt decred_controller CLK_LED DATA_AVAILABLE[0] DATA_AVAILABLE[1] DATA_AVAILABLE[2]
+ DATA_AVAILABLE[3] DATA_AVAILABLE[4] DATA_AVAILABLE[5] DATA_FROM_HASH[0] DATA_FROM_HASH[1]
+ DATA_FROM_HASH[2] DATA_FROM_HASH[3] DATA_FROM_HASH[4] DATA_FROM_HASH[5] DATA_FROM_HASH[6]
+ DATA_FROM_HASH[7] DATA_TO_HASH[0] DATA_TO_HASH[1] DATA_TO_HASH[2] DATA_TO_HASH[3]
+ DATA_TO_HASH[4] DATA_TO_HASH[5] DATA_TO_HASH[6] DATA_TO_HASH[7] EXT_RESET_N_fromHost
+ EXT_RESET_N_toClient HASH_ADDR[0] HASH_ADDR[1] HASH_ADDR[2] HASH_ADDR[3] HASH_ADDR[4]
+ HASH_ADDR[5] HASH_EN HASH_LED ID_fromClient ID_toHost IRQ_OUT_fromClient IRQ_OUT_toHost
+ M1_CLK_IN M1_CLK_SELECT MACRO_RD_SELECT[0] MACRO_RD_SELECT[1] MACRO_RD_SELECT[2]
+ MACRO_RD_SELECT[3] MACRO_RD_SELECT[4] MACRO_RD_SELECT[5] MACRO_WR_SELECT[0] MACRO_WR_SELECT[1]
+ MACRO_WR_SELECT[2] MACRO_WR_SELECT[3] MACRO_WR_SELECT[4] MACRO_WR_SELECT[5] MISO_fromClient
+ MISO_toHost MOSI_fromHost MOSI_toClient PLL_INPUT S1_CLK_IN S1_CLK_SELECT SCLK_fromHost
+ SCLK_toClient SCSN_fromHost SCSN_toClient THREAD_COUNT[0] THREAD_COUNT[1] THREAD_COUNT[2]
+ THREAD_COUNT[3] m1_clk_local one zero vccd1 vssd1 vccd2_uq0 vccd2 vssd2 vdda1_uq0
+ vdda1 vssa1 vdda2_uq0 vdda2 vssa2
X_2037_ _2036_/Y _1980_/A _2027_/B _2026_/A _1990_/A vssd1 vssd1 vccd1 vccd1 _2039_/A
+ sky130_fd_sc_hd__a41o_4
XFILLER_39_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2106_ _2099_/X _2106_/B vssd1 vssd1 vccd1 vccd1 _2497_/D sky130_fd_sc_hd__and2_4
XFILLER_22_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1270_ _1295_/A _1300_/B vssd1 vssd1 vccd1 vccd1 _1270_/Y sky130_fd_sc_hd__nand2_4
XFILLER_44_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1606_ _1603_/X _1605_/Y vssd1 vssd1 vccd1 vccd1 _2660_/D sky130_fd_sc_hd__nand2_4
X_2655_ _2655_/CLK _1691_/Y vssd1 vssd1 vccd1 vccd1 _1675_/A sky130_fd_sc_hd__dfxtp_4
X_2586_ _2695_/CLK _1895_/X vssd1 vssd1 vccd1 vccd1 HASH_ADDR[1] sky130_fd_sc_hd__dfxtp_4
XFILLER_59_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1399_ _1382_/A _1255_/B _1381_/X _1382_/C vssd1 vssd1 vccd1 vccd1 _1407_/B sky130_fd_sc_hd__and4_4
X_1537_ _1521_/X _1533_/X _1536_/X vssd1 vssd1 vccd1 vccd1 _1537_/Y sky130_fd_sc_hd__a21oi_4
X_1468_ _1468_/A vssd1 vssd1 vccd1 vccd1 _1694_/A sky130_fd_sc_hd__buf_2
XFILLER_50_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2440_ _2495_/CLK _2440_/D vssd1 vssd1 vccd1 vccd1 _1751_/A sky130_fd_sc_hd__dfxtp_4
X_1322_ _1321_/Y _1313_/A vssd1 vssd1 vccd1 vccd1 _1327_/A sky130_fd_sc_hd__nor2_4
XFILLER_56_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2371_ _2371_/A vssd1 vssd1 vccd1 vccd1 _2371_/Y sky130_fd_sc_hd__inv_2
X_1253_ _1414_/A _2671_/Q _1413_/A _1414_/C vssd1 vssd1 vccd1 vccd1 _1254_/D sky130_fd_sc_hd__nand4_4
Xclkbuf_1_0_0_m1_clk_local clkbuf_0_m1_clk_local/X vssd1 vssd1 vccd1 vccd1 clkbuf_1_0_0_m1_clk_local/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_5_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2707_ _2707_/CLK _1214_/Y vssd1 vssd1 vccd1 vccd1 _1203_/A sky130_fd_sc_hd__dfxtp_4
X_2569_ _2561_/CLK _2569_/D vssd1 vssd1 vccd1 vccd1 _2569_/Q sky130_fd_sc_hd__dfxtp_4
X_2638_ _2511_/CLK _2638_/D vssd1 vssd1 vccd1 vccd1 _1522_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_59_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_4 _1976_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1871_ _1871_/A _1871_/B vssd1 vssd1 vccd1 vccd1 _1871_/X sky130_fd_sc_hd__and2_4
X_1940_ _1941_/A _1940_/B vssd1 vssd1 vccd1 vccd1 _2560_/D sky130_fd_sc_hd__and2_4
X_2423_ _2517_/CLK _2422_/Q vssd1 vssd1 vccd1 vccd1 _2423_/Q sky130_fd_sc_hd__dfxtp_4
X_1305_ _1305_/A vssd1 vssd1 vccd1 vccd1 _1305_/Y sky130_fd_sc_hd__inv_2
XFILLER_56_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1236_ _2263_/B _1208_/A _1222_/X vssd1 vssd1 vccd1 vccd1 _1236_/Y sky130_fd_sc_hd__o21ai_4
X_2285_ _2190_/A _2479_/Q vssd1 vssd1 vccd1 vccd1 _2285_/Y sky130_fd_sc_hd__nor2_4
Xclkbuf_0_m1_clk_local m1_clk_local vssd1 vssd1 vccd1 vccd1 clkbuf_0_m1_clk_local/X
+ sky130_fd_sc_hd__clkbuf_16
X_2354_ _2353_/X vssd1 vssd1 vccd1 vccd1 _2354_/X sky130_fd_sc_hd__buf_2
XFILLER_64_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2070_ _2069_/X vssd1 vssd1 vccd1 vccd1 _2520_/D sky130_fd_sc_hd__inv_2
XFILLER_38_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_3_3_0_m1_clk_local clkbuf_3_3_0_m1_clk_local/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_7_0_m1_clk_local/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_61_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1854_ _1842_/A vssd1 vssd1 vccd1 vccd1 _1858_/A sky130_fd_sc_hd__buf_2
XFILLER_61_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1923_ _1921_/A _1923_/B vssd1 vssd1 vccd1 vccd1 _2570_/D sky130_fd_sc_hd__nor2_4
X_1785_ _1775_/X _1784_/X _1777_/X vssd1 vssd1 vccd1 vccd1 _1785_/X sky130_fd_sc_hd__o21a_4
X_2406_ SCSN_fromHost vssd1 vssd1 vccd1 vccd1 SCSN_toClient sky130_fd_sc_hd__buf_2
XFILLER_55_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1219_ _1219_/A vssd1 vssd1 vccd1 vccd1 _1225_/B sky130_fd_sc_hd__buf_2
XFILLER_37_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2337_ _2334_/X _2117_/X _2453_/Q vssd1 vssd1 vccd1 vccd1 _2337_/Y sky130_fd_sc_hd__nand3_4
X_2199_ _2199_/A _2220_/B vssd1 vssd1 vccd1 vccd1 _2199_/Y sky130_fd_sc_hd__nand2_4
X_2268_ _2222_/A _1887_/A _2494_/Q vssd1 vssd1 vccd1 vccd1 _2268_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_40_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1570_ _1635_/A _1635_/B _1637_/C vssd1 vssd1 vccd1 vccd1 _1573_/A sky130_fd_sc_hd__nand3_4
XFILLER_6_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2053_ _1983_/A vssd1 vssd1 vccd1 vccd1 _2053_/X sky130_fd_sc_hd__buf_2
X_2122_ _2114_/Y _2120_/Y _2121_/Y vssd1 vssd1 vccd1 vccd1 _2491_/D sky130_fd_sc_hd__o21ai_4
XFILLER_13_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1906_ _1875_/A vssd1 vssd1 vccd1 vccd1 _1921_/A sky130_fd_sc_hd__buf_2
X_1837_ _1833_/Y _1836_/Y vssd1 vssd1 vccd1 vccd1 _2625_/D sky130_fd_sc_hd__nor2_4
X_1768_ _1768_/A _1768_/B vssd1 vssd1 vccd1 vccd1 _1768_/Y sky130_fd_sc_hd__nand2_4
X_1699_ _1521_/X _1693_/Y _1618_/Y _1694_/Y _1698_/Y vssd1 vssd1 vccd1 vccd1 _2654_/D
+ sky130_fd_sc_hd__a41oi_4
XFILLER_1_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1622_ _1664_/C vssd1 vssd1 vccd1 vccd1 _1633_/D sky130_fd_sc_hd__inv_2
X_2671_ _2679_/CLK _2671_/D vssd1 vssd1 vccd1 vccd1 _2671_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1484_ _1480_/Y _1482_/Y _1483_/X vssd1 vssd1 vccd1 vccd1 _2666_/D sky130_fd_sc_hd__a21oi_4
X_1553_ _2494_/Q vssd1 vssd1 vccd1 vccd1 _2221_/B sky130_fd_sc_hd__buf_2
X_2036_ _2035_/X vssd1 vssd1 vccd1 vccd1 _2036_/Y sky130_fd_sc_hd__inv_2
X_2105_ _1840_/A _2105_/B vssd1 vssd1 vccd1 vccd1 _2498_/D sky130_fd_sc_hd__nand2_4
XFILLER_10_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1605_ _2239_/A _2660_/Q vssd1 vssd1 vccd1 vccd1 _1605_/Y sky130_fd_sc_hd__nand2_4
X_1536_ _1457_/X _1535_/X _1474_/X vssd1 vssd1 vccd1 vccd1 _1536_/X sky130_fd_sc_hd__a21o_4
X_2654_ _2514_/CLK _2654_/D vssd1 vssd1 vccd1 vccd1 _2654_/Q sky130_fd_sc_hd__dfxtp_4
X_2585_ _2582_/CLK _2585_/D vssd1 vssd1 vccd1 vccd1 HASH_ADDR[0] sky130_fd_sc_hd__dfxtp_4
X_1398_ _1394_/Y _1395_/Y _1397_/X vssd1 vssd1 vccd1 vccd1 _2679_/D sky130_fd_sc_hd__a21oi_4
X_1467_ _1460_/A _1450_/B _1462_/X vssd1 vssd1 vccd1 vccd1 _1467_/Y sky130_fd_sc_hd__o21ai_4
X_2019_ _2008_/A _2007_/X _1363_/C vssd1 vssd1 vccd1 vccd1 _2019_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_42_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1321_ _1247_/B vssd1 vssd1 vccd1 vccd1 _1321_/Y sky130_fd_sc_hd__inv_2
XFILLER_49_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1252_ _2674_/Q _1252_/B vssd1 vssd1 vccd1 vccd1 _1254_/C sky130_fd_sc_hd__nand2_4
X_2370_ _1243_/X _1675_/A _1235_/X _1608_/B _2369_/Y vssd1 vssd1 vccd1 vccd1 _2370_/Y
+ sky130_fd_sc_hd__o41ai_4
XFILLER_64_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_3_4_0_addressalyzerBlock.SPI_CLK clkbuf_3_5_0_addressalyzerBlock.SPI_CLK/A
+ vssd1 vssd1 vccd1 vccd1 clkbuf_4_9_0_addressalyzerBlock.SPI_CLK/A sky130_fd_sc_hd__clkbuf_1
X_2706_ _2707_/CLK _2706_/D vssd1 vssd1 vccd1 vccd1 _2706_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_32_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2499_ _2707_/CLK _2499_/D vssd1 vssd1 vccd1 vccd1 _2499_/Q sky130_fd_sc_hd__dfxtp_4
X_1519_ _1471_/X _1472_/X _1518_/X vssd1 vssd1 vccd1 vccd1 _1519_/X sky130_fd_sc_hd__a21o_4
X_2568_ _2561_/CLK _1928_/Y vssd1 vssd1 vccd1 vccd1 _1940_/B sky130_fd_sc_hd__dfxtp_4
XINSDIODE2_5 _1937_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2637_ _2443_/CLK _2637_/D vssd1 vssd1 vccd1 vccd1 _1794_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_23_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1870_ _1871_/A _2605_/Q vssd1 vssd1 vccd1 vccd1 _2599_/D sky130_fd_sc_hd__and2_4
XFILLER_43_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2353_ _1590_/A _2353_/B _2111_/X _2353_/D vssd1 vssd1 vccd1 vccd1 _2353_/X sky130_fd_sc_hd__and4_4
X_2422_ _2517_/CLK _2421_/Q vssd1 vssd1 vccd1 vccd1 _2422_/Q sky130_fd_sc_hd__dfxtp_4
X_1304_ _1956_/A _1282_/B _1304_/C vssd1 vssd1 vccd1 vccd1 _1304_/Y sky130_fd_sc_hd__nor3_4
X_1235_ _1207_/A vssd1 vssd1 vccd1 vccd1 _1235_/X sky130_fd_sc_hd__buf_2
X_2284_ _2281_/Y _2282_/Y _2283_/Y vssd1 vssd1 vccd1 vccd1 _2284_/X sky130_fd_sc_hd__a21o_4
XFILLER_37_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1999_ _2008_/A _2008_/B _2003_/A vssd1 vssd1 vccd1 vccd1 _2000_/B sky130_fd_sc_hd__nor3_4
XFILLER_20_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1922_ _1922_/A vssd1 vssd1 vccd1 vccd1 _1923_/B sky130_fd_sc_hd__inv_2
X_1853_ _1853_/A _2621_/Q vssd1 vssd1 vccd1 vccd1 _2613_/D sky130_fd_sc_hd__and2_4
X_1784_ _1489_/A vssd1 vssd1 vccd1 vccd1 _1784_/X sky130_fd_sc_hd__buf_2
XFILLER_57_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2405_ SCLK_fromHost vssd1 vssd1 vccd1 vccd1 SCLK_toClient sky130_fd_sc_hd__buf_2
X_2336_ _1672_/Y _2333_/X _2335_/Y vssd1 vssd1 vccd1 vccd1 _2454_/D sky130_fd_sc_hd__o21ai_4
X_1218_ _1216_/Y _1208_/X _1217_/Y vssd1 vssd1 vccd1 vccd1 _2706_/D sky130_fd_sc_hd__a21oi_4
X_2198_ _2222_/A _2198_/B vssd1 vssd1 vccd1 vccd1 _2200_/A sky130_fd_sc_hd__nand2_4
X_2267_ _1978_/B _1647_/X _2266_/Y vssd1 vssd1 vccd1 vccd1 _2267_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_20_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2052_ _2051_/X _2023_/B _2035_/X vssd1 vssd1 vccd1 vccd1 _2525_/D sky130_fd_sc_hd__and3_4
X_2121_ _2114_/Y _2117_/X _1649_/A vssd1 vssd1 vccd1 vccd1 _2121_/Y sky130_fd_sc_hd__nand3_4
X_1905_ _1901_/A _1904_/Y vssd1 vssd1 vccd1 vccd1 _1905_/Y sky130_fd_sc_hd__nor2_4
XFILLER_22_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1698_ _2654_/Q _1695_/X _1697_/X vssd1 vssd1 vccd1 vccd1 _1698_/Y sky130_fd_sc_hd__o21ai_4
X_1836_ _1836_/A _1974_/C vssd1 vssd1 vccd1 vccd1 _1836_/Y sky130_fd_sc_hd__xnor2_4
X_1767_ _1766_/X _2659_/Q _1770_/C vssd1 vssd1 vccd1 vccd1 _1767_/Y sky130_fd_sc_hd__nand3_4
XFILLER_45_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2319_ _2318_/Y vssd1 vssd1 vccd1 vccd1 _2319_/Y sky130_fd_sc_hd__inv_2
XFILLER_40_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2670_ _2670_/CLK _2670_/D vssd1 vssd1 vccd1 vccd1 _1413_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_8_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1552_ _2335_/C _1546_/X _1548_/X _1551_/Y vssd1 vssd1 vccd1 vccd1 _1552_/X sky130_fd_sc_hd__a211o_4
X_1621_ _1617_/X _1620_/Y _1492_/X vssd1 vssd1 vccd1 vccd1 _2659_/D sky130_fd_sc_hd__a21oi_4
X_2104_ _1840_/A _2104_/B vssd1 vssd1 vccd1 vccd1 _2499_/D sky130_fd_sc_hd__nand2_4
X_1483_ _1458_/X _1444_/A _1474_/X vssd1 vssd1 vccd1 vccd1 _1483_/X sky130_fd_sc_hd__a21o_4
XFILLER_50_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2035_ _1989_/D vssd1 vssd1 vccd1 vccd1 _2035_/X sky130_fd_sc_hd__buf_2
X_1819_ _1203_/B _1819_/B _1822_/B vssd1 vssd1 vccd1 vccd1 _1819_/Y sky130_fd_sc_hd__nand3_4
XFILLER_53_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1604_ _2165_/A vssd1 vssd1 vccd1 vccd1 _2239_/A sky130_fd_sc_hd__buf_2
X_1535_ _1595_/A vssd1 vssd1 vccd1 vccd1 _1535_/X sky130_fd_sc_hd__buf_2
X_2584_ _2581_/CLK _1899_/Y vssd1 vssd1 vccd1 vccd1 _1911_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_8_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2653_ _2495_/CLK _1711_/X vssd1 vssd1 vccd1 vccd1 _2653_/Q sky130_fd_sc_hd__dfxtp_4
X_1397_ _1259_/B _2679_/Q _1396_/X _1256_/Y _1298_/X vssd1 vssd1 vccd1 vccd1 _1397_/X
+ sky130_fd_sc_hd__a41o_4
X_1466_ _1459_/X _1465_/Y _2375_/A vssd1 vssd1 vccd1 vccd1 _1466_/Y sky130_fd_sc_hd__a21oi_4
X_2018_ _2017_/Y vssd1 vssd1 vccd1 vccd1 _2534_/D sky130_fd_sc_hd__inv_2
XFILLER_6_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1320_ _1320_/A vssd1 vssd1 vccd1 vccd1 _1320_/Y sky130_fd_sc_hd__inv_2
X_1251_ _2672_/Q vssd1 vssd1 vccd1 vccd1 _1254_/B sky130_fd_sc_hd__inv_2
X_2705_ _2705_/CLK _2705_/D vssd1 vssd1 vccd1 vccd1 _1220_/A sky130_fd_sc_hd__dfxtp_4
X_2636_ _2443_/CLK _2636_/D vssd1 vssd1 vccd1 vccd1 _2636_/Q sky130_fd_sc_hd__dfxtp_4
XINSDIODE2_6 _1936_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2498_ _2707_/CLK _2498_/D vssd1 vssd1 vccd1 vccd1 _2089_/A sky130_fd_sc_hd__dfxtp_4
X_1518_ _1516_/X _1508_/Y _1488_/X _1517_/Y _1469_/X vssd1 vssd1 vccd1 vccd1 _1518_/X
+ sky130_fd_sc_hd__o32a_4
X_2567_ _2581_/CLK _1930_/Y vssd1 vssd1 vccd1 vccd1 _2567_/Q sky130_fd_sc_hd__dfxtp_4
X_1449_ _1448_/Y vssd1 vssd1 vccd1 vccd1 _1450_/D sky130_fd_sc_hd__buf_2
XFILLER_55_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1303_ _1246_/Y _1247_/Y _1281_/C _1313_/A _1276_/Y vssd1 vssd1 vccd1 vccd1 _1304_/C
+ sky130_fd_sc_hd__o41a_4
X_2283_ _2395_/A _2187_/B _2187_/C vssd1 vssd1 vccd1 vccd1 _2283_/Y sky130_fd_sc_hd__nor3_4
X_2352_ _2351_/X vssd1 vssd1 vccd1 vccd1 _2352_/X sky130_fd_sc_hd__buf_2
X_2421_ _2420_/CLK _2421_/D vssd1 vssd1 vccd1 vccd1 _2421_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_64_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1234_ _1238_/C _1201_/A _1233_/X vssd1 vssd1 vccd1 vccd1 _1234_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_49_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2619_ _2621_/CLK _1846_/X vssd1 vssd1 vccd1 vccd1 _1856_/B sky130_fd_sc_hd__dfxtp_4
X_1998_ _2534_/Q vssd1 vssd1 vccd1 vccd1 _2008_/B sky130_fd_sc_hd__inv_2
XPHY_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1852_ _1853_/A _2622_/Q vssd1 vssd1 vccd1 vccd1 _2614_/D sky130_fd_sc_hd__and2_4
XFILLER_46_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1921_ _1921_/A _1921_/B vssd1 vssd1 vccd1 vccd1 _1921_/Y sky130_fd_sc_hd__nor2_4
X_1783_ _1964_/B _2634_/Q _1782_/X vssd1 vssd1 vccd1 vccd1 _1783_/X sky130_fd_sc_hd__o21a_4
XFILLER_6_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2404_ MOSI_fromHost vssd1 vssd1 vccd1 vccd1 MOSI_toClient sky130_fd_sc_hd__buf_2
XFILLER_57_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2335_ _2334_/X _2117_/X _2335_/C vssd1 vssd1 vccd1 vccd1 _2335_/Y sky130_fd_sc_hd__nand3_4
X_2266_ _2194_/X _1909_/A _2250_/B vssd1 vssd1 vccd1 vccd1 _2266_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_52_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1217_ _2165_/B _1209_/X _1212_/X vssd1 vssd1 vccd1 vccd1 _1217_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_37_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2197_ _2197_/A _2221_/B _2197_/C vssd1 vssd1 vccd1 vccd1 _2197_/Y sky130_fd_sc_hd__nand3_4
XFILLER_48_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2120_ _1829_/B _2115_/X _1694_/A vssd1 vssd1 vccd1 vccd1 _2120_/Y sky130_fd_sc_hd__nand3_4
X_2051_ _2057_/A _2057_/B _2057_/C _1988_/C _1988_/D vssd1 vssd1 vccd1 vccd1 _2051_/X
+ sky130_fd_sc_hd__a41o_4
XFILLER_30_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1904_ _1904_/A vssd1 vssd1 vccd1 vccd1 _1904_/Y sky130_fd_sc_hd__inv_2
X_1835_ _1966_/A _2542_/Q _1966_/B vssd1 vssd1 vccd1 vccd1 _1974_/C sky130_fd_sc_hd__nor3_4
XFILLER_15_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1697_ _1838_/A vssd1 vssd1 vccd1 vccd1 _1697_/X sky130_fd_sc_hd__buf_2
X_1766_ _1770_/B _1770_/D _1683_/D vssd1 vssd1 vccd1 vccd1 _1766_/X sky130_fd_sc_hd__a21o_4
X_2318_ _1656_/X _2112_/X vssd1 vssd1 vccd1 vccd1 _2318_/Y sky130_fd_sc_hd__nor2_4
X_2249_ _2249_/A _1546_/A vssd1 vssd1 vccd1 vccd1 _2249_/Y sky130_fd_sc_hd__nand2_4
XFILLER_65_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1620_ _2381_/B _1620_/B _2381_/C _1614_/Y vssd1 vssd1 vccd1 vccd1 _1620_/Y sky130_fd_sc_hd__nand4_4
X_1482_ _1481_/X _1470_/Y _1471_/X _1472_/X vssd1 vssd1 vccd1 vccd1 _1482_/Y sky130_fd_sc_hd__a22oi_4
XFILLER_8_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1551_ _2143_/A _1550_/Y vssd1 vssd1 vccd1 vccd1 _1551_/Y sky130_fd_sc_hd__nor2_4
X_2103_ _2099_/X MOSI_fromHost vssd1 vssd1 vccd1 vccd1 _2500_/D sky130_fd_sc_hd__and2_4
XFILLER_62_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2034_ _2034_/A vssd1 vssd1 vccd1 vccd1 _2034_/Y sky130_fd_sc_hd__inv_2
XFILLER_47_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1818_ _1747_/A vssd1 vssd1 vccd1 vccd1 _1818_/Y sky130_fd_sc_hd__inv_2
X_1749_ _1748_/Y vssd1 vssd1 vccd1 vccd1 _1749_/Y sky130_fd_sc_hd__inv_2
XFILLER_26_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_4_0_addressalyzerBlock.SPI_CLK clkbuf_4_5_0_addressalyzerBlock.SPI_CLK/A
+ vssd1 vssd1 vccd1 vccd1 _2443_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_3_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2652_ _2655_/CLK _1723_/Y vssd1 vssd1 vccd1 vccd1 _2652_/Q sky130_fd_sc_hd__dfxtp_4
X_1603_ _1585_/Y _1593_/Y _1602_/X vssd1 vssd1 vccd1 vccd1 _1603_/X sky130_fd_sc_hd__a21o_4
X_1465_ _1458_/X _1462_/X _1464_/X vssd1 vssd1 vccd1 vccd1 _1465_/Y sky130_fd_sc_hd__o21ai_4
X_1534_ _1442_/A vssd1 vssd1 vccd1 vccd1 _1595_/A sky130_fd_sc_hd__inv_2
X_2583_ _2679_/CLK _1901_/Y vssd1 vssd1 vccd1 vccd1 _1912_/B sky130_fd_sc_hd__dfxtp_4
X_2017_ _2017_/A _2005_/B _2016_/Y vssd1 vssd1 vccd1 vccd1 _2017_/Y sky130_fd_sc_hd__nand3_4
X_1396_ _1381_/X vssd1 vssd1 vccd1 vccd1 _1396_/X sky130_fd_sc_hd__buf_2
XFILLER_10_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1250_ _1382_/C vssd1 vssd1 vccd1 vccd1 _1254_/A sky130_fd_sc_hd__inv_2
XFILLER_24_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2704_ _2617_/CLK _2704_/D vssd1 vssd1 vccd1 vccd1 _1225_/A sky130_fd_sc_hd__dfxtp_4
Xclkbuf_4_8_0_m1_clk_local clkbuf_4_9_0_m1_clk_local/A vssd1 vssd1 vccd1 vccd1 _2527_/CLK
+ sky130_fd_sc_hd__clkbuf_1
X_2635_ _2443_/CLK _1803_/X vssd1 vssd1 vccd1 vccd1 _2635_/Q sky130_fd_sc_hd__dfxtp_4
X_1448_ _1478_/A vssd1 vssd1 vccd1 vccd1 _1448_/Y sky130_fd_sc_hd__inv_2
X_2566_ _2561_/CLK _1932_/Y vssd1 vssd1 vccd1 vccd1 _1942_/B sky130_fd_sc_hd__dfxtp_4
X_1517_ _1517_/A vssd1 vssd1 vccd1 vccd1 _1517_/Y sky130_fd_sc_hd__inv_2
X_2497_ _2655_/CLK _2497_/D vssd1 vssd1 vccd1 vccd1 _1770_/C sky130_fd_sc_hd__dfxtp_4
X_1379_ _1249_/A _1377_/Y _1378_/X vssd1 vssd1 vccd1 vccd1 _1385_/A sky130_fd_sc_hd__o21a_4
XFILLER_23_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2420_ _2420_/CLK _2419_/Q vssd1 vssd1 vccd1 vccd1 _2421_/D sky130_fd_sc_hd__dfxtp_4
X_1302_ _1956_/A _1302_/B _1302_/C vssd1 vssd1 vccd1 vccd1 _2697_/D sky130_fd_sc_hd__nor3_4
X_1233_ _1233_/A _1225_/B vssd1 vssd1 vccd1 vccd1 _1233_/X sky130_fd_sc_hd__or2_4
X_2282_ THREAD_COUNT[0] _2260_/A _2162_/A vssd1 vssd1 vccd1 vccd1 _2282_/Y sky130_fd_sc_hd__a21oi_4
X_2351_ _1527_/X _1535_/X _2111_/X _1631_/A _1668_/A vssd1 vssd1 vccd1 vccd1 _2351_/X
+ sky130_fd_sc_hd__a41o_4
XFILLER_29_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1997_ _1979_/Y vssd1 vssd1 vccd1 vccd1 _2008_/A sky130_fd_sc_hd__buf_2
X_2618_ _2621_/CLK _1847_/X vssd1 vssd1 vccd1 vccd1 _1857_/B sky130_fd_sc_hd__dfxtp_4
X_2549_ _2561_/CLK _2549_/D vssd1 vssd1 vccd1 vccd1 MACRO_WR_SELECT[4] sky130_fd_sc_hd__dfxtp_4
XFILLER_9_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0_addressalyzerBlock.SPI_CLK clkbuf_0_addressalyzerBlock.SPI_CLK/X vssd1
+ vssd1 vccd1 vccd1 clkbuf_1_0_0_addressalyzerBlock.SPI_CLK/X sky130_fd_sc_hd__clkbuf_1
XFILLER_34_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1851_ _1853_/A _2623_/Q vssd1 vssd1 vccd1 vccd1 _2615_/D sky130_fd_sc_hd__and2_4
X_1920_ _2469_/Q vssd1 vssd1 vccd1 vccd1 _1921_/B sky130_fd_sc_hd__inv_2
X_2403_ EXT_RESET_N_fromHost vssd1 vssd1 vccd1 vccd1 EXT_RESET_N_toClient sky130_fd_sc_hd__buf_2
X_1782_ _1775_/X _1481_/X _1777_/X vssd1 vssd1 vccd1 vccd1 _1782_/X sky130_fd_sc_hd__o21a_4
X_1216_ _1220_/A _1201_/X _1215_/X vssd1 vssd1 vccd1 vccd1 _1216_/Y sky130_fd_sc_hd__o21ai_4
X_2265_ _1500_/X _1594_/C _1255_/B _1592_/X vssd1 vssd1 vccd1 vccd1 _2265_/X sky130_fd_sc_hd__a2bb2o_4
X_2196_ HASH_LED _2220_/B vssd1 vssd1 vccd1 vccd1 _2197_/C sky130_fd_sc_hd__nand2_4
X_2334_ _2346_/A vssd1 vssd1 vccd1 vccd1 _2334_/X sky130_fd_sc_hd__buf_2
XFILLER_25_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2050_ _1988_/A vssd1 vssd1 vccd1 vccd1 _2057_/C sky130_fd_sc_hd__buf_2
XFILLER_10_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1834_ _1974_/A _2541_/Q vssd1 vssd1 vccd1 vccd1 _1966_/B sky130_fd_sc_hd__nand2_4
X_1903_ _1901_/A _1902_/Y vssd1 vssd1 vccd1 vccd1 _1903_/Y sky130_fd_sc_hd__nor2_4
X_1765_ _1765_/A _1765_/B _1765_/C _1765_/D vssd1 vssd1 vccd1 vccd1 _1770_/D sky130_fd_sc_hd__and4_4
X_1696_ _2353_/B vssd1 vssd1 vccd1 vccd1 _1838_/A sky130_fd_sc_hd__buf_2
XFILLER_57_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2317_ _1516_/X vssd1 vssd1 vccd1 vccd1 _2317_/X sky130_fd_sc_hd__buf_2
X_2179_ _2176_/Y _1560_/X _2178_/X vssd1 vssd1 vccd1 vccd1 _2179_/Y sky130_fd_sc_hd__a21boi_4
X_2248_ _2248_/A _2472_/Q vssd1 vssd1 vccd1 vccd1 _2250_/A sky130_fd_sc_hd__nand2_4
XFILLER_21_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1550_ _2462_/Q vssd1 vssd1 vccd1 vccd1 _1550_/Y sky130_fd_sc_hd__inv_2
X_1481_ _1481_/A vssd1 vssd1 vccd1 vccd1 _1481_/X sky130_fd_sc_hd__buf_2
X_2033_ _2031_/X _2032_/Y vssd1 vssd1 vccd1 vccd1 _2034_/A sky130_fd_sc_hd__nand2_4
XFILLER_39_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2102_ _2099_/X _2102_/B vssd1 vssd1 vccd1 vccd1 _2102_/X sky130_fd_sc_hd__and2_4
XFILLER_11_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1748_ _1668_/A _1828_/A vssd1 vssd1 vccd1 vccd1 _1748_/Y sky130_fd_sc_hd__nor2_4
X_1817_ _1798_/A _2501_/Q _1816_/X vssd1 vssd1 vccd1 vccd1 _2629_/D sky130_fd_sc_hd__o21a_4
X_1679_ _2653_/Q vssd1 vssd1 vccd1 vccd1 _1707_/A sky130_fd_sc_hd__buf_2
XFILLER_53_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1602_ _1594_/Y _2260_/A _1602_/C vssd1 vssd1 vccd1 vccd1 _1602_/X sky130_fd_sc_hd__or3_4
X_2651_ _2514_/CLK _2651_/D vssd1 vssd1 vccd1 vccd1 _2651_/Q sky130_fd_sc_hd__dfxtp_4
X_2582_ _2582_/CLK _1903_/Y vssd1 vssd1 vccd1 vccd1 _1913_/B sky130_fd_sc_hd__dfxtp_4
X_1464_ _1463_/X vssd1 vssd1 vccd1 vccd1 _1464_/X sky130_fd_sc_hd__buf_2
X_1395_ _2679_/Q vssd1 vssd1 vccd1 vccd1 _1395_/Y sky130_fd_sc_hd__inv_2
X_1533_ _1531_/X _1478_/X _1532_/Y _1469_/X vssd1 vssd1 vccd1 vccd1 _1533_/X sky130_fd_sc_hd__o22a_4
X_2016_ _2008_/A _2007_/X _2008_/B vssd1 vssd1 vccd1 vccd1 _2016_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_2_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2703_ _2617_/CLK _2703_/D vssd1 vssd1 vccd1 vccd1 _2703_/Q sky130_fd_sc_hd__dfxtp_4
X_1516_ _1515_/X vssd1 vssd1 vccd1 vccd1 _1516_/X sky130_fd_sc_hd__buf_2
X_2565_ _2581_/CLK _2565_/D vssd1 vssd1 vccd1 vccd1 _2565_/Q sky130_fd_sc_hd__dfxtp_4
X_2634_ _2443_/CLK _2634_/D vssd1 vssd1 vccd1 vccd1 _2634_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_59_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1378_ _1378_/A vssd1 vssd1 vccd1 vccd1 _1378_/X sky130_fd_sc_hd__buf_2
X_1447_ _1446_/Y vssd1 vssd1 vccd1 vccd1 _1478_/A sky130_fd_sc_hd__buf_2
XFILLER_4_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2496_ _2655_/CLK _2496_/D vssd1 vssd1 vccd1 vccd1 _2106_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_23_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1232_ _1230_/Y _1208_/X _1231_/Y vssd1 vssd1 vccd1 vccd1 _2703_/D sky130_fd_sc_hd__a21oi_4
X_1301_ _1305_/A _1268_/X _1300_/B vssd1 vssd1 vccd1 vccd1 _1302_/C sky130_fd_sc_hd__a21oi_4
X_2281_ _2265_/X _2279_/Y _2280_/X vssd1 vssd1 vccd1 vccd1 _2281_/Y sky130_fd_sc_hd__o21ai_4
X_2350_ _1978_/B _2341_/X _2137_/C _2331_/Y vssd1 vssd1 vccd1 vccd1 _2350_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_1_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1996_ _1996_/A _1995_/Y vssd1 vssd1 vccd1 vccd1 _2001_/A sky130_fd_sc_hd__nand2_4
X_2617_ _2617_/CLK _1849_/X vssd1 vssd1 vccd1 vccd1 _1858_/B sky130_fd_sc_hd__dfxtp_4
X_2548_ _2553_/CLK _2548_/D vssd1 vssd1 vccd1 vccd1 MACRO_WR_SELECT[3] sky130_fd_sc_hd__dfxtp_4
XFILLER_55_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2479_ _2707_/CLK _2479_/D vssd1 vssd1 vccd1 vccd1 _2479_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_18_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1850_ _1853_/A _1850_/B vssd1 vssd1 vccd1 vccd1 _1850_/X sky130_fd_sc_hd__and2_4
XFILLER_42_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1781_ _1964_/B _2635_/Q _1780_/X vssd1 vssd1 vccd1 vccd1 _1781_/X sky130_fd_sc_hd__o21a_4
XFILLER_41_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2402_ vssd1 vssd1 vccd1 vccd1 _2402_/HI zero sky130_fd_sc_hd__conb_1
X_2333_ _2346_/A vssd1 vssd1 vccd1 vccd1 _2333_/X sky130_fd_sc_hd__buf_2
X_2264_ _2262_/Y _2263_/Y vssd1 vssd1 vccd1 vccd1 _2480_/D sky130_fd_sc_hd__nand2_4
X_1215_ _2706_/Q _1203_/B vssd1 vssd1 vccd1 vccd1 _1215_/X sky130_fd_sc_hd__or2_4
XFILLER_37_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2195_ _2194_/X _2195_/B vssd1 vssd1 vccd1 vccd1 _2197_/A sky130_fd_sc_hd__nand2_4
XFILLER_60_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1979_ _1979_/A vssd1 vssd1 vccd1 vccd1 _1979_/Y sky130_fd_sc_hd__inv_2
XFILLER_29_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1902_ _2195_/B vssd1 vssd1 vccd1 vccd1 _1902_/Y sky130_fd_sc_hd__inv_2
XFILLER_30_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1764_ _1738_/Y _1751_/A _1717_/C _1761_/Y vssd1 vssd1 vccd1 vccd1 _1765_/D sky130_fd_sc_hd__a22oi_4
X_1833_ _1833_/A _2408_/Q _1833_/C vssd1 vssd1 vccd1 vccd1 _1833_/Y sky130_fd_sc_hd__nor3_4
X_2316_ _1934_/B _2305_/X _2137_/C _2307_/X vssd1 vssd1 vccd1 vccd1 _2463_/D sky130_fd_sc_hd__a2bb2o_4
X_1695_ _1685_/Y vssd1 vssd1 vccd1 vccd1 _1695_/X sky130_fd_sc_hd__buf_2
XFILLER_57_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2247_ _2247_/A _2221_/B _2247_/C vssd1 vssd1 vccd1 vccd1 _2251_/A sky130_fd_sc_hd__nand3_4
X_2178_ _1947_/A _2147_/B _1559_/X _2177_/Y vssd1 vssd1 vccd1 vccd1 _2178_/X sky130_fd_sc_hd__a211o_4
XFILLER_40_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_4_9_0_addressalyzerBlock.SPI_CLK clkbuf_4_9_0_addressalyzerBlock.SPI_CLK/A
+ vssd1 vssd1 vccd1 vccd1 _2705_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1480_ _1676_/D _1477_/Y _1479_/Y vssd1 vssd1 vccd1 vccd1 _1480_/Y sky130_fd_sc_hd__o21ai_4
X_2032_ _2026_/X _2012_/A _1990_/A _1990_/B vssd1 vssd1 vccd1 vccd1 _2032_/Y sky130_fd_sc_hd__nand4_4
XFILLER_47_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2101_ _2099_/X SCLK_fromHost vssd1 vssd1 vccd1 vccd1 _2101_/X sky130_fd_sc_hd__and2_4
X_1816_ _2629_/Q _2507_/Q _1815_/X vssd1 vssd1 vccd1 vccd1 _1816_/X sky130_fd_sc_hd__o21a_4
X_1747_ _1747_/A _1203_/B _1819_/B _1822_/B vssd1 vssd1 vccd1 vccd1 _1747_/Y sky130_fd_sc_hd__nand4_4
X_1678_ _2652_/Q _2651_/Q _1715_/A _1738_/A vssd1 vssd1 vccd1 vccd1 _1707_/D sky130_fd_sc_hd__and4_4
XFILLER_38_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1601_ _1600_/Y vssd1 vssd1 vccd1 vccd1 _1602_/C sky130_fd_sc_hd__inv_2
X_2581_ _2581_/CLK _1905_/Y vssd1 vssd1 vccd1 vccd1 _1914_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_8_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1532_ _1794_/A vssd1 vssd1 vccd1 vccd1 _1532_/Y sky130_fd_sc_hd__inv_2
X_2650_ _2495_/CLK _2650_/D vssd1 vssd1 vccd1 vccd1 _1715_/A sky130_fd_sc_hd__dfxtp_4
X_1463_ _1652_/A vssd1 vssd1 vccd1 vccd1 _1463_/X sky130_fd_sc_hd__buf_2
X_1394_ _1394_/A vssd1 vssd1 vccd1 vccd1 _1394_/Y sky130_fd_sc_hd__inv_2
XFILLER_4_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2015_ _2000_/B vssd1 vssd1 vccd1 vccd1 _2017_/A sky130_fd_sc_hd__inv_2
XFILLER_35_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_2_1_0_m1_clk_local clkbuf_1_0_0_m1_clk_local/X vssd1 vssd1 vccd1 vccd1 clkbuf_3_3_0_m1_clk_local/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_53_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2702_ _2705_/CLK _1237_/Y vssd1 vssd1 vccd1 vccd1 _1233_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_32_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_2_0_0_addressalyzerBlock.SPI_CLK clkbuf_1_0_0_addressalyzerBlock.SPI_CLK/X
+ vssd1 vssd1 vccd1 vccd1 clkbuf_3_1_0_addressalyzerBlock.SPI_CLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_20_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2564_ _2564_/CLK _1935_/X vssd1 vssd1 vccd1 vccd1 DATA_TO_HASH[7] sky130_fd_sc_hd__dfxtp_4
X_1515_ _1515_/A vssd1 vssd1 vccd1 vccd1 _1515_/X sky130_fd_sc_hd__buf_2
X_2495_ _2495_/CLK _2495_/D vssd1 vssd1 vccd1 vccd1 _2495_/Q sky130_fd_sc_hd__dfxtp_4
X_2633_ _2443_/CLK _2633_/D vssd1 vssd1 vccd1 vccd1 _2633_/Q sky130_fd_sc_hd__dfxtp_4
X_1377_ _1377_/A _1377_/B vssd1 vssd1 vccd1 vccd1 _1377_/Y sky130_fd_sc_hd__nor2_4
X_1446_ _2371_/A _1507_/A vssd1 vssd1 vccd1 vccd1 _1446_/Y sky130_fd_sc_hd__nor2_4
XFILLER_4_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1300_ _1285_/Y _1300_/B _1268_/X _2695_/Q vssd1 vssd1 vccd1 vccd1 _1302_/B sky130_fd_sc_hd__and4_4
X_1231_ _2481_/Q _1208_/A _1222_/X vssd1 vssd1 vccd1 vccd1 _1231_/Y sky130_fd_sc_hd__o21ai_4
X_2280_ _1414_/C _1656_/X _2158_/X _2112_/X _2154_/X vssd1 vssd1 vccd1 vccd1 _2280_/X
+ sky130_fd_sc_hd__a2111o_4
XFILLER_45_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1995_ CLK_LED vssd1 vssd1 vccd1 vccd1 _1995_/Y sky130_fd_sc_hd__inv_2
X_2616_ _2617_/CLK _1850_/X vssd1 vssd1 vccd1 vccd1 _1568_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_20_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2547_ _2699_/CLK _1961_/X vssd1 vssd1 vccd1 vccd1 MACRO_WR_SELECT[2] sky130_fd_sc_hd__dfxtp_4
X_1429_ _2671_/Q _1415_/Y vssd1 vssd1 vccd1 vccd1 _1429_/X sky130_fd_sc_hd__or2_4
X_2478_ _2478_/CLK _2295_/Y vssd1 vssd1 vccd1 vccd1 _1554_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_55_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_4_0_m1_clk_local clkbuf_4_5_0_m1_clk_local/A vssd1 vssd1 vccd1 vccd1 _2413_/CLK
+ sky130_fd_sc_hd__clkbuf_1
XPHY_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1780_ _1775_/X _1694_/A _1777_/X vssd1 vssd1 vccd1 vccd1 _1780_/X sky130_fd_sc_hd__o21a_4
X_2401_ vssd1 vssd1 vccd1 vccd1 one _2401_/LO sky130_fd_sc_hd__conb_1
XFILLER_34_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2332_ _2331_/Y vssd1 vssd1 vccd1 vccd1 _2346_/A sky130_fd_sc_hd__inv_2
X_2263_ _2239_/A _2263_/B vssd1 vssd1 vccd1 vccd1 _2263_/Y sky130_fd_sc_hd__nand2_4
X_1214_ _1204_/Y _1208_/X _1213_/Y vssd1 vssd1 vccd1 vccd1 _1214_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_37_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2194_ _2248_/A vssd1 vssd1 vccd1 vccd1 _2194_/X sky130_fd_sc_hd__buf_2
X_1978_ _1956_/A _1978_/B vssd1 vssd1 vccd1 vccd1 _1978_/Y sky130_fd_sc_hd__nor2_4
XFILLER_20_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1901_ _1901_/A _1901_/B vssd1 vssd1 vccd1 vccd1 _1901_/Y sky130_fd_sc_hd__nor2_4
XFILLER_15_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1832_ _1832_/A vssd1 vssd1 vccd1 vccd1 _1833_/C sky130_fd_sc_hd__inv_2
X_1694_ _1694_/A _2378_/B vssd1 vssd1 vccd1 vccd1 _1694_/Y sky130_fd_sc_hd__nand2_4
X_1763_ _2177_/B _2652_/Q _1712_/X _1758_/Y vssd1 vssd1 vccd1 vccd1 _1765_/C sky130_fd_sc_hd__a22oi_4
X_2315_ _1932_/B _2305_/X _1522_/A _2307_/X vssd1 vssd1 vccd1 vccd1 _2464_/D sky130_fd_sc_hd__a2bb2o_4
X_2246_ _2348_/C _2220_/B vssd1 vssd1 vccd1 vccd1 _2247_/C sky130_fd_sc_hd__nand2_4
X_2177_ _2272_/A _2177_/B vssd1 vssd1 vccd1 vccd1 _2177_/Y sky130_fd_sc_hd__nor2_4
Xclkbuf_4_14_0_addressalyzerBlock.SPI_CLK clkbuf_3_7_0_addressalyzerBlock.SPI_CLK/X
+ vssd1 vssd1 vccd1 vccd1 _2438_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_31_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2100_ _2099_/X _2100_/B vssd1 vssd1 vccd1 vccd1 _2100_/X sky130_fd_sc_hd__and2_4
XFILLER_62_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2031_ _1990_/B _2030_/X _1378_/X vssd1 vssd1 vccd1 vccd1 _2031_/X sky130_fd_sc_hd__o21a_4
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1815_ _1838_/A vssd1 vssd1 vccd1 vccd1 _1815_/X sky130_fd_sc_hd__buf_2
X_1746_ _1742_/Y _1744_/X _1745_/X vssd1 vssd1 vccd1 vccd1 _2648_/D sky130_fd_sc_hd__o21a_4
XFILLER_7_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1677_ _1676_/X vssd1 vssd1 vccd1 vccd1 _1683_/B sky130_fd_sc_hd__buf_2
X_2229_ _1439_/A _2611_/Q _1577_/A _2149_/X vssd1 vssd1 vccd1 vccd1 _2229_/X sky130_fd_sc_hd__o22a_4
XFILLER_53_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1531_ _1530_/X vssd1 vssd1 vccd1 vccd1 _1531_/X sky130_fd_sc_hd__buf_2
X_1600_ _2165_/A _1600_/B vssd1 vssd1 vccd1 vccd1 _1600_/Y sky130_fd_sc_hd__nor2_4
X_1462_ _1460_/Y _1444_/A _1444_/B _1486_/B _1450_/D vssd1 vssd1 vccd1 vccd1 _1462_/X
+ sky130_fd_sc_hd__o41a_4
X_2580_ _2582_/CLK _1908_/Y vssd1 vssd1 vccd1 vccd1 _1916_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_8_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1393_ _1392_/Y vssd1 vssd1 vccd1 vccd1 _1393_/Y sky130_fd_sc_hd__inv_2
X_2014_ _2014_/A _2014_/B _2014_/C vssd1 vssd1 vccd1 vccd1 _2014_/Y sky130_fd_sc_hd__nor3_4
XFILLER_50_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1729_ _1717_/C vssd1 vssd1 vccd1 vccd1 _1730_/A sky130_fd_sc_hd__inv_2
XFILLER_58_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2701_ _2707_/CLK _1245_/Y vssd1 vssd1 vccd1 vccd1 _1238_/C sky130_fd_sc_hd__dfxtp_4
X_2632_ _2511_/CLK _2632_/D vssd1 vssd1 vccd1 vccd1 _2632_/Q sky130_fd_sc_hd__dfxtp_4
X_2563_ _2695_/CLK _1936_/X vssd1 vssd1 vccd1 vccd1 DATA_TO_HASH[6] sky130_fd_sc_hd__dfxtp_4
X_1514_ _1510_/A vssd1 vssd1 vccd1 vccd1 _1515_/A sky130_fd_sc_hd__buf_2
X_1445_ _1540_/B vssd1 vssd1 vccd1 vccd1 _1460_/A sky130_fd_sc_hd__buf_2
X_2494_ _2494_/CLK _2494_/D vssd1 vssd1 vccd1 vccd1 _2494_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_55_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1376_ _1249_/B vssd1 vssd1 vccd1 vccd1 _1377_/A sky130_fd_sc_hd__inv_2
Xclkbuf_4_12_0_m1_clk_local clkbuf_3_6_0_m1_clk_local/X vssd1 vssd1 vccd1 vccd1 _2693_/CLK
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_23_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1230_ _1233_/A _1201_/A _1229_/X vssd1 vssd1 vccd1 vccd1 _1230_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_49_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1994_ _2534_/Q _1993_/Y _2000_/A _2536_/Q vssd1 vssd1 vccd1 vccd1 _1996_/A sky130_fd_sc_hd__nand4_4
X_2615_ _2617_/CLK _2615_/D vssd1 vssd1 vccd1 vccd1 _1653_/B sky130_fd_sc_hd__dfxtp_4
X_2546_ _2695_/CLK _1962_/X vssd1 vssd1 vccd1 vccd1 MACRO_WR_SELECT[1] sky130_fd_sc_hd__dfxtp_4
X_1428_ _2014_/A _1419_/A _1428_/C vssd1 vssd1 vccd1 vccd1 _1428_/Y sky130_fd_sc_hd__nor3_4
X_2477_ _2478_/CLK _2297_/Y vssd1 vssd1 vccd1 vccd1 _2477_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1359_ _1355_/B _1350_/Y _1358_/Y vssd1 vssd1 vccd1 vccd1 _2686_/D sky130_fd_sc_hd__o21a_4
XFILLER_28_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2400_ _2398_/Y _1235_/X _2399_/Y vssd1 vssd1 vccd1 vccd1 _2400_/Y sky130_fd_sc_hd__a21oi_4
X_2262_ _2241_/X _2261_/Y _2189_/X vssd1 vssd1 vccd1 vccd1 _2262_/Y sky130_fd_sc_hd__o21ai_4
X_1213_ _1662_/B _1209_/X _1212_/X vssd1 vssd1 vccd1 vccd1 _1213_/Y sky130_fd_sc_hd__o21ai_4
X_2331_ _2331_/A _1515_/X _1626_/Y _1508_/Y vssd1 vssd1 vccd1 vccd1 _2331_/Y sky130_fd_sc_hd__nor4_4
X_2193_ _1500_/A _2154_/X _1257_/A _1592_/X vssd1 vssd1 vccd1 vccd1 _2193_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_1_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1977_ _2447_/Q vssd1 vssd1 vccd1 vccd1 _1978_/B sky130_fd_sc_hd__inv_2
X_2529_ _2564_/CLK _2039_/X vssd1 vssd1 vccd1 vccd1 _1990_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_29_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1900_ _1900_/A vssd1 vssd1 vccd1 vccd1 _1901_/B sky130_fd_sc_hd__inv_2
X_1831_ _1203_/B _1822_/B _1830_/Y vssd1 vssd1 vccd1 vccd1 _2626_/D sky130_fd_sc_hd__o21a_4
X_1762_ _2652_/Q _2177_/B _1715_/A _1761_/Y vssd1 vssd1 vccd1 vccd1 _1765_/B sky130_fd_sc_hd__o22a_4
X_1693_ _2654_/Q _1692_/X _1689_/Y vssd1 vssd1 vccd1 vccd1 _1693_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_65_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2314_ _1929_/Y _2305_/X _1517_/A _2307_/X vssd1 vssd1 vccd1 vccd1 _2465_/D sky130_fd_sc_hd__a2bb2o_4
X_2245_ _2222_/A _2245_/B vssd1 vssd1 vccd1 vccd1 _2247_/A sky130_fd_sc_hd__nand2_4
X_2176_ _2172_/Y _2175_/Y vssd1 vssd1 vccd1 vccd1 _2176_/Y sky130_fd_sc_hd__nand2_4
XFILLER_31_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2030_ _2027_/A _2027_/B _2026_/A _1990_/A vssd1 vssd1 vccd1 vccd1 _2030_/X sky130_fd_sc_hd__and4_4
XFILLER_47_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1745_ _1707_/C _1685_/Y _1697_/X vssd1 vssd1 vccd1 vccd1 _1745_/X sky130_fd_sc_hd__o21a_4
X_1814_ _2629_/Q _1798_/A _1813_/X vssd1 vssd1 vccd1 vccd1 _2630_/D sky130_fd_sc_hd__o21a_4
XFILLER_15_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1676_ _1477_/Y _1652_/A _1540_/B _1676_/D vssd1 vssd1 vccd1 vccd1 _1676_/X sky130_fd_sc_hd__and4_4
XFILLER_7_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2159_ _2157_/Y _1656_/X _2158_/X _2112_/X _1594_/C vssd1 vssd1 vccd1 vccd1 _2159_/X
+ sky130_fd_sc_hd__a2111o_4
X_2228_ _2225_/Y _1560_/X _2227_/Y vssd1 vssd1 vccd1 vccd1 _2228_/Y sky130_fd_sc_hd__a21boi_4
XFILLER_42_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_3_0_0_addressalyzerBlock.SPI_CLK clkbuf_3_1_0_addressalyzerBlock.SPI_CLK/A
+ vssd1 vssd1 vccd1 vccd1 clkbuf_3_0_0_addressalyzerBlock.SPI_CLK/X sky130_fd_sc_hd__clkbuf_1
XFILLER_13_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1530_ _1499_/C vssd1 vssd1 vccd1 vccd1 _1530_/X sky130_fd_sc_hd__buf_2
X_1392_ _1392_/A _1392_/B vssd1 vssd1 vccd1 vccd1 _1392_/Y sky130_fd_sc_hd__nand2_4
X_1461_ _1444_/C vssd1 vssd1 vccd1 vccd1 _1486_/B sky130_fd_sc_hd__buf_2
X_2013_ _2532_/Q _2012_/X _1979_/A _2534_/Q _2000_/A vssd1 vssd1 vccd1 vccd1 _2014_/C
+ sky130_fd_sc_hd__a41oi_4
XFILLER_50_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1728_ _1485_/Y _1725_/Y _1618_/Y _1726_/Y _1727_/Y vssd1 vssd1 vccd1 vccd1 _2651_/D
+ sky130_fd_sc_hd__a41oi_4
XFILLER_12_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1659_ _1500_/X _2187_/B _1367_/A _1592_/X vssd1 vssd1 vccd1 vccd1 _1659_/Y sky130_fd_sc_hd__a2bb2oi_4
XFILLER_37_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2700_ _2695_/CLK _1284_/Y vssd1 vssd1 vccd1 vccd1 _2700_/Q sky130_fd_sc_hd__dfxtp_4
X_2631_ _2511_/CLK _2631_/D vssd1 vssd1 vccd1 vccd1 _2631_/Q sky130_fd_sc_hd__dfxtp_4
X_2562_ _2561_/CLK _1937_/X vssd1 vssd1 vccd1 vccd1 DATA_TO_HASH[5] sky130_fd_sc_hd__dfxtp_4
X_1375_ _1375_/A vssd1 vssd1 vccd1 vccd1 _1375_/Y sky130_fd_sc_hd__inv_2
X_1444_ _1444_/A _1444_/B _1444_/C vssd1 vssd1 vccd1 vccd1 _1450_/B sky130_fd_sc_hd__nor3_4
X_1513_ _1485_/Y _1509_/Y _1512_/X vssd1 vssd1 vccd1 vccd1 _1513_/X sky130_fd_sc_hd__a21o_4
X_2493_ _2493_/CLK _2493_/D vssd1 vssd1 vccd1 vccd1 _2493_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_63_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1993_ _1979_/Y _2003_/A vssd1 vssd1 vccd1 vccd1 _1993_/Y sky130_fd_sc_hd__nor2_4
X_2545_ _2545_/CLK _1963_/X vssd1 vssd1 vccd1 vccd1 MACRO_WR_SELECT[0] sky130_fd_sc_hd__dfxtp_4
X_2614_ _2621_/CLK _2614_/D vssd1 vssd1 vccd1 vccd1 _2614_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_9_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1358_ _1355_/B _1355_/A _1355_/C _1338_/X _1293_/X vssd1 vssd1 vccd1 vccd1 _1358_/Y
+ sky130_fd_sc_hd__a41oi_4
X_1427_ _1432_/A _2671_/Q _1414_/B _1432_/C _2672_/Q vssd1 vssd1 vccd1 vccd1 _1428_/C
+ sky130_fd_sc_hd__a41oi_4
X_2476_ _2478_/CLK _2476_/D vssd1 vssd1 vccd1 vccd1 _2476_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_18_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1289_ _1286_/X _2005_/B _1288_/Y vssd1 vssd1 vccd1 vccd1 _1289_/X sky130_fd_sc_hd__and3_4
XPHY_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2261_ _2259_/Y _2260_/Y _2162_/A vssd1 vssd1 vccd1 vccd1 _2261_/Y sky130_fd_sc_hd__a21oi_4
X_2192_ _2241_/A _2241_/B _2600_/Q _2241_/D vssd1 vssd1 vccd1 vccd1 _2192_/X sky130_fd_sc_hd__and4_4
X_1212_ _1222_/A vssd1 vssd1 vccd1 vccd1 _1212_/X sky130_fd_sc_hd__buf_2
XFILLER_1_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2330_ _1516_/X _2137_/Y _2319_/Y _1910_/B _2321_/X vssd1 vssd1 vccd1 vccd1 _2455_/D
+ sky130_fd_sc_hd__o32ai_4
XFILLER_52_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1976_ _1283_/B _1976_/B vssd1 vssd1 vccd1 vccd1 _1976_/X sky130_fd_sc_hd__and2_4
X_2528_ _2564_/CLK _2041_/Y vssd1 vssd1 vccd1 vccd1 _2528_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_29_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2459_ _2493_/CLK _2326_/Y vssd1 vssd1 vccd1 vccd1 _1900_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_61_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_4_0_0_m1_clk_local clkbuf_4_1_0_m1_clk_local/A vssd1 vssd1 vccd1 vccd1 _2582_/CLK
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_59_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1761_ _1761_/A vssd1 vssd1 vccd1 vccd1 _1761_/Y sky130_fd_sc_hd__inv_2
X_1830_ _1829_/Y vssd1 vssd1 vccd1 vccd1 _1830_/Y sky130_fd_sc_hd__inv_2
X_2313_ _1928_/B _2306_/X _1726_/A _2308_/X vssd1 vssd1 vccd1 vccd1 _2466_/D sky130_fd_sc_hd__a2bb2o_4
X_1692_ _1683_/B _1707_/A _1692_/C _1707_/D vssd1 vssd1 vccd1 vccd1 _1692_/X sky130_fd_sc_hd__and4_4
XFILLER_53_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2244_ _2170_/X _1751_/A _1562_/X vssd1 vssd1 vccd1 vccd1 _2244_/Y sky130_fd_sc_hd__a21oi_4
X_2175_ _1926_/B _2170_/X _2174_/Y vssd1 vssd1 vccd1 vccd1 _2175_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_31_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1959_ _1961_/A _2555_/Q vssd1 vssd1 vccd1 vccd1 _2549_/D sky130_fd_sc_hd__and2_4
XFILLER_48_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_3_6_0_m1_clk_local clkbuf_3_7_0_m1_clk_local/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_6_0_m1_clk_local/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_47_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1744_ _1707_/C _1683_/B _1743_/Y vssd1 vssd1 vccd1 vccd1 _1744_/X sky130_fd_sc_hd__o21a_4
XFILLER_7_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1813_ _2630_/Q _2507_/Q _1804_/X vssd1 vssd1 vccd1 vccd1 _1813_/X sky130_fd_sc_hd__o21a_4
X_1675_ _1675_/A vssd1 vssd1 vccd1 vccd1 _1683_/A sky130_fd_sc_hd__inv_2
X_2089_ _2089_/A vssd1 vssd1 vccd1 vccd1 _2104_/B sky130_fd_sc_hd__inv_2
X_2158_ _1542_/D vssd1 vssd1 vccd1 vccd1 _2158_/X sky130_fd_sc_hd__buf_2
X_2227_ _1952_/B _2170_/X _2226_/Y vssd1 vssd1 vccd1 vccd1 _2227_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_41_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1391_ _1394_/A _1257_/A _2679_/Q vssd1 vssd1 vccd1 vccd1 _1392_/B sky130_fd_sc_hd__nand3_4
X_1460_ _1460_/A vssd1 vssd1 vccd1 vccd1 _1460_/Y sky130_fd_sc_hd__inv_2
X_2012_ _2012_/A _2026_/A _2531_/Q _2012_/D vssd1 vssd1 vccd1 vccd1 _2012_/X sky130_fd_sc_hd__and4_4
XFILLER_50_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1658_ _1658_/A _1657_/X vssd1 vssd1 vccd1 vccd1 _1658_/Y sky130_fd_sc_hd__nand2_4
X_1727_ _1712_/X _1695_/X _1697_/X vssd1 vssd1 vccd1 vccd1 _1727_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_58_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1589_ _1594_/C vssd1 vssd1 vccd1 vccd1 _2187_/B sky130_fd_sc_hd__buf_2
XFILLER_41_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1512_ _1511_/X vssd1 vssd1 vccd1 vccd1 _1512_/X sky130_fd_sc_hd__buf_2
X_2561_ _2561_/CLK _1939_/X vssd1 vssd1 vccd1 vccd1 DATA_TO_HASH[4] sky130_fd_sc_hd__dfxtp_4
X_2492_ _2456_/CLK _2492_/D vssd1 vssd1 vccd1 vccd1 _2118_/C sky130_fd_sc_hd__dfxtp_4
X_2630_ _2511_/CLK _2630_/D vssd1 vssd1 vccd1 vccd1 _2630_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_55_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1374_ _1372_/Y _1330_/B _1373_/Y vssd1 vssd1 vccd1 vccd1 _1375_/A sky130_fd_sc_hd__nand3_4
X_1443_ _1637_/C _1496_/A _1497_/A _1571_/B vssd1 vssd1 vccd1 vccd1 _1444_/C sky130_fd_sc_hd__nand4_4
XFILLER_4_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1992_ _2531_/Q _1992_/B _2532_/Q _2012_/D vssd1 vssd1 vccd1 vccd1 _2003_/A sky130_fd_sc_hd__nand4_4
XFILLER_20_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2613_ _2621_/CLK _2613_/D vssd1 vssd1 vccd1 vccd1 _2613_/Q sky130_fd_sc_hd__dfxtp_4
X_2544_ _2514_/CLK _2544_/D vssd1 vssd1 vccd1 vccd1 _1618_/A sky130_fd_sc_hd__dfxtp_4
X_2475_ _2494_/CLK _2299_/Y vssd1 vssd1 vccd1 vccd1 _2475_/Q sky130_fd_sc_hd__dfxtp_4
X_1288_ _1282_/C _1305_/A _1268_/X _1282_/D vssd1 vssd1 vccd1 vccd1 _1288_/Y sky130_fd_sc_hd__nand4_4
X_1357_ _1345_/X _1355_/X _1356_/Y vssd1 vssd1 vccd1 vccd1 _1357_/X sky130_fd_sc_hd__o21a_4
X_1426_ _1414_/C vssd1 vssd1 vccd1 vccd1 _1432_/C sky130_fd_sc_hd__buf_2
XFILLER_28_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2260_ _2260_/A THREAD_COUNT[1] vssd1 vssd1 vccd1 vccd1 _2260_/Y sky130_fd_sc_hd__nand2_4
X_2191_ _2188_/X _2189_/X _2190_/Y vssd1 vssd1 vccd1 vccd1 _2191_/Y sky130_fd_sc_hd__a21oi_4
X_1211_ _2353_/B vssd1 vssd1 vccd1 vccd1 _1222_/A sky130_fd_sc_hd__buf_2
XFILLER_1_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1975_ _1975_/A vssd1 vssd1 vccd1 vccd1 _2540_/D sky130_fd_sc_hd__inv_2
X_2527_ _2527_/CLK _2045_/Y vssd1 vssd1 vccd1 vccd1 _1981_/A sky130_fd_sc_hd__dfxtp_4
X_1409_ _1401_/X _1396_/X _2058_/A vssd1 vssd1 vccd1 vccd1 _1409_/Y sky130_fd_sc_hd__a21oi_4
X_2458_ _2478_/CLK _2327_/Y vssd1 vssd1 vccd1 vccd1 _2195_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_43_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2389_ S1_CLK_IN vssd1 vssd1 vccd1 vccd1 _2389_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_4_0_0_addressalyzerBlock.SPI_CLK clkbuf_3_0_0_addressalyzerBlock.SPI_CLK/X
+ vssd1 vssd1 vccd1 vccd1 _2478_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_51_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1760_ _2443_/Q vssd1 vssd1 vccd1 vccd1 _2177_/B sky130_fd_sc_hd__inv_2
X_1691_ _1687_/Y _1690_/Y _1492_/X vssd1 vssd1 vccd1 vccd1 _1691_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_32_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2312_ _1926_/B _2306_/X _1784_/X _2308_/X vssd1 vssd1 vccd1 vccd1 _2467_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_65_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2243_ _1953_/A _2147_/B vssd1 vssd1 vccd1 vccd1 _2243_/Y sky130_fd_sc_hd__nand2_4
X_2174_ _2222_/A _2475_/Q _2494_/Q vssd1 vssd1 vccd1 vccd1 _2174_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_21_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1889_ _1378_/A vssd1 vssd1 vccd1 vccd1 _1915_/A sky130_fd_sc_hd__buf_2
X_1958_ _1961_/A _1958_/B vssd1 vssd1 vccd1 vccd1 _1958_/X sky130_fd_sc_hd__and2_4
Xclkbuf_3_5_0_addressalyzerBlock.SPI_CLK clkbuf_3_5_0_addressalyzerBlock.SPI_CLK/A
+ vssd1 vssd1 vccd1 vccd1 clkbuf_3_5_0_addressalyzerBlock.SPI_CLK/X sky130_fd_sc_hd__clkbuf_1
XFILLER_56_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1743_ _1464_/X _1450_/B _1460_/A _1707_/C _1488_/X vssd1 vssd1 vccd1 vccd1 _1743_/Y
+ sky130_fd_sc_hd__a41oi_4
X_1812_ _2630_/Q _1798_/A _1811_/X vssd1 vssd1 vccd1 vccd1 _2631_/D sky130_fd_sc_hd__o21a_4
XFILLER_7_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1674_ _1673_/Y vssd1 vssd1 vccd1 vccd1 _1674_/X sky130_fd_sc_hd__buf_2
X_2226_ _2194_/X _1761_/A _1559_/X vssd1 vssd1 vccd1 vccd1 _2226_/Y sky130_fd_sc_hd__a21oi_4
X_2088_ _1873_/A _2397_/A vssd1 vssd1 vccd1 vccd1 _2088_/X sky130_fd_sc_hd__and2_4
X_2157_ _2674_/Q vssd1 vssd1 vccd1 vccd1 _2157_/Y sky130_fd_sc_hd__inv_2
XFILLER_26_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1390_ _1257_/A _1389_/X _1378_/X vssd1 vssd1 vccd1 vccd1 _1392_/A sky130_fd_sc_hd__o21a_4
XFILLER_4_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2011_ _2528_/Q vssd1 vssd1 vccd1 vccd1 _2026_/A sky130_fd_sc_hd__buf_2
XFILLER_35_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1657_ _1321_/Y _1656_/X _1582_/X _1583_/X vssd1 vssd1 vccd1 vccd1 _1657_/X sky130_fd_sc_hd__a211o_4
X_1588_ _1587_/X vssd1 vssd1 vccd1 vccd1 _1594_/C sky130_fd_sc_hd__buf_2
X_1726_ _1726_/A _2378_/B vssd1 vssd1 vccd1 vccd1 _1726_/Y sky130_fd_sc_hd__nand2_4
X_2209_ _2206_/Y _2207_/Y _2208_/Y vssd1 vssd1 vccd1 vccd1 _2209_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_53_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1511_ _1542_/D vssd1 vssd1 vccd1 vccd1 _1511_/X sky130_fd_sc_hd__buf_2
X_1442_ _1442_/A vssd1 vssd1 vccd1 vccd1 _1571_/B sky130_fd_sc_hd__buf_2
X_2560_ _2561_/CLK _2560_/D vssd1 vssd1 vccd1 vccd1 DATA_TO_HASH[3] sky130_fd_sc_hd__dfxtp_4
X_2491_ _2443_/CLK _2491_/D vssd1 vssd1 vccd1 vccd1 _1649_/A sky130_fd_sc_hd__dfxtp_4
X_1373_ _1277_/A _1377_/B _1367_/A vssd1 vssd1 vccd1 vccd1 _1373_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_4_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2689_ _2559_/CLK _1344_/Y vssd1 vssd1 vccd1 vccd1 _1264_/B sky130_fd_sc_hd__dfxtp_4
X_1709_ _1702_/Y _1705_/Y _1708_/Y vssd1 vssd1 vccd1 vccd1 _1709_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_54_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2612_ _2612_/CLK _2612_/D vssd1 vssd1 vccd1 vccd1 _2612_/Q sky130_fd_sc_hd__dfxtp_4
X_1991_ _1990_/Y vssd1 vssd1 vccd1 vccd1 _2012_/D sky130_fd_sc_hd__inv_2
XFILLER_9_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1425_ _1414_/A vssd1 vssd1 vccd1 vccd1 _1432_/A sky130_fd_sc_hd__buf_2
X_2543_ _2413_/CLK _2543_/D vssd1 vssd1 vccd1 vccd1 _1966_/A sky130_fd_sc_hd__dfxtp_4
X_2474_ _2494_/CLK _2301_/Y vssd1 vssd1 vccd1 vccd1 _2198_/B sky130_fd_sc_hd__dfxtp_4
X_1356_ _1345_/X _1280_/A _1355_/B _1355_/C _1293_/X vssd1 vssd1 vccd1 vccd1 _1356_/Y
+ sky130_fd_sc_hd__a41oi_4
XFILLER_55_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1287_ _1274_/X vssd1 vssd1 vccd1 vccd1 _2005_/B sky130_fd_sc_hd__buf_2
XPHY_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2190_ _2190_/A _2190_/B vssd1 vssd1 vccd1 vccd1 _2190_/Y sky130_fd_sc_hd__nor2_4
X_1210_ _2331_/A vssd1 vssd1 vccd1 vccd1 _2353_/B sky130_fd_sc_hd__inv_2
XFILLER_1_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1974_ _1974_/A _1833_/Y _1974_/C vssd1 vssd1 vccd1 vccd1 _1975_/A sky130_fd_sc_hd__or3_4
X_2526_ _2527_/CLK _2047_/Y vssd1 vssd1 vccd1 vccd1 _1980_/A sky130_fd_sc_hd__dfxtp_4
X_1408_ _1293_/A vssd1 vssd1 vccd1 vccd1 _2058_/A sky130_fd_sc_hd__buf_2
X_2457_ _2494_/CLK _2457_/D vssd1 vssd1 vccd1 vccd1 _1904_/A sky130_fd_sc_hd__dfxtp_4
X_2388_ PLL_INPUT M1_CLK_SELECT _2387_/Y vssd1 vssd1 vccd1 vccd1 m1_clk_local sky130_fd_sc_hd__o21a_4
X_1339_ _1266_/A _1338_/X _1280_/B vssd1 vssd1 vccd1 vccd1 _1339_/Y sky130_fd_sc_hd__nand3_4
XFILLER_43_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1690_ _1688_/Y _1689_/Y _1675_/A vssd1 vssd1 vccd1 vccd1 _1690_/Y sky130_fd_sc_hd__o21ai_4
X_2242_ _1500_/A _2154_/X _1255_/A _1591_/Y vssd1 vssd1 vccd1 vccd1 _2242_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_25_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2311_ _1923_/B _2306_/X _1481_/X _2308_/X vssd1 vssd1 vccd1 vccd1 _2311_/X sky130_fd_sc_hd__a2bb2o_4
X_2173_ _2248_/A vssd1 vssd1 vccd1 vccd1 _2222_/A sky130_fd_sc_hd__buf_2
XFILLER_33_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1957_ _1915_/A vssd1 vssd1 vccd1 vccd1 _1961_/A sky130_fd_sc_hd__buf_2
X_2509_ _2508_/CLK _2509_/D vssd1 vssd1 vccd1 vccd1 _1828_/A sky130_fd_sc_hd__dfxtp_4
X_1888_ _1901_/A _1888_/B vssd1 vssd1 vccd1 vccd1 _2591_/D sky130_fd_sc_hd__nor2_4
XFILLER_56_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1811_ _2631_/Q _2507_/Q _1804_/X vssd1 vssd1 vccd1 vccd1 _1811_/X sky130_fd_sc_hd__o21a_4
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1673_ _2434_/Q vssd1 vssd1 vccd1 vccd1 _1673_/Y sky130_fd_sc_hd__inv_2
X_1742_ _1532_/Y _1674_/X _1695_/X vssd1 vssd1 vccd1 vccd1 _1742_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_38_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2225_ _2225_/A _2225_/B vssd1 vssd1 vccd1 vccd1 _2225_/Y sky130_fd_sc_hd__nand2_4
X_2156_ _2156_/A _2155_/X vssd1 vssd1 vccd1 vccd1 _2156_/Y sky130_fd_sc_hd__nand2_4
XFILLER_26_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2087_ _1873_/A IRQ_OUT_fromClient vssd1 vssd1 vccd1 vccd1 _2087_/X sky130_fd_sc_hd__and2_4
XFILLER_21_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2010_ _2009_/X _1981_/Y _1989_/D vssd1 vssd1 vccd1 vccd1 _2012_/A sky130_fd_sc_hd__nor3_4
XFILLER_50_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_3_2_0_m1_clk_local clkbuf_3_3_0_m1_clk_local/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_5_0_m1_clk_local/A
+ sky130_fd_sc_hd__clkbuf_1
X_1725_ _1712_/X _1724_/X _1720_/Y vssd1 vssd1 vccd1 vccd1 _1725_/Y sky130_fd_sc_hd__o21ai_4
X_1587_ _1587_/A vssd1 vssd1 vccd1 vccd1 _1587_/X sky130_fd_sc_hd__buf_2
X_1656_ _1499_/C vssd1 vssd1 vccd1 vccd1 _1656_/X sky130_fd_sc_hd__buf_2
X_2208_ _1263_/A _1530_/X _1515_/X _1581_/X _2139_/X vssd1 vssd1 vccd1 vccd1 _2208_/Y
+ sky130_fd_sc_hd__a2111oi_4
X_2139_ _1573_/A vssd1 vssd1 vccd1 vccd1 _2139_/X sky130_fd_sc_hd__buf_2
XFILLER_41_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1510_ _1510_/A vssd1 vssd1 vccd1 vccd1 _1542_/D sky130_fd_sc_hd__inv_2
X_1441_ _1541_/B vssd1 vssd1 vccd1 vccd1 _1444_/B sky130_fd_sc_hd__inv_2
X_2490_ _2493_/CLK _2128_/Y vssd1 vssd1 vccd1 vccd1 _2490_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_4_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1372_ _1367_/Y vssd1 vssd1 vccd1 vccd1 _1372_/Y sky130_fd_sc_hd__inv_2
XFILLER_23_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2688_ _2693_/CLK _2688_/D vssd1 vssd1 vccd1 vccd1 _1263_/A sky130_fd_sc_hd__dfxtp_4
X_1708_ _1708_/A _1450_/D vssd1 vssd1 vccd1 vccd1 _1708_/Y sky130_fd_sc_hd__nand2_4
X_1639_ _2143_/A _1638_/Y vssd1 vssd1 vccd1 vccd1 _1639_/Y sky130_fd_sc_hd__nor2_4
XFILLER_64_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1990_ _1990_/A _1990_/B vssd1 vssd1 vccd1 vccd1 _1990_/Y sky130_fd_sc_hd__nand2_4
X_2611_ _2621_/CLK _2611_/D vssd1 vssd1 vccd1 vccd1 _2611_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_55_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2542_ _2413_/CLK _1971_/X vssd1 vssd1 vccd1 vccd1 _2542_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_9_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1355_ _1355_/A _1355_/B _1355_/C _1338_/X vssd1 vssd1 vccd1 vccd1 _1355_/X sky130_fd_sc_hd__and4_4
X_1424_ _1424_/A vssd1 vssd1 vccd1 vccd1 _1424_/Y sky130_fd_sc_hd__inv_2
X_2473_ _2494_/CLK _2473_/D vssd1 vssd1 vccd1 vccd1 _1882_/A sky130_fd_sc_hd__dfxtp_4
X_1286_ _1285_/Y _2696_/Q _2695_/Q _1282_/D _1282_/C vssd1 vssd1 vccd1 vccd1 _1286_/X
+ sky130_fd_sc_hd__a41o_4
XPHY_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_4_5_0_addressalyzerBlock.SPI_CLK clkbuf_4_5_0_addressalyzerBlock.SPI_CLK/A
+ vssd1 vssd1 vccd1 vccd1 _2511_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_65_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1973_ _1969_/Y _1966_/B _1973_/C vssd1 vssd1 vccd1 vccd1 _1973_/X sky130_fd_sc_hd__and3_4
X_2525_ _2527_/CLK _2525_/D vssd1 vssd1 vccd1 vccd1 _1988_/D sky130_fd_sc_hd__dfxtp_4
X_1338_ _1266_/B vssd1 vssd1 vccd1 vccd1 _1338_/X sky130_fd_sc_hd__buf_2
X_1407_ _2014_/A _1407_/B _1407_/C vssd1 vssd1 vccd1 vccd1 _1407_/Y sky130_fd_sc_hd__nor3_4
X_2387_ _2387_/A M1_CLK_SELECT vssd1 vssd1 vccd1 vccd1 _2387_/Y sky130_fd_sc_hd__nand2_4
X_2456_ _2456_/CLK _2456_/D vssd1 vssd1 vccd1 vccd1 _2245_/B sky130_fd_sc_hd__dfxtp_4
X_1269_ _2697_/Q vssd1 vssd1 vccd1 vccd1 _1300_/B sky130_fd_sc_hd__buf_2
XPHY_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2241_ _2241_/A _2241_/B _2598_/Q _2241_/D vssd1 vssd1 vccd1 vccd1 _2241_/X sky130_fd_sc_hd__and4_4
XFILLER_38_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2310_ _1921_/B _2306_/X _1694_/A _2308_/X vssd1 vssd1 vccd1 vccd1 _2469_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_18_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2172_ _2169_/Y _1647_/X _2171_/Y vssd1 vssd1 vccd1 vccd1 _2172_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_65_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1956_ _1956_/A _1956_/B vssd1 vssd1 vccd1 vccd1 _2551_/D sky130_fd_sc_hd__nor2_4
XFILLER_33_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1887_ _1887_/A vssd1 vssd1 vccd1 vccd1 _1888_/B sky130_fd_sc_hd__inv_2
X_2508_ _2508_/CLK _2508_/D vssd1 vssd1 vccd1 vccd1 _2382_/C sky130_fd_sc_hd__dfxtp_4
XFILLER_56_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2439_ _2495_/CLK _2364_/X vssd1 vssd1 vccd1 vccd1 _1754_/B sky130_fd_sc_hd__dfxtp_4
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1810_ _2631_/Q _1798_/X _1809_/X vssd1 vssd1 vccd1 vccd1 _2632_/D sky130_fd_sc_hd__o21a_4
X_1741_ _1736_/Y _1739_/Y _1740_/X vssd1 vssd1 vccd1 vccd1 _1741_/X sky130_fd_sc_hd__o21a_4
X_1672_ _1452_/A vssd1 vssd1 vccd1 vccd1 _1672_/Y sky130_fd_sc_hd__inv_2
X_2155_ _1249_/A _1591_/A _1583_/X _1500_/A _2154_/X vssd1 vssd1 vccd1 vccd1 _2155_/X
+ sky130_fd_sc_hd__o32a_4
XFILLER_38_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2224_ _2224_/A _1548_/X _2223_/Y vssd1 vssd1 vccd1 vccd1 _2225_/B sky130_fd_sc_hd__nand3_4
XFILLER_61_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2086_ _1873_/A _2511_/Q vssd1 vssd1 vccd1 vccd1 _2086_/X sky130_fd_sc_hd__and2_4
XFILLER_21_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1939_ _1941_/A _2569_/Q vssd1 vssd1 vccd1 vccd1 _1939_/X sky130_fd_sc_hd__and2_4
XFILLER_16_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0_addressalyzerBlock.SPI_CLK clkbuf_0_addressalyzerBlock.SPI_CLK/X vssd1
+ vssd1 vccd1 vccd1 clkbuf_2_2_0_addressalyzerBlock.SPI_CLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_4_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1724_ _1676_/X _1717_/C _1717_/D _1707_/C vssd1 vssd1 vccd1 vccd1 _1724_/X sky130_fd_sc_hd__and4_4
X_1655_ _1582_/X _1535_/X _1583_/X _1637_/X _1654_/Y vssd1 vssd1 vccd1 vccd1 _1658_/A
+ sky130_fd_sc_hd__o32ai_4
X_1586_ _1635_/A _1635_/B _2163_/B vssd1 vssd1 vccd1 vccd1 _1587_/A sky130_fd_sc_hd__nand3_4
X_2207_ _1574_/X _2696_/Q _1544_/X vssd1 vssd1 vccd1 vccd1 _2207_/Y sky130_fd_sc_hd__a21oi_4
X_2069_ _2520_/Q _2067_/Y _2068_/Y vssd1 vssd1 vccd1 vccd1 _2069_/X sky130_fd_sc_hd__a21o_4
X_2138_ _1626_/Y _1598_/Y _2137_/Y _1956_/B _2126_/Y vssd1 vssd1 vccd1 vccd1 _2485_/D
+ sky130_fd_sc_hd__o32ai_4
XFILLER_41_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1371_ _1371_/A vssd1 vssd1 vccd1 vccd1 _1371_/Y sky130_fd_sc_hd__inv_2
X_1440_ _1676_/D vssd1 vssd1 vccd1 vccd1 _1444_/A sky130_fd_sc_hd__inv_2
XFILLER_4_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2687_ _2693_/CLK _1357_/X vssd1 vssd1 vccd1 vccd1 _2687_/Q sky130_fd_sc_hd__dfxtp_4
X_1638_ _1638_/A vssd1 vssd1 vccd1 vccd1 _1638_/Y sky130_fd_sc_hd__inv_2
X_1707_ _1707_/A _1683_/B _1707_/C _1707_/D vssd1 vssd1 vccd1 vccd1 _1708_/A sky130_fd_sc_hd__nand4_4
X_1569_ _1464_/X _1567_/Y _1568_/X vssd1 vssd1 vccd1 vccd1 _1569_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_39_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2610_ _2621_/CLK _1857_/X vssd1 vssd1 vccd1 vccd1 _2610_/Q sky130_fd_sc_hd__dfxtp_4
X_2472_ _2494_/CLK _2303_/Y vssd1 vssd1 vccd1 vccd1 _2472_/Q sky130_fd_sc_hd__dfxtp_4
X_2541_ _2413_/CLK _1973_/X vssd1 vssd1 vccd1 vccd1 _2541_/Q sky130_fd_sc_hd__dfxtp_4
X_1285_ _1281_/C _1281_/D vssd1 vssd1 vccd1 vccd1 _1285_/Y sky130_fd_sc_hd__nor2_4
X_1354_ _1353_/Y vssd1 vssd1 vccd1 vccd1 _2688_/D sky130_fd_sc_hd__inv_2
XFILLER_48_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1423_ _1419_/C _1419_/A _1422_/Y vssd1 vssd1 vccd1 vccd1 _1424_/A sky130_fd_sc_hd__o21ai_4
XFILLER_55_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_4_10_0_addressalyzerBlock.SPI_CLK clkbuf_3_5_0_addressalyzerBlock.SPI_CLK/X
+ vssd1 vssd1 vccd1 vccd1 _2621_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_42_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1972_ _1974_/A _2541_/Q vssd1 vssd1 vccd1 vccd1 _1973_/C sky130_fd_sc_hd__or2_4
X_2524_ _2527_/CLK _2524_/D vssd1 vssd1 vccd1 vccd1 _1988_/C sky130_fd_sc_hd__dfxtp_4
X_2455_ _2456_/CLK _2455_/D vssd1 vssd1 vccd1 vccd1 _1909_/A sky130_fd_sc_hd__dfxtp_4
X_1268_ _2696_/Q vssd1 vssd1 vccd1 vccd1 _1268_/X sky130_fd_sc_hd__buf_2
X_1337_ _1337_/A vssd1 vssd1 vccd1 vccd1 _1337_/Y sky130_fd_sc_hd__inv_2
X_1406_ _1401_/X _1396_/X _1255_/B vssd1 vssd1 vccd1 vccd1 _1407_/C sky130_fd_sc_hd__a21oi_4
XFILLER_29_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2386_ M1_CLK_IN vssd1 vssd1 vccd1 vccd1 _2387_/A sky130_fd_sc_hd__inv_2
XFILLER_51_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2240_ _2238_/Y _2239_/Y vssd1 vssd1 vccd1 vccd1 _2481_/D sky130_fd_sc_hd__nand2_4
X_2171_ _2170_/X _1900_/A _2250_/B vssd1 vssd1 vccd1 vccd1 _2171_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_25_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1955_ _2485_/Q vssd1 vssd1 vccd1 vccd1 _1956_/B sky130_fd_sc_hd__inv_2
X_1886_ _1875_/A vssd1 vssd1 vccd1 vccd1 _1901_/A sky130_fd_sc_hd__buf_2
X_2438_ _2438_/CLK _2438_/D vssd1 vssd1 vccd1 vccd1 _1664_/C sky130_fd_sc_hd__dfxtp_4
X_2507_ _2511_/CLK _2507_/D vssd1 vssd1 vccd1 vccd1 _2507_/Q sky130_fd_sc_hd__dfxtp_4
X_2369_ _1609_/Y _2369_/B _1613_/A vssd1 vssd1 vccd1 vccd1 _2369_/Y sky130_fd_sc_hd__nand3_4
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1671_ _1670_/Y vssd1 vssd1 vccd1 vccd1 _1671_/Y sky130_fd_sc_hd__inv_2
XFILLER_11_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1740_ _1717_/D _1685_/Y _1697_/X vssd1 vssd1 vccd1 vccd1 _1740_/X sky130_fd_sc_hd__o21a_4
XFILLER_53_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2154_ _1587_/A vssd1 vssd1 vccd1 vccd1 _2154_/X sky130_fd_sc_hd__buf_2
XFILLER_38_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2085_ _1873_/A _2503_/Q vssd1 vssd1 vccd1 vccd1 _2085_/X sky130_fd_sc_hd__and2_4
X_2223_ _2223_/A _1546_/A vssd1 vssd1 vccd1 vccd1 _2223_/Y sky130_fd_sc_hd__nand2_4
XFILLER_21_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1869_ _1871_/A _1869_/B vssd1 vssd1 vccd1 vccd1 _1869_/X sky130_fd_sc_hd__and2_4
X_1938_ _1915_/A vssd1 vssd1 vccd1 vccd1 _1941_/A sky130_fd_sc_hd__buf_2
XFILLER_29_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1654_ _1651_/Y _1653_/Y _1574_/X vssd1 vssd1 vccd1 vccd1 _1654_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_7_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1723_ _1719_/Y _1721_/Y _1722_/X vssd1 vssd1 vccd1 vccd1 _1723_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_58_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2206_ _1653_/A _2204_/Y _2205_/X vssd1 vssd1 vccd1 vccd1 _2206_/Y sky130_fd_sc_hd__o21ai_4
X_1585_ _1544_/X _1580_/Y _1584_/X vssd1 vssd1 vccd1 vccd1 _1585_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_66_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2068_ _2520_/Q _2067_/Y _1378_/X vssd1 vssd1 vccd1 vccd1 _2068_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_26_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2137_ _1829_/B _2115_/X _2137_/C vssd1 vssd1 vccd1 vccd1 _2137_/Y sky130_fd_sc_hd__nand3_4
XFILLER_1_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1370_ _1368_/X _1370_/B vssd1 vssd1 vccd1 vccd1 _1371_/A sky130_fd_sc_hd__nand2_4
XFILLER_4_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2686_ _2693_/CLK _2686_/D vssd1 vssd1 vccd1 vccd1 _1263_/C sky130_fd_sc_hd__dfxtp_4
X_1637_ _2241_/A _1282_/C _1637_/C _2241_/D vssd1 vssd1 vccd1 vccd1 _1637_/X sky130_fd_sc_hd__and4_4
X_1706_ _1692_/C vssd1 vssd1 vccd1 vccd1 _1707_/C sky130_fd_sc_hd__buf_2
X_1568_ _1568_/A _1439_/X vssd1 vssd1 vccd1 vccd1 _1568_/X sky130_fd_sc_hd__or2_4
X_1499_ _1510_/A _1581_/A _1499_/C vssd1 vssd1 vccd1 vccd1 _1500_/A sky130_fd_sc_hd__nand3_4
XFILLER_54_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1422_ _1419_/A _1419_/C _1298_/X vssd1 vssd1 vccd1 vccd1 _1422_/Y sky130_fd_sc_hd__a21oi_4
X_2540_ _2413_/CLK _2540_/D vssd1 vssd1 vccd1 vccd1 _1974_/A sky130_fd_sc_hd__dfxtp_4
X_2471_ _2494_/CLK _2471_/D vssd1 vssd1 vccd1 vccd1 _1887_/A sky130_fd_sc_hd__dfxtp_4
X_1284_ _1284_/A vssd1 vssd1 vccd1 vccd1 _1284_/Y sky130_fd_sc_hd__inv_2
XFILLER_55_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1353_ _1348_/X _1353_/B vssd1 vssd1 vccd1 vccd1 _1353_/Y sky130_fd_sc_hd__nand2_4
XFILLER_36_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2669_ _2670_/CLK _1436_/X vssd1 vssd1 vccd1 vccd1 _1414_/C sky130_fd_sc_hd__dfxtp_4
XFILLER_46_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1971_ _1969_/Y _1971_/B _1971_/C vssd1 vssd1 vccd1 vccd1 _1971_/X sky130_fd_sc_hd__and3_4
X_2523_ _2527_/CLK _2060_/X vssd1 vssd1 vccd1 vccd1 _1988_/A sky130_fd_sc_hd__dfxtp_4
X_1405_ _1298_/X vssd1 vssd1 vccd1 vccd1 _2014_/A sky130_fd_sc_hd__buf_2
X_2385_ EXT_RESET_N_fromHost vssd1 vssd1 vccd1 vccd1 _2385_/Y sky130_fd_sc_hd__inv_2
X_2454_ _2478_/CLK _2454_/D vssd1 vssd1 vccd1 vccd1 _2335_/C sky130_fd_sc_hd__dfxtp_4
X_1267_ _1246_/Y _1247_/Y _1281_/C _1313_/A vssd1 vssd1 vccd1 vccd1 _1305_/A sky130_fd_sc_hd__nor4_4
X_1336_ _1336_/A _1335_/Y vssd1 vssd1 vccd1 vccd1 _1337_/A sky130_fd_sc_hd__nand2_4
XFILLER_36_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_0_addressalyzerBlock.SPI_CLK _2391_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0_addressalyzerBlock.SPI_CLK/X
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_19_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2170_ _2248_/A vssd1 vssd1 vccd1 vccd1 _2170_/X sky130_fd_sc_hd__buf_2
X_1954_ _1946_/A _1954_/B vssd1 vssd1 vccd1 vccd1 _1954_/Y sky130_fd_sc_hd__nor2_4
XFILLER_18_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1885_ _1875_/X _1884_/Y vssd1 vssd1 vccd1 vccd1 _1885_/Y sky130_fd_sc_hd__nor2_4
Xclkbuf_2_1_0_addressalyzerBlock.SPI_CLK clkbuf_1_0_0_addressalyzerBlock.SPI_CLK/X
+ vssd1 vssd1 vccd1 vccd1 clkbuf_3_3_0_addressalyzerBlock.SPI_CLK/A sky130_fd_sc_hd__clkbuf_1
X_2368_ _2367_/X _1623_/Y _1840_/A vssd1 vssd1 vccd1 vccd1 _2438_/D sky130_fd_sc_hd__o21a_4
X_2437_ _2438_/CLK _2384_/Y vssd1 vssd1 vccd1 vccd1 _1632_/A sky130_fd_sc_hd__dfxtp_4
Xclkbuf_4_7_0_m1_clk_local clkbuf_4_7_0_m1_clk_local/A vssd1 vssd1 vccd1 vccd1 _2670_/CLK
+ sky130_fd_sc_hd__clkbuf_1
X_2506_ _2508_/CLK _2095_/X vssd1 vssd1 vccd1 vccd1 _1219_/A sky130_fd_sc_hd__dfxtp_4
X_1319_ _1317_/Y _1283_/B _1318_/Y vssd1 vssd1 vccd1 vccd1 _1320_/A sky130_fd_sc_hd__nand3_4
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2299_ _1489_/Y _2289_/X _2292_/X _1879_/B _2294_/X vssd1 vssd1 vccd1 vccd1 _2299_/Y
+ sky130_fd_sc_hd__o32ai_4
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1670_ _1666_/X _1667_/Y _1669_/Y vssd1 vssd1 vccd1 vccd1 _1670_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_30_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2222_ _2222_/A _1882_/A vssd1 vssd1 vccd1 vccd1 _2224_/A sky130_fd_sc_hd__nand2_4
XFILLER_23_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2153_ _2140_/Y _2151_/Y _2152_/Y vssd1 vssd1 vccd1 vccd1 _2156_/A sky130_fd_sc_hd__o21ai_4
X_2084_ _2375_/A _2084_/B vssd1 vssd1 vccd1 vccd1 _2514_/D sky130_fd_sc_hd__nor2_4
XFILLER_26_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1937_ _1915_/X _2570_/Q vssd1 vssd1 vccd1 vccd1 _1937_/X sky130_fd_sc_hd__and2_4
X_1868_ _1871_/A _1868_/B vssd1 vssd1 vccd1 vccd1 _1868_/X sky130_fd_sc_hd__and2_4
X_1799_ _2507_/Q vssd1 vssd1 vccd1 vccd1 _1799_/X sky130_fd_sc_hd__buf_2
XFILLER_44_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1653_ _1653_/A _1653_/B vssd1 vssd1 vccd1 vccd1 _1653_/Y sky130_fd_sc_hd__nand2_4
X_1584_ _1247_/A _1531_/X _1582_/X _1583_/X vssd1 vssd1 vccd1 vccd1 _1584_/X sky130_fd_sc_hd__a211o_4
X_1722_ _1243_/X vssd1 vssd1 vccd1 vccd1 _1722_/X sky130_fd_sc_hd__buf_2
X_2205_ _1439_/X _2612_/Q _1577_/A _2149_/X vssd1 vssd1 vccd1 vccd1 _2205_/X sky130_fd_sc_hd__o22a_4
XFILLER_66_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2067_ _2066_/Y _2067_/B vssd1 vssd1 vccd1 vccd1 _2067_/Y sky130_fd_sc_hd__nor2_4
XFILLER_34_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2136_ _2123_/X _2124_/X _2135_/Y _1954_/B _2127_/X vssd1 vssd1 vccd1 vccd1 _2486_/D
+ sky130_fd_sc_hd__o32ai_4
XFILLER_22_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1705_ _1705_/A vssd1 vssd1 vccd1 vccd1 _1705_/Y sky130_fd_sc_hd__inv_2
X_2685_ _2545_/CLK _2685_/D vssd1 vssd1 vccd1 vccd1 _1263_/D sky130_fd_sc_hd__dfxtp_4
X_1636_ _1572_/A vssd1 vssd1 vccd1 vccd1 _2241_/D sky130_fd_sc_hd__buf_2
X_1567_ _1557_/Y _1560_/X _1566_/X vssd1 vssd1 vccd1 vccd1 _1567_/Y sky130_fd_sc_hd__a21boi_4
XFILLER_66_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1498_ _1571_/B vssd1 vssd1 vccd1 vccd1 _1499_/C sky130_fd_sc_hd__buf_2
X_2119_ _2114_/Y _2116_/Y _2118_/Y vssd1 vssd1 vccd1 vccd1 _2492_/D sky130_fd_sc_hd__o21ai_4
XFILLER_13_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_15_0_addressalyzerBlock.SPI_CLK clkbuf_3_7_0_addressalyzerBlock.SPI_CLK/X
+ vssd1 vssd1 vccd1 vccd1 _2707_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_1_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1421_ _1421_/A vssd1 vssd1 vccd1 vccd1 _1421_/Y sky130_fd_sc_hd__inv_2
X_2470_ _2478_/CLK _2470_/D vssd1 vssd1 vccd1 vccd1 _2470_/Q sky130_fd_sc_hd__dfxtp_4
X_1283_ _1272_/X _1283_/B _1282_/Y vssd1 vssd1 vccd1 vccd1 _1284_/A sky130_fd_sc_hd__nand3_4
X_1352_ _1263_/A _1350_/Y _1345_/X _1355_/B vssd1 vssd1 vccd1 vccd1 _1353_/B sky130_fd_sc_hd__nand4_4
X_2668_ _2612_/CLK _1466_/Y vssd1 vssd1 vccd1 vccd1 _2668_/Q sky130_fd_sc_hd__dfxtp_4
X_2599_ _2705_/CLK _2599_/D vssd1 vssd1 vccd1 vccd1 _2599_/Q sky130_fd_sc_hd__dfxtp_4
X_1619_ _1618_/Y vssd1 vssd1 vccd1 vccd1 _1620_/B sky130_fd_sc_hd__inv_2
XFILLER_42_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1970_ _1974_/A _2541_/Q _2542_/Q vssd1 vssd1 vccd1 vccd1 _1971_/C sky130_fd_sc_hd__a21o_4
XFILLER_53_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2522_ _2527_/CLK _2522_/D vssd1 vssd1 vccd1 vccd1 _1984_/A sky130_fd_sc_hd__dfxtp_4
Xclkbuf_4_15_0_m1_clk_local clkbuf_3_7_0_m1_clk_local/X vssd1 vssd1 vccd1 vccd1 _2695_/CLK
+ sky130_fd_sc_hd__clkbuf_1
X_1335_ _1264_/A _1280_/A _1332_/X _1280_/B vssd1 vssd1 vccd1 vccd1 _1335_/Y sky130_fd_sc_hd__nand4_4
X_1404_ _1404_/A vssd1 vssd1 vccd1 vccd1 _1404_/Y sky130_fd_sc_hd__inv_2
X_2384_ _2091_/X _1633_/D _1478_/X vssd1 vssd1 vccd1 vccd1 _2384_/Y sky130_fd_sc_hd__nor3_4
X_2453_ _2478_/CLK _2453_/D vssd1 vssd1 vccd1 vccd1 _2453_/Q sky130_fd_sc_hd__dfxtp_4
X_1266_ _1266_/A _1266_/B _1266_/C _1280_/C vssd1 vssd1 vccd1 vccd1 _1313_/A sky130_fd_sc_hd__nand4_4
XFILLER_56_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1884_ _2472_/Q vssd1 vssd1 vccd1 vccd1 _1884_/Y sky130_fd_sc_hd__inv_2
X_1953_ _1953_/A vssd1 vssd1 vccd1 vccd1 _1954_/B sky130_fd_sc_hd__inv_2
X_2505_ _2508_/CLK _2505_/D vssd1 vssd1 vccd1 vccd1 _2094_/A sky130_fd_sc_hd__dfxtp_4
X_1318_ _1281_/D _1318_/B vssd1 vssd1 vccd1 vccd1 _1318_/Y sky130_fd_sc_hd__nand2_4
X_2436_ _2707_/CLK _2366_/Y vssd1 vssd1 vccd1 vccd1 _2365_/B sky130_fd_sc_hd__dfxtp_4
X_2367_ _1667_/B _1623_/B _2435_/Q vssd1 vssd1 vccd1 vccd1 _2367_/X sky130_fd_sc_hd__o21a_4
XFILLER_29_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2298_ _1700_/Y _2289_/X _2292_/X _1877_/B _2294_/X vssd1 vssd1 vccd1 vccd1 _2476_/D
+ sky130_fd_sc_hd__o32ai_4
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1249_ _1249_/A _1249_/B vssd1 vssd1 vccd1 vccd1 _1277_/A sky130_fd_sc_hd__nand2_4
XFILLER_24_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2152_ _1544_/X _1264_/A _1592_/X vssd1 vssd1 vccd1 vccd1 _2152_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_38_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2221_ _2221_/A _2221_/B _2221_/C vssd1 vssd1 vccd1 vccd1 _2225_/A sky130_fd_sc_hd__nand3_4
X_2083_ _2513_/Q vssd1 vssd1 vccd1 vccd1 _2084_/B sky130_fd_sc_hd__inv_2
X_1867_ _1871_/A _2608_/Q vssd1 vssd1 vccd1 vccd1 _2602_/D sky130_fd_sc_hd__and2_4
X_1936_ _1915_/X _2571_/Q vssd1 vssd1 vccd1 vccd1 _1936_/X sky130_fd_sc_hd__and2_4
X_1798_ _1798_/A vssd1 vssd1 vccd1 vccd1 _1798_/X sky130_fd_sc_hd__buf_2
X_2419_ _2420_/CLK _2419_/D vssd1 vssd1 vccd1 vccd1 _2419_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_16_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1721_ _1688_/Y _1720_/Y _2652_/Q vssd1 vssd1 vccd1 vccd1 _1721_/Y sky130_fd_sc_hd__o21ai_4
X_1652_ _1652_/A vssd1 vssd1 vccd1 vccd1 _1653_/A sky130_fd_sc_hd__buf_2
X_1583_ _1583_/A vssd1 vssd1 vccd1 vccd1 _1583_/X sky130_fd_sc_hd__buf_2
XFILLER_66_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2135_ _1829_/B _2115_/X _1522_/A vssd1 vssd1 vccd1 vccd1 _2135_/Y sky130_fd_sc_hd__nand3_4
X_2204_ _2201_/Y _1560_/X _2203_/Y vssd1 vssd1 vccd1 vccd1 _2204_/Y sky130_fd_sc_hd__a21boi_4
X_2066_ _2066_/A vssd1 vssd1 vccd1 vccd1 _2066_/Y sky130_fd_sc_hd__inv_2
XFILLER_34_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1919_ _1921_/A _1919_/B vssd1 vssd1 vccd1 vccd1 _1919_/Y sky130_fd_sc_hd__nor2_4
XFILLER_57_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2684_ _2564_/CLK _1371_/Y vssd1 vssd1 vccd1 vccd1 _2684_/Q sky130_fd_sc_hd__dfxtp_4
X_1704_ _1703_/Y _1464_/X _1692_/C _1707_/D vssd1 vssd1 vccd1 vccd1 _1705_/A sky130_fd_sc_hd__and4_4
X_1635_ _1635_/A _1635_/B vssd1 vssd1 vccd1 vccd1 _2241_/A sky130_fd_sc_hd__and2_4
X_1497_ _1497_/A vssd1 vssd1 vccd1 vccd1 _1581_/A sky130_fd_sc_hd__buf_2
X_1566_ _2118_/C _2147_/B _1562_/X _1565_/Y vssd1 vssd1 vccd1 vccd1 _1566_/X sky130_fd_sc_hd__a211o_4
XFILLER_66_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2049_ _1984_/A vssd1 vssd1 vccd1 vccd1 _2057_/B sky130_fd_sc_hd__buf_2
X_2118_ _2114_/Y _2117_/X _2118_/C vssd1 vssd1 vccd1 vccd1 _2118_/Y sky130_fd_sc_hd__nand3_4
XFILLER_45_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1351_ _1263_/C vssd1 vssd1 vccd1 vccd1 _1355_/B sky130_fd_sc_hd__buf_2
X_1420_ _1420_/A _1330_/B _1420_/C vssd1 vssd1 vccd1 vccd1 _1421_/A sky130_fd_sc_hd__nand3_4
X_1282_ _2700_/Q _1282_/B _1282_/C _1282_/D vssd1 vssd1 vccd1 vccd1 _1282_/Y sky130_fd_sc_hd__nand4_4
XFILLER_36_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2667_ _2612_/CLK _1476_/Y vssd1 vssd1 vccd1 vccd1 _1540_/B sky130_fd_sc_hd__dfxtp_4
X_1618_ _1618_/A _1618_/B vssd1 vssd1 vccd1 vccd1 _1618_/Y sky130_fd_sc_hd__nand2_4
X_2598_ _2621_/CLK _1871_/X vssd1 vssd1 vccd1 vccd1 _2598_/Q sky130_fd_sc_hd__dfxtp_4
X_1549_ _2493_/Q vssd1 vssd1 vccd1 vccd1 _2143_/A sky130_fd_sc_hd__buf_2
XFILLER_39_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_3_1_0_addressalyzerBlock.SPI_CLK clkbuf_3_1_0_addressalyzerBlock.SPI_CLK/A
+ vssd1 vssd1 vccd1 vccd1 clkbuf_4_2_0_addressalyzerBlock.SPI_CLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_1_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2521_ _2527_/CLK _2065_/Y vssd1 vssd1 vccd1 vccd1 _1983_/A sky130_fd_sc_hd__dfxtp_4
X_1334_ _1264_/A _1333_/X _1311_/X vssd1 vssd1 vccd1 vccd1 _1336_/A sky130_fd_sc_hd__o21a_4
X_1265_ _1265_/A vssd1 vssd1 vccd1 vccd1 _1280_/C sky130_fd_sc_hd__inv_2
X_1403_ _1403_/A _1402_/Y vssd1 vssd1 vccd1 vccd1 _1404_/A sky130_fd_sc_hd__nand2_4
XFILLER_46_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2383_ _1828_/Y _2429_/Q _2096_/X _2382_/X vssd1 vssd1 vccd1 vccd1 _2383_/X sky130_fd_sc_hd__a211o_4
X_2452_ _2478_/CLK _2452_/D vssd1 vssd1 vccd1 vccd1 ID_toHost sky130_fd_sc_hd__dfxtp_4
XFILLER_24_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_2_0_0_m1_clk_local clkbuf_1_0_0_m1_clk_local/X vssd1 vssd1 vccd1 vccd1 clkbuf_2_0_0_m1_clk_local/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_19_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1883_ _1875_/X _1882_/Y vssd1 vssd1 vccd1 vccd1 _1883_/Y sky130_fd_sc_hd__nor2_4
X_1952_ _1946_/A _1952_/B vssd1 vssd1 vccd1 vccd1 _1952_/Y sky130_fd_sc_hd__nor2_4
XFILLER_14_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2435_ _2707_/CLK _2376_/X vssd1 vssd1 vccd1 vccd1 _2435_/Q sky130_fd_sc_hd__dfxtp_4
X_2504_ _2508_/CLK _2098_/X vssd1 vssd1 vccd1 vccd1 _2504_/Q sky130_fd_sc_hd__dfxtp_4
X_1317_ _1313_/Y _1248_/B _1279_/Y vssd1 vssd1 vccd1 vccd1 _1317_/Y sky130_fd_sc_hd__nand3_4
X_1248_ _1248_/A _1248_/B vssd1 vssd1 vccd1 vccd1 _1281_/C sky130_fd_sc_hd__nand2_4
XFILLER_56_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2366_ _2365_/Y _1632_/Y _1722_/X vssd1 vssd1 vccd1 vccd1 _2366_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_2_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2297_ _2296_/Y _2289_/X _2292_/X _1643_/B _2294_/X vssd1 vssd1 vccd1 vccd1 _2297_/Y
+ sky130_fd_sc_hd__o32ai_4
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2151_ _2145_/X _2148_/Y _2150_/X vssd1 vssd1 vccd1 vccd1 _2151_/Y sky130_fd_sc_hd__a21oi_4
X_2082_ _1956_/A _2074_/A vssd1 vssd1 vccd1 vccd1 _2082_/Y sky130_fd_sc_hd__nor2_4
X_2220_ _1414_/A _2220_/B vssd1 vssd1 vccd1 vccd1 _2221_/C sky130_fd_sc_hd__nand2_4
XFILLER_53_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1866_ _1222_/A vssd1 vssd1 vccd1 vccd1 _1871_/A sky130_fd_sc_hd__buf_2
X_1935_ _1915_/X _1935_/B vssd1 vssd1 vccd1 vccd1 _1935_/X sky130_fd_sc_hd__and2_4
X_1797_ _2507_/Q vssd1 vssd1 vccd1 vccd1 _1798_/A sky130_fd_sc_hd__inv_2
X_2418_ _2420_/CLK _2418_/D vssd1 vssd1 vccd1 vccd1 _2419_/D sky130_fd_sc_hd__dfxtp_4
X_2349_ _1522_/Y _2334_/X _2348_/Y vssd1 vssd1 vccd1 vccd1 _2448_/D sky130_fd_sc_hd__o21ai_4
XFILLER_32_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_4_3_0_m1_clk_local clkbuf_4_3_0_m1_clk_local/A vssd1 vssd1 vccd1 vccd1 _2553_/CLK
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_16_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1651_ _1651_/A _1650_/Y vssd1 vssd1 vccd1 vccd1 _1651_/Y sky130_fd_sc_hd__nand2_4
X_1720_ _1712_/X _1714_/X _1717_/C _1717_/D _1488_/X vssd1 vssd1 vccd1 vccd1 _1720_/Y
+ sky130_fd_sc_hd__a41oi_4
X_1582_ _1581_/X vssd1 vssd1 vccd1 vccd1 _1582_/X sky130_fd_sc_hd__buf_2
XFILLER_3_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2065_ _2065_/A vssd1 vssd1 vccd1 vccd1 _2065_/Y sky130_fd_sc_hd__inv_2
X_2134_ _2123_/X _2124_/X _2133_/Y _1952_/B _2127_/X vssd1 vssd1 vccd1 vccd1 _2134_/Y
+ sky130_fd_sc_hd__o32ai_4
X_2203_ _1950_/B _1647_/X _2202_/Y vssd1 vssd1 vccd1 vccd1 _2203_/Y sky130_fd_sc_hd__o21ai_4
X_1849_ _1853_/A DATA_FROM_HASH[0] vssd1 vssd1 vccd1 vccd1 _1849_/X sky130_fd_sc_hd__and2_4
X_1918_ _2470_/Q vssd1 vssd1 vccd1 vccd1 _1919_/B sky130_fd_sc_hd__inv_2
XFILLER_27_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2683_ _2545_/CLK _1375_/Y vssd1 vssd1 vccd1 vccd1 _1369_/C sky130_fd_sc_hd__dfxtp_4
X_1703_ _1460_/Y _1444_/A _1444_/B _1486_/B vssd1 vssd1 vccd1 vccd1 _1703_/Y sky130_fd_sc_hd__nor4_4
X_1634_ _1628_/Y _1633_/Y _1492_/X vssd1 vssd1 vccd1 vccd1 _2658_/D sky130_fd_sc_hd__a21oi_4
XPHY_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1496_ _1496_/A vssd1 vssd1 vccd1 vccd1 _1510_/A sky130_fd_sc_hd__buf_2
X_1565_ _2272_/A _1565_/B vssd1 vssd1 vccd1 vccd1 _1565_/Y sky130_fd_sc_hd__nor2_4
XFILLER_66_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2048_ _1983_/Y _1985_/Y _2048_/C vssd1 vssd1 vccd1 vccd1 _2057_/A sky130_fd_sc_hd__nor3_4
X_2117_ _1776_/X vssd1 vssd1 vccd1 vccd1 _2117_/X sky130_fd_sc_hd__buf_2
XFILLER_22_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1281_ _1276_/Y _1246_/Y _1281_/C _1281_/D vssd1 vssd1 vccd1 vccd1 _1282_/B sky130_fd_sc_hd__nor4_4
X_1350_ _1350_/A _1277_/A _1277_/B _1277_/C vssd1 vssd1 vccd1 vccd1 _1350_/Y sky130_fd_sc_hd__nor4_4
XFILLER_51_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2597_ _2612_/CLK _2597_/D vssd1 vssd1 vccd1 vccd1 _2395_/A sky130_fd_sc_hd__dfxtp_4
X_2666_ _2438_/CLK _2666_/D vssd1 vssd1 vccd1 vccd1 _1676_/D sky130_fd_sc_hd__dfxtp_4
X_1617_ _1611_/Y _1615_/Y _1768_/A vssd1 vssd1 vccd1 vccd1 _1617_/X sky130_fd_sc_hd__a21o_4
XFILLER_8_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1479_ _1477_/Y _1676_/D _1478_/X vssd1 vssd1 vccd1 vccd1 _1479_/Y sky130_fd_sc_hd__a21oi_4
X_1548_ _2250_/B vssd1 vssd1 vccd1 vccd1 _1548_/X sky130_fd_sc_hd__buf_2
XFILLER_50_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1402_ _1255_/A _1401_/X _1255_/B _1396_/X vssd1 vssd1 vccd1 vccd1 _1402_/Y sky130_fd_sc_hd__nand4_4
X_2520_ _2527_/CLK _2520_/D vssd1 vssd1 vccd1 vccd1 _2520_/Q sky130_fd_sc_hd__dfxtp_4
X_2451_ _2493_/CLK _2451_/D vssd1 vssd1 vccd1 vccd1 _2451_/Q sky130_fd_sc_hd__dfxtp_4
X_1264_ _1264_/A _1264_/B vssd1 vssd1 vccd1 vccd1 _1265_/A sky130_fd_sc_hd__nand2_4
X_1333_ _1266_/A _1332_/X _1266_/B _1280_/B vssd1 vssd1 vccd1 vccd1 _1333_/X sky130_fd_sc_hd__and4_4
XFILLER_39_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2382_ _2381_/Y _1207_/A _2382_/C vssd1 vssd1 vccd1 vccd1 _2382_/X sky130_fd_sc_hd__and3_4
XFILLER_51_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2649_ _2495_/CLK _1741_/X vssd1 vssd1 vccd1 vccd1 _1738_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_35_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1882_ _1882_/A vssd1 vssd1 vccd1 vccd1 _1882_/Y sky130_fd_sc_hd__inv_2
X_1951_ _1951_/A vssd1 vssd1 vccd1 vccd1 _1952_/B sky130_fd_sc_hd__inv_2
XFILLER_14_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2365_ _1235_/X _2365_/B vssd1 vssd1 vccd1 vccd1 _2365_/Y sky130_fd_sc_hd__nand2_4
X_2434_ _2508_/CLK _2375_/Y vssd1 vssd1 vccd1 vccd1 _2434_/Q sky130_fd_sc_hd__dfxtp_4
X_2503_ _2655_/CLK _2100_/X vssd1 vssd1 vccd1 vccd1 _2503_/Q sky130_fd_sc_hd__dfxtp_4
X_1247_ _1247_/A _1247_/B vssd1 vssd1 vccd1 vccd1 _1247_/Y sky130_fd_sc_hd__nand2_4
X_1316_ _1315_/Y vssd1 vssd1 vccd1 vccd1 _2694_/D sky130_fd_sc_hd__inv_2
XFILLER_52_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2296_ _1468_/A vssd1 vssd1 vccd1 vccd1 _2296_/Y sky130_fd_sc_hd__inv_2
XFILLER_64_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_4_11_0_m1_clk_local clkbuf_3_5_0_m1_clk_local/X vssd1 vssd1 vccd1 vccd1 _2545_/CLK
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_24_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2150_ _1577_/A _2149_/X _1463_/X _2614_/Q vssd1 vssd1 vccd1 vccd1 _2150_/X sky130_fd_sc_hd__a2bb2o_4
X_2081_ _2074_/A _1986_/B _2080_/Y vssd1 vssd1 vccd1 vccd1 _2081_/X sky130_fd_sc_hd__o21a_4
XFILLER_61_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1934_ _1930_/A _1934_/B vssd1 vssd1 vccd1 vccd1 _2565_/D sky130_fd_sc_hd__nor2_4
XFILLER_14_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1865_ _1865_/A DATA_AVAILABLE[0] vssd1 vssd1 vccd1 vccd1 _2603_/D sky130_fd_sc_hd__and2_4
X_1796_ _1774_/A _2629_/Q _1795_/X vssd1 vssd1 vccd1 vccd1 _2637_/D sky130_fd_sc_hd__o21a_4
X_2417_ _2420_/CLK _2416_/Q vssd1 vssd1 vccd1 vccd1 _2418_/D sky130_fd_sc_hd__dfxtp_4
X_2348_ _2346_/A _2369_/B _2348_/C vssd1 vssd1 vccd1 vccd1 _2348_/Y sky130_fd_sc_hd__nand3_4
X_2279_ _2276_/Y _2277_/Y _2278_/Y vssd1 vssd1 vccd1 vccd1 _2279_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_44_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1581_ _1581_/A vssd1 vssd1 vccd1 vccd1 _1581_/X sky130_fd_sc_hd__buf_2
X_1650_ _1648_/Y _1649_/Y _1463_/X vssd1 vssd1 vccd1 vccd1 _1650_/Y sky130_fd_sc_hd__a21oi_4
X_2202_ _2194_/X _2442_/Q _1559_/X vssd1 vssd1 vccd1 vccd1 _2202_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_21_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2064_ _2053_/X _2055_/Y _2063_/Y vssd1 vssd1 vccd1 vccd1 _2065_/A sky130_fd_sc_hd__o21ai_4
XFILLER_34_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2133_ _1815_/X _1633_/A _1517_/A vssd1 vssd1 vccd1 vccd1 _2133_/Y sky130_fd_sc_hd__nand3_4
X_1917_ _1915_/X _1917_/B vssd1 vssd1 vccd1 vccd1 _1917_/X sky130_fd_sc_hd__and2_4
X_1848_ _1842_/A vssd1 vssd1 vccd1 vccd1 _1853_/A sky130_fd_sc_hd__buf_2
X_1779_ _1964_/B _2636_/Q _1778_/X vssd1 vssd1 vccd1 vccd1 _1779_/X sky130_fd_sc_hd__o21a_4
XFILLER_1_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_4_1_0_addressalyzerBlock.SPI_CLK clkbuf_3_0_0_addressalyzerBlock.SPI_CLK/X
+ vssd1 vssd1 vccd1 vccd1 _2456_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_16_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2682_ _2693_/CLK _2682_/D vssd1 vssd1 vccd1 vccd1 _1249_/A sky130_fd_sc_hd__dfxtp_4
X_1633_ _1633_/A _1632_/Y _1625_/C _1633_/D vssd1 vssd1 vccd1 vccd1 _1633_/Y sky130_fd_sc_hd__nand4_4
X_1564_ _2446_/Q vssd1 vssd1 vccd1 vccd1 _1565_/B sky130_fd_sc_hd__inv_2
X_1702_ _2653_/Q vssd1 vssd1 vccd1 vccd1 _1702_/Y sky130_fd_sc_hd__inv_2
XFILLER_66_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1495_ _2163_/B vssd1 vssd1 vccd1 vccd1 _2241_/B sky130_fd_sc_hd__buf_2
X_2047_ _2009_/X _2035_/X _2046_/Y vssd1 vssd1 vccd1 vccd1 _2047_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_39_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2116_ _1829_/B _2115_/X _1452_/X vssd1 vssd1 vccd1 vccd1 _2116_/Y sky130_fd_sc_hd__nand3_4
XFILLER_1_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_3_6_0_addressalyzerBlock.SPI_CLK clkbuf_3_7_0_addressalyzerBlock.SPI_CLK/A
+ vssd1 vssd1 vccd1 vccd1 clkbuf_3_6_0_addressalyzerBlock.SPI_CLK/X sky130_fd_sc_hd__clkbuf_1
XFILLER_9_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1280_ _1280_/A _1280_/B _1280_/C _1279_/Y vssd1 vssd1 vccd1 vccd1 _1281_/D sky130_fd_sc_hd__nand4_4
XFILLER_63_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2665_ _2438_/CLK _2665_/D vssd1 vssd1 vccd1 vccd1 _1541_/B sky130_fd_sc_hd__dfxtp_4
X_2596_ _2517_/CLK _2596_/D vssd1 vssd1 vccd1 vccd1 _1891_/B sky130_fd_sc_hd__dfxtp_4
X_1616_ _2659_/Q vssd1 vssd1 vccd1 vccd1 _1768_/A sky130_fd_sc_hd__inv_2
X_1547_ _2494_/Q vssd1 vssd1 vccd1 vccd1 _2250_/B sky130_fd_sc_hd__inv_2
X_1478_ _1478_/A vssd1 vssd1 vccd1 vccd1 _1478_/X sky130_fd_sc_hd__buf_2
XFILLER_27_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1401_ _1259_/B vssd1 vssd1 vccd1 vccd1 _1401_/X sky130_fd_sc_hd__buf_2
X_2381_ _2371_/Y _2381_/B _2381_/C vssd1 vssd1 vccd1 vccd1 _2381_/Y sky130_fd_sc_hd__nand3_4
X_2450_ _2494_/CLK _2450_/D vssd1 vssd1 vccd1 vccd1 HASH_LED sky130_fd_sc_hd__dfxtp_4
X_1332_ _1264_/B vssd1 vssd1 vccd1 vccd1 _1332_/X sky130_fd_sc_hd__buf_2
X_1263_ _1263_/A _2687_/Q _1263_/C _1263_/D vssd1 vssd1 vccd1 vccd1 _1266_/C sky130_fd_sc_hd__and4_4
XFILLER_51_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2648_ _2495_/CLK _2648_/D vssd1 vssd1 vccd1 vccd1 _1713_/D sky130_fd_sc_hd__dfxtp_4
X_2579_ _2582_/CLK _1910_/Y vssd1 vssd1 vccd1 vccd1 _1917_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_35_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1950_ _1946_/A _1950_/B vssd1 vssd1 vccd1 vccd1 _2554_/D sky130_fd_sc_hd__nor2_4
X_1881_ _1875_/X _1881_/B vssd1 vssd1 vccd1 vccd1 _1881_/Y sky130_fd_sc_hd__nor2_4
X_2502_ _2655_/CLK _2101_/X vssd1 vssd1 vccd1 vccd1 _2100_/B sky130_fd_sc_hd__dfxtp_4
X_1315_ _1315_/A _1315_/B vssd1 vssd1 vccd1 vccd1 _1315_/Y sky130_fd_sc_hd__nand2_4
XFILLER_51_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2433_ _2514_/CLK _2433_/D vssd1 vssd1 vccd1 vccd1 _1618_/B sky130_fd_sc_hd__dfxtp_4
X_2364_ _2272_/B _2351_/X _2137_/C _2353_/X vssd1 vssd1 vccd1 vccd1 _2364_/X sky130_fd_sc_hd__a2bb2o_4
X_1246_ _2695_/Q vssd1 vssd1 vccd1 vccd1 _1246_/Y sky130_fd_sc_hd__inv_2
X_2295_ _1672_/Y _2289_/X _2292_/X _1555_/B _2294_/X vssd1 vssd1 vccd1 vccd1 _2295_/Y
+ sky130_fd_sc_hd__o32ai_4
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2080_ _2074_/A _1986_/B _2058_/A vssd1 vssd1 vccd1 vccd1 _2080_/Y sky130_fd_sc_hd__a21oi_4
X_1933_ _2463_/Q vssd1 vssd1 vccd1 vccd1 _1934_/B sky130_fd_sc_hd__inv_2
X_1864_ _1865_/A DATA_AVAILABLE[1] vssd1 vssd1 vccd1 vccd1 _2604_/D sky130_fd_sc_hd__and2_4
X_1795_ _2647_/Q _2137_/C _1789_/X vssd1 vssd1 vccd1 vccd1 _1795_/X sky130_fd_sc_hd__o21a_4
X_2278_ _1263_/D _1530_/X _1515_/X _1581_/X _1577_/X vssd1 vssd1 vccd1 vccd1 _2278_/Y
+ sky130_fd_sc_hd__a2111oi_4
XFILLER_29_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2347_ _1517_/Y _2333_/X _2346_/Y vssd1 vssd1 vccd1 vccd1 _2449_/D sky130_fd_sc_hd__o21ai_4
X_2416_ _2420_/CLK _2415_/Q vssd1 vssd1 vccd1 vccd1 _2416_/Q sky130_fd_sc_hd__dfxtp_4
X_1229_ _2703_/Q _1225_/B vssd1 vssd1 vccd1 vccd1 _1229_/X sky130_fd_sc_hd__or2_4
XFILLER_25_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1580_ _1569_/Y _1575_/Y _1579_/Y vssd1 vssd1 vccd1 vccd1 _1580_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_7_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2132_ _2123_/X _2124_/X _2131_/Y _1950_/B _2127_/X vssd1 vssd1 vccd1 vccd1 _2488_/D
+ sky130_fd_sc_hd__o32ai_4
X_2201_ _2197_/Y _2200_/Y vssd1 vssd1 vccd1 vccd1 _2201_/Y sky130_fd_sc_hd__nand2_4
X_2063_ _2055_/Y _2053_/X _1298_/X vssd1 vssd1 vccd1 vccd1 _2063_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_19_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1847_ _1847_/A DATA_FROM_HASH[1] vssd1 vssd1 vccd1 vccd1 _1847_/X sky130_fd_sc_hd__and2_4
X_1916_ _1915_/X _1916_/B vssd1 vssd1 vccd1 vccd1 _2574_/D sky130_fd_sc_hd__and2_4
X_1778_ _1775_/X _1452_/X _1777_/X vssd1 vssd1 vccd1 vccd1 _1778_/X sky130_fd_sc_hd__o21a_4
XFILLER_57_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2681_ _2545_/CLK _2681_/D vssd1 vssd1 vccd1 vccd1 _1249_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_31_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1701_ _1700_/Y _1674_/X _1687_/B vssd1 vssd1 vccd1 vccd1 _1701_/Y sky130_fd_sc_hd__o21ai_4
XPHY_270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1494_ _1637_/C vssd1 vssd1 vccd1 vccd1 _2163_/B sky130_fd_sc_hd__inv_2
X_1632_ _1632_/A vssd1 vssd1 vccd1 vccd1 _1632_/Y sky130_fd_sc_hd__inv_2
X_1563_ _1546_/A vssd1 vssd1 vccd1 vccd1 _2272_/A sky130_fd_sc_hd__buf_2
XFILLER_54_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2115_ _1631_/A vssd1 vssd1 vccd1 vccd1 _2115_/X sky130_fd_sc_hd__buf_2
X_2046_ _2009_/X _2035_/X _1363_/C vssd1 vssd1 vccd1 vccd1 _2046_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_22_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_3_5_0_m1_clk_local clkbuf_3_4_0_m1_clk_local/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_5_0_m1_clk_local/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_63_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2664_ _2438_/CLK _2664_/D vssd1 vssd1 vccd1 vccd1 _1637_/C sky130_fd_sc_hd__dfxtp_4
XFILLER_8_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1477_ _1444_/B _1486_/B vssd1 vssd1 vccd1 vccd1 _1477_/Y sky130_fd_sc_hd__nor2_4
X_1615_ _2381_/B _1608_/B _2381_/C _1614_/Y vssd1 vssd1 vccd1 vccd1 _1615_/Y sky130_fd_sc_hd__nand4_4
X_2595_ _2670_/CLK _1879_/Y vssd1 vssd1 vccd1 vccd1 _2595_/Q sky130_fd_sc_hd__dfxtp_4
X_1546_ _1546_/A vssd1 vssd1 vccd1 vccd1 _1546_/X sky130_fd_sc_hd__buf_2
XFILLER_54_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2029_ _2531_/Q _2027_/X _2028_/Y vssd1 vssd1 vccd1 vccd1 _2029_/X sky130_fd_sc_hd__o21a_4
XFILLER_50_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1331_ _1330_/Y vssd1 vssd1 vccd1 vccd1 _2691_/D sky130_fd_sc_hd__inv_2
X_1400_ _1255_/A _1407_/B _1378_/X vssd1 vssd1 vccd1 vccd1 _1403_/A sky130_fd_sc_hd__o21a_4
X_2380_ _2096_/X _1683_/A _1618_/Y _2381_/B _2372_/X vssd1 vssd1 vccd1 vccd1 _2380_/Y
+ sky130_fd_sc_hd__o32ai_4
XFILLER_5_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1262_ _1277_/B vssd1 vssd1 vccd1 vccd1 _1266_/B sky130_fd_sc_hd__inv_2
XFILLER_17_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2647_ _2511_/CLK _2647_/D vssd1 vssd1 vccd1 vccd1 _2647_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1529_ _1521_/X _1524_/X _1528_/X vssd1 vssd1 vccd1 vccd1 _1529_/Y sky130_fd_sc_hd__a21oi_4
X_2578_ _2561_/CLK _1911_/X vssd1 vssd1 vccd1 vccd1 MACRO_RD_SELECT[5] sky130_fd_sc_hd__dfxtp_4
XFILLER_27_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1880_ _2198_/B vssd1 vssd1 vccd1 vccd1 _1881_/B sky130_fd_sc_hd__inv_2
X_2501_ _2655_/CLK _2102_/X vssd1 vssd1 vccd1 vccd1 _2501_/Q sky130_fd_sc_hd__dfxtp_4
X_1314_ _1248_/A _1313_/Y _1248_/B _1279_/Y vssd1 vssd1 vccd1 vccd1 _1315_/B sky130_fd_sc_hd__nand4_4
XFILLER_44_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2432_ _2707_/CLK _2380_/Y vssd1 vssd1 vccd1 vccd1 _1507_/A sky130_fd_sc_hd__dfxtp_4
X_2363_ _1751_/Y _2351_/X _1522_/A _2353_/X vssd1 vssd1 vccd1 vccd1 _2440_/D sky130_fd_sc_hd__a2bb2o_4
X_2294_ _2293_/X vssd1 vssd1 vccd1 vccd1 _2294_/X sky130_fd_sc_hd__buf_2
XFILLER_64_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1245_ _1238_/Y _1240_/Y _2375_/A vssd1 vssd1 vccd1 vccd1 _1245_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_20_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1863_ _1865_/A DATA_AVAILABLE[2] vssd1 vssd1 vccd1 vccd1 _2605_/D sky130_fd_sc_hd__and2_4
X_1932_ _1930_/A _1932_/B vssd1 vssd1 vccd1 vccd1 _1932_/Y sky130_fd_sc_hd__nor2_4
XFILLER_21_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1794_ _1794_/A vssd1 vssd1 vccd1 vccd1 _2137_/C sky130_fd_sc_hd__buf_2
X_2415_ _2420_/CLK _2414_/Q vssd1 vssd1 vccd1 vccd1 _2415_/Q sky130_fd_sc_hd__dfxtp_4
X_1228_ _1226_/Y _1208_/X _1227_/Y vssd1 vssd1 vccd1 vccd1 _2704_/D sky130_fd_sc_hd__a21oi_4
X_2277_ _1574_/X _1248_/B _1544_/X vssd1 vssd1 vccd1 vccd1 _2277_/Y sky130_fd_sc_hd__a21oi_4
X_2346_ _2346_/A _2369_/B _1432_/A vssd1 vssd1 vccd1 vccd1 _2346_/Y sky130_fd_sc_hd__nand3_4
XFILLER_52_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2062_ _2058_/A _1988_/B _2061_/Y vssd1 vssd1 vccd1 vccd1 _2522_/D sky130_fd_sc_hd__nor3_4
X_2131_ _1815_/X _1633_/A _2640_/Q vssd1 vssd1 vccd1 vccd1 _2131_/Y sky130_fd_sc_hd__nand3_4
X_2200_ _2200_/A _1548_/X _2199_/Y vssd1 vssd1 vccd1 vccd1 _2200_/Y sky130_fd_sc_hd__nand3_4
XFILLER_34_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_6_0_addressalyzerBlock.SPI_CLK clkbuf_4_7_0_addressalyzerBlock.SPI_CLK/A
+ vssd1 vssd1 vccd1 vccd1 _2495_/CLK sky130_fd_sc_hd__clkbuf_1
X_1846_ _1847_/A DATA_FROM_HASH[2] vssd1 vssd1 vccd1 vccd1 _1846_/X sky130_fd_sc_hd__and2_4
X_1915_ _1915_/A vssd1 vssd1 vccd1 vccd1 _1915_/X sky130_fd_sc_hd__buf_2
X_1777_ _1776_/X vssd1 vssd1 vccd1 vccd1 _1777_/X sky130_fd_sc_hd__buf_2
XFILLER_57_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2329_ _1516_/X _2135_/Y _2319_/Y _1908_/B _2321_/X vssd1 vssd1 vccd1 vccd1 _2456_/D
+ sky130_fd_sc_hd__o32ai_4
XFILLER_25_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2680_ _2679_/CLK _1393_/Y vssd1 vssd1 vccd1 vccd1 _1257_/A sky130_fd_sc_hd__dfxtp_4
X_1631_ _1631_/A vssd1 vssd1 vccd1 vccd1 _1633_/A sky130_fd_sc_hd__buf_2
X_1700_ _1481_/A vssd1 vssd1 vccd1 vccd1 _1700_/Y sky130_fd_sc_hd__inv_2
XPHY_260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1493_ _1487_/X _1491_/Y _1492_/X vssd1 vssd1 vccd1 vccd1 _2665_/D sky130_fd_sc_hd__a21oi_4
XFILLER_3_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1562_ _1559_/A vssd1 vssd1 vccd1 vccd1 _1562_/X sky130_fd_sc_hd__buf_2
XFILLER_66_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2045_ _2045_/A vssd1 vssd1 vccd1 vccd1 _2045_/Y sky130_fd_sc_hd__inv_2
XFILLER_39_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2114_ _2111_/X _2112_/X _2113_/X _2353_/D vssd1 vssd1 vccd1 vccd1 _2114_/Y sky130_fd_sc_hd__nand4_4
X_1829_ _1822_/Y _1829_/B _1828_/Y vssd1 vssd1 vccd1 vccd1 _1829_/Y sky130_fd_sc_hd__nand3_4
XFILLER_57_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2663_ _2438_/CLK _1520_/Y vssd1 vssd1 vccd1 vccd1 _1496_/A sky130_fd_sc_hd__dfxtp_4
X_1614_ _2429_/Q vssd1 vssd1 vccd1 vccd1 _1614_/Y sky130_fd_sc_hd__inv_2
X_2594_ _2517_/CLK _1881_/Y vssd1 vssd1 vccd1 vccd1 _2594_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_39_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1476_ _1467_/Y _1473_/Y _1475_/X vssd1 vssd1 vccd1 vccd1 _1476_/Y sky130_fd_sc_hd__a21oi_4
X_1545_ _2493_/Q vssd1 vssd1 vccd1 vccd1 _1546_/A sky130_fd_sc_hd__buf_2
X_2028_ _2026_/X _2012_/A _2531_/Q _2012_/D _1293_/X vssd1 vssd1 vccd1 vccd1 _2028_/Y
+ sky130_fd_sc_hd__a41oi_4
XFILLER_27_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1330_ _1330_/A _1330_/B _1329_/Y vssd1 vssd1 vccd1 vccd1 _1330_/Y sky130_fd_sc_hd__nand3_4
X_1261_ _2684_/Q _1369_/C vssd1 vssd1 vccd1 vccd1 _1277_/B sky130_fd_sc_hd__nand2_4
XFILLER_36_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2577_ _2699_/CLK _1912_/X vssd1 vssd1 vccd1 vccd1 MACRO_RD_SELECT[4] sky130_fd_sc_hd__dfxtp_4
X_2646_ _2508_/CLK _2646_/D vssd1 vssd1 vccd1 vccd1 _1768_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_59_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1459_ _1450_/Y _1453_/Y _1458_/X vssd1 vssd1 vccd1 vccd1 _1459_/X sky130_fd_sc_hd__a21o_4
X_1528_ _1457_/X _1527_/X _1474_/X vssd1 vssd1 vccd1 vccd1 _1528_/X sky130_fd_sc_hd__a21o_4
XFILLER_27_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2431_ _2514_/CLK _2370_/Y vssd1 vssd1 vccd1 vccd1 _1613_/A sky130_fd_sc_hd__dfxtp_4
X_2500_ _2655_/CLK _2500_/D vssd1 vssd1 vccd1 vccd1 _2102_/B sky130_fd_sc_hd__dfxtp_4
X_1313_ _1313_/A vssd1 vssd1 vccd1 vccd1 _1313_/Y sky130_fd_sc_hd__inv_2
XFILLER_56_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2293_ _2158_/X _1527_/X _1535_/X _1631_/A _1242_/A vssd1 vssd1 vccd1 vccd1 _2293_/X
+ sky130_fd_sc_hd__a41o_4
X_1244_ _1243_/X vssd1 vssd1 vccd1 vccd1 _2375_/A sky130_fd_sc_hd__buf_2
X_2362_ _1761_/Y _2352_/X _1517_/A _2354_/X vssd1 vssd1 vccd1 vccd1 _2441_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_24_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2629_ _2511_/CLK _2629_/D vssd1 vssd1 vccd1 vccd1 _2629_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_62_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1862_ _1865_/A DATA_AVAILABLE[3] vssd1 vssd1 vccd1 vccd1 _2606_/D sky130_fd_sc_hd__and2_4
XFILLER_61_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1931_ _2249_/A vssd1 vssd1 vccd1 vccd1 _1932_/B sky130_fd_sc_hd__inv_2
X_1793_ _1774_/A _2630_/Q _1792_/X vssd1 vssd1 vccd1 vccd1 _2638_/D sky130_fd_sc_hd__o21a_4
XFILLER_14_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2414_ _2420_/CLK _2414_/D vssd1 vssd1 vccd1 vccd1 _2414_/Q sky130_fd_sc_hd__dfxtp_4
X_1227_ _2482_/Q _1208_/A _1222_/X vssd1 vssd1 vccd1 vccd1 _1227_/Y sky130_fd_sc_hd__o21ai_4
X_2276_ _1653_/A _2274_/Y _2275_/X vssd1 vssd1 vccd1 vccd1 _2276_/Y sky130_fd_sc_hd__o21ai_4
X_2345_ _2300_/Y _2333_/X _2344_/Y vssd1 vssd1 vccd1 vccd1 _2450_/D sky130_fd_sc_hd__o21ai_4
XFILLER_52_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_11_0_addressalyzerBlock.SPI_CLK clkbuf_3_5_0_addressalyzerBlock.SPI_CLK/X
+ vssd1 vssd1 vccd1 vccd1 _2617_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2061_ _2055_/Y _2053_/X _2057_/B vssd1 vssd1 vccd1 vccd1 _2061_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_34_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2130_ _2123_/X _2124_/X _2129_/Y _1948_/B _2127_/X vssd1 vssd1 vccd1 vccd1 _2489_/D
+ sky130_fd_sc_hd__o32ai_4
XFILLER_34_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1914_ _1912_/A _1914_/B vssd1 vssd1 vccd1 vccd1 _1914_/X sky130_fd_sc_hd__and2_4
XFILLER_22_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1845_ _1847_/A DATA_FROM_HASH[3] vssd1 vssd1 vccd1 vccd1 _2620_/D sky130_fd_sc_hd__and2_4
X_1776_ _2353_/B vssd1 vssd1 vccd1 vccd1 _1776_/X sky130_fd_sc_hd__buf_2
XFILLER_8_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2328_ _1516_/X _2133_/Y _2319_/Y _1904_/Y _2321_/X vssd1 vssd1 vccd1 vccd1 _2457_/D
+ sky130_fd_sc_hd__o32ai_4
XFILLER_65_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2259_ _2242_/X _2257_/Y _2258_/X vssd1 vssd1 vccd1 vccd1 _2259_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_25_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1630_ _2353_/D vssd1 vssd1 vccd1 vccd1 _1631_/A sky130_fd_sc_hd__buf_2
XPHY_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1492_ _1243_/X vssd1 vssd1 vccd1 vccd1 _1492_/X sky130_fd_sc_hd__buf_2
X_1561_ _1546_/A vssd1 vssd1 vccd1 vccd1 _2147_/B sky130_fd_sc_hd__buf_2
XFILLER_54_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2044_ _2044_/A _2005_/B _2043_/Y vssd1 vssd1 vccd1 vccd1 _2045_/A sky130_fd_sc_hd__nand3_4
X_2113_ _1499_/C vssd1 vssd1 vccd1 vccd1 _2113_/X sky130_fd_sc_hd__buf_2
XFILLER_22_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1828_ _1828_/A vssd1 vssd1 vccd1 vccd1 _1828_/Y sky130_fd_sc_hd__inv_2
XFILLER_1_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1759_ _2651_/Q _1758_/Y _1702_/Y _1752_/A vssd1 vssd1 vccd1 vccd1 _1765_/A sky130_fd_sc_hd__o22a_4
XFILLER_57_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1544_ _1544_/A vssd1 vssd1 vccd1 vccd1 _1544_/X sky130_fd_sc_hd__buf_2
X_2662_ _2438_/CLK _1529_/Y vssd1 vssd1 vccd1 vccd1 _1497_/A sky130_fd_sc_hd__dfxtp_4
X_2593_ _2670_/CLK _1883_/Y vssd1 vssd1 vccd1 vccd1 _1894_/B sky130_fd_sc_hd__dfxtp_4
X_1613_ _1613_/A vssd1 vssd1 vccd1 vccd1 _2381_/C sky130_fd_sc_hd__inv_2
XFILLER_5_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1475_ _1458_/X _1460_/Y _1474_/X vssd1 vssd1 vccd1 vccd1 _1475_/X sky130_fd_sc_hd__a21o_4
XFILLER_27_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2027_ _2027_/A _2027_/B _2026_/X _2012_/D vssd1 vssd1 vccd1 vccd1 _2027_/X sky130_fd_sc_hd__and4_4
XFILLER_54_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1260_ _1277_/A _1277_/C vssd1 vssd1 vccd1 vccd1 _1266_/A sky130_fd_sc_hd__nor2_4
XFILLER_36_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_3_1_0_m1_clk_local clkbuf_2_0_0_m1_clk_local/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_3_0_m1_clk_local/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_32_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1527_ _1526_/X vssd1 vssd1 vccd1 vccd1 _1527_/X sky130_fd_sc_hd__buf_2
X_2576_ _2413_/CLK _2576_/D vssd1 vssd1 vccd1 vccd1 MACRO_RD_SELECT[3] sky130_fd_sc_hd__dfxtp_4
X_2645_ _2655_/CLK _2645_/D vssd1 vssd1 vccd1 vccd1 _2393_/A sky130_fd_sc_hd__dfxtp_4
X_1389_ _1259_/B _2679_/Q _1381_/X _1256_/Y vssd1 vssd1 vccd1 vccd1 _1389_/X sky130_fd_sc_hd__and4_4
X_1458_ _1457_/X vssd1 vssd1 vccd1 vccd1 _1458_/X sky130_fd_sc_hd__buf_2
XFILLER_42_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2430_ _2707_/CLK _2373_/Y vssd1 vssd1 vccd1 vccd1 _2371_/A sky130_fd_sc_hd__dfxtp_4
X_2361_ _1758_/Y _2352_/X _1726_/A _2354_/X vssd1 vssd1 vccd1 vccd1 _2361_/X sky130_fd_sc_hd__a2bb2o_4
X_1312_ _1248_/A _1310_/Y _1311_/X vssd1 vssd1 vccd1 vccd1 _1315_/A sky130_fd_sc_hd__o21a_4
X_1243_ _1668_/A vssd1 vssd1 vccd1 vccd1 _1243_/X sky130_fd_sc_hd__buf_2
XFILLER_2_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2292_ _2291_/Y vssd1 vssd1 vccd1 vccd1 _2292_/X sky130_fd_sc_hd__buf_2
XFILLER_20_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2559_ _2559_/CLK _1941_/X vssd1 vssd1 vccd1 vccd1 DATA_TO_HASH[2] sky130_fd_sc_hd__dfxtp_4
X_2628_ _2511_/CLK _2628_/D vssd1 vssd1 vccd1 vccd1 _1747_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_11_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1930_ _1930_/A _1929_/Y vssd1 vssd1 vccd1 vccd1 _1930_/Y sky130_fd_sc_hd__nor2_4
X_1861_ _1865_/A DATA_AVAILABLE[4] vssd1 vssd1 vccd1 vccd1 _2607_/D sky130_fd_sc_hd__and2_4
X_1792_ _2647_/Q _1522_/A _1789_/X vssd1 vssd1 vccd1 vccd1 _1792_/X sky130_fd_sc_hd__o21a_4
XFILLER_6_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2413_ _2413_/CLK _2412_/Q vssd1 vssd1 vccd1 vccd1 _2414_/D sky130_fd_sc_hd__dfxtp_4
X_2344_ _2334_/X _2369_/B HASH_LED vssd1 vssd1 vccd1 vccd1 _2344_/Y sky130_fd_sc_hd__nand3_4
X_1226_ _2703_/Q _1201_/X _1225_/X vssd1 vssd1 vccd1 vccd1 _1226_/Y sky130_fd_sc_hd__o21ai_4
X_2275_ _1439_/X _2609_/Q _1577_/A _2149_/X vssd1 vssd1 vccd1 vccd1 _2275_/X sky130_fd_sc_hd__o22a_4
XFILLER_37_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2060_ _2057_/C _1988_/B _2059_/Y vssd1 vssd1 vccd1 vccd1 _2060_/X sky130_fd_sc_hd__o21a_4
XFILLER_19_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1913_ _1912_/A _1913_/B vssd1 vssd1 vccd1 vccd1 _2576_/D sky130_fd_sc_hd__and2_4
X_1844_ _1847_/A DATA_FROM_HASH[4] vssd1 vssd1 vccd1 vccd1 _1844_/X sky130_fd_sc_hd__and2_4
X_1775_ _2647_/Q vssd1 vssd1 vccd1 vccd1 _1775_/X sky130_fd_sc_hd__buf_2
XFILLER_57_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2258_ _1414_/B _2113_/X _1511_/X _1526_/X _1587_/X vssd1 vssd1 vccd1 vccd1 _2258_/X
+ sky130_fd_sc_hd__a2111o_4
X_2327_ _2317_/X _2131_/Y _2320_/X _1902_/Y _2322_/X vssd1 vssd1 vccd1 vccd1 _2327_/Y
+ sky130_fd_sc_hd__o32ai_4
X_1209_ _1207_/A vssd1 vssd1 vccd1 vccd1 _1209_/X sky130_fd_sc_hd__buf_2
X_2189_ _2190_/A vssd1 vssd1 vccd1 vccd1 _2189_/X sky130_fd_sc_hd__buf_2
XFILLER_40_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1560_ _1559_/X vssd1 vssd1 vccd1 vccd1 _1560_/X sky130_fd_sc_hd__buf_2
XFILLER_66_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2112_ _1526_/X vssd1 vssd1 vccd1 vccd1 _2112_/X sky130_fd_sc_hd__buf_2
X_1491_ _1485_/Y _1490_/Y vssd1 vssd1 vccd1 vccd1 _1491_/Y sky130_fd_sc_hd__nand2_4
XFILLER_3_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2043_ _2009_/X _2035_/X _1981_/Y vssd1 vssd1 vccd1 vccd1 _2043_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_22_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1827_ _1838_/A vssd1 vssd1 vccd1 vccd1 _1829_/B sky130_fd_sc_hd__buf_2
X_1689_ _1683_/B _1683_/D _1478_/X vssd1 vssd1 vccd1 vccd1 _1689_/Y sky130_fd_sc_hd__a21oi_4
X_1758_ _2442_/Q vssd1 vssd1 vccd1 vccd1 _1758_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_2_2_0_addressalyzerBlock.SPI_CLK clkbuf_2_2_0_addressalyzerBlock.SPI_CLK/A
+ vssd1 vssd1 vccd1 vccd1 clkbuf_3_5_0_addressalyzerBlock.SPI_CLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_54_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2661_ _2438_/CLK _1537_/Y vssd1 vssd1 vccd1 vccd1 _1442_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_8_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1543_ _1539_/Y _1583_/A vssd1 vssd1 vccd1 vccd1 _1544_/A sky130_fd_sc_hd__nor2_4
X_1474_ _1668_/A vssd1 vssd1 vccd1 vccd1 _1474_/X sky130_fd_sc_hd__buf_2
X_1612_ _1507_/A vssd1 vssd1 vccd1 vccd1 _2381_/B sky130_fd_sc_hd__inv_2
X_2592_ _2670_/CLK _1885_/Y vssd1 vssd1 vccd1 vccd1 _1895_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_5_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2026_ _2026_/A vssd1 vssd1 vccd1 vccd1 _2026_/X sky130_fd_sc_hd__buf_2
XFILLER_54_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2644_ _2443_/CLK _1779_/X vssd1 vssd1 vccd1 vccd1 _1452_/A sky130_fd_sc_hd__dfxtp_4
X_2575_ _2559_/CLK _1914_/X vssd1 vssd1 vccd1 vccd1 MACRO_RD_SELECT[2] sky130_fd_sc_hd__dfxtp_4
X_1526_ _1571_/C vssd1 vssd1 vccd1 vccd1 _1526_/X sky130_fd_sc_hd__buf_2
X_1457_ _1455_/X _1457_/B vssd1 vssd1 vccd1 vccd1 _1457_/X sky130_fd_sc_hd__and2_4
X_1388_ _1377_/A _1377_/B _1387_/Y vssd1 vssd1 vccd1 vccd1 _2681_/D sky130_fd_sc_hd__a21oi_4
X_2009_ _1989_/A vssd1 vssd1 vccd1 vccd1 _2009_/X sky130_fd_sc_hd__buf_2
XFILLER_23_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1311_ _1378_/A vssd1 vssd1 vccd1 vccd1 _1311_/X sky130_fd_sc_hd__buf_2
X_2291_ _2291_/A vssd1 vssd1 vccd1 vccd1 _2291_/Y sky130_fd_sc_hd__inv_2
X_2360_ _2177_/B _2352_/X _1784_/X _2354_/X vssd1 vssd1 vccd1 vccd1 _2360_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_64_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1242_ _1242_/A vssd1 vssd1 vccd1 vccd1 _1668_/A sky130_fd_sc_hd__buf_2
XFILLER_24_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2627_ _2655_/CLK _1826_/Y vssd1 vssd1 vccd1 vccd1 _1819_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_21_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1509_ _1667_/B _1623_/B _1508_/Y vssd1 vssd1 vccd1 vccd1 _1509_/Y sky130_fd_sc_hd__o21ai_4
X_2558_ _2561_/CLK _1942_/X vssd1 vssd1 vccd1 vccd1 DATA_TO_HASH[1] sky130_fd_sc_hd__dfxtp_4
X_2489_ _2493_/CLK _2489_/D vssd1 vssd1 vccd1 vccd1 _1947_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_55_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1860_ _1842_/A vssd1 vssd1 vccd1 vccd1 _1865_/A sky130_fd_sc_hd__buf_2
XFILLER_36_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1791_ _1774_/A _2631_/Q _1790_/X vssd1 vssd1 vccd1 vccd1 _2639_/D sky130_fd_sc_hd__o21a_4
X_2343_ _1776_/X vssd1 vssd1 vccd1 vccd1 _2369_/B sky130_fd_sc_hd__buf_2
X_2412_ _2413_/CLK _2411_/Q vssd1 vssd1 vccd1 vccd1 _2412_/Q sky130_fd_sc_hd__dfxtp_4
X_2274_ _2270_/Y _1560_/X _2273_/X vssd1 vssd1 vccd1 vccd1 _2274_/Y sky130_fd_sc_hd__a21boi_4
X_1225_ _1225_/A _1225_/B vssd1 vssd1 vccd1 vccd1 _1225_/X sky130_fd_sc_hd__or2_4
XFILLER_52_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1989_ _1989_/A _1981_/Y _1989_/C _1989_/D vssd1 vssd1 vccd1 vccd1 _1992_/B sky130_fd_sc_hd__nor4_4
XFILLER_57_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1843_ _1847_/A DATA_FROM_HASH[5] vssd1 vssd1 vccd1 vccd1 _2622_/D sky130_fd_sc_hd__and2_4
X_1912_ _1912_/A _1912_/B vssd1 vssd1 vccd1 vccd1 _1912_/X sky130_fd_sc_hd__and2_4
XFILLER_8_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1774_ _1774_/A vssd1 vssd1 vccd1 vccd1 _1964_/B sky130_fd_sc_hd__buf_2
X_1208_ _1208_/A vssd1 vssd1 vccd1 vccd1 _1208_/X sky130_fd_sc_hd__buf_2
XFILLER_57_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2257_ _2254_/Y _2255_/Y _2256_/Y vssd1 vssd1 vccd1 vccd1 _2257_/Y sky130_fd_sc_hd__a21oi_4
X_2326_ _2317_/X _2129_/Y _2320_/X _1901_/B _2322_/X vssd1 vssd1 vccd1 vccd1 _2326_/Y
+ sky130_fd_sc_hd__o32ai_4
X_2188_ _2186_/Y _2162_/Y _2187_/Y vssd1 vssd1 vccd1 vccd1 _2188_/X sky130_fd_sc_hd__a21o_4
XFILLER_40_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1490_ _1541_/B _1488_/X _1486_/B _1489_/Y _1469_/X vssd1 vssd1 vccd1 vccd1 _1490_/Y
+ sky130_fd_sc_hd__o32ai_4
X_2042_ _2012_/A vssd1 vssd1 vccd1 vccd1 _2044_/A sky130_fd_sc_hd__inv_2
X_2111_ _1515_/A vssd1 vssd1 vccd1 vccd1 _2111_/X sky130_fd_sc_hd__buf_2
XFILLER_62_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1826_ _1826_/A vssd1 vssd1 vccd1 vccd1 _1826_/Y sky130_fd_sc_hd__inv_2
X_1757_ _1756_/X vssd1 vssd1 vccd1 vccd1 _1770_/B sky130_fd_sc_hd__inv_2
X_1688_ _1685_/Y vssd1 vssd1 vccd1 vccd1 _1688_/Y sky130_fd_sc_hd__inv_2
X_2309_ _1919_/B _2306_/X _1452_/X _2308_/X vssd1 vssd1 vccd1 vccd1 _2470_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_0_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2660_ _2705_/CLK _2660_/D vssd1 vssd1 vccd1 vccd1 _2660_/Q sky130_fd_sc_hd__dfxtp_4
X_1611_ _1608_/Y _1611_/B vssd1 vssd1 vccd1 vccd1 _1611_/Y sky130_fd_sc_hd__nor2_4
XFILLER_8_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1542_ _1637_/C _1635_/A _1635_/B _1542_/D vssd1 vssd1 vccd1 vccd1 _1583_/A sky130_fd_sc_hd__nand4_4
X_1473_ _1694_/A _1470_/Y _1471_/X _1472_/X vssd1 vssd1 vccd1 vccd1 _1473_/Y sky130_fd_sc_hd__a22oi_4
XFILLER_5_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2591_ _2582_/CLK _2591_/D vssd1 vssd1 vccd1 vccd1 _2591_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_54_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2025_ _1981_/A vssd1 vssd1 vccd1 vccd1 _2027_/B sky130_fd_sc_hd__buf_2
XFILLER_39_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1809_ _2632_/Q _1799_/X _1804_/X vssd1 vssd1 vccd1 vccd1 _1809_/X sky130_fd_sc_hd__o21a_4
XFILLER_58_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2643_ _2443_/CLK _1781_/X vssd1 vssd1 vccd1 vccd1 _1468_/A sky130_fd_sc_hd__dfxtp_4
X_2574_ _2582_/CLK _2574_/D vssd1 vssd1 vccd1 vccd1 MACRO_RD_SELECT[1] sky130_fd_sc_hd__dfxtp_4
X_1387_ _1377_/A _1377_/B _1363_/C vssd1 vssd1 vccd1 vccd1 _1387_/Y sky130_fd_sc_hd__o21ai_4
X_1525_ _1497_/A vssd1 vssd1 vccd1 vccd1 _1571_/C sky130_fd_sc_hd__inv_2
X_1456_ _1478_/A _1454_/Y _2429_/Q vssd1 vssd1 vccd1 vccd1 _1457_/B sky130_fd_sc_hd__nand3_4
X_2008_ _2008_/A _2008_/B _2006_/Y _2007_/X vssd1 vssd1 vccd1 vccd1 _2014_/B sky130_fd_sc_hd__nor4_4
XFILLER_55_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1310_ _1318_/B _1281_/D vssd1 vssd1 vccd1 vccd1 _1310_/Y sky130_fd_sc_hd__nor2_4
X_2290_ _1590_/A _2353_/B _1511_/X _2353_/D vssd1 vssd1 vccd1 vccd1 _2291_/A sky130_fd_sc_hd__and4_4
X_1241_ _2331_/A vssd1 vssd1 vccd1 vccd1 _1242_/A sky130_fd_sc_hd__buf_2
XFILLER_2_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2557_ _2413_/CLK _2557_/D vssd1 vssd1 vccd1 vccd1 DATA_TO_HASH[0] sky130_fd_sc_hd__dfxtp_4
X_2626_ _2655_/CLK _2626_/D vssd1 vssd1 vccd1 vccd1 _1822_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_55_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1439_ _1439_/A vssd1 vssd1 vccd1 vccd1 _1439_/X sky130_fd_sc_hd__buf_2
X_1508_ _1581_/A _1499_/C vssd1 vssd1 vccd1 vccd1 _1508_/Y sky130_fd_sc_hd__nand2_4
XFILLER_28_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2488_ _2493_/CLK _2488_/D vssd1 vssd1 vccd1 vccd1 _2488_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_62_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1790_ _2647_/Q _1517_/A _1789_/X vssd1 vssd1 vccd1 vccd1 _1790_/X sky130_fd_sc_hd__o21a_4
X_2411_ _2413_/CLK _1832_/A vssd1 vssd1 vccd1 vccd1 _2411_/Q sky130_fd_sc_hd__dfxtp_4
X_1224_ _1221_/Y _1208_/X _1223_/Y vssd1 vssd1 vccd1 vccd1 _2705_/D sky130_fd_sc_hd__a21oi_4
X_2273_ _2485_/Q _1546_/X _1559_/X _2272_/Y vssd1 vssd1 vccd1 vccd1 _2273_/X sky130_fd_sc_hd__a211o_4
X_2342_ _2169_/Y _2341_/X _1784_/X _2331_/Y vssd1 vssd1 vccd1 vccd1 _2451_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_52_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1988_ _1988_/A _1988_/B _1988_/C _1988_/D vssd1 vssd1 vccd1 vccd1 _1989_/D sky130_fd_sc_hd__nand4_4
X_2609_ _2621_/CLK _2609_/D vssd1 vssd1 vccd1 vccd1 _2609_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_2_3_0_m1_clk_local clkbuf_2_3_0_m1_clk_local/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_7_0_m1_clk_local/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_57_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_3_2_0_addressalyzerBlock.SPI_CLK clkbuf_3_3_0_addressalyzerBlock.SPI_CLK/A
+ vssd1 vssd1 vccd1 vccd1 clkbuf_4_5_0_addressalyzerBlock.SPI_CLK/A sky130_fd_sc_hd__clkbuf_1
X_1842_ _1842_/A vssd1 vssd1 vccd1 vccd1 _1847_/A sky130_fd_sc_hd__buf_2
X_1773_ _2647_/Q vssd1 vssd1 vccd1 vccd1 _1774_/A sky130_fd_sc_hd__inv_2
X_1911_ _1912_/A _1911_/B vssd1 vssd1 vccd1 vccd1 _1911_/X sky130_fd_sc_hd__and2_4
XFILLER_8_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1207_ _1207_/A vssd1 vssd1 vccd1 vccd1 _1208_/A sky130_fd_sc_hd__buf_2
X_2256_ _1263_/C _1530_/X _1515_/A _1581_/A _2139_/X vssd1 vssd1 vccd1 vccd1 _2256_/Y
+ sky130_fd_sc_hd__a2111oi_4
X_2187_ _2601_/Q _2187_/B _2187_/C vssd1 vssd1 vccd1 vccd1 _2187_/Y sky130_fd_sc_hd__nor3_4
X_2325_ _2317_/X _2125_/Y _2320_/X _2141_/B _2322_/X vssd1 vssd1 vccd1 vccd1 _2460_/D
+ sky130_fd_sc_hd__o32ai_4
XFILLER_43_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2041_ _2014_/A _1992_/B _2041_/C vssd1 vssd1 vccd1 vccd1 _2041_/Y sky130_fd_sc_hd__nor3_4
XFILLER_47_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2110_ _1521_/X _1533_/X _1536_/X vssd1 vssd1 vccd1 vccd1 _2493_/D sky130_fd_sc_hd__a21oi_4
XFILLER_62_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1825_ _1819_/B _1823_/Y _1824_/Y vssd1 vssd1 vccd1 vccd1 _1826_/A sky130_fd_sc_hd__a21o_4
X_1756_ _1738_/A _1751_/Y _1753_/Y _1754_/X _1755_/X vssd1 vssd1 vccd1 vccd1 _1756_/X
+ sky130_fd_sc_hd__a2111o_4
Xclkbuf_4_6_0_m1_clk_local clkbuf_4_7_0_m1_clk_local/A vssd1 vssd1 vccd1 vccd1 _2517_/CLK
+ sky130_fd_sc_hd__clkbuf_1
X_2308_ _2307_/X vssd1 vssd1 vccd1 vccd1 _2308_/X sky130_fd_sc_hd__buf_2
X_1687_ _1684_/Y _1687_/B vssd1 vssd1 vccd1 vccd1 _1687_/Y sky130_fd_sc_hd__nand2_4
X_2239_ _2239_/A _2481_/Q vssd1 vssd1 vccd1 vccd1 _2239_/Y sky130_fd_sc_hd__nand2_4
XFILLER_38_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1610_ _1623_/B _1613_/A _1609_/Y vssd1 vssd1 vccd1 vccd1 _1611_/B sky130_fd_sc_hd__o21a_4
X_2590_ _2517_/CLK _1891_/X vssd1 vssd1 vccd1 vccd1 HASH_ADDR[5] sky130_fd_sc_hd__dfxtp_4
XFILLER_8_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1541_ _1676_/D _1541_/B vssd1 vssd1 vccd1 vccd1 _1635_/B sky130_fd_sc_hd__nor2_4
X_1472_ _1457_/B vssd1 vssd1 vccd1 vccd1 _1472_/X sky130_fd_sc_hd__buf_2
X_2024_ _2009_/X _1989_/D vssd1 vssd1 vccd1 vccd1 _2027_/A sky130_fd_sc_hd__nor2_4
XFILLER_35_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1808_ _2632_/Q _1798_/X _1807_/X vssd1 vssd1 vccd1 vccd1 _2633_/D sky130_fd_sc_hd__o21a_4
X_1739_ _1737_/Y _1738_/Y _1733_/X vssd1 vssd1 vccd1 vccd1 _1739_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_65_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1524_ _1522_/Y _1469_/X _1590_/A _1509_/Y vssd1 vssd1 vccd1 vccd1 _1524_/X sky130_fd_sc_hd__o22a_4
X_2573_ _2582_/CLK _1917_/X vssd1 vssd1 vccd1 vccd1 MACRO_RD_SELECT[0] sky130_fd_sc_hd__dfxtp_4
X_2642_ _2443_/CLK _1783_/X vssd1 vssd1 vccd1 vccd1 _1481_/A sky130_fd_sc_hd__dfxtp_4
X_1386_ _1385_/Y vssd1 vssd1 vccd1 vccd1 _2682_/D sky130_fd_sc_hd__inv_2
X_1455_ _1446_/Y _1454_/Y _1205_/Y vssd1 vssd1 vccd1 vccd1 _1455_/X sky130_fd_sc_hd__a21o_4
X_2007_ _2003_/A vssd1 vssd1 vccd1 vccd1 _2007_/X sky130_fd_sc_hd__buf_2
XFILLER_35_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1240_ _2479_/Q _1240_/B vssd1 vssd1 vccd1 vccd1 _1240_/Y sky130_fd_sc_hd__nand2_4
XFILLER_2_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1507_ _1507_/A vssd1 vssd1 vccd1 vccd1 _1623_/B sky130_fd_sc_hd__buf_2
X_2556_ _2581_/CLK _1946_/Y vssd1 vssd1 vccd1 vccd1 _1958_/B sky130_fd_sc_hd__dfxtp_4
X_2487_ _2493_/CLK _2134_/Y vssd1 vssd1 vccd1 vccd1 _1951_/A sky130_fd_sc_hd__dfxtp_4
X_2625_ _2413_/CLK _2625_/D vssd1 vssd1 vccd1 vccd1 _1836_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_55_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1369_ _1355_/A _2684_/Q _1369_/C vssd1 vssd1 vccd1 vccd1 _1370_/B sky130_fd_sc_hd__nand3_4
X_1438_ _1652_/A vssd1 vssd1 vccd1 vccd1 _1439_/A sky130_fd_sc_hd__inv_2
XFILLER_62_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2341_ _1512_/X _1582_/X _1531_/X _2115_/X _2096_/A vssd1 vssd1 vccd1 vccd1 _2341_/X
+ sky130_fd_sc_hd__a41o_4
X_2410_ _2413_/CLK _1833_/A vssd1 vssd1 vccd1 vccd1 _1832_/A sky130_fd_sc_hd__dfxtp_4
X_1223_ _2190_/B _1209_/X _1222_/X vssd1 vssd1 vccd1 vccd1 _1223_/Y sky130_fd_sc_hd__o21ai_4
X_2272_ _2272_/A _2272_/B vssd1 vssd1 vccd1 vccd1 _2272_/Y sky130_fd_sc_hd__nor2_4
XFILLER_60_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1987_ _1983_/Y _1987_/B _1985_/Y _2048_/C vssd1 vssd1 vccd1 vccd1 _1988_/B sky130_fd_sc_hd__nor4_4
XFILLER_20_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2608_ _2621_/CLK _1859_/X vssd1 vssd1 vccd1 vccd1 _2608_/Q sky130_fd_sc_hd__dfxtp_4
X_2539_ _2553_/CLK _1976_/X vssd1 vssd1 vccd1 vccd1 HASH_EN sky130_fd_sc_hd__dfxtp_4
XPHY_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1910_ _1921_/A _1910_/B vssd1 vssd1 vccd1 vccd1 _1910_/Y sky130_fd_sc_hd__nor2_4
X_1841_ _1840_/A DATA_FROM_HASH[6] vssd1 vssd1 vccd1 vccd1 _1841_/X sky130_fd_sc_hd__and2_4
XFILLER_8_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1772_ _1770_/Y _1771_/Y _1722_/X vssd1 vssd1 vccd1 vccd1 _2645_/D sky130_fd_sc_hd__a21oi_4
X_2324_ _2317_/X _2120_/Y _2320_/X _1638_/Y _2322_/X vssd1 vssd1 vccd1 vccd1 _2461_/D
+ sky130_fd_sc_hd__o32ai_4
Xclkbuf_4_14_0_m1_clk_local clkbuf_3_7_0_m1_clk_local/X vssd1 vssd1 vccd1 vccd1 _2699_/CLK
+ sky130_fd_sc_hd__clkbuf_1
X_2255_ _1574_/A _1248_/A _1544_/A vssd1 vssd1 vccd1 vccd1 _2255_/Y sky130_fd_sc_hd__a21oi_4
X_2186_ _2168_/Y _2184_/Y _2185_/X vssd1 vssd1 vccd1 vccd1 _2186_/Y sky130_fd_sc_hd__o21ai_4
X_1206_ _1205_/Y vssd1 vssd1 vccd1 vccd1 _1207_/A sky130_fd_sc_hd__buf_2
XFILLER_56_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2040_ _2027_/A _2027_/B _2026_/X vssd1 vssd1 vccd1 vccd1 _2041_/C sky130_fd_sc_hd__a21oi_4
XFILLER_62_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1824_ _1819_/B _1823_/Y _1748_/Y vssd1 vssd1 vccd1 vccd1 _1824_/Y sky130_fd_sc_hd__o21ai_4
X_1686_ _1685_/Y vssd1 vssd1 vccd1 vccd1 _1687_/B sky130_fd_sc_hd__buf_2
X_1755_ _2654_/Q _1755_/B vssd1 vssd1 vccd1 vccd1 _1755_/X sky130_fd_sc_hd__xor2_4
X_2238_ _2217_/X _2237_/Y _2189_/X vssd1 vssd1 vccd1 vccd1 _2238_/Y sky130_fd_sc_hd__o21ai_4
X_2307_ _1539_/A _2287_/Y _1512_/X vssd1 vssd1 vccd1 vccd1 _2307_/X sky130_fd_sc_hd__and3_4
XFILLER_38_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2169_ _2451_/Q vssd1 vssd1 vccd1 vccd1 _2169_/Y sky130_fd_sc_hd__inv_2
XFILLER_21_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1540_ _2668_/Q _1540_/B vssd1 vssd1 vccd1 vccd1 _1635_/A sky130_fd_sc_hd__nor2_4
XFILLER_39_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1471_ _1455_/X vssd1 vssd1 vccd1 vccd1 _1471_/X sky130_fd_sc_hd__buf_2
XFILLER_10_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2023_ _2021_/X _2023_/B _2007_/X vssd1 vssd1 vccd1 vccd1 _2023_/X sky130_fd_sc_hd__and3_4
XFILLER_54_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1807_ _2633_/Q _1799_/X _1804_/X vssd1 vssd1 vccd1 vccd1 _1807_/X sky130_fd_sc_hd__o21a_4
XFILLER_49_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1669_ _1666_/X _2165_/A _2096_/A vssd1 vssd1 vccd1 vccd1 _1669_/Y sky130_fd_sc_hd__a21oi_4
X_1738_ _1738_/A vssd1 vssd1 vccd1 vccd1 _1738_/Y sky130_fd_sc_hd__inv_2
XFILLER_45_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1523_ _1497_/A _1571_/B vssd1 vssd1 vccd1 vccd1 _1590_/A sky130_fd_sc_hd__nor2_4
X_1454_ _1618_/B _2434_/Q vssd1 vssd1 vccd1 vccd1 _1454_/Y sky130_fd_sc_hd__nor2_4
X_2572_ _2670_/CLK _1919_/Y vssd1 vssd1 vccd1 vccd1 _1935_/B sky130_fd_sc_hd__dfxtp_4
X_2641_ _2443_/CLK _1786_/X vssd1 vssd1 vccd1 vccd1 _1489_/A sky130_fd_sc_hd__dfxtp_4
X_1385_ _1385_/A _1384_/Y vssd1 vssd1 vccd1 vccd1 _1385_/Y sky130_fd_sc_hd__nand2_4
XFILLER_27_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2006_ _2000_/A vssd1 vssd1 vccd1 vccd1 _2006_/Y sky130_fd_sc_hd__inv_2
XFILLER_58_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2624_ _2617_/CLK _2624_/D vssd1 vssd1 vccd1 vccd1 _1850_/B sky130_fd_sc_hd__dfxtp_4
X_1437_ _2668_/Q vssd1 vssd1 vccd1 vccd1 _1652_/A sky130_fd_sc_hd__buf_2
X_1506_ _2371_/A vssd1 vssd1 vccd1 vccd1 _1667_/B sky130_fd_sc_hd__buf_2
X_2486_ _2493_/CLK _2486_/D vssd1 vssd1 vccd1 vccd1 _1953_/A sky130_fd_sc_hd__dfxtp_4
Xclkbuf_4_2_0_addressalyzerBlock.SPI_CLK clkbuf_4_2_0_addressalyzerBlock.SPI_CLK/A
+ vssd1 vssd1 vccd1 vccd1 _2494_/CLK sky130_fd_sc_hd__clkbuf_1
X_2555_ _2553_/CLK _1948_/Y vssd1 vssd1 vccd1 vccd1 _2555_/Q sky130_fd_sc_hd__dfxtp_4
X_1368_ _2684_/Q _1367_/Y _1311_/X vssd1 vssd1 vccd1 vccd1 _1368_/X sky130_fd_sc_hd__o21a_4
X_1299_ _1298_/X vssd1 vssd1 vccd1 vccd1 _1956_/A sky130_fd_sc_hd__buf_2
XFILLER_61_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_3_7_0_addressalyzerBlock.SPI_CLK clkbuf_3_7_0_addressalyzerBlock.SPI_CLK/A
+ vssd1 vssd1 vccd1 vccd1 clkbuf_3_7_0_addressalyzerBlock.SPI_CLK/X sky130_fd_sc_hd__clkbuf_1
XFILLER_10_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2340_ _1700_/Y _2333_/X _2339_/Y vssd1 vssd1 vccd1 vccd1 _2452_/D sky130_fd_sc_hd__o21ai_4
X_2271_ _1754_/B vssd1 vssd1 vccd1 vccd1 _2272_/B sky130_fd_sc_hd__inv_2
X_1222_ _1222_/A vssd1 vssd1 vccd1 vccd1 _1222_/X sky130_fd_sc_hd__buf_2
XFILLER_37_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1986_ _2515_/Q _1986_/B _1986_/C _1986_/D vssd1 vssd1 vccd1 vccd1 _2048_/C sky130_fd_sc_hd__nand4_4
X_2607_ _2612_/CLK _2607_/D vssd1 vssd1 vccd1 vccd1 _1868_/B sky130_fd_sc_hd__dfxtp_4
X_2538_ _2693_/CLK _1978_/Y vssd1 vssd1 vccd1 vccd1 _1976_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_28_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2469_ _2456_/CLK _2469_/D vssd1 vssd1 vccd1 vccd1 _2469_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1840_ _1840_/A DATA_FROM_HASH[7] vssd1 vssd1 vccd1 vccd1 _2624_/D sky130_fd_sc_hd__and2_4
XFILLER_42_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1771_ _1768_/A _2393_/A vssd1 vssd1 vccd1 vccd1 _1771_/Y sky130_fd_sc_hd__nand2_4
X_2254_ _1463_/X _2252_/Y _2253_/X vssd1 vssd1 vccd1 vccd1 _2254_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_40_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2323_ _2317_/X _2116_/Y _2320_/X _1550_/Y _2322_/X vssd1 vssd1 vccd1 vccd1 _2462_/D
+ sky130_fd_sc_hd__o32ai_4
X_2185_ _1419_/C _1656_/X _2158_/X _2112_/X _1594_/C vssd1 vssd1 vccd1 vccd1 _2185_/X
+ sky130_fd_sc_hd__a2111o_4
X_1205_ _1618_/A vssd1 vssd1 vccd1 vccd1 _1205_/Y sky130_fd_sc_hd__inv_2
XFILLER_40_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1969_ _1833_/Y _1974_/C vssd1 vssd1 vccd1 vccd1 _1969_/Y sky130_fd_sc_hd__nor2_4
XFILLER_48_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1823_ _1822_/Y vssd1 vssd1 vccd1 vccd1 _1823_/Y sky130_fd_sc_hd__inv_2
X_1685_ _1471_/X _1472_/X _1620_/B vssd1 vssd1 vccd1 vccd1 _1685_/Y sky130_fd_sc_hd__a21oi_4
X_1754_ _1713_/D _1754_/B vssd1 vssd1 vccd1 vccd1 _1754_/X sky130_fd_sc_hd__xor2_4
X_2237_ _2235_/Y _2236_/Y _2162_/A vssd1 vssd1 vccd1 vccd1 _2237_/Y sky130_fd_sc_hd__a21oi_4
X_2306_ _2305_/X vssd1 vssd1 vccd1 vccd1 _2306_/X sky130_fd_sc_hd__buf_2
XFILLER_53_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2168_ _1377_/A _2111_/X _1591_/A _1577_/X _2167_/X vssd1 vssd1 vccd1 vccd1 _2168_/Y
+ sky130_fd_sc_hd__o41ai_4
XFILLER_38_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2099_ _1222_/A vssd1 vssd1 vccd1 vccd1 _2099_/X sky130_fd_sc_hd__buf_2
XFILLER_21_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1470_ _1469_/X vssd1 vssd1 vccd1 vccd1 _1470_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2022_ _1274_/X vssd1 vssd1 vccd1 vccd1 _2023_/B sky130_fd_sc_hd__buf_2
X_1806_ _2633_/Q _1798_/X _1805_/X vssd1 vssd1 vccd1 vccd1 _2634_/D sky130_fd_sc_hd__o21a_4
X_1599_ _2187_/C _1598_/Y _1587_/X vssd1 vssd1 vccd1 vccd1 _1600_/B sky130_fd_sc_hd__a21oi_4
X_1668_ _1668_/A vssd1 vssd1 vccd1 vccd1 _2096_/A sky130_fd_sc_hd__buf_2
X_1737_ _1714_/X vssd1 vssd1 vccd1 vccd1 _1737_/Y sky130_fd_sc_hd__inv_2
XFILLER_53_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_4_2_0_m1_clk_local clkbuf_4_3_0_m1_clk_local/A vssd1 vssd1 vccd1 vccd1 _2561_/CLK
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_49_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2640_ _2443_/CLK _2640_/D vssd1 vssd1 vccd1 vccd1 _2640_/Q sky130_fd_sc_hd__dfxtp_4
X_1453_ _1618_/B _2378_/B _1452_/X vssd1 vssd1 vccd1 vccd1 _1453_/Y sky130_fd_sc_hd__o21ai_4
X_2571_ _2581_/CLK _1921_/Y vssd1 vssd1 vccd1 vccd1 _2571_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_4_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1522_ _1522_/A vssd1 vssd1 vccd1 vccd1 _1522_/Y sky130_fd_sc_hd__inv_2
X_2005_ _2004_/X _2005_/B _1996_/A vssd1 vssd1 vccd1 vccd1 _2005_/X sky130_fd_sc_hd__and3_4
X_1384_ _1249_/A _1394_/A _1249_/B _1384_/D vssd1 vssd1 vccd1 vccd1 _1384_/Y sky130_fd_sc_hd__nand4_4
XFILLER_50_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2623_ _2617_/CLK _1841_/X vssd1 vssd1 vccd1 vccd1 _2623_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_9_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2554_ _2553_/CLK _2554_/D vssd1 vssd1 vccd1 vccd1 _1960_/B sky130_fd_sc_hd__dfxtp_4
X_1367_ _1367_/A _1277_/A _1377_/B vssd1 vssd1 vccd1 vccd1 _1367_/Y sky130_fd_sc_hd__nor3_4
X_1505_ _1501_/X _1503_/Y _1504_/X vssd1 vssd1 vccd1 vccd1 _2664_/D sky130_fd_sc_hd__a21oi_4
X_1436_ _1432_/A _1432_/C _1435_/Y vssd1 vssd1 vccd1 vccd1 _1436_/X sky130_fd_sc_hd__o21a_4
X_2485_ _2493_/CLK _2485_/D vssd1 vssd1 vccd1 vccd1 _2485_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_55_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1298_ _1293_/A vssd1 vssd1 vccd1 vccd1 _1298_/X sky130_fd_sc_hd__buf_2
XFILLER_11_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1221_ _1225_/A _1201_/X _1220_/X vssd1 vssd1 vccd1 vccd1 _1221_/Y sky130_fd_sc_hd__o21ai_4
X_2270_ _2267_/Y _2270_/B vssd1 vssd1 vccd1 vccd1 _2270_/Y sky130_fd_sc_hd__nand2_4
XFILLER_60_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1985_ _2066_/A _2520_/Q vssd1 vssd1 vccd1 vccd1 _1985_/Y sky130_fd_sc_hd__nand2_4
X_2537_ _2545_/CLK _2002_/Y vssd1 vssd1 vccd1 vccd1 CLK_LED sky130_fd_sc_hd__dfxtp_4
X_2606_ _2621_/CLK _2606_/D vssd1 vssd1 vccd1 vccd1 _1869_/B sky130_fd_sc_hd__dfxtp_4
X_2399_ _2660_/Q _1208_/A _1222_/X vssd1 vssd1 vccd1 vccd1 _2399_/Y sky130_fd_sc_hd__o21ai_4
X_1419_ _1419_/A _2674_/Q _1419_/C vssd1 vssd1 vccd1 vccd1 _1420_/C sky130_fd_sc_hd__nand3_4
X_2468_ _2456_/CLK _2311_/X vssd1 vssd1 vccd1 vccd1 _1922_/A sky130_fd_sc_hd__dfxtp_4
XPHY_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1770_ _2659_/Q _1770_/B _1770_/C _1770_/D vssd1 vssd1 vccd1 vccd1 _1770_/Y sky130_fd_sc_hd__nand4_4
X_2253_ _1439_/A _2610_/Q _1573_/A _2149_/A vssd1 vssd1 vccd1 vccd1 _2253_/X sky130_fd_sc_hd__o22a_4
X_2184_ _2181_/Y _2182_/Y _2183_/Y vssd1 vssd1 vccd1 vccd1 _2184_/Y sky130_fd_sc_hd__a21oi_4
X_1204_ _2706_/Q _1201_/X _1203_/X vssd1 vssd1 vccd1 vccd1 _1204_/Y sky130_fd_sc_hd__o21ai_4
X_2322_ _2321_/X vssd1 vssd1 vccd1 vccd1 _2322_/X sky130_fd_sc_hd__buf_2
XFILLER_18_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1899_ _1901_/A _2141_/B vssd1 vssd1 vccd1 vccd1 _1899_/Y sky130_fd_sc_hd__nor2_4
X_1968_ _1833_/Y _1974_/C _1967_/Y vssd1 vssd1 vccd1 vccd1 _2543_/D sky130_fd_sc_hd__nor3_4
XFILLER_17_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1822_ _1219_/A _1822_/B vssd1 vssd1 vccd1 vccd1 _1822_/Y sky130_fd_sc_hd__nand2_4
X_1753_ _1707_/A _1753_/B vssd1 vssd1 vccd1 vccd1 _1753_/Y sky130_fd_sc_hd__nor2_4
X_1684_ _1672_/Y _1674_/X _1683_/Y vssd1 vssd1 vccd1 vccd1 _1684_/Y sky130_fd_sc_hd__o21ai_4
X_2236_ _2260_/A THREAD_COUNT[2] vssd1 vssd1 vccd1 vccd1 _2236_/Y sky130_fd_sc_hd__nand2_4
X_2167_ _1500_/A _1587_/A vssd1 vssd1 vccd1 vccd1 _2167_/X sky130_fd_sc_hd__or2_4
X_2305_ _1512_/X _1527_/X _1531_/X _1631_/A _1242_/A vssd1 vssd1 vccd1 vccd1 _2305_/X
+ sky130_fd_sc_hd__a41o_4
XFILLER_53_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2098_ _1243_/X SCSN_fromHost vssd1 vssd1 vccd1 vccd1 _2098_/X sky130_fd_sc_hd__or2_4
Xclkbuf_4_10_0_m1_clk_local clkbuf_3_5_0_m1_clk_local/X vssd1 vssd1 vccd1 vccd1 _2679_/CLK
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_56_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2021_ _2012_/A _2026_/A _2531_/Q _2012_/D _2532_/Q vssd1 vssd1 vccd1 vccd1 _2021_/X
+ sky130_fd_sc_hd__a41o_4
XFILLER_50_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1805_ _2634_/Q _1799_/X _1804_/X vssd1 vssd1 vccd1 vccd1 _1805_/X sky130_fd_sc_hd__o21a_4
X_1736_ _1522_/Y _1674_/X _1687_/B vssd1 vssd1 vccd1 vccd1 _1736_/Y sky130_fd_sc_hd__o21ai_4
X_1667_ _1632_/A _1667_/B _2435_/Q vssd1 vssd1 vccd1 vccd1 _1667_/Y sky130_fd_sc_hd__nor3_4
X_1598_ _1571_/C _1510_/A _1571_/B vssd1 vssd1 vccd1 vccd1 _1598_/Y sky130_fd_sc_hd__nand3_4
XFILLER_26_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2219_ _2194_/X _1904_/A vssd1 vssd1 vccd1 vccd1 _2221_/A sky130_fd_sc_hd__nand2_4
XFILLER_41_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2570_ _2582_/CLK _2570_/D vssd1 vssd1 vccd1 vccd1 _2570_/Q sky130_fd_sc_hd__dfxtp_4
X_1383_ _1382_/X vssd1 vssd1 vccd1 vccd1 _1394_/A sky130_fd_sc_hd__buf_2
X_1521_ _1485_/Y vssd1 vssd1 vccd1 vccd1 _1521_/X sky130_fd_sc_hd__buf_2
XFILLER_4_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1452_ _1452_/A vssd1 vssd1 vccd1 vccd1 _1452_/X sky130_fd_sc_hd__buf_2
X_2004_ _2003_/Y _1979_/A _2534_/Q _2000_/A _2536_/Q vssd1 vssd1 vccd1 vccd1 _2004_/X
+ sky130_fd_sc_hd__a41o_4
XFILLER_23_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2699_ _2699_/CLK _1289_/X vssd1 vssd1 vccd1 vccd1 _1282_/C sky130_fd_sc_hd__dfxtp_4
Xclkbuf_4_7_0_addressalyzerBlock.SPI_CLK clkbuf_4_7_0_addressalyzerBlock.SPI_CLK/A
+ vssd1 vssd1 vccd1 vccd1 _2655_/CLK sky130_fd_sc_hd__clkbuf_1
X_1719_ _1719_/A _1687_/B vssd1 vssd1 vccd1 vccd1 _1719_/Y sky130_fd_sc_hd__nand2_4
XFILLER_58_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2622_ _2621_/CLK _2622_/D vssd1 vssd1 vccd1 vccd1 _2622_/Q sky130_fd_sc_hd__dfxtp_4
X_1504_ _1458_/X _2241_/B _1474_/X vssd1 vssd1 vccd1 vccd1 _1504_/X sky130_fd_sc_hd__a21o_4
X_2553_ _2553_/CLK _1952_/Y vssd1 vssd1 vccd1 vccd1 _2553_/Q sky130_fd_sc_hd__dfxtp_4
X_2484_ _2705_/CLK _2166_/Y vssd1 vssd1 vccd1 vccd1 _2165_/B sky130_fd_sc_hd__dfxtp_4
X_1366_ _1277_/C vssd1 vssd1 vccd1 vccd1 _1377_/B sky130_fd_sc_hd__buf_2
X_1435_ _1432_/A _1432_/C _2058_/A vssd1 vssd1 vccd1 vccd1 _1435_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_28_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1297_ _1297_/A vssd1 vssd1 vccd1 vccd1 _1297_/Y sky130_fd_sc_hd__inv_2
XFILLER_11_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1220_ _1220_/A _1225_/B vssd1 vssd1 vccd1 vccd1 _1220_/X sky130_fd_sc_hd__or2_4
XFILLER_33_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1984_ _1984_/A vssd1 vssd1 vccd1 vccd1 _1987_/B sky130_fd_sc_hd__inv_2
XFILLER_20_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2536_ _2564_/CLK _2005_/X vssd1 vssd1 vccd1 vccd1 _2536_/Q sky130_fd_sc_hd__dfxtp_4
X_2605_ _2612_/CLK _2605_/D vssd1 vssd1 vccd1 vccd1 _2605_/Q sky130_fd_sc_hd__dfxtp_4
X_2467_ _2456_/CLK _2467_/D vssd1 vssd1 vccd1 vccd1 _1925_/A sky130_fd_sc_hd__dfxtp_4
X_1349_ _1263_/D vssd1 vssd1 vccd1 vccd1 _1350_/A sky130_fd_sc_hd__inv_2
X_2398_ _1203_/A _1201_/A _2397_/X vssd1 vssd1 vccd1 vccd1 _2398_/Y sky130_fd_sc_hd__o21ai_4
X_1418_ _1254_/B _1254_/D vssd1 vssd1 vccd1 vccd1 _1419_/A sky130_fd_sc_hd__nor2_4
XFILLER_28_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2321_ _2158_/X _1535_/X _1582_/X _2353_/D _1242_/A vssd1 vssd1 vccd1 vccd1 _2321_/X
+ sky130_fd_sc_hd__a41o_4
XFILLER_6_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2183_ _1332_/X _2113_/X _1515_/X _1581_/X _1577_/X vssd1 vssd1 vccd1 vccd1 _2183_/Y
+ sky130_fd_sc_hd__a2111oi_4
X_1203_ _1203_/A _1203_/B vssd1 vssd1 vccd1 vccd1 _1203_/X sky130_fd_sc_hd__or2_4
XFILLER_26_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2252_ _2243_/Y _2244_/Y _2251_/Y _1562_/X vssd1 vssd1 vccd1 vccd1 _2252_/Y sky130_fd_sc_hd__a22oi_4
XFILLER_25_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1967_ _1971_/B _1966_/A _1966_/Y vssd1 vssd1 vccd1 vccd1 _1967_/Y sky130_fd_sc_hd__a21oi_4
X_1898_ _2460_/Q vssd1 vssd1 vccd1 vccd1 _2141_/B sky130_fd_sc_hd__inv_2
X_2519_ _2527_/CLK _2072_/Y vssd1 vssd1 vccd1 vccd1 _2066_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_56_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1683_ _1683_/A _1683_/B _1448_/Y _1683_/D vssd1 vssd1 vccd1 vccd1 _1683_/Y sky130_fd_sc_hd__nand4_4
X_1821_ _1818_/Y _1819_/Y _1820_/Y vssd1 vssd1 vccd1 vccd1 _2628_/D sky130_fd_sc_hd__a21oi_4
X_1752_ _1752_/A vssd1 vssd1 vccd1 vccd1 _1753_/B sky130_fd_sc_hd__inv_2
X_2304_ _1532_/Y _2288_/Y _2291_/Y _1888_/B _2293_/X vssd1 vssd1 vccd1 vccd1 _2471_/D
+ sky130_fd_sc_hd__o32ai_4
XFILLER_57_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2235_ _2218_/Y _2233_/Y _2234_/X vssd1 vssd1 vccd1 vccd1 _2235_/Y sky130_fd_sc_hd__o21ai_4
X_2166_ _2239_/A _2164_/Y _2165_/Y vssd1 vssd1 vccd1 vccd1 _2166_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_38_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2097_ _2096_/X _2504_/Q vssd1 vssd1 vccd1 vccd1 _2505_/D sky130_fd_sc_hd__or2_4
XFILLER_21_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2020_ _2008_/A _2007_/X _2019_/Y vssd1 vssd1 vccd1 vccd1 _2533_/D sky130_fd_sc_hd__a21oi_4
XFILLER_47_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1666_ _1664_/C _1478_/A _1664_/Y _1665_/Y vssd1 vssd1 vccd1 vccd1 _1666_/X sky130_fd_sc_hd__a211o_4
X_1804_ _1838_/A vssd1 vssd1 vccd1 vccd1 _1804_/X sky130_fd_sc_hd__buf_2
X_1735_ _1732_/Y _1734_/X _1722_/X vssd1 vssd1 vccd1 vccd1 _2650_/D sky130_fd_sc_hd__a21oi_4
X_1597_ _2190_/A vssd1 vssd1 vccd1 vccd1 _2165_/A sky130_fd_sc_hd__inv_2
X_2149_ _2149_/A vssd1 vssd1 vccd1 vccd1 _2149_/X sky130_fd_sc_hd__buf_2
X_2218_ _1395_/Y _2111_/X _1591_/A _1577_/X _2167_/X vssd1 vssd1 vccd1 vccd1 _2218_/Y
+ sky130_fd_sc_hd__o41ai_4
XFILLER_41_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0_m1_clk_local clkbuf_0_m1_clk_local/X vssd1 vssd1 vccd1 vccd1 clkbuf_2_3_0_m1_clk_local/A
+ sky130_fd_sc_hd__clkbuf_1
X_1520_ _1513_/X _1519_/X _1492_/X vssd1 vssd1 vccd1 vccd1 _1520_/Y sky130_fd_sc_hd__a21oi_4
X_1382_ _1382_/A _1381_/X _1382_/C _1256_/Y vssd1 vssd1 vccd1 vccd1 _1382_/X sky130_fd_sc_hd__and4_4
Xclkbuf_4_12_0_addressalyzerBlock.SPI_CLK clkbuf_3_6_0_addressalyzerBlock.SPI_CLK/X
+ vssd1 vssd1 vccd1 vccd1 _2514_/CLK sky130_fd_sc_hd__clkbuf_1
X_1451_ _2434_/Q vssd1 vssd1 vccd1 vccd1 _2378_/B sky130_fd_sc_hd__buf_2
X_2003_ _2003_/A vssd1 vssd1 vccd1 vccd1 _2003_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2698_ _2699_/CLK _1297_/Y vssd1 vssd1 vccd1 vccd1 _1295_/A sky130_fd_sc_hd__dfxtp_4
X_1649_ _1649_/A _2147_/B vssd1 vssd1 vccd1 vccd1 _1649_/Y sky130_fd_sc_hd__nand2_4
X_1718_ _2652_/Q _1478_/X _1717_/Y _1489_/Y _1673_/Y vssd1 vssd1 vccd1 vccd1 _1719_/A
+ sky130_fd_sc_hd__o32ai_4
XFILLER_58_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2621_ _2621_/CLK _1844_/X vssd1 vssd1 vccd1 vccd1 _2621_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_56_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2483_ _2705_/CLK _2191_/Y vssd1 vssd1 vccd1 vccd1 _2190_/B sky130_fd_sc_hd__dfxtp_4
X_1503_ _1726_/A _1470_/Y _1471_/X _1472_/X vssd1 vssd1 vccd1 vccd1 _1503_/Y sky130_fd_sc_hd__a22oi_4
X_2552_ _2553_/CLK _1954_/Y vssd1 vssd1 vccd1 vccd1 _2552_/Q sky130_fd_sc_hd__dfxtp_4
X_1296_ _1294_/Y _1296_/B vssd1 vssd1 vccd1 vccd1 _1297_/A sky130_fd_sc_hd__nand2_4
XFILLER_55_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1365_ _1369_/C vssd1 vssd1 vccd1 vccd1 _1367_/A sky130_fd_sc_hd__inv_2
X_1434_ _1434_/A vssd1 vssd1 vccd1 vccd1 _2670_/D sky130_fd_sc_hd__inv_2
XFILLER_63_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_3_4_0_m1_clk_local clkbuf_3_4_0_m1_clk_local/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_9_0_m1_clk_local/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_37_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2604_ _2621_/CLK _2604_/D vssd1 vssd1 vccd1 vccd1 _1871_/B sky130_fd_sc_hd__dfxtp_4
X_1983_ _1983_/A vssd1 vssd1 vccd1 vccd1 _1983_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2535_ _2564_/CLK _2014_/Y vssd1 vssd1 vccd1 vccd1 _2000_/A sky130_fd_sc_hd__dfxtp_4
X_1417_ _1415_/Y _1419_/C _2672_/Q _2671_/Q _2674_/Q vssd1 vssd1 vccd1 vccd1 _1420_/A
+ sky130_fd_sc_hd__a41o_4
X_2466_ _2478_/CLK _2466_/D vssd1 vssd1 vccd1 vccd1 _2199_/A sky130_fd_sc_hd__dfxtp_4
X_1279_ _1247_/Y vssd1 vssd1 vccd1 vccd1 _1279_/Y sky130_fd_sc_hd__inv_2
X_1348_ _1263_/A _1347_/X _1311_/X vssd1 vssd1 vccd1 vccd1 _1348_/X sky130_fd_sc_hd__o21a_4
X_2397_ _2397_/A _1225_/B vssd1 vssd1 vccd1 vccd1 _2397_/X sky130_fd_sc_hd__or2_4
XFILLER_36_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2320_ _2319_/Y vssd1 vssd1 vccd1 vccd1 _2320_/X sky130_fd_sc_hd__buf_2
X_2251_ _2251_/A _2251_/B vssd1 vssd1 vccd1 vccd1 _2251_/Y sky130_fd_sc_hd__nand2_4
XFILLER_65_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2182_ _1574_/X _2697_/Q _1544_/X vssd1 vssd1 vccd1 vccd1 _2182_/Y sky130_fd_sc_hd__a21oi_4
X_1202_ _1219_/A vssd1 vssd1 vccd1 vccd1 _1203_/B sky130_fd_sc_hd__buf_2
X_1966_ _1966_/A _1966_/B vssd1 vssd1 vccd1 vccd1 _1966_/Y sky130_fd_sc_hd__nor2_4
X_1897_ _1912_/A _2591_/Q vssd1 vssd1 vccd1 vccd1 _2585_/D sky130_fd_sc_hd__and2_4
X_2518_ _2670_/CLK _2077_/X vssd1 vssd1 vccd1 vccd1 _1986_/D sky130_fd_sc_hd__dfxtp_4
X_2449_ _2494_/CLK _2449_/D vssd1 vssd1 vccd1 vccd1 _1414_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_24_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1820_ _1747_/Y _1748_/Y vssd1 vssd1 vccd1 vccd1 _1820_/Y sky130_fd_sc_hd__nand2_4
XFILLER_15_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1751_ _1751_/A vssd1 vssd1 vccd1 vccd1 _1751_/Y sky130_fd_sc_hd__inv_2
X_1682_ _1681_/X vssd1 vssd1 vccd1 vccd1 _1683_/D sky130_fd_sc_hd__buf_2
X_2234_ _2671_/Q _2113_/X _1511_/X _1526_/X _1587_/X vssd1 vssd1 vccd1 vccd1 _2234_/X
+ sky130_fd_sc_hd__a2111o_4
X_2303_ _1522_/Y _2288_/Y _2291_/Y _1884_/Y _2293_/X vssd1 vssd1 vccd1 vccd1 _2303_/Y
+ sky130_fd_sc_hd__o32ai_4
X_2165_ _2165_/A _2165_/B vssd1 vssd1 vccd1 vccd1 _2165_/Y sky130_fd_sc_hd__nand2_4
X_2096_ _2096_/A vssd1 vssd1 vccd1 vccd1 _2096_/X sky130_fd_sc_hd__buf_2
XFILLER_21_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1949_ _2488_/Q vssd1 vssd1 vccd1 vccd1 _1950_/B sky130_fd_sc_hd__inv_2
XFILLER_56_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1803_ _2634_/Q _1798_/X _1802_/X vssd1 vssd1 vccd1 vccd1 _1803_/X sky130_fd_sc_hd__o21a_4
X_1596_ _1595_/Y _1587_/X vssd1 vssd1 vccd1 vccd1 _2260_/A sky130_fd_sc_hd__nor2_4
X_1665_ _2371_/A _1623_/B _1625_/C vssd1 vssd1 vccd1 vccd1 _1665_/Y sky130_fd_sc_hd__nor3_4
X_1734_ _1733_/X _1695_/X _1730_/A vssd1 vssd1 vccd1 vccd1 _1734_/X sky130_fd_sc_hd__a21o_4
XFILLER_58_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2217_ _2241_/A _2241_/B _2599_/Q _2241_/D vssd1 vssd1 vccd1 vccd1 _2217_/X sky130_fd_sc_hd__and4_4
XFILLER_38_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2079_ _2079_/A _2023_/B _2074_/Y vssd1 vssd1 vccd1 vccd1 _2079_/X sky130_fd_sc_hd__and3_4
X_2148_ _2146_/Y _2147_/Y _1463_/X vssd1 vssd1 vccd1 vccd1 _2148_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_49_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1450_ _1439_/X _1450_/B _1460_/A _1450_/D vssd1 vssd1 vccd1 vccd1 _1450_/Y sky130_fd_sc_hd__nand4_4
X_1381_ _1381_/A vssd1 vssd1 vccd1 vccd1 _1381_/X sky130_fd_sc_hd__buf_2
X_2002_ _2002_/A vssd1 vssd1 vccd1 vccd1 _2002_/Y sky130_fd_sc_hd__inv_2
XFILLER_50_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2697_ _2559_/CLK _2697_/D vssd1 vssd1 vccd1 vccd1 _2697_/Q sky130_fd_sc_hd__dfxtp_4
X_1579_ _2700_/Q _1577_/X _2187_/C vssd1 vssd1 vccd1 vccd1 _1579_/Y sky130_fd_sc_hd__nor3_4
X_1648_ _1647_/X _1755_/B _1562_/X vssd1 vssd1 vccd1 vccd1 _1648_/Y sky130_fd_sc_hd__a21oi_4
X_1717_ _1712_/X _1714_/X _1717_/C _1717_/D vssd1 vssd1 vccd1 vccd1 _1717_/Y sky130_fd_sc_hd__nand4_4
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2620_ _2621_/CLK _2620_/D vssd1 vssd1 vccd1 vccd1 _1855_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_32_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2551_ _2545_/CLK _2551_/D vssd1 vssd1 vccd1 vccd1 _2551_/Q sky130_fd_sc_hd__dfxtp_4
X_2482_ _2617_/CLK _2216_/Y vssd1 vssd1 vccd1 vccd1 _2482_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_49_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1433_ _1431_/X _1330_/B _1432_/Y vssd1 vssd1 vccd1 vccd1 _1434_/A sky130_fd_sc_hd__nand3_4
X_1502_ _2640_/Q vssd1 vssd1 vccd1 vccd1 _1726_/A sky130_fd_sc_hd__buf_2
X_1295_ _1295_/A _1305_/A _1300_/B _1268_/X vssd1 vssd1 vccd1 vccd1 _1296_/B sky130_fd_sc_hd__nand4_4
X_1364_ _1363_/Y vssd1 vssd1 vccd1 vccd1 _2685_/D sky130_fd_sc_hd__inv_2
XFILLER_11_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_2_3_0_addressalyzerBlock.SPI_CLK clkbuf_2_2_0_addressalyzerBlock.SPI_CLK/A
+ vssd1 vssd1 vccd1 vccd1 clkbuf_3_7_0_addressalyzerBlock.SPI_CLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_6_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1982_ _2528_/Q vssd1 vssd1 vccd1 vccd1 _1989_/C sky130_fd_sc_hd__inv_2
XFILLER_45_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2603_ _2621_/CLK _2603_/D vssd1 vssd1 vccd1 vccd1 _1873_/B sky130_fd_sc_hd__dfxtp_4
X_2534_ _2545_/CLK _2534_/D vssd1 vssd1 vccd1 vccd1 _2534_/Q sky130_fd_sc_hd__dfxtp_4
X_1347_ _1280_/A _1345_/X _1263_/C _1355_/C vssd1 vssd1 vccd1 vccd1 _1347_/X sky130_fd_sc_hd__and4_4
X_2396_ _2601_/Q _2602_/Q _2396_/C _2396_/D vssd1 vssd1 vccd1 vccd1 IRQ_OUT_toHost
+ sky130_fd_sc_hd__or4_4
X_1416_ _1252_/B vssd1 vssd1 vccd1 vccd1 _1419_/C sky130_fd_sc_hd__buf_2
X_2465_ _2456_/CLK _2465_/D vssd1 vssd1 vccd1 vccd1 _2223_/A sky130_fd_sc_hd__dfxtp_4
X_1278_ _1266_/C vssd1 vssd1 vccd1 vccd1 _1280_/B sky130_fd_sc_hd__buf_2
XFILLER_51_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1201_ _1201_/A vssd1 vssd1 vccd1 vccd1 _1201_/X sky130_fd_sc_hd__buf_2
XFILLER_2_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2250_ _2250_/A _2250_/B _2249_/Y vssd1 vssd1 vccd1 vccd1 _2251_/B sky130_fd_sc_hd__nand3_4
XFILLER_65_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2181_ _1653_/A _2179_/Y _2180_/X vssd1 vssd1 vccd1 vccd1 _2181_/Y sky130_fd_sc_hd__o21ai_4
X_1965_ _1974_/A _2541_/Q _2542_/Q vssd1 vssd1 vccd1 vccd1 _1971_/B sky130_fd_sc_hd__nand3_4
X_2517_ _2517_/CLK _2079_/X vssd1 vssd1 vccd1 vccd1 _1986_/C sky130_fd_sc_hd__dfxtp_4
X_1896_ _1915_/A vssd1 vssd1 vccd1 vccd1 _1912_/A sky130_fd_sc_hd__buf_2
XFILLER_0_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2379_ _2377_/Y _2378_/Y _2091_/X vssd1 vssd1 vccd1 vccd1 _2433_/D sky130_fd_sc_hd__a21oi_4
X_2448_ _2494_/CLK _2448_/D vssd1 vssd1 vccd1 vccd1 _2348_/C sky130_fd_sc_hd__dfxtp_4
XFILLER_33_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1750_ _1747_/Y _1749_/Y vssd1 vssd1 vccd1 vccd1 _2647_/D sky130_fd_sc_hd__nor2_4
X_1681_ _1707_/D _2654_/Q _1707_/A _1692_/C vssd1 vssd1 vccd1 vccd1 _1681_/X sky130_fd_sc_hd__and4_4
X_2233_ _2230_/Y _2231_/Y _2232_/Y vssd1 vssd1 vccd1 vccd1 _2233_/Y sky130_fd_sc_hd__a21oi_4
X_2164_ _2160_/Y _2162_/Y _2163_/X vssd1 vssd1 vccd1 vccd1 _2164_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_38_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2302_ _1517_/Y _2288_/Y _2291_/Y _1882_/Y _2293_/X vssd1 vssd1 vccd1 vccd1 _2473_/D
+ sky130_fd_sc_hd__o32ai_4
XFILLER_65_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2095_ _1212_/X _2084_/B _2105_/B _2514_/Q vssd1 vssd1 vccd1 vccd1 _2095_/X sky130_fd_sc_hd__and4_4
X_1879_ _1875_/X _1879_/B vssd1 vssd1 vccd1 vccd1 _1879_/Y sky130_fd_sc_hd__nor2_4
X_1948_ _1946_/A _1948_/B vssd1 vssd1 vccd1 vccd1 _1948_/Y sky130_fd_sc_hd__nor2_4
XFILLER_44_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1802_ _2635_/Q _1799_/X _1789_/X vssd1 vssd1 vccd1 vccd1 _1802_/X sky130_fd_sc_hd__o21a_4
X_1733_ _1703_/Y _1464_/X _1738_/A _1692_/C _1488_/X vssd1 vssd1 vccd1 vccd1 _1733_/X
+ sky130_fd_sc_hd__a41o_4
X_1595_ _1595_/A _1515_/A _1581_/A vssd1 vssd1 vccd1 vccd1 _1595_/Y sky130_fd_sc_hd__nand3_4
X_1664_ _1632_/A _2435_/Q _1664_/C vssd1 vssd1 vccd1 vccd1 _1664_/Y sky130_fd_sc_hd__nor3_4
XFILLER_7_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2216_ _2214_/Y _2216_/B vssd1 vssd1 vccd1 vccd1 _2216_/Y sky130_fd_sc_hd__nand2_4
XFILLER_53_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2147_ _2490_/Q _2147_/B vssd1 vssd1 vccd1 vccd1 _2147_/Y sky130_fd_sc_hd__nand2_4
X_2078_ _2074_/A _1986_/B _1986_/C vssd1 vssd1 vccd1 vccd1 _2079_/A sky130_fd_sc_hd__a21o_4
XFILLER_30_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1380_ _1254_/B _1254_/C _1254_/D vssd1 vssd1 vccd1 vccd1 _1382_/A sky130_fd_sc_hd__nor3_4
X_2001_ _2001_/A _1330_/B _2000_/Y vssd1 vssd1 vccd1 vccd1 _2002_/A sky130_fd_sc_hd__nand3_4
XFILLER_35_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2696_ _2559_/CLK _1304_/Y vssd1 vssd1 vccd1 vccd1 _2696_/Q sky130_fd_sc_hd__dfxtp_4
X_1716_ _1738_/A vssd1 vssd1 vccd1 vccd1 _1717_/D sky130_fd_sc_hd__buf_2
X_1578_ _2149_/A vssd1 vssd1 vccd1 vccd1 _2187_/C sky130_fd_sc_hd__buf_2
X_1647_ _2248_/A vssd1 vssd1 vccd1 vccd1 _1647_/X sky130_fd_sc_hd__buf_2
XFILLER_26_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2550_ _2564_/CLK _1958_/X vssd1 vssd1 vccd1 vccd1 MACRO_WR_SELECT[5] sky130_fd_sc_hd__dfxtp_4
X_2481_ _2617_/CLK _2481_/D vssd1 vssd1 vccd1 vccd1 _2481_/Q sky130_fd_sc_hd__dfxtp_4
X_1363_ _1360_/X _1361_/Y _1363_/C vssd1 vssd1 vccd1 vccd1 _1363_/Y sky130_fd_sc_hd__nand3_4
X_1501_ _2241_/B _1500_/X _1486_/Y vssd1 vssd1 vccd1 vccd1 _1501_/X sky130_fd_sc_hd__a21o_4
X_1432_ _1432_/A _1414_/B _1432_/C vssd1 vssd1 vccd1 vccd1 _1432_/Y sky130_fd_sc_hd__nand3_4
XFILLER_63_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1294_ _1290_/Y _1291_/Y _1293_/X vssd1 vssd1 vccd1 vccd1 _1294_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_23_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2679_ _2679_/CLK _2679_/D vssd1 vssd1 vccd1 vccd1 _2679_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_10_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1981_ _1981_/A vssd1 vssd1 vccd1 vccd1 _1981_/Y sky130_fd_sc_hd__inv_2
XFILLER_61_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2533_ _2564_/CLK _2533_/D vssd1 vssd1 vccd1 vccd1 _1979_/A sky130_fd_sc_hd__dfxtp_4
X_2602_ _2612_/CLK _2602_/D vssd1 vssd1 vccd1 vccd1 _2602_/Q sky130_fd_sc_hd__dfxtp_4
X_1346_ _1263_/D vssd1 vssd1 vccd1 vccd1 _1355_/C sky130_fd_sc_hd__buf_2
X_2395_ _2395_/A _2598_/Q _2599_/Q _2600_/Q vssd1 vssd1 vccd1 vccd1 _2396_/D sky130_fd_sc_hd__or4_4
X_1415_ _1414_/Y vssd1 vssd1 vccd1 vccd1 _1415_/Y sky130_fd_sc_hd__inv_2
X_2464_ _2456_/CLK _2464_/D vssd1 vssd1 vccd1 vccd1 _2249_/A sky130_fd_sc_hd__dfxtp_4
X_1277_ _1277_/A _1277_/B _1277_/C vssd1 vssd1 vccd1 vccd1 _1280_/A sky130_fd_sc_hd__nor3_4
XFILLER_51_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2180_ _1439_/X _2613_/Q _2139_/X _2149_/X vssd1 vssd1 vccd1 vccd1 _2180_/X sky130_fd_sc_hd__o22a_4
X_1200_ _1219_/A vssd1 vssd1 vccd1 vccd1 _1201_/A sky130_fd_sc_hd__inv_2
XFILLER_65_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1964_ _2375_/A _1964_/B vssd1 vssd1 vccd1 vccd1 _2544_/D sky130_fd_sc_hd__nor2_4
X_1895_ _1890_/X _1895_/B vssd1 vssd1 vccd1 vccd1 _1895_/X sky130_fd_sc_hd__and2_4
Xclkbuf_3_0_0_m1_clk_local clkbuf_2_0_0_m1_clk_local/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_1_0_m1_clk_local/A
+ sky130_fd_sc_hd__clkbuf_1
X_2516_ _2517_/CLK _2081_/X vssd1 vssd1 vccd1 vccd1 _1986_/B sky130_fd_sc_hd__dfxtp_4
X_2447_ _2493_/CLK _2350_/X vssd1 vssd1 vccd1 vccd1 _2447_/Q sky130_fd_sc_hd__dfxtp_4
X_1329_ _1313_/A _1321_/Y vssd1 vssd1 vccd1 vccd1 _1329_/Y sky130_fd_sc_hd__nand2_4
XFILLER_56_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2378_ _1240_/B _2378_/B vssd1 vssd1 vccd1 vccd1 _2378_/Y sky130_fd_sc_hd__nand2_4
XFILLER_33_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2301_ _2300_/Y _2289_/X _2292_/X _1881_/B _2294_/X vssd1 vssd1 vccd1 vccd1 _2301_/Y
+ sky130_fd_sc_hd__o32ai_4
X_1680_ _1713_/D vssd1 vssd1 vccd1 vccd1 _1692_/C sky130_fd_sc_hd__buf_2
XFILLER_65_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2232_ _1345_/X _1530_/X _1515_/A _1581_/X _2139_/X vssd1 vssd1 vccd1 vccd1 _2232_/Y
+ sky130_fd_sc_hd__a2111oi_4
X_2163_ _2241_/A _2163_/B _2602_/Q _2241_/D vssd1 vssd1 vccd1 vccd1 _2163_/X sky130_fd_sc_hd__and4_4
XFILLER_38_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2094_ _2094_/A vssd1 vssd1 vccd1 vccd1 _2105_/B sky130_fd_sc_hd__inv_2
XFILLER_0_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1878_ _2475_/Q vssd1 vssd1 vccd1 vccd1 _1879_/B sky130_fd_sc_hd__inv_2
XFILLER_21_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1947_ _1947_/A vssd1 vssd1 vccd1 vccd1 _1948_/B sky130_fd_sc_hd__inv_2
XFILLER_52_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1663_ _1602_/C _1661_/Y _1662_/Y vssd1 vssd1 vccd1 vccd1 _2657_/D sky130_fd_sc_hd__o21ai_4
X_1801_ _2635_/Q _1798_/X _1800_/X vssd1 vssd1 vccd1 vccd1 _2636_/D sky130_fd_sc_hd__o21a_4
X_1732_ _1731_/Y _1687_/B vssd1 vssd1 vccd1 vccd1 _1732_/Y sky130_fd_sc_hd__nand2_4
X_1594_ _1381_/X _1500_/X _1594_/C vssd1 vssd1 vccd1 vccd1 _1594_/Y sky130_fd_sc_hd__nor3_4
X_2215_ _2239_/A _2482_/Q vssd1 vssd1 vccd1 vccd1 _2216_/B sky130_fd_sc_hd__nand2_4
XFILLER_53_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2077_ _2076_/X _2023_/B _2067_/B vssd1 vssd1 vccd1 vccd1 _2077_/X sky130_fd_sc_hd__and3_4
X_2146_ _1647_/X _1752_/A _1562_/X vssd1 vssd1 vccd1 vccd1 _2146_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_34_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2000_ _2000_/A _2000_/B _2536_/Q CLK_LED vssd1 vssd1 vccd1 vccd1 _2000_/Y sky130_fd_sc_hd__nand4_4
XFILLER_50_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_3_3_0_addressalyzerBlock.SPI_CLK clkbuf_3_3_0_addressalyzerBlock.SPI_CLK/A
+ vssd1 vssd1 vccd1 vccd1 clkbuf_4_7_0_addressalyzerBlock.SPI_CLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_16_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2695_ _2695_/CLK _2695_/D vssd1 vssd1 vccd1 vccd1 _2695_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_4_9_0_m1_clk_local clkbuf_4_9_0_m1_clk_local/A vssd1 vssd1 vccd1 vccd1 _2564_/CLK
+ sky130_fd_sc_hd__clkbuf_1
X_1715_ _1715_/A vssd1 vssd1 vccd1 vccd1 _1717_/C sky130_fd_sc_hd__buf_2
X_1646_ _2493_/Q vssd1 vssd1 vccd1 vccd1 _2248_/A sky130_fd_sc_hd__inv_2
X_1577_ _1577_/A vssd1 vssd1 vccd1 vccd1 _1577_/X sky130_fd_sc_hd__buf_2
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2129_ _1815_/X _1633_/A _1784_/X vssd1 vssd1 vccd1 vccd1 _2129_/Y sky130_fd_sc_hd__nand3_4
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2480_ _2705_/CLK _2480_/D vssd1 vssd1 vccd1 vccd1 _2263_/B sky130_fd_sc_hd__dfxtp_4
X_1500_ _1500_/A vssd1 vssd1 vccd1 vccd1 _1500_/X sky130_fd_sc_hd__buf_2
XFILLER_9_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1293_ _1293_/A vssd1 vssd1 vccd1 vccd1 _1293_/X sky130_fd_sc_hd__buf_2
X_1362_ _1274_/X vssd1 vssd1 vccd1 vccd1 _1363_/C sky130_fd_sc_hd__buf_2
X_1431_ _1414_/A _1432_/C _1414_/B vssd1 vssd1 vccd1 vccd1 _1431_/X sky130_fd_sc_hd__a21o_4
XFILLER_51_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2678_ _2527_/CLK _1404_/Y vssd1 vssd1 vccd1 vccd1 _1255_/A sky130_fd_sc_hd__dfxtp_4
X_1629_ _1626_/A vssd1 vssd1 vccd1 vccd1 _2353_/D sky130_fd_sc_hd__buf_2
XFILLER_36_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1980_ _1980_/A vssd1 vssd1 vccd1 vccd1 _1989_/A sky130_fd_sc_hd__inv_2
XFILLER_9_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2532_ _2564_/CLK _2023_/X vssd1 vssd1 vccd1 vccd1 _2532_/Q sky130_fd_sc_hd__dfxtp_4
X_2601_ _2612_/CLK _1868_/X vssd1 vssd1 vccd1 vccd1 _2601_/Q sky130_fd_sc_hd__dfxtp_4
X_2463_ _2456_/CLK _2463_/D vssd1 vssd1 vccd1 vccd1 _2463_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_9_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1276_ _2696_/Q vssd1 vssd1 vccd1 vccd1 _1276_/Y sky130_fd_sc_hd__inv_2
X_1345_ _2687_/Q vssd1 vssd1 vccd1 vccd1 _1345_/X sky130_fd_sc_hd__buf_2
X_2394_ _2393_/A _2392_/Y _2393_/Y vssd1 vssd1 vccd1 vccd1 MISO_toHost sky130_fd_sc_hd__a21oi_4
X_1414_ _1414_/A _1414_/B _1414_/C vssd1 vssd1 vccd1 vccd1 _1414_/Y sky130_fd_sc_hd__nand3_4
XPHY_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1963_ _1283_/B _2551_/Q vssd1 vssd1 vccd1 vccd1 _1963_/X sky130_fd_sc_hd__and2_4
X_1894_ _1890_/X _1894_/B vssd1 vssd1 vccd1 vccd1 _2587_/D sky130_fd_sc_hd__and2_4
X_2515_ _2670_/CLK _2082_/Y vssd1 vssd1 vccd1 vccd1 _2515_/Q sky130_fd_sc_hd__dfxtp_4
X_2446_ _2443_/CLK _2355_/X vssd1 vssd1 vccd1 vccd1 _2446_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_56_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1328_ _1274_/X vssd1 vssd1 vccd1 vccd1 _1330_/B sky130_fd_sc_hd__buf_2
X_1259_ _1381_/A _1259_/B _1256_/Y _1384_/D vssd1 vssd1 vccd1 vccd1 _1277_/C sky130_fd_sc_hd__nand4_4
X_2377_ _1608_/Y vssd1 vssd1 vccd1 vccd1 _2377_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2231_ _1574_/A _2695_/Q _1544_/A vssd1 vssd1 vccd1 vccd1 _2231_/Y sky130_fd_sc_hd__a21oi_4
X_2300_ _1726_/A vssd1 vssd1 vccd1 vccd1 _2300_/Y sky130_fd_sc_hd__inv_2
XFILLER_65_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2162_ _2162_/A vssd1 vssd1 vccd1 vccd1 _2162_/Y sky130_fd_sc_hd__inv_2
X_2093_ _2091_/X _2094_/A _2514_/Q _2084_/B vssd1 vssd1 vccd1 vccd1 _2507_/D sky130_fd_sc_hd__nor4_4
XFILLER_17_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1946_ _1946_/A _1945_/Y vssd1 vssd1 vccd1 vccd1 _1946_/Y sky130_fd_sc_hd__nor2_4
X_1877_ _1875_/X _1877_/B vssd1 vssd1 vccd1 vccd1 _2596_/D sky130_fd_sc_hd__nor2_4
X_2429_ _2508_/CLK _2383_/X vssd1 vssd1 vccd1 vccd1 _2429_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_56_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1800_ _2636_/Q _1799_/X _1789_/X vssd1 vssd1 vccd1 vccd1 _1800_/X sky130_fd_sc_hd__o21a_4
XPHY_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1662_ _2165_/A _1662_/B vssd1 vssd1 vccd1 vccd1 _1662_/Y sky130_fd_sc_hd__nand2_4
XFILLER_7_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1731_ _1517_/Y _1674_/X _1730_/Y vssd1 vssd1 vccd1 vccd1 _1731_/Y sky130_fd_sc_hd__o21ai_4
X_2214_ _2192_/X _2213_/Y _2189_/X vssd1 vssd1 vccd1 vccd1 _2214_/Y sky130_fd_sc_hd__o21ai_4
X_1593_ _1500_/X _2187_/B _2684_/Q _1592_/X vssd1 vssd1 vccd1 vccd1 _1593_/Y sky130_fd_sc_hd__a2bb2oi_4
X_2076_ _1986_/D _2075_/Y vssd1 vssd1 vccd1 vccd1 _2076_/X sky130_fd_sc_hd__or2_4
X_2145_ _2142_/X _2144_/X _2495_/Q vssd1 vssd1 vccd1 vccd1 _2145_/X sky130_fd_sc_hd__a21o_4
XFILLER_19_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1929_ _2223_/A vssd1 vssd1 vccd1 vccd1 _1929_/Y sky130_fd_sc_hd__inv_2
XFILLER_39_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2694_ _2693_/CLK _2694_/D vssd1 vssd1 vccd1 vccd1 _1248_/A sky130_fd_sc_hd__dfxtp_4
X_1576_ _1573_/A vssd1 vssd1 vccd1 vccd1 _1577_/A sky130_fd_sc_hd__buf_2
X_1714_ _1714_/A vssd1 vssd1 vccd1 vccd1 _1714_/X sky130_fd_sc_hd__buf_2
X_1645_ _1640_/X _1644_/X _2495_/Q vssd1 vssd1 vccd1 vccd1 _1651_/A sky130_fd_sc_hd__a21o_4
XFILLER_54_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2059_ _2053_/X _2055_/Y _2057_/B _2057_/C _1293_/X vssd1 vssd1 vccd1 vccd1 _2059_/Y
+ sky130_fd_sc_hd__a41oi_4
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2128_ _2123_/X _2124_/X _2125_/Y _1945_/Y _2127_/X vssd1 vssd1 vccd1 vccd1 _2128_/Y
+ sky130_fd_sc_hd__o32ai_4
XFILLER_26_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1430_ _1429_/X _2005_/B _1254_/D vssd1 vssd1 vccd1 vccd1 _2671_/D sky130_fd_sc_hd__and3_4
XFILLER_31_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1361_ _1350_/Y vssd1 vssd1 vccd1 vccd1 _1361_/Y sky130_fd_sc_hd__inv_2
XFILLER_48_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1292_ _1273_/A vssd1 vssd1 vccd1 vccd1 _1293_/A sky130_fd_sc_hd__buf_2
XFILLER_63_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2677_ _2527_/CLK _1407_/Y vssd1 vssd1 vccd1 vccd1 _1255_/B sky130_fd_sc_hd__dfxtp_4
X_1628_ _1623_/Y _1625_/Y _1627_/X vssd1 vssd1 vccd1 vccd1 _1628_/Y sky130_fd_sc_hd__o21ai_4
X_1559_ _1559_/A vssd1 vssd1 vccd1 vccd1 _1559_/X sky130_fd_sc_hd__buf_2
XFILLER_52_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2600_ _2621_/CLK _1869_/X vssd1 vssd1 vccd1 vccd1 _2600_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_9_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2531_ _2564_/CLK _2029_/X vssd1 vssd1 vccd1 vccd1 _2531_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_47_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2393_ _2393_/A MISO_fromClient vssd1 vssd1 vccd1 vccd1 _2393_/Y sky130_fd_sc_hd__nor2_4
X_1413_ _1413_/A vssd1 vssd1 vccd1 vccd1 _1414_/B sky130_fd_sc_hd__buf_2
X_2462_ _2456_/CLK _2462_/D vssd1 vssd1 vccd1 vccd1 _2462_/Q sky130_fd_sc_hd__dfxtp_4
X_1344_ _1343_/Y vssd1 vssd1 vccd1 vccd1 _1344_/Y sky130_fd_sc_hd__inv_2
X_1275_ _1274_/X vssd1 vssd1 vccd1 vccd1 _1283_/B sky130_fd_sc_hd__buf_2
XFILLER_36_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1962_ _1961_/A _2552_/Q vssd1 vssd1 vccd1 vccd1 _1962_/X sky130_fd_sc_hd__and2_4
X_1893_ _1890_/X _2594_/Q vssd1 vssd1 vccd1 vccd1 _2588_/D sky130_fd_sc_hd__and2_4
X_2376_ _1240_/B _2365_/B _2096_/X _1665_/Y vssd1 vssd1 vccd1 vccd1 _2376_/X sky130_fd_sc_hd__a211o_4
X_2514_ _2514_/CLK _2514_/D vssd1 vssd1 vccd1 vccd1 _2514_/Q sky130_fd_sc_hd__dfxtp_4
X_2445_ _2443_/CLK _2358_/Y vssd1 vssd1 vccd1 vccd1 _1755_/B sky130_fd_sc_hd__dfxtp_4
X_1327_ _1327_/A vssd1 vssd1 vccd1 vccd1 _1330_/A sky130_fd_sc_hd__inv_2
XFILLER_56_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1258_ _1257_/Y vssd1 vssd1 vccd1 vccd1 _1384_/D sky130_fd_sc_hd__inv_2
XPHY_207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2230_ _1653_/A _2228_/Y _2229_/X vssd1 vssd1 vccd1 vccd1 _2230_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_46_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2161_ _1600_/B vssd1 vssd1 vccd1 vccd1 _2162_/A sky130_fd_sc_hd__buf_2
XFILLER_38_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2092_ _2091_/X _2499_/Q _2104_/B vssd1 vssd1 vccd1 vccd1 _2508_/D sky130_fd_sc_hd__nor3_4
XFILLER_0_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1945_ _2490_/Q vssd1 vssd1 vccd1 vccd1 _1945_/Y sky130_fd_sc_hd__inv_2
X_1876_ _2476_/Q vssd1 vssd1 vccd1 vccd1 _1877_/B sky130_fd_sc_hd__inv_2
XFILLER_29_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2428_ _2494_/CLK _2427_/Q vssd1 vssd1 vccd1 vccd1 _2331_/A sky130_fd_sc_hd__dfxtp_4
X_2359_ _1753_/B _2352_/X _1481_/X _2354_/X vssd1 vssd1 vccd1 vccd1 _2444_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_52_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_4_3_0_addressalyzerBlock.SPI_CLK clkbuf_4_2_0_addressalyzerBlock.SPI_CLK/A
+ vssd1 vssd1 vccd1 vccd1 _2493_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1661_ _1658_/Y _1659_/Y _1660_/Y vssd1 vssd1 vccd1 vccd1 _1661_/Y sky130_fd_sc_hd__a21oi_4
X_1592_ _1591_/Y vssd1 vssd1 vccd1 vccd1 _1592_/X sky130_fd_sc_hd__buf_2
XFILLER_11_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1730_ _1730_/A _1714_/X _1717_/D _1448_/Y vssd1 vssd1 vccd1 vccd1 _1730_/Y sky130_fd_sc_hd__nand4_4
X_2213_ _2211_/Y _2212_/Y _2162_/A vssd1 vssd1 vccd1 vccd1 _2213_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_38_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2144_ _1922_/A _1546_/X _2221_/B _2143_/Y vssd1 vssd1 vccd1 vccd1 _2144_/X sky130_fd_sc_hd__a211o_4
XFILLER_34_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2075_ _2074_/Y vssd1 vssd1 vccd1 vccd1 _2075_/Y sky130_fd_sc_hd__inv_2
XFILLER_26_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1859_ _1858_/A DATA_AVAILABLE[5] vssd1 vssd1 vccd1 vccd1 _1859_/X sky130_fd_sc_hd__and2_4
X_1928_ _1930_/A _1928_/B vssd1 vssd1 vccd1 vccd1 _1928_/Y sky130_fd_sc_hd__nor2_4
Xclkbuf_2_2_0_m1_clk_local clkbuf_2_3_0_m1_clk_local/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_4_0_m1_clk_local/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_39_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1713_ _1450_/B _1652_/A _1460_/A _1713_/D vssd1 vssd1 vccd1 vccd1 _1714_/A sky130_fd_sc_hd__and4_4
X_2693_ _2693_/CLK _1320_/Y vssd1 vssd1 vccd1 vccd1 _1248_/B sky130_fd_sc_hd__dfxtp_4
X_1575_ _1574_/X vssd1 vssd1 vccd1 vccd1 _1575_/Y sky130_fd_sc_hd__inv_2
X_1644_ _2469_/Q _2272_/A _2494_/Q _1643_/Y vssd1 vssd1 vccd1 vccd1 _1644_/X sky130_fd_sc_hd__a211o_4
XFILLER_58_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2127_ _2126_/Y vssd1 vssd1 vccd1 vccd1 _2127_/X sky130_fd_sc_hd__buf_2
XFILLER_26_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2058_ _2058_/A _2056_/Y _2058_/C vssd1 vssd1 vccd1 vccd1 _2524_/D sky130_fd_sc_hd__nor3_4
XFILLER_34_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1360_ _1355_/A _1338_/X _1355_/C vssd1 vssd1 vccd1 vccd1 _1360_/X sky130_fd_sc_hd__a21o_4
X_1291_ _1295_/A vssd1 vssd1 vccd1 vccd1 _1291_/Y sky130_fd_sc_hd__inv_2
XFILLER_63_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2676_ _2679_/CLK _1410_/X vssd1 vssd1 vccd1 vccd1 _1381_/A sky130_fd_sc_hd__dfxtp_4
X_1627_ _1626_/Y _1450_/D _1768_/B _1667_/B vssd1 vssd1 vccd1 vccd1 _1627_/X sky130_fd_sc_hd__a2bb2o_4
X_1489_ _1489_/A vssd1 vssd1 vccd1 vccd1 _1489_/Y sky130_fd_sc_hd__inv_2
X_1558_ _2495_/Q vssd1 vssd1 vccd1 vccd1 _1559_/A sky130_fd_sc_hd__inv_2
XFILLER_54_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_5_0_m1_clk_local clkbuf_4_5_0_m1_clk_local/A vssd1 vssd1 vccd1 vccd1 _2420_/CLK
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_10_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2530_ _2564_/CLK _2034_/Y vssd1 vssd1 vccd1 vccd1 _1990_/B sky130_fd_sc_hd__dfxtp_4
XFILLER_13_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1343_ _1332_/X _1340_/Y _1342_/Y vssd1 vssd1 vccd1 vccd1 _1343_/Y sky130_fd_sc_hd__o21ai_4
X_2392_ _2392_/A vssd1 vssd1 vccd1 vccd1 _2392_/Y sky130_fd_sc_hd__inv_2
X_1412_ _2014_/A _1401_/X _1412_/C vssd1 vssd1 vccd1 vccd1 _1412_/Y sky130_fd_sc_hd__nor3_4
X_2461_ _2456_/CLK _2461_/D vssd1 vssd1 vccd1 vccd1 _1638_/A sky130_fd_sc_hd__dfxtp_4
X_1274_ _1378_/A vssd1 vssd1 vccd1 vccd1 _1274_/X sky130_fd_sc_hd__buf_2
XFILLER_36_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2659_ _2655_/CLK _2659_/D vssd1 vssd1 vccd1 vccd1 _2659_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_63_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1892_ _1890_/X _2595_/Q vssd1 vssd1 vccd1 vccd1 _1892_/X sky130_fd_sc_hd__and2_4
X_1961_ _1961_/A _2553_/Q vssd1 vssd1 vccd1 vccd1 _1961_/X sky130_fd_sc_hd__and2_4
X_2513_ _2655_/CLK _2085_/X vssd1 vssd1 vccd1 vccd1 _2513_/Q sky130_fd_sc_hd__dfxtp_4
X_1326_ _1325_/Y vssd1 vssd1 vccd1 vccd1 _2692_/D sky130_fd_sc_hd__inv_2
XFILLER_56_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2375_ _2375_/A _2375_/B vssd1 vssd1 vccd1 vccd1 _2375_/Y sky130_fd_sc_hd__nor2_4
X_2444_ _2495_/CLK _2444_/D vssd1 vssd1 vccd1 vccd1 _1752_/A sky130_fd_sc_hd__dfxtp_4
X_1257_ _1257_/A _2679_/Q vssd1 vssd1 vccd1 vccd1 _1257_/Y sky130_fd_sc_hd__nand2_4
XFILLER_24_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XINSDIODE2_0 DATA_AVAILABLE[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2160_ _2156_/Y _2159_/X vssd1 vssd1 vccd1 vccd1 _2160_/Y sky130_fd_sc_hd__nand2_4
XFILLER_2_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2091_ _2096_/A vssd1 vssd1 vccd1 vccd1 _2091_/X sky130_fd_sc_hd__buf_2
X_1875_ _1875_/A vssd1 vssd1 vccd1 vccd1 _1875_/X sky130_fd_sc_hd__buf_2
X_1944_ _1875_/A vssd1 vssd1 vccd1 vccd1 _1946_/A sky130_fd_sc_hd__buf_2
X_2427_ _2494_/CLK _2425_/Q vssd1 vssd1 vccd1 vccd1 _2427_/Q sky130_fd_sc_hd__dfxtp_4
X_1309_ _1248_/B vssd1 vssd1 vccd1 vccd1 _1318_/B sky130_fd_sc_hd__inv_2
XFILLER_29_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2289_ _2288_/Y vssd1 vssd1 vccd1 vccd1 _2289_/X sky130_fd_sc_hd__buf_2
X_2358_ _2296_/Y _2357_/A _2357_/Y vssd1 vssd1 vccd1 vccd1 _2358_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_52_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1591_ _1591_/A _1583_/A vssd1 vssd1 vccd1 vccd1 _1591_/Y sky130_fd_sc_hd__nor2_4
X_1660_ _1254_/A _1531_/X _1512_/X _1527_/X _2187_/B vssd1 vssd1 vccd1 vccd1 _1660_/Y
+ sky130_fd_sc_hd__a2111oi_4
X_2212_ _2260_/A THREAD_COUNT[3] vssd1 vssd1 vccd1 vccd1 _2212_/Y sky130_fd_sc_hd__nand2_4
X_2143_ _2143_/A _1877_/B vssd1 vssd1 vccd1 vccd1 _2143_/Y sky130_fd_sc_hd__nor2_4
XFILLER_46_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2074_ _2074_/A _1986_/B _1986_/C vssd1 vssd1 vccd1 vccd1 _2074_/Y sky130_fd_sc_hd__nand3_4
X_1858_ _1858_/A _1858_/B vssd1 vssd1 vccd1 vccd1 _2609_/D sky130_fd_sc_hd__and2_4
X_1927_ _2199_/A vssd1 vssd1 vccd1 vccd1 _1928_/B sky130_fd_sc_hd__inv_2
XFILLER_1_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1789_ _1776_/X vssd1 vssd1 vccd1 vccd1 _1789_/X sky130_fd_sc_hd__buf_2
XFILLER_55_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2692_ _2559_/CLK _2692_/D vssd1 vssd1 vccd1 vccd1 _1247_/A sky130_fd_sc_hd__dfxtp_4
XPHY_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1712_ _2651_/Q vssd1 vssd1 vccd1 vccd1 _1712_/X sky130_fd_sc_hd__buf_2
XFILLER_6_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1643_ _2220_/B _1643_/B vssd1 vssd1 vccd1 vccd1 _1643_/Y sky130_fd_sc_hd__nor2_4
X_1574_ _1574_/A vssd1 vssd1 vccd1 vccd1 _1574_/X sky130_fd_sc_hd__buf_2
Xclkbuf_4_13_0_m1_clk_local clkbuf_3_6_0_m1_clk_local/X vssd1 vssd1 vccd1 vccd1 _2559_/CLK
+ sky130_fd_sc_hd__clkbuf_1
X_2057_ _2057_/A _2057_/B _2057_/C _1988_/C vssd1 vssd1 vccd1 vccd1 _2058_/C sky130_fd_sc_hd__and4_4
X_2126_ _2114_/Y _1776_/X vssd1 vssd1 vccd1 vccd1 _2126_/Y sky130_fd_sc_hd__nand2_4
XFILLER_26_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1290_ _1300_/B _1285_/Y _2696_/Q _2695_/Q vssd1 vssd1 vccd1 vccd1 _1290_/Y sky130_fd_sc_hd__nand4_4
XFILLER_0_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1626_ _1626_/A vssd1 vssd1 vccd1 vccd1 _1626_/Y sky130_fd_sc_hd__inv_2
X_2675_ _2679_/CLK _1412_/Y vssd1 vssd1 vccd1 vccd1 _1382_/C sky130_fd_sc_hd__dfxtp_4
XFILLER_39_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1488_ _1478_/A vssd1 vssd1 vccd1 vccd1 _1488_/X sky130_fd_sc_hd__buf_2
X_1557_ _1552_/X _1556_/X vssd1 vssd1 vccd1 vccd1 _1557_/Y sky130_fd_sc_hd__nand2_4
X_2109_ _1521_/X _1524_/X _1528_/X vssd1 vssd1 vccd1 vccd1 _2494_/D sky130_fd_sc_hd__a21oi_4
XFILLER_27_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2460_ _2456_/CLK _2460_/D vssd1 vssd1 vccd1 vccd1 _2460_/Q sky130_fd_sc_hd__dfxtp_4
X_1342_ _1332_/X _1355_/A _1338_/X _1280_/B _1293_/A vssd1 vssd1 vccd1 vccd1 _1342_/Y
+ sky130_fd_sc_hd__a41oi_4
X_1411_ _1382_/C _1382_/A vssd1 vssd1 vccd1 vccd1 _1412_/C sky130_fd_sc_hd__nor2_4
X_1273_ _1273_/A vssd1 vssd1 vccd1 vccd1 _1378_/A sky130_fd_sc_hd__inv_2
X_2391_ _1836_/A S1_CLK_SELECT _2390_/Y vssd1 vssd1 vccd1 vccd1 _2391_/X sky130_fd_sc_hd__o21a_4
XFILLER_51_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2589_ _2559_/CLK _1892_/X vssd1 vssd1 vccd1 vccd1 HASH_ADDR[4] sky130_fd_sc_hd__dfxtp_4
X_2658_ _2438_/CLK _2658_/D vssd1 vssd1 vccd1 vccd1 _1626_/A sky130_fd_sc_hd__dfxtp_4
X_1609_ _1240_/B _2382_/C vssd1 vssd1 vccd1 vccd1 _1609_/Y sky130_fd_sc_hd__nor2_4
XFILLER_47_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1891_ _1890_/X _1891_/B vssd1 vssd1 vccd1 vccd1 _1891_/X sky130_fd_sc_hd__and2_4
X_1960_ _1961_/A _1960_/B vssd1 vssd1 vccd1 vccd1 _2548_/D sky130_fd_sc_hd__and2_4
XFILLER_21_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2512_ _2612_/CLK _2086_/X vssd1 vssd1 vccd1 vccd1 _2396_/C sky130_fd_sc_hd__dfxtp_4
X_2443_ _2443_/CLK _2360_/X vssd1 vssd1 vccd1 vccd1 _2443_/Q sky130_fd_sc_hd__dfxtp_4
X_1325_ _1323_/X _1324_/Y vssd1 vssd1 vccd1 vccd1 _1325_/Y sky130_fd_sc_hd__nand2_4
X_1256_ _1255_/Y vssd1 vssd1 vccd1 vccd1 _1256_/Y sky130_fd_sc_hd__inv_2
X_2374_ _1828_/A _2429_/Q _1209_/X _2378_/B vssd1 vssd1 vccd1 vccd1 _2375_/B sky130_fd_sc_hd__a22oi_4
XPHY_209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_1 DATA_FROM_HASH[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_8_0_addressalyzerBlock.SPI_CLK clkbuf_4_9_0_addressalyzerBlock.SPI_CLK/A
+ vssd1 vssd1 vccd1 vccd1 _2612_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_30_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2090_ _1212_/X _2104_/B _2499_/Q vssd1 vssd1 vccd1 vccd1 _2509_/D sky130_fd_sc_hd__and3_4
XFILLER_2_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1874_ _1293_/A vssd1 vssd1 vccd1 vccd1 _1875_/A sky130_fd_sc_hd__buf_2
X_1943_ _1941_/A _2565_/Q vssd1 vssd1 vccd1 vccd1 _2557_/D sky130_fd_sc_hd__and2_4
XFILLER_9_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2426_ _2670_/CLK _2385_/Y vssd1 vssd1 vccd1 vccd1 _2407_/D sky130_fd_sc_hd__dfxtp_4
X_1308_ _1307_/Y vssd1 vssd1 vccd1 vccd1 _2695_/D sky130_fd_sc_hd__inv_2
XFILLER_44_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1239_ _1618_/A vssd1 vssd1 vccd1 vccd1 _1240_/B sky130_fd_sc_hd__buf_2
X_2288_ _2287_/Y vssd1 vssd1 vccd1 vccd1 _2288_/Y sky130_fd_sc_hd__inv_2
X_2357_ _2357_/A _2369_/B _1755_/B vssd1 vssd1 vccd1 vccd1 _2357_/Y sky130_fd_sc_hd__nand3_4
XFILLER_60_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1590_ _1590_/A vssd1 vssd1 vccd1 vccd1 _1591_/A sky130_fd_sc_hd__inv_2
X_2211_ _2193_/X _2209_/Y _2210_/X vssd1 vssd1 vccd1 vccd1 _2211_/Y sky130_fd_sc_hd__o21ai_4
X_2073_ _2515_/Q vssd1 vssd1 vccd1 vccd1 _2074_/A sky130_fd_sc_hd__buf_2
X_2142_ ID_toHost _1546_/X _1548_/X _2141_/Y vssd1 vssd1 vccd1 vccd1 _2142_/X sky130_fd_sc_hd__a211o_4
X_1857_ _1858_/A _1857_/B vssd1 vssd1 vccd1 vccd1 _1857_/X sky130_fd_sc_hd__and2_4
X_1788_ _1774_/A _2632_/Q _1787_/X vssd1 vssd1 vccd1 vccd1 _2640_/D sky130_fd_sc_hd__o21a_4
X_1926_ _1930_/A _1926_/B vssd1 vssd1 vccd1 vccd1 _2569_/D sky130_fd_sc_hd__nor2_4
XFILLER_29_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2409_ _2413_/CLK _2408_/Q vssd1 vssd1 vccd1 vccd1 _1833_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_40_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2691_ _2559_/CLK _2691_/D vssd1 vssd1 vccd1 vccd1 _1247_/B sky130_fd_sc_hd__dfxtp_4
XPHY_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1642_ _2477_/Q vssd1 vssd1 vccd1 vccd1 _1643_/B sky130_fd_sc_hd__inv_2
X_1711_ _1701_/Y _1709_/Y _1710_/X vssd1 vssd1 vccd1 vccd1 _1711_/X sky130_fd_sc_hd__o21a_4
X_1573_ _1573_/A _2149_/A vssd1 vssd1 vccd1 vccd1 _1574_/A sky130_fd_sc_hd__nor2_4
XFILLER_66_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2056_ _2053_/X _2055_/Y _2057_/B _2057_/C _1988_/C vssd1 vssd1 vccd1 vccd1 _2056_/Y
+ sky130_fd_sc_hd__a41oi_4
X_2125_ _1815_/X _1633_/A _1481_/X vssd1 vssd1 vccd1 vccd1 _2125_/Y sky130_fd_sc_hd__nand3_4
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1909_ _1909_/A vssd1 vssd1 vccd1 vccd1 _1910_/B sky130_fd_sc_hd__inv_2
XFILLER_22_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1625_ _1632_/A _1664_/C _1625_/C vssd1 vssd1 vccd1 vccd1 _1625_/Y sky130_fd_sc_hd__nor3_4
X_2674_ _2679_/CLK _1421_/Y vssd1 vssd1 vccd1 vccd1 _2674_/Q sky130_fd_sc_hd__dfxtp_4
X_1556_ _2470_/Q _1546_/X _2221_/B _1555_/Y vssd1 vssd1 vccd1 vccd1 _1556_/X sky130_fd_sc_hd__a211o_4
X_1487_ _1485_/Y _1486_/Y _1444_/B vssd1 vssd1 vccd1 vccd1 _1487_/X sky130_fd_sc_hd__a21o_4
XFILLER_54_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2039_ _2039_/A _2023_/B _2039_/C vssd1 vssd1 vccd1 vccd1 _2039_/X sky130_fd_sc_hd__and3_4
X_2108_ _1513_/X _1519_/X _2091_/X vssd1 vssd1 vccd1 vccd1 _2495_/D sky130_fd_sc_hd__a21oi_4
XFILLER_6_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1410_ _1396_/X _1401_/X _1409_/Y vssd1 vssd1 vccd1 vccd1 _1410_/X sky130_fd_sc_hd__o21a_4
XFILLER_5_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1272_ _1305_/A _1282_/C _1268_/X _1282_/D _2700_/Q vssd1 vssd1 vccd1 vccd1 _1272_/X
+ sky130_fd_sc_hd__a41o_4
X_1341_ _1266_/A vssd1 vssd1 vccd1 vccd1 _1355_/A sky130_fd_sc_hd__buf_2
XFILLER_3_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2390_ _2389_/Y S1_CLK_SELECT vssd1 vssd1 vccd1 vccd1 _2390_/Y sky130_fd_sc_hd__nand2_4
XFILLER_51_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2657_ _2612_/CLK _2657_/D vssd1 vssd1 vccd1 vccd1 _1662_/B sky130_fd_sc_hd__dfxtp_4
X_1539_ _1539_/A vssd1 vssd1 vccd1 vccd1 _1539_/Y sky130_fd_sc_hd__inv_2
X_1608_ _1240_/B _1608_/B vssd1 vssd1 vccd1 vccd1 _1608_/Y sky130_fd_sc_hd__nor2_4
X_2588_ _2517_/CLK _2588_/D vssd1 vssd1 vccd1 vccd1 HASH_ADDR[3] sky130_fd_sc_hd__dfxtp_4
XFILLER_47_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_1_0_m1_clk_local clkbuf_4_1_0_m1_clk_local/A vssd1 vssd1 vccd1 vccd1 _2581_/CLK
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_58_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1890_ _1915_/A vssd1 vssd1 vccd1 vccd1 _1890_/X sky130_fd_sc_hd__buf_2
XFILLER_45_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2373_ _2096_/X _1235_/X _2381_/C _2371_/Y _2372_/X vssd1 vssd1 vccd1 vccd1 _2373_/Y
+ sky130_fd_sc_hd__o32ai_4
XFILLER_5_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2511_ _2511_/CLK _2087_/X vssd1 vssd1 vccd1 vccd1 _2511_/Q sky130_fd_sc_hd__dfxtp_4
X_2442_ _2495_/CLK _2361_/X vssd1 vssd1 vccd1 vccd1 _2442_/Q sky130_fd_sc_hd__dfxtp_4
X_1324_ _1313_/Y _1247_/A _1247_/B vssd1 vssd1 vccd1 vccd1 _1324_/Y sky130_fd_sc_hd__nand3_4
XFILLER_56_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1255_ _1255_/A _1255_/B vssd1 vssd1 vccd1 vccd1 _1255_/Y sky130_fd_sc_hd__nand2_4
Xclkbuf_4_13_0_addressalyzerBlock.SPI_CLK clkbuf_3_6_0_addressalyzerBlock.SPI_CLK/X
+ vssd1 vssd1 vccd1 vccd1 _2508_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_24_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_2 DATA_FROM_HASH[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_3_7_0_m1_clk_local clkbuf_3_7_0_m1_clk_local/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_7_0_m1_clk_local/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_23_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1942_ _1941_/A _1942_/B vssd1 vssd1 vccd1 vccd1 _1942_/X sky130_fd_sc_hd__and2_4
XFILLER_21_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1873_ _1873_/A _1873_/B vssd1 vssd1 vccd1 vccd1 _2597_/D sky130_fd_sc_hd__and2_4
XFILLER_9_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2425_ _2670_/CLK _2424_/Q vssd1 vssd1 vccd1 vccd1 _2425_/Q sky130_fd_sc_hd__dfxtp_4
X_2356_ _2353_/X vssd1 vssd1 vccd1 vccd1 _2357_/A sky130_fd_sc_hd__inv_2
X_1307_ _1305_/Y _1283_/B _1306_/Y vssd1 vssd1 vccd1 vccd1 _1307_/Y sky130_fd_sc_hd__nand3_4
XFILLER_56_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1238_ _1201_/X _1209_/X _1238_/C vssd1 vssd1 vccd1 vccd1 _1238_/Y sky130_fd_sc_hd__nand3_4
XFILLER_37_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2287_ _1242_/A _1626_/Y vssd1 vssd1 vccd1 vccd1 _2287_/Y sky130_fd_sc_hd__nor2_4
XFILLER_60_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2210_ _2672_/Q _2113_/X _1511_/X _1526_/X _2154_/X vssd1 vssd1 vccd1 vccd1 _2210_/X
+ sky130_fd_sc_hd__a2111o_4
XFILLER_53_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2072_ _2066_/Y _2067_/B _2071_/Y vssd1 vssd1 vccd1 vccd1 _2072_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_34_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2141_ _2143_/A _2141_/B vssd1 vssd1 vccd1 vccd1 _2141_/Y sky130_fd_sc_hd__nor2_4
XFILLER_19_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1925_ _1925_/A vssd1 vssd1 vccd1 vccd1 _1926_/B sky130_fd_sc_hd__inv_2
X_1856_ _1858_/A _1856_/B vssd1 vssd1 vccd1 vccd1 _2611_/D sky130_fd_sc_hd__and2_4
X_1787_ _1775_/X _2640_/Q _1777_/X vssd1 vssd1 vccd1 vccd1 _1787_/X sky130_fd_sc_hd__o21a_4
XFILLER_57_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2408_ _2517_/CLK _1273_/A vssd1 vssd1 vccd1 vccd1 _2408_/Q sky130_fd_sc_hd__dfxtp_4
X_2339_ _2334_/X _2117_/X ID_toHost vssd1 vssd1 vccd1 vccd1 _2339_/Y sky130_fd_sc_hd__nand3_4
XFILLER_40_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2690_ _2559_/CLK _1337_/Y vssd1 vssd1 vccd1 vccd1 _1264_/A sky130_fd_sc_hd__dfxtp_4
X_1572_ _1572_/A vssd1 vssd1 vccd1 vccd1 _2149_/A sky130_fd_sc_hd__inv_2
XFILLER_6_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1710_ _1707_/A _1695_/X _1697_/X vssd1 vssd1 vccd1 vccd1 _1710_/X sky130_fd_sc_hd__o21a_4
X_1641_ _2493_/Q vssd1 vssd1 vccd1 vccd1 _2220_/B sky130_fd_sc_hd__buf_2
X_2124_ _1598_/Y vssd1 vssd1 vccd1 vccd1 _2124_/X sky130_fd_sc_hd__buf_2
XFILLER_66_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2055_ _1985_/Y _2067_/B vssd1 vssd1 vccd1 vccd1 _2055_/Y sky130_fd_sc_hd__nor2_4
XFILLER_34_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1839_ _1842_/A vssd1 vssd1 vccd1 vccd1 _1840_/A sky130_fd_sc_hd__buf_2
X_1908_ _1921_/A _1908_/B vssd1 vssd1 vccd1 vccd1 _1908_/Y sky130_fd_sc_hd__nor2_4
XFILLER_1_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1624_ _2435_/Q vssd1 vssd1 vccd1 vccd1 _1625_/C sky130_fd_sc_hd__inv_2
X_2673_ _2679_/CLK _1424_/Y vssd1 vssd1 vccd1 vccd1 _1252_/B sky130_fd_sc_hd__dfxtp_4
X_1555_ _2143_/A _1555_/B vssd1 vssd1 vccd1 vccd1 _1555_/Y sky130_fd_sc_hd__nor2_4
XFILLER_54_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1486_ _1450_/D _1486_/B vssd1 vssd1 vccd1 vccd1 _1486_/Y sky130_fd_sc_hd__nand2_4
X_2107_ _1212_/X ID_fromClient vssd1 vssd1 vccd1 vccd1 _2496_/D sky130_fd_sc_hd__and2_4
X_2038_ _2027_/B _2027_/A _2026_/X _1990_/A vssd1 vssd1 vccd1 vccd1 _2039_/C sky130_fd_sc_hd__nand4_4
XFILLER_45_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1340_ _1339_/Y vssd1 vssd1 vccd1 vccd1 _1340_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1271_ _1270_/Y vssd1 vssd1 vccd1 vccd1 _1282_/D sky130_fd_sc_hd__inv_2
XFILLER_36_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2656_ _2707_/CLK _1671_/Y vssd1 vssd1 vccd1 vccd1 _2190_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_59_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1538_ _1497_/A _1595_/A vssd1 vssd1 vccd1 vccd1 _1539_/A sky130_fd_sc_hd__nor2_4
X_1469_ _1454_/Y vssd1 vssd1 vccd1 vccd1 _1469_/X sky130_fd_sc_hd__buf_2
X_2587_ _2517_/CLK _2587_/D vssd1 vssd1 vccd1 vccd1 HASH_ADDR[2] sky130_fd_sc_hd__dfxtp_4
X_1607_ _1618_/B vssd1 vssd1 vccd1 vccd1 _1608_/B sky130_fd_sc_hd__inv_2
XFILLER_27_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2510_ _2707_/CLK _2088_/X vssd1 vssd1 vccd1 vccd1 _2392_/A sky130_fd_sc_hd__dfxtp_4
X_1323_ _1247_/A _1327_/A _1311_/X vssd1 vssd1 vccd1 vccd1 _1323_/X sky130_fd_sc_hd__o21a_4
XFILLER_38_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2372_ _1207_/A _2382_/C _2096_/A vssd1 vssd1 vccd1 vccd1 _2372_/X sky130_fd_sc_hd__a21o_4
X_2441_ _2443_/CLK _2441_/D vssd1 vssd1 vccd1 vccd1 _1761_/A sky130_fd_sc_hd__dfxtp_4
X_1254_ _1254_/A _1254_/B _1254_/C _1254_/D vssd1 vssd1 vccd1 vccd1 _1259_/B sky130_fd_sc_hd__nor4_4
XFILLER_32_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2708_ _2705_/CLK _2400_/Y vssd1 vssd1 vccd1 vccd1 _2397_/A sky130_fd_sc_hd__dfxtp_4
X_2639_ _2511_/CLK _2639_/D vssd1 vssd1 vccd1 vccd1 _1517_/A sky130_fd_sc_hd__dfxtp_4
XINSDIODE2_3 EXT_RESET_N_fromHost vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1872_ _1222_/A vssd1 vssd1 vccd1 vccd1 _1873_/A sky130_fd_sc_hd__buf_2
X_1941_ _1941_/A _2567_/Q vssd1 vssd1 vccd1 vccd1 _1941_/X sky130_fd_sc_hd__and2_4
XFILLER_14_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1306_ _1281_/C _1281_/D _1246_/Y vssd1 vssd1 vccd1 vccd1 _1306_/Y sky130_fd_sc_hd__o21ai_4
X_2286_ _2284_/X _2189_/X _2285_/Y vssd1 vssd1 vccd1 vccd1 _2479_/D sky130_fd_sc_hd__a21oi_4
X_2424_ _2517_/CLK _2423_/Q vssd1 vssd1 vccd1 vccd1 _2424_/Q sky130_fd_sc_hd__dfxtp_4
X_2355_ _1565_/B _2352_/X _1452_/X _2354_/X vssd1 vssd1 vccd1 vccd1 _2355_/X sky130_fd_sc_hd__a2bb2o_4
X_1237_ _1234_/Y _1235_/X _1236_/Y vssd1 vssd1 vccd1 vccd1 _1237_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_52_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2140_ _1295_/A _2139_/X _2187_/C _1539_/Y _1583_/X vssd1 vssd1 vccd1 vccd1 _2140_/Y
+ sky130_fd_sc_hd__o32ai_4
XFILLER_38_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2071_ _2066_/Y _2067_/B _1363_/C vssd1 vssd1 vccd1 vccd1 _2071_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_34_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1855_ _1858_/A _1855_/B vssd1 vssd1 vccd1 vccd1 _2612_/D sky130_fd_sc_hd__and2_4
X_1924_ _1875_/A vssd1 vssd1 vccd1 vccd1 _1930_/A sky130_fd_sc_hd__buf_2
X_1786_ _1964_/B _2633_/Q _1785_/X vssd1 vssd1 vccd1 vccd1 _1786_/X sky130_fd_sc_hd__o21a_4
X_2407_ _2670_/CLK _2407_/D vssd1 vssd1 vccd1 vccd1 _1273_/A sky130_fd_sc_hd__dfxtp_4
X_2338_ _2296_/Y _2333_/X _2337_/Y vssd1 vssd1 vccd1 vccd1 _2453_/D sky130_fd_sc_hd__o21ai_4
X_2269_ _1934_/B _2170_/X _2268_/Y vssd1 vssd1 vccd1 vccd1 _2270_/B sky130_fd_sc_hd__o21ai_4
XFILLER_4_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1571_ _1510_/A _1571_/B _1571_/C vssd1 vssd1 vccd1 vccd1 _1572_/A sky130_fd_sc_hd__nor3_4
XFILLER_6_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1640_ _2453_/Q _2272_/A _1548_/X _1639_/Y vssd1 vssd1 vccd1 vccd1 _1640_/X sky130_fd_sc_hd__a211o_4
XFILLER_66_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2123_ _1626_/Y vssd1 vssd1 vccd1 vccd1 _2123_/X sky130_fd_sc_hd__buf_2
X_2054_ _2048_/C vssd1 vssd1 vccd1 vccd1 _2067_/B sky130_fd_sc_hd__buf_2
XFILLER_34_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1838_ _1838_/A vssd1 vssd1 vccd1 vccd1 _1842_/A sky130_fd_sc_hd__buf_2
X_1907_ _2245_/B vssd1 vssd1 vccd1 vccd1 _1908_/B sky130_fd_sc_hd__inv_2
XFILLER_66_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1769_ _1767_/Y _1768_/Y _1722_/X vssd1 vssd1 vccd1 vccd1 _2646_/D sky130_fd_sc_hd__a21oi_4
XFILLER_13_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2672_ _2679_/CLK _1428_/Y vssd1 vssd1 vccd1 vccd1 _2672_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1623_ _1667_/B _1623_/B _1633_/D vssd1 vssd1 vccd1 vccd1 _1623_/Y sky130_fd_sc_hd__nor3_4
X_1485_ _1457_/X vssd1 vssd1 vccd1 vccd1 _1485_/Y sky130_fd_sc_hd__inv_2
X_1554_ _1554_/A vssd1 vssd1 vccd1 vccd1 _1555_/B sky130_fd_sc_hd__inv_2
.ends


magic
tech sky130A
magscale 1 2
timestamp 1608074288
<< locali >>
rect 312093 382007 312127 382449
rect 306849 360723 306883 365789
rect 195805 276403 195839 276505
rect 206017 276335 206051 276505
rect 216413 276403 216447 276505
rect 226625 276335 226659 276505
rect 237021 276403 237055 276573
rect 247141 276335 247175 276573
rect 208995 276301 209053 276335
rect 229603 276301 229661 276335
rect 257629 276131 257663 276301
rect 260515 276233 260665 276267
rect 269773 275927 269807 276165
rect 292221 275995 292255 276165
rect 291979 275961 292255 275995
rect 558561 105995 558595 113305
rect 558745 92803 558779 102969
rect 264989 71383 265023 71825
<< viali >>
rect 312093 382449 312127 382483
rect 312093 381973 312127 382007
rect 306849 365789 306883 365823
rect 306849 360689 306883 360723
rect 237021 276573 237055 276607
rect 195805 276505 195839 276539
rect 195805 276369 195839 276403
rect 206017 276505 206051 276539
rect 216413 276505 216447 276539
rect 216413 276369 216447 276403
rect 226625 276505 226659 276539
rect 237021 276369 237055 276403
rect 247141 276573 247175 276607
rect 206017 276301 206051 276335
rect 208961 276301 208995 276335
rect 209053 276301 209087 276335
rect 226625 276301 226659 276335
rect 229569 276301 229603 276335
rect 229661 276301 229695 276335
rect 247141 276301 247175 276335
rect 257629 276301 257663 276335
rect 260481 276233 260515 276267
rect 260665 276233 260699 276267
rect 257629 276097 257663 276131
rect 269773 276165 269807 276199
rect 292221 276165 292255 276199
rect 291945 275961 291979 275995
rect 269773 275893 269807 275927
rect 558561 113305 558595 113339
rect 558561 105961 558595 105995
rect 558745 102969 558779 103003
rect 558745 92769 558779 92803
rect 264989 71825 265023 71859
rect 264989 71349 265023 71383
<< metal1 >>
rect 8018 700612 8024 700664
rect 8076 700652 8082 700664
rect 8202 700652 8208 700664
rect 8076 700624 8208 700652
rect 8076 700612 8082 700624
rect 8202 700612 8208 700624
rect 8260 700652 8266 700664
rect 72970 700652 72976 700664
rect 8260 700624 72976 700652
rect 8260 700612 8266 700624
rect 72970 700612 72976 700624
rect 73028 700652 73034 700664
rect 137830 700652 137836 700664
rect 73028 700624 137836 700652
rect 73028 700612 73034 700624
rect 137830 700612 137836 700624
rect 137888 700652 137894 700664
rect 202782 700652 202788 700664
rect 137888 700624 202788 700652
rect 137888 700612 137894 700624
rect 202782 700612 202788 700624
rect 202840 700612 202846 700664
rect 267642 700612 267648 700664
rect 267700 700652 267706 700664
rect 332502 700652 332508 700664
rect 267700 700624 332508 700652
rect 267700 700612 267706 700624
rect 332502 700612 332508 700624
rect 332560 700652 332566 700664
rect 397454 700652 397460 700664
rect 332560 700624 397460 700652
rect 332560 700612 332566 700624
rect 397454 700612 397460 700624
rect 397512 700652 397518 700664
rect 462314 700652 462320 700664
rect 397512 700624 462320 700652
rect 397512 700612 397518 700624
rect 462314 700612 462320 700624
rect 462372 700652 462378 700664
rect 527174 700652 527180 700664
rect 462372 700624 527180 700652
rect 462372 700612 462378 700624
rect 527174 700612 527180 700624
rect 527232 700612 527238 700664
rect 24302 700544 24308 700596
rect 24360 700584 24366 700596
rect 24946 700584 24952 700596
rect 24360 700556 24952 700584
rect 24360 700544 24366 700556
rect 24946 700544 24952 700556
rect 25004 700544 25010 700596
rect 218974 700000 218980 700052
rect 219032 700040 219038 700052
rect 272978 700040 272984 700052
rect 219032 700012 272984 700040
rect 219032 700000 219038 700012
rect 272978 700000 272984 700012
rect 273036 700000 273042 700052
rect 295794 700000 295800 700052
rect 295852 700040 295858 700052
rect 429838 700040 429844 700052
rect 295852 700012 429844 700040
rect 295852 700000 295858 700012
rect 429838 700000 429844 700012
rect 429896 700000 429902 700052
rect 154114 699932 154120 699984
rect 154172 699972 154178 699984
rect 268562 699972 268568 699984
rect 154172 699944 268568 699972
rect 154172 699932 154178 699944
rect 268562 699932 268568 699944
rect 268620 699932 268626 699984
rect 304626 699932 304632 699984
rect 304684 699972 304690 699984
rect 494790 699972 494796 699984
rect 304684 699944 494796 699972
rect 304684 699932 304690 699944
rect 494790 699932 494796 699944
rect 494848 699932 494854 699984
rect 527174 699932 527180 699984
rect 527232 699972 527238 699984
rect 579890 699972 579896 699984
rect 527232 699944 579896 699972
rect 527232 699932 527238 699944
rect 579890 699932 579896 699944
rect 579948 699932 579954 699984
rect 89162 699864 89168 699916
rect 89220 699904 89226 699916
rect 277394 699904 277400 699916
rect 89220 699876 277400 699904
rect 89220 699864 89226 699876
rect 277394 699864 277400 699876
rect 277452 699864 277458 699916
rect 288434 699864 288440 699916
rect 288492 699904 288498 699916
rect 559650 699904 559656 699916
rect 288492 699876 559656 699904
rect 288492 699864 288498 699876
rect 559650 699864 559656 699876
rect 559708 699864 559714 699916
rect 314194 674160 314200 674212
rect 314252 674200 314258 674212
rect 578510 674200 578516 674212
rect 314252 674172 578516 674200
rect 314252 674160 314258 674172
rect 578510 674160 578516 674172
rect 578568 674160 578574 674212
rect 2958 653488 2964 653540
rect 3016 653528 3022 653540
rect 8018 653528 8024 653540
rect 3016 653500 8024 653528
rect 3016 653488 3022 653500
rect 8018 653488 8024 653500
rect 8076 653488 8082 653540
rect 310514 627104 310520 627156
rect 310572 627144 310578 627156
rect 578786 627144 578792 627156
rect 310572 627116 578792 627144
rect 310572 627104 310578 627116
rect 578786 627104 578792 627116
rect 578844 627104 578850 627156
rect 193858 586440 193864 586492
rect 193916 586480 193922 586492
rect 292758 586480 292764 586492
rect 193916 586452 292764 586480
rect 193916 586440 193922 586452
rect 292758 586440 292764 586452
rect 292816 586440 292822 586492
rect 265986 586372 265992 586424
rect 266044 586412 266050 586424
rect 313642 586412 313648 586424
rect 266044 586384 313648 586412
rect 266044 586372 266050 586384
rect 313642 586372 313648 586384
rect 313700 586372 313706 586424
rect 242066 586304 242072 586356
rect 242124 586344 242130 586356
rect 307478 586344 307484 586356
rect 242124 586316 307484 586344
rect 242124 586304 242130 586316
rect 307478 586304 307484 586316
rect 307536 586304 307542 586356
rect 217962 586236 217968 586288
rect 218020 586276 218026 586288
rect 306834 586276 306840 586288
rect 218020 586248 306840 586276
rect 218020 586236 218026 586248
rect 306834 586236 306840 586248
rect 306892 586276 306898 586288
rect 307570 586276 307576 586288
rect 306892 586248 307576 586276
rect 306892 586236 306898 586248
rect 307570 586236 307576 586248
rect 307628 586236 307634 586288
rect 276658 586168 276664 586220
rect 276716 586208 276722 586220
rect 365438 586208 365444 586220
rect 276716 586180 365444 586208
rect 276716 586168 276722 586180
rect 365438 586168 365444 586180
rect 365496 586168 365502 586220
rect 291378 586100 291384 586152
rect 291436 586140 291442 586152
rect 341518 586140 341524 586152
rect 291436 586112 341524 586140
rect 291436 586100 291442 586112
rect 341518 586100 341524 586112
rect 341576 586100 341582 586152
rect 169754 586032 169760 586084
rect 169812 586072 169818 586084
rect 294414 586072 294420 586084
rect 169812 586044 294420 586072
rect 169812 586032 169818 586044
rect 294414 586032 294420 586044
rect 294472 586032 294478 586084
rect 73522 585964 73528 586016
rect 73580 586004 73586 586016
rect 275922 586004 275928 586016
rect 73580 585976 275928 586004
rect 73580 585964 73586 585976
rect 275922 585964 275928 585976
rect 275980 586004 275986 586016
rect 276658 586004 276664 586016
rect 275980 585976 276664 586004
rect 275980 585964 275986 585976
rect 276658 585964 276664 585976
rect 276716 585964 276722 586016
rect 307570 585964 307576 586016
rect 307628 586004 307634 586016
rect 509878 586004 509884 586016
rect 307628 585976 509884 586004
rect 307628 585964 307634 585976
rect 509878 585964 509884 585976
rect 509936 585964 509942 586016
rect 49602 585896 49608 585948
rect 49660 585936 49666 585948
rect 291378 585936 291384 585948
rect 49660 585908 291384 585936
rect 49660 585896 49666 585908
rect 291378 585896 291384 585908
rect 291436 585896 291442 585948
rect 313642 585896 313648 585948
rect 313700 585936 313706 585948
rect 557902 585936 557908 585948
rect 313700 585908 557908 585936
rect 313700 585896 313706 585908
rect 557902 585896 557908 585908
rect 557960 585896 557966 585948
rect 26510 582360 26516 582412
rect 26568 582400 26574 582412
rect 267090 582400 267096 582412
rect 26568 582372 267096 582400
rect 26568 582360 26574 582372
rect 267090 582360 267096 582372
rect 267148 582360 267154 582412
rect 24762 582292 24768 582344
rect 24820 582332 24826 582344
rect 286226 582332 286232 582344
rect 24820 582304 286232 582332
rect 24820 582292 24826 582304
rect 286226 582292 286232 582304
rect 286284 582292 286290 582344
rect 319806 582292 319812 582344
rect 319864 582332 319870 582344
rect 558638 582332 558644 582344
rect 319864 582304 558644 582332
rect 319864 582292 319870 582304
rect 558638 582292 558644 582304
rect 558696 582292 558702 582344
rect 27246 582224 27252 582276
rect 27304 582264 27310 582276
rect 314930 582264 314936 582276
rect 27304 582236 314936 582264
rect 27304 582224 27310 582236
rect 314930 582224 314936 582236
rect 314988 582224 314994 582276
rect 318610 582224 318616 582276
rect 318668 582264 318674 582276
rect 560846 582264 560852 582276
rect 318668 582236 560852 582264
rect 318668 582224 318674 582236
rect 560846 582224 560852 582236
rect 560904 582224 560910 582276
rect 314286 579980 314292 580032
rect 314344 580020 314350 580032
rect 314930 580020 314936 580032
rect 314344 579992 314936 580020
rect 314344 579980 314350 579992
rect 314930 579980 314936 579992
rect 314988 579980 314994 580032
rect 319806 580020 319812 580032
rect 317984 579992 319812 580020
rect 317414 579912 317420 579964
rect 317472 579952 317478 579964
rect 317984 579952 318012 579992
rect 319806 579980 319812 579992
rect 319864 579980 319870 580032
rect 558546 579980 558552 580032
rect 558604 580020 558610 580032
rect 578786 580020 578792 580032
rect 558604 579992 578792 580020
rect 558604 579980 558610 579992
rect 578786 579980 578792 579992
rect 578844 579980 578850 580032
rect 317472 579924 318012 579952
rect 317472 579912 317478 579924
rect 26510 574104 26516 574116
rect 25056 574076 26516 574104
rect 24854 573996 24860 574048
rect 24912 574036 24918 574048
rect 25056 574036 25084 574076
rect 26510 574064 26516 574076
rect 26568 574064 26574 574116
rect 313550 574064 313556 574116
rect 313608 574104 313614 574116
rect 317414 574104 317420 574116
rect 313608 574076 317420 574104
rect 313608 574064 313614 574076
rect 317414 574064 317420 574076
rect 317472 574064 317478 574116
rect 24912 574008 25084 574036
rect 24912 573996 24918 574008
rect 311618 571140 311624 571192
rect 311676 571180 311682 571192
rect 313550 571180 313556 571192
rect 311676 571152 313556 571180
rect 311676 571140 311682 571152
rect 313550 571140 313556 571152
rect 313608 571140 313614 571192
rect 269298 547612 269304 547664
rect 269356 547652 269362 547664
rect 291286 547652 291292 547664
rect 269356 547624 291292 547652
rect 269356 547612 269362 547624
rect 291286 547612 291292 547624
rect 291344 547612 291350 547664
rect 286226 545300 286232 545352
rect 286284 545340 286290 545352
rect 315022 545340 315028 545352
rect 286284 545312 315028 545340
rect 286284 545300 286290 545312
rect 315022 545300 315028 545312
rect 315080 545300 315086 545352
rect 267090 531972 267096 532024
rect 267148 532012 267154 532024
rect 269298 532012 269304 532024
rect 267148 531984 269304 532012
rect 267148 531972 267154 531984
rect 269298 531972 269304 531984
rect 269356 531972 269362 532024
rect 269298 529932 269304 529984
rect 269356 529972 269362 529984
rect 269356 529944 269436 529972
rect 269356 529932 269362 529944
rect 269408 529904 269436 529944
rect 272334 529904 272340 529916
rect 269408 529876 272340 529904
rect 272334 529864 272340 529876
rect 272392 529864 272398 529916
rect 272334 523948 272340 524000
rect 272392 523988 272398 524000
rect 274450 523988 274456 524000
rect 272392 523960 274456 523988
rect 272392 523948 272398 523960
rect 274450 523948 274456 523960
rect 274508 523948 274514 524000
rect 558638 516604 558644 516656
rect 558696 516644 558702 516656
rect 560018 516644 560024 516656
rect 558696 516616 560024 516644
rect 558696 516604 558702 516616
rect 560018 516604 560024 516616
rect 560076 516604 560082 516656
rect 274450 514428 274456 514480
rect 274508 514468 274514 514480
rect 278590 514468 278596 514480
rect 274508 514440 278596 514468
rect 274508 514428 274514 514440
rect 278590 514428 278596 514440
rect 278648 514428 278654 514480
rect 278590 513272 278596 513324
rect 278648 513312 278654 513324
rect 282546 513312 282552 513324
rect 278648 513284 282552 513312
rect 278648 513272 278654 513284
rect 282546 513272 282552 513284
rect 282604 513272 282610 513324
rect 269298 511504 269304 511556
rect 269356 511544 269362 511556
rect 309318 511544 309324 511556
rect 269356 511516 309324 511544
rect 269356 511504 269362 511516
rect 309318 511504 309324 511516
rect 309376 511504 309382 511556
rect 282638 509328 282644 509380
rect 282696 509368 282702 509380
rect 315022 509368 315028 509380
rect 282696 509340 315028 509368
rect 282696 509328 282702 509340
rect 315022 509328 315028 509340
rect 315080 509328 315086 509380
rect 558638 485800 558644 485852
rect 558696 485840 558702 485852
rect 578786 485840 578792 485852
rect 558696 485812 578792 485840
rect 558696 485800 558702 485812
rect 578786 485800 578792 485812
rect 578844 485800 578850 485852
rect 558730 438676 558736 438728
rect 558788 438716 558794 438728
rect 578786 438716 578792 438728
rect 558788 438688 578792 438716
rect 558788 438676 558794 438688
rect 578786 438676 578792 438688
rect 578844 438676 578850 438728
rect 560018 421880 560024 421932
rect 560076 421920 560082 421932
rect 560846 421920 560852 421932
rect 560076 421892 560852 421920
rect 560076 421880 560082 421892
rect 560846 421880 560852 421892
rect 560904 421880 560910 421932
rect 269298 404812 269304 404864
rect 269356 404852 269362 404864
rect 286318 404852 286324 404864
rect 269356 404824 286324 404852
rect 269356 404812 269362 404824
rect 286318 404812 286324 404824
rect 286376 404812 286382 404864
rect 299474 401888 299480 401940
rect 299532 401928 299538 401940
rect 315022 401928 315028 401940
rect 299532 401900 315028 401928
rect 299532 401888 299538 401900
rect 315022 401888 315028 401900
rect 315080 401888 315086 401940
rect 558822 397468 558828 397520
rect 558880 397508 558886 397520
rect 560018 397508 560024 397520
rect 558880 397480 560024 397508
rect 558880 397468 558886 397480
rect 560018 397468 560024 397480
rect 560076 397468 560082 397520
rect 270586 386316 270592 386368
rect 270644 386356 270650 386368
rect 558822 386356 558828 386368
rect 270644 386328 558828 386356
rect 270644 386316 270650 386328
rect 558822 386316 558828 386328
rect 558880 386316 558886 386368
rect 24854 386248 24860 386300
rect 24912 386288 24918 386300
rect 298830 386288 298836 386300
rect 24912 386260 298836 386288
rect 24912 386248 24918 386260
rect 298830 386248 298836 386260
rect 298888 386248 298894 386300
rect 270034 386180 270040 386232
rect 270092 386220 270098 386232
rect 270586 386220 270592 386232
rect 270092 386192 270592 386220
rect 270092 386180 270098 386192
rect 270586 386180 270592 386192
rect 270644 386180 270650 386232
rect 298830 385908 298836 385960
rect 298888 385948 298894 385960
rect 299474 385948 299480 385960
rect 298888 385920 299480 385948
rect 298888 385908 298894 385920
rect 299474 385908 299480 385920
rect 299532 385908 299538 385960
rect 286318 385636 286324 385688
rect 286376 385676 286382 385688
rect 293678 385676 293684 385688
rect 286376 385648 293684 385676
rect 286376 385636 286382 385648
rect 293678 385636 293684 385648
rect 293736 385676 293742 385688
rect 560846 385676 560852 385688
rect 293736 385648 560852 385676
rect 293736 385636 293742 385648
rect 560846 385636 560852 385648
rect 560904 385636 560910 385688
rect 87690 382644 87696 382696
rect 87748 382684 87754 382696
rect 294414 382684 294420 382696
rect 87748 382656 294420 382684
rect 87748 382644 87754 382656
rect 294414 382644 294420 382656
rect 294472 382644 294478 382696
rect 135898 382576 135904 382628
rect 135956 382616 135962 382628
rect 276382 382616 276388 382628
rect 135956 382588 276388 382616
rect 135956 382576 135962 382588
rect 276382 382576 276388 382588
rect 276440 382576 276446 382628
rect 256050 382508 256056 382560
rect 256108 382548 256114 382560
rect 300118 382548 300124 382560
rect 256108 382520 300124 382548
rect 256108 382508 256114 382520
rect 300118 382508 300124 382520
rect 300176 382508 300182 382560
rect 312081 382483 312139 382489
rect 312081 382449 312093 382483
rect 312127 382480 312139 382483
rect 313550 382480 313556 382492
rect 312127 382452 313556 382480
rect 312127 382449 312139 382452
rect 312081 382443 312139 382449
rect 313550 382440 313556 382452
rect 313608 382480 313614 382492
rect 331490 382480 331496 382492
rect 313608 382452 331496 382480
rect 313608 382440 313614 382452
rect 331490 382440 331496 382452
rect 331548 382440 331554 382492
rect 232130 382372 232136 382424
rect 232188 382412 232194 382424
rect 313734 382412 313740 382424
rect 232188 382384 313740 382412
rect 232188 382372 232194 382384
rect 313734 382372 313740 382384
rect 313792 382372 313798 382424
rect 270770 382304 270776 382356
rect 270828 382344 270834 382356
rect 355594 382344 355600 382356
rect 270828 382316 355600 382344
rect 270828 382304 270834 382316
rect 355594 382304 355600 382316
rect 355652 382304 355658 382356
rect 208026 382236 208032 382288
rect 208084 382276 208090 382288
rect 313550 382276 313556 382288
rect 208084 382248 313556 382276
rect 208084 382236 208090 382248
rect 313550 382236 313556 382248
rect 313608 382236 313614 382288
rect 111794 382168 111800 382220
rect 111852 382208 111858 382220
rect 274450 382208 274456 382220
rect 111852 382180 274456 382208
rect 111852 382168 111858 382180
rect 274450 382168 274456 382180
rect 274508 382208 274514 382220
rect 403618 382208 403624 382220
rect 274508 382180 403624 382208
rect 274508 382168 274514 382180
rect 403618 382168 403624 382180
rect 403676 382168 403682 382220
rect 183922 382100 183928 382152
rect 183980 382140 183986 382152
rect 270678 382140 270684 382152
rect 183980 382112 270684 382140
rect 183980 382100 183986 382112
rect 270678 382100 270684 382112
rect 270736 382140 270742 382152
rect 475930 382140 475936 382152
rect 270736 382112 475936 382140
rect 270736 382100 270742 382112
rect 475930 382100 475936 382112
rect 475988 382100 475994 382152
rect 63770 382032 63776 382084
rect 63828 382072 63834 382084
rect 270770 382072 270776 382084
rect 63828 382044 270776 382072
rect 63828 382032 63834 382044
rect 270770 382032 270776 382044
rect 270828 382032 270834 382084
rect 313550 382032 313556 382084
rect 313608 382072 313614 382084
rect 313826 382072 313832 382084
rect 313608 382044 313832 382072
rect 313608 382032 313614 382044
rect 313826 382032 313832 382044
rect 313884 382072 313890 382084
rect 499850 382072 499856 382084
rect 313884 382044 499856 382072
rect 313884 382032 313890 382044
rect 499850 382032 499856 382044
rect 499908 382032 499914 382084
rect 39666 381964 39672 382016
rect 39724 382004 39730 382016
rect 312081 382007 312139 382013
rect 312081 382004 312093 382007
rect 39724 381976 312093 382004
rect 39724 381964 39730 381976
rect 312081 381973 312093 381976
rect 312127 381973 312139 382007
rect 312081 381967 312139 381973
rect 313734 381964 313740 382016
rect 313792 382004 313798 382016
rect 523954 382004 523960 382016
rect 313792 381976 523960 382004
rect 313792 381964 313798 381976
rect 523954 381964 523960 381976
rect 524012 381964 524018 382016
rect 306834 365820 306840 365832
rect 306795 365792 306840 365820
rect 306834 365780 306840 365792
rect 306892 365780 306898 365832
rect 306837 360723 306895 360729
rect 306837 360689 306849 360723
rect 306883 360720 306895 360723
rect 306926 360720 306932 360732
rect 306883 360692 306932 360720
rect 306883 360689 306895 360692
rect 306837 360683 306895 360689
rect 306926 360680 306932 360692
rect 306984 360680 306990 360732
rect 309134 359116 309140 359168
rect 309192 359156 309198 359168
rect 310514 359156 310520 359168
rect 309192 359128 310520 359156
rect 309192 359116 309198 359128
rect 310514 359116 310520 359128
rect 310572 359116 310578 359168
rect 277394 358504 277400 358556
rect 277452 358544 277458 358556
rect 292574 358544 292580 358556
rect 277452 358516 292580 358544
rect 277452 358504 277458 358516
rect 292574 358504 292580 358516
rect 292632 358504 292638 358556
rect 3786 358436 3792 358488
rect 3844 358476 3850 358488
rect 278406 358476 278412 358488
rect 3844 358448 278412 358476
rect 3844 358436 3850 358448
rect 278406 358436 278412 358448
rect 278464 358436 278470 358488
rect 294966 358436 294972 358488
rect 295024 358476 295030 358488
rect 295794 358476 295800 358488
rect 295024 358448 295800 358476
rect 295024 358436 295030 358448
rect 295794 358436 295800 358448
rect 295852 358436 295858 358488
rect 3694 358368 3700 358420
rect 3752 358408 3758 358420
rect 280798 358408 280804 358420
rect 3752 358380 280804 358408
rect 3752 358368 3758 358380
rect 280798 358368 280804 358380
rect 280856 358368 280862 358420
rect 273070 357688 273076 357740
rect 273128 357728 273134 357740
rect 311342 357728 311348 357740
rect 273128 357700 311348 357728
rect 273128 357688 273134 357700
rect 311342 357688 311348 357700
rect 311400 357688 311406 357740
rect 270402 354016 270408 354068
rect 270460 354056 270466 354068
rect 579338 354056 579344 354068
rect 270460 354028 579344 354056
rect 270460 354016 270466 354028
rect 579338 354016 579344 354028
rect 579396 354016 579402 354068
rect 270494 353948 270500 354000
rect 270552 353988 270558 354000
rect 579154 353988 579160 354000
rect 270552 353960 579160 353988
rect 270552 353948 270558 353960
rect 579154 353948 579160 353960
rect 579212 353948 579218 354000
rect 314010 344360 314016 344412
rect 314068 344400 314074 344412
rect 558638 344400 558644 344412
rect 314068 344372 558644 344400
rect 314068 344360 314074 344372
rect 558638 344360 558644 344372
rect 558696 344360 558702 344412
rect 314010 341436 314016 341488
rect 314068 341476 314074 341488
rect 579246 341476 579252 341488
rect 314068 341448 579252 341476
rect 314068 341436 314074 341448
rect 579246 341436 579252 341448
rect 579304 341436 579310 341488
rect 268562 339940 268568 339992
rect 268620 339980 268626 339992
rect 270218 339980 270224 339992
rect 268620 339952 270224 339980
rect 268620 339940 268626 339952
rect 270218 339940 270224 339952
rect 270276 339940 270282 339992
rect 3970 332596 3976 332648
rect 4028 332636 4034 332648
rect 269390 332636 269396 332648
rect 4028 332608 269396 332636
rect 4028 332596 4034 332608
rect 269390 332596 269396 332608
rect 269448 332596 269454 332648
rect 24854 328244 24860 328296
rect 24912 328284 24918 328296
rect 269390 328284 269396 328296
rect 24912 328256 269396 328284
rect 24912 328244 24918 328256
rect 269390 328244 269396 328256
rect 269448 328244 269454 328296
rect 24946 325252 24952 325304
rect 25004 325292 25010 325304
rect 269390 325292 269396 325304
rect 25004 325264 269396 325292
rect 25004 325252 25010 325264
rect 269390 325252 269396 325264
rect 269448 325252 269454 325304
rect 313642 323892 313648 323944
rect 313700 323932 313706 323944
rect 314010 323932 314016 323944
rect 313700 323904 314016 323932
rect 313700 323892 313706 323904
rect 314010 323892 314016 323904
rect 314068 323892 314074 323944
rect 313642 323756 313648 323808
rect 313700 323796 313706 323808
rect 558546 323796 558552 323808
rect 313700 323768 558552 323796
rect 313700 323756 313706 323768
rect 558546 323756 558552 323768
rect 558604 323756 558610 323808
rect 3602 317908 3608 317960
rect 3660 317948 3666 317960
rect 311526 317948 311532 317960
rect 3660 317920 311532 317948
rect 3660 317908 3666 317920
rect 311526 317908 311532 317920
rect 311584 317908 311590 317960
rect 309134 314712 309140 314764
rect 309192 314752 309198 314764
rect 310514 314752 310520 314764
rect 309192 314724 310520 314752
rect 309192 314712 309198 314724
rect 310514 314712 310520 314724
rect 310572 314712 310578 314764
rect 3878 313488 3884 313540
rect 3936 313528 3942 313540
rect 304350 313528 304356 313540
rect 3936 313500 304356 313528
rect 3936 313488 3942 313500
rect 304350 313488 304356 313500
rect 304408 313488 304414 313540
rect 283190 313420 283196 313472
rect 283248 313460 283254 313472
rect 558730 313460 558736 313472
rect 283248 313432 558736 313460
rect 283248 313420 283254 313432
rect 558730 313420 558736 313432
rect 558788 313420 558794 313472
rect 272978 313352 272984 313404
rect 273036 313392 273042 313404
rect 297358 313392 297364 313404
rect 273036 313364 297364 313392
rect 273036 313352 273042 313364
rect 297358 313352 297364 313364
rect 297416 313352 297422 313404
rect 98546 312740 98552 312792
rect 98604 312780 98610 312792
rect 278590 312780 278596 312792
rect 98604 312752 278596 312780
rect 98604 312740 98610 312752
rect 278590 312740 278596 312752
rect 278648 312740 278654 312792
rect 306742 309136 306748 309188
rect 306800 309176 306806 309188
rect 307110 309176 307116 309188
rect 306800 309148 307116 309176
rect 306800 309136 306806 309148
rect 307110 309136 307116 309148
rect 307168 309136 307174 309188
rect 306558 298732 306564 298784
rect 306616 298772 306622 298784
rect 306834 298772 306840 298784
rect 306616 298744 306840 298772
rect 306616 298732 306622 298744
rect 306834 298732 306840 298744
rect 306892 298732 306898 298784
rect 306742 281120 306748 281172
rect 306800 281160 306806 281172
rect 306926 281160 306932 281172
rect 306800 281132 306932 281160
rect 306800 281120 306806 281132
rect 306926 281120 306932 281132
rect 306984 281120 306990 281172
rect 97994 276700 98000 276752
rect 98052 276740 98058 276752
rect 98546 276740 98552 276752
rect 98052 276712 98552 276740
rect 98052 276700 98058 276712
rect 98546 276700 98552 276712
rect 98604 276700 98610 276752
rect 237009 276607 237067 276613
rect 237009 276573 237021 276607
rect 237055 276604 237067 276607
rect 247129 276607 247187 276613
rect 247129 276604 247141 276607
rect 237055 276576 247141 276604
rect 237055 276573 237067 276576
rect 237009 276567 237067 276573
rect 247129 276573 247141 276576
rect 247175 276573 247187 276607
rect 247129 276567 247187 276573
rect 195793 276539 195851 276545
rect 195793 276505 195805 276539
rect 195839 276536 195851 276539
rect 206005 276539 206063 276545
rect 206005 276536 206017 276539
rect 195839 276508 206017 276536
rect 195839 276505 195851 276508
rect 195793 276499 195851 276505
rect 206005 276505 206017 276508
rect 206051 276505 206063 276539
rect 206005 276499 206063 276505
rect 216401 276539 216459 276545
rect 216401 276505 216413 276539
rect 216447 276536 216459 276539
rect 226613 276539 226671 276545
rect 226613 276536 226625 276539
rect 216447 276508 226625 276536
rect 216447 276505 216459 276508
rect 216401 276499 216459 276505
rect 226613 276505 226625 276508
rect 226659 276505 226671 276539
rect 226613 276499 226671 276505
rect 247328 276440 257568 276468
rect 194226 276360 194232 276412
rect 194284 276400 194290 276412
rect 195793 276403 195851 276409
rect 195793 276400 195805 276403
rect 194284 276372 195805 276400
rect 194284 276360 194290 276372
rect 195793 276369 195805 276372
rect 195839 276369 195851 276403
rect 216401 276403 216459 276409
rect 216401 276400 216413 276403
rect 195793 276363 195851 276369
rect 211172 276372 216413 276400
rect 206005 276335 206063 276341
rect 206005 276301 206017 276335
rect 206051 276332 206063 276335
rect 208949 276335 209007 276341
rect 208949 276332 208961 276335
rect 206051 276304 208961 276332
rect 206051 276301 206063 276304
rect 206005 276295 206063 276301
rect 208949 276301 208961 276304
rect 208995 276301 209007 276335
rect 208949 276295 209007 276301
rect 209041 276335 209099 276341
rect 209041 276301 209053 276335
rect 209087 276332 209099 276335
rect 211172 276332 211200 276372
rect 216401 276369 216413 276372
rect 216447 276369 216459 276403
rect 237009 276403 237067 276409
rect 237009 276400 237021 276403
rect 216401 276363 216459 276369
rect 231780 276372 237021 276400
rect 209087 276304 211200 276332
rect 226613 276335 226671 276341
rect 209087 276301 209099 276304
rect 209041 276295 209099 276301
rect 226613 276301 226625 276335
rect 226659 276332 226671 276335
rect 229557 276335 229615 276341
rect 229557 276332 229569 276335
rect 226659 276304 229569 276332
rect 226659 276301 226671 276304
rect 226613 276295 226671 276301
rect 229557 276301 229569 276304
rect 229603 276301 229615 276335
rect 229557 276295 229615 276301
rect 229649 276335 229707 276341
rect 229649 276301 229661 276335
rect 229695 276332 229707 276335
rect 231780 276332 231808 276372
rect 237009 276369 237021 276372
rect 237055 276369 237067 276403
rect 237009 276363 237067 276369
rect 229695 276304 231808 276332
rect 247129 276335 247187 276341
rect 229695 276301 229707 276304
rect 229649 276295 229707 276301
rect 247129 276301 247141 276335
rect 247175 276332 247187 276335
rect 247328 276332 247356 276440
rect 257540 276400 257568 276440
rect 257540 276372 257660 276400
rect 257632 276341 257660 276372
rect 247175 276304 247356 276332
rect 257617 276335 257675 276341
rect 247175 276301 247187 276304
rect 247129 276295 247187 276301
rect 257617 276301 257629 276335
rect 257663 276301 257675 276335
rect 257617 276295 257675 276301
rect 266354 276292 266360 276344
rect 266412 276332 266418 276344
rect 313642 276332 313648 276344
rect 266412 276304 313648 276332
rect 266412 276292 266418 276304
rect 313642 276292 313648 276304
rect 313700 276292 313706 276344
rect 242434 276224 242440 276276
rect 242492 276264 242498 276276
rect 260469 276267 260527 276273
rect 260469 276264 260481 276267
rect 242492 276236 260481 276264
rect 242492 276224 242498 276236
rect 260469 276233 260481 276236
rect 260515 276233 260527 276267
rect 260469 276227 260527 276233
rect 260653 276267 260711 276273
rect 260653 276233 260665 276267
rect 260699 276264 260711 276267
rect 306926 276264 306932 276276
rect 260699 276236 306932 276264
rect 260699 276233 260711 276236
rect 260653 276227 260711 276233
rect 306926 276224 306932 276236
rect 306984 276224 306990 276276
rect 269761 276199 269819 276205
rect 269761 276196 269773 276199
rect 260668 276168 269773 276196
rect 257617 276131 257675 276137
rect 257617 276097 257629 276131
rect 257663 276128 257675 276131
rect 260668 276128 260696 276168
rect 269761 276165 269773 276168
rect 269807 276165 269819 276199
rect 269761 276159 269819 276165
rect 292209 276199 292267 276205
rect 292209 276165 292221 276199
rect 292255 276196 292267 276199
rect 295150 276196 295156 276208
rect 292255 276168 295156 276196
rect 292255 276165 292267 276168
rect 292209 276159 292267 276165
rect 295150 276156 295156 276168
rect 295208 276196 295214 276208
rect 461946 276196 461952 276208
rect 295208 276168 461952 276196
rect 295208 276156 295214 276168
rect 461946 276156 461952 276168
rect 462004 276156 462010 276208
rect 486050 276128 486056 276140
rect 257663 276100 260696 276128
rect 295812 276100 486056 276128
rect 257663 276097 257675 276100
rect 257617 276091 257675 276097
rect 170122 275952 170128 276004
rect 170180 275992 170186 276004
rect 291933 275995 291991 276001
rect 291933 275992 291945 275995
rect 170180 275964 291945 275992
rect 170180 275952 170186 275964
rect 291933 275961 291945 275964
rect 291979 275961 291991 275995
rect 291933 275955 291991 275961
rect 269761 275927 269819 275933
rect 269761 275893 269773 275927
rect 269807 275924 269819 275927
rect 292114 275924 292120 275936
rect 269807 275896 292120 275924
rect 269807 275893 269819 275896
rect 269761 275887 269819 275893
rect 292114 275884 292120 275896
rect 292172 275924 292178 275936
rect 295812 275924 295840 276100
rect 486050 276088 486056 276100
rect 486108 276088 486114 276140
rect 306926 276020 306932 276072
rect 306984 276060 306990 276072
rect 534258 276060 534264 276072
rect 306984 276032 534264 276060
rect 306984 276020 306990 276032
rect 534258 276020 534264 276032
rect 534316 276020 534322 276072
rect 313642 275952 313648 276004
rect 313700 275992 313706 276004
rect 558178 275992 558184 276004
rect 313700 275964 558184 275992
rect 313700 275952 313706 275964
rect 558178 275952 558184 275964
rect 558236 275952 558242 276004
rect 292172 275896 295840 275924
rect 292172 275884 292178 275896
rect 295886 275476 295892 275528
rect 295944 275516 295950 275528
rect 341794 275516 341800 275528
rect 295944 275488 341800 275516
rect 295944 275476 295950 275488
rect 341794 275476 341800 275488
rect 341852 275476 341858 275528
rect 218330 275408 218336 275460
rect 218388 275448 218394 275460
rect 306742 275448 306748 275460
rect 218388 275420 306748 275448
rect 218388 275408 218394 275420
rect 306742 275408 306748 275420
rect 306800 275408 306806 275460
rect 73522 275340 73528 275392
rect 73580 275380 73586 275392
rect 275830 275380 275836 275392
rect 73580 275352 275836 275380
rect 73580 275340 73586 275352
rect 275830 275340 275836 275352
rect 275888 275380 275894 275392
rect 365714 275380 365720 275392
rect 275888 275352 365720 275380
rect 275888 275340 275894 275352
rect 365714 275340 365720 275352
rect 365772 275340 365778 275392
rect 49970 275272 49976 275324
rect 50028 275312 50034 275324
rect 295886 275312 295892 275324
rect 50028 275284 295892 275312
rect 50028 275272 50034 275284
rect 295886 275272 295892 275284
rect 295944 275272 295950 275324
rect 306742 275272 306748 275324
rect 306800 275312 306806 275324
rect 510154 275312 510160 275324
rect 306800 275284 510160 275312
rect 306800 275272 306806 275284
rect 510154 275272 510160 275284
rect 510212 275272 510218 275324
rect 289998 272416 290004 272468
rect 290056 272456 290062 272468
rect 290642 272456 290648 272468
rect 290056 272428 290648 272456
rect 290056 272416 290062 272428
rect 290642 272416 290648 272428
rect 290700 272456 290706 272468
rect 560846 272456 560852 272468
rect 290700 272428 560852 272456
rect 290700 272416 290706 272428
rect 560846 272416 560852 272428
rect 560904 272416 560910 272468
rect 27246 272348 27252 272400
rect 27304 272388 27310 272400
rect 313918 272388 313924 272400
rect 27304 272360 313924 272388
rect 27304 272348 27310 272360
rect 313918 272348 313924 272360
rect 313976 272348 313982 272400
rect 24946 272008 24952 272060
rect 25004 272048 25010 272060
rect 276014 272048 276020 272060
rect 25004 272020 276020 272048
rect 25004 272008 25010 272020
rect 276014 272008 276020 272020
rect 276072 272008 276078 272060
rect 24762 271940 24768 271992
rect 24820 271980 24826 271992
rect 276198 271980 276204 271992
rect 24820 271952 276204 271980
rect 24820 271940 24826 271952
rect 276198 271940 276204 271952
rect 276256 271940 276262 271992
rect 310514 271940 310520 271992
rect 310572 271980 310578 271992
rect 558546 271980 558552 271992
rect 310572 271952 558552 271980
rect 310572 271940 310578 271952
rect 558546 271940 558552 271952
rect 558604 271940 558610 271992
rect 309778 271464 309784 271516
rect 309836 271504 309842 271516
rect 310514 271504 310520 271516
rect 309836 271476 310520 271504
rect 309836 271464 309842 271476
rect 310514 271464 310520 271476
rect 310572 271464 310578 271516
rect 276198 270852 276204 270904
rect 276256 270892 276262 270904
rect 286318 270892 286324 270904
rect 276256 270864 286324 270892
rect 276256 270852 276262 270864
rect 286318 270852 286324 270864
rect 286376 270852 286382 270904
rect 313918 270784 313924 270836
rect 313976 270824 313982 270836
rect 315022 270824 315028 270836
rect 313976 270796 315028 270824
rect 313976 270784 313982 270796
rect 315022 270784 315028 270796
rect 315080 270784 315086 270836
rect 269022 238416 269028 238468
rect 269080 238456 269086 238468
rect 290642 238456 290648 238468
rect 269080 238428 290648 238456
rect 269080 238416 269086 238428
rect 290642 238416 290648 238428
rect 290700 238416 290706 238468
rect 286318 235492 286324 235544
rect 286376 235532 286382 235544
rect 315022 235532 315028 235544
rect 286376 235504 315028 235532
rect 286376 235492 286382 235504
rect 315022 235492 315028 235504
rect 315080 235492 315086 235544
rect 558546 209108 558552 209160
rect 558604 209148 558610 209160
rect 560754 209148 560760 209160
rect 558604 209120 560760 209148
rect 558604 209108 558610 209120
rect 560754 209108 560760 209120
rect 560812 209108 560818 209160
rect 268010 203056 268016 203108
rect 268068 203096 268074 203108
rect 309778 203096 309784 203108
rect 268068 203068 309784 203096
rect 268068 203056 268074 203068
rect 309778 203056 309784 203068
rect 309836 203056 309842 203108
rect 276014 202308 276020 202360
rect 276072 202348 276078 202360
rect 282638 202348 282644 202360
rect 276072 202320 282644 202348
rect 276072 202308 276078 202320
rect 282638 202308 282644 202320
rect 282696 202308 282702 202360
rect 282638 200132 282644 200184
rect 282696 200172 282702 200184
rect 315022 200172 315028 200184
rect 282696 200144 315028 200172
rect 282696 200132 282702 200144
rect 315022 200132 315028 200144
rect 315080 200132 315086 200184
rect 269298 130228 269304 130280
rect 269356 130268 269362 130280
rect 270586 130268 270592 130280
rect 269356 130240 270592 130268
rect 269356 130228 269362 130240
rect 270586 130228 270592 130240
rect 270644 130268 270650 130280
rect 286594 130268 286600 130280
rect 270644 130240 286600 130268
rect 270644 130228 270650 130240
rect 286594 130228 286600 130240
rect 286652 130228 286658 130280
rect 286594 126624 286600 126676
rect 286652 126664 286658 126676
rect 286652 126636 287100 126664
rect 286652 126624 286658 126636
rect 287072 126596 287100 126636
rect 292850 126596 292856 126608
rect 287072 126568 292856 126596
rect 292850 126556 292856 126568
rect 292908 126556 292914 126608
rect 292942 122204 292948 122256
rect 293000 122244 293006 122256
rect 297358 122244 297364 122256
rect 293000 122216 297364 122244
rect 293000 122204 293006 122216
rect 297358 122204 297364 122216
rect 297416 122204 297422 122256
rect 297358 118124 297364 118176
rect 297416 118164 297422 118176
rect 298830 118164 298836 118176
rect 297416 118136 298836 118164
rect 297416 118124 297422 118136
rect 298830 118124 298836 118136
rect 298888 118124 298894 118176
rect 558454 116288 558460 116340
rect 558512 116328 558518 116340
rect 558638 116328 558644 116340
rect 558512 116300 558644 116328
rect 558512 116288 558518 116300
rect 558638 116288 558644 116300
rect 558696 116288 558702 116340
rect 298830 115948 298836 116000
rect 298888 115988 298894 116000
rect 300946 115988 300952 116000
rect 298888 115960 300952 115988
rect 298888 115948 298894 115960
rect 300946 115948 300952 115960
rect 301004 115948 301010 116000
rect 558546 113336 558552 113348
rect 558507 113308 558552 113336
rect 558546 113296 558552 113308
rect 558604 113296 558610 113348
rect 300946 108944 300952 108996
rect 301004 108984 301010 108996
rect 301004 108956 301820 108984
rect 301004 108944 301010 108956
rect 301792 108916 301820 108956
rect 303246 108916 303252 108928
rect 301792 108888 303252 108916
rect 303246 108876 303252 108888
rect 303304 108876 303310 108928
rect 558549 105995 558607 106001
rect 558549 105961 558561 105995
rect 558595 105992 558607 105995
rect 558730 105992 558736 106004
rect 558595 105964 558736 105992
rect 558595 105961 558607 105964
rect 558549 105955 558607 105961
rect 558730 105952 558736 105964
rect 558788 105952 558794 106004
rect 303246 102960 303252 103012
rect 303304 103000 303310 103012
rect 304902 103000 304908 103012
rect 303304 102972 304908 103000
rect 303304 102960 303310 102972
rect 304902 102960 304908 102972
rect 304960 102960 304966 103012
rect 558730 103000 558736 103012
rect 558691 102972 558736 103000
rect 558730 102960 558736 102972
rect 558788 102960 558794 103012
rect 304902 98540 304908 98592
rect 304960 98580 304966 98592
rect 308214 98580 308220 98592
rect 304960 98552 308220 98580
rect 304960 98540 304966 98552
rect 308214 98540 308220 98552
rect 308272 98540 308278 98592
rect 308214 96636 308220 96688
rect 308272 96676 308278 96688
rect 310606 96676 310612 96688
rect 308272 96648 310612 96676
rect 308272 96636 308278 96648
rect 310606 96636 310612 96648
rect 310664 96636 310670 96688
rect 269298 94868 269304 94920
rect 269356 94908 269362 94920
rect 286226 94908 286232 94920
rect 269356 94880 286232 94908
rect 269356 94868 269362 94880
rect 286226 94868 286232 94880
rect 286284 94868 286290 94920
rect 558733 92803 558791 92809
rect 558733 92769 558745 92803
rect 558779 92800 558791 92803
rect 558822 92800 558828 92812
rect 558779 92772 558828 92800
rect 558779 92769 558791 92772
rect 558733 92763 558791 92769
rect 558822 92760 558828 92772
rect 558880 92760 558886 92812
rect 299566 91264 299572 91316
rect 299624 91304 299630 91316
rect 315022 91304 315028 91316
rect 299624 91276 315028 91304
rect 299624 91264 299630 91276
rect 315022 91264 315028 91276
rect 315080 91264 315086 91316
rect 310606 91196 310612 91248
rect 310664 91236 310670 91248
rect 314194 91236 314200 91248
rect 310664 91208 314200 91236
rect 310664 91196 310670 91208
rect 314194 91196 314200 91208
rect 314252 91196 314258 91248
rect 558822 85524 558828 85536
rect 558748 85496 558828 85524
rect 558748 85332 558776 85496
rect 558822 85484 558828 85496
rect 558880 85484 558886 85536
rect 558730 85280 558736 85332
rect 558788 85280 558794 85332
rect 314194 82356 314200 82408
rect 314252 82396 314258 82408
rect 316402 82396 316408 82408
rect 314252 82368 316408 82396
rect 314252 82356 314258 82368
rect 316402 82356 316408 82368
rect 316460 82356 316466 82408
rect 316402 77256 316408 77308
rect 316460 77296 316466 77308
rect 319806 77296 319812 77308
rect 316460 77268 319812 77296
rect 316460 77256 316466 77268
rect 319806 77256 319812 77268
rect 319864 77256 319870 77308
rect 24946 75964 24952 76016
rect 25004 76004 25010 76016
rect 299566 76004 299572 76016
rect 25004 75976 299572 76004
rect 25004 75964 25010 75976
rect 299566 75964 299572 75976
rect 299624 75964 299630 76016
rect 319806 75964 319812 76016
rect 319864 76004 319870 76016
rect 558730 76004 558736 76016
rect 319864 75976 558736 76004
rect 319864 75964 319870 75976
rect 558730 75964 558736 75976
rect 558788 75964 558794 76016
rect 286226 75896 286232 75948
rect 286284 75936 286290 75948
rect 560846 75936 560852 75948
rect 286284 75908 560852 75936
rect 286284 75896 286290 75908
rect 560846 75896 560852 75908
rect 560904 75896 560910 75948
rect 313734 72292 313740 72344
rect 313792 72332 313798 72344
rect 313792 72304 313872 72332
rect 313792 72292 313798 72304
rect 313550 72196 313556 72208
rect 313463 72168 313556 72196
rect 313550 72156 313556 72168
rect 313608 72196 313614 72208
rect 313734 72196 313740 72208
rect 313608 72168 313740 72196
rect 313608 72156 313614 72168
rect 313734 72156 313740 72168
rect 313792 72156 313798 72208
rect 39666 72088 39672 72140
rect 39724 72128 39730 72140
rect 313568 72128 313596 72156
rect 39724 72100 313596 72128
rect 313844 72128 313872 72304
rect 313918 72128 313924 72140
rect 313844 72100 313924 72128
rect 39724 72088 39730 72100
rect 313918 72088 313924 72100
rect 313976 72128 313982 72140
rect 523954 72128 523960 72140
rect 313976 72100 523960 72128
rect 313976 72088 313982 72100
rect 523954 72088 523960 72100
rect 524012 72088 524018 72140
rect 256050 72020 256056 72072
rect 256108 72060 256114 72072
rect 299474 72060 299480 72072
rect 256108 72032 299480 72060
rect 256108 72020 256114 72032
rect 299474 72020 299480 72032
rect 299532 72060 299538 72072
rect 548058 72060 548064 72072
rect 299532 72032 548064 72060
rect 299532 72020 299538 72032
rect 548058 72020 548064 72032
rect 548116 72020 548122 72072
rect 270310 71952 270316 72004
rect 270368 71992 270374 72004
rect 270678 71992 270684 72004
rect 270368 71964 270684 71992
rect 270368 71952 270374 71964
rect 270678 71952 270684 71964
rect 270736 71992 270742 72004
rect 475930 71992 475936 72004
rect 270736 71964 475936 71992
rect 270736 71952 270742 71964
rect 475930 71952 475936 71964
rect 475988 71952 475994 72004
rect 87690 71884 87696 71936
rect 87748 71924 87754 71936
rect 288434 71924 288440 71936
rect 87748 71896 288440 71924
rect 87748 71884 87754 71896
rect 288434 71884 288440 71896
rect 288492 71884 288498 71936
rect 313550 71884 313556 71936
rect 313608 71924 313614 71936
rect 313826 71924 313832 71936
rect 313608 71896 313832 71924
rect 313608 71884 313614 71896
rect 313826 71884 313832 71896
rect 313884 71924 313890 71936
rect 499850 71924 499856 71936
rect 313884 71896 499856 71924
rect 313884 71884 313890 71896
rect 499850 71884 499856 71896
rect 499908 71884 499914 71936
rect 111794 71816 111800 71868
rect 111852 71856 111858 71868
rect 264977 71859 265035 71865
rect 264977 71856 264989 71859
rect 111852 71828 264989 71856
rect 111852 71816 111858 71828
rect 264977 71825 264989 71828
rect 265023 71825 265035 71859
rect 264977 71819 265035 71825
rect 276658 71816 276664 71868
rect 276716 71856 276722 71868
rect 427722 71856 427728 71868
rect 276716 71828 427728 71856
rect 276716 71816 276722 71828
rect 427722 71816 427728 71828
rect 427780 71816 427786 71868
rect 160002 71748 160008 71800
rect 160060 71788 160066 71800
rect 273070 71788 273076 71800
rect 160060 71760 273076 71788
rect 160060 71748 160066 71760
rect 273070 71748 273076 71760
rect 273128 71748 273134 71800
rect 275186 71748 275192 71800
rect 275244 71788 275250 71800
rect 403618 71788 403624 71800
rect 275244 71760 403624 71788
rect 275244 71748 275250 71760
rect 403618 71748 403624 71760
rect 403676 71748 403682 71800
rect 208026 71680 208032 71732
rect 208084 71720 208090 71732
rect 313550 71720 313556 71732
rect 208084 71692 313556 71720
rect 208084 71680 208090 71692
rect 313550 71680 313556 71692
rect 313608 71680 313614 71732
rect 183922 71612 183928 71664
rect 183980 71652 183986 71664
rect 270310 71652 270316 71664
rect 183980 71624 270316 71652
rect 183980 71612 183986 71624
rect 270310 71612 270316 71624
rect 270368 71612 270374 71664
rect 288434 71612 288440 71664
rect 288492 71652 288498 71664
rect 379514 71652 379520 71664
rect 288492 71624 379520 71652
rect 288492 71612 288498 71624
rect 379514 71612 379520 71624
rect 379572 71612 379578 71664
rect 63770 71544 63776 71596
rect 63828 71584 63834 71596
rect 270770 71584 270776 71596
rect 63828 71556 270776 71584
rect 63828 71544 63834 71556
rect 270770 71544 270776 71556
rect 270828 71584 270834 71596
rect 355594 71584 355600 71596
rect 270828 71556 355600 71584
rect 270828 71544 270834 71556
rect 355594 71544 355600 71556
rect 355652 71544 355658 71596
rect 232130 71476 232136 71528
rect 232188 71516 232194 71528
rect 313918 71516 313924 71528
rect 232188 71488 313924 71516
rect 232188 71476 232194 71488
rect 313918 71476 313924 71488
rect 313976 71476 313982 71528
rect 135898 71408 135904 71460
rect 135956 71448 135962 71460
rect 275922 71448 275928 71460
rect 135956 71420 275928 71448
rect 135956 71408 135962 71420
rect 275922 71408 275928 71420
rect 275980 71448 275986 71460
rect 276658 71448 276664 71460
rect 275980 71420 276664 71448
rect 275980 71408 275986 71420
rect 276658 71408 276664 71420
rect 276716 71408 276722 71460
rect 313734 71408 313740 71460
rect 313792 71448 313798 71460
rect 331490 71448 331496 71460
rect 313792 71420 331496 71448
rect 313792 71408 313798 71420
rect 331490 71408 331496 71420
rect 331548 71408 331554 71460
rect 264977 71383 265035 71389
rect 264977 71349 264989 71383
rect 265023 71380 265035 71383
rect 275186 71380 275192 71392
rect 265023 71352 275192 71380
rect 265023 71349 265035 71352
rect 264977 71343 265035 71349
rect 275186 71340 275192 71352
rect 275244 71340 275250 71392
<< via1 >>
rect 8024 700612 8076 700664
rect 8208 700612 8260 700664
rect 72976 700612 73028 700664
rect 137836 700612 137888 700664
rect 202788 700612 202840 700664
rect 267648 700612 267700 700664
rect 332508 700612 332560 700664
rect 397460 700612 397512 700664
rect 462320 700612 462372 700664
rect 527180 700612 527232 700664
rect 24308 700544 24360 700596
rect 24952 700544 25004 700596
rect 218980 700000 219032 700052
rect 272984 700000 273036 700052
rect 295800 700000 295852 700052
rect 429844 700000 429896 700052
rect 154120 699932 154172 699984
rect 268568 699932 268620 699984
rect 304632 699932 304684 699984
rect 494796 699932 494848 699984
rect 527180 699932 527232 699984
rect 579896 699932 579948 699984
rect 89168 699864 89220 699916
rect 277400 699864 277452 699916
rect 288440 699864 288492 699916
rect 559656 699864 559708 699916
rect 314200 674160 314252 674212
rect 578516 674160 578568 674212
rect 2964 653488 3016 653540
rect 8024 653488 8076 653540
rect 310520 627104 310572 627156
rect 578792 627104 578844 627156
rect 193864 586440 193916 586492
rect 292764 586440 292816 586492
rect 265992 586372 266044 586424
rect 313648 586372 313700 586424
rect 242072 586304 242124 586356
rect 307484 586304 307536 586356
rect 217968 586236 218020 586288
rect 306840 586236 306892 586288
rect 307576 586236 307628 586288
rect 276664 586168 276716 586220
rect 365444 586168 365496 586220
rect 291384 586100 291436 586152
rect 341524 586100 341576 586152
rect 169760 586032 169812 586084
rect 294420 586032 294472 586084
rect 73528 585964 73580 586016
rect 275928 585964 275980 586016
rect 276664 585964 276716 586016
rect 307576 585964 307628 586016
rect 509884 585964 509936 586016
rect 49608 585896 49660 585948
rect 291384 585896 291436 585948
rect 313648 585896 313700 585948
rect 557908 585896 557960 585948
rect 26516 582360 26568 582412
rect 267096 582360 267148 582412
rect 24768 582292 24820 582344
rect 286232 582292 286284 582344
rect 319812 582292 319864 582344
rect 558644 582292 558696 582344
rect 27252 582224 27304 582276
rect 314936 582224 314988 582276
rect 318616 582224 318668 582276
rect 560852 582224 560904 582276
rect 314292 579980 314344 580032
rect 314936 579980 314988 580032
rect 317420 579912 317472 579964
rect 319812 579980 319864 580032
rect 558552 579980 558604 580032
rect 578792 579980 578844 580032
rect 24860 573996 24912 574048
rect 26516 574064 26568 574116
rect 313556 574064 313608 574116
rect 317420 574064 317472 574116
rect 311624 571140 311676 571192
rect 313556 571140 313608 571192
rect 269304 547612 269356 547664
rect 291292 547612 291344 547664
rect 286232 545300 286284 545352
rect 315028 545300 315080 545352
rect 267096 531972 267148 532024
rect 269304 531972 269356 532024
rect 269304 529932 269356 529984
rect 272340 529864 272392 529916
rect 272340 523948 272392 524000
rect 274456 523948 274508 524000
rect 558644 516604 558696 516656
rect 560024 516604 560076 516656
rect 274456 514428 274508 514480
rect 278596 514428 278648 514480
rect 278596 513272 278648 513324
rect 282552 513272 282604 513324
rect 269304 511504 269356 511556
rect 309324 511504 309376 511556
rect 282644 509328 282696 509380
rect 315028 509328 315080 509380
rect 558644 485800 558696 485852
rect 578792 485800 578844 485852
rect 558736 438676 558788 438728
rect 578792 438676 578844 438728
rect 560024 421880 560076 421932
rect 560852 421880 560904 421932
rect 269304 404812 269356 404864
rect 286324 404812 286376 404864
rect 299480 401888 299532 401940
rect 315028 401888 315080 401940
rect 558828 397468 558880 397520
rect 560024 397468 560076 397520
rect 270592 386316 270644 386368
rect 558828 386316 558880 386368
rect 24860 386248 24912 386300
rect 298836 386248 298888 386300
rect 270040 386180 270092 386232
rect 270592 386180 270644 386232
rect 298836 385908 298888 385960
rect 299480 385908 299532 385960
rect 286324 385636 286376 385688
rect 293684 385636 293736 385688
rect 560852 385636 560904 385688
rect 87696 382644 87748 382696
rect 294420 382644 294472 382696
rect 135904 382576 135956 382628
rect 276388 382576 276440 382628
rect 256056 382508 256108 382560
rect 300124 382508 300176 382560
rect 313556 382440 313608 382492
rect 331496 382440 331548 382492
rect 232136 382372 232188 382424
rect 313740 382372 313792 382424
rect 270776 382304 270828 382356
rect 355600 382304 355652 382356
rect 208032 382236 208084 382288
rect 313556 382236 313608 382288
rect 111800 382168 111852 382220
rect 274456 382168 274508 382220
rect 403624 382168 403676 382220
rect 183928 382100 183980 382152
rect 270684 382100 270736 382152
rect 475936 382100 475988 382152
rect 63776 382032 63828 382084
rect 270776 382032 270828 382084
rect 313556 382032 313608 382084
rect 313832 382032 313884 382084
rect 499856 382032 499908 382084
rect 39672 381964 39724 382016
rect 313740 381964 313792 382016
rect 523960 381964 524012 382016
rect 306840 365823 306892 365832
rect 306840 365789 306849 365823
rect 306849 365789 306883 365823
rect 306883 365789 306892 365823
rect 306840 365780 306892 365789
rect 306932 360680 306984 360732
rect 309140 359116 309192 359168
rect 310520 359116 310572 359168
rect 277400 358504 277452 358556
rect 292580 358504 292632 358556
rect 3792 358436 3844 358488
rect 278412 358436 278464 358488
rect 294972 358436 295024 358488
rect 295800 358436 295852 358488
rect 3700 358368 3752 358420
rect 280804 358368 280856 358420
rect 273076 357688 273128 357740
rect 311348 357688 311400 357740
rect 270408 354016 270460 354068
rect 579344 354016 579396 354068
rect 270500 353948 270552 354000
rect 579160 353948 579212 354000
rect 314016 344360 314068 344412
rect 558644 344360 558696 344412
rect 314016 341436 314068 341488
rect 579252 341436 579304 341488
rect 268568 339940 268620 339992
rect 270224 339940 270276 339992
rect 3976 332596 4028 332648
rect 269396 332596 269448 332648
rect 24860 328244 24912 328296
rect 269396 328244 269448 328296
rect 24952 325252 25004 325304
rect 269396 325252 269448 325304
rect 313648 323892 313700 323944
rect 314016 323892 314068 323944
rect 313648 323756 313700 323808
rect 558552 323756 558604 323808
rect 3608 317908 3660 317960
rect 311532 317908 311584 317960
rect 309140 314712 309192 314764
rect 310520 314712 310572 314764
rect 3884 313488 3936 313540
rect 304356 313488 304408 313540
rect 283196 313420 283248 313472
rect 558736 313420 558788 313472
rect 272984 313352 273036 313404
rect 297364 313352 297416 313404
rect 98552 312740 98604 312792
rect 278596 312740 278648 312792
rect 306748 309136 306800 309188
rect 307116 309136 307168 309188
rect 306564 298732 306616 298784
rect 306840 298732 306892 298784
rect 306748 281120 306800 281172
rect 306932 281120 306984 281172
rect 98000 276700 98052 276752
rect 98552 276700 98604 276752
rect 194232 276360 194284 276412
rect 266360 276292 266412 276344
rect 313648 276292 313700 276344
rect 242440 276224 242492 276276
rect 306932 276224 306984 276276
rect 295156 276156 295208 276208
rect 461952 276156 462004 276208
rect 170128 275952 170180 276004
rect 292120 275884 292172 275936
rect 486056 276088 486108 276140
rect 306932 276020 306984 276072
rect 534264 276020 534316 276072
rect 313648 275952 313700 276004
rect 558184 275952 558236 276004
rect 295892 275476 295944 275528
rect 341800 275476 341852 275528
rect 218336 275408 218388 275460
rect 306748 275408 306800 275460
rect 73528 275340 73580 275392
rect 275836 275340 275888 275392
rect 365720 275340 365772 275392
rect 49976 275272 50028 275324
rect 295892 275272 295944 275324
rect 306748 275272 306800 275324
rect 510160 275272 510212 275324
rect 290004 272416 290056 272468
rect 290648 272416 290700 272468
rect 560852 272416 560904 272468
rect 27252 272348 27304 272400
rect 313924 272348 313976 272400
rect 24952 272008 25004 272060
rect 276020 272008 276072 272060
rect 24768 271940 24820 271992
rect 276204 271940 276256 271992
rect 310520 271940 310572 271992
rect 558552 271940 558604 271992
rect 309784 271464 309836 271516
rect 310520 271464 310572 271516
rect 276204 270852 276256 270904
rect 286324 270852 286376 270904
rect 313924 270784 313976 270836
rect 315028 270784 315080 270836
rect 269028 238416 269080 238468
rect 290648 238416 290700 238468
rect 286324 235492 286376 235544
rect 315028 235492 315080 235544
rect 558552 209108 558604 209160
rect 560760 209108 560812 209160
rect 268016 203056 268068 203108
rect 309784 203056 309836 203108
rect 276020 202308 276072 202360
rect 282644 202308 282696 202360
rect 282644 200132 282696 200184
rect 315028 200132 315080 200184
rect 269304 130228 269356 130280
rect 270592 130228 270644 130280
rect 286600 130228 286652 130280
rect 286600 126624 286652 126676
rect 292856 126556 292908 126608
rect 292948 122204 293000 122256
rect 297364 122204 297416 122256
rect 297364 118124 297416 118176
rect 298836 118124 298888 118176
rect 558460 116288 558512 116340
rect 558644 116288 558696 116340
rect 298836 115948 298888 116000
rect 300952 115948 301004 116000
rect 558552 113339 558604 113348
rect 558552 113305 558561 113339
rect 558561 113305 558595 113339
rect 558595 113305 558604 113339
rect 558552 113296 558604 113305
rect 300952 108944 301004 108996
rect 303252 108876 303304 108928
rect 558736 105952 558788 106004
rect 303252 102960 303304 103012
rect 304908 102960 304960 103012
rect 558736 103003 558788 103012
rect 558736 102969 558745 103003
rect 558745 102969 558779 103003
rect 558779 102969 558788 103003
rect 558736 102960 558788 102969
rect 304908 98540 304960 98592
rect 308220 98540 308272 98592
rect 308220 96636 308272 96688
rect 310612 96636 310664 96688
rect 269304 94868 269356 94920
rect 286232 94868 286284 94920
rect 558828 92760 558880 92812
rect 299572 91264 299624 91316
rect 315028 91264 315080 91316
rect 310612 91196 310664 91248
rect 314200 91196 314252 91248
rect 558828 85484 558880 85536
rect 558736 85280 558788 85332
rect 314200 82356 314252 82408
rect 316408 82356 316460 82408
rect 316408 77256 316460 77308
rect 319812 77256 319864 77308
rect 24952 75964 25004 76016
rect 299572 75964 299624 76016
rect 319812 75964 319864 76016
rect 558736 75964 558788 76016
rect 286232 75896 286284 75948
rect 560852 75896 560904 75948
rect 313740 72292 313792 72344
rect 313556 72156 313608 72208
rect 313740 72156 313792 72208
rect 39672 72088 39724 72140
rect 313924 72088 313976 72140
rect 523960 72088 524012 72140
rect 256056 72020 256108 72072
rect 299480 72020 299532 72072
rect 548064 72020 548116 72072
rect 270316 71952 270368 72004
rect 270684 71952 270736 72004
rect 475936 71952 475988 72004
rect 87696 71884 87748 71936
rect 288440 71884 288492 71936
rect 313556 71884 313608 71936
rect 313832 71884 313884 71936
rect 499856 71884 499908 71936
rect 111800 71816 111852 71868
rect 276664 71816 276716 71868
rect 427728 71816 427780 71868
rect 160008 71748 160060 71800
rect 273076 71748 273128 71800
rect 275192 71748 275244 71800
rect 403624 71748 403676 71800
rect 208032 71680 208084 71732
rect 313556 71680 313608 71732
rect 183928 71612 183980 71664
rect 270316 71612 270368 71664
rect 288440 71612 288492 71664
rect 379520 71612 379572 71664
rect 63776 71544 63828 71596
rect 270776 71544 270828 71596
rect 355600 71544 355652 71596
rect 232136 71476 232188 71528
rect 313924 71476 313976 71528
rect 135904 71408 135956 71460
rect 275928 71408 275980 71460
rect 276664 71408 276716 71460
rect 313740 71408 313792 71460
rect 331496 71408 331548 71460
rect 275192 71340 275244 71392
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 8128 703474 8156 703520
rect 8128 703446 8248 703474
rect 8220 700670 8248 703446
rect 8024 700664 8076 700670
rect 8024 700606 8076 700612
rect 8208 700664 8260 700670
rect 8208 700606 8260 700612
rect 3606 667992 3662 668001
rect 3606 667927 3662 667936
rect 2962 653576 3018 653585
rect 2962 653511 2964 653520
rect 3016 653511 3018 653520
rect 2964 653482 3016 653488
rect 2976 596057 3004 653482
rect 2962 596048 3018 596057
rect 2962 595983 3018 595992
rect 2976 538665 3004 595983
rect 2962 538656 3018 538665
rect 2962 538591 3018 538600
rect 2976 481137 3004 538591
rect 2962 481128 3018 481137
rect 2962 481063 3018 481072
rect 2976 423745 3004 481063
rect 2962 423736 3018 423745
rect 2962 423671 3018 423680
rect 3620 317966 3648 667927
rect 8036 653546 8064 700606
rect 24320 700602 24348 703520
rect 72988 700670 73016 703520
rect 72976 700664 73028 700670
rect 72976 700606 73028 700612
rect 24308 700596 24360 700602
rect 24308 700538 24360 700544
rect 24952 700596 25004 700602
rect 24952 700538 25004 700544
rect 8024 653540 8076 653546
rect 8024 653482 8076 653488
rect 3698 610464 3754 610473
rect 3698 610399 3754 610408
rect 3712 609521 3740 610399
rect 3698 609512 3754 609521
rect 3698 609447 3754 609456
rect 24768 582344 24820 582350
rect 24768 582286 24820 582292
rect 3698 553072 3754 553081
rect 3698 553007 3754 553016
rect 3712 358426 3740 553007
rect 24780 545601 24808 582286
rect 24860 574048 24912 574054
rect 24860 573990 24912 573996
rect 24766 545592 24822 545601
rect 24766 545527 24822 545536
rect 24872 509969 24900 573990
rect 24858 509960 24914 509969
rect 24858 509895 24914 509904
rect 3790 495544 3846 495553
rect 3790 495479 3846 495488
rect 3804 358494 3832 495479
rect 3974 438016 4030 438025
rect 3974 437951 4030 437960
rect 3882 423736 3938 423745
rect 3882 423671 3938 423680
rect 3792 358488 3844 358494
rect 3792 358430 3844 358436
rect 3700 358420 3752 358426
rect 3700 358362 3752 358368
rect 3608 317960 3660 317966
rect 3608 317902 3660 317908
rect 3896 313546 3924 423671
rect 3988 332654 4016 437951
rect 24858 402112 24914 402121
rect 24858 402047 24914 402056
rect 24872 386306 24900 402047
rect 24860 386300 24912 386306
rect 24860 386242 24912 386248
rect 3976 332648 4028 332654
rect 3976 332590 4028 332596
rect 24860 328296 24912 328302
rect 24860 328238 24912 328244
rect 3884 313540 3936 313546
rect 3884 313482 3936 313488
rect 24768 271992 24820 271998
rect 24768 271934 24820 271940
rect 24780 234705 24808 271934
rect 24766 234696 24822 234705
rect 24766 234631 24822 234640
rect 24872 128081 24900 328238
rect 24964 325310 24992 700538
rect 89180 699922 89208 703520
rect 137848 700670 137876 703520
rect 137836 700664 137888 700670
rect 137836 700606 137888 700612
rect 154132 699990 154160 703520
rect 202800 700670 202828 703520
rect 202788 700664 202840 700670
rect 202788 700606 202840 700612
rect 218992 700058 219020 703520
rect 267660 700670 267688 703520
rect 267648 700664 267700 700670
rect 300136 700641 300164 703520
rect 332520 700670 332548 703520
rect 332508 700664 332560 700670
rect 267648 700606 267700 700612
rect 300122 700632 300178 700641
rect 332508 700606 332560 700612
rect 300122 700567 300178 700576
rect 218980 700052 219032 700058
rect 218980 699994 219032 700000
rect 272984 700052 273036 700058
rect 272984 699994 273036 700000
rect 295800 700052 295852 700058
rect 295800 699994 295852 700000
rect 154120 699984 154172 699990
rect 154120 699926 154172 699932
rect 268568 699984 268620 699990
rect 268568 699926 268620 699932
rect 89168 699916 89220 699922
rect 89168 699858 89220 699864
rect 193864 586492 193916 586498
rect 193864 586434 193916 586440
rect 169760 586084 169812 586090
rect 169760 586026 169812 586032
rect 73528 586016 73580 586022
rect 73528 585958 73580 585964
rect 49608 585948 49660 585954
rect 49608 585890 49660 585896
rect 49620 583930 49648 585890
rect 73540 583930 73568 585958
rect 169772 583930 169800 586026
rect 193876 583930 193904 586434
rect 265992 586424 266044 586430
rect 265992 586366 266044 586372
rect 242072 586356 242124 586362
rect 242072 586298 242124 586304
rect 217968 586288 218020 586294
rect 217968 586230 218020 586236
rect 217980 583930 218008 586230
rect 242084 583930 242112 586298
rect 266004 583930 266032 586366
rect 49620 583902 49680 583930
rect 73540 583902 73600 583930
rect 169772 583902 169832 583930
rect 193876 583902 193936 583930
rect 217980 583902 218040 583930
rect 242084 583902 242144 583930
rect 266004 583902 266064 583930
rect 26516 582412 26568 582418
rect 26516 582354 26568 582360
rect 267096 582412 267148 582418
rect 267096 582354 267148 582360
rect 26528 574122 26556 582354
rect 27252 582276 27304 582282
rect 27252 582218 27304 582224
rect 27264 581233 27292 582218
rect 27250 581224 27306 581233
rect 27250 581159 27306 581168
rect 26516 574116 26568 574122
rect 26516 574058 26568 574064
rect 267108 532030 267136 582354
rect 267096 532024 267148 532030
rect 267096 531966 267148 531972
rect 39376 383982 39712 384010
rect 63480 383982 63816 384010
rect 87400 383982 87736 384010
rect 111504 383982 111840 384010
rect 135608 383982 135944 384010
rect 183816 383982 183968 384010
rect 207736 383982 208072 384010
rect 231840 383982 232176 384010
rect 255944 383982 256096 384010
rect 39684 382022 39712 383982
rect 63788 382090 63816 383982
rect 87708 382702 87736 383982
rect 87696 382696 87748 382702
rect 87696 382638 87748 382644
rect 111812 382226 111840 383982
rect 135916 382634 135944 383982
rect 135904 382628 135956 382634
rect 135904 382570 135956 382576
rect 111800 382220 111852 382226
rect 111800 382162 111852 382168
rect 183940 382158 183968 383982
rect 208044 382294 208072 383982
rect 232148 382430 232176 383982
rect 256068 382566 256096 383982
rect 256056 382560 256108 382566
rect 256056 382502 256108 382508
rect 232136 382424 232188 382430
rect 232136 382366 232188 382372
rect 208032 382288 208084 382294
rect 208032 382230 208084 382236
rect 183928 382152 183980 382158
rect 183928 382094 183980 382100
rect 63776 382084 63828 382090
rect 63776 382026 63828 382032
rect 39672 382016 39724 382022
rect 39672 381958 39724 381964
rect 268580 339998 268608 699926
rect 269304 547664 269356 547670
rect 269302 547632 269304 547641
rect 269356 547632 269358 547641
rect 269302 547567 269358 547576
rect 269304 532024 269356 532030
rect 269304 531966 269356 531972
rect 269316 529990 269344 531966
rect 269304 529984 269356 529990
rect 269304 529926 269356 529932
rect 272340 529916 272392 529922
rect 272340 529858 272392 529864
rect 272352 524006 272380 529858
rect 272340 524000 272392 524006
rect 272340 523942 272392 523948
rect 269302 512000 269358 512009
rect 269302 511935 269358 511944
rect 269316 511562 269344 511935
rect 269304 511556 269356 511562
rect 269304 511498 269356 511504
rect 270038 440736 270094 440745
rect 270038 440671 270094 440680
rect 269302 405376 269358 405385
rect 269302 405311 269358 405320
rect 269316 404870 269344 405311
rect 269304 404864 269356 404870
rect 269304 404806 269356 404812
rect 270052 386238 270080 440671
rect 270592 386368 270644 386374
rect 270592 386310 270644 386316
rect 270604 386238 270632 386310
rect 270040 386232 270092 386238
rect 270040 386174 270092 386180
rect 270592 386232 270644 386238
rect 270592 386174 270644 386180
rect 270408 354068 270460 354074
rect 270408 354010 270460 354016
rect 270420 345817 270448 354010
rect 270500 354000 270552 354006
rect 270500 353942 270552 353948
rect 270406 345808 270462 345817
rect 270406 345743 270462 345752
rect 268658 341864 268714 341873
rect 268658 341799 268714 341808
rect 268568 339992 268620 339998
rect 268568 339934 268620 339940
rect 24952 325304 25004 325310
rect 24952 325246 25004 325252
rect 98552 312792 98604 312798
rect 98552 312734 98604 312740
rect 98564 276758 98592 312734
rect 98000 276752 98052 276758
rect 98000 276694 98052 276700
rect 98552 276752 98604 276758
rect 98552 276694 98604 276700
rect 73528 275392 73580 275398
rect 73528 275334 73580 275340
rect 49976 275324 50028 275330
rect 49976 275266 50028 275272
rect 49988 273578 50016 275266
rect 49680 273550 50016 273578
rect 73540 273578 73568 275334
rect 98012 273578 98040 276694
rect 194232 276412 194284 276418
rect 194232 276354 194284 276360
rect 170128 276004 170180 276010
rect 170128 275946 170180 275952
rect 170140 273578 170168 275946
rect 194244 273578 194272 276354
rect 266360 276344 266412 276350
rect 266360 276286 266412 276292
rect 242440 276276 242492 276282
rect 242440 276218 242492 276224
rect 218336 275460 218388 275466
rect 218336 275402 218388 275408
rect 218348 273578 218376 275402
rect 242452 273578 242480 276218
rect 266372 273578 266400 276286
rect 73540 273550 73600 273578
rect 97704 273550 98040 273578
rect 169832 273550 170168 273578
rect 193936 273550 194272 273578
rect 218040 273550 218376 273578
rect 242144 273550 242480 273578
rect 266064 273550 266400 273578
rect 27252 272400 27304 272406
rect 27252 272342 27304 272348
rect 24952 272060 25004 272066
rect 24952 272002 25004 272008
rect 24964 199073 24992 272002
rect 27264 270881 27292 272342
rect 27250 270872 27306 270881
rect 27250 270807 27306 270816
rect 268016 203108 268068 203114
rect 268016 203050 268068 203056
rect 268028 201793 268056 203050
rect 268014 201784 268070 201793
rect 268014 201719 268070 201728
rect 24950 199064 25006 199073
rect 24950 198999 25006 199008
rect 268672 166161 268700 341799
rect 270224 339992 270276 339998
rect 270224 339934 270276 339940
rect 270236 339697 270264 339934
rect 270222 339688 270278 339697
rect 270222 339623 270278 339632
rect 269396 332648 269448 332654
rect 269396 332590 269448 332596
rect 269408 332353 269436 332590
rect 269394 332344 269450 332353
rect 269394 332279 269450 332288
rect 269394 328400 269450 328409
rect 269394 328335 269450 328344
rect 269408 328302 269436 328335
rect 269396 328296 269448 328302
rect 269396 328238 269448 328244
rect 269396 325304 269448 325310
rect 269394 325272 269396 325281
rect 269448 325272 269450 325281
rect 269394 325207 269450 325216
rect 270512 322289 270540 353942
rect 270498 322280 270554 322289
rect 270498 322215 270554 322224
rect 270604 318345 270632 386174
rect 270776 382356 270828 382362
rect 270776 382298 270828 382304
rect 270684 382152 270736 382158
rect 270684 382094 270736 382100
rect 270696 335481 270724 382094
rect 270788 382090 270816 382298
rect 270776 382084 270828 382090
rect 270776 382026 270828 382032
rect 270788 352753 270816 382026
rect 270774 352744 270830 352753
rect 270774 352679 270830 352688
rect 270682 335472 270738 335481
rect 270682 335407 270738 335416
rect 270590 318336 270646 318345
rect 270590 318271 270646 318280
rect 269028 238468 269080 238474
rect 269028 238410 269080 238416
rect 269040 237425 269068 238410
rect 269026 237416 269082 237425
rect 269026 237351 269082 237360
rect 268658 166152 268714 166161
rect 268658 166087 268714 166096
rect 269302 130520 269358 130529
rect 269302 130455 269358 130464
rect 269316 130286 269344 130455
rect 270604 130286 270632 318271
rect 269304 130280 269356 130286
rect 269304 130222 269356 130228
rect 270592 130280 270644 130286
rect 270592 130222 270644 130228
rect 24858 128072 24914 128081
rect 24858 128007 24914 128016
rect 269302 95160 269358 95169
rect 269302 95095 269358 95104
rect 269316 94926 269344 95095
rect 269304 94920 269356 94926
rect 269304 94862 269356 94868
rect 24950 92440 25006 92449
rect 24950 92375 25006 92384
rect 24964 76022 24992 92375
rect 24952 76016 25004 76022
rect 24952 75958 25004 75964
rect 39376 73630 39712 73658
rect 63480 73630 63816 73658
rect 87400 73630 87736 73658
rect 111504 73630 111840 73658
rect 135608 73630 135944 73658
rect 159712 73630 160048 73658
rect 183816 73630 183968 73658
rect 207736 73630 208072 73658
rect 231840 73630 232176 73658
rect 255944 73630 256096 73658
rect 39684 72146 39712 73630
rect 39672 72140 39724 72146
rect 39672 72082 39724 72088
rect 63788 71602 63816 73630
rect 87708 71942 87736 73630
rect 87696 71936 87748 71942
rect 87696 71878 87748 71884
rect 111812 71874 111840 73630
rect 111800 71868 111852 71874
rect 111800 71810 111852 71816
rect 63776 71596 63828 71602
rect 63776 71538 63828 71544
rect 135916 71466 135944 73630
rect 160020 71806 160048 73630
rect 160008 71800 160060 71806
rect 160008 71742 160060 71748
rect 183940 71670 183968 73630
rect 208044 71738 208072 73630
rect 208032 71732 208084 71738
rect 208032 71674 208084 71680
rect 183928 71664 183980 71670
rect 183928 71606 183980 71612
rect 232148 71534 232176 73630
rect 256068 72078 256096 73630
rect 256056 72072 256108 72078
rect 256056 72014 256108 72020
rect 270696 72010 270724 335407
rect 270316 72004 270368 72010
rect 270316 71946 270368 71952
rect 270684 72004 270736 72010
rect 270684 71946 270736 71952
rect 270328 71670 270356 71946
rect 270316 71664 270368 71670
rect 270316 71606 270368 71612
rect 270788 71602 270816 352679
rect 272996 313410 273024 699994
rect 277400 699916 277452 699922
rect 277400 699858 277452 699864
rect 288440 699916 288492 699922
rect 288440 699858 288492 699864
rect 276664 586220 276716 586226
rect 276664 586162 276716 586168
rect 276676 586022 276704 586162
rect 275928 586016 275980 586022
rect 275928 585958 275980 585964
rect 276664 586016 276716 586022
rect 276664 585958 276716 585964
rect 274456 524000 274508 524006
rect 274456 523942 274508 523948
rect 274468 514486 274496 523942
rect 274456 514480 274508 514486
rect 274456 514422 274508 514428
rect 274456 382220 274508 382226
rect 274456 382162 274508 382168
rect 273076 357740 273128 357746
rect 273076 357682 273128 357688
rect 272984 313404 273036 313410
rect 272984 313346 273036 313352
rect 273088 71806 273116 357682
rect 274468 354929 274496 382162
rect 275940 354929 275968 585958
rect 276388 382628 276440 382634
rect 276388 382570 276440 382576
rect 276400 382129 276428 382570
rect 276386 382120 276442 382129
rect 276386 382055 276442 382064
rect 277412 358562 277440 699858
rect 286232 582344 286284 582350
rect 286232 582286 286284 582292
rect 286244 545358 286272 582286
rect 286232 545352 286284 545358
rect 286232 545294 286284 545300
rect 278596 514480 278648 514486
rect 278596 514422 278648 514428
rect 278608 513330 278636 514422
rect 278596 513324 278648 513330
rect 278596 513266 278648 513272
rect 282552 513324 282604 513330
rect 282552 513266 282604 513272
rect 282564 509402 282592 513266
rect 282564 509386 282684 509402
rect 282564 509380 282696 509386
rect 282564 509374 282644 509380
rect 282644 509322 282696 509328
rect 282656 359417 282684 509322
rect 282642 359408 282698 359417
rect 282642 359343 282698 359352
rect 277400 358556 277452 358562
rect 277400 358498 277452 358504
rect 278412 358488 278464 358494
rect 278412 358430 278464 358436
rect 278424 355436 278452 358430
rect 280804 358420 280856 358426
rect 280804 358362 280856 358368
rect 280816 355436 280844 358362
rect 282656 355314 282684 359343
rect 286244 359281 286272 545294
rect 286324 404864 286376 404870
rect 286324 404806 286376 404812
rect 286336 385694 286364 404806
rect 286324 385688 286376 385694
rect 286324 385630 286376 385636
rect 285586 359272 285642 359281
rect 285586 359207 285642 359216
rect 286230 359272 286286 359281
rect 286230 359207 286286 359216
rect 285600 355436 285628 359207
rect 288452 355314 288480 699858
rect 292764 586492 292816 586498
rect 292764 586434 292816 586440
rect 291384 586152 291436 586158
rect 292776 586129 292804 586434
rect 294418 586256 294474 586265
rect 294418 586191 294474 586200
rect 291384 586094 291436 586100
rect 292762 586120 292818 586129
rect 291396 585954 291424 586094
rect 294432 586090 294460 586191
rect 292762 586055 292818 586064
rect 294420 586084 294472 586090
rect 294420 586026 294472 586032
rect 291384 585948 291436 585954
rect 291384 585890 291436 585896
rect 291292 547664 291344 547670
rect 291292 547606 291344 547612
rect 291304 546825 291332 547606
rect 291290 546816 291346 546825
rect 291290 546751 291346 546760
rect 282656 355286 283222 355314
rect 287822 355286 288480 355314
rect 291396 354929 291424 585890
rect 293684 385688 293736 385694
rect 293684 385630 293736 385636
rect 293696 384305 293724 385630
rect 293682 384296 293738 384305
rect 293682 384231 293738 384240
rect 294420 382696 294472 382702
rect 294420 382638 294472 382644
rect 294432 382265 294460 382638
rect 294418 382256 294474 382265
rect 294418 382191 294474 382200
rect 292580 358556 292632 358562
rect 292580 358498 292632 358504
rect 292592 355436 292620 358498
rect 295812 358494 295840 699994
rect 304632 699984 304684 699990
rect 364996 699961 365024 703520
rect 397472 700670 397500 703520
rect 397460 700664 397512 700670
rect 397460 700606 397512 700612
rect 429856 700058 429884 703520
rect 462332 700670 462360 703520
rect 462320 700664 462372 700670
rect 462320 700606 462372 700612
rect 429844 700052 429896 700058
rect 429844 699994 429896 700000
rect 494808 699990 494836 703520
rect 527192 700670 527220 703520
rect 527180 700664 527232 700670
rect 527180 700606 527232 700612
rect 527192 699990 527220 700606
rect 494796 699984 494848 699990
rect 304632 699926 304684 699932
rect 364982 699952 365038 699961
rect 299480 401940 299532 401946
rect 299480 401882 299532 401888
rect 298836 386300 298888 386306
rect 298836 386242 298888 386248
rect 298848 385966 298876 386242
rect 299492 385966 299520 401882
rect 298836 385960 298888 385966
rect 298836 385902 298888 385908
rect 299480 385960 299532 385966
rect 299480 385902 299532 385908
rect 294972 358488 295024 358494
rect 294972 358430 295024 358436
rect 295800 358488 295852 358494
rect 295800 358430 295852 358436
rect 294984 355436 295012 358430
rect 274086 354920 274142 354929
rect 273838 354878 274086 354906
rect 274086 354855 274142 354864
rect 274454 354920 274510 354929
rect 274454 354855 274510 354864
rect 275926 354920 275982 354929
rect 290462 354920 290518 354929
rect 275982 354878 276046 354906
rect 290214 354878 290462 354906
rect 275926 354855 275982 354864
rect 290462 354855 290518 354864
rect 291382 354920 291438 354929
rect 297638 354920 297694 354929
rect 297390 354878 297638 354906
rect 291382 354855 291438 354864
rect 298848 354906 298876 385902
rect 300124 382560 300176 382566
rect 300124 382502 300176 382508
rect 300136 381993 300164 382502
rect 300122 381984 300178 381993
rect 300122 381919 300178 381928
rect 300136 381313 300164 381919
rect 300122 381304 300178 381313
rect 300122 381239 300178 381248
rect 304644 355450 304672 699926
rect 494796 699926 494848 699932
rect 527180 699984 527232 699990
rect 527180 699926 527232 699932
rect 559668 699922 559696 703520
rect 579896 699984 579948 699990
rect 579896 699926 579948 699932
rect 364982 699887 365038 699896
rect 559656 699916 559708 699922
rect 559656 699858 559708 699864
rect 579908 698057 579936 699926
rect 579894 698048 579950 698057
rect 579894 697983 579950 697992
rect 578514 674656 578570 674665
rect 578514 674591 578570 674600
rect 578528 674218 578556 674591
rect 314200 674212 314252 674218
rect 314200 674154 314252 674160
rect 578516 674212 578568 674218
rect 578516 674154 578568 674160
rect 310520 627156 310572 627162
rect 310520 627098 310572 627104
rect 307484 586356 307536 586362
rect 307484 586298 307536 586304
rect 306840 586288 306892 586294
rect 306840 586230 306892 586236
rect 306852 365838 306880 586230
rect 307496 585993 307524 586298
rect 307576 586288 307628 586294
rect 307576 586230 307628 586236
rect 307588 586022 307616 586230
rect 307576 586016 307628 586022
rect 307482 585984 307538 585993
rect 307576 585958 307628 585964
rect 307482 585919 307538 585928
rect 309322 511592 309378 511601
rect 309322 511527 309324 511536
rect 309376 511527 309378 511536
rect 309324 511498 309376 511504
rect 309336 504937 309364 511498
rect 309322 504928 309378 504937
rect 309322 504863 309378 504872
rect 309966 473784 310022 473793
rect 309966 473719 310022 473728
rect 309980 463729 310008 473719
rect 309966 463720 310022 463729
rect 309966 463655 310022 463664
rect 309966 432576 310022 432585
rect 309966 432511 310022 432520
rect 309980 422521 310008 432511
rect 309966 422512 310022 422521
rect 309966 422447 310022 422456
rect 309782 412176 309838 412185
rect 309782 412111 309838 412120
rect 309796 402121 309824 412111
rect 309782 402112 309838 402121
rect 309782 402047 309838 402056
rect 309782 391504 309838 391513
rect 309782 391439 309838 391448
rect 309796 381313 309824 391439
rect 309782 381304 309838 381313
rect 309782 381239 309838 381248
rect 309414 370968 309470 370977
rect 309414 370903 309470 370912
rect 306840 365832 306892 365838
rect 306840 365774 306892 365780
rect 309428 360913 309456 370903
rect 309414 360904 309470 360913
rect 309414 360839 309470 360848
rect 306932 360732 306984 360738
rect 306932 360674 306984 360680
rect 304382 355422 304672 355450
rect 306470 355328 306526 355337
rect 306944 355314 306972 360674
rect 310532 359174 310560 627098
rect 313648 586424 313700 586430
rect 313648 586366 313700 586372
rect 313660 585954 313688 586366
rect 313648 585948 313700 585954
rect 313648 585890 313700 585896
rect 313556 574116 313608 574122
rect 313556 574058 313608 574064
rect 313568 571198 313596 574058
rect 311624 571192 311676 571198
rect 311624 571134 311676 571140
rect 313556 571192 313608 571198
rect 313556 571134 313608 571140
rect 311636 566681 311664 571134
rect 311622 566672 311678 566681
rect 311622 566607 311678 566616
rect 313556 382492 313608 382498
rect 313556 382434 313608 382440
rect 313568 382378 313596 382434
rect 313476 382350 313596 382378
rect 313476 381970 313504 382350
rect 313556 382288 313608 382294
rect 313556 382230 313608 382236
rect 313568 382090 313596 382230
rect 313556 382084 313608 382090
rect 313556 382026 313608 382032
rect 313476 381942 313596 381970
rect 309140 359168 309192 359174
rect 309140 359110 309192 359116
rect 310520 359168 310572 359174
rect 310520 359110 310572 359116
rect 309152 355436 309180 359110
rect 311348 357740 311400 357746
rect 311348 357682 311400 357688
rect 311360 355436 311388 357682
rect 306526 355286 306972 355314
rect 306470 355263 306526 355272
rect 299478 354920 299534 354929
rect 298848 354878 299478 354906
rect 297638 354855 297694 354864
rect 299534 354878 299598 354906
rect 299478 354855 299534 354864
rect 313568 347993 313596 381942
rect 313554 347984 313610 347993
rect 313554 347919 313610 347928
rect 311532 317960 311584 317966
rect 311532 317902 311584 317908
rect 311544 317121 311572 317902
rect 311530 317112 311586 317121
rect 311530 317047 311586 317056
rect 274086 316296 274142 316305
rect 273838 316254 274086 316282
rect 292854 316296 292910 316305
rect 274086 316231 274142 316240
rect 292132 316254 292854 316282
rect 290646 315752 290702 315761
rect 290646 315687 290702 315696
rect 276110 315616 276166 315625
rect 275940 315574 276110 315602
rect 275834 276720 275890 276729
rect 275834 276655 275890 276664
rect 275848 275398 275876 276655
rect 275836 275392 275888 275398
rect 275836 275334 275888 275340
rect 275190 72040 275246 72049
rect 275190 71975 275246 71984
rect 275204 71806 275232 71975
rect 273076 71800 273128 71806
rect 273076 71742 273128 71748
rect 275192 71800 275244 71806
rect 275192 71742 275244 71748
rect 270776 71596 270828 71602
rect 270776 71538 270828 71544
rect 232136 71528 232188 71534
rect 232136 71470 232188 71476
rect 135904 71460 135956 71466
rect 135904 71402 135956 71408
rect 275204 71398 275232 71742
rect 275940 71466 275968 315574
rect 290660 315602 290688 315687
rect 276166 315574 276230 315602
rect 276110 315551 276166 315560
rect 276124 315491 276152 315551
rect 278608 312798 278636 315588
rect 280816 313177 280844 315588
rect 283208 313478 283236 315588
rect 283196 313472 283248 313478
rect 283196 313414 283248 313420
rect 280802 313168 280858 313177
rect 280802 313103 280858 313112
rect 278596 312792 278648 312798
rect 278596 312734 278648 312740
rect 285600 312089 285628 315588
rect 287992 313449 288020 315588
rect 290016 315574 290688 315602
rect 287978 313440 288034 313449
rect 287978 313375 288034 313384
rect 288438 313440 288494 313449
rect 288438 313375 288494 313384
rect 285586 312080 285642 312089
rect 285586 312015 285642 312024
rect 286230 312080 286286 312089
rect 286230 312015 286286 312024
rect 276018 272232 276074 272241
rect 276018 272167 276074 272176
rect 276032 272066 276060 272167
rect 276202 272096 276258 272105
rect 276020 272060 276072 272066
rect 276202 272031 276258 272040
rect 276020 272002 276072 272008
rect 276032 202366 276060 272002
rect 276216 271998 276244 272031
rect 276204 271992 276256 271998
rect 276204 271934 276256 271940
rect 276216 270910 276244 271934
rect 276204 270904 276256 270910
rect 276204 270846 276256 270852
rect 276020 202360 276072 202366
rect 276020 202302 276072 202308
rect 282644 202360 282696 202366
rect 282644 202302 282696 202308
rect 282656 200190 282684 202302
rect 282644 200184 282696 200190
rect 282644 200126 282696 200132
rect 286244 94926 286272 312015
rect 286324 270904 286376 270910
rect 286324 270846 286376 270852
rect 286336 235550 286364 270846
rect 286324 235544 286376 235550
rect 286324 235486 286376 235492
rect 286600 130280 286652 130286
rect 286600 130222 286652 130228
rect 286612 126682 286640 130222
rect 286600 126676 286652 126682
rect 286600 126618 286652 126624
rect 286232 94920 286284 94926
rect 286232 94862 286284 94868
rect 286244 75954 286272 94862
rect 286232 75948 286284 75954
rect 286232 75890 286284 75896
rect 288452 71942 288480 313375
rect 290016 272474 290044 315574
rect 292132 275942 292160 316254
rect 295246 316296 295302 316305
rect 294998 316254 295246 316282
rect 292854 316231 292910 316240
rect 295168 276214 295196 316254
rect 300030 316296 300086 316305
rect 295246 316231 295302 316240
rect 299492 316254 300030 316282
rect 297376 313410 297404 315588
rect 297364 313404 297416 313410
rect 297364 313346 297416 313352
rect 295156 276208 295208 276214
rect 295156 276150 295208 276156
rect 292120 275936 292172 275942
rect 292120 275878 292172 275884
rect 295892 275528 295944 275534
rect 295892 275470 295944 275476
rect 295904 275369 295932 275470
rect 295890 275360 295946 275369
rect 295890 275295 295892 275304
rect 295944 275295 295946 275304
rect 295892 275266 295944 275272
rect 290004 272468 290056 272474
rect 290004 272410 290056 272416
rect 290648 272468 290700 272474
rect 290648 272410 290700 272416
rect 290660 238474 290688 272410
rect 290648 238468 290700 238474
rect 290648 238410 290700 238416
rect 292856 126608 292908 126614
rect 292856 126550 292908 126556
rect 292868 125066 292896 126550
rect 292868 125038 292988 125066
rect 292960 122262 292988 125038
rect 292948 122256 293000 122262
rect 292948 122198 293000 122204
rect 297364 122256 297416 122262
rect 297364 122198 297416 122204
rect 297376 118182 297404 122198
rect 297364 118176 297416 118182
rect 297364 118118 297416 118124
rect 298836 118176 298888 118182
rect 298836 118118 298888 118124
rect 298848 116006 298876 118118
rect 298836 116000 298888 116006
rect 298836 115942 298888 115948
rect 299492 72078 299520 316254
rect 300030 316231 300086 316240
rect 309414 316296 309470 316305
rect 309414 316231 309470 316240
rect 306654 315616 306710 315625
rect 304368 313546 304396 315588
rect 309428 315602 309456 316231
rect 306710 315588 306774 315602
rect 309166 315588 309456 315602
rect 306710 315574 306788 315588
rect 306654 315551 306710 315560
rect 304356 313540 304408 313546
rect 304356 313482 304408 313488
rect 306760 309194 306788 315574
rect 309152 315574 309456 315588
rect 309152 314770 309180 315574
rect 309140 314764 309192 314770
rect 309140 314706 309192 314712
rect 310520 314764 310572 314770
rect 310520 314706 310572 314712
rect 306748 309188 306800 309194
rect 306748 309130 306800 309136
rect 307116 309188 307168 309194
rect 307116 309130 307168 309136
rect 307128 301730 307156 309130
rect 306852 301702 307156 301730
rect 306852 298790 306880 301702
rect 306564 298784 306616 298790
rect 306564 298726 306616 298732
rect 306840 298784 306892 298790
rect 306840 298726 306892 298732
rect 306576 288561 306604 298726
rect 306562 288552 306618 288561
rect 306562 288487 306618 288496
rect 306746 288552 306802 288561
rect 306746 288487 306802 288496
rect 306760 281178 306788 288487
rect 306748 281172 306800 281178
rect 306748 281114 306800 281120
rect 306932 281172 306984 281178
rect 306932 281114 306984 281120
rect 306746 276720 306802 276729
rect 306746 276655 306802 276664
rect 306760 275466 306788 276655
rect 306944 276282 306972 281114
rect 306932 276276 306984 276282
rect 306932 276218 306984 276224
rect 306944 276078 306972 276218
rect 306932 276072 306984 276078
rect 306932 276014 306984 276020
rect 306748 275460 306800 275466
rect 306748 275402 306800 275408
rect 306760 275330 306788 275402
rect 306748 275324 306800 275330
rect 306748 275266 306800 275272
rect 310532 271998 310560 314706
rect 310520 271992 310572 271998
rect 310520 271934 310572 271940
rect 310532 271522 310560 271934
rect 309784 271516 309836 271522
rect 309784 271458 309836 271464
rect 310520 271516 310572 271522
rect 310520 271458 310572 271464
rect 309796 203114 309824 271458
rect 309784 203108 309836 203114
rect 309784 203050 309836 203056
rect 300952 116000 301004 116006
rect 300952 115942 301004 115948
rect 300964 109002 300992 115942
rect 300952 108996 301004 109002
rect 300952 108938 301004 108944
rect 303252 108928 303304 108934
rect 303252 108870 303304 108876
rect 303264 103018 303292 108870
rect 303252 103012 303304 103018
rect 303252 102954 303304 102960
rect 304908 103012 304960 103018
rect 304908 102954 304960 102960
rect 304920 98598 304948 102954
rect 304908 98592 304960 98598
rect 304908 98534 304960 98540
rect 308220 98592 308272 98598
rect 308220 98534 308272 98540
rect 308232 96694 308260 98534
rect 308220 96688 308272 96694
rect 308220 96630 308272 96636
rect 310612 96688 310664 96694
rect 310612 96630 310664 96636
rect 299570 92712 299626 92721
rect 299570 92647 299626 92656
rect 299584 91322 299612 92647
rect 299572 91316 299624 91322
rect 299572 91258 299624 91264
rect 299584 76022 299612 91258
rect 310624 91254 310652 96630
rect 310612 91248 310664 91254
rect 310612 91190 310664 91196
rect 299572 76016 299624 76022
rect 299572 75958 299624 75964
rect 313568 72214 313596 347919
rect 313660 323950 313688 585890
rect 313740 382424 313792 382430
rect 313740 382366 313792 382372
rect 313752 382022 313780 382366
rect 313832 382084 313884 382090
rect 313832 382026 313884 382032
rect 313740 382016 313792 382022
rect 313740 381958 313792 381964
rect 313752 330721 313780 381958
rect 313738 330712 313794 330721
rect 313738 330647 313794 330656
rect 313648 323944 313700 323950
rect 313648 323886 313700 323892
rect 313648 323808 313700 323814
rect 313648 323750 313700 323756
rect 313660 323649 313688 323750
rect 313646 323640 313702 323649
rect 313646 323575 313702 323584
rect 313646 320648 313702 320657
rect 313646 320583 313702 320592
rect 313660 276350 313688 320583
rect 313648 276344 313700 276350
rect 313648 276286 313700 276292
rect 313660 276010 313688 276286
rect 313648 276004 313700 276010
rect 313648 275946 313700 275952
rect 313752 72350 313780 330647
rect 313844 327049 313872 382026
rect 313922 351792 313978 351801
rect 313922 351727 313978 351736
rect 313830 327040 313886 327049
rect 313830 326975 313886 326984
rect 313740 72344 313792 72350
rect 313740 72286 313792 72292
rect 313556 72208 313608 72214
rect 313556 72150 313608 72156
rect 313740 72208 313792 72214
rect 313740 72150 313792 72156
rect 299480 72072 299532 72078
rect 299480 72014 299532 72020
rect 288440 71936 288492 71942
rect 288440 71878 288492 71884
rect 313556 71936 313608 71942
rect 313556 71878 313608 71884
rect 276664 71868 276716 71874
rect 276664 71810 276716 71816
rect 276676 71466 276704 71810
rect 288452 71670 288480 71878
rect 313568 71738 313596 71878
rect 313556 71732 313608 71738
rect 313556 71674 313608 71680
rect 288440 71664 288492 71670
rect 288440 71606 288492 71612
rect 313752 71466 313780 72150
rect 313844 71942 313872 326975
rect 313936 272406 313964 351727
rect 314014 344448 314070 344457
rect 314014 344383 314016 344392
rect 314068 344383 314070 344392
rect 314016 344354 314068 344360
rect 314016 341488 314068 341494
rect 314016 341430 314068 341436
rect 314028 341193 314056 341430
rect 314014 341184 314070 341193
rect 314014 341119 314070 341128
rect 314212 338065 314240 674154
rect 579908 651137 579936 697983
rect 579894 651128 579950 651137
rect 579894 651063 579950 651072
rect 578790 627736 578846 627745
rect 578790 627671 578846 627680
rect 578804 627162 578832 627671
rect 578792 627156 578844 627162
rect 578792 627098 578844 627104
rect 579908 604217 579936 651063
rect 579894 604208 579950 604217
rect 579894 604143 579950 604152
rect 461674 586256 461730 586265
rect 365444 586220 365496 586226
rect 461674 586191 461730 586200
rect 365444 586162 365496 586168
rect 341524 586152 341576 586158
rect 341524 586094 341576 586100
rect 341536 583930 341564 586094
rect 365456 583930 365484 586162
rect 461688 583930 461716 586191
rect 485778 586120 485834 586129
rect 485778 586055 485834 586064
rect 485792 583930 485820 586055
rect 509884 586016 509936 586022
rect 509884 585958 509936 585964
rect 533986 585984 534042 585993
rect 509896 583930 509924 585958
rect 533986 585919 534042 585928
rect 557908 585948 557960 585954
rect 534000 583930 534028 585919
rect 557908 585890 557960 585896
rect 557920 583930 557948 585890
rect 341536 583902 341826 583930
rect 365456 583902 365746 583930
rect 461688 583902 461978 583930
rect 485792 583902 486082 583930
rect 509896 583902 510186 583930
rect 534000 583902 534290 583930
rect 557920 583902 558210 583930
rect 319812 582344 319864 582350
rect 319812 582286 319864 582292
rect 558644 582344 558696 582350
rect 558644 582286 558696 582292
rect 314936 582276 314988 582282
rect 314936 582218 314988 582224
rect 318616 582276 318668 582282
rect 318616 582218 318668 582224
rect 314948 580530 314976 582218
rect 315026 580544 315082 580553
rect 314948 580502 315026 580530
rect 314948 580038 314976 580502
rect 315026 580479 315082 580488
rect 314292 580032 314344 580038
rect 314292 579974 314344 579980
rect 314936 580032 314988 580038
rect 314936 579974 314988 579980
rect 314304 351801 314332 579974
rect 317420 579964 317472 579970
rect 317420 579906 317472 579912
rect 317432 574122 317460 579906
rect 317420 574116 317472 574122
rect 317420 574058 317472 574064
rect 318628 546825 318656 582218
rect 319824 580038 319852 582286
rect 319812 580032 319864 580038
rect 319812 579974 319864 579980
rect 558552 580032 558604 580038
rect 558552 579974 558604 579980
rect 318614 546816 318670 546825
rect 318614 546751 318670 546760
rect 315028 545352 315080 545358
rect 315028 545294 315080 545300
rect 315040 545193 315068 545294
rect 315026 545184 315082 545193
rect 315026 545119 315082 545128
rect 315026 509416 315082 509425
rect 315026 509351 315028 509360
rect 315080 509351 315082 509360
rect 315028 509322 315080 509328
rect 315026 402384 315082 402393
rect 315026 402319 315082 402328
rect 315040 401946 315068 402319
rect 315028 401940 315080 401946
rect 315028 401882 315080 401888
rect 331508 382498 331536 383996
rect 331496 382492 331548 382498
rect 331496 382434 331548 382440
rect 355612 382362 355640 383996
rect 355600 382356 355652 382362
rect 355600 382298 355652 382304
rect 379532 382265 379560 383996
rect 379518 382256 379574 382265
rect 403636 382226 403664 383996
rect 379518 382191 379574 382200
rect 403624 382220 403676 382226
rect 403624 382162 403676 382168
rect 427740 382129 427768 383996
rect 475948 382158 475976 383996
rect 475936 382152 475988 382158
rect 427726 382120 427782 382129
rect 475936 382094 475988 382100
rect 499868 382090 499896 383996
rect 427726 382055 427782 382064
rect 499856 382084 499908 382090
rect 499856 382026 499908 382032
rect 523972 382022 524000 383996
rect 523960 382016 524012 382022
rect 548076 381993 548104 383996
rect 523960 381958 524012 381964
rect 548062 381984 548118 381993
rect 548062 381919 548118 381928
rect 314290 351792 314346 351801
rect 314290 351727 314346 351736
rect 314198 338056 314254 338065
rect 314198 337991 314254 338000
rect 314016 323944 314068 323950
rect 314016 323886 314068 323892
rect 314028 320657 314056 323886
rect 558564 323814 558592 579974
rect 558656 516662 558684 582286
rect 560852 582276 560904 582282
rect 560852 582218 560904 582224
rect 560864 547777 560892 582218
rect 578790 580816 578846 580825
rect 578790 580751 578846 580760
rect 578804 580038 578832 580751
rect 578792 580032 578844 580038
rect 578792 579974 578844 579980
rect 579908 557297 579936 604143
rect 579894 557288 579950 557297
rect 579894 557223 579950 557232
rect 560850 547768 560906 547777
rect 560850 547703 560906 547712
rect 579158 533896 579214 533905
rect 579158 533831 579214 533840
rect 558644 516656 558696 516662
rect 558644 516598 558696 516604
rect 560024 516656 560076 516662
rect 560024 516598 560076 516604
rect 560036 512145 560064 516598
rect 560022 512136 560078 512145
rect 560022 512071 560078 512080
rect 578790 486840 578846 486849
rect 578790 486775 578846 486784
rect 578804 485858 578832 486775
rect 558644 485852 558696 485858
rect 558644 485794 558696 485800
rect 578792 485852 578844 485858
rect 578792 485794 578844 485800
rect 558656 344418 558684 485794
rect 560850 440736 560906 440745
rect 560850 440671 560906 440680
rect 558736 438728 558788 438734
rect 558736 438670 558788 438676
rect 558644 344412 558696 344418
rect 558644 344354 558696 344360
rect 558552 323808 558604 323814
rect 558552 323750 558604 323756
rect 314014 320648 314070 320657
rect 314014 320583 314070 320592
rect 558748 313478 558776 438670
rect 560864 421938 560892 440671
rect 578790 439920 578846 439929
rect 578790 439855 578846 439864
rect 578804 438734 578832 439855
rect 578792 438728 578844 438734
rect 578792 438670 578844 438676
rect 560024 421932 560076 421938
rect 560024 421874 560076 421880
rect 560852 421932 560904 421938
rect 560852 421874 560904 421880
rect 560036 397526 560064 421874
rect 560850 405376 560906 405385
rect 560850 405311 560906 405320
rect 558828 397520 558880 397526
rect 558828 397462 558880 397468
rect 560024 397520 560076 397526
rect 560024 397462 560076 397468
rect 558840 386374 558868 397462
rect 558828 386368 558880 386374
rect 558828 386310 558880 386316
rect 560864 385694 560892 405311
rect 560852 385688 560904 385694
rect 560852 385630 560904 385636
rect 579172 354006 579200 533831
rect 579908 510377 579936 557223
rect 579894 510368 579950 510377
rect 579894 510303 579950 510312
rect 579908 463457 579936 510303
rect 579894 463448 579950 463457
rect 579894 463383 579950 463392
rect 579908 416537 579936 463383
rect 579894 416528 579950 416537
rect 579894 416463 579950 416472
rect 579908 415177 579936 416463
rect 579250 415168 579306 415177
rect 579250 415103 579306 415112
rect 579894 415168 579950 415177
rect 579894 415103 579950 415112
rect 579160 354000 579212 354006
rect 579160 353942 579212 353948
rect 579264 341494 579292 415103
rect 579342 393000 579398 393009
rect 579342 392935 579398 392944
rect 579356 354074 579384 392935
rect 579344 354068 579396 354074
rect 579344 354010 579396 354016
rect 579252 341488 579304 341494
rect 579252 341430 579304 341436
rect 558736 313472 558788 313478
rect 558736 313414 558788 313420
rect 461952 276208 462004 276214
rect 461952 276150 462004 276156
rect 341800 275528 341852 275534
rect 341800 275470 341852 275476
rect 341812 273564 341840 275470
rect 365720 275392 365772 275398
rect 365720 275334 365772 275340
rect 365732 273564 365760 275334
rect 461964 273564 461992 276150
rect 486056 276140 486108 276146
rect 486056 276082 486108 276088
rect 486068 273564 486096 276082
rect 534264 276072 534316 276078
rect 534264 276014 534316 276020
rect 510160 275324 510212 275330
rect 510160 275266 510212 275272
rect 510172 273564 510200 275266
rect 534276 273564 534304 276014
rect 558184 276004 558236 276010
rect 558184 275946 558236 275952
rect 558196 273564 558224 275946
rect 560852 272468 560904 272474
rect 560852 272410 560904 272416
rect 313924 272400 313976 272406
rect 313924 272342 313976 272348
rect 313936 270842 313964 272342
rect 558552 271992 558604 271998
rect 558552 271934 558604 271940
rect 313924 270836 313976 270842
rect 313924 270778 313976 270784
rect 315028 270836 315080 270842
rect 315028 270778 315080 270784
rect 315040 270337 315068 270778
rect 315026 270328 315082 270337
rect 315026 270263 315082 270272
rect 315028 235544 315080 235550
rect 315028 235486 315080 235492
rect 315040 234705 315068 235486
rect 315026 234696 315082 234705
rect 315026 234631 315082 234640
rect 558564 209166 558592 271934
rect 560864 237425 560892 272410
rect 560850 237416 560906 237425
rect 560850 237351 560906 237360
rect 558552 209160 558604 209166
rect 558552 209102 558604 209108
rect 560760 209160 560812 209166
rect 560760 209102 560812 209108
rect 560772 207482 560800 209102
rect 560772 207454 560892 207482
rect 560864 201793 560892 207454
rect 560850 201784 560906 201793
rect 560850 201719 560906 201728
rect 315028 200184 315080 200190
rect 315028 200126 315080 200132
rect 315040 199073 315068 200126
rect 315026 199064 315082 199073
rect 315026 198999 315082 199008
rect 558918 130520 558974 130529
rect 558748 130478 558918 130506
rect 558748 128602 558776 130478
rect 558918 130455 558974 130464
rect 558656 128574 558776 128602
rect 558656 116346 558684 128574
rect 558460 116340 558512 116346
rect 558460 116282 558512 116288
rect 558644 116340 558696 116346
rect 558644 116282 558696 116288
rect 558472 116226 558500 116282
rect 558472 116198 558592 116226
rect 558564 113354 558592 116198
rect 558552 113348 558604 113354
rect 558552 113290 558604 113296
rect 558736 106004 558788 106010
rect 558736 105946 558788 105952
rect 558748 103018 558776 105946
rect 558736 103012 558788 103018
rect 558736 102954 558788 102960
rect 560850 95160 560906 95169
rect 560850 95095 560906 95104
rect 558828 92812 558880 92818
rect 558828 92754 558880 92760
rect 315026 92440 315082 92449
rect 315026 92375 315082 92384
rect 315040 91322 315068 92375
rect 315028 91316 315080 91322
rect 315028 91258 315080 91264
rect 314200 91248 314252 91254
rect 314200 91190 314252 91196
rect 314212 82414 314240 91190
rect 558840 85542 558868 92754
rect 558828 85536 558880 85542
rect 558828 85478 558880 85484
rect 558736 85332 558788 85338
rect 558736 85274 558788 85280
rect 314200 82408 314252 82414
rect 314200 82350 314252 82356
rect 316408 82408 316460 82414
rect 316408 82350 316460 82356
rect 316420 77314 316448 82350
rect 316408 77308 316460 77314
rect 316408 77250 316460 77256
rect 319812 77308 319864 77314
rect 319812 77250 319864 77256
rect 319824 76022 319852 77250
rect 558748 76022 558776 85274
rect 319812 76016 319864 76022
rect 319812 75958 319864 75964
rect 558736 76016 558788 76022
rect 558736 75958 558788 75964
rect 560864 75954 560892 95095
rect 560852 75948 560904 75954
rect 560852 75890 560904 75896
rect 313924 72140 313976 72146
rect 313924 72082 313976 72088
rect 313832 71936 313884 71942
rect 313832 71878 313884 71884
rect 313936 71534 313964 72082
rect 313924 71528 313976 71534
rect 313924 71470 313976 71476
rect 331508 71466 331536 73644
rect 355612 71602 355640 73644
rect 379532 71670 379560 73644
rect 403636 71806 403664 73644
rect 427740 71874 427768 73644
rect 475948 72010 475976 73644
rect 475936 72004 475988 72010
rect 475936 71946 475988 71952
rect 499868 71942 499896 73644
rect 523972 72146 524000 73644
rect 523960 72140 524012 72146
rect 523960 72082 524012 72088
rect 548076 72078 548104 73644
rect 548064 72072 548116 72078
rect 548064 72014 548116 72020
rect 499856 71936 499908 71942
rect 499856 71878 499908 71884
rect 427728 71868 427780 71874
rect 427728 71810 427780 71816
rect 403624 71800 403676 71806
rect 403624 71742 403676 71748
rect 379520 71664 379572 71670
rect 379520 71606 379572 71612
rect 355600 71596 355652 71602
rect 355600 71538 355652 71544
rect 275928 71460 275980 71466
rect 275928 71402 275980 71408
rect 276664 71460 276716 71466
rect 276664 71402 276716 71408
rect 313740 71460 313792 71466
rect 313740 71402 313792 71408
rect 331496 71460 331548 71466
rect 331496 71402 331548 71408
rect 275192 71392 275244 71398
rect 275192 71334 275244 71340
rect 583390 3632 583446 3641
rect 583390 3567 583446 3576
rect 583404 480 583432 3567
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8822 -960 8934 480
rect 10018 -960 10130 480
rect 11214 -960 11326 480
rect 12410 -960 12522 480
rect 13606 -960 13718 480
rect 14802 -960 14914 480
rect 15998 -960 16110 480
rect 17194 -960 17306 480
rect 18298 -960 18410 480
rect 19494 -960 19606 480
rect 20690 -960 20802 480
rect 21886 -960 21998 480
rect 23082 -960 23194 480
rect 24278 -960 24390 480
rect 25474 -960 25586 480
rect 26670 -960 26782 480
rect 27866 -960 27978 480
rect 29062 -960 29174 480
rect 30258 -960 30370 480
rect 31454 -960 31566 480
rect 32650 -960 32762 480
rect 33846 -960 33958 480
rect 34950 -960 35062 480
rect 36146 -960 36258 480
rect 37342 -960 37454 480
rect 38538 -960 38650 480
rect 39734 -960 39846 480
rect 40930 -960 41042 480
rect 42126 -960 42238 480
rect 43322 -960 43434 480
rect 44518 -960 44630 480
rect 45714 -960 45826 480
rect 46910 -960 47022 480
rect 48106 -960 48218 480
rect 49302 -960 49414 480
rect 50498 -960 50610 480
rect 51602 -960 51714 480
rect 52798 -960 52910 480
rect 53994 -960 54106 480
rect 55190 -960 55302 480
rect 56386 -960 56498 480
rect 57582 -960 57694 480
rect 58778 -960 58890 480
rect 59974 -960 60086 480
rect 61170 -960 61282 480
rect 62366 -960 62478 480
rect 63562 -960 63674 480
rect 64758 -960 64870 480
rect 65954 -960 66066 480
rect 67150 -960 67262 480
rect 68254 -960 68366 480
rect 69450 -960 69562 480
rect 70646 -960 70758 480
rect 71842 -960 71954 480
rect 73038 -960 73150 480
rect 74234 -960 74346 480
rect 75430 -960 75542 480
rect 76626 -960 76738 480
rect 77822 -960 77934 480
rect 79018 -960 79130 480
rect 80214 -960 80326 480
rect 81410 -960 81522 480
rect 82606 -960 82718 480
rect 83802 -960 83914 480
rect 84906 -960 85018 480
rect 86102 -960 86214 480
rect 87298 -960 87410 480
rect 88494 -960 88606 480
rect 89690 -960 89802 480
rect 90886 -960 90998 480
rect 92082 -960 92194 480
rect 93278 -960 93390 480
rect 94474 -960 94586 480
rect 95670 -960 95782 480
rect 96866 -960 96978 480
rect 98062 -960 98174 480
rect 99258 -960 99370 480
rect 100454 -960 100566 480
rect 101558 -960 101670 480
rect 102754 -960 102866 480
rect 103950 -960 104062 480
rect 105146 -960 105258 480
rect 106342 -960 106454 480
rect 107538 -960 107650 480
rect 108734 -960 108846 480
rect 109930 -960 110042 480
rect 111126 -960 111238 480
rect 112322 -960 112434 480
rect 113518 -960 113630 480
rect 114714 -960 114826 480
rect 115910 -960 116022 480
rect 117106 -960 117218 480
rect 118210 -960 118322 480
rect 119406 -960 119518 480
rect 120602 -960 120714 480
rect 121798 -960 121910 480
rect 122994 -960 123106 480
rect 124190 -960 124302 480
rect 125386 -960 125498 480
rect 126582 -960 126694 480
rect 127778 -960 127890 480
rect 128974 -960 129086 480
rect 130170 -960 130282 480
rect 131366 -960 131478 480
rect 132562 -960 132674 480
rect 133758 -960 133870 480
rect 134862 -960 134974 480
rect 136058 -960 136170 480
rect 137254 -960 137366 480
rect 138450 -960 138562 480
rect 139646 -960 139758 480
rect 140842 -960 140954 480
rect 142038 -960 142150 480
rect 143234 -960 143346 480
rect 144430 -960 144542 480
rect 145626 -960 145738 480
rect 146822 -960 146934 480
rect 148018 -960 148130 480
rect 149214 -960 149326 480
rect 150410 -960 150522 480
rect 151514 -960 151626 480
rect 152710 -960 152822 480
rect 153906 -960 154018 480
rect 155102 -960 155214 480
rect 156298 -960 156410 480
rect 157494 -960 157606 480
rect 158690 -960 158802 480
rect 159886 -960 159998 480
rect 161082 -960 161194 480
rect 162278 -960 162390 480
rect 163474 -960 163586 480
rect 164670 -960 164782 480
rect 165866 -960 165978 480
rect 167062 -960 167174 480
rect 168166 -960 168278 480
rect 169362 -960 169474 480
rect 170558 -960 170670 480
rect 171754 -960 171866 480
rect 172950 -960 173062 480
rect 174146 -960 174258 480
rect 175342 -960 175454 480
rect 176538 -960 176650 480
rect 177734 -960 177846 480
rect 178930 -960 179042 480
rect 180126 -960 180238 480
rect 181322 -960 181434 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184818 -960 184930 480
rect 186014 -960 186126 480
rect 187210 -960 187322 480
rect 188406 -960 188518 480
rect 189602 -960 189714 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197974 -960 198086 480
rect 199170 -960 199282 480
rect 200366 -960 200478 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206254 -960 206366 480
rect 207450 -960 207562 480
rect 208646 -960 208758 480
rect 209842 -960 209954 480
rect 211038 -960 211150 480
rect 212234 -960 212346 480
rect 213430 -960 213542 480
rect 214626 -960 214738 480
rect 215822 -960 215934 480
rect 217018 -960 217130 480
rect 218122 -960 218234 480
rect 219318 -960 219430 480
rect 220514 -960 220626 480
rect 221710 -960 221822 480
rect 222906 -960 223018 480
rect 224102 -960 224214 480
rect 225298 -960 225410 480
rect 226494 -960 226606 480
rect 227690 -960 227802 480
rect 228886 -960 228998 480
rect 230082 -960 230194 480
rect 231278 -960 231390 480
rect 232474 -960 232586 480
rect 233670 -960 233782 480
rect 234774 -960 234886 480
rect 235970 -960 236082 480
rect 237166 -960 237278 480
rect 238362 -960 238474 480
rect 239558 -960 239670 480
rect 240754 -960 240866 480
rect 241950 -960 242062 480
rect 243146 -960 243258 480
rect 244342 -960 244454 480
rect 245538 -960 245650 480
rect 246734 -960 246846 480
rect 247930 -960 248042 480
rect 249126 -960 249238 480
rect 250322 -960 250434 480
rect 251426 -960 251538 480
rect 252622 -960 252734 480
rect 253818 -960 253930 480
rect 255014 -960 255126 480
rect 256210 -960 256322 480
rect 257406 -960 257518 480
rect 258602 -960 258714 480
rect 259798 -960 259910 480
rect 260994 -960 261106 480
rect 262190 -960 262302 480
rect 263386 -960 263498 480
rect 264582 -960 264694 480
rect 265778 -960 265890 480
rect 266974 -960 267086 480
rect 268078 -960 268190 480
rect 269274 -960 269386 480
rect 270470 -960 270582 480
rect 271666 -960 271778 480
rect 272862 -960 272974 480
rect 274058 -960 274170 480
rect 275254 -960 275366 480
rect 276450 -960 276562 480
rect 277646 -960 277758 480
rect 278842 -960 278954 480
rect 280038 -960 280150 480
rect 281234 -960 281346 480
rect 282430 -960 282542 480
rect 283626 -960 283738 480
rect 284730 -960 284842 480
rect 285926 -960 286038 480
rect 287122 -960 287234 480
rect 288318 -960 288430 480
rect 289514 -960 289626 480
rect 290710 -960 290822 480
rect 291906 -960 292018 480
rect 293102 -960 293214 480
rect 294298 -960 294410 480
rect 295494 -960 295606 480
rect 296690 -960 296802 480
rect 297886 -960 297998 480
rect 299082 -960 299194 480
rect 300278 -960 300390 480
rect 301382 -960 301494 480
rect 302578 -960 302690 480
rect 303774 -960 303886 480
rect 304970 -960 305082 480
rect 306166 -960 306278 480
rect 307362 -960 307474 480
rect 308558 -960 308670 480
rect 309754 -960 309866 480
rect 310950 -960 311062 480
rect 312146 -960 312258 480
rect 313342 -960 313454 480
rect 314538 -960 314650 480
rect 315734 -960 315846 480
rect 316930 -960 317042 480
rect 318034 -960 318146 480
rect 319230 -960 319342 480
rect 320426 -960 320538 480
rect 321622 -960 321734 480
rect 322818 -960 322930 480
rect 324014 -960 324126 480
rect 325210 -960 325322 480
rect 326406 -960 326518 480
rect 327602 -960 327714 480
rect 328798 -960 328910 480
rect 329994 -960 330106 480
rect 331190 -960 331302 480
rect 332386 -960 332498 480
rect 333582 -960 333694 480
rect 334686 -960 334798 480
rect 335882 -960 335994 480
rect 337078 -960 337190 480
rect 338274 -960 338386 480
rect 339470 -960 339582 480
rect 340666 -960 340778 480
rect 341862 -960 341974 480
rect 343058 -960 343170 480
rect 344254 -960 344366 480
rect 345450 -960 345562 480
rect 346646 -960 346758 480
rect 347842 -960 347954 480
rect 349038 -960 349150 480
rect 350234 -960 350346 480
rect 351338 -960 351450 480
rect 352534 -960 352646 480
rect 353730 -960 353842 480
rect 354926 -960 355038 480
rect 356122 -960 356234 480
rect 357318 -960 357430 480
rect 358514 -960 358626 480
rect 359710 -960 359822 480
rect 360906 -960 361018 480
rect 362102 -960 362214 480
rect 363298 -960 363410 480
rect 364494 -960 364606 480
rect 365690 -960 365802 480
rect 366886 -960 366998 480
rect 367990 -960 368102 480
rect 369186 -960 369298 480
rect 370382 -960 370494 480
rect 371578 -960 371690 480
rect 372774 -960 372886 480
rect 373970 -960 374082 480
rect 375166 -960 375278 480
rect 376362 -960 376474 480
rect 377558 -960 377670 480
rect 378754 -960 378866 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384642 -960 384754 480
rect 385838 -960 385950 480
rect 387034 -960 387146 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395406 -960 395518 480
rect 396602 -960 396714 480
rect 397798 -960 397910 480
rect 398994 -960 399106 480
rect 400190 -960 400302 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403686 -960 403798 480
rect 404882 -960 404994 480
rect 406078 -960 406190 480
rect 407274 -960 407386 480
rect 408470 -960 408582 480
rect 409666 -960 409778 480
rect 410862 -960 410974 480
rect 412058 -960 412170 480
rect 413254 -960 413366 480
rect 414450 -960 414562 480
rect 415646 -960 415758 480
rect 416842 -960 416954 480
rect 417946 -960 418058 480
rect 419142 -960 419254 480
rect 420338 -960 420450 480
rect 421534 -960 421646 480
rect 422730 -960 422842 480
rect 423926 -960 424038 480
rect 425122 -960 425234 480
rect 426318 -960 426430 480
rect 427514 -960 427626 480
rect 428710 -960 428822 480
rect 429906 -960 430018 480
rect 431102 -960 431214 480
rect 432298 -960 432410 480
rect 433494 -960 433606 480
rect 434598 -960 434710 480
rect 435794 -960 435906 480
rect 436990 -960 437102 480
rect 438186 -960 438298 480
rect 439382 -960 439494 480
rect 440578 -960 440690 480
rect 441774 -960 441886 480
rect 442970 -960 443082 480
rect 444166 -960 444278 480
rect 445362 -960 445474 480
rect 446558 -960 446670 480
rect 447754 -960 447866 480
rect 448950 -960 449062 480
rect 450146 -960 450258 480
rect 451250 -960 451362 480
rect 452446 -960 452558 480
rect 453642 -960 453754 480
rect 454838 -960 454950 480
rect 456034 -960 456146 480
rect 457230 -960 457342 480
rect 458426 -960 458538 480
rect 459622 -960 459734 480
rect 460818 -960 460930 480
rect 462014 -960 462126 480
rect 463210 -960 463322 480
rect 464406 -960 464518 480
rect 465602 -960 465714 480
rect 466798 -960 466910 480
rect 467902 -960 468014 480
rect 469098 -960 469210 480
rect 470294 -960 470406 480
rect 471490 -960 471602 480
rect 472686 -960 472798 480
rect 473882 -960 473994 480
rect 475078 -960 475190 480
rect 476274 -960 476386 480
rect 477470 -960 477582 480
rect 478666 -960 478778 480
rect 479862 -960 479974 480
rect 481058 -960 481170 480
rect 482254 -960 482366 480
rect 483450 -960 483562 480
rect 484554 -960 484666 480
rect 485750 -960 485862 480
rect 486946 -960 487058 480
rect 488142 -960 488254 480
rect 489338 -960 489450 480
rect 490534 -960 490646 480
rect 491730 -960 491842 480
rect 492926 -960 493038 480
rect 494122 -960 494234 480
rect 495318 -960 495430 480
rect 496514 -960 496626 480
rect 497710 -960 497822 480
rect 498906 -960 499018 480
rect 500102 -960 500214 480
rect 501206 -960 501318 480
rect 502402 -960 502514 480
rect 503598 -960 503710 480
rect 504794 -960 504906 480
rect 505990 -960 506102 480
rect 507186 -960 507298 480
rect 508382 -960 508494 480
rect 509578 -960 509690 480
rect 510774 -960 510886 480
rect 511970 -960 512082 480
rect 513166 -960 513278 480
rect 514362 -960 514474 480
rect 515558 -960 515670 480
rect 516754 -960 516866 480
rect 517858 -960 517970 480
rect 519054 -960 519166 480
rect 520250 -960 520362 480
rect 521446 -960 521558 480
rect 522642 -960 522754 480
rect 523838 -960 523950 480
rect 525034 -960 525146 480
rect 526230 -960 526342 480
rect 527426 -960 527538 480
rect 528622 -960 528734 480
rect 529818 -960 529930 480
rect 531014 -960 531126 480
rect 532210 -960 532322 480
rect 533406 -960 533518 480
rect 534510 -960 534622 480
rect 535706 -960 535818 480
rect 536902 -960 537014 480
rect 538098 -960 538210 480
rect 539294 -960 539406 480
rect 540490 -960 540602 480
rect 541686 -960 541798 480
rect 542882 -960 542994 480
rect 544078 -960 544190 480
rect 545274 -960 545386 480
rect 546470 -960 546582 480
rect 547666 -960 547778 480
rect 548862 -960 548974 480
rect 550058 -960 550170 480
rect 551162 -960 551274 480
rect 552358 -960 552470 480
rect 553554 -960 553666 480
rect 554750 -960 554862 480
rect 555946 -960 556058 480
rect 557142 -960 557254 480
rect 558338 -960 558450 480
rect 559534 -960 559646 480
rect 560730 -960 560842 480
rect 561926 -960 562038 480
rect 563122 -960 563234 480
rect 564318 -960 564430 480
rect 565514 -960 565626 480
rect 566710 -960 566822 480
rect 567814 -960 567926 480
rect 569010 -960 569122 480
rect 570206 -960 570318 480
rect 571402 -960 571514 480
rect 572598 -960 572710 480
rect 573794 -960 573906 480
rect 574990 -960 575102 480
rect 576186 -960 576298 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3606 667936 3662 667992
rect 2962 653540 3018 653576
rect 2962 653520 2964 653540
rect 2964 653520 3016 653540
rect 3016 653520 3018 653540
rect 2962 595992 3018 596048
rect 2962 538600 3018 538656
rect 2962 481072 3018 481128
rect 2962 423680 3018 423736
rect 3698 610408 3754 610464
rect 3698 609456 3754 609512
rect 3698 553016 3754 553072
rect 24766 545536 24822 545592
rect 24858 509904 24914 509960
rect 3790 495488 3846 495544
rect 3974 437960 4030 438016
rect 3882 423680 3938 423736
rect 24858 402056 24914 402112
rect 24766 234640 24822 234696
rect 300122 700576 300178 700632
rect 27250 581168 27306 581224
rect 269302 547612 269304 547632
rect 269304 547612 269356 547632
rect 269356 547612 269358 547632
rect 269302 547576 269358 547612
rect 269302 511944 269358 512000
rect 270038 440680 270094 440736
rect 269302 405320 269358 405376
rect 270406 345752 270462 345808
rect 268658 341808 268714 341864
rect 27250 270816 27306 270872
rect 268014 201728 268070 201784
rect 24950 199008 25006 199064
rect 270222 339632 270278 339688
rect 269394 332288 269450 332344
rect 269394 328344 269450 328400
rect 269394 325252 269396 325272
rect 269396 325252 269448 325272
rect 269448 325252 269450 325272
rect 269394 325216 269450 325252
rect 270498 322224 270554 322280
rect 270774 352688 270830 352744
rect 270682 335416 270738 335472
rect 270590 318280 270646 318336
rect 269026 237360 269082 237416
rect 268658 166096 268714 166152
rect 269302 130464 269358 130520
rect 24858 128016 24914 128072
rect 269302 95104 269358 95160
rect 24950 92384 25006 92440
rect 276386 382064 276442 382120
rect 282642 359352 282698 359408
rect 285586 359216 285642 359272
rect 286230 359216 286286 359272
rect 294418 586200 294474 586256
rect 292762 586064 292818 586120
rect 291290 546760 291346 546816
rect 293682 384240 293738 384296
rect 294418 382200 294474 382256
rect 274086 354864 274142 354920
rect 274454 354864 274510 354920
rect 275926 354864 275982 354920
rect 290462 354864 290518 354920
rect 291382 354864 291438 354920
rect 297638 354864 297694 354920
rect 300122 381928 300178 381984
rect 300122 381248 300178 381304
rect 364982 699896 365038 699952
rect 579894 697992 579950 698048
rect 578514 674600 578570 674656
rect 307482 585928 307538 585984
rect 309322 511556 309378 511592
rect 309322 511536 309324 511556
rect 309324 511536 309376 511556
rect 309376 511536 309378 511556
rect 309322 504872 309378 504928
rect 309966 473728 310022 473784
rect 309966 463664 310022 463720
rect 309966 432520 310022 432576
rect 309966 422456 310022 422512
rect 309782 412120 309838 412176
rect 309782 402056 309838 402112
rect 309782 391448 309838 391504
rect 309782 381248 309838 381304
rect 309414 370912 309470 370968
rect 309414 360848 309470 360904
rect 306470 355272 306526 355328
rect 311622 566616 311678 566672
rect 299478 354864 299534 354920
rect 313554 347928 313610 347984
rect 311530 317056 311586 317112
rect 274086 316240 274142 316296
rect 290646 315696 290702 315752
rect 275834 276664 275890 276720
rect 275190 71984 275246 72040
rect 276110 315560 276166 315616
rect 280802 313112 280858 313168
rect 287978 313384 288034 313440
rect 288438 313384 288494 313440
rect 285586 312024 285642 312080
rect 286230 312024 286286 312080
rect 276018 272176 276074 272232
rect 276202 272040 276258 272096
rect 292854 316240 292910 316296
rect 295246 316240 295302 316296
rect 295890 275324 295946 275360
rect 295890 275304 295892 275324
rect 295892 275304 295944 275324
rect 295944 275304 295946 275324
rect 300030 316240 300086 316296
rect 309414 316240 309470 316296
rect 306654 315560 306710 315616
rect 306562 288496 306618 288552
rect 306746 288496 306802 288552
rect 306746 276664 306802 276720
rect 299570 92656 299626 92712
rect 313738 330656 313794 330712
rect 313646 323584 313702 323640
rect 313646 320592 313702 320648
rect 313922 351736 313978 351792
rect 313830 326984 313886 327040
rect 314014 344412 314070 344448
rect 314014 344392 314016 344412
rect 314016 344392 314068 344412
rect 314068 344392 314070 344412
rect 314014 341128 314070 341184
rect 579894 651072 579950 651128
rect 578790 627680 578846 627736
rect 579894 604152 579950 604208
rect 461674 586200 461730 586256
rect 485778 586064 485834 586120
rect 533986 585928 534042 585984
rect 315026 580488 315082 580544
rect 318614 546760 318670 546816
rect 315026 545128 315082 545184
rect 315026 509380 315082 509416
rect 315026 509360 315028 509380
rect 315028 509360 315080 509380
rect 315080 509360 315082 509380
rect 315026 402328 315082 402384
rect 379518 382200 379574 382256
rect 427726 382064 427782 382120
rect 548062 381928 548118 381984
rect 314290 351736 314346 351792
rect 314198 338000 314254 338056
rect 578790 580760 578846 580816
rect 579894 557232 579950 557288
rect 560850 547712 560906 547768
rect 579158 533840 579214 533896
rect 560022 512080 560078 512136
rect 578790 486784 578846 486840
rect 560850 440680 560906 440736
rect 314014 320592 314070 320648
rect 578790 439864 578846 439920
rect 560850 405320 560906 405376
rect 579894 510312 579950 510368
rect 579894 463392 579950 463448
rect 579894 416472 579950 416528
rect 579250 415112 579306 415168
rect 579894 415112 579950 415168
rect 579342 392944 579398 393000
rect 315026 270272 315082 270328
rect 315026 234640 315082 234696
rect 560850 237360 560906 237416
rect 560850 201728 560906 201784
rect 315026 199008 315082 199064
rect 558918 130464 558974 130520
rect 560850 95104 560906 95160
rect 315026 92384 315082 92440
rect 583390 3576 583446 3632
<< metal3 >>
rect 299054 700572 299060 700636
rect 299124 700634 299130 700636
rect 300117 700634 300183 700637
rect 299124 700632 300183 700634
rect 299124 700576 300122 700632
rect 300178 700576 300183 700632
rect 299124 700574 300183 700576
rect 299124 700572 299130 700574
rect 300117 700571 300183 700574
rect 275134 699892 275140 699956
rect 275204 699954 275210 699956
rect 364977 699954 365043 699957
rect 275204 699952 365043 699954
rect 275204 699896 364982 699952
rect 365038 699896 365043 699952
rect 275204 699894 365043 699896
rect 275204 699892 275210 699894
rect 364977 699891 365043 699894
rect 579889 698050 579955 698053
rect 583520 698050 584960 698140
rect 579889 698048 584960 698050
rect 579889 697992 579894 698048
rect 579950 697992 584960 698048
rect 579889 697990 584960 697992
rect 579889 697987 579955 697990
rect 583520 697900 584960 697990
rect -960 696540 480 696780
rect 583520 686204 584960 686444
rect -960 682124 480 682364
rect 578509 674658 578575 674661
rect 583520 674658 584960 674748
rect 578509 674656 584960 674658
rect 578509 674600 578514 674656
rect 578570 674600 584960 674656
rect 578509 674598 584960 674600
rect 578509 674595 578575 674598
rect 583520 674508 584960 674598
rect -960 667994 480 668084
rect 3601 667994 3667 667997
rect -960 667992 3667 667994
rect -960 667936 3606 667992
rect 3662 667936 3667 667992
rect -960 667934 3667 667936
rect -960 667844 480 667934
rect 3601 667931 3667 667934
rect 583520 662676 584960 662916
rect -960 653578 480 653668
rect 2957 653578 3023 653581
rect -960 653576 3023 653578
rect -960 653520 2962 653576
rect 3018 653520 3023 653576
rect -960 653518 3023 653520
rect -960 653428 480 653518
rect 2957 653515 3023 653518
rect 579889 651130 579955 651133
rect 583520 651130 584960 651220
rect 579889 651128 584960 651130
rect 579889 651072 579894 651128
rect 579950 651072 584960 651128
rect 579889 651070 584960 651072
rect 579889 651067 579955 651070
rect 583520 650980 584960 651070
rect 583520 639284 584960 639524
rect -960 639012 480 639252
rect 578785 627738 578851 627741
rect 583520 627738 584960 627828
rect 578785 627736 584960 627738
rect 578785 627680 578790 627736
rect 578846 627680 584960 627736
rect 578785 627678 584960 627680
rect 578785 627675 578851 627678
rect 583520 627588 584960 627678
rect -960 624732 480 624972
rect 583520 615756 584960 615996
rect -960 610466 480 610556
rect 3693 610466 3759 610469
rect -960 610464 3759 610466
rect -960 610408 3698 610464
rect 3754 610408 3759 610464
rect -960 610406 3759 610408
rect -960 610316 480 610406
rect 3693 610403 3759 610406
rect 3693 609514 3759 609517
rect 310646 609514 310652 609516
rect 3693 609512 310652 609514
rect 3693 609456 3698 609512
rect 3754 609456 310652 609512
rect 3693 609454 310652 609456
rect 3693 609451 3759 609454
rect 310646 609452 310652 609454
rect 310716 609452 310722 609516
rect 579889 604210 579955 604213
rect 583520 604210 584960 604300
rect 579889 604208 584960 604210
rect 579889 604152 579894 604208
rect 579950 604152 584960 604208
rect 579889 604150 584960 604152
rect 579889 604147 579955 604150
rect 583520 604060 584960 604150
rect -960 596050 480 596140
rect 2957 596050 3023 596053
rect -960 596048 3023 596050
rect -960 595992 2962 596048
rect 3018 595992 3023 596048
rect -960 595990 3023 595992
rect -960 595900 480 595990
rect 2957 595987 3023 595990
rect 583520 592364 584960 592604
rect 294413 586258 294479 586261
rect 295742 586258 295748 586260
rect 294413 586256 295748 586258
rect 294413 586200 294418 586256
rect 294474 586200 295748 586256
rect 294413 586198 295748 586200
rect 294413 586195 294479 586198
rect 295742 586196 295748 586198
rect 295812 586258 295818 586260
rect 461669 586258 461735 586261
rect 295812 586256 461735 586258
rect 295812 586200 461674 586256
rect 461730 586200 461735 586256
rect 295812 586198 461735 586200
rect 295812 586196 295818 586198
rect 461669 586195 461735 586198
rect 292757 586124 292823 586125
rect 292757 586120 292804 586124
rect 292868 586122 292874 586124
rect 485773 586122 485839 586125
rect 292868 586120 485839 586122
rect 292757 586064 292762 586120
rect 292868 586064 485778 586120
rect 485834 586064 485839 586120
rect 292757 586060 292804 586064
rect 292868 586062 485839 586064
rect 292868 586060 292874 586062
rect 292757 586059 292823 586060
rect 485773 586059 485839 586062
rect 306598 585924 306604 585988
rect 306668 585986 306674 585988
rect 307477 585986 307543 585989
rect 533981 585986 534047 585989
rect 306668 585984 534047 585986
rect 306668 585928 307482 585984
rect 307538 585928 533986 585984
rect 534042 585928 534047 585984
rect 306668 585926 534047 585928
rect 306668 585924 306674 585926
rect 307477 585923 307543 585926
rect 533981 585923 534047 585926
rect -960 581620 480 581860
rect 27245 581226 27311 581229
rect 27245 581224 27354 581226
rect 27245 581168 27250 581224
rect 27306 581168 27354 581224
rect 27245 581163 27354 581168
rect 27294 580584 27354 581163
rect 578785 580818 578851 580821
rect 583520 580818 584960 580908
rect 578785 580816 584960 580818
rect 578785 580760 578790 580816
rect 578846 580760 584960 580816
rect 578785 580758 584960 580760
rect 578785 580755 578851 580758
rect 583520 580668 584960 580758
rect 315021 580546 315087 580549
rect 318934 580546 318994 580584
rect 315021 580544 318994 580546
rect 315021 580488 315026 580544
rect 315082 580488 318994 580544
rect 315021 580486 318994 580488
rect 315021 580483 315087 580486
rect 583520 568836 584960 569076
rect -960 567204 480 567444
rect 310462 566612 310468 566676
rect 310532 566674 310538 566676
rect 311617 566674 311683 566677
rect 310532 566672 311683 566674
rect 310532 566616 311622 566672
rect 311678 566616 311683 566672
rect 310532 566614 311683 566616
rect 310532 566612 310538 566614
rect 311617 566611 311683 566614
rect 579889 557290 579955 557293
rect 583520 557290 584960 557380
rect 579889 557288 584960 557290
rect 579889 557232 579894 557288
rect 579950 557232 584960 557288
rect 579889 557230 584960 557232
rect 579889 557227 579955 557230
rect 583520 557140 584960 557230
rect -960 553074 480 553164
rect 3693 553074 3759 553077
rect -960 553072 3759 553074
rect -960 553016 3698 553072
rect 3754 553016 3759 553072
rect -960 553014 3759 553016
rect -960 552924 480 553014
rect 3693 553011 3759 553014
rect 560845 547770 560911 547773
rect 558870 547768 560911 547770
rect 558870 547712 560850 547768
rect 560906 547712 560911 547768
rect 558870 547710 560911 547712
rect 558870 547702 558930 547710
rect 560845 547707 560911 547710
rect 266524 547642 266922 547702
rect 558716 547642 558930 547702
rect 266862 547634 266922 547642
rect 269297 547634 269363 547637
rect 266862 547632 269363 547634
rect 266862 547576 269302 547632
rect 269358 547576 269363 547632
rect 266862 547574 269363 547576
rect 269297 547571 269363 547574
rect 291285 546818 291351 546821
rect 293534 546818 293540 546820
rect 291285 546816 293540 546818
rect 291285 546760 291290 546816
rect 291346 546760 293540 546816
rect 291285 546758 293540 546760
rect 291285 546755 291351 546758
rect 293534 546756 293540 546758
rect 293604 546818 293610 546820
rect 318609 546818 318675 546821
rect 293604 546816 318675 546818
rect 293604 546760 318614 546816
rect 318670 546760 318675 546816
rect 293604 546758 318675 546760
rect 293604 546756 293610 546758
rect 318609 546755 318675 546758
rect 24761 545594 24827 545597
rect 24761 545592 26802 545594
rect 24761 545536 24766 545592
rect 24822 545536 26802 545592
rect 24761 545534 26802 545536
rect 24761 545531 24827 545534
rect 26742 544952 26802 545534
rect 583520 545444 584960 545684
rect 315021 545186 315087 545189
rect 315021 545184 318994 545186
rect 315021 545128 315026 545184
rect 315082 545128 318994 545184
rect 315021 545126 318994 545128
rect 315021 545123 315087 545126
rect 318934 544952 318994 545126
rect -960 538658 480 538748
rect 2957 538658 3023 538661
rect -960 538656 3023 538658
rect -960 538600 2962 538656
rect 3018 538600 3023 538656
rect -960 538598 3023 538600
rect -960 538508 480 538598
rect 2957 538595 3023 538598
rect 579153 533898 579219 533901
rect 583520 533898 584960 533988
rect 579153 533896 584960 533898
rect 579153 533840 579158 533896
rect 579214 533840 584960 533896
rect 579153 533838 584960 533840
rect 579153 533835 579219 533838
rect 583520 533748 584960 533838
rect -960 524092 480 524332
rect 583520 521916 584960 522156
rect 560017 512138 560083 512141
rect 558870 512136 560083 512138
rect 558870 512080 560022 512136
rect 560078 512080 560083 512136
rect 558870 512078 560083 512080
rect 558870 512070 558930 512078
rect 560017 512075 560083 512078
rect 266524 512010 266922 512070
rect 558716 512010 558930 512070
rect 266862 512002 266922 512010
rect 269297 512002 269363 512005
rect 266862 512000 269363 512002
rect 266862 511944 269302 512000
rect 269358 511944 269363 512000
rect 266862 511942 269363 511944
rect 269297 511939 269363 511942
rect 309317 511594 309383 511597
rect 310462 511594 310468 511596
rect 309317 511592 310468 511594
rect 309317 511536 309322 511592
rect 309378 511536 310468 511592
rect 309317 511534 310468 511536
rect 309317 511531 309383 511534
rect 310462 511532 310468 511534
rect 310532 511532 310538 511596
rect 579889 510370 579955 510373
rect 583520 510370 584960 510460
rect 579889 510368 584960 510370
rect 579889 510312 579894 510368
rect 579950 510312 584960 510368
rect 579889 510310 584960 510312
rect 579889 510307 579955 510310
rect 583520 510220 584960 510310
rect -960 509812 480 510052
rect 24853 509962 24919 509965
rect 24853 509960 26802 509962
rect 24853 509904 24858 509960
rect 24914 509904 26802 509960
rect 24853 509902 26802 509904
rect 24853 509899 24919 509902
rect 26742 509320 26802 509902
rect 315021 509418 315087 509421
rect 315021 509416 318994 509418
rect 315021 509360 315026 509416
rect 315082 509360 318994 509416
rect 315021 509358 318994 509360
rect 315021 509355 315087 509358
rect 318934 509320 318994 509358
rect 309317 504932 309383 504933
rect 309317 504930 309364 504932
rect 309272 504928 309364 504930
rect 309272 504872 309322 504928
rect 309272 504870 309364 504872
rect 309317 504868 309364 504870
rect 309428 504868 309434 504932
rect 309317 504867 309383 504868
rect 583520 498524 584960 498764
rect 309358 497660 309364 497724
rect 309428 497660 309434 497724
rect 309366 497450 309426 497660
rect 309542 497450 309548 497452
rect 309366 497390 309548 497450
rect 309542 497388 309548 497390
rect 309612 497388 309618 497452
rect -960 495546 480 495636
rect 3785 495546 3851 495549
rect -960 495544 3851 495546
rect -960 495488 3790 495544
rect 3846 495488 3851 495544
rect -960 495486 3851 495488
rect -960 495396 480 495486
rect 3785 495483 3851 495486
rect 578785 486842 578851 486845
rect 583520 486842 584960 486932
rect 578785 486840 584960 486842
rect 578785 486784 578790 486840
rect 578846 486784 584960 486840
rect 578785 486782 584960 486784
rect 578785 486779 578851 486782
rect 583520 486692 584960 486782
rect 309726 484196 309732 484260
rect 309796 484196 309802 484260
rect 309734 484122 309794 484196
rect 309910 484122 309916 484124
rect 309734 484062 309916 484122
rect 309910 484060 309916 484062
rect 309980 484060 309986 484124
rect -960 481130 480 481220
rect 2957 481130 3023 481133
rect -960 481128 3023 481130
rect -960 481072 2962 481128
rect 3018 481072 3023 481128
rect -960 481070 3023 481072
rect -960 480980 480 481070
rect 2957 481067 3023 481070
rect 583520 474996 584960 475236
rect 309910 473860 309916 473924
rect 309980 473860 309986 473924
rect 309918 473789 309978 473860
rect 309918 473784 310027 473789
rect 309918 473728 309966 473784
rect 310022 473728 310027 473784
rect 309918 473726 310027 473728
rect 309961 473723 310027 473726
rect -960 466700 480 466940
rect 309961 463722 310027 463725
rect 310094 463722 310100 463724
rect 309961 463720 310100 463722
rect 309961 463664 309966 463720
rect 310022 463664 310100 463720
rect 309961 463662 310100 463664
rect 309961 463659 310027 463662
rect 310094 463660 310100 463662
rect 310164 463660 310170 463724
rect 579889 463450 579955 463453
rect 583520 463450 584960 463540
rect 579889 463448 584960 463450
rect 579889 463392 579894 463448
rect 579950 463392 584960 463448
rect 579889 463390 584960 463392
rect 579889 463387 579955 463390
rect 583520 463300 584960 463390
rect 309542 458492 309548 458556
rect 309612 458554 309618 458556
rect 310094 458554 310100 458556
rect 309612 458494 310100 458554
rect 309612 458492 309618 458494
rect 310094 458492 310100 458494
rect 310164 458492 310170 458556
rect -960 452284 480 452524
rect 583520 451604 584960 451844
rect 309542 445980 309548 446044
rect 309612 446042 309618 446044
rect 310094 446042 310100 446044
rect 309612 445982 310100 446042
rect 309612 445980 309618 445982
rect 310094 445980 310100 445982
rect 310164 445980 310170 446044
rect 266524 440746 267106 440806
rect 558716 440746 559298 440806
rect 267046 440738 267106 440746
rect 270033 440738 270099 440741
rect 267046 440736 270099 440738
rect 267046 440680 270038 440736
rect 270094 440680 270099 440736
rect 267046 440678 270099 440680
rect 559238 440738 559298 440746
rect 560845 440738 560911 440741
rect 559238 440736 560911 440738
rect 559238 440680 560850 440736
rect 560906 440680 560911 440736
rect 559238 440678 560911 440680
rect 270033 440675 270099 440678
rect 560845 440675 560911 440678
rect 578785 439922 578851 439925
rect 583520 439922 584960 440012
rect 578785 439920 584960 439922
rect 578785 439864 578790 439920
rect 578846 439864 584960 439920
rect 578785 439862 584960 439864
rect 578785 439859 578851 439862
rect 583520 439772 584960 439862
rect -960 438018 480 438108
rect 3969 438018 4035 438021
rect -960 438016 4035 438018
rect -960 437960 3974 438016
rect 4030 437960 4035 438016
rect -960 437958 4035 437960
rect -960 437868 480 437958
rect 3969 437955 4035 437958
rect 310094 435780 310100 435844
rect 310164 435780 310170 435844
rect 310102 435708 310162 435780
rect 310094 435644 310100 435708
rect 310164 435644 310170 435708
rect 309961 432580 310027 432581
rect 309910 432516 309916 432580
rect 309980 432578 310027 432580
rect 309980 432576 310072 432578
rect 310022 432520 310072 432576
rect 309980 432518 310072 432520
rect 309980 432516 310027 432518
rect 309961 432515 310027 432516
rect 583520 428076 584960 428316
rect -960 423738 480 423828
rect 2957 423738 3023 423741
rect 3877 423738 3943 423741
rect -960 423736 3943 423738
rect -960 423680 2962 423736
rect 3018 423680 3882 423736
rect 3938 423680 3943 423736
rect -960 423678 3943 423680
rect -960 423588 480 423678
rect 2957 423675 3023 423678
rect 3877 423675 3943 423678
rect 309726 422452 309732 422516
rect 309796 422514 309802 422516
rect 309961 422514 310027 422517
rect 309796 422512 310027 422514
rect 309796 422456 309966 422512
rect 310022 422456 310027 422512
rect 309796 422454 310027 422456
rect 309796 422452 309802 422454
rect 309961 422451 310027 422454
rect 579889 416530 579955 416533
rect 583520 416530 584960 416620
rect 579889 416528 584960 416530
rect 579889 416472 579894 416528
rect 579950 416472 584960 416528
rect 579889 416470 584960 416472
rect 579889 416467 579955 416470
rect 583520 416380 584960 416470
rect 309726 415244 309732 415308
rect 309796 415244 309802 415308
rect 309734 415034 309794 415244
rect 579245 415170 579311 415173
rect 579889 415170 579955 415173
rect 579245 415168 579955 415170
rect 579245 415112 579250 415168
rect 579306 415112 579894 415168
rect 579950 415112 579955 415168
rect 579245 415110 579955 415112
rect 579245 415107 579311 415110
rect 579889 415107 579955 415110
rect 309910 415034 309916 415036
rect 309734 414974 309916 415034
rect 309910 414972 309916 414974
rect 309980 414972 309986 415036
rect 309777 412178 309843 412181
rect 309910 412178 309916 412180
rect 309777 412176 309916 412178
rect 309777 412120 309782 412176
rect 309838 412120 309916 412176
rect 309777 412118 309916 412120
rect 309777 412115 309843 412118
rect 309910 412116 309916 412118
rect 309980 412116 309986 412180
rect -960 409172 480 409412
rect 266524 405386 266922 405446
rect 558716 405386 559298 405446
rect 266862 405378 266922 405386
rect 269297 405378 269363 405381
rect 266862 405376 269363 405378
rect 266862 405320 269302 405376
rect 269358 405320 269363 405376
rect 266862 405318 269363 405320
rect 559238 405378 559298 405386
rect 560845 405378 560911 405381
rect 559238 405376 560911 405378
rect 559238 405320 560850 405376
rect 560906 405320 560911 405376
rect 559238 405318 560911 405320
rect 269297 405315 269363 405318
rect 560845 405315 560911 405318
rect 583520 404684 584960 404924
rect 24853 402114 24919 402117
rect 26742 402114 26802 402696
rect 315021 402386 315087 402389
rect 318934 402386 318994 402696
rect 315021 402384 318994 402386
rect 315021 402328 315026 402384
rect 315082 402328 318994 402384
rect 315021 402326 318994 402328
rect 315021 402323 315087 402326
rect 309777 402114 309843 402117
rect 24853 402112 26802 402114
rect 24853 402056 24858 402112
rect 24914 402056 26802 402112
rect 24853 402054 26802 402056
rect 309734 402112 309843 402114
rect 309734 402056 309782 402112
rect 309838 402056 309843 402112
rect 24853 402051 24919 402054
rect 309734 402051 309843 402056
rect 309734 401980 309794 402051
rect 309726 401916 309732 401980
rect 309796 401916 309802 401980
rect -960 394892 480 395132
rect 309726 394572 309732 394636
rect 309796 394572 309802 394636
rect 309734 394362 309794 394572
rect 309910 394362 309916 394364
rect 309734 394302 309916 394362
rect 309910 394300 309916 394302
rect 309980 394300 309986 394364
rect 579337 393002 579403 393005
rect 583520 393002 584960 393092
rect 579337 393000 584960 393002
rect 579337 392944 579342 393000
rect 579398 392944 584960 393000
rect 579337 392942 584960 392944
rect 579337 392939 579403 392942
rect 583520 392852 584960 392942
rect 309777 391506 309843 391509
rect 309910 391506 309916 391508
rect 309777 391504 309916 391506
rect 309777 391448 309782 391504
rect 309838 391448 309916 391504
rect 309777 391446 309916 391448
rect 309777 391443 309843 391446
rect 309910 391444 309916 391446
rect 309980 391444 309986 391508
rect 293677 384300 293743 384301
rect 293677 384296 293724 384300
rect 293788 384298 293794 384300
rect 293677 384240 293682 384296
rect 293677 384236 293724 384240
rect 293788 384238 293834 384298
rect 293788 384236 293794 384238
rect 293677 384235 293743 384236
rect 294413 382258 294479 382261
rect 295006 382258 295012 382260
rect 294413 382256 295012 382258
rect 294413 382200 294418 382256
rect 294474 382200 295012 382256
rect 294413 382198 295012 382200
rect 294413 382195 294479 382198
rect 295006 382196 295012 382198
rect 295076 382258 295082 382260
rect 379513 382258 379579 382261
rect 295076 382256 379579 382258
rect 295076 382200 379518 382256
rect 379574 382200 379579 382256
rect 295076 382198 379579 382200
rect 295076 382196 295082 382198
rect 379513 382195 379579 382198
rect 276238 382060 276244 382124
rect 276308 382122 276314 382124
rect 276381 382122 276447 382125
rect 427721 382122 427787 382125
rect 276308 382120 427787 382122
rect 276308 382064 276386 382120
rect 276442 382064 427726 382120
rect 427782 382064 427787 382120
rect 276308 382062 427787 382064
rect 276308 382060 276314 382062
rect 276381 382059 276447 382062
rect 427721 382059 427787 382062
rect 300117 381986 300183 381989
rect 548057 381986 548123 381989
rect 300117 381984 548123 381986
rect 300117 381928 300122 381984
rect 300178 381928 548062 381984
rect 548118 381928 548123 381984
rect 300117 381926 548123 381928
rect 300117 381923 300183 381926
rect 548057 381923 548123 381926
rect 300117 381308 300183 381309
rect 309777 381308 309843 381309
rect 300117 381304 300164 381308
rect 300228 381306 300234 381308
rect 309726 381306 309732 381308
rect 300117 381248 300122 381304
rect 300117 381244 300164 381248
rect 300228 381246 300274 381306
rect 309686 381246 309732 381306
rect 309796 381304 309843 381308
rect 309838 381248 309843 381304
rect 300228 381244 300234 381246
rect 309726 381244 309732 381246
rect 309796 381244 309843 381248
rect 300117 381243 300183 381244
rect 309777 381243 309843 381244
rect 583520 381156 584960 381396
rect -960 380476 480 380716
rect 309726 374098 309732 374100
rect 309550 374038 309732 374098
rect 309550 373828 309610 374038
rect 309726 374036 309732 374038
rect 309796 374036 309802 374100
rect 309542 373764 309548 373828
rect 309612 373764 309618 373828
rect 309409 370970 309475 370973
rect 309542 370970 309548 370972
rect 309409 370968 309548 370970
rect 309409 370912 309414 370968
rect 309470 370912 309548 370968
rect 309409 370910 309548 370912
rect 309409 370907 309475 370910
rect 309542 370908 309548 370910
rect 309612 370908 309618 370972
rect 583520 369460 584960 369700
rect -960 366060 480 366300
rect 309409 360906 309475 360909
rect 309366 360904 309475 360906
rect 309366 360848 309414 360904
rect 309470 360848 309475 360904
rect 309366 360843 309475 360848
rect 309366 360772 309426 360843
rect 309358 360708 309364 360772
rect 309428 360708 309434 360772
rect 276422 359348 276428 359412
rect 276492 359410 276498 359412
rect 282637 359410 282703 359413
rect 276492 359408 282703 359410
rect 276492 359352 282642 359408
rect 282698 359352 282703 359408
rect 276492 359350 282703 359352
rect 276492 359348 276498 359350
rect 282637 359347 282703 359350
rect 276606 359212 276612 359276
rect 276676 359274 276682 359276
rect 285581 359274 285647 359277
rect 286225 359274 286291 359277
rect 276676 359272 286291 359274
rect 276676 359216 285586 359272
rect 285642 359216 286230 359272
rect 286286 359216 286291 359272
rect 276676 359214 286291 359216
rect 276676 359212 276682 359214
rect 285581 359211 285647 359214
rect 286225 359211 286291 359214
rect 583520 357764 584960 358004
rect 306465 355332 306531 355333
rect 306414 355330 306420 355332
rect 306374 355270 306420 355330
rect 306484 355328 306531 355332
rect 306526 355272 306531 355328
rect 306414 355268 306420 355270
rect 306484 355268 306531 355272
rect 306465 355267 306531 355268
rect 274081 354922 274147 354925
rect 274449 354924 274515 354925
rect 275921 354924 275987 354925
rect 274398 354922 274404 354924
rect 274081 354920 274404 354922
rect 274468 354922 274515 354924
rect 274468 354920 274596 354922
rect 274081 354864 274086 354920
rect 274142 354864 274404 354920
rect 274510 354864 274596 354920
rect 274081 354862 274404 354864
rect 274081 354859 274147 354862
rect 274398 354860 274404 354862
rect 274468 354862 274596 354864
rect 274468 354860 274515 354862
rect 275870 354860 275876 354924
rect 275940 354922 275987 354924
rect 290457 354922 290523 354925
rect 291377 354922 291443 354925
rect 295926 354922 295932 354924
rect 275940 354920 276032 354922
rect 275982 354864 276032 354920
rect 275940 354862 276032 354864
rect 290457 354920 295932 354922
rect 290457 354864 290462 354920
rect 290518 354864 291382 354920
rect 291438 354864 295932 354920
rect 290457 354862 295932 354864
rect 275940 354860 275987 354862
rect 274449 354859 274515 354860
rect 275921 354859 275987 354860
rect 290457 354859 290523 354862
rect 291377 354859 291443 354862
rect 295926 354860 295932 354862
rect 295996 354860 296002 354924
rect 297633 354922 297699 354925
rect 299473 354924 299539 354925
rect 298686 354922 298692 354924
rect 297633 354920 298692 354922
rect 297633 354864 297638 354920
rect 297694 354864 298692 354920
rect 297633 354862 298692 354864
rect 297633 354859 297699 354862
rect 298686 354860 298692 354862
rect 298756 354860 298762 354924
rect 299422 354860 299428 354924
rect 299492 354922 299539 354924
rect 299492 354920 299584 354922
rect 299534 354864 299584 354920
rect 299492 354862 299584 354864
rect 299492 354860 299539 354862
rect 299473 354859 299539 354860
rect 292798 353636 292804 353700
rect 292868 353698 292874 353700
rect 294270 353698 294276 353700
rect 292868 353638 294276 353698
rect 292868 353636 292874 353638
rect 294270 353636 294276 353638
rect 294340 353636 294346 353700
rect 270769 352746 270835 352749
rect 272014 352746 272074 352988
rect 270769 352744 272074 352746
rect 270769 352688 270774 352744
rect 270830 352688 272074 352744
rect 270769 352686 272074 352688
rect 270769 352683 270835 352686
rect -960 351780 480 352020
rect 313917 351794 313983 351797
rect 314285 351794 314351 351797
rect 311942 351792 314351 351794
rect 311942 351736 313922 351792
rect 313978 351736 314290 351792
rect 314346 351736 314351 351792
rect 311942 351734 314351 351736
rect 311942 351356 312002 351734
rect 313917 351731 313983 351734
rect 314285 351731 314351 351734
rect 313549 347986 313615 347989
rect 311942 347984 313615 347986
rect 311942 347928 313554 347984
rect 313610 347928 313615 347984
rect 311942 347926 313615 347928
rect 311942 347820 312002 347926
rect 313549 347923 313615 347926
rect 583520 345932 584960 346172
rect 270401 345810 270467 345813
rect 272014 345810 272074 345916
rect 270401 345808 272074 345810
rect 270401 345752 270406 345808
rect 270462 345752 272074 345808
rect 270401 345750 272074 345752
rect 270401 345747 270467 345750
rect 314009 344450 314075 344453
rect 311942 344448 314075 344450
rect 311942 344392 314014 344448
rect 314070 344392 314075 344448
rect 311942 344390 314075 344392
rect 311942 344284 312002 344390
rect 314009 344387 314075 344390
rect 268653 341866 268719 341869
rect 272014 341866 272074 342380
rect 268653 341864 272074 341866
rect 268653 341808 268658 341864
rect 268714 341808 272074 341864
rect 268653 341806 272074 341808
rect 268653 341803 268719 341806
rect 314009 341186 314075 341189
rect 311942 341184 314075 341186
rect 311942 341128 314014 341184
rect 314070 341128 314075 341184
rect 311942 341126 314075 341128
rect 311942 340748 312002 341126
rect 314009 341123 314075 341126
rect 270217 339690 270283 339693
rect 270217 339688 272074 339690
rect 270217 339632 270222 339688
rect 270278 339632 272074 339688
rect 270217 339630 272074 339632
rect 270217 339627 270283 339630
rect 272014 339116 272074 339630
rect 314193 338058 314259 338061
rect 311942 338056 314259 338058
rect 311942 338000 314198 338056
rect 314254 338000 314259 338056
rect 311942 337998 314259 338000
rect -960 337364 480 337604
rect 311942 337484 312002 337998
rect 314193 337995 314259 337998
rect 270677 335474 270743 335477
rect 272014 335474 272074 335580
rect 270677 335472 272074 335474
rect 270677 335416 270682 335472
rect 270738 335416 272074 335472
rect 270677 335414 272074 335416
rect 270677 335411 270743 335414
rect 583520 334236 584960 334476
rect 311390 333844 311450 333948
rect 311382 333780 311388 333844
rect 311452 333780 311458 333844
rect 269389 332346 269455 332349
rect 269389 332344 272074 332346
rect 269389 332288 269394 332344
rect 269450 332288 272074 332344
rect 269389 332286 272074 332288
rect 269389 332283 269455 332286
rect 272014 332044 272074 332286
rect 313733 330714 313799 330717
rect 311942 330712 313799 330714
rect 311942 330656 313738 330712
rect 313794 330656 313799 330712
rect 311942 330654 313799 330656
rect 311942 330412 312002 330654
rect 313733 330651 313799 330654
rect 269389 328402 269455 328405
rect 272014 328402 272074 328508
rect 269389 328400 272074 328402
rect 269389 328344 269394 328400
rect 269450 328344 272074 328400
rect 269389 328342 272074 328344
rect 269389 328339 269455 328342
rect 313825 327042 313891 327045
rect 311942 327040 313891 327042
rect 311942 326984 313830 327040
rect 313886 326984 313891 327040
rect 311942 326982 313891 326984
rect 311942 326876 312002 326982
rect 313825 326979 313891 326982
rect 269389 325274 269455 325277
rect 269389 325272 272074 325274
rect 269389 325216 269394 325272
rect 269450 325216 272074 325272
rect 269389 325214 272074 325216
rect 269389 325211 269455 325214
rect 272014 324972 272074 325214
rect 313641 323642 313707 323645
rect 311942 323640 313707 323642
rect 311942 323584 313646 323640
rect 313702 323584 313707 323640
rect 311942 323582 313707 323584
rect 311942 323340 312002 323582
rect 313641 323579 313707 323582
rect -960 322948 480 323188
rect 583520 322540 584960 322780
rect 270493 322282 270559 322285
rect 270493 322280 272074 322282
rect 270493 322224 270498 322280
rect 270554 322224 272074 322280
rect 270493 322222 272074 322224
rect 270493 322219 270559 322222
rect 272014 321708 272074 322222
rect 313641 320650 313707 320653
rect 314009 320650 314075 320653
rect 311942 320648 314075 320650
rect 311942 320592 313646 320648
rect 313702 320592 314014 320648
rect 314070 320592 314075 320648
rect 311942 320590 314075 320592
rect 311942 320076 312002 320590
rect 313641 320587 313707 320590
rect 314009 320587 314075 320590
rect 270585 318338 270651 318341
rect 270585 318336 272074 318338
rect 270585 318280 270590 318336
rect 270646 318280 272074 318336
rect 270585 318278 272074 318280
rect 270585 318275 270651 318278
rect 272014 318172 272074 318278
rect 311525 317114 311591 317117
rect 311525 317112 311634 317114
rect 311525 317056 311530 317112
rect 311586 317056 311634 317112
rect 311525 317051 311634 317056
rect 311574 316540 311634 317051
rect 274081 316298 274147 316301
rect 275134 316298 275140 316300
rect 274081 316296 275140 316298
rect 274081 316240 274086 316296
rect 274142 316240 275140 316296
rect 274081 316238 275140 316240
rect 274081 316235 274147 316238
rect 275134 316236 275140 316238
rect 275204 316236 275210 316300
rect 292849 316298 292915 316301
rect 294270 316298 294276 316300
rect 292849 316296 294276 316298
rect 292849 316240 292854 316296
rect 292910 316240 294276 316296
rect 292849 316238 294276 316240
rect 292849 316235 292915 316238
rect 294270 316236 294276 316238
rect 294340 316236 294346 316300
rect 295241 316298 295307 316301
rect 295742 316298 295748 316300
rect 295241 316296 295748 316298
rect 295241 316240 295246 316296
rect 295302 316240 295748 316296
rect 295241 316238 295748 316240
rect 295241 316235 295307 316238
rect 295742 316236 295748 316238
rect 295812 316236 295818 316300
rect 300025 316298 300091 316301
rect 300158 316298 300164 316300
rect 300025 316296 300164 316298
rect 300025 316240 300030 316296
rect 300086 316240 300164 316296
rect 300025 316238 300164 316240
rect 300025 316235 300091 316238
rect 300158 316236 300164 316238
rect 300228 316236 300234 316300
rect 309409 316298 309475 316301
rect 309726 316298 309732 316300
rect 309409 316296 309732 316298
rect 309409 316240 309414 316296
rect 309470 316240 309732 316296
rect 309409 316238 309732 316240
rect 309409 316235 309475 316238
rect 309726 316236 309732 316238
rect 309796 316236 309802 316300
rect 290641 315754 290707 315757
rect 293534 315754 293540 315756
rect 290641 315752 293540 315754
rect 290641 315696 290646 315752
rect 290702 315696 293540 315752
rect 290641 315694 293540 315696
rect 290641 315691 290707 315694
rect 293534 315692 293540 315694
rect 293604 315692 293610 315756
rect 276105 315618 276171 315621
rect 306649 315620 306715 315621
rect 276238 315618 276244 315620
rect 276105 315616 276244 315618
rect 276105 315560 276110 315616
rect 276166 315560 276244 315616
rect 276105 315558 276244 315560
rect 276105 315555 276171 315558
rect 276238 315556 276244 315558
rect 276308 315556 276314 315620
rect 306598 315618 306604 315620
rect 306558 315558 306604 315618
rect 306668 315616 306715 315620
rect 306710 315560 306715 315616
rect 306598 315556 306604 315558
rect 306668 315556 306715 315560
rect 306649 315555 306715 315556
rect 287973 313442 288039 313445
rect 288433 313442 288499 313445
rect 295006 313442 295012 313444
rect 287973 313440 295012 313442
rect 287973 313384 287978 313440
rect 288034 313384 288438 313440
rect 288494 313384 295012 313440
rect 287973 313382 295012 313384
rect 287973 313379 288039 313382
rect 288433 313379 288499 313382
rect 295006 313380 295012 313382
rect 295076 313380 295082 313444
rect 280797 313170 280863 313173
rect 299054 313170 299060 313172
rect 280797 313168 299060 313170
rect 280797 313112 280802 313168
rect 280858 313112 299060 313168
rect 280797 313110 299060 313112
rect 280797 313107 280863 313110
rect 299054 313108 299060 313110
rect 299124 313108 299130 313172
rect 285581 312082 285647 312085
rect 286225 312082 286291 312085
rect 293718 312082 293724 312084
rect 285581 312080 293724 312082
rect 285581 312024 285586 312080
rect 285642 312024 286230 312080
rect 286286 312024 293724 312080
rect 285581 312022 293724 312024
rect 285581 312019 285647 312022
rect 286225 312019 286291 312022
rect 293718 312020 293724 312022
rect 293788 312020 293794 312084
rect 583520 310708 584960 310948
rect -960 308668 480 308908
rect 583520 299012 584960 299252
rect -960 294252 480 294492
rect 306557 288554 306623 288557
rect 306741 288554 306807 288557
rect 306557 288552 306807 288554
rect 306557 288496 306562 288552
rect 306618 288496 306746 288552
rect 306802 288496 306807 288552
rect 306557 288494 306807 288496
rect 306557 288491 306623 288494
rect 306741 288491 306807 288494
rect 583520 287316 584960 287556
rect -960 279972 480 280212
rect 275829 276724 275895 276725
rect 275829 276720 275876 276724
rect 275940 276722 275946 276724
rect 275829 276664 275834 276720
rect 275829 276660 275876 276664
rect 275940 276662 275986 276722
rect 275940 276660 275946 276662
rect 306414 276660 306420 276724
rect 306484 276722 306490 276724
rect 306741 276722 306807 276725
rect 306484 276720 306807 276722
rect 306484 276664 306746 276720
rect 306802 276664 306807 276720
rect 306484 276662 306807 276664
rect 306484 276660 306490 276662
rect 275829 276659 275895 276660
rect 306741 276659 306807 276662
rect 583520 275620 584960 275860
rect 295885 275364 295951 275365
rect 295885 275360 295932 275364
rect 295996 275362 296002 275364
rect 295885 275304 295890 275360
rect 295885 275300 295932 275304
rect 295996 275302 296042 275362
rect 295996 275300 296002 275302
rect 295885 275299 295951 275300
rect 276013 272234 276079 272237
rect 276422 272234 276428 272236
rect 276013 272232 276428 272234
rect 276013 272176 276018 272232
rect 276074 272176 276428 272232
rect 276013 272174 276428 272176
rect 276013 272171 276079 272174
rect 276422 272172 276428 272174
rect 276492 272172 276498 272236
rect 276197 272098 276263 272101
rect 276606 272098 276612 272100
rect 276197 272096 276612 272098
rect 276197 272040 276202 272096
rect 276258 272040 276612 272096
rect 276197 272038 276612 272040
rect 276197 272035 276263 272038
rect 276606 272036 276612 272038
rect 276676 272036 276682 272100
rect 27245 270874 27311 270877
rect 27245 270872 27354 270874
rect 27245 270816 27250 270872
rect 27306 270816 27354 270872
rect 27245 270811 27354 270816
rect 27294 270300 27354 270811
rect 315021 270330 315087 270333
rect 315021 270328 318964 270330
rect 315021 270272 315026 270328
rect 315082 270272 318964 270328
rect 315021 270270 318964 270272
rect 315021 270267 315087 270270
rect -960 265556 480 265796
rect 583520 263788 584960 264028
rect 583520 252092 584960 252332
rect -960 251140 480 251380
rect 583520 240396 584960 240636
rect 269021 237418 269087 237421
rect 560845 237418 560911 237421
rect 266524 237416 269087 237418
rect 266524 237360 269026 237416
rect 269082 237360 269087 237416
rect 266524 237358 269087 237360
rect 558716 237416 560911 237418
rect 558716 237360 560850 237416
rect 560906 237360 560911 237416
rect 558716 237358 560911 237360
rect 269021 237355 269087 237358
rect 560845 237355 560911 237358
rect -960 236860 480 237100
rect 24761 234698 24827 234701
rect 315021 234698 315087 234701
rect 24761 234696 26772 234698
rect 24761 234640 24766 234696
rect 24822 234640 26772 234696
rect 24761 234638 26772 234640
rect 315021 234696 318964 234698
rect 315021 234640 315026 234696
rect 315082 234640 318964 234696
rect 315021 234638 318964 234640
rect 24761 234635 24827 234638
rect 315021 234635 315087 234638
rect 583520 228700 584960 228940
rect -960 222444 480 222684
rect 583520 216868 584960 217108
rect -960 208028 480 208268
rect 583520 205172 584960 205412
rect 268009 201786 268075 201789
rect 560845 201786 560911 201789
rect 266524 201784 268075 201786
rect 266524 201728 268014 201784
rect 268070 201728 268075 201784
rect 266524 201726 268075 201728
rect 558716 201784 560911 201786
rect 558716 201728 560850 201784
rect 560906 201728 560911 201784
rect 558716 201726 560911 201728
rect 268009 201723 268075 201726
rect 560845 201723 560911 201726
rect 24945 199066 25011 199069
rect 315021 199066 315087 199069
rect 24945 199064 26772 199066
rect 24945 199008 24950 199064
rect 25006 199008 26772 199064
rect 24945 199006 26772 199008
rect 315021 199064 318964 199066
rect 315021 199008 315026 199064
rect 315082 199008 318964 199064
rect 315021 199006 318964 199008
rect 24945 199003 25011 199006
rect 315021 199003 315087 199006
rect -960 193748 480 193988
rect 583520 193476 584960 193716
rect 583520 181780 584960 182020
rect -960 179332 480 179572
rect 583520 169948 584960 170188
rect 268653 166154 268719 166157
rect 266524 166152 268719 166154
rect 266524 166096 268658 166152
rect 268714 166096 268719 166152
rect 266524 166094 268719 166096
rect 268653 166091 268719 166094
rect -960 164916 480 165156
rect 583520 158252 584960 158492
rect -960 150636 480 150876
rect 583520 146556 584960 146796
rect -960 136220 480 136460
rect 583520 134724 584960 134964
rect 269297 130522 269363 130525
rect 558913 130522 558979 130525
rect 266524 130520 269363 130522
rect 266524 130464 269302 130520
rect 269358 130464 269363 130520
rect 266524 130462 269363 130464
rect 558716 130520 558979 130522
rect 558716 130464 558918 130520
rect 558974 130464 558979 130520
rect 558716 130462 558979 130464
rect 269297 130459 269363 130462
rect 558913 130459 558979 130462
rect 24853 128074 24919 128077
rect 24853 128072 26772 128074
rect 24853 128016 24858 128072
rect 24914 128016 26772 128072
rect 24853 128014 26772 128016
rect 24853 128011 24919 128014
rect 583520 123028 584960 123268
rect -960 121940 480 122180
rect 583520 111332 584960 111572
rect -960 107524 480 107764
rect 583520 99636 584960 99876
rect 269297 95162 269363 95165
rect 560845 95162 560911 95165
rect 266524 95160 269363 95162
rect 266524 95104 269302 95160
rect 269358 95104 269363 95160
rect 266524 95102 269363 95104
rect 558716 95160 560911 95162
rect 558716 95104 560850 95160
rect 560906 95104 560911 95160
rect 558716 95102 560911 95104
rect 269297 95099 269363 95102
rect 560845 95099 560911 95102
rect -960 93108 480 93348
rect 299422 92652 299428 92716
rect 299492 92714 299498 92716
rect 299565 92714 299631 92717
rect 299492 92712 299631 92714
rect 299492 92656 299570 92712
rect 299626 92656 299631 92712
rect 299492 92654 299631 92656
rect 299492 92652 299498 92654
rect 299565 92651 299631 92654
rect 24945 92442 25011 92445
rect 315021 92442 315087 92445
rect 24945 92440 26772 92442
rect 24945 92384 24950 92440
rect 25006 92384 26772 92440
rect 24945 92382 26772 92384
rect 315021 92440 318964 92442
rect 315021 92384 315026 92440
rect 315082 92384 318964 92440
rect 315021 92382 318964 92384
rect 24945 92379 25011 92382
rect 315021 92379 315087 92382
rect 583520 87804 584960 88044
rect -960 78828 480 79068
rect 583520 76108 584960 76348
rect 274398 71980 274404 72044
rect 274468 72042 274474 72044
rect 275185 72042 275251 72045
rect 274468 72040 275251 72042
rect 274468 71984 275190 72040
rect 275246 71984 275251 72040
rect 274468 71982 275251 71984
rect 274468 71980 274474 71982
rect 275185 71979 275251 71982
rect -960 64412 480 64652
rect 583520 64412 584960 64652
rect 583520 52716 584960 52956
rect -960 49996 480 50236
rect 583520 40884 584960 41124
rect -960 35716 480 35956
rect 583520 29188 584960 29428
rect -960 21300 480 21540
rect 583520 17492 584960 17732
rect -960 7020 480 7260
rect 583520 5796 584960 6036
rect 298686 3572 298692 3636
rect 298756 3634 298762 3636
rect 583385 3634 583451 3637
rect 298756 3632 583451 3634
rect 298756 3576 583390 3632
rect 583446 3576 583451 3632
rect 298756 3574 583451 3576
rect 298756 3572 298762 3574
rect 583385 3571 583451 3574
<< via3 >>
rect 299060 700572 299124 700636
rect 275140 699892 275204 699956
rect 310652 609452 310716 609516
rect 295748 586196 295812 586260
rect 292804 586120 292868 586124
rect 292804 586064 292818 586120
rect 292818 586064 292868 586120
rect 292804 586060 292868 586064
rect 306604 585924 306668 585988
rect 310468 566612 310532 566676
rect 293540 546756 293604 546820
rect 310468 511532 310532 511596
rect 309364 504928 309428 504932
rect 309364 504872 309378 504928
rect 309378 504872 309428 504928
rect 309364 504868 309428 504872
rect 309364 497660 309428 497724
rect 309548 497388 309612 497452
rect 309732 484196 309796 484260
rect 309916 484060 309980 484124
rect 309916 473860 309980 473924
rect 310100 463660 310164 463724
rect 309548 458492 309612 458556
rect 310100 458492 310164 458556
rect 309548 445980 309612 446044
rect 310100 445980 310164 446044
rect 310100 435780 310164 435844
rect 310100 435644 310164 435708
rect 309916 432576 309980 432580
rect 309916 432520 309966 432576
rect 309966 432520 309980 432576
rect 309916 432516 309980 432520
rect 309732 422452 309796 422516
rect 309732 415244 309796 415308
rect 309916 414972 309980 415036
rect 309916 412116 309980 412180
rect 309732 401916 309796 401980
rect 309732 394572 309796 394636
rect 309916 394300 309980 394364
rect 309916 391444 309980 391508
rect 293724 384296 293788 384300
rect 293724 384240 293738 384296
rect 293738 384240 293788 384296
rect 293724 384236 293788 384240
rect 295012 382196 295076 382260
rect 276244 382060 276308 382124
rect 300164 381304 300228 381308
rect 300164 381248 300178 381304
rect 300178 381248 300228 381304
rect 300164 381244 300228 381248
rect 309732 381304 309796 381308
rect 309732 381248 309782 381304
rect 309782 381248 309796 381304
rect 309732 381244 309796 381248
rect 309732 374036 309796 374100
rect 309548 373764 309612 373828
rect 309548 370908 309612 370972
rect 309364 360708 309428 360772
rect 276428 359348 276492 359412
rect 276612 359212 276676 359276
rect 306420 355328 306484 355332
rect 306420 355272 306470 355328
rect 306470 355272 306484 355328
rect 306420 355268 306484 355272
rect 274404 354920 274468 354924
rect 274404 354864 274454 354920
rect 274454 354864 274468 354920
rect 274404 354860 274468 354864
rect 275876 354920 275940 354924
rect 275876 354864 275926 354920
rect 275926 354864 275940 354920
rect 275876 354860 275940 354864
rect 295932 354860 295996 354924
rect 298692 354860 298756 354924
rect 299428 354920 299492 354924
rect 299428 354864 299478 354920
rect 299478 354864 299492 354920
rect 299428 354860 299492 354864
rect 292804 353636 292868 353700
rect 294276 353636 294340 353700
rect 311388 333780 311452 333844
rect 275140 316236 275204 316300
rect 294276 316236 294340 316300
rect 295748 316236 295812 316300
rect 300164 316236 300228 316300
rect 309732 316236 309796 316300
rect 293540 315692 293604 315756
rect 276244 315556 276308 315620
rect 306604 315616 306668 315620
rect 306604 315560 306654 315616
rect 306654 315560 306668 315616
rect 306604 315556 306668 315560
rect 295012 313380 295076 313444
rect 299060 313108 299124 313172
rect 293724 312020 293788 312084
rect 275876 276720 275940 276724
rect 275876 276664 275890 276720
rect 275890 276664 275940 276720
rect 275876 276660 275940 276664
rect 306420 276660 306484 276724
rect 295932 275360 295996 275364
rect 295932 275304 295946 275360
rect 295946 275304 295996 275360
rect 295932 275300 295996 275304
rect 276428 272172 276492 272236
rect 276612 272036 276676 272100
rect 299428 92652 299492 92716
rect 274404 71980 274468 72044
rect 298692 3572 298756 3636
<< metal4 >>
rect -8576 711418 -7976 711440
rect -8576 711182 -8394 711418
rect -8158 711182 -7976 711418
rect -8576 711098 -7976 711182
rect -8576 710862 -8394 711098
rect -8158 710862 -7976 711098
rect -8576 -6926 -7976 710862
rect 591900 711418 592500 711440
rect 591900 711182 592082 711418
rect 592318 711182 592500 711418
rect 591900 711098 592500 711182
rect 591900 710862 592082 711098
rect 592318 710862 592500 711098
rect -7636 710478 -7036 710500
rect -7636 710242 -7454 710478
rect -7218 710242 -7036 710478
rect -7636 710158 -7036 710242
rect -7636 709922 -7454 710158
rect -7218 709922 -7036 710158
rect -7636 -5986 -7036 709922
rect 590960 710478 591560 710500
rect 590960 710242 591142 710478
rect 591378 710242 591560 710478
rect 590960 710158 591560 710242
rect 590960 709922 591142 710158
rect 591378 709922 591560 710158
rect -6696 709538 -6096 709560
rect -6696 709302 -6514 709538
rect -6278 709302 -6096 709538
rect -6696 709218 -6096 709302
rect -6696 708982 -6514 709218
rect -6278 708982 -6096 709218
rect -6696 -5046 -6096 708982
rect 590020 709538 590620 709560
rect 590020 709302 590202 709538
rect 590438 709302 590620 709538
rect 590020 709218 590620 709302
rect 590020 708982 590202 709218
rect 590438 708982 590620 709218
rect -5756 708598 -5156 708620
rect -5756 708362 -5574 708598
rect -5338 708362 -5156 708598
rect -5756 708278 -5156 708362
rect -5756 708042 -5574 708278
rect -5338 708042 -5156 708278
rect -5756 -4106 -5156 708042
rect 589080 708598 589680 708620
rect 589080 708362 589262 708598
rect 589498 708362 589680 708598
rect 589080 708278 589680 708362
rect 589080 708042 589262 708278
rect 589498 708042 589680 708278
rect -4816 707658 -4216 707680
rect -4816 707422 -4634 707658
rect -4398 707422 -4216 707658
rect -4816 707338 -4216 707422
rect -4816 707102 -4634 707338
rect -4398 707102 -4216 707338
rect -4816 -3166 -4216 707102
rect 588140 707658 588740 707680
rect 588140 707422 588322 707658
rect 588558 707422 588740 707658
rect 588140 707338 588740 707422
rect 588140 707102 588322 707338
rect 588558 707102 588740 707338
rect -3876 706718 -3276 706740
rect -3876 706482 -3694 706718
rect -3458 706482 -3276 706718
rect -3876 706398 -3276 706482
rect -3876 706162 -3694 706398
rect -3458 706162 -3276 706398
rect -3876 -2226 -3276 706162
rect 587200 706718 587800 706740
rect 587200 706482 587382 706718
rect 587618 706482 587800 706718
rect 587200 706398 587800 706482
rect 587200 706162 587382 706398
rect 587618 706162 587800 706398
rect -2936 705778 -2336 705800
rect -2936 705542 -2754 705778
rect -2518 705542 -2336 705778
rect -2936 705458 -2336 705542
rect -2936 705222 -2754 705458
rect -2518 705222 -2336 705458
rect -2936 668454 -2336 705222
rect -2936 668218 -2754 668454
rect -2518 668218 -2336 668454
rect -2936 668134 -2336 668218
rect -2936 667898 -2754 668134
rect -2518 667898 -2336 668134
rect -2936 632454 -2336 667898
rect -2936 632218 -2754 632454
rect -2518 632218 -2336 632454
rect -2936 632134 -2336 632218
rect -2936 631898 -2754 632134
rect -2518 631898 -2336 632134
rect -2936 596454 -2336 631898
rect -2936 596218 -2754 596454
rect -2518 596218 -2336 596454
rect -2936 596134 -2336 596218
rect -2936 595898 -2754 596134
rect -2518 595898 -2336 596134
rect -2936 560454 -2336 595898
rect -2936 560218 -2754 560454
rect -2518 560218 -2336 560454
rect -2936 560134 -2336 560218
rect -2936 559898 -2754 560134
rect -2518 559898 -2336 560134
rect -2936 524454 -2336 559898
rect -2936 524218 -2754 524454
rect -2518 524218 -2336 524454
rect -2936 524134 -2336 524218
rect -2936 523898 -2754 524134
rect -2518 523898 -2336 524134
rect -2936 488454 -2336 523898
rect -2936 488218 -2754 488454
rect -2518 488218 -2336 488454
rect -2936 488134 -2336 488218
rect -2936 487898 -2754 488134
rect -2518 487898 -2336 488134
rect -2936 452454 -2336 487898
rect -2936 452218 -2754 452454
rect -2518 452218 -2336 452454
rect -2936 452134 -2336 452218
rect -2936 451898 -2754 452134
rect -2518 451898 -2336 452134
rect -2936 416454 -2336 451898
rect -2936 416218 -2754 416454
rect -2518 416218 -2336 416454
rect -2936 416134 -2336 416218
rect -2936 415898 -2754 416134
rect -2518 415898 -2336 416134
rect -2936 380454 -2336 415898
rect -2936 380218 -2754 380454
rect -2518 380218 -2336 380454
rect -2936 380134 -2336 380218
rect -2936 379898 -2754 380134
rect -2518 379898 -2336 380134
rect -2936 344454 -2336 379898
rect -2936 344218 -2754 344454
rect -2518 344218 -2336 344454
rect -2936 344134 -2336 344218
rect -2936 343898 -2754 344134
rect -2518 343898 -2336 344134
rect -2936 308454 -2336 343898
rect -2936 308218 -2754 308454
rect -2518 308218 -2336 308454
rect -2936 308134 -2336 308218
rect -2936 307898 -2754 308134
rect -2518 307898 -2336 308134
rect -2936 272454 -2336 307898
rect -2936 272218 -2754 272454
rect -2518 272218 -2336 272454
rect -2936 272134 -2336 272218
rect -2936 271898 -2754 272134
rect -2518 271898 -2336 272134
rect -2936 236454 -2336 271898
rect -2936 236218 -2754 236454
rect -2518 236218 -2336 236454
rect -2936 236134 -2336 236218
rect -2936 235898 -2754 236134
rect -2518 235898 -2336 236134
rect -2936 200454 -2336 235898
rect -2936 200218 -2754 200454
rect -2518 200218 -2336 200454
rect -2936 200134 -2336 200218
rect -2936 199898 -2754 200134
rect -2518 199898 -2336 200134
rect -2936 164454 -2336 199898
rect -2936 164218 -2754 164454
rect -2518 164218 -2336 164454
rect -2936 164134 -2336 164218
rect -2936 163898 -2754 164134
rect -2518 163898 -2336 164134
rect -2936 128454 -2336 163898
rect -2936 128218 -2754 128454
rect -2518 128218 -2336 128454
rect -2936 128134 -2336 128218
rect -2936 127898 -2754 128134
rect -2518 127898 -2336 128134
rect -2936 92454 -2336 127898
rect -2936 92218 -2754 92454
rect -2518 92218 -2336 92454
rect -2936 92134 -2336 92218
rect -2936 91898 -2754 92134
rect -2518 91898 -2336 92134
rect -2936 56454 -2336 91898
rect -2936 56218 -2754 56454
rect -2518 56218 -2336 56454
rect -2936 56134 -2336 56218
rect -2936 55898 -2754 56134
rect -2518 55898 -2336 56134
rect -2936 20454 -2336 55898
rect -2936 20218 -2754 20454
rect -2518 20218 -2336 20454
rect -2936 20134 -2336 20218
rect -2936 19898 -2754 20134
rect -2518 19898 -2336 20134
rect -2936 -1286 -2336 19898
rect -1996 704838 -1396 704860
rect -1996 704602 -1814 704838
rect -1578 704602 -1396 704838
rect -1996 704518 -1396 704602
rect -1996 704282 -1814 704518
rect -1578 704282 -1396 704518
rect -1996 686454 -1396 704282
rect -1996 686218 -1814 686454
rect -1578 686218 -1396 686454
rect -1996 686134 -1396 686218
rect -1996 685898 -1814 686134
rect -1578 685898 -1396 686134
rect -1996 650454 -1396 685898
rect -1996 650218 -1814 650454
rect -1578 650218 -1396 650454
rect -1996 650134 -1396 650218
rect -1996 649898 -1814 650134
rect -1578 649898 -1396 650134
rect -1996 614454 -1396 649898
rect -1996 614218 -1814 614454
rect -1578 614218 -1396 614454
rect -1996 614134 -1396 614218
rect -1996 613898 -1814 614134
rect -1578 613898 -1396 614134
rect -1996 578454 -1396 613898
rect -1996 578218 -1814 578454
rect -1578 578218 -1396 578454
rect -1996 578134 -1396 578218
rect -1996 577898 -1814 578134
rect -1578 577898 -1396 578134
rect -1996 542454 -1396 577898
rect -1996 542218 -1814 542454
rect -1578 542218 -1396 542454
rect -1996 542134 -1396 542218
rect -1996 541898 -1814 542134
rect -1578 541898 -1396 542134
rect -1996 506454 -1396 541898
rect -1996 506218 -1814 506454
rect -1578 506218 -1396 506454
rect -1996 506134 -1396 506218
rect -1996 505898 -1814 506134
rect -1578 505898 -1396 506134
rect -1996 470454 -1396 505898
rect -1996 470218 -1814 470454
rect -1578 470218 -1396 470454
rect -1996 470134 -1396 470218
rect -1996 469898 -1814 470134
rect -1578 469898 -1396 470134
rect -1996 434454 -1396 469898
rect -1996 434218 -1814 434454
rect -1578 434218 -1396 434454
rect -1996 434134 -1396 434218
rect -1996 433898 -1814 434134
rect -1578 433898 -1396 434134
rect -1996 398454 -1396 433898
rect -1996 398218 -1814 398454
rect -1578 398218 -1396 398454
rect -1996 398134 -1396 398218
rect -1996 397898 -1814 398134
rect -1578 397898 -1396 398134
rect -1996 362454 -1396 397898
rect -1996 362218 -1814 362454
rect -1578 362218 -1396 362454
rect -1996 362134 -1396 362218
rect -1996 361898 -1814 362134
rect -1578 361898 -1396 362134
rect -1996 326454 -1396 361898
rect -1996 326218 -1814 326454
rect -1578 326218 -1396 326454
rect -1996 326134 -1396 326218
rect -1996 325898 -1814 326134
rect -1578 325898 -1396 326134
rect -1996 290454 -1396 325898
rect -1996 290218 -1814 290454
rect -1578 290218 -1396 290454
rect -1996 290134 -1396 290218
rect -1996 289898 -1814 290134
rect -1578 289898 -1396 290134
rect -1996 254454 -1396 289898
rect -1996 254218 -1814 254454
rect -1578 254218 -1396 254454
rect -1996 254134 -1396 254218
rect -1996 253898 -1814 254134
rect -1578 253898 -1396 254134
rect -1996 218454 -1396 253898
rect -1996 218218 -1814 218454
rect -1578 218218 -1396 218454
rect -1996 218134 -1396 218218
rect -1996 217898 -1814 218134
rect -1578 217898 -1396 218134
rect -1996 182454 -1396 217898
rect -1996 182218 -1814 182454
rect -1578 182218 -1396 182454
rect -1996 182134 -1396 182218
rect -1996 181898 -1814 182134
rect -1578 181898 -1396 182134
rect -1996 146454 -1396 181898
rect -1996 146218 -1814 146454
rect -1578 146218 -1396 146454
rect -1996 146134 -1396 146218
rect -1996 145898 -1814 146134
rect -1578 145898 -1396 146134
rect -1996 110454 -1396 145898
rect -1996 110218 -1814 110454
rect -1578 110218 -1396 110454
rect -1996 110134 -1396 110218
rect -1996 109898 -1814 110134
rect -1578 109898 -1396 110134
rect -1996 74454 -1396 109898
rect -1996 74218 -1814 74454
rect -1578 74218 -1396 74454
rect -1996 74134 -1396 74218
rect -1996 73898 -1814 74134
rect -1578 73898 -1396 74134
rect -1996 38454 -1396 73898
rect -1996 38218 -1814 38454
rect -1578 38218 -1396 38454
rect -1996 38134 -1396 38218
rect -1996 37898 -1814 38134
rect -1578 37898 -1396 38134
rect -1996 2454 -1396 37898
rect -1996 2218 -1814 2454
rect -1578 2218 -1396 2454
rect -1996 2134 -1396 2218
rect -1996 1898 -1814 2134
rect -1578 1898 -1396 2134
rect -1996 -346 -1396 1898
rect -1996 -582 -1814 -346
rect -1578 -582 -1396 -346
rect -1996 -666 -1396 -582
rect -1996 -902 -1814 -666
rect -1578 -902 -1396 -666
rect -1996 -924 -1396 -902
rect 804 704838 1404 705800
rect 804 704602 986 704838
rect 1222 704602 1404 704838
rect 804 704518 1404 704602
rect 804 704282 986 704518
rect 1222 704282 1404 704518
rect 804 686454 1404 704282
rect 804 686218 986 686454
rect 1222 686218 1404 686454
rect 804 686134 1404 686218
rect 804 685898 986 686134
rect 1222 685898 1404 686134
rect 804 650454 1404 685898
rect 804 650218 986 650454
rect 1222 650218 1404 650454
rect 804 650134 1404 650218
rect 804 649898 986 650134
rect 1222 649898 1404 650134
rect 804 614454 1404 649898
rect 804 614218 986 614454
rect 1222 614218 1404 614454
rect 804 614134 1404 614218
rect 804 613898 986 614134
rect 1222 613898 1404 614134
rect 804 578454 1404 613898
rect 804 578218 986 578454
rect 1222 578218 1404 578454
rect 804 578134 1404 578218
rect 804 577898 986 578134
rect 1222 577898 1404 578134
rect 804 542454 1404 577898
rect 804 542218 986 542454
rect 1222 542218 1404 542454
rect 804 542134 1404 542218
rect 804 541898 986 542134
rect 1222 541898 1404 542134
rect 804 506454 1404 541898
rect 804 506218 986 506454
rect 1222 506218 1404 506454
rect 804 506134 1404 506218
rect 804 505898 986 506134
rect 1222 505898 1404 506134
rect 804 470454 1404 505898
rect 804 470218 986 470454
rect 1222 470218 1404 470454
rect 804 470134 1404 470218
rect 804 469898 986 470134
rect 1222 469898 1404 470134
rect 804 434454 1404 469898
rect 804 434218 986 434454
rect 1222 434218 1404 434454
rect 804 434134 1404 434218
rect 804 433898 986 434134
rect 1222 433898 1404 434134
rect 804 398454 1404 433898
rect 804 398218 986 398454
rect 1222 398218 1404 398454
rect 804 398134 1404 398218
rect 804 397898 986 398134
rect 1222 397898 1404 398134
rect 804 362454 1404 397898
rect 804 362218 986 362454
rect 1222 362218 1404 362454
rect 804 362134 1404 362218
rect 804 361898 986 362134
rect 1222 361898 1404 362134
rect 804 326454 1404 361898
rect 804 326218 986 326454
rect 1222 326218 1404 326454
rect 804 326134 1404 326218
rect 804 325898 986 326134
rect 1222 325898 1404 326134
rect 804 290454 1404 325898
rect 804 290218 986 290454
rect 1222 290218 1404 290454
rect 804 290134 1404 290218
rect 804 289898 986 290134
rect 1222 289898 1404 290134
rect 804 254454 1404 289898
rect 804 254218 986 254454
rect 1222 254218 1404 254454
rect 804 254134 1404 254218
rect 804 253898 986 254134
rect 1222 253898 1404 254134
rect 804 218454 1404 253898
rect 804 218218 986 218454
rect 1222 218218 1404 218454
rect 804 218134 1404 218218
rect 804 217898 986 218134
rect 1222 217898 1404 218134
rect 804 182454 1404 217898
rect 804 182218 986 182454
rect 1222 182218 1404 182454
rect 804 182134 1404 182218
rect 804 181898 986 182134
rect 1222 181898 1404 182134
rect 804 146454 1404 181898
rect 804 146218 986 146454
rect 1222 146218 1404 146454
rect 804 146134 1404 146218
rect 804 145898 986 146134
rect 1222 145898 1404 146134
rect 804 110454 1404 145898
rect 804 110218 986 110454
rect 1222 110218 1404 110454
rect 804 110134 1404 110218
rect 804 109898 986 110134
rect 1222 109898 1404 110134
rect 804 74454 1404 109898
rect 804 74218 986 74454
rect 1222 74218 1404 74454
rect 804 74134 1404 74218
rect 804 73898 986 74134
rect 1222 73898 1404 74134
rect 804 38454 1404 73898
rect 804 38218 986 38454
rect 1222 38218 1404 38454
rect 804 38134 1404 38218
rect 804 37898 986 38134
rect 1222 37898 1404 38134
rect 804 2454 1404 37898
rect 804 2218 986 2454
rect 1222 2218 1404 2454
rect 804 2134 1404 2218
rect 804 1898 986 2134
rect 1222 1898 1404 2134
rect 804 -346 1404 1898
rect 804 -582 986 -346
rect 1222 -582 1404 -346
rect 804 -666 1404 -582
rect 804 -902 986 -666
rect 1222 -902 1404 -666
rect -2936 -1522 -2754 -1286
rect -2518 -1522 -2336 -1286
rect -2936 -1606 -2336 -1522
rect -2936 -1842 -2754 -1606
rect -2518 -1842 -2336 -1606
rect -2936 -1864 -2336 -1842
rect 804 -1864 1404 -902
rect 18804 705778 19404 705800
rect 18804 705542 18986 705778
rect 19222 705542 19404 705778
rect 18804 705458 19404 705542
rect 18804 705222 18986 705458
rect 19222 705222 19404 705458
rect 18804 668454 19404 705222
rect 18804 668218 18986 668454
rect 19222 668218 19404 668454
rect 18804 668134 19404 668218
rect 18804 667898 18986 668134
rect 19222 667898 19404 668134
rect 18804 632454 19404 667898
rect 18804 632218 18986 632454
rect 19222 632218 19404 632454
rect 18804 632134 19404 632218
rect 18804 631898 18986 632134
rect 19222 631898 19404 632134
rect 18804 596454 19404 631898
rect 18804 596218 18986 596454
rect 19222 596218 19404 596454
rect 18804 596134 19404 596218
rect 18804 595898 18986 596134
rect 19222 595898 19404 596134
rect 18804 560454 19404 595898
rect 36804 704838 37404 705800
rect 36804 704602 36986 704838
rect 37222 704602 37404 704838
rect 36804 704518 37404 704602
rect 36804 704282 36986 704518
rect 37222 704282 37404 704518
rect 36804 686454 37404 704282
rect 36804 686218 36986 686454
rect 37222 686218 37404 686454
rect 36804 686134 37404 686218
rect 36804 685898 36986 686134
rect 37222 685898 37404 686134
rect 36804 650454 37404 685898
rect 36804 650218 36986 650454
rect 37222 650218 37404 650454
rect 36804 650134 37404 650218
rect 36804 649898 36986 650134
rect 37222 649898 37404 650134
rect 36804 614454 37404 649898
rect 36804 614218 36986 614454
rect 37222 614218 37404 614454
rect 36804 614134 37404 614218
rect 36804 613898 36986 614134
rect 37222 613898 37404 614134
rect 36804 584916 37404 613898
rect 54804 705778 55404 705800
rect 54804 705542 54986 705778
rect 55222 705542 55404 705778
rect 54804 705458 55404 705542
rect 54804 705222 54986 705458
rect 55222 705222 55404 705458
rect 54804 668454 55404 705222
rect 54804 668218 54986 668454
rect 55222 668218 55404 668454
rect 54804 668134 55404 668218
rect 54804 667898 54986 668134
rect 55222 667898 55404 668134
rect 54804 632454 55404 667898
rect 54804 632218 54986 632454
rect 55222 632218 55404 632454
rect 54804 632134 55404 632218
rect 54804 631898 54986 632134
rect 55222 631898 55404 632134
rect 54804 596454 55404 631898
rect 54804 596218 54986 596454
rect 55222 596218 55404 596454
rect 54804 596134 55404 596218
rect 54804 595898 54986 596134
rect 55222 595898 55404 596134
rect 54804 584916 55404 595898
rect 72804 704838 73404 705800
rect 72804 704602 72986 704838
rect 73222 704602 73404 704838
rect 72804 704518 73404 704602
rect 72804 704282 72986 704518
rect 73222 704282 73404 704518
rect 72804 686454 73404 704282
rect 72804 686218 72986 686454
rect 73222 686218 73404 686454
rect 72804 686134 73404 686218
rect 72804 685898 72986 686134
rect 73222 685898 73404 686134
rect 72804 650454 73404 685898
rect 72804 650218 72986 650454
rect 73222 650218 73404 650454
rect 72804 650134 73404 650218
rect 72804 649898 72986 650134
rect 73222 649898 73404 650134
rect 72804 614454 73404 649898
rect 72804 614218 72986 614454
rect 73222 614218 73404 614454
rect 72804 614134 73404 614218
rect 72804 613898 72986 614134
rect 73222 613898 73404 614134
rect 72804 584916 73404 613898
rect 90804 705778 91404 705800
rect 90804 705542 90986 705778
rect 91222 705542 91404 705778
rect 90804 705458 91404 705542
rect 90804 705222 90986 705458
rect 91222 705222 91404 705458
rect 90804 668454 91404 705222
rect 90804 668218 90986 668454
rect 91222 668218 91404 668454
rect 90804 668134 91404 668218
rect 90804 667898 90986 668134
rect 91222 667898 91404 668134
rect 90804 632454 91404 667898
rect 90804 632218 90986 632454
rect 91222 632218 91404 632454
rect 90804 632134 91404 632218
rect 90804 631898 90986 632134
rect 91222 631898 91404 632134
rect 90804 596454 91404 631898
rect 90804 596218 90986 596454
rect 91222 596218 91404 596454
rect 90804 596134 91404 596218
rect 90804 595898 90986 596134
rect 91222 595898 91404 596134
rect 90804 584916 91404 595898
rect 108804 704838 109404 705800
rect 108804 704602 108986 704838
rect 109222 704602 109404 704838
rect 108804 704518 109404 704602
rect 108804 704282 108986 704518
rect 109222 704282 109404 704518
rect 108804 686454 109404 704282
rect 108804 686218 108986 686454
rect 109222 686218 109404 686454
rect 108804 686134 109404 686218
rect 108804 685898 108986 686134
rect 109222 685898 109404 686134
rect 108804 650454 109404 685898
rect 108804 650218 108986 650454
rect 109222 650218 109404 650454
rect 108804 650134 109404 650218
rect 108804 649898 108986 650134
rect 109222 649898 109404 650134
rect 108804 614454 109404 649898
rect 108804 614218 108986 614454
rect 109222 614218 109404 614454
rect 108804 614134 109404 614218
rect 108804 613898 108986 614134
rect 109222 613898 109404 614134
rect 108804 584916 109404 613898
rect 126804 705778 127404 705800
rect 126804 705542 126986 705778
rect 127222 705542 127404 705778
rect 126804 705458 127404 705542
rect 126804 705222 126986 705458
rect 127222 705222 127404 705458
rect 126804 668454 127404 705222
rect 126804 668218 126986 668454
rect 127222 668218 127404 668454
rect 126804 668134 127404 668218
rect 126804 667898 126986 668134
rect 127222 667898 127404 668134
rect 126804 632454 127404 667898
rect 126804 632218 126986 632454
rect 127222 632218 127404 632454
rect 126804 632134 127404 632218
rect 126804 631898 126986 632134
rect 127222 631898 127404 632134
rect 126804 596454 127404 631898
rect 126804 596218 126986 596454
rect 127222 596218 127404 596454
rect 126804 596134 127404 596218
rect 126804 595898 126986 596134
rect 127222 595898 127404 596134
rect 126804 584916 127404 595898
rect 144804 704838 145404 705800
rect 144804 704602 144986 704838
rect 145222 704602 145404 704838
rect 144804 704518 145404 704602
rect 144804 704282 144986 704518
rect 145222 704282 145404 704518
rect 144804 686454 145404 704282
rect 144804 686218 144986 686454
rect 145222 686218 145404 686454
rect 144804 686134 145404 686218
rect 144804 685898 144986 686134
rect 145222 685898 145404 686134
rect 144804 650454 145404 685898
rect 144804 650218 144986 650454
rect 145222 650218 145404 650454
rect 144804 650134 145404 650218
rect 144804 649898 144986 650134
rect 145222 649898 145404 650134
rect 144804 614454 145404 649898
rect 144804 614218 144986 614454
rect 145222 614218 145404 614454
rect 144804 614134 145404 614218
rect 144804 613898 144986 614134
rect 145222 613898 145404 614134
rect 144804 584916 145404 613898
rect 162804 705778 163404 705800
rect 162804 705542 162986 705778
rect 163222 705542 163404 705778
rect 162804 705458 163404 705542
rect 162804 705222 162986 705458
rect 163222 705222 163404 705458
rect 162804 668454 163404 705222
rect 162804 668218 162986 668454
rect 163222 668218 163404 668454
rect 162804 668134 163404 668218
rect 162804 667898 162986 668134
rect 163222 667898 163404 668134
rect 162804 632454 163404 667898
rect 162804 632218 162986 632454
rect 163222 632218 163404 632454
rect 162804 632134 163404 632218
rect 162804 631898 162986 632134
rect 163222 631898 163404 632134
rect 162804 596454 163404 631898
rect 162804 596218 162986 596454
rect 163222 596218 163404 596454
rect 162804 596134 163404 596218
rect 162804 595898 162986 596134
rect 163222 595898 163404 596134
rect 162804 584916 163404 595898
rect 180804 704838 181404 705800
rect 180804 704602 180986 704838
rect 181222 704602 181404 704838
rect 180804 704518 181404 704602
rect 180804 704282 180986 704518
rect 181222 704282 181404 704518
rect 180804 686454 181404 704282
rect 180804 686218 180986 686454
rect 181222 686218 181404 686454
rect 180804 686134 181404 686218
rect 180804 685898 180986 686134
rect 181222 685898 181404 686134
rect 180804 650454 181404 685898
rect 180804 650218 180986 650454
rect 181222 650218 181404 650454
rect 180804 650134 181404 650218
rect 180804 649898 180986 650134
rect 181222 649898 181404 650134
rect 180804 614454 181404 649898
rect 180804 614218 180986 614454
rect 181222 614218 181404 614454
rect 180804 614134 181404 614218
rect 180804 613898 180986 614134
rect 181222 613898 181404 614134
rect 180804 584916 181404 613898
rect 198804 705778 199404 705800
rect 198804 705542 198986 705778
rect 199222 705542 199404 705778
rect 198804 705458 199404 705542
rect 198804 705222 198986 705458
rect 199222 705222 199404 705458
rect 198804 668454 199404 705222
rect 198804 668218 198986 668454
rect 199222 668218 199404 668454
rect 198804 668134 199404 668218
rect 198804 667898 198986 668134
rect 199222 667898 199404 668134
rect 198804 632454 199404 667898
rect 198804 632218 198986 632454
rect 199222 632218 199404 632454
rect 198804 632134 199404 632218
rect 198804 631898 198986 632134
rect 199222 631898 199404 632134
rect 198804 596454 199404 631898
rect 198804 596218 198986 596454
rect 199222 596218 199404 596454
rect 198804 596134 199404 596218
rect 198804 595898 198986 596134
rect 199222 595898 199404 596134
rect 198804 584916 199404 595898
rect 216804 704838 217404 705800
rect 216804 704602 216986 704838
rect 217222 704602 217404 704838
rect 216804 704518 217404 704602
rect 216804 704282 216986 704518
rect 217222 704282 217404 704518
rect 216804 686454 217404 704282
rect 216804 686218 216986 686454
rect 217222 686218 217404 686454
rect 216804 686134 217404 686218
rect 216804 685898 216986 686134
rect 217222 685898 217404 686134
rect 216804 650454 217404 685898
rect 216804 650218 216986 650454
rect 217222 650218 217404 650454
rect 216804 650134 217404 650218
rect 216804 649898 216986 650134
rect 217222 649898 217404 650134
rect 216804 614454 217404 649898
rect 216804 614218 216986 614454
rect 217222 614218 217404 614454
rect 216804 614134 217404 614218
rect 216804 613898 216986 614134
rect 217222 613898 217404 614134
rect 216804 584916 217404 613898
rect 234804 705778 235404 705800
rect 234804 705542 234986 705778
rect 235222 705542 235404 705778
rect 234804 705458 235404 705542
rect 234804 705222 234986 705458
rect 235222 705222 235404 705458
rect 234804 668454 235404 705222
rect 234804 668218 234986 668454
rect 235222 668218 235404 668454
rect 234804 668134 235404 668218
rect 234804 667898 234986 668134
rect 235222 667898 235404 668134
rect 234804 632454 235404 667898
rect 234804 632218 234986 632454
rect 235222 632218 235404 632454
rect 234804 632134 235404 632218
rect 234804 631898 234986 632134
rect 235222 631898 235404 632134
rect 234804 596454 235404 631898
rect 234804 596218 234986 596454
rect 235222 596218 235404 596454
rect 234804 596134 235404 596218
rect 234804 595898 234986 596134
rect 235222 595898 235404 596134
rect 234804 584916 235404 595898
rect 252804 704838 253404 705800
rect 252804 704602 252986 704838
rect 253222 704602 253404 704838
rect 252804 704518 253404 704602
rect 252804 704282 252986 704518
rect 253222 704282 253404 704518
rect 252804 686454 253404 704282
rect 252804 686218 252986 686454
rect 253222 686218 253404 686454
rect 252804 686134 253404 686218
rect 252804 685898 252986 686134
rect 253222 685898 253404 686134
rect 252804 650454 253404 685898
rect 252804 650218 252986 650454
rect 253222 650218 253404 650454
rect 252804 650134 253404 650218
rect 252804 649898 252986 650134
rect 253222 649898 253404 650134
rect 252804 614454 253404 649898
rect 252804 614218 252986 614454
rect 253222 614218 253404 614454
rect 252804 614134 253404 614218
rect 252804 613898 252986 614134
rect 253222 613898 253404 614134
rect 252804 584916 253404 613898
rect 270804 705778 271404 705800
rect 270804 705542 270986 705778
rect 271222 705542 271404 705778
rect 270804 705458 271404 705542
rect 270804 705222 270986 705458
rect 271222 705222 271404 705458
rect 270804 668454 271404 705222
rect 288804 704838 289404 705800
rect 288804 704602 288986 704838
rect 289222 704602 289404 704838
rect 288804 704518 289404 704602
rect 288804 704282 288986 704518
rect 289222 704282 289404 704518
rect 275139 699956 275205 699957
rect 275139 699892 275140 699956
rect 275204 699892 275205 699956
rect 275139 699891 275205 699892
rect 270804 668218 270986 668454
rect 271222 668218 271404 668454
rect 270804 668134 271404 668218
rect 270804 667898 270986 668134
rect 271222 667898 271404 668134
rect 270804 632454 271404 667898
rect 270804 632218 270986 632454
rect 271222 632218 271404 632454
rect 270804 632134 271404 632218
rect 270804 631898 270986 632134
rect 271222 631898 271404 632134
rect 270804 596454 271404 631898
rect 270804 596218 270986 596454
rect 271222 596218 271404 596454
rect 270804 596134 271404 596218
rect 270804 595898 270986 596134
rect 271222 595898 271404 596134
rect 262128 578454 262448 578476
rect 262128 578218 262170 578454
rect 262406 578218 262448 578454
rect 262128 578134 262448 578218
rect 262128 577898 262170 578134
rect 262406 577898 262448 578134
rect 262128 577876 262448 577898
rect 18804 560218 18986 560454
rect 19222 560218 19404 560454
rect 18804 560134 19404 560218
rect 18804 559898 18986 560134
rect 19222 559898 19404 560134
rect 18804 524454 19404 559898
rect 246768 560454 247088 560476
rect 246768 560218 246810 560454
rect 247046 560218 247088 560454
rect 246768 560134 247088 560218
rect 246768 559898 246810 560134
rect 247046 559898 247088 560134
rect 246768 559876 247088 559898
rect 270804 560454 271404 595898
rect 270804 560218 270986 560454
rect 271222 560218 271404 560454
rect 270804 560134 271404 560218
rect 270804 559898 270986 560134
rect 271222 559898 271404 560134
rect 262128 542454 262448 542476
rect 262128 542218 262170 542454
rect 262406 542218 262448 542454
rect 262128 542134 262448 542218
rect 262128 541898 262170 542134
rect 262406 541898 262448 542134
rect 262128 541876 262448 541898
rect 18804 524218 18986 524454
rect 19222 524218 19404 524454
rect 18804 524134 19404 524218
rect 18804 523898 18986 524134
rect 19222 523898 19404 524134
rect 18804 488454 19404 523898
rect 246768 524454 247088 524476
rect 246768 524218 246810 524454
rect 247046 524218 247088 524454
rect 246768 524134 247088 524218
rect 246768 523898 246810 524134
rect 247046 523898 247088 524134
rect 246768 523876 247088 523898
rect 270804 524454 271404 559898
rect 270804 524218 270986 524454
rect 271222 524218 271404 524454
rect 270804 524134 271404 524218
rect 270804 523898 270986 524134
rect 271222 523898 271404 524134
rect 262128 506454 262448 506476
rect 262128 506218 262170 506454
rect 262406 506218 262448 506454
rect 262128 506134 262448 506218
rect 262128 505898 262170 506134
rect 262406 505898 262448 506134
rect 262128 505876 262448 505898
rect 18804 488218 18986 488454
rect 19222 488218 19404 488454
rect 18804 488134 19404 488218
rect 18804 487898 18986 488134
rect 19222 487898 19404 488134
rect 18804 452454 19404 487898
rect 246768 488454 247088 488476
rect 246768 488218 246810 488454
rect 247046 488218 247088 488454
rect 246768 488134 247088 488218
rect 246768 487898 246810 488134
rect 247046 487898 247088 488134
rect 246768 487876 247088 487898
rect 270804 488454 271404 523898
rect 270804 488218 270986 488454
rect 271222 488218 271404 488454
rect 270804 488134 271404 488218
rect 270804 487898 270986 488134
rect 271222 487898 271404 488134
rect 262128 470454 262448 470476
rect 262128 470218 262170 470454
rect 262406 470218 262448 470454
rect 262128 470134 262448 470218
rect 262128 469898 262170 470134
rect 262406 469898 262448 470134
rect 262128 469876 262448 469898
rect 18804 452218 18986 452454
rect 19222 452218 19404 452454
rect 18804 452134 19404 452218
rect 18804 451898 18986 452134
rect 19222 451898 19404 452134
rect 18804 416454 19404 451898
rect 246768 452454 247088 452476
rect 246768 452218 246810 452454
rect 247046 452218 247088 452454
rect 246768 452134 247088 452218
rect 246768 451898 246810 452134
rect 247046 451898 247088 452134
rect 246768 451876 247088 451898
rect 270804 452454 271404 487898
rect 270804 452218 270986 452454
rect 271222 452218 271404 452454
rect 270804 452134 271404 452218
rect 270804 451898 270986 452134
rect 271222 451898 271404 452134
rect 262128 434454 262448 434476
rect 262128 434218 262170 434454
rect 262406 434218 262448 434454
rect 262128 434134 262448 434218
rect 262128 433898 262170 434134
rect 262406 433898 262448 434134
rect 262128 433876 262448 433898
rect 18804 416218 18986 416454
rect 19222 416218 19404 416454
rect 18804 416134 19404 416218
rect 18804 415898 18986 416134
rect 19222 415898 19404 416134
rect 18804 380454 19404 415898
rect 246768 416454 247088 416476
rect 246768 416218 246810 416454
rect 247046 416218 247088 416454
rect 246768 416134 247088 416218
rect 246768 415898 246810 416134
rect 247046 415898 247088 416134
rect 246768 415876 247088 415898
rect 270804 416454 271404 451898
rect 270804 416218 270986 416454
rect 271222 416218 271404 416454
rect 270804 416134 271404 416218
rect 270804 415898 270986 416134
rect 271222 415898 271404 416134
rect 262128 398454 262448 398476
rect 262128 398218 262170 398454
rect 262406 398218 262448 398454
rect 262128 398134 262448 398218
rect 262128 397898 262170 398134
rect 262406 397898 262448 398134
rect 262128 397876 262448 397898
rect 18804 380218 18986 380454
rect 19222 380218 19404 380454
rect 18804 380134 19404 380218
rect 18804 379898 18986 380134
rect 19222 379898 19404 380134
rect 18804 344454 19404 379898
rect 18804 344218 18986 344454
rect 19222 344218 19404 344454
rect 18804 344134 19404 344218
rect 18804 343898 18986 344134
rect 19222 343898 19404 344134
rect 18804 308454 19404 343898
rect 18804 308218 18986 308454
rect 19222 308218 19404 308454
rect 18804 308134 19404 308218
rect 18804 307898 18986 308134
rect 19222 307898 19404 308134
rect 18804 272454 19404 307898
rect 36804 362454 37404 382916
rect 36804 362218 36986 362454
rect 37222 362218 37404 362454
rect 36804 362134 37404 362218
rect 36804 361898 36986 362134
rect 37222 361898 37404 362134
rect 36804 326454 37404 361898
rect 36804 326218 36986 326454
rect 37222 326218 37404 326454
rect 36804 326134 37404 326218
rect 36804 325898 36986 326134
rect 37222 325898 37404 326134
rect 36804 290454 37404 325898
rect 36804 290218 36986 290454
rect 37222 290218 37404 290454
rect 36804 290134 37404 290218
rect 36804 289898 36986 290134
rect 37222 289898 37404 290134
rect 36804 274600 37404 289898
rect 54804 380454 55404 382916
rect 54804 380218 54986 380454
rect 55222 380218 55404 380454
rect 54804 380134 55404 380218
rect 54804 379898 54986 380134
rect 55222 379898 55404 380134
rect 54804 344454 55404 379898
rect 54804 344218 54986 344454
rect 55222 344218 55404 344454
rect 54804 344134 55404 344218
rect 54804 343898 54986 344134
rect 55222 343898 55404 344134
rect 54804 308454 55404 343898
rect 54804 308218 54986 308454
rect 55222 308218 55404 308454
rect 54804 308134 55404 308218
rect 54804 307898 54986 308134
rect 55222 307898 55404 308134
rect 54804 274600 55404 307898
rect 72804 362454 73404 382916
rect 72804 362218 72986 362454
rect 73222 362218 73404 362454
rect 72804 362134 73404 362218
rect 72804 361898 72986 362134
rect 73222 361898 73404 362134
rect 72804 326454 73404 361898
rect 72804 326218 72986 326454
rect 73222 326218 73404 326454
rect 72804 326134 73404 326218
rect 72804 325898 72986 326134
rect 73222 325898 73404 326134
rect 72804 290454 73404 325898
rect 72804 290218 72986 290454
rect 73222 290218 73404 290454
rect 72804 290134 73404 290218
rect 72804 289898 72986 290134
rect 73222 289898 73404 290134
rect 72804 274600 73404 289898
rect 90804 380454 91404 382916
rect 90804 380218 90986 380454
rect 91222 380218 91404 380454
rect 90804 380134 91404 380218
rect 90804 379898 90986 380134
rect 91222 379898 91404 380134
rect 90804 344454 91404 379898
rect 90804 344218 90986 344454
rect 91222 344218 91404 344454
rect 90804 344134 91404 344218
rect 90804 343898 90986 344134
rect 91222 343898 91404 344134
rect 90804 308454 91404 343898
rect 90804 308218 90986 308454
rect 91222 308218 91404 308454
rect 90804 308134 91404 308218
rect 90804 307898 90986 308134
rect 91222 307898 91404 308134
rect 90804 274600 91404 307898
rect 108804 362454 109404 382916
rect 108804 362218 108986 362454
rect 109222 362218 109404 362454
rect 108804 362134 109404 362218
rect 108804 361898 108986 362134
rect 109222 361898 109404 362134
rect 108804 326454 109404 361898
rect 108804 326218 108986 326454
rect 109222 326218 109404 326454
rect 108804 326134 109404 326218
rect 108804 325898 108986 326134
rect 109222 325898 109404 326134
rect 108804 290454 109404 325898
rect 108804 290218 108986 290454
rect 109222 290218 109404 290454
rect 108804 290134 109404 290218
rect 108804 289898 108986 290134
rect 109222 289898 109404 290134
rect 108804 274600 109404 289898
rect 126804 380454 127404 382916
rect 126804 380218 126986 380454
rect 127222 380218 127404 380454
rect 126804 380134 127404 380218
rect 126804 379898 126986 380134
rect 127222 379898 127404 380134
rect 126804 344454 127404 379898
rect 126804 344218 126986 344454
rect 127222 344218 127404 344454
rect 126804 344134 127404 344218
rect 126804 343898 126986 344134
rect 127222 343898 127404 344134
rect 126804 308454 127404 343898
rect 126804 308218 126986 308454
rect 127222 308218 127404 308454
rect 126804 308134 127404 308218
rect 126804 307898 126986 308134
rect 127222 307898 127404 308134
rect 126804 274600 127404 307898
rect 144804 362454 145404 382916
rect 144804 362218 144986 362454
rect 145222 362218 145404 362454
rect 144804 362134 145404 362218
rect 144804 361898 144986 362134
rect 145222 361898 145404 362134
rect 144804 326454 145404 361898
rect 144804 326218 144986 326454
rect 145222 326218 145404 326454
rect 144804 326134 145404 326218
rect 144804 325898 144986 326134
rect 145222 325898 145404 326134
rect 144804 290454 145404 325898
rect 144804 290218 144986 290454
rect 145222 290218 145404 290454
rect 144804 290134 145404 290218
rect 144804 289898 144986 290134
rect 145222 289898 145404 290134
rect 144804 274600 145404 289898
rect 162804 380454 163404 382916
rect 162804 380218 162986 380454
rect 163222 380218 163404 380454
rect 162804 380134 163404 380218
rect 162804 379898 162986 380134
rect 163222 379898 163404 380134
rect 162804 344454 163404 379898
rect 162804 344218 162986 344454
rect 163222 344218 163404 344454
rect 162804 344134 163404 344218
rect 162804 343898 162986 344134
rect 163222 343898 163404 344134
rect 162804 308454 163404 343898
rect 162804 308218 162986 308454
rect 163222 308218 163404 308454
rect 162804 308134 163404 308218
rect 162804 307898 162986 308134
rect 163222 307898 163404 308134
rect 162804 274600 163404 307898
rect 180804 362454 181404 382916
rect 180804 362218 180986 362454
rect 181222 362218 181404 362454
rect 180804 362134 181404 362218
rect 180804 361898 180986 362134
rect 181222 361898 181404 362134
rect 180804 326454 181404 361898
rect 180804 326218 180986 326454
rect 181222 326218 181404 326454
rect 180804 326134 181404 326218
rect 180804 325898 180986 326134
rect 181222 325898 181404 326134
rect 180804 290454 181404 325898
rect 180804 290218 180986 290454
rect 181222 290218 181404 290454
rect 180804 290134 181404 290218
rect 180804 289898 180986 290134
rect 181222 289898 181404 290134
rect 180804 274600 181404 289898
rect 198804 380454 199404 382916
rect 198804 380218 198986 380454
rect 199222 380218 199404 380454
rect 198804 380134 199404 380218
rect 198804 379898 198986 380134
rect 199222 379898 199404 380134
rect 198804 344454 199404 379898
rect 198804 344218 198986 344454
rect 199222 344218 199404 344454
rect 198804 344134 199404 344218
rect 198804 343898 198986 344134
rect 199222 343898 199404 344134
rect 198804 308454 199404 343898
rect 198804 308218 198986 308454
rect 199222 308218 199404 308454
rect 198804 308134 199404 308218
rect 198804 307898 198986 308134
rect 199222 307898 199404 308134
rect 198804 274600 199404 307898
rect 216804 362454 217404 382916
rect 216804 362218 216986 362454
rect 217222 362218 217404 362454
rect 216804 362134 217404 362218
rect 216804 361898 216986 362134
rect 217222 361898 217404 362134
rect 216804 326454 217404 361898
rect 216804 326218 216986 326454
rect 217222 326218 217404 326454
rect 216804 326134 217404 326218
rect 216804 325898 216986 326134
rect 217222 325898 217404 326134
rect 216804 290454 217404 325898
rect 216804 290218 216986 290454
rect 217222 290218 217404 290454
rect 216804 290134 217404 290218
rect 216804 289898 216986 290134
rect 217222 289898 217404 290134
rect 216804 274600 217404 289898
rect 234804 380454 235404 382916
rect 234804 380218 234986 380454
rect 235222 380218 235404 380454
rect 234804 380134 235404 380218
rect 234804 379898 234986 380134
rect 235222 379898 235404 380134
rect 234804 344454 235404 379898
rect 234804 344218 234986 344454
rect 235222 344218 235404 344454
rect 234804 344134 235404 344218
rect 234804 343898 234986 344134
rect 235222 343898 235404 344134
rect 234804 308454 235404 343898
rect 234804 308218 234986 308454
rect 235222 308218 235404 308454
rect 234804 308134 235404 308218
rect 234804 307898 234986 308134
rect 235222 307898 235404 308134
rect 234804 274600 235404 307898
rect 252804 362454 253404 382916
rect 252804 362218 252986 362454
rect 253222 362218 253404 362454
rect 252804 362134 253404 362218
rect 252804 361898 252986 362134
rect 253222 361898 253404 362134
rect 252804 326454 253404 361898
rect 270804 380454 271404 415898
rect 270804 380218 270986 380454
rect 271222 380218 271404 380454
rect 270804 380134 271404 380218
rect 270804 379898 270986 380134
rect 271222 379898 271404 380134
rect 270804 356560 271404 379898
rect 274403 354924 274469 354925
rect 274403 354860 274404 354924
rect 274468 354860 274469 354924
rect 274403 354859 274469 354860
rect 252804 326218 252986 326454
rect 253222 326218 253404 326454
rect 252804 326134 253404 326218
rect 252804 325898 252986 326134
rect 253222 325898 253404 326134
rect 252804 290454 253404 325898
rect 252804 290218 252986 290454
rect 253222 290218 253404 290454
rect 252804 290134 253404 290218
rect 252804 289898 252986 290134
rect 253222 289898 253404 290134
rect 252804 274600 253404 289898
rect 270804 308454 271404 314560
rect 270804 308218 270986 308454
rect 271222 308218 271404 308454
rect 270804 308134 271404 308218
rect 270804 307898 270986 308134
rect 271222 307898 271404 308134
rect 18804 272218 18986 272454
rect 19222 272218 19404 272454
rect 18804 272134 19404 272218
rect 18804 271898 18986 272134
rect 19222 271898 19404 272134
rect 18804 236454 19404 271898
rect 270804 272454 271404 307898
rect 270804 272218 270986 272454
rect 271222 272218 271404 272454
rect 270804 272134 271404 272218
rect 270804 271898 270986 272134
rect 271222 271898 271404 272134
rect 262128 254454 262448 254476
rect 262128 254218 262170 254454
rect 262406 254218 262448 254454
rect 262128 254134 262448 254218
rect 262128 253898 262170 254134
rect 262406 253898 262448 254134
rect 262128 253876 262448 253898
rect 18804 236218 18986 236454
rect 19222 236218 19404 236454
rect 18804 236134 19404 236218
rect 18804 235898 18986 236134
rect 19222 235898 19404 236134
rect 18804 200454 19404 235898
rect 246768 236454 247088 236476
rect 246768 236218 246810 236454
rect 247046 236218 247088 236454
rect 246768 236134 247088 236218
rect 246768 235898 246810 236134
rect 247046 235898 247088 236134
rect 246768 235876 247088 235898
rect 270804 236454 271404 271898
rect 270804 236218 270986 236454
rect 271222 236218 271404 236454
rect 270804 236134 271404 236218
rect 270804 235898 270986 236134
rect 271222 235898 271404 236134
rect 262128 218454 262448 218476
rect 262128 218218 262170 218454
rect 262406 218218 262448 218454
rect 262128 218134 262448 218218
rect 262128 217898 262170 218134
rect 262406 217898 262448 218134
rect 262128 217876 262448 217898
rect 18804 200218 18986 200454
rect 19222 200218 19404 200454
rect 18804 200134 19404 200218
rect 18804 199898 18986 200134
rect 19222 199898 19404 200134
rect 18804 164454 19404 199898
rect 246768 200454 247088 200476
rect 246768 200218 246810 200454
rect 247046 200218 247088 200454
rect 246768 200134 247088 200218
rect 246768 199898 246810 200134
rect 247046 199898 247088 200134
rect 246768 199876 247088 199898
rect 270804 200454 271404 235898
rect 270804 200218 270986 200454
rect 271222 200218 271404 200454
rect 270804 200134 271404 200218
rect 270804 199898 270986 200134
rect 271222 199898 271404 200134
rect 262128 182454 262448 182476
rect 262128 182218 262170 182454
rect 262406 182218 262448 182454
rect 262128 182134 262448 182218
rect 262128 181898 262170 182134
rect 262406 181898 262448 182134
rect 262128 181876 262448 181898
rect 18804 164218 18986 164454
rect 19222 164218 19404 164454
rect 18804 164134 19404 164218
rect 18804 163898 18986 164134
rect 19222 163898 19404 164134
rect 18804 128454 19404 163898
rect 246768 164454 247088 164476
rect 246768 164218 246810 164454
rect 247046 164218 247088 164454
rect 246768 164134 247088 164218
rect 246768 163898 246810 164134
rect 247046 163898 247088 164134
rect 246768 163876 247088 163898
rect 270804 164454 271404 199898
rect 270804 164218 270986 164454
rect 271222 164218 271404 164454
rect 270804 164134 271404 164218
rect 270804 163898 270986 164134
rect 271222 163898 271404 164134
rect 262128 146454 262448 146476
rect 262128 146218 262170 146454
rect 262406 146218 262448 146454
rect 262128 146134 262448 146218
rect 262128 145898 262170 146134
rect 262406 145898 262448 146134
rect 262128 145876 262448 145898
rect 18804 128218 18986 128454
rect 19222 128218 19404 128454
rect 18804 128134 19404 128218
rect 18804 127898 18986 128134
rect 19222 127898 19404 128134
rect 18804 92454 19404 127898
rect 246768 128454 247088 128476
rect 246768 128218 246810 128454
rect 247046 128218 247088 128454
rect 246768 128134 247088 128218
rect 246768 127898 246810 128134
rect 247046 127898 247088 128134
rect 246768 127876 247088 127898
rect 270804 128454 271404 163898
rect 270804 128218 270986 128454
rect 271222 128218 271404 128454
rect 270804 128134 271404 128218
rect 270804 127898 270986 128134
rect 271222 127898 271404 128134
rect 262128 110454 262448 110476
rect 262128 110218 262170 110454
rect 262406 110218 262448 110454
rect 262128 110134 262448 110218
rect 262128 109898 262170 110134
rect 262406 109898 262448 110134
rect 262128 109876 262448 109898
rect 18804 92218 18986 92454
rect 19222 92218 19404 92454
rect 18804 92134 19404 92218
rect 18804 91898 18986 92134
rect 19222 91898 19404 92134
rect 18804 56454 19404 91898
rect 246768 92454 247088 92476
rect 246768 92218 246810 92454
rect 247046 92218 247088 92454
rect 246768 92134 247088 92218
rect 246768 91898 246810 92134
rect 247046 91898 247088 92134
rect 246768 91876 247088 91898
rect 270804 92454 271404 127898
rect 270804 92218 270986 92454
rect 271222 92218 271404 92454
rect 270804 92134 271404 92218
rect 270804 91898 270986 92134
rect 271222 91898 271404 92134
rect 18804 56218 18986 56454
rect 19222 56218 19404 56454
rect 18804 56134 19404 56218
rect 18804 55898 18986 56134
rect 19222 55898 19404 56134
rect 18804 20454 19404 55898
rect 18804 20218 18986 20454
rect 19222 20218 19404 20454
rect 18804 20134 19404 20218
rect 18804 19898 18986 20134
rect 19222 19898 19404 20134
rect 18804 -1286 19404 19898
rect 18804 -1522 18986 -1286
rect 19222 -1522 19404 -1286
rect 18804 -1606 19404 -1522
rect 18804 -1842 18986 -1606
rect 19222 -1842 19404 -1606
rect 18804 -1864 19404 -1842
rect 36804 38454 37404 72600
rect 36804 38218 36986 38454
rect 37222 38218 37404 38454
rect 36804 38134 37404 38218
rect 36804 37898 36986 38134
rect 37222 37898 37404 38134
rect 36804 2454 37404 37898
rect 36804 2218 36986 2454
rect 37222 2218 37404 2454
rect 36804 2134 37404 2218
rect 36804 1898 36986 2134
rect 37222 1898 37404 2134
rect 36804 -346 37404 1898
rect 36804 -582 36986 -346
rect 37222 -582 37404 -346
rect 36804 -666 37404 -582
rect 36804 -902 36986 -666
rect 37222 -902 37404 -666
rect 36804 -1864 37404 -902
rect 54804 56454 55404 72600
rect 54804 56218 54986 56454
rect 55222 56218 55404 56454
rect 54804 56134 55404 56218
rect 54804 55898 54986 56134
rect 55222 55898 55404 56134
rect 54804 20454 55404 55898
rect 54804 20218 54986 20454
rect 55222 20218 55404 20454
rect 54804 20134 55404 20218
rect 54804 19898 54986 20134
rect 55222 19898 55404 20134
rect 54804 -1286 55404 19898
rect 54804 -1522 54986 -1286
rect 55222 -1522 55404 -1286
rect 54804 -1606 55404 -1522
rect 54804 -1842 54986 -1606
rect 55222 -1842 55404 -1606
rect 54804 -1864 55404 -1842
rect 72804 38454 73404 72600
rect 72804 38218 72986 38454
rect 73222 38218 73404 38454
rect 72804 38134 73404 38218
rect 72804 37898 72986 38134
rect 73222 37898 73404 38134
rect 72804 2454 73404 37898
rect 72804 2218 72986 2454
rect 73222 2218 73404 2454
rect 72804 2134 73404 2218
rect 72804 1898 72986 2134
rect 73222 1898 73404 2134
rect 72804 -346 73404 1898
rect 72804 -582 72986 -346
rect 73222 -582 73404 -346
rect 72804 -666 73404 -582
rect 72804 -902 72986 -666
rect 73222 -902 73404 -666
rect 72804 -1864 73404 -902
rect 90804 56454 91404 72600
rect 90804 56218 90986 56454
rect 91222 56218 91404 56454
rect 90804 56134 91404 56218
rect 90804 55898 90986 56134
rect 91222 55898 91404 56134
rect 90804 20454 91404 55898
rect 90804 20218 90986 20454
rect 91222 20218 91404 20454
rect 90804 20134 91404 20218
rect 90804 19898 90986 20134
rect 91222 19898 91404 20134
rect 90804 -1286 91404 19898
rect 90804 -1522 90986 -1286
rect 91222 -1522 91404 -1286
rect 90804 -1606 91404 -1522
rect 90804 -1842 90986 -1606
rect 91222 -1842 91404 -1606
rect 90804 -1864 91404 -1842
rect 108804 38454 109404 72600
rect 108804 38218 108986 38454
rect 109222 38218 109404 38454
rect 108804 38134 109404 38218
rect 108804 37898 108986 38134
rect 109222 37898 109404 38134
rect 108804 2454 109404 37898
rect 108804 2218 108986 2454
rect 109222 2218 109404 2454
rect 108804 2134 109404 2218
rect 108804 1898 108986 2134
rect 109222 1898 109404 2134
rect 108804 -346 109404 1898
rect 108804 -582 108986 -346
rect 109222 -582 109404 -346
rect 108804 -666 109404 -582
rect 108804 -902 108986 -666
rect 109222 -902 109404 -666
rect 108804 -1864 109404 -902
rect 126804 56454 127404 72600
rect 126804 56218 126986 56454
rect 127222 56218 127404 56454
rect 126804 56134 127404 56218
rect 126804 55898 126986 56134
rect 127222 55898 127404 56134
rect 126804 20454 127404 55898
rect 126804 20218 126986 20454
rect 127222 20218 127404 20454
rect 126804 20134 127404 20218
rect 126804 19898 126986 20134
rect 127222 19898 127404 20134
rect 126804 -1286 127404 19898
rect 126804 -1522 126986 -1286
rect 127222 -1522 127404 -1286
rect 126804 -1606 127404 -1522
rect 126804 -1842 126986 -1606
rect 127222 -1842 127404 -1606
rect 126804 -1864 127404 -1842
rect 144804 38454 145404 72600
rect 144804 38218 144986 38454
rect 145222 38218 145404 38454
rect 144804 38134 145404 38218
rect 144804 37898 144986 38134
rect 145222 37898 145404 38134
rect 144804 2454 145404 37898
rect 144804 2218 144986 2454
rect 145222 2218 145404 2454
rect 144804 2134 145404 2218
rect 144804 1898 144986 2134
rect 145222 1898 145404 2134
rect 144804 -346 145404 1898
rect 144804 -582 144986 -346
rect 145222 -582 145404 -346
rect 144804 -666 145404 -582
rect 144804 -902 144986 -666
rect 145222 -902 145404 -666
rect 144804 -1864 145404 -902
rect 162804 56454 163404 72600
rect 162804 56218 162986 56454
rect 163222 56218 163404 56454
rect 162804 56134 163404 56218
rect 162804 55898 162986 56134
rect 163222 55898 163404 56134
rect 162804 20454 163404 55898
rect 162804 20218 162986 20454
rect 163222 20218 163404 20454
rect 162804 20134 163404 20218
rect 162804 19898 162986 20134
rect 163222 19898 163404 20134
rect 162804 -1286 163404 19898
rect 162804 -1522 162986 -1286
rect 163222 -1522 163404 -1286
rect 162804 -1606 163404 -1522
rect 162804 -1842 162986 -1606
rect 163222 -1842 163404 -1606
rect 162804 -1864 163404 -1842
rect 180804 38454 181404 72600
rect 180804 38218 180986 38454
rect 181222 38218 181404 38454
rect 180804 38134 181404 38218
rect 180804 37898 180986 38134
rect 181222 37898 181404 38134
rect 180804 2454 181404 37898
rect 180804 2218 180986 2454
rect 181222 2218 181404 2454
rect 180804 2134 181404 2218
rect 180804 1898 180986 2134
rect 181222 1898 181404 2134
rect 180804 -346 181404 1898
rect 180804 -582 180986 -346
rect 181222 -582 181404 -346
rect 180804 -666 181404 -582
rect 180804 -902 180986 -666
rect 181222 -902 181404 -666
rect 180804 -1864 181404 -902
rect 198804 56454 199404 72600
rect 198804 56218 198986 56454
rect 199222 56218 199404 56454
rect 198804 56134 199404 56218
rect 198804 55898 198986 56134
rect 199222 55898 199404 56134
rect 198804 20454 199404 55898
rect 198804 20218 198986 20454
rect 199222 20218 199404 20454
rect 198804 20134 199404 20218
rect 198804 19898 198986 20134
rect 199222 19898 199404 20134
rect 198804 -1286 199404 19898
rect 198804 -1522 198986 -1286
rect 199222 -1522 199404 -1286
rect 198804 -1606 199404 -1522
rect 198804 -1842 198986 -1606
rect 199222 -1842 199404 -1606
rect 198804 -1864 199404 -1842
rect 216804 38454 217404 72600
rect 216804 38218 216986 38454
rect 217222 38218 217404 38454
rect 216804 38134 217404 38218
rect 216804 37898 216986 38134
rect 217222 37898 217404 38134
rect 216804 2454 217404 37898
rect 216804 2218 216986 2454
rect 217222 2218 217404 2454
rect 216804 2134 217404 2218
rect 216804 1898 216986 2134
rect 217222 1898 217404 2134
rect 216804 -346 217404 1898
rect 216804 -582 216986 -346
rect 217222 -582 217404 -346
rect 216804 -666 217404 -582
rect 216804 -902 216986 -666
rect 217222 -902 217404 -666
rect 216804 -1864 217404 -902
rect 234804 56454 235404 72600
rect 234804 56218 234986 56454
rect 235222 56218 235404 56454
rect 234804 56134 235404 56218
rect 234804 55898 234986 56134
rect 235222 55898 235404 56134
rect 234804 20454 235404 55898
rect 234804 20218 234986 20454
rect 235222 20218 235404 20454
rect 234804 20134 235404 20218
rect 234804 19898 234986 20134
rect 235222 19898 235404 20134
rect 234804 -1286 235404 19898
rect 234804 -1522 234986 -1286
rect 235222 -1522 235404 -1286
rect 234804 -1606 235404 -1522
rect 234804 -1842 234986 -1606
rect 235222 -1842 235404 -1606
rect 234804 -1864 235404 -1842
rect 252804 38454 253404 72600
rect 252804 38218 252986 38454
rect 253222 38218 253404 38454
rect 252804 38134 253404 38218
rect 252804 37898 252986 38134
rect 253222 37898 253404 38134
rect 252804 2454 253404 37898
rect 252804 2218 252986 2454
rect 253222 2218 253404 2454
rect 252804 2134 253404 2218
rect 252804 1898 252986 2134
rect 253222 1898 253404 2134
rect 252804 -346 253404 1898
rect 252804 -582 252986 -346
rect 253222 -582 253404 -346
rect 252804 -666 253404 -582
rect 252804 -902 252986 -666
rect 253222 -902 253404 -666
rect 252804 -1864 253404 -902
rect 270804 56454 271404 91898
rect 274406 72045 274466 354859
rect 275142 316301 275202 699891
rect 288804 686454 289404 704282
rect 306804 705778 307404 705800
rect 306804 705542 306986 705778
rect 307222 705542 307404 705778
rect 306804 705458 307404 705542
rect 306804 705222 306986 705458
rect 307222 705222 307404 705458
rect 299059 700636 299125 700637
rect 299059 700572 299060 700636
rect 299124 700572 299125 700636
rect 299059 700571 299125 700572
rect 288804 686218 288986 686454
rect 289222 686218 289404 686454
rect 288804 686134 289404 686218
rect 288804 685898 288986 686134
rect 289222 685898 289404 686134
rect 288804 650454 289404 685898
rect 288804 650218 288986 650454
rect 289222 650218 289404 650454
rect 288804 650134 289404 650218
rect 288804 649898 288986 650134
rect 289222 649898 289404 650134
rect 288804 614454 289404 649898
rect 288804 614218 288986 614454
rect 289222 614218 289404 614454
rect 288804 614134 289404 614218
rect 288804 613898 288986 614134
rect 289222 613898 289404 614134
rect 288804 578454 289404 613898
rect 295747 586260 295813 586261
rect 295747 586196 295748 586260
rect 295812 586196 295813 586260
rect 295747 586195 295813 586196
rect 292803 586124 292869 586125
rect 292803 586060 292804 586124
rect 292868 586060 292869 586124
rect 292803 586059 292869 586060
rect 288804 578218 288986 578454
rect 289222 578218 289404 578454
rect 288804 578134 289404 578218
rect 288804 577898 288986 578134
rect 289222 577898 289404 578134
rect 288804 542454 289404 577898
rect 288804 542218 288986 542454
rect 289222 542218 289404 542454
rect 288804 542134 289404 542218
rect 288804 541898 288986 542134
rect 289222 541898 289404 542134
rect 288804 506454 289404 541898
rect 288804 506218 288986 506454
rect 289222 506218 289404 506454
rect 288804 506134 289404 506218
rect 288804 505898 288986 506134
rect 289222 505898 289404 506134
rect 288804 470454 289404 505898
rect 288804 470218 288986 470454
rect 289222 470218 289404 470454
rect 288804 470134 289404 470218
rect 288804 469898 288986 470134
rect 289222 469898 289404 470134
rect 288804 434454 289404 469898
rect 288804 434218 288986 434454
rect 289222 434218 289404 434454
rect 288804 434134 289404 434218
rect 288804 433898 288986 434134
rect 289222 433898 289404 434134
rect 288804 398454 289404 433898
rect 288804 398218 288986 398454
rect 289222 398218 289404 398454
rect 288804 398134 289404 398218
rect 288804 397898 288986 398134
rect 289222 397898 289404 398134
rect 276243 382124 276309 382125
rect 276243 382060 276244 382124
rect 276308 382060 276309 382124
rect 276243 382059 276309 382060
rect 275875 354924 275941 354925
rect 275875 354860 275876 354924
rect 275940 354860 275941 354924
rect 275875 354859 275941 354860
rect 275139 316300 275205 316301
rect 275139 316236 275140 316300
rect 275204 316236 275205 316300
rect 275139 316235 275205 316236
rect 275878 276725 275938 354859
rect 276246 315621 276306 382059
rect 288804 362454 289404 397898
rect 288804 362218 288986 362454
rect 289222 362218 289404 362454
rect 288804 362134 289404 362218
rect 288804 361898 288986 362134
rect 289222 361898 289404 362134
rect 276427 359412 276493 359413
rect 276427 359348 276428 359412
rect 276492 359348 276493 359412
rect 276427 359347 276493 359348
rect 276243 315620 276309 315621
rect 276243 315556 276244 315620
rect 276308 315556 276309 315620
rect 276243 315555 276309 315556
rect 275875 276724 275941 276725
rect 275875 276660 275876 276724
rect 275940 276660 275941 276724
rect 275875 276659 275941 276660
rect 276430 272237 276490 359347
rect 276611 359276 276677 359277
rect 276611 359212 276612 359276
rect 276676 359212 276677 359276
rect 276611 359211 276677 359212
rect 276427 272236 276493 272237
rect 276427 272172 276428 272236
rect 276492 272172 276493 272236
rect 276427 272171 276493 272172
rect 276614 272101 276674 359211
rect 288804 356560 289404 361898
rect 292806 353701 292866 586059
rect 293539 546820 293605 546821
rect 293539 546756 293540 546820
rect 293604 546756 293605 546820
rect 293539 546755 293605 546756
rect 292803 353700 292869 353701
rect 292803 353636 292804 353700
rect 292868 353636 292869 353700
rect 292803 353635 292869 353636
rect 292112 344454 292432 344476
rect 292112 344218 292154 344454
rect 292390 344218 292432 344454
rect 292112 344134 292432 344218
rect 292112 343898 292154 344134
rect 292390 343898 292432 344134
rect 292112 343876 292432 343898
rect 293542 315757 293602 546755
rect 293723 384300 293789 384301
rect 293723 384236 293724 384300
rect 293788 384236 293789 384300
rect 293723 384235 293789 384236
rect 293539 315756 293605 315757
rect 293539 315692 293540 315756
rect 293604 315692 293605 315756
rect 293539 315691 293605 315692
rect 288804 290454 289404 314560
rect 293726 312085 293786 384235
rect 295011 382260 295077 382261
rect 295011 382196 295012 382260
rect 295076 382196 295077 382260
rect 295011 382195 295077 382196
rect 294275 353700 294341 353701
rect 294275 353636 294276 353700
rect 294340 353636 294341 353700
rect 294275 353635 294341 353636
rect 294278 316301 294338 353635
rect 294275 316300 294341 316301
rect 294275 316236 294276 316300
rect 294340 316236 294341 316300
rect 294275 316235 294341 316236
rect 295014 313445 295074 382195
rect 295750 316301 295810 586195
rect 295931 354924 295997 354925
rect 295931 354860 295932 354924
rect 295996 354860 295997 354924
rect 295931 354859 295997 354860
rect 298691 354924 298757 354925
rect 298691 354860 298692 354924
rect 298756 354860 298757 354924
rect 298691 354859 298757 354860
rect 295747 316300 295813 316301
rect 295747 316236 295748 316300
rect 295812 316236 295813 316300
rect 295747 316235 295813 316236
rect 295011 313444 295077 313445
rect 295011 313380 295012 313444
rect 295076 313380 295077 313444
rect 295011 313379 295077 313380
rect 293723 312084 293789 312085
rect 293723 312020 293724 312084
rect 293788 312020 293789 312084
rect 293723 312019 293789 312020
rect 288804 290218 288986 290454
rect 289222 290218 289404 290454
rect 288804 290134 289404 290218
rect 288804 289898 288986 290134
rect 289222 289898 289404 290134
rect 276611 272100 276677 272101
rect 276611 272036 276612 272100
rect 276676 272036 276677 272100
rect 276611 272035 276677 272036
rect 288804 254454 289404 289898
rect 295934 275365 295994 354859
rect 295931 275364 295997 275365
rect 295931 275300 295932 275364
rect 295996 275300 295997 275364
rect 295931 275299 295997 275300
rect 288804 254218 288986 254454
rect 289222 254218 289404 254454
rect 288804 254134 289404 254218
rect 288804 253898 288986 254134
rect 289222 253898 289404 254134
rect 288804 218454 289404 253898
rect 288804 218218 288986 218454
rect 289222 218218 289404 218454
rect 288804 218134 289404 218218
rect 288804 217898 288986 218134
rect 289222 217898 289404 218134
rect 288804 182454 289404 217898
rect 288804 182218 288986 182454
rect 289222 182218 289404 182454
rect 288804 182134 289404 182218
rect 288804 181898 288986 182134
rect 289222 181898 289404 182134
rect 288804 146454 289404 181898
rect 288804 146218 288986 146454
rect 289222 146218 289404 146454
rect 288804 146134 289404 146218
rect 288804 145898 288986 146134
rect 289222 145898 289404 146134
rect 288804 110454 289404 145898
rect 288804 110218 288986 110454
rect 289222 110218 289404 110454
rect 288804 110134 289404 110218
rect 288804 109898 288986 110134
rect 289222 109898 289404 110134
rect 288804 74454 289404 109898
rect 288804 74218 288986 74454
rect 289222 74218 289404 74454
rect 288804 74134 289404 74218
rect 288804 73898 288986 74134
rect 289222 73898 289404 74134
rect 274403 72044 274469 72045
rect 274403 71980 274404 72044
rect 274468 71980 274469 72044
rect 274403 71979 274469 71980
rect 270804 56218 270986 56454
rect 271222 56218 271404 56454
rect 270804 56134 271404 56218
rect 270804 55898 270986 56134
rect 271222 55898 271404 56134
rect 270804 20454 271404 55898
rect 270804 20218 270986 20454
rect 271222 20218 271404 20454
rect 270804 20134 271404 20218
rect 270804 19898 270986 20134
rect 271222 19898 271404 20134
rect 270804 -1286 271404 19898
rect 270804 -1522 270986 -1286
rect 271222 -1522 271404 -1286
rect 270804 -1606 271404 -1522
rect 270804 -1842 270986 -1606
rect 271222 -1842 271404 -1606
rect 270804 -1864 271404 -1842
rect 288804 38454 289404 73898
rect 288804 38218 288986 38454
rect 289222 38218 289404 38454
rect 288804 38134 289404 38218
rect 288804 37898 288986 38134
rect 289222 37898 289404 38134
rect 288804 2454 289404 37898
rect 298694 3637 298754 354859
rect 299062 313173 299122 700571
rect 306804 668454 307404 705222
rect 306804 668218 306986 668454
rect 307222 668218 307404 668454
rect 306804 668134 307404 668218
rect 306804 667898 306986 668134
rect 307222 667898 307404 668134
rect 306804 632454 307404 667898
rect 306804 632218 306986 632454
rect 307222 632218 307404 632454
rect 306804 632134 307404 632218
rect 306804 631898 306986 632134
rect 307222 631898 307404 632134
rect 306804 596454 307404 631898
rect 324804 704838 325404 705800
rect 324804 704602 324986 704838
rect 325222 704602 325404 704838
rect 324804 704518 325404 704602
rect 324804 704282 324986 704518
rect 325222 704282 325404 704518
rect 324804 686454 325404 704282
rect 324804 686218 324986 686454
rect 325222 686218 325404 686454
rect 324804 686134 325404 686218
rect 324804 685898 324986 686134
rect 325222 685898 325404 686134
rect 324804 650454 325404 685898
rect 324804 650218 324986 650454
rect 325222 650218 325404 650454
rect 324804 650134 325404 650218
rect 324804 649898 324986 650134
rect 325222 649898 325404 650134
rect 324804 614454 325404 649898
rect 324804 614218 324986 614454
rect 325222 614218 325404 614454
rect 324804 614134 325404 614218
rect 324804 613898 324986 614134
rect 325222 613898 325404 614134
rect 310651 609516 310717 609517
rect 310651 609452 310652 609516
rect 310716 609452 310717 609516
rect 310651 609451 310717 609452
rect 306804 596218 306986 596454
rect 307222 596218 307404 596454
rect 306804 596134 307404 596218
rect 306804 595898 306986 596134
rect 307222 595898 307404 596134
rect 306603 585988 306669 585989
rect 306603 585924 306604 585988
rect 306668 585924 306669 585988
rect 306603 585923 306669 585924
rect 300163 381308 300229 381309
rect 300163 381244 300164 381308
rect 300228 381244 300229 381308
rect 300163 381243 300229 381244
rect 299427 354924 299493 354925
rect 299427 354860 299428 354924
rect 299492 354860 299493 354924
rect 299427 354859 299493 354860
rect 299059 313172 299125 313173
rect 299059 313108 299060 313172
rect 299124 313108 299125 313172
rect 299059 313107 299125 313108
rect 299430 92717 299490 354859
rect 300166 316301 300226 381243
rect 306419 355332 306485 355333
rect 306419 355268 306420 355332
rect 306484 355268 306485 355332
rect 306419 355267 306485 355268
rect 300163 316300 300229 316301
rect 300163 316236 300164 316300
rect 300228 316236 300229 316300
rect 300163 316235 300229 316236
rect 306422 276725 306482 355267
rect 306606 315621 306666 585923
rect 306804 560454 307404 595898
rect 310467 566676 310533 566677
rect 310467 566612 310468 566676
rect 310532 566612 310533 566676
rect 310467 566611 310533 566612
rect 306804 560218 306986 560454
rect 307222 560218 307404 560454
rect 306804 560134 307404 560218
rect 306804 559898 306986 560134
rect 307222 559898 307404 560134
rect 306804 524454 307404 559898
rect 306804 524218 306986 524454
rect 307222 524218 307404 524454
rect 306804 524134 307404 524218
rect 306804 523898 306986 524134
rect 307222 523898 307404 524134
rect 306804 488454 307404 523898
rect 310470 511597 310530 566611
rect 310467 511596 310533 511597
rect 310467 511532 310468 511596
rect 310532 511532 310533 511596
rect 310467 511531 310533 511532
rect 309363 504932 309429 504933
rect 309363 504868 309364 504932
rect 309428 504868 309429 504932
rect 309363 504867 309429 504868
rect 309366 497725 309426 504867
rect 309363 497724 309429 497725
rect 309363 497660 309364 497724
rect 309428 497660 309429 497724
rect 309363 497659 309429 497660
rect 309547 497452 309613 497453
rect 309547 497388 309548 497452
rect 309612 497388 309613 497452
rect 309547 497387 309613 497388
rect 306804 488218 306986 488454
rect 307222 488218 307404 488454
rect 306804 488134 307404 488218
rect 306804 487898 306986 488134
rect 307222 487898 307404 488134
rect 306804 452454 307404 487898
rect 309550 487250 309610 497387
rect 309550 487190 309794 487250
rect 309734 484261 309794 487190
rect 309731 484260 309797 484261
rect 309731 484196 309732 484260
rect 309796 484196 309797 484260
rect 309731 484195 309797 484196
rect 309915 484124 309981 484125
rect 309915 484060 309916 484124
rect 309980 484060 309981 484124
rect 309915 484059 309981 484060
rect 309918 473925 309978 484059
rect 309915 473924 309981 473925
rect 309915 473860 309916 473924
rect 309980 473860 309981 473924
rect 309915 473859 309981 473860
rect 310099 463724 310165 463725
rect 310099 463660 310100 463724
rect 310164 463660 310165 463724
rect 310099 463659 310165 463660
rect 310102 458557 310162 463659
rect 309547 458556 309613 458557
rect 309547 458492 309548 458556
rect 309612 458492 309613 458556
rect 309547 458491 309613 458492
rect 310099 458556 310165 458557
rect 310099 458492 310100 458556
rect 310164 458492 310165 458556
rect 310099 458491 310165 458492
rect 306804 452218 306986 452454
rect 307222 452218 307404 452454
rect 306804 452134 307404 452218
rect 306804 451898 306986 452134
rect 307222 451898 307404 452134
rect 306804 416454 307404 451898
rect 309550 446045 309610 458491
rect 309547 446044 309613 446045
rect 309547 445980 309548 446044
rect 309612 445980 309613 446044
rect 309547 445979 309613 445980
rect 310099 446044 310165 446045
rect 310099 445980 310100 446044
rect 310164 445980 310165 446044
rect 310099 445979 310165 445980
rect 310102 435845 310162 445979
rect 310099 435844 310165 435845
rect 310099 435780 310100 435844
rect 310164 435780 310165 435844
rect 310099 435779 310165 435780
rect 310099 435708 310165 435709
rect 310099 435644 310100 435708
rect 310164 435644 310165 435708
rect 310099 435643 310165 435644
rect 310102 432850 310162 435643
rect 309918 432790 310162 432850
rect 309918 432581 309978 432790
rect 309915 432580 309981 432581
rect 309915 432516 309916 432580
rect 309980 432516 309981 432580
rect 309915 432515 309981 432516
rect 309731 422516 309797 422517
rect 309731 422452 309732 422516
rect 309796 422452 309797 422516
rect 309731 422451 309797 422452
rect 306804 416218 306986 416454
rect 307222 416218 307404 416454
rect 306804 416134 307404 416218
rect 306804 415898 306986 416134
rect 307222 415898 307404 416134
rect 306804 380454 307404 415898
rect 309734 415309 309794 422451
rect 309731 415308 309797 415309
rect 309731 415244 309732 415308
rect 309796 415244 309797 415308
rect 309731 415243 309797 415244
rect 309915 415036 309981 415037
rect 309915 414972 309916 415036
rect 309980 414972 309981 415036
rect 309915 414971 309981 414972
rect 309918 412181 309978 414971
rect 309915 412180 309981 412181
rect 309915 412116 309916 412180
rect 309980 412116 309981 412180
rect 309915 412115 309981 412116
rect 309731 401980 309797 401981
rect 309731 401916 309732 401980
rect 309796 401916 309797 401980
rect 309731 401915 309797 401916
rect 309734 394637 309794 401915
rect 309731 394636 309797 394637
rect 309731 394572 309732 394636
rect 309796 394572 309797 394636
rect 309731 394571 309797 394572
rect 309915 394364 309981 394365
rect 309915 394300 309916 394364
rect 309980 394300 309981 394364
rect 309915 394299 309981 394300
rect 309918 391509 309978 394299
rect 309915 391508 309981 391509
rect 309915 391444 309916 391508
rect 309980 391444 309981 391508
rect 309915 391443 309981 391444
rect 309731 381308 309797 381309
rect 309731 381244 309732 381308
rect 309796 381244 309797 381308
rect 309731 381243 309797 381244
rect 306804 380218 306986 380454
rect 307222 380218 307404 380454
rect 306804 380134 307404 380218
rect 306804 379898 306986 380134
rect 307222 379898 307404 380134
rect 306804 356560 307404 379898
rect 309734 374101 309794 381243
rect 309731 374100 309797 374101
rect 309731 374036 309732 374100
rect 309796 374036 309797 374100
rect 309731 374035 309797 374036
rect 309547 373828 309613 373829
rect 309547 373764 309548 373828
rect 309612 373764 309613 373828
rect 309547 373763 309613 373764
rect 309550 370973 309610 373763
rect 309547 370972 309613 370973
rect 309547 370908 309548 370972
rect 309612 370908 309613 370972
rect 309547 370907 309613 370908
rect 309363 360772 309429 360773
rect 309363 360708 309364 360772
rect 309428 360708 309429 360772
rect 309363 360707 309429 360708
rect 309366 355330 309426 360707
rect 309366 355270 309610 355330
rect 309550 342410 309610 355270
rect 309550 342350 309794 342410
rect 309734 332890 309794 342350
rect 310654 334250 310714 609451
rect 324804 584916 325404 613898
rect 342804 705778 343404 705800
rect 342804 705542 342986 705778
rect 343222 705542 343404 705778
rect 342804 705458 343404 705542
rect 342804 705222 342986 705458
rect 343222 705222 343404 705458
rect 342804 668454 343404 705222
rect 342804 668218 342986 668454
rect 343222 668218 343404 668454
rect 342804 668134 343404 668218
rect 342804 667898 342986 668134
rect 343222 667898 343404 668134
rect 342804 632454 343404 667898
rect 342804 632218 342986 632454
rect 343222 632218 343404 632454
rect 342804 632134 343404 632218
rect 342804 631898 342986 632134
rect 343222 631898 343404 632134
rect 342804 596454 343404 631898
rect 342804 596218 342986 596454
rect 343222 596218 343404 596454
rect 342804 596134 343404 596218
rect 342804 595898 342986 596134
rect 343222 595898 343404 596134
rect 342804 584916 343404 595898
rect 360804 704838 361404 705800
rect 360804 704602 360986 704838
rect 361222 704602 361404 704838
rect 360804 704518 361404 704602
rect 360804 704282 360986 704518
rect 361222 704282 361404 704518
rect 360804 686454 361404 704282
rect 360804 686218 360986 686454
rect 361222 686218 361404 686454
rect 360804 686134 361404 686218
rect 360804 685898 360986 686134
rect 361222 685898 361404 686134
rect 360804 650454 361404 685898
rect 360804 650218 360986 650454
rect 361222 650218 361404 650454
rect 360804 650134 361404 650218
rect 360804 649898 360986 650134
rect 361222 649898 361404 650134
rect 360804 614454 361404 649898
rect 360804 614218 360986 614454
rect 361222 614218 361404 614454
rect 360804 614134 361404 614218
rect 360804 613898 360986 614134
rect 361222 613898 361404 614134
rect 360804 584916 361404 613898
rect 378804 705778 379404 705800
rect 378804 705542 378986 705778
rect 379222 705542 379404 705778
rect 378804 705458 379404 705542
rect 378804 705222 378986 705458
rect 379222 705222 379404 705458
rect 378804 668454 379404 705222
rect 378804 668218 378986 668454
rect 379222 668218 379404 668454
rect 378804 668134 379404 668218
rect 378804 667898 378986 668134
rect 379222 667898 379404 668134
rect 378804 632454 379404 667898
rect 378804 632218 378986 632454
rect 379222 632218 379404 632454
rect 378804 632134 379404 632218
rect 378804 631898 378986 632134
rect 379222 631898 379404 632134
rect 378804 596454 379404 631898
rect 378804 596218 378986 596454
rect 379222 596218 379404 596454
rect 378804 596134 379404 596218
rect 378804 595898 378986 596134
rect 379222 595898 379404 596134
rect 378804 584916 379404 595898
rect 396804 704838 397404 705800
rect 396804 704602 396986 704838
rect 397222 704602 397404 704838
rect 396804 704518 397404 704602
rect 396804 704282 396986 704518
rect 397222 704282 397404 704518
rect 396804 686454 397404 704282
rect 396804 686218 396986 686454
rect 397222 686218 397404 686454
rect 396804 686134 397404 686218
rect 396804 685898 396986 686134
rect 397222 685898 397404 686134
rect 396804 650454 397404 685898
rect 396804 650218 396986 650454
rect 397222 650218 397404 650454
rect 396804 650134 397404 650218
rect 396804 649898 396986 650134
rect 397222 649898 397404 650134
rect 396804 614454 397404 649898
rect 396804 614218 396986 614454
rect 397222 614218 397404 614454
rect 396804 614134 397404 614218
rect 396804 613898 396986 614134
rect 397222 613898 397404 614134
rect 396804 584916 397404 613898
rect 414804 705778 415404 705800
rect 414804 705542 414986 705778
rect 415222 705542 415404 705778
rect 414804 705458 415404 705542
rect 414804 705222 414986 705458
rect 415222 705222 415404 705458
rect 414804 668454 415404 705222
rect 414804 668218 414986 668454
rect 415222 668218 415404 668454
rect 414804 668134 415404 668218
rect 414804 667898 414986 668134
rect 415222 667898 415404 668134
rect 414804 632454 415404 667898
rect 414804 632218 414986 632454
rect 415222 632218 415404 632454
rect 414804 632134 415404 632218
rect 414804 631898 414986 632134
rect 415222 631898 415404 632134
rect 414804 596454 415404 631898
rect 414804 596218 414986 596454
rect 415222 596218 415404 596454
rect 414804 596134 415404 596218
rect 414804 595898 414986 596134
rect 415222 595898 415404 596134
rect 414804 584916 415404 595898
rect 432804 704838 433404 705800
rect 432804 704602 432986 704838
rect 433222 704602 433404 704838
rect 432804 704518 433404 704602
rect 432804 704282 432986 704518
rect 433222 704282 433404 704518
rect 432804 686454 433404 704282
rect 432804 686218 432986 686454
rect 433222 686218 433404 686454
rect 432804 686134 433404 686218
rect 432804 685898 432986 686134
rect 433222 685898 433404 686134
rect 432804 650454 433404 685898
rect 432804 650218 432986 650454
rect 433222 650218 433404 650454
rect 432804 650134 433404 650218
rect 432804 649898 432986 650134
rect 433222 649898 433404 650134
rect 432804 614454 433404 649898
rect 432804 614218 432986 614454
rect 433222 614218 433404 614454
rect 432804 614134 433404 614218
rect 432804 613898 432986 614134
rect 433222 613898 433404 614134
rect 432804 584916 433404 613898
rect 450804 705778 451404 705800
rect 450804 705542 450986 705778
rect 451222 705542 451404 705778
rect 450804 705458 451404 705542
rect 450804 705222 450986 705458
rect 451222 705222 451404 705458
rect 450804 668454 451404 705222
rect 450804 668218 450986 668454
rect 451222 668218 451404 668454
rect 450804 668134 451404 668218
rect 450804 667898 450986 668134
rect 451222 667898 451404 668134
rect 450804 632454 451404 667898
rect 450804 632218 450986 632454
rect 451222 632218 451404 632454
rect 450804 632134 451404 632218
rect 450804 631898 450986 632134
rect 451222 631898 451404 632134
rect 450804 596454 451404 631898
rect 450804 596218 450986 596454
rect 451222 596218 451404 596454
rect 450804 596134 451404 596218
rect 450804 595898 450986 596134
rect 451222 595898 451404 596134
rect 450804 584916 451404 595898
rect 468804 704838 469404 705800
rect 468804 704602 468986 704838
rect 469222 704602 469404 704838
rect 468804 704518 469404 704602
rect 468804 704282 468986 704518
rect 469222 704282 469404 704518
rect 468804 686454 469404 704282
rect 468804 686218 468986 686454
rect 469222 686218 469404 686454
rect 468804 686134 469404 686218
rect 468804 685898 468986 686134
rect 469222 685898 469404 686134
rect 468804 650454 469404 685898
rect 468804 650218 468986 650454
rect 469222 650218 469404 650454
rect 468804 650134 469404 650218
rect 468804 649898 468986 650134
rect 469222 649898 469404 650134
rect 468804 614454 469404 649898
rect 468804 614218 468986 614454
rect 469222 614218 469404 614454
rect 468804 614134 469404 614218
rect 468804 613898 468986 614134
rect 469222 613898 469404 614134
rect 468804 584916 469404 613898
rect 486804 705778 487404 705800
rect 486804 705542 486986 705778
rect 487222 705542 487404 705778
rect 486804 705458 487404 705542
rect 486804 705222 486986 705458
rect 487222 705222 487404 705458
rect 486804 668454 487404 705222
rect 486804 668218 486986 668454
rect 487222 668218 487404 668454
rect 486804 668134 487404 668218
rect 486804 667898 486986 668134
rect 487222 667898 487404 668134
rect 486804 632454 487404 667898
rect 486804 632218 486986 632454
rect 487222 632218 487404 632454
rect 486804 632134 487404 632218
rect 486804 631898 486986 632134
rect 487222 631898 487404 632134
rect 486804 596454 487404 631898
rect 486804 596218 486986 596454
rect 487222 596218 487404 596454
rect 486804 596134 487404 596218
rect 486804 595898 486986 596134
rect 487222 595898 487404 596134
rect 486804 584916 487404 595898
rect 504804 704838 505404 705800
rect 504804 704602 504986 704838
rect 505222 704602 505404 704838
rect 504804 704518 505404 704602
rect 504804 704282 504986 704518
rect 505222 704282 505404 704518
rect 504804 686454 505404 704282
rect 504804 686218 504986 686454
rect 505222 686218 505404 686454
rect 504804 686134 505404 686218
rect 504804 685898 504986 686134
rect 505222 685898 505404 686134
rect 504804 650454 505404 685898
rect 504804 650218 504986 650454
rect 505222 650218 505404 650454
rect 504804 650134 505404 650218
rect 504804 649898 504986 650134
rect 505222 649898 505404 650134
rect 504804 614454 505404 649898
rect 504804 614218 504986 614454
rect 505222 614218 505404 614454
rect 504804 614134 505404 614218
rect 504804 613898 504986 614134
rect 505222 613898 505404 614134
rect 504804 584916 505404 613898
rect 522804 705778 523404 705800
rect 522804 705542 522986 705778
rect 523222 705542 523404 705778
rect 522804 705458 523404 705542
rect 522804 705222 522986 705458
rect 523222 705222 523404 705458
rect 522804 668454 523404 705222
rect 522804 668218 522986 668454
rect 523222 668218 523404 668454
rect 522804 668134 523404 668218
rect 522804 667898 522986 668134
rect 523222 667898 523404 668134
rect 522804 632454 523404 667898
rect 522804 632218 522986 632454
rect 523222 632218 523404 632454
rect 522804 632134 523404 632218
rect 522804 631898 522986 632134
rect 523222 631898 523404 632134
rect 522804 596454 523404 631898
rect 522804 596218 522986 596454
rect 523222 596218 523404 596454
rect 522804 596134 523404 596218
rect 522804 595898 522986 596134
rect 523222 595898 523404 596134
rect 522804 584916 523404 595898
rect 540804 704838 541404 705800
rect 540804 704602 540986 704838
rect 541222 704602 541404 704838
rect 540804 704518 541404 704602
rect 540804 704282 540986 704518
rect 541222 704282 541404 704518
rect 540804 686454 541404 704282
rect 540804 686218 540986 686454
rect 541222 686218 541404 686454
rect 540804 686134 541404 686218
rect 540804 685898 540986 686134
rect 541222 685898 541404 686134
rect 540804 650454 541404 685898
rect 540804 650218 540986 650454
rect 541222 650218 541404 650454
rect 540804 650134 541404 650218
rect 540804 649898 540986 650134
rect 541222 649898 541404 650134
rect 540804 614454 541404 649898
rect 540804 614218 540986 614454
rect 541222 614218 541404 614454
rect 540804 614134 541404 614218
rect 540804 613898 540986 614134
rect 541222 613898 541404 614134
rect 540804 584916 541404 613898
rect 558804 705778 559404 705800
rect 558804 705542 558986 705778
rect 559222 705542 559404 705778
rect 558804 705458 559404 705542
rect 558804 705222 558986 705458
rect 559222 705222 559404 705458
rect 558804 668454 559404 705222
rect 558804 668218 558986 668454
rect 559222 668218 559404 668454
rect 558804 668134 559404 668218
rect 558804 667898 558986 668134
rect 559222 667898 559404 668134
rect 558804 632454 559404 667898
rect 558804 632218 558986 632454
rect 559222 632218 559404 632454
rect 558804 632134 559404 632218
rect 558804 631898 558986 632134
rect 559222 631898 559404 632134
rect 558804 596454 559404 631898
rect 558804 596218 558986 596454
rect 559222 596218 559404 596454
rect 558804 596134 559404 596218
rect 558804 595898 558986 596134
rect 559222 595898 559404 596134
rect 558804 584916 559404 595898
rect 576804 704838 577404 705800
rect 586260 705778 586860 705800
rect 586260 705542 586442 705778
rect 586678 705542 586860 705778
rect 586260 705458 586860 705542
rect 586260 705222 586442 705458
rect 586678 705222 586860 705458
rect 576804 704602 576986 704838
rect 577222 704602 577404 704838
rect 576804 704518 577404 704602
rect 576804 704282 576986 704518
rect 577222 704282 577404 704518
rect 576804 686454 577404 704282
rect 576804 686218 576986 686454
rect 577222 686218 577404 686454
rect 576804 686134 577404 686218
rect 576804 685898 576986 686134
rect 577222 685898 577404 686134
rect 576804 650454 577404 685898
rect 576804 650218 576986 650454
rect 577222 650218 577404 650454
rect 576804 650134 577404 650218
rect 576804 649898 576986 650134
rect 577222 649898 577404 650134
rect 576804 614454 577404 649898
rect 576804 614218 576986 614454
rect 577222 614218 577404 614454
rect 576804 614134 577404 614218
rect 576804 613898 576986 614134
rect 577222 613898 577404 614134
rect 554256 578454 554576 578476
rect 554256 578218 554298 578454
rect 554534 578218 554576 578454
rect 554256 578134 554576 578218
rect 554256 577898 554298 578134
rect 554534 577898 554576 578134
rect 554256 577876 554576 577898
rect 576804 578454 577404 613898
rect 576804 578218 576986 578454
rect 577222 578218 577404 578454
rect 576804 578134 577404 578218
rect 576804 577898 576986 578134
rect 577222 577898 577404 578134
rect 538896 560454 539216 560476
rect 538896 560218 538938 560454
rect 539174 560218 539216 560454
rect 538896 560134 539216 560218
rect 538896 559898 538938 560134
rect 539174 559898 539216 560134
rect 538896 559876 539216 559898
rect 554256 542454 554576 542476
rect 554256 542218 554298 542454
rect 554534 542218 554576 542454
rect 554256 542134 554576 542218
rect 554256 541898 554298 542134
rect 554534 541898 554576 542134
rect 554256 541876 554576 541898
rect 576804 542454 577404 577898
rect 576804 542218 576986 542454
rect 577222 542218 577404 542454
rect 576804 542134 577404 542218
rect 576804 541898 576986 542134
rect 577222 541898 577404 542134
rect 538896 524454 539216 524476
rect 538896 524218 538938 524454
rect 539174 524218 539216 524454
rect 538896 524134 539216 524218
rect 538896 523898 538938 524134
rect 539174 523898 539216 524134
rect 538896 523876 539216 523898
rect 554256 506454 554576 506476
rect 554256 506218 554298 506454
rect 554534 506218 554576 506454
rect 554256 506134 554576 506218
rect 554256 505898 554298 506134
rect 554534 505898 554576 506134
rect 554256 505876 554576 505898
rect 576804 506454 577404 541898
rect 576804 506218 576986 506454
rect 577222 506218 577404 506454
rect 576804 506134 577404 506218
rect 576804 505898 576986 506134
rect 577222 505898 577404 506134
rect 538896 488454 539216 488476
rect 538896 488218 538938 488454
rect 539174 488218 539216 488454
rect 538896 488134 539216 488218
rect 538896 487898 538938 488134
rect 539174 487898 539216 488134
rect 538896 487876 539216 487898
rect 554256 470454 554576 470476
rect 554256 470218 554298 470454
rect 554534 470218 554576 470454
rect 554256 470134 554576 470218
rect 554256 469898 554298 470134
rect 554534 469898 554576 470134
rect 554256 469876 554576 469898
rect 576804 470454 577404 505898
rect 576804 470218 576986 470454
rect 577222 470218 577404 470454
rect 576804 470134 577404 470218
rect 576804 469898 576986 470134
rect 577222 469898 577404 470134
rect 538896 452454 539216 452476
rect 538896 452218 538938 452454
rect 539174 452218 539216 452454
rect 538896 452134 539216 452218
rect 538896 451898 538938 452134
rect 539174 451898 539216 452134
rect 538896 451876 539216 451898
rect 554256 434454 554576 434476
rect 554256 434218 554298 434454
rect 554534 434218 554576 434454
rect 554256 434134 554576 434218
rect 554256 433898 554298 434134
rect 554534 433898 554576 434134
rect 554256 433876 554576 433898
rect 576804 434454 577404 469898
rect 576804 434218 576986 434454
rect 577222 434218 577404 434454
rect 576804 434134 577404 434218
rect 576804 433898 576986 434134
rect 577222 433898 577404 434134
rect 538896 416454 539216 416476
rect 538896 416218 538938 416454
rect 539174 416218 539216 416454
rect 538896 416134 539216 416218
rect 538896 415898 538938 416134
rect 539174 415898 539216 416134
rect 538896 415876 539216 415898
rect 554256 398454 554576 398476
rect 554256 398218 554298 398454
rect 554534 398218 554576 398454
rect 554256 398134 554576 398218
rect 554256 397898 554298 398134
rect 554534 397898 554576 398134
rect 554256 397876 554576 397898
rect 576804 398454 577404 433898
rect 576804 398218 576986 398454
rect 577222 398218 577404 398454
rect 576804 398134 577404 398218
rect 576804 397898 576986 398134
rect 577222 397898 577404 398134
rect 324804 362454 325404 382916
rect 324804 362218 324986 362454
rect 325222 362218 325404 362454
rect 324804 362134 325404 362218
rect 324804 361898 324986 362134
rect 325222 361898 325404 362134
rect 310654 334190 311450 334250
rect 311390 333845 311450 334190
rect 311387 333844 311453 333845
rect 311387 333780 311388 333844
rect 311452 333780 311453 333844
rect 311387 333779 311453 333780
rect 309550 332830 309794 332890
rect 307472 326454 307792 326476
rect 307472 326218 307514 326454
rect 307750 326218 307792 326454
rect 307472 326134 307792 326218
rect 307472 325898 307514 326134
rect 307750 325898 307792 326134
rect 307472 325876 307792 325898
rect 309550 322010 309610 332830
rect 324804 326454 325404 361898
rect 324804 326218 324986 326454
rect 325222 326218 325404 326454
rect 324804 326134 325404 326218
rect 324804 325898 324986 326134
rect 325222 325898 325404 326134
rect 309550 321950 309794 322010
rect 309734 316301 309794 321950
rect 309731 316300 309797 316301
rect 309731 316236 309732 316300
rect 309796 316236 309797 316300
rect 309731 316235 309797 316236
rect 306603 315620 306669 315621
rect 306603 315556 306604 315620
rect 306668 315556 306669 315620
rect 306603 315555 306669 315556
rect 306804 308454 307404 314560
rect 306804 308218 306986 308454
rect 307222 308218 307404 308454
rect 306804 308134 307404 308218
rect 306804 307898 306986 308134
rect 307222 307898 307404 308134
rect 306419 276724 306485 276725
rect 306419 276660 306420 276724
rect 306484 276660 306485 276724
rect 306419 276659 306485 276660
rect 306804 272454 307404 307898
rect 324804 290454 325404 325898
rect 324804 290218 324986 290454
rect 325222 290218 325404 290454
rect 324804 290134 325404 290218
rect 324804 289898 324986 290134
rect 325222 289898 325404 290134
rect 324804 274600 325404 289898
rect 342804 380454 343404 382916
rect 342804 380218 342986 380454
rect 343222 380218 343404 380454
rect 342804 380134 343404 380218
rect 342804 379898 342986 380134
rect 343222 379898 343404 380134
rect 342804 344454 343404 379898
rect 342804 344218 342986 344454
rect 343222 344218 343404 344454
rect 342804 344134 343404 344218
rect 342804 343898 342986 344134
rect 343222 343898 343404 344134
rect 342804 308454 343404 343898
rect 342804 308218 342986 308454
rect 343222 308218 343404 308454
rect 342804 308134 343404 308218
rect 342804 307898 342986 308134
rect 343222 307898 343404 308134
rect 342804 274600 343404 307898
rect 360804 362454 361404 382916
rect 360804 362218 360986 362454
rect 361222 362218 361404 362454
rect 360804 362134 361404 362218
rect 360804 361898 360986 362134
rect 361222 361898 361404 362134
rect 360804 326454 361404 361898
rect 360804 326218 360986 326454
rect 361222 326218 361404 326454
rect 360804 326134 361404 326218
rect 360804 325898 360986 326134
rect 361222 325898 361404 326134
rect 360804 290454 361404 325898
rect 360804 290218 360986 290454
rect 361222 290218 361404 290454
rect 360804 290134 361404 290218
rect 360804 289898 360986 290134
rect 361222 289898 361404 290134
rect 360804 274600 361404 289898
rect 378804 380454 379404 382916
rect 378804 380218 378986 380454
rect 379222 380218 379404 380454
rect 378804 380134 379404 380218
rect 378804 379898 378986 380134
rect 379222 379898 379404 380134
rect 378804 344454 379404 379898
rect 378804 344218 378986 344454
rect 379222 344218 379404 344454
rect 378804 344134 379404 344218
rect 378804 343898 378986 344134
rect 379222 343898 379404 344134
rect 378804 308454 379404 343898
rect 378804 308218 378986 308454
rect 379222 308218 379404 308454
rect 378804 308134 379404 308218
rect 378804 307898 378986 308134
rect 379222 307898 379404 308134
rect 378804 274600 379404 307898
rect 396804 362454 397404 382916
rect 396804 362218 396986 362454
rect 397222 362218 397404 362454
rect 396804 362134 397404 362218
rect 396804 361898 396986 362134
rect 397222 361898 397404 362134
rect 396804 326454 397404 361898
rect 396804 326218 396986 326454
rect 397222 326218 397404 326454
rect 396804 326134 397404 326218
rect 396804 325898 396986 326134
rect 397222 325898 397404 326134
rect 396804 290454 397404 325898
rect 396804 290218 396986 290454
rect 397222 290218 397404 290454
rect 396804 290134 397404 290218
rect 396804 289898 396986 290134
rect 397222 289898 397404 290134
rect 396804 274600 397404 289898
rect 414804 380454 415404 382916
rect 414804 380218 414986 380454
rect 415222 380218 415404 380454
rect 414804 380134 415404 380218
rect 414804 379898 414986 380134
rect 415222 379898 415404 380134
rect 414804 344454 415404 379898
rect 414804 344218 414986 344454
rect 415222 344218 415404 344454
rect 414804 344134 415404 344218
rect 414804 343898 414986 344134
rect 415222 343898 415404 344134
rect 414804 308454 415404 343898
rect 414804 308218 414986 308454
rect 415222 308218 415404 308454
rect 414804 308134 415404 308218
rect 414804 307898 414986 308134
rect 415222 307898 415404 308134
rect 414804 274600 415404 307898
rect 432804 362454 433404 382916
rect 432804 362218 432986 362454
rect 433222 362218 433404 362454
rect 432804 362134 433404 362218
rect 432804 361898 432986 362134
rect 433222 361898 433404 362134
rect 432804 326454 433404 361898
rect 432804 326218 432986 326454
rect 433222 326218 433404 326454
rect 432804 326134 433404 326218
rect 432804 325898 432986 326134
rect 433222 325898 433404 326134
rect 432804 290454 433404 325898
rect 432804 290218 432986 290454
rect 433222 290218 433404 290454
rect 432804 290134 433404 290218
rect 432804 289898 432986 290134
rect 433222 289898 433404 290134
rect 432804 274600 433404 289898
rect 450804 380454 451404 382916
rect 450804 380218 450986 380454
rect 451222 380218 451404 380454
rect 450804 380134 451404 380218
rect 450804 379898 450986 380134
rect 451222 379898 451404 380134
rect 450804 344454 451404 379898
rect 450804 344218 450986 344454
rect 451222 344218 451404 344454
rect 450804 344134 451404 344218
rect 450804 343898 450986 344134
rect 451222 343898 451404 344134
rect 450804 308454 451404 343898
rect 450804 308218 450986 308454
rect 451222 308218 451404 308454
rect 450804 308134 451404 308218
rect 450804 307898 450986 308134
rect 451222 307898 451404 308134
rect 450804 274600 451404 307898
rect 468804 362454 469404 382916
rect 468804 362218 468986 362454
rect 469222 362218 469404 362454
rect 468804 362134 469404 362218
rect 468804 361898 468986 362134
rect 469222 361898 469404 362134
rect 468804 326454 469404 361898
rect 468804 326218 468986 326454
rect 469222 326218 469404 326454
rect 468804 326134 469404 326218
rect 468804 325898 468986 326134
rect 469222 325898 469404 326134
rect 468804 290454 469404 325898
rect 468804 290218 468986 290454
rect 469222 290218 469404 290454
rect 468804 290134 469404 290218
rect 468804 289898 468986 290134
rect 469222 289898 469404 290134
rect 468804 274600 469404 289898
rect 486804 380454 487404 382916
rect 486804 380218 486986 380454
rect 487222 380218 487404 380454
rect 486804 380134 487404 380218
rect 486804 379898 486986 380134
rect 487222 379898 487404 380134
rect 486804 344454 487404 379898
rect 486804 344218 486986 344454
rect 487222 344218 487404 344454
rect 486804 344134 487404 344218
rect 486804 343898 486986 344134
rect 487222 343898 487404 344134
rect 486804 308454 487404 343898
rect 486804 308218 486986 308454
rect 487222 308218 487404 308454
rect 486804 308134 487404 308218
rect 486804 307898 486986 308134
rect 487222 307898 487404 308134
rect 486804 274600 487404 307898
rect 504804 362454 505404 382916
rect 504804 362218 504986 362454
rect 505222 362218 505404 362454
rect 504804 362134 505404 362218
rect 504804 361898 504986 362134
rect 505222 361898 505404 362134
rect 504804 326454 505404 361898
rect 504804 326218 504986 326454
rect 505222 326218 505404 326454
rect 504804 326134 505404 326218
rect 504804 325898 504986 326134
rect 505222 325898 505404 326134
rect 504804 290454 505404 325898
rect 504804 290218 504986 290454
rect 505222 290218 505404 290454
rect 504804 290134 505404 290218
rect 504804 289898 504986 290134
rect 505222 289898 505404 290134
rect 504804 274600 505404 289898
rect 522804 380454 523404 382916
rect 522804 380218 522986 380454
rect 523222 380218 523404 380454
rect 522804 380134 523404 380218
rect 522804 379898 522986 380134
rect 523222 379898 523404 380134
rect 522804 344454 523404 379898
rect 522804 344218 522986 344454
rect 523222 344218 523404 344454
rect 522804 344134 523404 344218
rect 522804 343898 522986 344134
rect 523222 343898 523404 344134
rect 522804 308454 523404 343898
rect 522804 308218 522986 308454
rect 523222 308218 523404 308454
rect 522804 308134 523404 308218
rect 522804 307898 522986 308134
rect 523222 307898 523404 308134
rect 522804 274600 523404 307898
rect 540804 362454 541404 382916
rect 540804 362218 540986 362454
rect 541222 362218 541404 362454
rect 540804 362134 541404 362218
rect 540804 361898 540986 362134
rect 541222 361898 541404 362134
rect 540804 326454 541404 361898
rect 540804 326218 540986 326454
rect 541222 326218 541404 326454
rect 540804 326134 541404 326218
rect 540804 325898 540986 326134
rect 541222 325898 541404 326134
rect 540804 290454 541404 325898
rect 540804 290218 540986 290454
rect 541222 290218 541404 290454
rect 540804 290134 541404 290218
rect 540804 289898 540986 290134
rect 541222 289898 541404 290134
rect 540804 274600 541404 289898
rect 558804 380454 559404 382916
rect 558804 380218 558986 380454
rect 559222 380218 559404 380454
rect 558804 380134 559404 380218
rect 558804 379898 558986 380134
rect 559222 379898 559404 380134
rect 558804 344454 559404 379898
rect 558804 344218 558986 344454
rect 559222 344218 559404 344454
rect 558804 344134 559404 344218
rect 558804 343898 558986 344134
rect 559222 343898 559404 344134
rect 558804 308454 559404 343898
rect 558804 308218 558986 308454
rect 559222 308218 559404 308454
rect 558804 308134 559404 308218
rect 558804 307898 558986 308134
rect 559222 307898 559404 308134
rect 558804 274600 559404 307898
rect 576804 362454 577404 397898
rect 576804 362218 576986 362454
rect 577222 362218 577404 362454
rect 576804 362134 577404 362218
rect 576804 361898 576986 362134
rect 577222 361898 577404 362134
rect 576804 326454 577404 361898
rect 576804 326218 576986 326454
rect 577222 326218 577404 326454
rect 576804 326134 577404 326218
rect 576804 325898 576986 326134
rect 577222 325898 577404 326134
rect 576804 290454 577404 325898
rect 576804 290218 576986 290454
rect 577222 290218 577404 290454
rect 576804 290134 577404 290218
rect 576804 289898 576986 290134
rect 577222 289898 577404 290134
rect 306804 272218 306986 272454
rect 307222 272218 307404 272454
rect 306804 272134 307404 272218
rect 306804 271898 306986 272134
rect 307222 271898 307404 272134
rect 306804 236454 307404 271898
rect 554256 254454 554576 254476
rect 554256 254218 554298 254454
rect 554534 254218 554576 254454
rect 554256 254134 554576 254218
rect 554256 253898 554298 254134
rect 554534 253898 554576 254134
rect 554256 253876 554576 253898
rect 576804 254454 577404 289898
rect 576804 254218 576986 254454
rect 577222 254218 577404 254454
rect 576804 254134 577404 254218
rect 576804 253898 576986 254134
rect 577222 253898 577404 254134
rect 306804 236218 306986 236454
rect 307222 236218 307404 236454
rect 306804 236134 307404 236218
rect 306804 235898 306986 236134
rect 307222 235898 307404 236134
rect 306804 200454 307404 235898
rect 538896 236454 539216 236476
rect 538896 236218 538938 236454
rect 539174 236218 539216 236454
rect 538896 236134 539216 236218
rect 538896 235898 538938 236134
rect 539174 235898 539216 236134
rect 538896 235876 539216 235898
rect 554256 218454 554576 218476
rect 554256 218218 554298 218454
rect 554534 218218 554576 218454
rect 554256 218134 554576 218218
rect 554256 217898 554298 218134
rect 554534 217898 554576 218134
rect 554256 217876 554576 217898
rect 576804 218454 577404 253898
rect 576804 218218 576986 218454
rect 577222 218218 577404 218454
rect 576804 218134 577404 218218
rect 576804 217898 576986 218134
rect 577222 217898 577404 218134
rect 306804 200218 306986 200454
rect 307222 200218 307404 200454
rect 306804 200134 307404 200218
rect 306804 199898 306986 200134
rect 307222 199898 307404 200134
rect 306804 164454 307404 199898
rect 538896 200454 539216 200476
rect 538896 200218 538938 200454
rect 539174 200218 539216 200454
rect 538896 200134 539216 200218
rect 538896 199898 538938 200134
rect 539174 199898 539216 200134
rect 538896 199876 539216 199898
rect 554256 182454 554576 182476
rect 554256 182218 554298 182454
rect 554534 182218 554576 182454
rect 554256 182134 554576 182218
rect 554256 181898 554298 182134
rect 554534 181898 554576 182134
rect 554256 181876 554576 181898
rect 576804 182454 577404 217898
rect 576804 182218 576986 182454
rect 577222 182218 577404 182454
rect 576804 182134 577404 182218
rect 576804 181898 576986 182134
rect 577222 181898 577404 182134
rect 306804 164218 306986 164454
rect 307222 164218 307404 164454
rect 306804 164134 307404 164218
rect 306804 163898 306986 164134
rect 307222 163898 307404 164134
rect 306804 128454 307404 163898
rect 538896 164454 539216 164476
rect 538896 164218 538938 164454
rect 539174 164218 539216 164454
rect 538896 164134 539216 164218
rect 538896 163898 538938 164134
rect 539174 163898 539216 164134
rect 538896 163876 539216 163898
rect 554256 146454 554576 146476
rect 554256 146218 554298 146454
rect 554534 146218 554576 146454
rect 554256 146134 554576 146218
rect 554256 145898 554298 146134
rect 554534 145898 554576 146134
rect 554256 145876 554576 145898
rect 576804 146454 577404 181898
rect 576804 146218 576986 146454
rect 577222 146218 577404 146454
rect 576804 146134 577404 146218
rect 576804 145898 576986 146134
rect 577222 145898 577404 146134
rect 306804 128218 306986 128454
rect 307222 128218 307404 128454
rect 306804 128134 307404 128218
rect 306804 127898 306986 128134
rect 307222 127898 307404 128134
rect 299427 92716 299493 92717
rect 299427 92652 299428 92716
rect 299492 92652 299493 92716
rect 299427 92651 299493 92652
rect 306804 92454 307404 127898
rect 538896 128454 539216 128476
rect 538896 128218 538938 128454
rect 539174 128218 539216 128454
rect 538896 128134 539216 128218
rect 538896 127898 538938 128134
rect 539174 127898 539216 128134
rect 538896 127876 539216 127898
rect 554256 110454 554576 110476
rect 554256 110218 554298 110454
rect 554534 110218 554576 110454
rect 554256 110134 554576 110218
rect 554256 109898 554298 110134
rect 554534 109898 554576 110134
rect 554256 109876 554576 109898
rect 576804 110454 577404 145898
rect 576804 110218 576986 110454
rect 577222 110218 577404 110454
rect 576804 110134 577404 110218
rect 576804 109898 576986 110134
rect 577222 109898 577404 110134
rect 306804 92218 306986 92454
rect 307222 92218 307404 92454
rect 306804 92134 307404 92218
rect 306804 91898 306986 92134
rect 307222 91898 307404 92134
rect 306804 56454 307404 91898
rect 538896 92454 539216 92476
rect 538896 92218 538938 92454
rect 539174 92218 539216 92454
rect 538896 92134 539216 92218
rect 538896 91898 538938 92134
rect 539174 91898 539216 92134
rect 538896 91876 539216 91898
rect 576804 74454 577404 109898
rect 576804 74218 576986 74454
rect 577222 74218 577404 74454
rect 576804 74134 577404 74218
rect 576804 73898 576986 74134
rect 577222 73898 577404 74134
rect 306804 56218 306986 56454
rect 307222 56218 307404 56454
rect 306804 56134 307404 56218
rect 306804 55898 306986 56134
rect 307222 55898 307404 56134
rect 306804 20454 307404 55898
rect 306804 20218 306986 20454
rect 307222 20218 307404 20454
rect 306804 20134 307404 20218
rect 306804 19898 306986 20134
rect 307222 19898 307404 20134
rect 298691 3636 298757 3637
rect 298691 3572 298692 3636
rect 298756 3572 298757 3636
rect 298691 3571 298757 3572
rect 288804 2218 288986 2454
rect 289222 2218 289404 2454
rect 288804 2134 289404 2218
rect 288804 1898 288986 2134
rect 289222 1898 289404 2134
rect 288804 -346 289404 1898
rect 288804 -582 288986 -346
rect 289222 -582 289404 -346
rect 288804 -666 289404 -582
rect 288804 -902 288986 -666
rect 289222 -902 289404 -666
rect 288804 -1864 289404 -902
rect 306804 -1286 307404 19898
rect 306804 -1522 306986 -1286
rect 307222 -1522 307404 -1286
rect 306804 -1606 307404 -1522
rect 306804 -1842 306986 -1606
rect 307222 -1842 307404 -1606
rect 306804 -1864 307404 -1842
rect 324804 38454 325404 72600
rect 324804 38218 324986 38454
rect 325222 38218 325404 38454
rect 324804 38134 325404 38218
rect 324804 37898 324986 38134
rect 325222 37898 325404 38134
rect 324804 2454 325404 37898
rect 324804 2218 324986 2454
rect 325222 2218 325404 2454
rect 324804 2134 325404 2218
rect 324804 1898 324986 2134
rect 325222 1898 325404 2134
rect 324804 -346 325404 1898
rect 324804 -582 324986 -346
rect 325222 -582 325404 -346
rect 324804 -666 325404 -582
rect 324804 -902 324986 -666
rect 325222 -902 325404 -666
rect 324804 -1864 325404 -902
rect 342804 56454 343404 72600
rect 342804 56218 342986 56454
rect 343222 56218 343404 56454
rect 342804 56134 343404 56218
rect 342804 55898 342986 56134
rect 343222 55898 343404 56134
rect 342804 20454 343404 55898
rect 342804 20218 342986 20454
rect 343222 20218 343404 20454
rect 342804 20134 343404 20218
rect 342804 19898 342986 20134
rect 343222 19898 343404 20134
rect 342804 -1286 343404 19898
rect 342804 -1522 342986 -1286
rect 343222 -1522 343404 -1286
rect 342804 -1606 343404 -1522
rect 342804 -1842 342986 -1606
rect 343222 -1842 343404 -1606
rect 342804 -1864 343404 -1842
rect 360804 38454 361404 72600
rect 360804 38218 360986 38454
rect 361222 38218 361404 38454
rect 360804 38134 361404 38218
rect 360804 37898 360986 38134
rect 361222 37898 361404 38134
rect 360804 2454 361404 37898
rect 360804 2218 360986 2454
rect 361222 2218 361404 2454
rect 360804 2134 361404 2218
rect 360804 1898 360986 2134
rect 361222 1898 361404 2134
rect 360804 -346 361404 1898
rect 360804 -582 360986 -346
rect 361222 -582 361404 -346
rect 360804 -666 361404 -582
rect 360804 -902 360986 -666
rect 361222 -902 361404 -666
rect 360804 -1864 361404 -902
rect 378804 56454 379404 72600
rect 378804 56218 378986 56454
rect 379222 56218 379404 56454
rect 378804 56134 379404 56218
rect 378804 55898 378986 56134
rect 379222 55898 379404 56134
rect 378804 20454 379404 55898
rect 378804 20218 378986 20454
rect 379222 20218 379404 20454
rect 378804 20134 379404 20218
rect 378804 19898 378986 20134
rect 379222 19898 379404 20134
rect 378804 -1286 379404 19898
rect 378804 -1522 378986 -1286
rect 379222 -1522 379404 -1286
rect 378804 -1606 379404 -1522
rect 378804 -1842 378986 -1606
rect 379222 -1842 379404 -1606
rect 378804 -1864 379404 -1842
rect 396804 38454 397404 72600
rect 396804 38218 396986 38454
rect 397222 38218 397404 38454
rect 396804 38134 397404 38218
rect 396804 37898 396986 38134
rect 397222 37898 397404 38134
rect 396804 2454 397404 37898
rect 396804 2218 396986 2454
rect 397222 2218 397404 2454
rect 396804 2134 397404 2218
rect 396804 1898 396986 2134
rect 397222 1898 397404 2134
rect 396804 -346 397404 1898
rect 396804 -582 396986 -346
rect 397222 -582 397404 -346
rect 396804 -666 397404 -582
rect 396804 -902 396986 -666
rect 397222 -902 397404 -666
rect 396804 -1864 397404 -902
rect 414804 56454 415404 72600
rect 414804 56218 414986 56454
rect 415222 56218 415404 56454
rect 414804 56134 415404 56218
rect 414804 55898 414986 56134
rect 415222 55898 415404 56134
rect 414804 20454 415404 55898
rect 414804 20218 414986 20454
rect 415222 20218 415404 20454
rect 414804 20134 415404 20218
rect 414804 19898 414986 20134
rect 415222 19898 415404 20134
rect 414804 -1286 415404 19898
rect 414804 -1522 414986 -1286
rect 415222 -1522 415404 -1286
rect 414804 -1606 415404 -1522
rect 414804 -1842 414986 -1606
rect 415222 -1842 415404 -1606
rect 414804 -1864 415404 -1842
rect 432804 38454 433404 72600
rect 432804 38218 432986 38454
rect 433222 38218 433404 38454
rect 432804 38134 433404 38218
rect 432804 37898 432986 38134
rect 433222 37898 433404 38134
rect 432804 2454 433404 37898
rect 432804 2218 432986 2454
rect 433222 2218 433404 2454
rect 432804 2134 433404 2218
rect 432804 1898 432986 2134
rect 433222 1898 433404 2134
rect 432804 -346 433404 1898
rect 432804 -582 432986 -346
rect 433222 -582 433404 -346
rect 432804 -666 433404 -582
rect 432804 -902 432986 -666
rect 433222 -902 433404 -666
rect 432804 -1864 433404 -902
rect 450804 56454 451404 72600
rect 450804 56218 450986 56454
rect 451222 56218 451404 56454
rect 450804 56134 451404 56218
rect 450804 55898 450986 56134
rect 451222 55898 451404 56134
rect 450804 20454 451404 55898
rect 450804 20218 450986 20454
rect 451222 20218 451404 20454
rect 450804 20134 451404 20218
rect 450804 19898 450986 20134
rect 451222 19898 451404 20134
rect 450804 -1286 451404 19898
rect 450804 -1522 450986 -1286
rect 451222 -1522 451404 -1286
rect 450804 -1606 451404 -1522
rect 450804 -1842 450986 -1606
rect 451222 -1842 451404 -1606
rect 450804 -1864 451404 -1842
rect 468804 38454 469404 72600
rect 468804 38218 468986 38454
rect 469222 38218 469404 38454
rect 468804 38134 469404 38218
rect 468804 37898 468986 38134
rect 469222 37898 469404 38134
rect 468804 2454 469404 37898
rect 468804 2218 468986 2454
rect 469222 2218 469404 2454
rect 468804 2134 469404 2218
rect 468804 1898 468986 2134
rect 469222 1898 469404 2134
rect 468804 -346 469404 1898
rect 468804 -582 468986 -346
rect 469222 -582 469404 -346
rect 468804 -666 469404 -582
rect 468804 -902 468986 -666
rect 469222 -902 469404 -666
rect 468804 -1864 469404 -902
rect 486804 56454 487404 72600
rect 486804 56218 486986 56454
rect 487222 56218 487404 56454
rect 486804 56134 487404 56218
rect 486804 55898 486986 56134
rect 487222 55898 487404 56134
rect 486804 20454 487404 55898
rect 486804 20218 486986 20454
rect 487222 20218 487404 20454
rect 486804 20134 487404 20218
rect 486804 19898 486986 20134
rect 487222 19898 487404 20134
rect 486804 -1286 487404 19898
rect 486804 -1522 486986 -1286
rect 487222 -1522 487404 -1286
rect 486804 -1606 487404 -1522
rect 486804 -1842 486986 -1606
rect 487222 -1842 487404 -1606
rect 486804 -1864 487404 -1842
rect 504804 38454 505404 72600
rect 504804 38218 504986 38454
rect 505222 38218 505404 38454
rect 504804 38134 505404 38218
rect 504804 37898 504986 38134
rect 505222 37898 505404 38134
rect 504804 2454 505404 37898
rect 504804 2218 504986 2454
rect 505222 2218 505404 2454
rect 504804 2134 505404 2218
rect 504804 1898 504986 2134
rect 505222 1898 505404 2134
rect 504804 -346 505404 1898
rect 504804 -582 504986 -346
rect 505222 -582 505404 -346
rect 504804 -666 505404 -582
rect 504804 -902 504986 -666
rect 505222 -902 505404 -666
rect 504804 -1864 505404 -902
rect 522804 56454 523404 72600
rect 522804 56218 522986 56454
rect 523222 56218 523404 56454
rect 522804 56134 523404 56218
rect 522804 55898 522986 56134
rect 523222 55898 523404 56134
rect 522804 20454 523404 55898
rect 522804 20218 522986 20454
rect 523222 20218 523404 20454
rect 522804 20134 523404 20218
rect 522804 19898 522986 20134
rect 523222 19898 523404 20134
rect 522804 -1286 523404 19898
rect 522804 -1522 522986 -1286
rect 523222 -1522 523404 -1286
rect 522804 -1606 523404 -1522
rect 522804 -1842 522986 -1606
rect 523222 -1842 523404 -1606
rect 522804 -1864 523404 -1842
rect 540804 38454 541404 72600
rect 540804 38218 540986 38454
rect 541222 38218 541404 38454
rect 540804 38134 541404 38218
rect 540804 37898 540986 38134
rect 541222 37898 541404 38134
rect 540804 2454 541404 37898
rect 540804 2218 540986 2454
rect 541222 2218 541404 2454
rect 540804 2134 541404 2218
rect 540804 1898 540986 2134
rect 541222 1898 541404 2134
rect 540804 -346 541404 1898
rect 540804 -582 540986 -346
rect 541222 -582 541404 -346
rect 540804 -666 541404 -582
rect 540804 -902 540986 -666
rect 541222 -902 541404 -666
rect 540804 -1864 541404 -902
rect 558804 56454 559404 72600
rect 558804 56218 558986 56454
rect 559222 56218 559404 56454
rect 558804 56134 559404 56218
rect 558804 55898 558986 56134
rect 559222 55898 559404 56134
rect 558804 20454 559404 55898
rect 558804 20218 558986 20454
rect 559222 20218 559404 20454
rect 558804 20134 559404 20218
rect 558804 19898 558986 20134
rect 559222 19898 559404 20134
rect 558804 -1286 559404 19898
rect 558804 -1522 558986 -1286
rect 559222 -1522 559404 -1286
rect 558804 -1606 559404 -1522
rect 558804 -1842 558986 -1606
rect 559222 -1842 559404 -1606
rect 558804 -1864 559404 -1842
rect 576804 38454 577404 73898
rect 576804 38218 576986 38454
rect 577222 38218 577404 38454
rect 576804 38134 577404 38218
rect 576804 37898 576986 38134
rect 577222 37898 577404 38134
rect 576804 2454 577404 37898
rect 576804 2218 576986 2454
rect 577222 2218 577404 2454
rect 576804 2134 577404 2218
rect 576804 1898 576986 2134
rect 577222 1898 577404 2134
rect 576804 -346 577404 1898
rect 576804 -582 576986 -346
rect 577222 -582 577404 -346
rect 576804 -666 577404 -582
rect 576804 -902 576986 -666
rect 577222 -902 577404 -666
rect 576804 -1864 577404 -902
rect 585320 704838 585920 704860
rect 585320 704602 585502 704838
rect 585738 704602 585920 704838
rect 585320 704518 585920 704602
rect 585320 704282 585502 704518
rect 585738 704282 585920 704518
rect 585320 686454 585920 704282
rect 585320 686218 585502 686454
rect 585738 686218 585920 686454
rect 585320 686134 585920 686218
rect 585320 685898 585502 686134
rect 585738 685898 585920 686134
rect 585320 650454 585920 685898
rect 585320 650218 585502 650454
rect 585738 650218 585920 650454
rect 585320 650134 585920 650218
rect 585320 649898 585502 650134
rect 585738 649898 585920 650134
rect 585320 614454 585920 649898
rect 585320 614218 585502 614454
rect 585738 614218 585920 614454
rect 585320 614134 585920 614218
rect 585320 613898 585502 614134
rect 585738 613898 585920 614134
rect 585320 578454 585920 613898
rect 585320 578218 585502 578454
rect 585738 578218 585920 578454
rect 585320 578134 585920 578218
rect 585320 577898 585502 578134
rect 585738 577898 585920 578134
rect 585320 542454 585920 577898
rect 585320 542218 585502 542454
rect 585738 542218 585920 542454
rect 585320 542134 585920 542218
rect 585320 541898 585502 542134
rect 585738 541898 585920 542134
rect 585320 506454 585920 541898
rect 585320 506218 585502 506454
rect 585738 506218 585920 506454
rect 585320 506134 585920 506218
rect 585320 505898 585502 506134
rect 585738 505898 585920 506134
rect 585320 470454 585920 505898
rect 585320 470218 585502 470454
rect 585738 470218 585920 470454
rect 585320 470134 585920 470218
rect 585320 469898 585502 470134
rect 585738 469898 585920 470134
rect 585320 434454 585920 469898
rect 585320 434218 585502 434454
rect 585738 434218 585920 434454
rect 585320 434134 585920 434218
rect 585320 433898 585502 434134
rect 585738 433898 585920 434134
rect 585320 398454 585920 433898
rect 585320 398218 585502 398454
rect 585738 398218 585920 398454
rect 585320 398134 585920 398218
rect 585320 397898 585502 398134
rect 585738 397898 585920 398134
rect 585320 362454 585920 397898
rect 585320 362218 585502 362454
rect 585738 362218 585920 362454
rect 585320 362134 585920 362218
rect 585320 361898 585502 362134
rect 585738 361898 585920 362134
rect 585320 326454 585920 361898
rect 585320 326218 585502 326454
rect 585738 326218 585920 326454
rect 585320 326134 585920 326218
rect 585320 325898 585502 326134
rect 585738 325898 585920 326134
rect 585320 290454 585920 325898
rect 585320 290218 585502 290454
rect 585738 290218 585920 290454
rect 585320 290134 585920 290218
rect 585320 289898 585502 290134
rect 585738 289898 585920 290134
rect 585320 254454 585920 289898
rect 585320 254218 585502 254454
rect 585738 254218 585920 254454
rect 585320 254134 585920 254218
rect 585320 253898 585502 254134
rect 585738 253898 585920 254134
rect 585320 218454 585920 253898
rect 585320 218218 585502 218454
rect 585738 218218 585920 218454
rect 585320 218134 585920 218218
rect 585320 217898 585502 218134
rect 585738 217898 585920 218134
rect 585320 182454 585920 217898
rect 585320 182218 585502 182454
rect 585738 182218 585920 182454
rect 585320 182134 585920 182218
rect 585320 181898 585502 182134
rect 585738 181898 585920 182134
rect 585320 146454 585920 181898
rect 585320 146218 585502 146454
rect 585738 146218 585920 146454
rect 585320 146134 585920 146218
rect 585320 145898 585502 146134
rect 585738 145898 585920 146134
rect 585320 110454 585920 145898
rect 585320 110218 585502 110454
rect 585738 110218 585920 110454
rect 585320 110134 585920 110218
rect 585320 109898 585502 110134
rect 585738 109898 585920 110134
rect 585320 74454 585920 109898
rect 585320 74218 585502 74454
rect 585738 74218 585920 74454
rect 585320 74134 585920 74218
rect 585320 73898 585502 74134
rect 585738 73898 585920 74134
rect 585320 38454 585920 73898
rect 585320 38218 585502 38454
rect 585738 38218 585920 38454
rect 585320 38134 585920 38218
rect 585320 37898 585502 38134
rect 585738 37898 585920 38134
rect 585320 2454 585920 37898
rect 585320 2218 585502 2454
rect 585738 2218 585920 2454
rect 585320 2134 585920 2218
rect 585320 1898 585502 2134
rect 585738 1898 585920 2134
rect 585320 -346 585920 1898
rect 585320 -582 585502 -346
rect 585738 -582 585920 -346
rect 585320 -666 585920 -582
rect 585320 -902 585502 -666
rect 585738 -902 585920 -666
rect 585320 -924 585920 -902
rect 586260 668454 586860 705222
rect 586260 668218 586442 668454
rect 586678 668218 586860 668454
rect 586260 668134 586860 668218
rect 586260 667898 586442 668134
rect 586678 667898 586860 668134
rect 586260 632454 586860 667898
rect 586260 632218 586442 632454
rect 586678 632218 586860 632454
rect 586260 632134 586860 632218
rect 586260 631898 586442 632134
rect 586678 631898 586860 632134
rect 586260 596454 586860 631898
rect 586260 596218 586442 596454
rect 586678 596218 586860 596454
rect 586260 596134 586860 596218
rect 586260 595898 586442 596134
rect 586678 595898 586860 596134
rect 586260 560454 586860 595898
rect 586260 560218 586442 560454
rect 586678 560218 586860 560454
rect 586260 560134 586860 560218
rect 586260 559898 586442 560134
rect 586678 559898 586860 560134
rect 586260 524454 586860 559898
rect 586260 524218 586442 524454
rect 586678 524218 586860 524454
rect 586260 524134 586860 524218
rect 586260 523898 586442 524134
rect 586678 523898 586860 524134
rect 586260 488454 586860 523898
rect 586260 488218 586442 488454
rect 586678 488218 586860 488454
rect 586260 488134 586860 488218
rect 586260 487898 586442 488134
rect 586678 487898 586860 488134
rect 586260 452454 586860 487898
rect 586260 452218 586442 452454
rect 586678 452218 586860 452454
rect 586260 452134 586860 452218
rect 586260 451898 586442 452134
rect 586678 451898 586860 452134
rect 586260 416454 586860 451898
rect 586260 416218 586442 416454
rect 586678 416218 586860 416454
rect 586260 416134 586860 416218
rect 586260 415898 586442 416134
rect 586678 415898 586860 416134
rect 586260 380454 586860 415898
rect 586260 380218 586442 380454
rect 586678 380218 586860 380454
rect 586260 380134 586860 380218
rect 586260 379898 586442 380134
rect 586678 379898 586860 380134
rect 586260 344454 586860 379898
rect 586260 344218 586442 344454
rect 586678 344218 586860 344454
rect 586260 344134 586860 344218
rect 586260 343898 586442 344134
rect 586678 343898 586860 344134
rect 586260 308454 586860 343898
rect 586260 308218 586442 308454
rect 586678 308218 586860 308454
rect 586260 308134 586860 308218
rect 586260 307898 586442 308134
rect 586678 307898 586860 308134
rect 586260 272454 586860 307898
rect 586260 272218 586442 272454
rect 586678 272218 586860 272454
rect 586260 272134 586860 272218
rect 586260 271898 586442 272134
rect 586678 271898 586860 272134
rect 586260 236454 586860 271898
rect 586260 236218 586442 236454
rect 586678 236218 586860 236454
rect 586260 236134 586860 236218
rect 586260 235898 586442 236134
rect 586678 235898 586860 236134
rect 586260 200454 586860 235898
rect 586260 200218 586442 200454
rect 586678 200218 586860 200454
rect 586260 200134 586860 200218
rect 586260 199898 586442 200134
rect 586678 199898 586860 200134
rect 586260 164454 586860 199898
rect 586260 164218 586442 164454
rect 586678 164218 586860 164454
rect 586260 164134 586860 164218
rect 586260 163898 586442 164134
rect 586678 163898 586860 164134
rect 586260 128454 586860 163898
rect 586260 128218 586442 128454
rect 586678 128218 586860 128454
rect 586260 128134 586860 128218
rect 586260 127898 586442 128134
rect 586678 127898 586860 128134
rect 586260 92454 586860 127898
rect 586260 92218 586442 92454
rect 586678 92218 586860 92454
rect 586260 92134 586860 92218
rect 586260 91898 586442 92134
rect 586678 91898 586860 92134
rect 586260 56454 586860 91898
rect 586260 56218 586442 56454
rect 586678 56218 586860 56454
rect 586260 56134 586860 56218
rect 586260 55898 586442 56134
rect 586678 55898 586860 56134
rect 586260 20454 586860 55898
rect 586260 20218 586442 20454
rect 586678 20218 586860 20454
rect 586260 20134 586860 20218
rect 586260 19898 586442 20134
rect 586678 19898 586860 20134
rect 586260 -1286 586860 19898
rect 586260 -1522 586442 -1286
rect 586678 -1522 586860 -1286
rect 586260 -1606 586860 -1522
rect 586260 -1842 586442 -1606
rect 586678 -1842 586860 -1606
rect 586260 -1864 586860 -1842
rect -3876 -2462 -3694 -2226
rect -3458 -2462 -3276 -2226
rect -3876 -2546 -3276 -2462
rect -3876 -2782 -3694 -2546
rect -3458 -2782 -3276 -2546
rect -3876 -2804 -3276 -2782
rect 587200 -2226 587800 706162
rect 587200 -2462 587382 -2226
rect 587618 -2462 587800 -2226
rect 587200 -2546 587800 -2462
rect 587200 -2782 587382 -2546
rect 587618 -2782 587800 -2546
rect 587200 -2804 587800 -2782
rect -4816 -3402 -4634 -3166
rect -4398 -3402 -4216 -3166
rect -4816 -3486 -4216 -3402
rect -4816 -3722 -4634 -3486
rect -4398 -3722 -4216 -3486
rect -4816 -3744 -4216 -3722
rect 588140 -3166 588740 707102
rect 588140 -3402 588322 -3166
rect 588558 -3402 588740 -3166
rect 588140 -3486 588740 -3402
rect 588140 -3722 588322 -3486
rect 588558 -3722 588740 -3486
rect 588140 -3744 588740 -3722
rect -5756 -4342 -5574 -4106
rect -5338 -4342 -5156 -4106
rect -5756 -4426 -5156 -4342
rect -5756 -4662 -5574 -4426
rect -5338 -4662 -5156 -4426
rect -5756 -4684 -5156 -4662
rect 589080 -4106 589680 708042
rect 589080 -4342 589262 -4106
rect 589498 -4342 589680 -4106
rect 589080 -4426 589680 -4342
rect 589080 -4662 589262 -4426
rect 589498 -4662 589680 -4426
rect 589080 -4684 589680 -4662
rect -6696 -5282 -6514 -5046
rect -6278 -5282 -6096 -5046
rect -6696 -5366 -6096 -5282
rect -6696 -5602 -6514 -5366
rect -6278 -5602 -6096 -5366
rect -6696 -5624 -6096 -5602
rect 590020 -5046 590620 708982
rect 590020 -5282 590202 -5046
rect 590438 -5282 590620 -5046
rect 590020 -5366 590620 -5282
rect 590020 -5602 590202 -5366
rect 590438 -5602 590620 -5366
rect 590020 -5624 590620 -5602
rect -7636 -6222 -7454 -5986
rect -7218 -6222 -7036 -5986
rect -7636 -6306 -7036 -6222
rect -7636 -6542 -7454 -6306
rect -7218 -6542 -7036 -6306
rect -7636 -6564 -7036 -6542
rect 590960 -5986 591560 709922
rect 590960 -6222 591142 -5986
rect 591378 -6222 591560 -5986
rect 590960 -6306 591560 -6222
rect 590960 -6542 591142 -6306
rect 591378 -6542 591560 -6306
rect 590960 -6564 591560 -6542
rect -8576 -7162 -8394 -6926
rect -8158 -7162 -7976 -6926
rect -8576 -7246 -7976 -7162
rect -8576 -7482 -8394 -7246
rect -8158 -7482 -7976 -7246
rect -8576 -7504 -7976 -7482
rect 591900 -6926 592500 710862
rect 591900 -7162 592082 -6926
rect 592318 -7162 592500 -6926
rect 591900 -7246 592500 -7162
rect 591900 -7482 592082 -7246
rect 592318 -7482 592500 -7246
rect 591900 -7504 592500 -7482
<< via4 >>
rect -8394 711182 -8158 711418
rect -8394 710862 -8158 711098
rect 592082 711182 592318 711418
rect 592082 710862 592318 711098
rect -7454 710242 -7218 710478
rect -7454 709922 -7218 710158
rect 591142 710242 591378 710478
rect 591142 709922 591378 710158
rect -6514 709302 -6278 709538
rect -6514 708982 -6278 709218
rect 590202 709302 590438 709538
rect 590202 708982 590438 709218
rect -5574 708362 -5338 708598
rect -5574 708042 -5338 708278
rect 589262 708362 589498 708598
rect 589262 708042 589498 708278
rect -4634 707422 -4398 707658
rect -4634 707102 -4398 707338
rect 588322 707422 588558 707658
rect 588322 707102 588558 707338
rect -3694 706482 -3458 706718
rect -3694 706162 -3458 706398
rect 587382 706482 587618 706718
rect 587382 706162 587618 706398
rect -2754 705542 -2518 705778
rect -2754 705222 -2518 705458
rect -2754 668218 -2518 668454
rect -2754 667898 -2518 668134
rect -2754 632218 -2518 632454
rect -2754 631898 -2518 632134
rect -2754 596218 -2518 596454
rect -2754 595898 -2518 596134
rect -2754 560218 -2518 560454
rect -2754 559898 -2518 560134
rect -2754 524218 -2518 524454
rect -2754 523898 -2518 524134
rect -2754 488218 -2518 488454
rect -2754 487898 -2518 488134
rect -2754 452218 -2518 452454
rect -2754 451898 -2518 452134
rect -2754 416218 -2518 416454
rect -2754 415898 -2518 416134
rect -2754 380218 -2518 380454
rect -2754 379898 -2518 380134
rect -2754 344218 -2518 344454
rect -2754 343898 -2518 344134
rect -2754 308218 -2518 308454
rect -2754 307898 -2518 308134
rect -2754 272218 -2518 272454
rect -2754 271898 -2518 272134
rect -2754 236218 -2518 236454
rect -2754 235898 -2518 236134
rect -2754 200218 -2518 200454
rect -2754 199898 -2518 200134
rect -2754 164218 -2518 164454
rect -2754 163898 -2518 164134
rect -2754 128218 -2518 128454
rect -2754 127898 -2518 128134
rect -2754 92218 -2518 92454
rect -2754 91898 -2518 92134
rect -2754 56218 -2518 56454
rect -2754 55898 -2518 56134
rect -2754 20218 -2518 20454
rect -2754 19898 -2518 20134
rect -1814 704602 -1578 704838
rect -1814 704282 -1578 704518
rect -1814 686218 -1578 686454
rect -1814 685898 -1578 686134
rect -1814 650218 -1578 650454
rect -1814 649898 -1578 650134
rect -1814 614218 -1578 614454
rect -1814 613898 -1578 614134
rect -1814 578218 -1578 578454
rect -1814 577898 -1578 578134
rect -1814 542218 -1578 542454
rect -1814 541898 -1578 542134
rect -1814 506218 -1578 506454
rect -1814 505898 -1578 506134
rect -1814 470218 -1578 470454
rect -1814 469898 -1578 470134
rect -1814 434218 -1578 434454
rect -1814 433898 -1578 434134
rect -1814 398218 -1578 398454
rect -1814 397898 -1578 398134
rect -1814 362218 -1578 362454
rect -1814 361898 -1578 362134
rect -1814 326218 -1578 326454
rect -1814 325898 -1578 326134
rect -1814 290218 -1578 290454
rect -1814 289898 -1578 290134
rect -1814 254218 -1578 254454
rect -1814 253898 -1578 254134
rect -1814 218218 -1578 218454
rect -1814 217898 -1578 218134
rect -1814 182218 -1578 182454
rect -1814 181898 -1578 182134
rect -1814 146218 -1578 146454
rect -1814 145898 -1578 146134
rect -1814 110218 -1578 110454
rect -1814 109898 -1578 110134
rect -1814 74218 -1578 74454
rect -1814 73898 -1578 74134
rect -1814 38218 -1578 38454
rect -1814 37898 -1578 38134
rect -1814 2218 -1578 2454
rect -1814 1898 -1578 2134
rect -1814 -582 -1578 -346
rect -1814 -902 -1578 -666
rect 986 704602 1222 704838
rect 986 704282 1222 704518
rect 986 686218 1222 686454
rect 986 685898 1222 686134
rect 986 650218 1222 650454
rect 986 649898 1222 650134
rect 986 614218 1222 614454
rect 986 613898 1222 614134
rect 986 578218 1222 578454
rect 986 577898 1222 578134
rect 986 542218 1222 542454
rect 986 541898 1222 542134
rect 986 506218 1222 506454
rect 986 505898 1222 506134
rect 986 470218 1222 470454
rect 986 469898 1222 470134
rect 986 434218 1222 434454
rect 986 433898 1222 434134
rect 986 398218 1222 398454
rect 986 397898 1222 398134
rect 986 362218 1222 362454
rect 986 361898 1222 362134
rect 986 326218 1222 326454
rect 986 325898 1222 326134
rect 986 290218 1222 290454
rect 986 289898 1222 290134
rect 986 254218 1222 254454
rect 986 253898 1222 254134
rect 986 218218 1222 218454
rect 986 217898 1222 218134
rect 986 182218 1222 182454
rect 986 181898 1222 182134
rect 986 146218 1222 146454
rect 986 145898 1222 146134
rect 986 110218 1222 110454
rect 986 109898 1222 110134
rect 986 74218 1222 74454
rect 986 73898 1222 74134
rect 986 38218 1222 38454
rect 986 37898 1222 38134
rect 986 2218 1222 2454
rect 986 1898 1222 2134
rect 986 -582 1222 -346
rect 986 -902 1222 -666
rect -2754 -1522 -2518 -1286
rect -2754 -1842 -2518 -1606
rect 18986 705542 19222 705778
rect 18986 705222 19222 705458
rect 18986 668218 19222 668454
rect 18986 667898 19222 668134
rect 18986 632218 19222 632454
rect 18986 631898 19222 632134
rect 18986 596218 19222 596454
rect 18986 595898 19222 596134
rect 36986 704602 37222 704838
rect 36986 704282 37222 704518
rect 36986 686218 37222 686454
rect 36986 685898 37222 686134
rect 36986 650218 37222 650454
rect 36986 649898 37222 650134
rect 36986 614218 37222 614454
rect 36986 613898 37222 614134
rect 54986 705542 55222 705778
rect 54986 705222 55222 705458
rect 54986 668218 55222 668454
rect 54986 667898 55222 668134
rect 54986 632218 55222 632454
rect 54986 631898 55222 632134
rect 54986 596218 55222 596454
rect 54986 595898 55222 596134
rect 72986 704602 73222 704838
rect 72986 704282 73222 704518
rect 72986 686218 73222 686454
rect 72986 685898 73222 686134
rect 72986 650218 73222 650454
rect 72986 649898 73222 650134
rect 72986 614218 73222 614454
rect 72986 613898 73222 614134
rect 90986 705542 91222 705778
rect 90986 705222 91222 705458
rect 90986 668218 91222 668454
rect 90986 667898 91222 668134
rect 90986 632218 91222 632454
rect 90986 631898 91222 632134
rect 90986 596218 91222 596454
rect 90986 595898 91222 596134
rect 108986 704602 109222 704838
rect 108986 704282 109222 704518
rect 108986 686218 109222 686454
rect 108986 685898 109222 686134
rect 108986 650218 109222 650454
rect 108986 649898 109222 650134
rect 108986 614218 109222 614454
rect 108986 613898 109222 614134
rect 126986 705542 127222 705778
rect 126986 705222 127222 705458
rect 126986 668218 127222 668454
rect 126986 667898 127222 668134
rect 126986 632218 127222 632454
rect 126986 631898 127222 632134
rect 126986 596218 127222 596454
rect 126986 595898 127222 596134
rect 144986 704602 145222 704838
rect 144986 704282 145222 704518
rect 144986 686218 145222 686454
rect 144986 685898 145222 686134
rect 144986 650218 145222 650454
rect 144986 649898 145222 650134
rect 144986 614218 145222 614454
rect 144986 613898 145222 614134
rect 162986 705542 163222 705778
rect 162986 705222 163222 705458
rect 162986 668218 163222 668454
rect 162986 667898 163222 668134
rect 162986 632218 163222 632454
rect 162986 631898 163222 632134
rect 162986 596218 163222 596454
rect 162986 595898 163222 596134
rect 180986 704602 181222 704838
rect 180986 704282 181222 704518
rect 180986 686218 181222 686454
rect 180986 685898 181222 686134
rect 180986 650218 181222 650454
rect 180986 649898 181222 650134
rect 180986 614218 181222 614454
rect 180986 613898 181222 614134
rect 198986 705542 199222 705778
rect 198986 705222 199222 705458
rect 198986 668218 199222 668454
rect 198986 667898 199222 668134
rect 198986 632218 199222 632454
rect 198986 631898 199222 632134
rect 198986 596218 199222 596454
rect 198986 595898 199222 596134
rect 216986 704602 217222 704838
rect 216986 704282 217222 704518
rect 216986 686218 217222 686454
rect 216986 685898 217222 686134
rect 216986 650218 217222 650454
rect 216986 649898 217222 650134
rect 216986 614218 217222 614454
rect 216986 613898 217222 614134
rect 234986 705542 235222 705778
rect 234986 705222 235222 705458
rect 234986 668218 235222 668454
rect 234986 667898 235222 668134
rect 234986 632218 235222 632454
rect 234986 631898 235222 632134
rect 234986 596218 235222 596454
rect 234986 595898 235222 596134
rect 252986 704602 253222 704838
rect 252986 704282 253222 704518
rect 252986 686218 253222 686454
rect 252986 685898 253222 686134
rect 252986 650218 253222 650454
rect 252986 649898 253222 650134
rect 252986 614218 253222 614454
rect 252986 613898 253222 614134
rect 270986 705542 271222 705778
rect 270986 705222 271222 705458
rect 288986 704602 289222 704838
rect 288986 704282 289222 704518
rect 270986 668218 271222 668454
rect 270986 667898 271222 668134
rect 270986 632218 271222 632454
rect 270986 631898 271222 632134
rect 270986 596218 271222 596454
rect 270986 595898 271222 596134
rect 262170 578218 262406 578454
rect 262170 577898 262406 578134
rect 18986 560218 19222 560454
rect 18986 559898 19222 560134
rect 246810 560218 247046 560454
rect 246810 559898 247046 560134
rect 270986 560218 271222 560454
rect 270986 559898 271222 560134
rect 262170 542218 262406 542454
rect 262170 541898 262406 542134
rect 18986 524218 19222 524454
rect 18986 523898 19222 524134
rect 246810 524218 247046 524454
rect 246810 523898 247046 524134
rect 270986 524218 271222 524454
rect 270986 523898 271222 524134
rect 262170 506218 262406 506454
rect 262170 505898 262406 506134
rect 18986 488218 19222 488454
rect 18986 487898 19222 488134
rect 246810 488218 247046 488454
rect 246810 487898 247046 488134
rect 270986 488218 271222 488454
rect 270986 487898 271222 488134
rect 262170 470218 262406 470454
rect 262170 469898 262406 470134
rect 18986 452218 19222 452454
rect 18986 451898 19222 452134
rect 246810 452218 247046 452454
rect 246810 451898 247046 452134
rect 270986 452218 271222 452454
rect 270986 451898 271222 452134
rect 262170 434218 262406 434454
rect 262170 433898 262406 434134
rect 18986 416218 19222 416454
rect 18986 415898 19222 416134
rect 246810 416218 247046 416454
rect 246810 415898 247046 416134
rect 270986 416218 271222 416454
rect 270986 415898 271222 416134
rect 262170 398218 262406 398454
rect 262170 397898 262406 398134
rect 18986 380218 19222 380454
rect 18986 379898 19222 380134
rect 18986 344218 19222 344454
rect 18986 343898 19222 344134
rect 18986 308218 19222 308454
rect 18986 307898 19222 308134
rect 36986 362218 37222 362454
rect 36986 361898 37222 362134
rect 36986 326218 37222 326454
rect 36986 325898 37222 326134
rect 36986 290218 37222 290454
rect 36986 289898 37222 290134
rect 54986 380218 55222 380454
rect 54986 379898 55222 380134
rect 54986 344218 55222 344454
rect 54986 343898 55222 344134
rect 54986 308218 55222 308454
rect 54986 307898 55222 308134
rect 72986 362218 73222 362454
rect 72986 361898 73222 362134
rect 72986 326218 73222 326454
rect 72986 325898 73222 326134
rect 72986 290218 73222 290454
rect 72986 289898 73222 290134
rect 90986 380218 91222 380454
rect 90986 379898 91222 380134
rect 90986 344218 91222 344454
rect 90986 343898 91222 344134
rect 90986 308218 91222 308454
rect 90986 307898 91222 308134
rect 108986 362218 109222 362454
rect 108986 361898 109222 362134
rect 108986 326218 109222 326454
rect 108986 325898 109222 326134
rect 108986 290218 109222 290454
rect 108986 289898 109222 290134
rect 126986 380218 127222 380454
rect 126986 379898 127222 380134
rect 126986 344218 127222 344454
rect 126986 343898 127222 344134
rect 126986 308218 127222 308454
rect 126986 307898 127222 308134
rect 144986 362218 145222 362454
rect 144986 361898 145222 362134
rect 144986 326218 145222 326454
rect 144986 325898 145222 326134
rect 144986 290218 145222 290454
rect 144986 289898 145222 290134
rect 162986 380218 163222 380454
rect 162986 379898 163222 380134
rect 162986 344218 163222 344454
rect 162986 343898 163222 344134
rect 162986 308218 163222 308454
rect 162986 307898 163222 308134
rect 180986 362218 181222 362454
rect 180986 361898 181222 362134
rect 180986 326218 181222 326454
rect 180986 325898 181222 326134
rect 180986 290218 181222 290454
rect 180986 289898 181222 290134
rect 198986 380218 199222 380454
rect 198986 379898 199222 380134
rect 198986 344218 199222 344454
rect 198986 343898 199222 344134
rect 198986 308218 199222 308454
rect 198986 307898 199222 308134
rect 216986 362218 217222 362454
rect 216986 361898 217222 362134
rect 216986 326218 217222 326454
rect 216986 325898 217222 326134
rect 216986 290218 217222 290454
rect 216986 289898 217222 290134
rect 234986 380218 235222 380454
rect 234986 379898 235222 380134
rect 234986 344218 235222 344454
rect 234986 343898 235222 344134
rect 234986 308218 235222 308454
rect 234986 307898 235222 308134
rect 252986 362218 253222 362454
rect 252986 361898 253222 362134
rect 270986 380218 271222 380454
rect 270986 379898 271222 380134
rect 252986 326218 253222 326454
rect 252986 325898 253222 326134
rect 252986 290218 253222 290454
rect 252986 289898 253222 290134
rect 270986 308218 271222 308454
rect 270986 307898 271222 308134
rect 18986 272218 19222 272454
rect 18986 271898 19222 272134
rect 270986 272218 271222 272454
rect 270986 271898 271222 272134
rect 262170 254218 262406 254454
rect 262170 253898 262406 254134
rect 18986 236218 19222 236454
rect 18986 235898 19222 236134
rect 246810 236218 247046 236454
rect 246810 235898 247046 236134
rect 270986 236218 271222 236454
rect 270986 235898 271222 236134
rect 262170 218218 262406 218454
rect 262170 217898 262406 218134
rect 18986 200218 19222 200454
rect 18986 199898 19222 200134
rect 246810 200218 247046 200454
rect 246810 199898 247046 200134
rect 270986 200218 271222 200454
rect 270986 199898 271222 200134
rect 262170 182218 262406 182454
rect 262170 181898 262406 182134
rect 18986 164218 19222 164454
rect 18986 163898 19222 164134
rect 246810 164218 247046 164454
rect 246810 163898 247046 164134
rect 270986 164218 271222 164454
rect 270986 163898 271222 164134
rect 262170 146218 262406 146454
rect 262170 145898 262406 146134
rect 18986 128218 19222 128454
rect 18986 127898 19222 128134
rect 246810 128218 247046 128454
rect 246810 127898 247046 128134
rect 270986 128218 271222 128454
rect 270986 127898 271222 128134
rect 262170 110218 262406 110454
rect 262170 109898 262406 110134
rect 18986 92218 19222 92454
rect 18986 91898 19222 92134
rect 246810 92218 247046 92454
rect 246810 91898 247046 92134
rect 270986 92218 271222 92454
rect 270986 91898 271222 92134
rect 18986 56218 19222 56454
rect 18986 55898 19222 56134
rect 18986 20218 19222 20454
rect 18986 19898 19222 20134
rect 18986 -1522 19222 -1286
rect 18986 -1842 19222 -1606
rect 36986 38218 37222 38454
rect 36986 37898 37222 38134
rect 36986 2218 37222 2454
rect 36986 1898 37222 2134
rect 36986 -582 37222 -346
rect 36986 -902 37222 -666
rect 54986 56218 55222 56454
rect 54986 55898 55222 56134
rect 54986 20218 55222 20454
rect 54986 19898 55222 20134
rect 54986 -1522 55222 -1286
rect 54986 -1842 55222 -1606
rect 72986 38218 73222 38454
rect 72986 37898 73222 38134
rect 72986 2218 73222 2454
rect 72986 1898 73222 2134
rect 72986 -582 73222 -346
rect 72986 -902 73222 -666
rect 90986 56218 91222 56454
rect 90986 55898 91222 56134
rect 90986 20218 91222 20454
rect 90986 19898 91222 20134
rect 90986 -1522 91222 -1286
rect 90986 -1842 91222 -1606
rect 108986 38218 109222 38454
rect 108986 37898 109222 38134
rect 108986 2218 109222 2454
rect 108986 1898 109222 2134
rect 108986 -582 109222 -346
rect 108986 -902 109222 -666
rect 126986 56218 127222 56454
rect 126986 55898 127222 56134
rect 126986 20218 127222 20454
rect 126986 19898 127222 20134
rect 126986 -1522 127222 -1286
rect 126986 -1842 127222 -1606
rect 144986 38218 145222 38454
rect 144986 37898 145222 38134
rect 144986 2218 145222 2454
rect 144986 1898 145222 2134
rect 144986 -582 145222 -346
rect 144986 -902 145222 -666
rect 162986 56218 163222 56454
rect 162986 55898 163222 56134
rect 162986 20218 163222 20454
rect 162986 19898 163222 20134
rect 162986 -1522 163222 -1286
rect 162986 -1842 163222 -1606
rect 180986 38218 181222 38454
rect 180986 37898 181222 38134
rect 180986 2218 181222 2454
rect 180986 1898 181222 2134
rect 180986 -582 181222 -346
rect 180986 -902 181222 -666
rect 198986 56218 199222 56454
rect 198986 55898 199222 56134
rect 198986 20218 199222 20454
rect 198986 19898 199222 20134
rect 198986 -1522 199222 -1286
rect 198986 -1842 199222 -1606
rect 216986 38218 217222 38454
rect 216986 37898 217222 38134
rect 216986 2218 217222 2454
rect 216986 1898 217222 2134
rect 216986 -582 217222 -346
rect 216986 -902 217222 -666
rect 234986 56218 235222 56454
rect 234986 55898 235222 56134
rect 234986 20218 235222 20454
rect 234986 19898 235222 20134
rect 234986 -1522 235222 -1286
rect 234986 -1842 235222 -1606
rect 252986 38218 253222 38454
rect 252986 37898 253222 38134
rect 252986 2218 253222 2454
rect 252986 1898 253222 2134
rect 252986 -582 253222 -346
rect 252986 -902 253222 -666
rect 306986 705542 307222 705778
rect 306986 705222 307222 705458
rect 288986 686218 289222 686454
rect 288986 685898 289222 686134
rect 288986 650218 289222 650454
rect 288986 649898 289222 650134
rect 288986 614218 289222 614454
rect 288986 613898 289222 614134
rect 288986 578218 289222 578454
rect 288986 577898 289222 578134
rect 288986 542218 289222 542454
rect 288986 541898 289222 542134
rect 288986 506218 289222 506454
rect 288986 505898 289222 506134
rect 288986 470218 289222 470454
rect 288986 469898 289222 470134
rect 288986 434218 289222 434454
rect 288986 433898 289222 434134
rect 288986 398218 289222 398454
rect 288986 397898 289222 398134
rect 288986 362218 289222 362454
rect 288986 361898 289222 362134
rect 292154 344218 292390 344454
rect 292154 343898 292390 344134
rect 288986 290218 289222 290454
rect 288986 289898 289222 290134
rect 288986 254218 289222 254454
rect 288986 253898 289222 254134
rect 288986 218218 289222 218454
rect 288986 217898 289222 218134
rect 288986 182218 289222 182454
rect 288986 181898 289222 182134
rect 288986 146218 289222 146454
rect 288986 145898 289222 146134
rect 288986 110218 289222 110454
rect 288986 109898 289222 110134
rect 288986 74218 289222 74454
rect 288986 73898 289222 74134
rect 270986 56218 271222 56454
rect 270986 55898 271222 56134
rect 270986 20218 271222 20454
rect 270986 19898 271222 20134
rect 270986 -1522 271222 -1286
rect 270986 -1842 271222 -1606
rect 288986 38218 289222 38454
rect 288986 37898 289222 38134
rect 306986 668218 307222 668454
rect 306986 667898 307222 668134
rect 306986 632218 307222 632454
rect 306986 631898 307222 632134
rect 324986 704602 325222 704838
rect 324986 704282 325222 704518
rect 324986 686218 325222 686454
rect 324986 685898 325222 686134
rect 324986 650218 325222 650454
rect 324986 649898 325222 650134
rect 324986 614218 325222 614454
rect 324986 613898 325222 614134
rect 306986 596218 307222 596454
rect 306986 595898 307222 596134
rect 306986 560218 307222 560454
rect 306986 559898 307222 560134
rect 306986 524218 307222 524454
rect 306986 523898 307222 524134
rect 306986 488218 307222 488454
rect 306986 487898 307222 488134
rect 306986 452218 307222 452454
rect 306986 451898 307222 452134
rect 306986 416218 307222 416454
rect 306986 415898 307222 416134
rect 306986 380218 307222 380454
rect 306986 379898 307222 380134
rect 342986 705542 343222 705778
rect 342986 705222 343222 705458
rect 342986 668218 343222 668454
rect 342986 667898 343222 668134
rect 342986 632218 343222 632454
rect 342986 631898 343222 632134
rect 342986 596218 343222 596454
rect 342986 595898 343222 596134
rect 360986 704602 361222 704838
rect 360986 704282 361222 704518
rect 360986 686218 361222 686454
rect 360986 685898 361222 686134
rect 360986 650218 361222 650454
rect 360986 649898 361222 650134
rect 360986 614218 361222 614454
rect 360986 613898 361222 614134
rect 378986 705542 379222 705778
rect 378986 705222 379222 705458
rect 378986 668218 379222 668454
rect 378986 667898 379222 668134
rect 378986 632218 379222 632454
rect 378986 631898 379222 632134
rect 378986 596218 379222 596454
rect 378986 595898 379222 596134
rect 396986 704602 397222 704838
rect 396986 704282 397222 704518
rect 396986 686218 397222 686454
rect 396986 685898 397222 686134
rect 396986 650218 397222 650454
rect 396986 649898 397222 650134
rect 396986 614218 397222 614454
rect 396986 613898 397222 614134
rect 414986 705542 415222 705778
rect 414986 705222 415222 705458
rect 414986 668218 415222 668454
rect 414986 667898 415222 668134
rect 414986 632218 415222 632454
rect 414986 631898 415222 632134
rect 414986 596218 415222 596454
rect 414986 595898 415222 596134
rect 432986 704602 433222 704838
rect 432986 704282 433222 704518
rect 432986 686218 433222 686454
rect 432986 685898 433222 686134
rect 432986 650218 433222 650454
rect 432986 649898 433222 650134
rect 432986 614218 433222 614454
rect 432986 613898 433222 614134
rect 450986 705542 451222 705778
rect 450986 705222 451222 705458
rect 450986 668218 451222 668454
rect 450986 667898 451222 668134
rect 450986 632218 451222 632454
rect 450986 631898 451222 632134
rect 450986 596218 451222 596454
rect 450986 595898 451222 596134
rect 468986 704602 469222 704838
rect 468986 704282 469222 704518
rect 468986 686218 469222 686454
rect 468986 685898 469222 686134
rect 468986 650218 469222 650454
rect 468986 649898 469222 650134
rect 468986 614218 469222 614454
rect 468986 613898 469222 614134
rect 486986 705542 487222 705778
rect 486986 705222 487222 705458
rect 486986 668218 487222 668454
rect 486986 667898 487222 668134
rect 486986 632218 487222 632454
rect 486986 631898 487222 632134
rect 486986 596218 487222 596454
rect 486986 595898 487222 596134
rect 504986 704602 505222 704838
rect 504986 704282 505222 704518
rect 504986 686218 505222 686454
rect 504986 685898 505222 686134
rect 504986 650218 505222 650454
rect 504986 649898 505222 650134
rect 504986 614218 505222 614454
rect 504986 613898 505222 614134
rect 522986 705542 523222 705778
rect 522986 705222 523222 705458
rect 522986 668218 523222 668454
rect 522986 667898 523222 668134
rect 522986 632218 523222 632454
rect 522986 631898 523222 632134
rect 522986 596218 523222 596454
rect 522986 595898 523222 596134
rect 540986 704602 541222 704838
rect 540986 704282 541222 704518
rect 540986 686218 541222 686454
rect 540986 685898 541222 686134
rect 540986 650218 541222 650454
rect 540986 649898 541222 650134
rect 540986 614218 541222 614454
rect 540986 613898 541222 614134
rect 558986 705542 559222 705778
rect 558986 705222 559222 705458
rect 558986 668218 559222 668454
rect 558986 667898 559222 668134
rect 558986 632218 559222 632454
rect 558986 631898 559222 632134
rect 558986 596218 559222 596454
rect 558986 595898 559222 596134
rect 586442 705542 586678 705778
rect 586442 705222 586678 705458
rect 576986 704602 577222 704838
rect 576986 704282 577222 704518
rect 576986 686218 577222 686454
rect 576986 685898 577222 686134
rect 576986 650218 577222 650454
rect 576986 649898 577222 650134
rect 576986 614218 577222 614454
rect 576986 613898 577222 614134
rect 554298 578218 554534 578454
rect 554298 577898 554534 578134
rect 576986 578218 577222 578454
rect 576986 577898 577222 578134
rect 538938 560218 539174 560454
rect 538938 559898 539174 560134
rect 554298 542218 554534 542454
rect 554298 541898 554534 542134
rect 576986 542218 577222 542454
rect 576986 541898 577222 542134
rect 538938 524218 539174 524454
rect 538938 523898 539174 524134
rect 554298 506218 554534 506454
rect 554298 505898 554534 506134
rect 576986 506218 577222 506454
rect 576986 505898 577222 506134
rect 538938 488218 539174 488454
rect 538938 487898 539174 488134
rect 554298 470218 554534 470454
rect 554298 469898 554534 470134
rect 576986 470218 577222 470454
rect 576986 469898 577222 470134
rect 538938 452218 539174 452454
rect 538938 451898 539174 452134
rect 554298 434218 554534 434454
rect 554298 433898 554534 434134
rect 576986 434218 577222 434454
rect 576986 433898 577222 434134
rect 538938 416218 539174 416454
rect 538938 415898 539174 416134
rect 554298 398218 554534 398454
rect 554298 397898 554534 398134
rect 576986 398218 577222 398454
rect 576986 397898 577222 398134
rect 324986 362218 325222 362454
rect 324986 361898 325222 362134
rect 307514 326218 307750 326454
rect 307514 325898 307750 326134
rect 324986 326218 325222 326454
rect 324986 325898 325222 326134
rect 306986 308218 307222 308454
rect 306986 307898 307222 308134
rect 324986 290218 325222 290454
rect 324986 289898 325222 290134
rect 342986 380218 343222 380454
rect 342986 379898 343222 380134
rect 342986 344218 343222 344454
rect 342986 343898 343222 344134
rect 342986 308218 343222 308454
rect 342986 307898 343222 308134
rect 360986 362218 361222 362454
rect 360986 361898 361222 362134
rect 360986 326218 361222 326454
rect 360986 325898 361222 326134
rect 360986 290218 361222 290454
rect 360986 289898 361222 290134
rect 378986 380218 379222 380454
rect 378986 379898 379222 380134
rect 378986 344218 379222 344454
rect 378986 343898 379222 344134
rect 378986 308218 379222 308454
rect 378986 307898 379222 308134
rect 396986 362218 397222 362454
rect 396986 361898 397222 362134
rect 396986 326218 397222 326454
rect 396986 325898 397222 326134
rect 396986 290218 397222 290454
rect 396986 289898 397222 290134
rect 414986 380218 415222 380454
rect 414986 379898 415222 380134
rect 414986 344218 415222 344454
rect 414986 343898 415222 344134
rect 414986 308218 415222 308454
rect 414986 307898 415222 308134
rect 432986 362218 433222 362454
rect 432986 361898 433222 362134
rect 432986 326218 433222 326454
rect 432986 325898 433222 326134
rect 432986 290218 433222 290454
rect 432986 289898 433222 290134
rect 450986 380218 451222 380454
rect 450986 379898 451222 380134
rect 450986 344218 451222 344454
rect 450986 343898 451222 344134
rect 450986 308218 451222 308454
rect 450986 307898 451222 308134
rect 468986 362218 469222 362454
rect 468986 361898 469222 362134
rect 468986 326218 469222 326454
rect 468986 325898 469222 326134
rect 468986 290218 469222 290454
rect 468986 289898 469222 290134
rect 486986 380218 487222 380454
rect 486986 379898 487222 380134
rect 486986 344218 487222 344454
rect 486986 343898 487222 344134
rect 486986 308218 487222 308454
rect 486986 307898 487222 308134
rect 504986 362218 505222 362454
rect 504986 361898 505222 362134
rect 504986 326218 505222 326454
rect 504986 325898 505222 326134
rect 504986 290218 505222 290454
rect 504986 289898 505222 290134
rect 522986 380218 523222 380454
rect 522986 379898 523222 380134
rect 522986 344218 523222 344454
rect 522986 343898 523222 344134
rect 522986 308218 523222 308454
rect 522986 307898 523222 308134
rect 540986 362218 541222 362454
rect 540986 361898 541222 362134
rect 540986 326218 541222 326454
rect 540986 325898 541222 326134
rect 540986 290218 541222 290454
rect 540986 289898 541222 290134
rect 558986 380218 559222 380454
rect 558986 379898 559222 380134
rect 558986 344218 559222 344454
rect 558986 343898 559222 344134
rect 558986 308218 559222 308454
rect 558986 307898 559222 308134
rect 576986 362218 577222 362454
rect 576986 361898 577222 362134
rect 576986 326218 577222 326454
rect 576986 325898 577222 326134
rect 576986 290218 577222 290454
rect 576986 289898 577222 290134
rect 306986 272218 307222 272454
rect 306986 271898 307222 272134
rect 554298 254218 554534 254454
rect 554298 253898 554534 254134
rect 576986 254218 577222 254454
rect 576986 253898 577222 254134
rect 306986 236218 307222 236454
rect 306986 235898 307222 236134
rect 538938 236218 539174 236454
rect 538938 235898 539174 236134
rect 554298 218218 554534 218454
rect 554298 217898 554534 218134
rect 576986 218218 577222 218454
rect 576986 217898 577222 218134
rect 306986 200218 307222 200454
rect 306986 199898 307222 200134
rect 538938 200218 539174 200454
rect 538938 199898 539174 200134
rect 554298 182218 554534 182454
rect 554298 181898 554534 182134
rect 576986 182218 577222 182454
rect 576986 181898 577222 182134
rect 306986 164218 307222 164454
rect 306986 163898 307222 164134
rect 538938 164218 539174 164454
rect 538938 163898 539174 164134
rect 554298 146218 554534 146454
rect 554298 145898 554534 146134
rect 576986 146218 577222 146454
rect 576986 145898 577222 146134
rect 306986 128218 307222 128454
rect 306986 127898 307222 128134
rect 538938 128218 539174 128454
rect 538938 127898 539174 128134
rect 554298 110218 554534 110454
rect 554298 109898 554534 110134
rect 576986 110218 577222 110454
rect 576986 109898 577222 110134
rect 306986 92218 307222 92454
rect 306986 91898 307222 92134
rect 538938 92218 539174 92454
rect 538938 91898 539174 92134
rect 576986 74218 577222 74454
rect 576986 73898 577222 74134
rect 306986 56218 307222 56454
rect 306986 55898 307222 56134
rect 306986 20218 307222 20454
rect 306986 19898 307222 20134
rect 288986 2218 289222 2454
rect 288986 1898 289222 2134
rect 288986 -582 289222 -346
rect 288986 -902 289222 -666
rect 306986 -1522 307222 -1286
rect 306986 -1842 307222 -1606
rect 324986 38218 325222 38454
rect 324986 37898 325222 38134
rect 324986 2218 325222 2454
rect 324986 1898 325222 2134
rect 324986 -582 325222 -346
rect 324986 -902 325222 -666
rect 342986 56218 343222 56454
rect 342986 55898 343222 56134
rect 342986 20218 343222 20454
rect 342986 19898 343222 20134
rect 342986 -1522 343222 -1286
rect 342986 -1842 343222 -1606
rect 360986 38218 361222 38454
rect 360986 37898 361222 38134
rect 360986 2218 361222 2454
rect 360986 1898 361222 2134
rect 360986 -582 361222 -346
rect 360986 -902 361222 -666
rect 378986 56218 379222 56454
rect 378986 55898 379222 56134
rect 378986 20218 379222 20454
rect 378986 19898 379222 20134
rect 378986 -1522 379222 -1286
rect 378986 -1842 379222 -1606
rect 396986 38218 397222 38454
rect 396986 37898 397222 38134
rect 396986 2218 397222 2454
rect 396986 1898 397222 2134
rect 396986 -582 397222 -346
rect 396986 -902 397222 -666
rect 414986 56218 415222 56454
rect 414986 55898 415222 56134
rect 414986 20218 415222 20454
rect 414986 19898 415222 20134
rect 414986 -1522 415222 -1286
rect 414986 -1842 415222 -1606
rect 432986 38218 433222 38454
rect 432986 37898 433222 38134
rect 432986 2218 433222 2454
rect 432986 1898 433222 2134
rect 432986 -582 433222 -346
rect 432986 -902 433222 -666
rect 450986 56218 451222 56454
rect 450986 55898 451222 56134
rect 450986 20218 451222 20454
rect 450986 19898 451222 20134
rect 450986 -1522 451222 -1286
rect 450986 -1842 451222 -1606
rect 468986 38218 469222 38454
rect 468986 37898 469222 38134
rect 468986 2218 469222 2454
rect 468986 1898 469222 2134
rect 468986 -582 469222 -346
rect 468986 -902 469222 -666
rect 486986 56218 487222 56454
rect 486986 55898 487222 56134
rect 486986 20218 487222 20454
rect 486986 19898 487222 20134
rect 486986 -1522 487222 -1286
rect 486986 -1842 487222 -1606
rect 504986 38218 505222 38454
rect 504986 37898 505222 38134
rect 504986 2218 505222 2454
rect 504986 1898 505222 2134
rect 504986 -582 505222 -346
rect 504986 -902 505222 -666
rect 522986 56218 523222 56454
rect 522986 55898 523222 56134
rect 522986 20218 523222 20454
rect 522986 19898 523222 20134
rect 522986 -1522 523222 -1286
rect 522986 -1842 523222 -1606
rect 540986 38218 541222 38454
rect 540986 37898 541222 38134
rect 540986 2218 541222 2454
rect 540986 1898 541222 2134
rect 540986 -582 541222 -346
rect 540986 -902 541222 -666
rect 558986 56218 559222 56454
rect 558986 55898 559222 56134
rect 558986 20218 559222 20454
rect 558986 19898 559222 20134
rect 558986 -1522 559222 -1286
rect 558986 -1842 559222 -1606
rect 576986 38218 577222 38454
rect 576986 37898 577222 38134
rect 576986 2218 577222 2454
rect 576986 1898 577222 2134
rect 576986 -582 577222 -346
rect 576986 -902 577222 -666
rect 585502 704602 585738 704838
rect 585502 704282 585738 704518
rect 585502 686218 585738 686454
rect 585502 685898 585738 686134
rect 585502 650218 585738 650454
rect 585502 649898 585738 650134
rect 585502 614218 585738 614454
rect 585502 613898 585738 614134
rect 585502 578218 585738 578454
rect 585502 577898 585738 578134
rect 585502 542218 585738 542454
rect 585502 541898 585738 542134
rect 585502 506218 585738 506454
rect 585502 505898 585738 506134
rect 585502 470218 585738 470454
rect 585502 469898 585738 470134
rect 585502 434218 585738 434454
rect 585502 433898 585738 434134
rect 585502 398218 585738 398454
rect 585502 397898 585738 398134
rect 585502 362218 585738 362454
rect 585502 361898 585738 362134
rect 585502 326218 585738 326454
rect 585502 325898 585738 326134
rect 585502 290218 585738 290454
rect 585502 289898 585738 290134
rect 585502 254218 585738 254454
rect 585502 253898 585738 254134
rect 585502 218218 585738 218454
rect 585502 217898 585738 218134
rect 585502 182218 585738 182454
rect 585502 181898 585738 182134
rect 585502 146218 585738 146454
rect 585502 145898 585738 146134
rect 585502 110218 585738 110454
rect 585502 109898 585738 110134
rect 585502 74218 585738 74454
rect 585502 73898 585738 74134
rect 585502 38218 585738 38454
rect 585502 37898 585738 38134
rect 585502 2218 585738 2454
rect 585502 1898 585738 2134
rect 585502 -582 585738 -346
rect 585502 -902 585738 -666
rect 586442 668218 586678 668454
rect 586442 667898 586678 668134
rect 586442 632218 586678 632454
rect 586442 631898 586678 632134
rect 586442 596218 586678 596454
rect 586442 595898 586678 596134
rect 586442 560218 586678 560454
rect 586442 559898 586678 560134
rect 586442 524218 586678 524454
rect 586442 523898 586678 524134
rect 586442 488218 586678 488454
rect 586442 487898 586678 488134
rect 586442 452218 586678 452454
rect 586442 451898 586678 452134
rect 586442 416218 586678 416454
rect 586442 415898 586678 416134
rect 586442 380218 586678 380454
rect 586442 379898 586678 380134
rect 586442 344218 586678 344454
rect 586442 343898 586678 344134
rect 586442 308218 586678 308454
rect 586442 307898 586678 308134
rect 586442 272218 586678 272454
rect 586442 271898 586678 272134
rect 586442 236218 586678 236454
rect 586442 235898 586678 236134
rect 586442 200218 586678 200454
rect 586442 199898 586678 200134
rect 586442 164218 586678 164454
rect 586442 163898 586678 164134
rect 586442 128218 586678 128454
rect 586442 127898 586678 128134
rect 586442 92218 586678 92454
rect 586442 91898 586678 92134
rect 586442 56218 586678 56454
rect 586442 55898 586678 56134
rect 586442 20218 586678 20454
rect 586442 19898 586678 20134
rect 586442 -1522 586678 -1286
rect 586442 -1842 586678 -1606
rect -3694 -2462 -3458 -2226
rect -3694 -2782 -3458 -2546
rect 587382 -2462 587618 -2226
rect 587382 -2782 587618 -2546
rect -4634 -3402 -4398 -3166
rect -4634 -3722 -4398 -3486
rect 588322 -3402 588558 -3166
rect 588322 -3722 588558 -3486
rect -5574 -4342 -5338 -4106
rect -5574 -4662 -5338 -4426
rect 589262 -4342 589498 -4106
rect 589262 -4662 589498 -4426
rect -6514 -5282 -6278 -5046
rect -6514 -5602 -6278 -5366
rect 590202 -5282 590438 -5046
rect 590202 -5602 590438 -5366
rect -7454 -6222 -7218 -5986
rect -7454 -6542 -7218 -6306
rect 591142 -6222 591378 -5986
rect 591142 -6542 591378 -6306
rect -8394 -7162 -8158 -6926
rect -8394 -7482 -8158 -7246
rect 592082 -7162 592318 -6926
rect 592082 -7482 592318 -7246
<< metal5 >>
rect -8576 711440 -7976 711442
rect 591900 711440 592500 711442
rect -8576 711418 592500 711440
rect -8576 711182 -8394 711418
rect -8158 711182 592082 711418
rect 592318 711182 592500 711418
rect -8576 711098 592500 711182
rect -8576 710862 -8394 711098
rect -8158 710862 592082 711098
rect 592318 710862 592500 711098
rect -8576 710840 592500 710862
rect -8576 710838 -7976 710840
rect 591900 710838 592500 710840
rect -7636 710500 -7036 710502
rect 590960 710500 591560 710502
rect -7636 710478 591560 710500
rect -7636 710242 -7454 710478
rect -7218 710242 591142 710478
rect 591378 710242 591560 710478
rect -7636 710158 591560 710242
rect -7636 709922 -7454 710158
rect -7218 709922 591142 710158
rect 591378 709922 591560 710158
rect -7636 709900 591560 709922
rect -7636 709898 -7036 709900
rect 590960 709898 591560 709900
rect -6696 709560 -6096 709562
rect 590020 709560 590620 709562
rect -6696 709538 590620 709560
rect -6696 709302 -6514 709538
rect -6278 709302 590202 709538
rect 590438 709302 590620 709538
rect -6696 709218 590620 709302
rect -6696 708982 -6514 709218
rect -6278 708982 590202 709218
rect 590438 708982 590620 709218
rect -6696 708960 590620 708982
rect -6696 708958 -6096 708960
rect 590020 708958 590620 708960
rect -5756 708620 -5156 708622
rect 589080 708620 589680 708622
rect -5756 708598 589680 708620
rect -5756 708362 -5574 708598
rect -5338 708362 589262 708598
rect 589498 708362 589680 708598
rect -5756 708278 589680 708362
rect -5756 708042 -5574 708278
rect -5338 708042 589262 708278
rect 589498 708042 589680 708278
rect -5756 708020 589680 708042
rect -5756 708018 -5156 708020
rect 589080 708018 589680 708020
rect -4816 707680 -4216 707682
rect 588140 707680 588740 707682
rect -4816 707658 588740 707680
rect -4816 707422 -4634 707658
rect -4398 707422 588322 707658
rect 588558 707422 588740 707658
rect -4816 707338 588740 707422
rect -4816 707102 -4634 707338
rect -4398 707102 588322 707338
rect 588558 707102 588740 707338
rect -4816 707080 588740 707102
rect -4816 707078 -4216 707080
rect 588140 707078 588740 707080
rect -3876 706740 -3276 706742
rect 587200 706740 587800 706742
rect -3876 706718 587800 706740
rect -3876 706482 -3694 706718
rect -3458 706482 587382 706718
rect 587618 706482 587800 706718
rect -3876 706398 587800 706482
rect -3876 706162 -3694 706398
rect -3458 706162 587382 706398
rect 587618 706162 587800 706398
rect -3876 706140 587800 706162
rect -3876 706138 -3276 706140
rect 587200 706138 587800 706140
rect -2936 705800 -2336 705802
rect 18804 705800 19404 705802
rect 54804 705800 55404 705802
rect 90804 705800 91404 705802
rect 126804 705800 127404 705802
rect 162804 705800 163404 705802
rect 198804 705800 199404 705802
rect 234804 705800 235404 705802
rect 270804 705800 271404 705802
rect 306804 705800 307404 705802
rect 342804 705800 343404 705802
rect 378804 705800 379404 705802
rect 414804 705800 415404 705802
rect 450804 705800 451404 705802
rect 486804 705800 487404 705802
rect 522804 705800 523404 705802
rect 558804 705800 559404 705802
rect 586260 705800 586860 705802
rect -2936 705778 586860 705800
rect -2936 705542 -2754 705778
rect -2518 705542 18986 705778
rect 19222 705542 54986 705778
rect 55222 705542 90986 705778
rect 91222 705542 126986 705778
rect 127222 705542 162986 705778
rect 163222 705542 198986 705778
rect 199222 705542 234986 705778
rect 235222 705542 270986 705778
rect 271222 705542 306986 705778
rect 307222 705542 342986 705778
rect 343222 705542 378986 705778
rect 379222 705542 414986 705778
rect 415222 705542 450986 705778
rect 451222 705542 486986 705778
rect 487222 705542 522986 705778
rect 523222 705542 558986 705778
rect 559222 705542 586442 705778
rect 586678 705542 586860 705778
rect -2936 705458 586860 705542
rect -2936 705222 -2754 705458
rect -2518 705222 18986 705458
rect 19222 705222 54986 705458
rect 55222 705222 90986 705458
rect 91222 705222 126986 705458
rect 127222 705222 162986 705458
rect 163222 705222 198986 705458
rect 199222 705222 234986 705458
rect 235222 705222 270986 705458
rect 271222 705222 306986 705458
rect 307222 705222 342986 705458
rect 343222 705222 378986 705458
rect 379222 705222 414986 705458
rect 415222 705222 450986 705458
rect 451222 705222 486986 705458
rect 487222 705222 522986 705458
rect 523222 705222 558986 705458
rect 559222 705222 586442 705458
rect 586678 705222 586860 705458
rect -2936 705200 586860 705222
rect -2936 705198 -2336 705200
rect 18804 705198 19404 705200
rect 54804 705198 55404 705200
rect 90804 705198 91404 705200
rect 126804 705198 127404 705200
rect 162804 705198 163404 705200
rect 198804 705198 199404 705200
rect 234804 705198 235404 705200
rect 270804 705198 271404 705200
rect 306804 705198 307404 705200
rect 342804 705198 343404 705200
rect 378804 705198 379404 705200
rect 414804 705198 415404 705200
rect 450804 705198 451404 705200
rect 486804 705198 487404 705200
rect 522804 705198 523404 705200
rect 558804 705198 559404 705200
rect 586260 705198 586860 705200
rect -1996 704860 -1396 704862
rect 804 704860 1404 704862
rect 36804 704860 37404 704862
rect 72804 704860 73404 704862
rect 108804 704860 109404 704862
rect 144804 704860 145404 704862
rect 180804 704860 181404 704862
rect 216804 704860 217404 704862
rect 252804 704860 253404 704862
rect 288804 704860 289404 704862
rect 324804 704860 325404 704862
rect 360804 704860 361404 704862
rect 396804 704860 397404 704862
rect 432804 704860 433404 704862
rect 468804 704860 469404 704862
rect 504804 704860 505404 704862
rect 540804 704860 541404 704862
rect 576804 704860 577404 704862
rect 585320 704860 585920 704862
rect -1996 704838 585920 704860
rect -1996 704602 -1814 704838
rect -1578 704602 986 704838
rect 1222 704602 36986 704838
rect 37222 704602 72986 704838
rect 73222 704602 108986 704838
rect 109222 704602 144986 704838
rect 145222 704602 180986 704838
rect 181222 704602 216986 704838
rect 217222 704602 252986 704838
rect 253222 704602 288986 704838
rect 289222 704602 324986 704838
rect 325222 704602 360986 704838
rect 361222 704602 396986 704838
rect 397222 704602 432986 704838
rect 433222 704602 468986 704838
rect 469222 704602 504986 704838
rect 505222 704602 540986 704838
rect 541222 704602 576986 704838
rect 577222 704602 585502 704838
rect 585738 704602 585920 704838
rect -1996 704518 585920 704602
rect -1996 704282 -1814 704518
rect -1578 704282 986 704518
rect 1222 704282 36986 704518
rect 37222 704282 72986 704518
rect 73222 704282 108986 704518
rect 109222 704282 144986 704518
rect 145222 704282 180986 704518
rect 181222 704282 216986 704518
rect 217222 704282 252986 704518
rect 253222 704282 288986 704518
rect 289222 704282 324986 704518
rect 325222 704282 360986 704518
rect 361222 704282 396986 704518
rect 397222 704282 432986 704518
rect 433222 704282 468986 704518
rect 469222 704282 504986 704518
rect 505222 704282 540986 704518
rect 541222 704282 576986 704518
rect 577222 704282 585502 704518
rect 585738 704282 585920 704518
rect -1996 704260 585920 704282
rect -1996 704258 -1396 704260
rect 804 704258 1404 704260
rect 36804 704258 37404 704260
rect 72804 704258 73404 704260
rect 108804 704258 109404 704260
rect 144804 704258 145404 704260
rect 180804 704258 181404 704260
rect 216804 704258 217404 704260
rect 252804 704258 253404 704260
rect 288804 704258 289404 704260
rect 324804 704258 325404 704260
rect 360804 704258 361404 704260
rect 396804 704258 397404 704260
rect 432804 704258 433404 704260
rect 468804 704258 469404 704260
rect 504804 704258 505404 704260
rect 540804 704258 541404 704260
rect 576804 704258 577404 704260
rect 585320 704258 585920 704260
rect -1996 686476 -1396 686478
rect 804 686476 1404 686478
rect 36804 686476 37404 686478
rect 72804 686476 73404 686478
rect 108804 686476 109404 686478
rect 144804 686476 145404 686478
rect 180804 686476 181404 686478
rect 216804 686476 217404 686478
rect 252804 686476 253404 686478
rect 288804 686476 289404 686478
rect 324804 686476 325404 686478
rect 360804 686476 361404 686478
rect 396804 686476 397404 686478
rect 432804 686476 433404 686478
rect 468804 686476 469404 686478
rect 504804 686476 505404 686478
rect 540804 686476 541404 686478
rect 576804 686476 577404 686478
rect 585320 686476 585920 686478
rect -2936 686454 586860 686476
rect -2936 686218 -1814 686454
rect -1578 686218 986 686454
rect 1222 686218 36986 686454
rect 37222 686218 72986 686454
rect 73222 686218 108986 686454
rect 109222 686218 144986 686454
rect 145222 686218 180986 686454
rect 181222 686218 216986 686454
rect 217222 686218 252986 686454
rect 253222 686218 288986 686454
rect 289222 686218 324986 686454
rect 325222 686218 360986 686454
rect 361222 686218 396986 686454
rect 397222 686218 432986 686454
rect 433222 686218 468986 686454
rect 469222 686218 504986 686454
rect 505222 686218 540986 686454
rect 541222 686218 576986 686454
rect 577222 686218 585502 686454
rect 585738 686218 586860 686454
rect -2936 686134 586860 686218
rect -2936 685898 -1814 686134
rect -1578 685898 986 686134
rect 1222 685898 36986 686134
rect 37222 685898 72986 686134
rect 73222 685898 108986 686134
rect 109222 685898 144986 686134
rect 145222 685898 180986 686134
rect 181222 685898 216986 686134
rect 217222 685898 252986 686134
rect 253222 685898 288986 686134
rect 289222 685898 324986 686134
rect 325222 685898 360986 686134
rect 361222 685898 396986 686134
rect 397222 685898 432986 686134
rect 433222 685898 468986 686134
rect 469222 685898 504986 686134
rect 505222 685898 540986 686134
rect 541222 685898 576986 686134
rect 577222 685898 585502 686134
rect 585738 685898 586860 686134
rect -2936 685876 586860 685898
rect -1996 685874 -1396 685876
rect 804 685874 1404 685876
rect 36804 685874 37404 685876
rect 72804 685874 73404 685876
rect 108804 685874 109404 685876
rect 144804 685874 145404 685876
rect 180804 685874 181404 685876
rect 216804 685874 217404 685876
rect 252804 685874 253404 685876
rect 288804 685874 289404 685876
rect 324804 685874 325404 685876
rect 360804 685874 361404 685876
rect 396804 685874 397404 685876
rect 432804 685874 433404 685876
rect 468804 685874 469404 685876
rect 504804 685874 505404 685876
rect 540804 685874 541404 685876
rect 576804 685874 577404 685876
rect 585320 685874 585920 685876
rect -2936 668476 -2336 668478
rect 18804 668476 19404 668478
rect 54804 668476 55404 668478
rect 90804 668476 91404 668478
rect 126804 668476 127404 668478
rect 162804 668476 163404 668478
rect 198804 668476 199404 668478
rect 234804 668476 235404 668478
rect 270804 668476 271404 668478
rect 306804 668476 307404 668478
rect 342804 668476 343404 668478
rect 378804 668476 379404 668478
rect 414804 668476 415404 668478
rect 450804 668476 451404 668478
rect 486804 668476 487404 668478
rect 522804 668476 523404 668478
rect 558804 668476 559404 668478
rect 586260 668476 586860 668478
rect -2936 668454 586860 668476
rect -2936 668218 -2754 668454
rect -2518 668218 18986 668454
rect 19222 668218 54986 668454
rect 55222 668218 90986 668454
rect 91222 668218 126986 668454
rect 127222 668218 162986 668454
rect 163222 668218 198986 668454
rect 199222 668218 234986 668454
rect 235222 668218 270986 668454
rect 271222 668218 306986 668454
rect 307222 668218 342986 668454
rect 343222 668218 378986 668454
rect 379222 668218 414986 668454
rect 415222 668218 450986 668454
rect 451222 668218 486986 668454
rect 487222 668218 522986 668454
rect 523222 668218 558986 668454
rect 559222 668218 586442 668454
rect 586678 668218 586860 668454
rect -2936 668134 586860 668218
rect -2936 667898 -2754 668134
rect -2518 667898 18986 668134
rect 19222 667898 54986 668134
rect 55222 667898 90986 668134
rect 91222 667898 126986 668134
rect 127222 667898 162986 668134
rect 163222 667898 198986 668134
rect 199222 667898 234986 668134
rect 235222 667898 270986 668134
rect 271222 667898 306986 668134
rect 307222 667898 342986 668134
rect 343222 667898 378986 668134
rect 379222 667898 414986 668134
rect 415222 667898 450986 668134
rect 451222 667898 486986 668134
rect 487222 667898 522986 668134
rect 523222 667898 558986 668134
rect 559222 667898 586442 668134
rect 586678 667898 586860 668134
rect -2936 667876 586860 667898
rect -2936 667874 -2336 667876
rect 18804 667874 19404 667876
rect 54804 667874 55404 667876
rect 90804 667874 91404 667876
rect 126804 667874 127404 667876
rect 162804 667874 163404 667876
rect 198804 667874 199404 667876
rect 234804 667874 235404 667876
rect 270804 667874 271404 667876
rect 306804 667874 307404 667876
rect 342804 667874 343404 667876
rect 378804 667874 379404 667876
rect 414804 667874 415404 667876
rect 450804 667874 451404 667876
rect 486804 667874 487404 667876
rect 522804 667874 523404 667876
rect 558804 667874 559404 667876
rect 586260 667874 586860 667876
rect -1996 650476 -1396 650478
rect 804 650476 1404 650478
rect 36804 650476 37404 650478
rect 72804 650476 73404 650478
rect 108804 650476 109404 650478
rect 144804 650476 145404 650478
rect 180804 650476 181404 650478
rect 216804 650476 217404 650478
rect 252804 650476 253404 650478
rect 288804 650476 289404 650478
rect 324804 650476 325404 650478
rect 360804 650476 361404 650478
rect 396804 650476 397404 650478
rect 432804 650476 433404 650478
rect 468804 650476 469404 650478
rect 504804 650476 505404 650478
rect 540804 650476 541404 650478
rect 576804 650476 577404 650478
rect 585320 650476 585920 650478
rect -2936 650454 586860 650476
rect -2936 650218 -1814 650454
rect -1578 650218 986 650454
rect 1222 650218 36986 650454
rect 37222 650218 72986 650454
rect 73222 650218 108986 650454
rect 109222 650218 144986 650454
rect 145222 650218 180986 650454
rect 181222 650218 216986 650454
rect 217222 650218 252986 650454
rect 253222 650218 288986 650454
rect 289222 650218 324986 650454
rect 325222 650218 360986 650454
rect 361222 650218 396986 650454
rect 397222 650218 432986 650454
rect 433222 650218 468986 650454
rect 469222 650218 504986 650454
rect 505222 650218 540986 650454
rect 541222 650218 576986 650454
rect 577222 650218 585502 650454
rect 585738 650218 586860 650454
rect -2936 650134 586860 650218
rect -2936 649898 -1814 650134
rect -1578 649898 986 650134
rect 1222 649898 36986 650134
rect 37222 649898 72986 650134
rect 73222 649898 108986 650134
rect 109222 649898 144986 650134
rect 145222 649898 180986 650134
rect 181222 649898 216986 650134
rect 217222 649898 252986 650134
rect 253222 649898 288986 650134
rect 289222 649898 324986 650134
rect 325222 649898 360986 650134
rect 361222 649898 396986 650134
rect 397222 649898 432986 650134
rect 433222 649898 468986 650134
rect 469222 649898 504986 650134
rect 505222 649898 540986 650134
rect 541222 649898 576986 650134
rect 577222 649898 585502 650134
rect 585738 649898 586860 650134
rect -2936 649876 586860 649898
rect -1996 649874 -1396 649876
rect 804 649874 1404 649876
rect 36804 649874 37404 649876
rect 72804 649874 73404 649876
rect 108804 649874 109404 649876
rect 144804 649874 145404 649876
rect 180804 649874 181404 649876
rect 216804 649874 217404 649876
rect 252804 649874 253404 649876
rect 288804 649874 289404 649876
rect 324804 649874 325404 649876
rect 360804 649874 361404 649876
rect 396804 649874 397404 649876
rect 432804 649874 433404 649876
rect 468804 649874 469404 649876
rect 504804 649874 505404 649876
rect 540804 649874 541404 649876
rect 576804 649874 577404 649876
rect 585320 649874 585920 649876
rect -2936 632476 -2336 632478
rect 18804 632476 19404 632478
rect 54804 632476 55404 632478
rect 90804 632476 91404 632478
rect 126804 632476 127404 632478
rect 162804 632476 163404 632478
rect 198804 632476 199404 632478
rect 234804 632476 235404 632478
rect 270804 632476 271404 632478
rect 306804 632476 307404 632478
rect 342804 632476 343404 632478
rect 378804 632476 379404 632478
rect 414804 632476 415404 632478
rect 450804 632476 451404 632478
rect 486804 632476 487404 632478
rect 522804 632476 523404 632478
rect 558804 632476 559404 632478
rect 586260 632476 586860 632478
rect -2936 632454 586860 632476
rect -2936 632218 -2754 632454
rect -2518 632218 18986 632454
rect 19222 632218 54986 632454
rect 55222 632218 90986 632454
rect 91222 632218 126986 632454
rect 127222 632218 162986 632454
rect 163222 632218 198986 632454
rect 199222 632218 234986 632454
rect 235222 632218 270986 632454
rect 271222 632218 306986 632454
rect 307222 632218 342986 632454
rect 343222 632218 378986 632454
rect 379222 632218 414986 632454
rect 415222 632218 450986 632454
rect 451222 632218 486986 632454
rect 487222 632218 522986 632454
rect 523222 632218 558986 632454
rect 559222 632218 586442 632454
rect 586678 632218 586860 632454
rect -2936 632134 586860 632218
rect -2936 631898 -2754 632134
rect -2518 631898 18986 632134
rect 19222 631898 54986 632134
rect 55222 631898 90986 632134
rect 91222 631898 126986 632134
rect 127222 631898 162986 632134
rect 163222 631898 198986 632134
rect 199222 631898 234986 632134
rect 235222 631898 270986 632134
rect 271222 631898 306986 632134
rect 307222 631898 342986 632134
rect 343222 631898 378986 632134
rect 379222 631898 414986 632134
rect 415222 631898 450986 632134
rect 451222 631898 486986 632134
rect 487222 631898 522986 632134
rect 523222 631898 558986 632134
rect 559222 631898 586442 632134
rect 586678 631898 586860 632134
rect -2936 631876 586860 631898
rect -2936 631874 -2336 631876
rect 18804 631874 19404 631876
rect 54804 631874 55404 631876
rect 90804 631874 91404 631876
rect 126804 631874 127404 631876
rect 162804 631874 163404 631876
rect 198804 631874 199404 631876
rect 234804 631874 235404 631876
rect 270804 631874 271404 631876
rect 306804 631874 307404 631876
rect 342804 631874 343404 631876
rect 378804 631874 379404 631876
rect 414804 631874 415404 631876
rect 450804 631874 451404 631876
rect 486804 631874 487404 631876
rect 522804 631874 523404 631876
rect 558804 631874 559404 631876
rect 586260 631874 586860 631876
rect -1996 614476 -1396 614478
rect 804 614476 1404 614478
rect 36804 614476 37404 614478
rect 72804 614476 73404 614478
rect 108804 614476 109404 614478
rect 144804 614476 145404 614478
rect 180804 614476 181404 614478
rect 216804 614476 217404 614478
rect 252804 614476 253404 614478
rect 288804 614476 289404 614478
rect 324804 614476 325404 614478
rect 360804 614476 361404 614478
rect 396804 614476 397404 614478
rect 432804 614476 433404 614478
rect 468804 614476 469404 614478
rect 504804 614476 505404 614478
rect 540804 614476 541404 614478
rect 576804 614476 577404 614478
rect 585320 614476 585920 614478
rect -2936 614454 586860 614476
rect -2936 614218 -1814 614454
rect -1578 614218 986 614454
rect 1222 614218 36986 614454
rect 37222 614218 72986 614454
rect 73222 614218 108986 614454
rect 109222 614218 144986 614454
rect 145222 614218 180986 614454
rect 181222 614218 216986 614454
rect 217222 614218 252986 614454
rect 253222 614218 288986 614454
rect 289222 614218 324986 614454
rect 325222 614218 360986 614454
rect 361222 614218 396986 614454
rect 397222 614218 432986 614454
rect 433222 614218 468986 614454
rect 469222 614218 504986 614454
rect 505222 614218 540986 614454
rect 541222 614218 576986 614454
rect 577222 614218 585502 614454
rect 585738 614218 586860 614454
rect -2936 614134 586860 614218
rect -2936 613898 -1814 614134
rect -1578 613898 986 614134
rect 1222 613898 36986 614134
rect 37222 613898 72986 614134
rect 73222 613898 108986 614134
rect 109222 613898 144986 614134
rect 145222 613898 180986 614134
rect 181222 613898 216986 614134
rect 217222 613898 252986 614134
rect 253222 613898 288986 614134
rect 289222 613898 324986 614134
rect 325222 613898 360986 614134
rect 361222 613898 396986 614134
rect 397222 613898 432986 614134
rect 433222 613898 468986 614134
rect 469222 613898 504986 614134
rect 505222 613898 540986 614134
rect 541222 613898 576986 614134
rect 577222 613898 585502 614134
rect 585738 613898 586860 614134
rect -2936 613876 586860 613898
rect -1996 613874 -1396 613876
rect 804 613874 1404 613876
rect 36804 613874 37404 613876
rect 72804 613874 73404 613876
rect 108804 613874 109404 613876
rect 144804 613874 145404 613876
rect 180804 613874 181404 613876
rect 216804 613874 217404 613876
rect 252804 613874 253404 613876
rect 288804 613874 289404 613876
rect 324804 613874 325404 613876
rect 360804 613874 361404 613876
rect 396804 613874 397404 613876
rect 432804 613874 433404 613876
rect 468804 613874 469404 613876
rect 504804 613874 505404 613876
rect 540804 613874 541404 613876
rect 576804 613874 577404 613876
rect 585320 613874 585920 613876
rect -2936 596476 -2336 596478
rect 18804 596476 19404 596478
rect 54804 596476 55404 596478
rect 90804 596476 91404 596478
rect 126804 596476 127404 596478
rect 162804 596476 163404 596478
rect 198804 596476 199404 596478
rect 234804 596476 235404 596478
rect 270804 596476 271404 596478
rect 306804 596476 307404 596478
rect 342804 596476 343404 596478
rect 378804 596476 379404 596478
rect 414804 596476 415404 596478
rect 450804 596476 451404 596478
rect 486804 596476 487404 596478
rect 522804 596476 523404 596478
rect 558804 596476 559404 596478
rect 586260 596476 586860 596478
rect -2936 596454 586860 596476
rect -2936 596218 -2754 596454
rect -2518 596218 18986 596454
rect 19222 596218 54986 596454
rect 55222 596218 90986 596454
rect 91222 596218 126986 596454
rect 127222 596218 162986 596454
rect 163222 596218 198986 596454
rect 199222 596218 234986 596454
rect 235222 596218 270986 596454
rect 271222 596218 306986 596454
rect 307222 596218 342986 596454
rect 343222 596218 378986 596454
rect 379222 596218 414986 596454
rect 415222 596218 450986 596454
rect 451222 596218 486986 596454
rect 487222 596218 522986 596454
rect 523222 596218 558986 596454
rect 559222 596218 586442 596454
rect 586678 596218 586860 596454
rect -2936 596134 586860 596218
rect -2936 595898 -2754 596134
rect -2518 595898 18986 596134
rect 19222 595898 54986 596134
rect 55222 595898 90986 596134
rect 91222 595898 126986 596134
rect 127222 595898 162986 596134
rect 163222 595898 198986 596134
rect 199222 595898 234986 596134
rect 235222 595898 270986 596134
rect 271222 595898 306986 596134
rect 307222 595898 342986 596134
rect 343222 595898 378986 596134
rect 379222 595898 414986 596134
rect 415222 595898 450986 596134
rect 451222 595898 486986 596134
rect 487222 595898 522986 596134
rect 523222 595898 558986 596134
rect 559222 595898 586442 596134
rect 586678 595898 586860 596134
rect -2936 595876 586860 595898
rect -2936 595874 -2336 595876
rect 18804 595874 19404 595876
rect 54804 595874 55404 595876
rect 90804 595874 91404 595876
rect 126804 595874 127404 595876
rect 162804 595874 163404 595876
rect 198804 595874 199404 595876
rect 234804 595874 235404 595876
rect 270804 595874 271404 595876
rect 306804 595874 307404 595876
rect 342804 595874 343404 595876
rect 378804 595874 379404 595876
rect 414804 595874 415404 595876
rect 450804 595874 451404 595876
rect 486804 595874 487404 595876
rect 522804 595874 523404 595876
rect 558804 595874 559404 595876
rect 586260 595874 586860 595876
rect -1996 578476 -1396 578478
rect 804 578476 1404 578478
rect 262128 578476 262448 578478
rect 288804 578476 289404 578478
rect 554256 578476 554576 578478
rect 576804 578476 577404 578478
rect 585320 578476 585920 578478
rect -2936 578454 586860 578476
rect -2936 578218 -1814 578454
rect -1578 578218 986 578454
rect 1222 578218 262170 578454
rect 262406 578218 288986 578454
rect 289222 578218 554298 578454
rect 554534 578218 576986 578454
rect 577222 578218 585502 578454
rect 585738 578218 586860 578454
rect -2936 578134 586860 578218
rect -2936 577898 -1814 578134
rect -1578 577898 986 578134
rect 1222 577898 262170 578134
rect 262406 577898 288986 578134
rect 289222 577898 554298 578134
rect 554534 577898 576986 578134
rect 577222 577898 585502 578134
rect 585738 577898 586860 578134
rect -2936 577876 586860 577898
rect -1996 577874 -1396 577876
rect 804 577874 1404 577876
rect 262128 577874 262448 577876
rect 288804 577874 289404 577876
rect 554256 577874 554576 577876
rect 576804 577874 577404 577876
rect 585320 577874 585920 577876
rect -2936 560476 -2336 560478
rect 18804 560476 19404 560478
rect 246768 560476 247088 560478
rect 270804 560476 271404 560478
rect 306804 560476 307404 560478
rect 538896 560476 539216 560478
rect 586260 560476 586860 560478
rect -2936 560454 586860 560476
rect -2936 560218 -2754 560454
rect -2518 560218 18986 560454
rect 19222 560218 246810 560454
rect 247046 560218 270986 560454
rect 271222 560218 306986 560454
rect 307222 560218 538938 560454
rect 539174 560218 586442 560454
rect 586678 560218 586860 560454
rect -2936 560134 586860 560218
rect -2936 559898 -2754 560134
rect -2518 559898 18986 560134
rect 19222 559898 246810 560134
rect 247046 559898 270986 560134
rect 271222 559898 306986 560134
rect 307222 559898 538938 560134
rect 539174 559898 586442 560134
rect 586678 559898 586860 560134
rect -2936 559876 586860 559898
rect -2936 559874 -2336 559876
rect 18804 559874 19404 559876
rect 246768 559874 247088 559876
rect 270804 559874 271404 559876
rect 306804 559874 307404 559876
rect 538896 559874 539216 559876
rect 586260 559874 586860 559876
rect -1996 542476 -1396 542478
rect 804 542476 1404 542478
rect 262128 542476 262448 542478
rect 288804 542476 289404 542478
rect 554256 542476 554576 542478
rect 576804 542476 577404 542478
rect 585320 542476 585920 542478
rect -2936 542454 586860 542476
rect -2936 542218 -1814 542454
rect -1578 542218 986 542454
rect 1222 542218 262170 542454
rect 262406 542218 288986 542454
rect 289222 542218 554298 542454
rect 554534 542218 576986 542454
rect 577222 542218 585502 542454
rect 585738 542218 586860 542454
rect -2936 542134 586860 542218
rect -2936 541898 -1814 542134
rect -1578 541898 986 542134
rect 1222 541898 262170 542134
rect 262406 541898 288986 542134
rect 289222 541898 554298 542134
rect 554534 541898 576986 542134
rect 577222 541898 585502 542134
rect 585738 541898 586860 542134
rect -2936 541876 586860 541898
rect -1996 541874 -1396 541876
rect 804 541874 1404 541876
rect 262128 541874 262448 541876
rect 288804 541874 289404 541876
rect 554256 541874 554576 541876
rect 576804 541874 577404 541876
rect 585320 541874 585920 541876
rect -2936 524476 -2336 524478
rect 18804 524476 19404 524478
rect 246768 524476 247088 524478
rect 270804 524476 271404 524478
rect 306804 524476 307404 524478
rect 538896 524476 539216 524478
rect 586260 524476 586860 524478
rect -2936 524454 586860 524476
rect -2936 524218 -2754 524454
rect -2518 524218 18986 524454
rect 19222 524218 246810 524454
rect 247046 524218 270986 524454
rect 271222 524218 306986 524454
rect 307222 524218 538938 524454
rect 539174 524218 586442 524454
rect 586678 524218 586860 524454
rect -2936 524134 586860 524218
rect -2936 523898 -2754 524134
rect -2518 523898 18986 524134
rect 19222 523898 246810 524134
rect 247046 523898 270986 524134
rect 271222 523898 306986 524134
rect 307222 523898 538938 524134
rect 539174 523898 586442 524134
rect 586678 523898 586860 524134
rect -2936 523876 586860 523898
rect -2936 523874 -2336 523876
rect 18804 523874 19404 523876
rect 246768 523874 247088 523876
rect 270804 523874 271404 523876
rect 306804 523874 307404 523876
rect 538896 523874 539216 523876
rect 586260 523874 586860 523876
rect -1996 506476 -1396 506478
rect 804 506476 1404 506478
rect 262128 506476 262448 506478
rect 288804 506476 289404 506478
rect 554256 506476 554576 506478
rect 576804 506476 577404 506478
rect 585320 506476 585920 506478
rect -2936 506454 586860 506476
rect -2936 506218 -1814 506454
rect -1578 506218 986 506454
rect 1222 506218 262170 506454
rect 262406 506218 288986 506454
rect 289222 506218 554298 506454
rect 554534 506218 576986 506454
rect 577222 506218 585502 506454
rect 585738 506218 586860 506454
rect -2936 506134 586860 506218
rect -2936 505898 -1814 506134
rect -1578 505898 986 506134
rect 1222 505898 262170 506134
rect 262406 505898 288986 506134
rect 289222 505898 554298 506134
rect 554534 505898 576986 506134
rect 577222 505898 585502 506134
rect 585738 505898 586860 506134
rect -2936 505876 586860 505898
rect -1996 505874 -1396 505876
rect 804 505874 1404 505876
rect 262128 505874 262448 505876
rect 288804 505874 289404 505876
rect 554256 505874 554576 505876
rect 576804 505874 577404 505876
rect 585320 505874 585920 505876
rect -2936 488476 -2336 488478
rect 18804 488476 19404 488478
rect 246768 488476 247088 488478
rect 270804 488476 271404 488478
rect 306804 488476 307404 488478
rect 538896 488476 539216 488478
rect 586260 488476 586860 488478
rect -2936 488454 586860 488476
rect -2936 488218 -2754 488454
rect -2518 488218 18986 488454
rect 19222 488218 246810 488454
rect 247046 488218 270986 488454
rect 271222 488218 306986 488454
rect 307222 488218 538938 488454
rect 539174 488218 586442 488454
rect 586678 488218 586860 488454
rect -2936 488134 586860 488218
rect -2936 487898 -2754 488134
rect -2518 487898 18986 488134
rect 19222 487898 246810 488134
rect 247046 487898 270986 488134
rect 271222 487898 306986 488134
rect 307222 487898 538938 488134
rect 539174 487898 586442 488134
rect 586678 487898 586860 488134
rect -2936 487876 586860 487898
rect -2936 487874 -2336 487876
rect 18804 487874 19404 487876
rect 246768 487874 247088 487876
rect 270804 487874 271404 487876
rect 306804 487874 307404 487876
rect 538896 487874 539216 487876
rect 586260 487874 586860 487876
rect -1996 470476 -1396 470478
rect 804 470476 1404 470478
rect 262128 470476 262448 470478
rect 288804 470476 289404 470478
rect 554256 470476 554576 470478
rect 576804 470476 577404 470478
rect 585320 470476 585920 470478
rect -2936 470454 586860 470476
rect -2936 470218 -1814 470454
rect -1578 470218 986 470454
rect 1222 470218 262170 470454
rect 262406 470218 288986 470454
rect 289222 470218 554298 470454
rect 554534 470218 576986 470454
rect 577222 470218 585502 470454
rect 585738 470218 586860 470454
rect -2936 470134 586860 470218
rect -2936 469898 -1814 470134
rect -1578 469898 986 470134
rect 1222 469898 262170 470134
rect 262406 469898 288986 470134
rect 289222 469898 554298 470134
rect 554534 469898 576986 470134
rect 577222 469898 585502 470134
rect 585738 469898 586860 470134
rect -2936 469876 586860 469898
rect -1996 469874 -1396 469876
rect 804 469874 1404 469876
rect 262128 469874 262448 469876
rect 288804 469874 289404 469876
rect 554256 469874 554576 469876
rect 576804 469874 577404 469876
rect 585320 469874 585920 469876
rect -2936 452476 -2336 452478
rect 18804 452476 19404 452478
rect 246768 452476 247088 452478
rect 270804 452476 271404 452478
rect 306804 452476 307404 452478
rect 538896 452476 539216 452478
rect 586260 452476 586860 452478
rect -2936 452454 586860 452476
rect -2936 452218 -2754 452454
rect -2518 452218 18986 452454
rect 19222 452218 246810 452454
rect 247046 452218 270986 452454
rect 271222 452218 306986 452454
rect 307222 452218 538938 452454
rect 539174 452218 586442 452454
rect 586678 452218 586860 452454
rect -2936 452134 586860 452218
rect -2936 451898 -2754 452134
rect -2518 451898 18986 452134
rect 19222 451898 246810 452134
rect 247046 451898 270986 452134
rect 271222 451898 306986 452134
rect 307222 451898 538938 452134
rect 539174 451898 586442 452134
rect 586678 451898 586860 452134
rect -2936 451876 586860 451898
rect -2936 451874 -2336 451876
rect 18804 451874 19404 451876
rect 246768 451874 247088 451876
rect 270804 451874 271404 451876
rect 306804 451874 307404 451876
rect 538896 451874 539216 451876
rect 586260 451874 586860 451876
rect -1996 434476 -1396 434478
rect 804 434476 1404 434478
rect 262128 434476 262448 434478
rect 288804 434476 289404 434478
rect 554256 434476 554576 434478
rect 576804 434476 577404 434478
rect 585320 434476 585920 434478
rect -2936 434454 586860 434476
rect -2936 434218 -1814 434454
rect -1578 434218 986 434454
rect 1222 434218 262170 434454
rect 262406 434218 288986 434454
rect 289222 434218 554298 434454
rect 554534 434218 576986 434454
rect 577222 434218 585502 434454
rect 585738 434218 586860 434454
rect -2936 434134 586860 434218
rect -2936 433898 -1814 434134
rect -1578 433898 986 434134
rect 1222 433898 262170 434134
rect 262406 433898 288986 434134
rect 289222 433898 554298 434134
rect 554534 433898 576986 434134
rect 577222 433898 585502 434134
rect 585738 433898 586860 434134
rect -2936 433876 586860 433898
rect -1996 433874 -1396 433876
rect 804 433874 1404 433876
rect 262128 433874 262448 433876
rect 288804 433874 289404 433876
rect 554256 433874 554576 433876
rect 576804 433874 577404 433876
rect 585320 433874 585920 433876
rect -2936 416476 -2336 416478
rect 18804 416476 19404 416478
rect 246768 416476 247088 416478
rect 270804 416476 271404 416478
rect 306804 416476 307404 416478
rect 538896 416476 539216 416478
rect 586260 416476 586860 416478
rect -2936 416454 586860 416476
rect -2936 416218 -2754 416454
rect -2518 416218 18986 416454
rect 19222 416218 246810 416454
rect 247046 416218 270986 416454
rect 271222 416218 306986 416454
rect 307222 416218 538938 416454
rect 539174 416218 586442 416454
rect 586678 416218 586860 416454
rect -2936 416134 586860 416218
rect -2936 415898 -2754 416134
rect -2518 415898 18986 416134
rect 19222 415898 246810 416134
rect 247046 415898 270986 416134
rect 271222 415898 306986 416134
rect 307222 415898 538938 416134
rect 539174 415898 586442 416134
rect 586678 415898 586860 416134
rect -2936 415876 586860 415898
rect -2936 415874 -2336 415876
rect 18804 415874 19404 415876
rect 246768 415874 247088 415876
rect 270804 415874 271404 415876
rect 306804 415874 307404 415876
rect 538896 415874 539216 415876
rect 586260 415874 586860 415876
rect -1996 398476 -1396 398478
rect 804 398476 1404 398478
rect 262128 398476 262448 398478
rect 288804 398476 289404 398478
rect 554256 398476 554576 398478
rect 576804 398476 577404 398478
rect 585320 398476 585920 398478
rect -2936 398454 586860 398476
rect -2936 398218 -1814 398454
rect -1578 398218 986 398454
rect 1222 398218 262170 398454
rect 262406 398218 288986 398454
rect 289222 398218 554298 398454
rect 554534 398218 576986 398454
rect 577222 398218 585502 398454
rect 585738 398218 586860 398454
rect -2936 398134 586860 398218
rect -2936 397898 -1814 398134
rect -1578 397898 986 398134
rect 1222 397898 262170 398134
rect 262406 397898 288986 398134
rect 289222 397898 554298 398134
rect 554534 397898 576986 398134
rect 577222 397898 585502 398134
rect 585738 397898 586860 398134
rect -2936 397876 586860 397898
rect -1996 397874 -1396 397876
rect 804 397874 1404 397876
rect 262128 397874 262448 397876
rect 288804 397874 289404 397876
rect 554256 397874 554576 397876
rect 576804 397874 577404 397876
rect 585320 397874 585920 397876
rect -2936 380476 -2336 380478
rect 18804 380476 19404 380478
rect 54804 380476 55404 380478
rect 90804 380476 91404 380478
rect 126804 380476 127404 380478
rect 162804 380476 163404 380478
rect 198804 380476 199404 380478
rect 234804 380476 235404 380478
rect 270804 380476 271404 380478
rect 306804 380476 307404 380478
rect 342804 380476 343404 380478
rect 378804 380476 379404 380478
rect 414804 380476 415404 380478
rect 450804 380476 451404 380478
rect 486804 380476 487404 380478
rect 522804 380476 523404 380478
rect 558804 380476 559404 380478
rect 586260 380476 586860 380478
rect -2936 380454 586860 380476
rect -2936 380218 -2754 380454
rect -2518 380218 18986 380454
rect 19222 380218 54986 380454
rect 55222 380218 90986 380454
rect 91222 380218 126986 380454
rect 127222 380218 162986 380454
rect 163222 380218 198986 380454
rect 199222 380218 234986 380454
rect 235222 380218 270986 380454
rect 271222 380218 306986 380454
rect 307222 380218 342986 380454
rect 343222 380218 378986 380454
rect 379222 380218 414986 380454
rect 415222 380218 450986 380454
rect 451222 380218 486986 380454
rect 487222 380218 522986 380454
rect 523222 380218 558986 380454
rect 559222 380218 586442 380454
rect 586678 380218 586860 380454
rect -2936 380134 586860 380218
rect -2936 379898 -2754 380134
rect -2518 379898 18986 380134
rect 19222 379898 54986 380134
rect 55222 379898 90986 380134
rect 91222 379898 126986 380134
rect 127222 379898 162986 380134
rect 163222 379898 198986 380134
rect 199222 379898 234986 380134
rect 235222 379898 270986 380134
rect 271222 379898 306986 380134
rect 307222 379898 342986 380134
rect 343222 379898 378986 380134
rect 379222 379898 414986 380134
rect 415222 379898 450986 380134
rect 451222 379898 486986 380134
rect 487222 379898 522986 380134
rect 523222 379898 558986 380134
rect 559222 379898 586442 380134
rect 586678 379898 586860 380134
rect -2936 379876 586860 379898
rect -2936 379874 -2336 379876
rect 18804 379874 19404 379876
rect 54804 379874 55404 379876
rect 90804 379874 91404 379876
rect 126804 379874 127404 379876
rect 162804 379874 163404 379876
rect 198804 379874 199404 379876
rect 234804 379874 235404 379876
rect 270804 379874 271404 379876
rect 306804 379874 307404 379876
rect 342804 379874 343404 379876
rect 378804 379874 379404 379876
rect 414804 379874 415404 379876
rect 450804 379874 451404 379876
rect 486804 379874 487404 379876
rect 522804 379874 523404 379876
rect 558804 379874 559404 379876
rect 586260 379874 586860 379876
rect -1996 362476 -1396 362478
rect 804 362476 1404 362478
rect 36804 362476 37404 362478
rect 72804 362476 73404 362478
rect 108804 362476 109404 362478
rect 144804 362476 145404 362478
rect 180804 362476 181404 362478
rect 216804 362476 217404 362478
rect 252804 362476 253404 362478
rect 288804 362476 289404 362478
rect 324804 362476 325404 362478
rect 360804 362476 361404 362478
rect 396804 362476 397404 362478
rect 432804 362476 433404 362478
rect 468804 362476 469404 362478
rect 504804 362476 505404 362478
rect 540804 362476 541404 362478
rect 576804 362476 577404 362478
rect 585320 362476 585920 362478
rect -2936 362454 586860 362476
rect -2936 362218 -1814 362454
rect -1578 362218 986 362454
rect 1222 362218 36986 362454
rect 37222 362218 72986 362454
rect 73222 362218 108986 362454
rect 109222 362218 144986 362454
rect 145222 362218 180986 362454
rect 181222 362218 216986 362454
rect 217222 362218 252986 362454
rect 253222 362218 288986 362454
rect 289222 362218 324986 362454
rect 325222 362218 360986 362454
rect 361222 362218 396986 362454
rect 397222 362218 432986 362454
rect 433222 362218 468986 362454
rect 469222 362218 504986 362454
rect 505222 362218 540986 362454
rect 541222 362218 576986 362454
rect 577222 362218 585502 362454
rect 585738 362218 586860 362454
rect -2936 362134 586860 362218
rect -2936 361898 -1814 362134
rect -1578 361898 986 362134
rect 1222 361898 36986 362134
rect 37222 361898 72986 362134
rect 73222 361898 108986 362134
rect 109222 361898 144986 362134
rect 145222 361898 180986 362134
rect 181222 361898 216986 362134
rect 217222 361898 252986 362134
rect 253222 361898 288986 362134
rect 289222 361898 324986 362134
rect 325222 361898 360986 362134
rect 361222 361898 396986 362134
rect 397222 361898 432986 362134
rect 433222 361898 468986 362134
rect 469222 361898 504986 362134
rect 505222 361898 540986 362134
rect 541222 361898 576986 362134
rect 577222 361898 585502 362134
rect 585738 361898 586860 362134
rect -2936 361876 586860 361898
rect -1996 361874 -1396 361876
rect 804 361874 1404 361876
rect 36804 361874 37404 361876
rect 72804 361874 73404 361876
rect 108804 361874 109404 361876
rect 144804 361874 145404 361876
rect 180804 361874 181404 361876
rect 216804 361874 217404 361876
rect 252804 361874 253404 361876
rect 288804 361874 289404 361876
rect 324804 361874 325404 361876
rect 360804 361874 361404 361876
rect 396804 361874 397404 361876
rect 432804 361874 433404 361876
rect 468804 361874 469404 361876
rect 504804 361874 505404 361876
rect 540804 361874 541404 361876
rect 576804 361874 577404 361876
rect 585320 361874 585920 361876
rect -2936 344476 -2336 344478
rect 18804 344476 19404 344478
rect 54804 344476 55404 344478
rect 90804 344476 91404 344478
rect 126804 344476 127404 344478
rect 162804 344476 163404 344478
rect 198804 344476 199404 344478
rect 234804 344476 235404 344478
rect 292112 344476 292432 344478
rect 342804 344476 343404 344478
rect 378804 344476 379404 344478
rect 414804 344476 415404 344478
rect 450804 344476 451404 344478
rect 486804 344476 487404 344478
rect 522804 344476 523404 344478
rect 558804 344476 559404 344478
rect 586260 344476 586860 344478
rect -2936 344454 586860 344476
rect -2936 344218 -2754 344454
rect -2518 344218 18986 344454
rect 19222 344218 54986 344454
rect 55222 344218 90986 344454
rect 91222 344218 126986 344454
rect 127222 344218 162986 344454
rect 163222 344218 198986 344454
rect 199222 344218 234986 344454
rect 235222 344218 292154 344454
rect 292390 344218 342986 344454
rect 343222 344218 378986 344454
rect 379222 344218 414986 344454
rect 415222 344218 450986 344454
rect 451222 344218 486986 344454
rect 487222 344218 522986 344454
rect 523222 344218 558986 344454
rect 559222 344218 586442 344454
rect 586678 344218 586860 344454
rect -2936 344134 586860 344218
rect -2936 343898 -2754 344134
rect -2518 343898 18986 344134
rect 19222 343898 54986 344134
rect 55222 343898 90986 344134
rect 91222 343898 126986 344134
rect 127222 343898 162986 344134
rect 163222 343898 198986 344134
rect 199222 343898 234986 344134
rect 235222 343898 292154 344134
rect 292390 343898 342986 344134
rect 343222 343898 378986 344134
rect 379222 343898 414986 344134
rect 415222 343898 450986 344134
rect 451222 343898 486986 344134
rect 487222 343898 522986 344134
rect 523222 343898 558986 344134
rect 559222 343898 586442 344134
rect 586678 343898 586860 344134
rect -2936 343876 586860 343898
rect -2936 343874 -2336 343876
rect 18804 343874 19404 343876
rect 54804 343874 55404 343876
rect 90804 343874 91404 343876
rect 126804 343874 127404 343876
rect 162804 343874 163404 343876
rect 198804 343874 199404 343876
rect 234804 343874 235404 343876
rect 292112 343874 292432 343876
rect 342804 343874 343404 343876
rect 378804 343874 379404 343876
rect 414804 343874 415404 343876
rect 450804 343874 451404 343876
rect 486804 343874 487404 343876
rect 522804 343874 523404 343876
rect 558804 343874 559404 343876
rect 586260 343874 586860 343876
rect -1996 326476 -1396 326478
rect 804 326476 1404 326478
rect 36804 326476 37404 326478
rect 72804 326476 73404 326478
rect 108804 326476 109404 326478
rect 144804 326476 145404 326478
rect 180804 326476 181404 326478
rect 216804 326476 217404 326478
rect 252804 326476 253404 326478
rect 307472 326476 307792 326478
rect 324804 326476 325404 326478
rect 360804 326476 361404 326478
rect 396804 326476 397404 326478
rect 432804 326476 433404 326478
rect 468804 326476 469404 326478
rect 504804 326476 505404 326478
rect 540804 326476 541404 326478
rect 576804 326476 577404 326478
rect 585320 326476 585920 326478
rect -2936 326454 586860 326476
rect -2936 326218 -1814 326454
rect -1578 326218 986 326454
rect 1222 326218 36986 326454
rect 37222 326218 72986 326454
rect 73222 326218 108986 326454
rect 109222 326218 144986 326454
rect 145222 326218 180986 326454
rect 181222 326218 216986 326454
rect 217222 326218 252986 326454
rect 253222 326218 307514 326454
rect 307750 326218 324986 326454
rect 325222 326218 360986 326454
rect 361222 326218 396986 326454
rect 397222 326218 432986 326454
rect 433222 326218 468986 326454
rect 469222 326218 504986 326454
rect 505222 326218 540986 326454
rect 541222 326218 576986 326454
rect 577222 326218 585502 326454
rect 585738 326218 586860 326454
rect -2936 326134 586860 326218
rect -2936 325898 -1814 326134
rect -1578 325898 986 326134
rect 1222 325898 36986 326134
rect 37222 325898 72986 326134
rect 73222 325898 108986 326134
rect 109222 325898 144986 326134
rect 145222 325898 180986 326134
rect 181222 325898 216986 326134
rect 217222 325898 252986 326134
rect 253222 325898 307514 326134
rect 307750 325898 324986 326134
rect 325222 325898 360986 326134
rect 361222 325898 396986 326134
rect 397222 325898 432986 326134
rect 433222 325898 468986 326134
rect 469222 325898 504986 326134
rect 505222 325898 540986 326134
rect 541222 325898 576986 326134
rect 577222 325898 585502 326134
rect 585738 325898 586860 326134
rect -2936 325876 586860 325898
rect -1996 325874 -1396 325876
rect 804 325874 1404 325876
rect 36804 325874 37404 325876
rect 72804 325874 73404 325876
rect 108804 325874 109404 325876
rect 144804 325874 145404 325876
rect 180804 325874 181404 325876
rect 216804 325874 217404 325876
rect 252804 325874 253404 325876
rect 307472 325874 307792 325876
rect 324804 325874 325404 325876
rect 360804 325874 361404 325876
rect 396804 325874 397404 325876
rect 432804 325874 433404 325876
rect 468804 325874 469404 325876
rect 504804 325874 505404 325876
rect 540804 325874 541404 325876
rect 576804 325874 577404 325876
rect 585320 325874 585920 325876
rect -2936 308476 -2336 308478
rect 18804 308476 19404 308478
rect 54804 308476 55404 308478
rect 90804 308476 91404 308478
rect 126804 308476 127404 308478
rect 162804 308476 163404 308478
rect 198804 308476 199404 308478
rect 234804 308476 235404 308478
rect 270804 308476 271404 308478
rect 306804 308476 307404 308478
rect 342804 308476 343404 308478
rect 378804 308476 379404 308478
rect 414804 308476 415404 308478
rect 450804 308476 451404 308478
rect 486804 308476 487404 308478
rect 522804 308476 523404 308478
rect 558804 308476 559404 308478
rect 586260 308476 586860 308478
rect -2936 308454 586860 308476
rect -2936 308218 -2754 308454
rect -2518 308218 18986 308454
rect 19222 308218 54986 308454
rect 55222 308218 90986 308454
rect 91222 308218 126986 308454
rect 127222 308218 162986 308454
rect 163222 308218 198986 308454
rect 199222 308218 234986 308454
rect 235222 308218 270986 308454
rect 271222 308218 306986 308454
rect 307222 308218 342986 308454
rect 343222 308218 378986 308454
rect 379222 308218 414986 308454
rect 415222 308218 450986 308454
rect 451222 308218 486986 308454
rect 487222 308218 522986 308454
rect 523222 308218 558986 308454
rect 559222 308218 586442 308454
rect 586678 308218 586860 308454
rect -2936 308134 586860 308218
rect -2936 307898 -2754 308134
rect -2518 307898 18986 308134
rect 19222 307898 54986 308134
rect 55222 307898 90986 308134
rect 91222 307898 126986 308134
rect 127222 307898 162986 308134
rect 163222 307898 198986 308134
rect 199222 307898 234986 308134
rect 235222 307898 270986 308134
rect 271222 307898 306986 308134
rect 307222 307898 342986 308134
rect 343222 307898 378986 308134
rect 379222 307898 414986 308134
rect 415222 307898 450986 308134
rect 451222 307898 486986 308134
rect 487222 307898 522986 308134
rect 523222 307898 558986 308134
rect 559222 307898 586442 308134
rect 586678 307898 586860 308134
rect -2936 307876 586860 307898
rect -2936 307874 -2336 307876
rect 18804 307874 19404 307876
rect 54804 307874 55404 307876
rect 90804 307874 91404 307876
rect 126804 307874 127404 307876
rect 162804 307874 163404 307876
rect 198804 307874 199404 307876
rect 234804 307874 235404 307876
rect 270804 307874 271404 307876
rect 306804 307874 307404 307876
rect 342804 307874 343404 307876
rect 378804 307874 379404 307876
rect 414804 307874 415404 307876
rect 450804 307874 451404 307876
rect 486804 307874 487404 307876
rect 522804 307874 523404 307876
rect 558804 307874 559404 307876
rect 586260 307874 586860 307876
rect -1996 290476 -1396 290478
rect 804 290476 1404 290478
rect 36804 290476 37404 290478
rect 72804 290476 73404 290478
rect 108804 290476 109404 290478
rect 144804 290476 145404 290478
rect 180804 290476 181404 290478
rect 216804 290476 217404 290478
rect 252804 290476 253404 290478
rect 288804 290476 289404 290478
rect 324804 290476 325404 290478
rect 360804 290476 361404 290478
rect 396804 290476 397404 290478
rect 432804 290476 433404 290478
rect 468804 290476 469404 290478
rect 504804 290476 505404 290478
rect 540804 290476 541404 290478
rect 576804 290476 577404 290478
rect 585320 290476 585920 290478
rect -2936 290454 586860 290476
rect -2936 290218 -1814 290454
rect -1578 290218 986 290454
rect 1222 290218 36986 290454
rect 37222 290218 72986 290454
rect 73222 290218 108986 290454
rect 109222 290218 144986 290454
rect 145222 290218 180986 290454
rect 181222 290218 216986 290454
rect 217222 290218 252986 290454
rect 253222 290218 288986 290454
rect 289222 290218 324986 290454
rect 325222 290218 360986 290454
rect 361222 290218 396986 290454
rect 397222 290218 432986 290454
rect 433222 290218 468986 290454
rect 469222 290218 504986 290454
rect 505222 290218 540986 290454
rect 541222 290218 576986 290454
rect 577222 290218 585502 290454
rect 585738 290218 586860 290454
rect -2936 290134 586860 290218
rect -2936 289898 -1814 290134
rect -1578 289898 986 290134
rect 1222 289898 36986 290134
rect 37222 289898 72986 290134
rect 73222 289898 108986 290134
rect 109222 289898 144986 290134
rect 145222 289898 180986 290134
rect 181222 289898 216986 290134
rect 217222 289898 252986 290134
rect 253222 289898 288986 290134
rect 289222 289898 324986 290134
rect 325222 289898 360986 290134
rect 361222 289898 396986 290134
rect 397222 289898 432986 290134
rect 433222 289898 468986 290134
rect 469222 289898 504986 290134
rect 505222 289898 540986 290134
rect 541222 289898 576986 290134
rect 577222 289898 585502 290134
rect 585738 289898 586860 290134
rect -2936 289876 586860 289898
rect -1996 289874 -1396 289876
rect 804 289874 1404 289876
rect 36804 289874 37404 289876
rect 72804 289874 73404 289876
rect 108804 289874 109404 289876
rect 144804 289874 145404 289876
rect 180804 289874 181404 289876
rect 216804 289874 217404 289876
rect 252804 289874 253404 289876
rect 288804 289874 289404 289876
rect 324804 289874 325404 289876
rect 360804 289874 361404 289876
rect 396804 289874 397404 289876
rect 432804 289874 433404 289876
rect 468804 289874 469404 289876
rect 504804 289874 505404 289876
rect 540804 289874 541404 289876
rect 576804 289874 577404 289876
rect 585320 289874 585920 289876
rect -2936 272476 -2336 272478
rect 18804 272476 19404 272478
rect 270804 272476 271404 272478
rect 306804 272476 307404 272478
rect 586260 272476 586860 272478
rect -2936 272454 586860 272476
rect -2936 272218 -2754 272454
rect -2518 272218 18986 272454
rect 19222 272218 270986 272454
rect 271222 272218 306986 272454
rect 307222 272218 586442 272454
rect 586678 272218 586860 272454
rect -2936 272134 586860 272218
rect -2936 271898 -2754 272134
rect -2518 271898 18986 272134
rect 19222 271898 270986 272134
rect 271222 271898 306986 272134
rect 307222 271898 586442 272134
rect 586678 271898 586860 272134
rect -2936 271876 586860 271898
rect -2936 271874 -2336 271876
rect 18804 271874 19404 271876
rect 270804 271874 271404 271876
rect 306804 271874 307404 271876
rect 586260 271874 586860 271876
rect -1996 254476 -1396 254478
rect 804 254476 1404 254478
rect 262128 254476 262448 254478
rect 288804 254476 289404 254478
rect 554256 254476 554576 254478
rect 576804 254476 577404 254478
rect 585320 254476 585920 254478
rect -2936 254454 586860 254476
rect -2936 254218 -1814 254454
rect -1578 254218 986 254454
rect 1222 254218 262170 254454
rect 262406 254218 288986 254454
rect 289222 254218 554298 254454
rect 554534 254218 576986 254454
rect 577222 254218 585502 254454
rect 585738 254218 586860 254454
rect -2936 254134 586860 254218
rect -2936 253898 -1814 254134
rect -1578 253898 986 254134
rect 1222 253898 262170 254134
rect 262406 253898 288986 254134
rect 289222 253898 554298 254134
rect 554534 253898 576986 254134
rect 577222 253898 585502 254134
rect 585738 253898 586860 254134
rect -2936 253876 586860 253898
rect -1996 253874 -1396 253876
rect 804 253874 1404 253876
rect 262128 253874 262448 253876
rect 288804 253874 289404 253876
rect 554256 253874 554576 253876
rect 576804 253874 577404 253876
rect 585320 253874 585920 253876
rect -2936 236476 -2336 236478
rect 18804 236476 19404 236478
rect 246768 236476 247088 236478
rect 270804 236476 271404 236478
rect 306804 236476 307404 236478
rect 538896 236476 539216 236478
rect 586260 236476 586860 236478
rect -2936 236454 586860 236476
rect -2936 236218 -2754 236454
rect -2518 236218 18986 236454
rect 19222 236218 246810 236454
rect 247046 236218 270986 236454
rect 271222 236218 306986 236454
rect 307222 236218 538938 236454
rect 539174 236218 586442 236454
rect 586678 236218 586860 236454
rect -2936 236134 586860 236218
rect -2936 235898 -2754 236134
rect -2518 235898 18986 236134
rect 19222 235898 246810 236134
rect 247046 235898 270986 236134
rect 271222 235898 306986 236134
rect 307222 235898 538938 236134
rect 539174 235898 586442 236134
rect 586678 235898 586860 236134
rect -2936 235876 586860 235898
rect -2936 235874 -2336 235876
rect 18804 235874 19404 235876
rect 246768 235874 247088 235876
rect 270804 235874 271404 235876
rect 306804 235874 307404 235876
rect 538896 235874 539216 235876
rect 586260 235874 586860 235876
rect -1996 218476 -1396 218478
rect 804 218476 1404 218478
rect 262128 218476 262448 218478
rect 288804 218476 289404 218478
rect 554256 218476 554576 218478
rect 576804 218476 577404 218478
rect 585320 218476 585920 218478
rect -2936 218454 586860 218476
rect -2936 218218 -1814 218454
rect -1578 218218 986 218454
rect 1222 218218 262170 218454
rect 262406 218218 288986 218454
rect 289222 218218 554298 218454
rect 554534 218218 576986 218454
rect 577222 218218 585502 218454
rect 585738 218218 586860 218454
rect -2936 218134 586860 218218
rect -2936 217898 -1814 218134
rect -1578 217898 986 218134
rect 1222 217898 262170 218134
rect 262406 217898 288986 218134
rect 289222 217898 554298 218134
rect 554534 217898 576986 218134
rect 577222 217898 585502 218134
rect 585738 217898 586860 218134
rect -2936 217876 586860 217898
rect -1996 217874 -1396 217876
rect 804 217874 1404 217876
rect 262128 217874 262448 217876
rect 288804 217874 289404 217876
rect 554256 217874 554576 217876
rect 576804 217874 577404 217876
rect 585320 217874 585920 217876
rect -2936 200476 -2336 200478
rect 18804 200476 19404 200478
rect 246768 200476 247088 200478
rect 270804 200476 271404 200478
rect 306804 200476 307404 200478
rect 538896 200476 539216 200478
rect 586260 200476 586860 200478
rect -2936 200454 586860 200476
rect -2936 200218 -2754 200454
rect -2518 200218 18986 200454
rect 19222 200218 246810 200454
rect 247046 200218 270986 200454
rect 271222 200218 306986 200454
rect 307222 200218 538938 200454
rect 539174 200218 586442 200454
rect 586678 200218 586860 200454
rect -2936 200134 586860 200218
rect -2936 199898 -2754 200134
rect -2518 199898 18986 200134
rect 19222 199898 246810 200134
rect 247046 199898 270986 200134
rect 271222 199898 306986 200134
rect 307222 199898 538938 200134
rect 539174 199898 586442 200134
rect 586678 199898 586860 200134
rect -2936 199876 586860 199898
rect -2936 199874 -2336 199876
rect 18804 199874 19404 199876
rect 246768 199874 247088 199876
rect 270804 199874 271404 199876
rect 306804 199874 307404 199876
rect 538896 199874 539216 199876
rect 586260 199874 586860 199876
rect -1996 182476 -1396 182478
rect 804 182476 1404 182478
rect 262128 182476 262448 182478
rect 288804 182476 289404 182478
rect 554256 182476 554576 182478
rect 576804 182476 577404 182478
rect 585320 182476 585920 182478
rect -2936 182454 586860 182476
rect -2936 182218 -1814 182454
rect -1578 182218 986 182454
rect 1222 182218 262170 182454
rect 262406 182218 288986 182454
rect 289222 182218 554298 182454
rect 554534 182218 576986 182454
rect 577222 182218 585502 182454
rect 585738 182218 586860 182454
rect -2936 182134 586860 182218
rect -2936 181898 -1814 182134
rect -1578 181898 986 182134
rect 1222 181898 262170 182134
rect 262406 181898 288986 182134
rect 289222 181898 554298 182134
rect 554534 181898 576986 182134
rect 577222 181898 585502 182134
rect 585738 181898 586860 182134
rect -2936 181876 586860 181898
rect -1996 181874 -1396 181876
rect 804 181874 1404 181876
rect 262128 181874 262448 181876
rect 288804 181874 289404 181876
rect 554256 181874 554576 181876
rect 576804 181874 577404 181876
rect 585320 181874 585920 181876
rect -2936 164476 -2336 164478
rect 18804 164476 19404 164478
rect 246768 164476 247088 164478
rect 270804 164476 271404 164478
rect 306804 164476 307404 164478
rect 538896 164476 539216 164478
rect 586260 164476 586860 164478
rect -2936 164454 586860 164476
rect -2936 164218 -2754 164454
rect -2518 164218 18986 164454
rect 19222 164218 246810 164454
rect 247046 164218 270986 164454
rect 271222 164218 306986 164454
rect 307222 164218 538938 164454
rect 539174 164218 586442 164454
rect 586678 164218 586860 164454
rect -2936 164134 586860 164218
rect -2936 163898 -2754 164134
rect -2518 163898 18986 164134
rect 19222 163898 246810 164134
rect 247046 163898 270986 164134
rect 271222 163898 306986 164134
rect 307222 163898 538938 164134
rect 539174 163898 586442 164134
rect 586678 163898 586860 164134
rect -2936 163876 586860 163898
rect -2936 163874 -2336 163876
rect 18804 163874 19404 163876
rect 246768 163874 247088 163876
rect 270804 163874 271404 163876
rect 306804 163874 307404 163876
rect 538896 163874 539216 163876
rect 586260 163874 586860 163876
rect -1996 146476 -1396 146478
rect 804 146476 1404 146478
rect 262128 146476 262448 146478
rect 288804 146476 289404 146478
rect 554256 146476 554576 146478
rect 576804 146476 577404 146478
rect 585320 146476 585920 146478
rect -2936 146454 586860 146476
rect -2936 146218 -1814 146454
rect -1578 146218 986 146454
rect 1222 146218 262170 146454
rect 262406 146218 288986 146454
rect 289222 146218 554298 146454
rect 554534 146218 576986 146454
rect 577222 146218 585502 146454
rect 585738 146218 586860 146454
rect -2936 146134 586860 146218
rect -2936 145898 -1814 146134
rect -1578 145898 986 146134
rect 1222 145898 262170 146134
rect 262406 145898 288986 146134
rect 289222 145898 554298 146134
rect 554534 145898 576986 146134
rect 577222 145898 585502 146134
rect 585738 145898 586860 146134
rect -2936 145876 586860 145898
rect -1996 145874 -1396 145876
rect 804 145874 1404 145876
rect 262128 145874 262448 145876
rect 288804 145874 289404 145876
rect 554256 145874 554576 145876
rect 576804 145874 577404 145876
rect 585320 145874 585920 145876
rect -2936 128476 -2336 128478
rect 18804 128476 19404 128478
rect 246768 128476 247088 128478
rect 270804 128476 271404 128478
rect 306804 128476 307404 128478
rect 538896 128476 539216 128478
rect 586260 128476 586860 128478
rect -2936 128454 586860 128476
rect -2936 128218 -2754 128454
rect -2518 128218 18986 128454
rect 19222 128218 246810 128454
rect 247046 128218 270986 128454
rect 271222 128218 306986 128454
rect 307222 128218 538938 128454
rect 539174 128218 586442 128454
rect 586678 128218 586860 128454
rect -2936 128134 586860 128218
rect -2936 127898 -2754 128134
rect -2518 127898 18986 128134
rect 19222 127898 246810 128134
rect 247046 127898 270986 128134
rect 271222 127898 306986 128134
rect 307222 127898 538938 128134
rect 539174 127898 586442 128134
rect 586678 127898 586860 128134
rect -2936 127876 586860 127898
rect -2936 127874 -2336 127876
rect 18804 127874 19404 127876
rect 246768 127874 247088 127876
rect 270804 127874 271404 127876
rect 306804 127874 307404 127876
rect 538896 127874 539216 127876
rect 586260 127874 586860 127876
rect -1996 110476 -1396 110478
rect 804 110476 1404 110478
rect 262128 110476 262448 110478
rect 288804 110476 289404 110478
rect 554256 110476 554576 110478
rect 576804 110476 577404 110478
rect 585320 110476 585920 110478
rect -2936 110454 586860 110476
rect -2936 110218 -1814 110454
rect -1578 110218 986 110454
rect 1222 110218 262170 110454
rect 262406 110218 288986 110454
rect 289222 110218 554298 110454
rect 554534 110218 576986 110454
rect 577222 110218 585502 110454
rect 585738 110218 586860 110454
rect -2936 110134 586860 110218
rect -2936 109898 -1814 110134
rect -1578 109898 986 110134
rect 1222 109898 262170 110134
rect 262406 109898 288986 110134
rect 289222 109898 554298 110134
rect 554534 109898 576986 110134
rect 577222 109898 585502 110134
rect 585738 109898 586860 110134
rect -2936 109876 586860 109898
rect -1996 109874 -1396 109876
rect 804 109874 1404 109876
rect 262128 109874 262448 109876
rect 288804 109874 289404 109876
rect 554256 109874 554576 109876
rect 576804 109874 577404 109876
rect 585320 109874 585920 109876
rect -2936 92476 -2336 92478
rect 18804 92476 19404 92478
rect 246768 92476 247088 92478
rect 270804 92476 271404 92478
rect 306804 92476 307404 92478
rect 538896 92476 539216 92478
rect 586260 92476 586860 92478
rect -2936 92454 586860 92476
rect -2936 92218 -2754 92454
rect -2518 92218 18986 92454
rect 19222 92218 246810 92454
rect 247046 92218 270986 92454
rect 271222 92218 306986 92454
rect 307222 92218 538938 92454
rect 539174 92218 586442 92454
rect 586678 92218 586860 92454
rect -2936 92134 586860 92218
rect -2936 91898 -2754 92134
rect -2518 91898 18986 92134
rect 19222 91898 246810 92134
rect 247046 91898 270986 92134
rect 271222 91898 306986 92134
rect 307222 91898 538938 92134
rect 539174 91898 586442 92134
rect 586678 91898 586860 92134
rect -2936 91876 586860 91898
rect -2936 91874 -2336 91876
rect 18804 91874 19404 91876
rect 246768 91874 247088 91876
rect 270804 91874 271404 91876
rect 306804 91874 307404 91876
rect 538896 91874 539216 91876
rect 586260 91874 586860 91876
rect -1996 74476 -1396 74478
rect 804 74476 1404 74478
rect 288804 74476 289404 74478
rect 576804 74476 577404 74478
rect 585320 74476 585920 74478
rect -2936 74454 586860 74476
rect -2936 74218 -1814 74454
rect -1578 74218 986 74454
rect 1222 74218 288986 74454
rect 289222 74218 576986 74454
rect 577222 74218 585502 74454
rect 585738 74218 586860 74454
rect -2936 74134 586860 74218
rect -2936 73898 -1814 74134
rect -1578 73898 986 74134
rect 1222 73898 288986 74134
rect 289222 73898 576986 74134
rect 577222 73898 585502 74134
rect 585738 73898 586860 74134
rect -2936 73876 586860 73898
rect -1996 73874 -1396 73876
rect 804 73874 1404 73876
rect 288804 73874 289404 73876
rect 576804 73874 577404 73876
rect 585320 73874 585920 73876
rect -2936 56476 -2336 56478
rect 18804 56476 19404 56478
rect 54804 56476 55404 56478
rect 90804 56476 91404 56478
rect 126804 56476 127404 56478
rect 162804 56476 163404 56478
rect 198804 56476 199404 56478
rect 234804 56476 235404 56478
rect 270804 56476 271404 56478
rect 306804 56476 307404 56478
rect 342804 56476 343404 56478
rect 378804 56476 379404 56478
rect 414804 56476 415404 56478
rect 450804 56476 451404 56478
rect 486804 56476 487404 56478
rect 522804 56476 523404 56478
rect 558804 56476 559404 56478
rect 586260 56476 586860 56478
rect -2936 56454 586860 56476
rect -2936 56218 -2754 56454
rect -2518 56218 18986 56454
rect 19222 56218 54986 56454
rect 55222 56218 90986 56454
rect 91222 56218 126986 56454
rect 127222 56218 162986 56454
rect 163222 56218 198986 56454
rect 199222 56218 234986 56454
rect 235222 56218 270986 56454
rect 271222 56218 306986 56454
rect 307222 56218 342986 56454
rect 343222 56218 378986 56454
rect 379222 56218 414986 56454
rect 415222 56218 450986 56454
rect 451222 56218 486986 56454
rect 487222 56218 522986 56454
rect 523222 56218 558986 56454
rect 559222 56218 586442 56454
rect 586678 56218 586860 56454
rect -2936 56134 586860 56218
rect -2936 55898 -2754 56134
rect -2518 55898 18986 56134
rect 19222 55898 54986 56134
rect 55222 55898 90986 56134
rect 91222 55898 126986 56134
rect 127222 55898 162986 56134
rect 163222 55898 198986 56134
rect 199222 55898 234986 56134
rect 235222 55898 270986 56134
rect 271222 55898 306986 56134
rect 307222 55898 342986 56134
rect 343222 55898 378986 56134
rect 379222 55898 414986 56134
rect 415222 55898 450986 56134
rect 451222 55898 486986 56134
rect 487222 55898 522986 56134
rect 523222 55898 558986 56134
rect 559222 55898 586442 56134
rect 586678 55898 586860 56134
rect -2936 55876 586860 55898
rect -2936 55874 -2336 55876
rect 18804 55874 19404 55876
rect 54804 55874 55404 55876
rect 90804 55874 91404 55876
rect 126804 55874 127404 55876
rect 162804 55874 163404 55876
rect 198804 55874 199404 55876
rect 234804 55874 235404 55876
rect 270804 55874 271404 55876
rect 306804 55874 307404 55876
rect 342804 55874 343404 55876
rect 378804 55874 379404 55876
rect 414804 55874 415404 55876
rect 450804 55874 451404 55876
rect 486804 55874 487404 55876
rect 522804 55874 523404 55876
rect 558804 55874 559404 55876
rect 586260 55874 586860 55876
rect -1996 38476 -1396 38478
rect 804 38476 1404 38478
rect 36804 38476 37404 38478
rect 72804 38476 73404 38478
rect 108804 38476 109404 38478
rect 144804 38476 145404 38478
rect 180804 38476 181404 38478
rect 216804 38476 217404 38478
rect 252804 38476 253404 38478
rect 288804 38476 289404 38478
rect 324804 38476 325404 38478
rect 360804 38476 361404 38478
rect 396804 38476 397404 38478
rect 432804 38476 433404 38478
rect 468804 38476 469404 38478
rect 504804 38476 505404 38478
rect 540804 38476 541404 38478
rect 576804 38476 577404 38478
rect 585320 38476 585920 38478
rect -2936 38454 586860 38476
rect -2936 38218 -1814 38454
rect -1578 38218 986 38454
rect 1222 38218 36986 38454
rect 37222 38218 72986 38454
rect 73222 38218 108986 38454
rect 109222 38218 144986 38454
rect 145222 38218 180986 38454
rect 181222 38218 216986 38454
rect 217222 38218 252986 38454
rect 253222 38218 288986 38454
rect 289222 38218 324986 38454
rect 325222 38218 360986 38454
rect 361222 38218 396986 38454
rect 397222 38218 432986 38454
rect 433222 38218 468986 38454
rect 469222 38218 504986 38454
rect 505222 38218 540986 38454
rect 541222 38218 576986 38454
rect 577222 38218 585502 38454
rect 585738 38218 586860 38454
rect -2936 38134 586860 38218
rect -2936 37898 -1814 38134
rect -1578 37898 986 38134
rect 1222 37898 36986 38134
rect 37222 37898 72986 38134
rect 73222 37898 108986 38134
rect 109222 37898 144986 38134
rect 145222 37898 180986 38134
rect 181222 37898 216986 38134
rect 217222 37898 252986 38134
rect 253222 37898 288986 38134
rect 289222 37898 324986 38134
rect 325222 37898 360986 38134
rect 361222 37898 396986 38134
rect 397222 37898 432986 38134
rect 433222 37898 468986 38134
rect 469222 37898 504986 38134
rect 505222 37898 540986 38134
rect 541222 37898 576986 38134
rect 577222 37898 585502 38134
rect 585738 37898 586860 38134
rect -2936 37876 586860 37898
rect -1996 37874 -1396 37876
rect 804 37874 1404 37876
rect 36804 37874 37404 37876
rect 72804 37874 73404 37876
rect 108804 37874 109404 37876
rect 144804 37874 145404 37876
rect 180804 37874 181404 37876
rect 216804 37874 217404 37876
rect 252804 37874 253404 37876
rect 288804 37874 289404 37876
rect 324804 37874 325404 37876
rect 360804 37874 361404 37876
rect 396804 37874 397404 37876
rect 432804 37874 433404 37876
rect 468804 37874 469404 37876
rect 504804 37874 505404 37876
rect 540804 37874 541404 37876
rect 576804 37874 577404 37876
rect 585320 37874 585920 37876
rect -2936 20476 -2336 20478
rect 18804 20476 19404 20478
rect 54804 20476 55404 20478
rect 90804 20476 91404 20478
rect 126804 20476 127404 20478
rect 162804 20476 163404 20478
rect 198804 20476 199404 20478
rect 234804 20476 235404 20478
rect 270804 20476 271404 20478
rect 306804 20476 307404 20478
rect 342804 20476 343404 20478
rect 378804 20476 379404 20478
rect 414804 20476 415404 20478
rect 450804 20476 451404 20478
rect 486804 20476 487404 20478
rect 522804 20476 523404 20478
rect 558804 20476 559404 20478
rect 586260 20476 586860 20478
rect -2936 20454 586860 20476
rect -2936 20218 -2754 20454
rect -2518 20218 18986 20454
rect 19222 20218 54986 20454
rect 55222 20218 90986 20454
rect 91222 20218 126986 20454
rect 127222 20218 162986 20454
rect 163222 20218 198986 20454
rect 199222 20218 234986 20454
rect 235222 20218 270986 20454
rect 271222 20218 306986 20454
rect 307222 20218 342986 20454
rect 343222 20218 378986 20454
rect 379222 20218 414986 20454
rect 415222 20218 450986 20454
rect 451222 20218 486986 20454
rect 487222 20218 522986 20454
rect 523222 20218 558986 20454
rect 559222 20218 586442 20454
rect 586678 20218 586860 20454
rect -2936 20134 586860 20218
rect -2936 19898 -2754 20134
rect -2518 19898 18986 20134
rect 19222 19898 54986 20134
rect 55222 19898 90986 20134
rect 91222 19898 126986 20134
rect 127222 19898 162986 20134
rect 163222 19898 198986 20134
rect 199222 19898 234986 20134
rect 235222 19898 270986 20134
rect 271222 19898 306986 20134
rect 307222 19898 342986 20134
rect 343222 19898 378986 20134
rect 379222 19898 414986 20134
rect 415222 19898 450986 20134
rect 451222 19898 486986 20134
rect 487222 19898 522986 20134
rect 523222 19898 558986 20134
rect 559222 19898 586442 20134
rect 586678 19898 586860 20134
rect -2936 19876 586860 19898
rect -2936 19874 -2336 19876
rect 18804 19874 19404 19876
rect 54804 19874 55404 19876
rect 90804 19874 91404 19876
rect 126804 19874 127404 19876
rect 162804 19874 163404 19876
rect 198804 19874 199404 19876
rect 234804 19874 235404 19876
rect 270804 19874 271404 19876
rect 306804 19874 307404 19876
rect 342804 19874 343404 19876
rect 378804 19874 379404 19876
rect 414804 19874 415404 19876
rect 450804 19874 451404 19876
rect 486804 19874 487404 19876
rect 522804 19874 523404 19876
rect 558804 19874 559404 19876
rect 586260 19874 586860 19876
rect -1996 2476 -1396 2478
rect 804 2476 1404 2478
rect 36804 2476 37404 2478
rect 72804 2476 73404 2478
rect 108804 2476 109404 2478
rect 144804 2476 145404 2478
rect 180804 2476 181404 2478
rect 216804 2476 217404 2478
rect 252804 2476 253404 2478
rect 288804 2476 289404 2478
rect 324804 2476 325404 2478
rect 360804 2476 361404 2478
rect 396804 2476 397404 2478
rect 432804 2476 433404 2478
rect 468804 2476 469404 2478
rect 504804 2476 505404 2478
rect 540804 2476 541404 2478
rect 576804 2476 577404 2478
rect 585320 2476 585920 2478
rect -2936 2454 586860 2476
rect -2936 2218 -1814 2454
rect -1578 2218 986 2454
rect 1222 2218 36986 2454
rect 37222 2218 72986 2454
rect 73222 2218 108986 2454
rect 109222 2218 144986 2454
rect 145222 2218 180986 2454
rect 181222 2218 216986 2454
rect 217222 2218 252986 2454
rect 253222 2218 288986 2454
rect 289222 2218 324986 2454
rect 325222 2218 360986 2454
rect 361222 2218 396986 2454
rect 397222 2218 432986 2454
rect 433222 2218 468986 2454
rect 469222 2218 504986 2454
rect 505222 2218 540986 2454
rect 541222 2218 576986 2454
rect 577222 2218 585502 2454
rect 585738 2218 586860 2454
rect -2936 2134 586860 2218
rect -2936 1898 -1814 2134
rect -1578 1898 986 2134
rect 1222 1898 36986 2134
rect 37222 1898 72986 2134
rect 73222 1898 108986 2134
rect 109222 1898 144986 2134
rect 145222 1898 180986 2134
rect 181222 1898 216986 2134
rect 217222 1898 252986 2134
rect 253222 1898 288986 2134
rect 289222 1898 324986 2134
rect 325222 1898 360986 2134
rect 361222 1898 396986 2134
rect 397222 1898 432986 2134
rect 433222 1898 468986 2134
rect 469222 1898 504986 2134
rect 505222 1898 540986 2134
rect 541222 1898 576986 2134
rect 577222 1898 585502 2134
rect 585738 1898 586860 2134
rect -2936 1876 586860 1898
rect -1996 1874 -1396 1876
rect 804 1874 1404 1876
rect 36804 1874 37404 1876
rect 72804 1874 73404 1876
rect 108804 1874 109404 1876
rect 144804 1874 145404 1876
rect 180804 1874 181404 1876
rect 216804 1874 217404 1876
rect 252804 1874 253404 1876
rect 288804 1874 289404 1876
rect 324804 1874 325404 1876
rect 360804 1874 361404 1876
rect 396804 1874 397404 1876
rect 432804 1874 433404 1876
rect 468804 1874 469404 1876
rect 504804 1874 505404 1876
rect 540804 1874 541404 1876
rect 576804 1874 577404 1876
rect 585320 1874 585920 1876
rect -1996 -324 -1396 -322
rect 804 -324 1404 -322
rect 36804 -324 37404 -322
rect 72804 -324 73404 -322
rect 108804 -324 109404 -322
rect 144804 -324 145404 -322
rect 180804 -324 181404 -322
rect 216804 -324 217404 -322
rect 252804 -324 253404 -322
rect 288804 -324 289404 -322
rect 324804 -324 325404 -322
rect 360804 -324 361404 -322
rect 396804 -324 397404 -322
rect 432804 -324 433404 -322
rect 468804 -324 469404 -322
rect 504804 -324 505404 -322
rect 540804 -324 541404 -322
rect 576804 -324 577404 -322
rect 585320 -324 585920 -322
rect -1996 -346 585920 -324
rect -1996 -582 -1814 -346
rect -1578 -582 986 -346
rect 1222 -582 36986 -346
rect 37222 -582 72986 -346
rect 73222 -582 108986 -346
rect 109222 -582 144986 -346
rect 145222 -582 180986 -346
rect 181222 -582 216986 -346
rect 217222 -582 252986 -346
rect 253222 -582 288986 -346
rect 289222 -582 324986 -346
rect 325222 -582 360986 -346
rect 361222 -582 396986 -346
rect 397222 -582 432986 -346
rect 433222 -582 468986 -346
rect 469222 -582 504986 -346
rect 505222 -582 540986 -346
rect 541222 -582 576986 -346
rect 577222 -582 585502 -346
rect 585738 -582 585920 -346
rect -1996 -666 585920 -582
rect -1996 -902 -1814 -666
rect -1578 -902 986 -666
rect 1222 -902 36986 -666
rect 37222 -902 72986 -666
rect 73222 -902 108986 -666
rect 109222 -902 144986 -666
rect 145222 -902 180986 -666
rect 181222 -902 216986 -666
rect 217222 -902 252986 -666
rect 253222 -902 288986 -666
rect 289222 -902 324986 -666
rect 325222 -902 360986 -666
rect 361222 -902 396986 -666
rect 397222 -902 432986 -666
rect 433222 -902 468986 -666
rect 469222 -902 504986 -666
rect 505222 -902 540986 -666
rect 541222 -902 576986 -666
rect 577222 -902 585502 -666
rect 585738 -902 585920 -666
rect -1996 -924 585920 -902
rect -1996 -926 -1396 -924
rect 804 -926 1404 -924
rect 36804 -926 37404 -924
rect 72804 -926 73404 -924
rect 108804 -926 109404 -924
rect 144804 -926 145404 -924
rect 180804 -926 181404 -924
rect 216804 -926 217404 -924
rect 252804 -926 253404 -924
rect 288804 -926 289404 -924
rect 324804 -926 325404 -924
rect 360804 -926 361404 -924
rect 396804 -926 397404 -924
rect 432804 -926 433404 -924
rect 468804 -926 469404 -924
rect 504804 -926 505404 -924
rect 540804 -926 541404 -924
rect 576804 -926 577404 -924
rect 585320 -926 585920 -924
rect -2936 -1264 -2336 -1262
rect 18804 -1264 19404 -1262
rect 54804 -1264 55404 -1262
rect 90804 -1264 91404 -1262
rect 126804 -1264 127404 -1262
rect 162804 -1264 163404 -1262
rect 198804 -1264 199404 -1262
rect 234804 -1264 235404 -1262
rect 270804 -1264 271404 -1262
rect 306804 -1264 307404 -1262
rect 342804 -1264 343404 -1262
rect 378804 -1264 379404 -1262
rect 414804 -1264 415404 -1262
rect 450804 -1264 451404 -1262
rect 486804 -1264 487404 -1262
rect 522804 -1264 523404 -1262
rect 558804 -1264 559404 -1262
rect 586260 -1264 586860 -1262
rect -2936 -1286 586860 -1264
rect -2936 -1522 -2754 -1286
rect -2518 -1522 18986 -1286
rect 19222 -1522 54986 -1286
rect 55222 -1522 90986 -1286
rect 91222 -1522 126986 -1286
rect 127222 -1522 162986 -1286
rect 163222 -1522 198986 -1286
rect 199222 -1522 234986 -1286
rect 235222 -1522 270986 -1286
rect 271222 -1522 306986 -1286
rect 307222 -1522 342986 -1286
rect 343222 -1522 378986 -1286
rect 379222 -1522 414986 -1286
rect 415222 -1522 450986 -1286
rect 451222 -1522 486986 -1286
rect 487222 -1522 522986 -1286
rect 523222 -1522 558986 -1286
rect 559222 -1522 586442 -1286
rect 586678 -1522 586860 -1286
rect -2936 -1606 586860 -1522
rect -2936 -1842 -2754 -1606
rect -2518 -1842 18986 -1606
rect 19222 -1842 54986 -1606
rect 55222 -1842 90986 -1606
rect 91222 -1842 126986 -1606
rect 127222 -1842 162986 -1606
rect 163222 -1842 198986 -1606
rect 199222 -1842 234986 -1606
rect 235222 -1842 270986 -1606
rect 271222 -1842 306986 -1606
rect 307222 -1842 342986 -1606
rect 343222 -1842 378986 -1606
rect 379222 -1842 414986 -1606
rect 415222 -1842 450986 -1606
rect 451222 -1842 486986 -1606
rect 487222 -1842 522986 -1606
rect 523222 -1842 558986 -1606
rect 559222 -1842 586442 -1606
rect 586678 -1842 586860 -1606
rect -2936 -1864 586860 -1842
rect -2936 -1866 -2336 -1864
rect 18804 -1866 19404 -1864
rect 54804 -1866 55404 -1864
rect 90804 -1866 91404 -1864
rect 126804 -1866 127404 -1864
rect 162804 -1866 163404 -1864
rect 198804 -1866 199404 -1864
rect 234804 -1866 235404 -1864
rect 270804 -1866 271404 -1864
rect 306804 -1866 307404 -1864
rect 342804 -1866 343404 -1864
rect 378804 -1866 379404 -1864
rect 414804 -1866 415404 -1864
rect 450804 -1866 451404 -1864
rect 486804 -1866 487404 -1864
rect 522804 -1866 523404 -1864
rect 558804 -1866 559404 -1864
rect 586260 -1866 586860 -1864
rect -3876 -2204 -3276 -2202
rect 587200 -2204 587800 -2202
rect -3876 -2226 587800 -2204
rect -3876 -2462 -3694 -2226
rect -3458 -2462 587382 -2226
rect 587618 -2462 587800 -2226
rect -3876 -2546 587800 -2462
rect -3876 -2782 -3694 -2546
rect -3458 -2782 587382 -2546
rect 587618 -2782 587800 -2546
rect -3876 -2804 587800 -2782
rect -3876 -2806 -3276 -2804
rect 587200 -2806 587800 -2804
rect -4816 -3144 -4216 -3142
rect 588140 -3144 588740 -3142
rect -4816 -3166 588740 -3144
rect -4816 -3402 -4634 -3166
rect -4398 -3402 588322 -3166
rect 588558 -3402 588740 -3166
rect -4816 -3486 588740 -3402
rect -4816 -3722 -4634 -3486
rect -4398 -3722 588322 -3486
rect 588558 -3722 588740 -3486
rect -4816 -3744 588740 -3722
rect -4816 -3746 -4216 -3744
rect 588140 -3746 588740 -3744
rect -5756 -4084 -5156 -4082
rect 589080 -4084 589680 -4082
rect -5756 -4106 589680 -4084
rect -5756 -4342 -5574 -4106
rect -5338 -4342 589262 -4106
rect 589498 -4342 589680 -4106
rect -5756 -4426 589680 -4342
rect -5756 -4662 -5574 -4426
rect -5338 -4662 589262 -4426
rect 589498 -4662 589680 -4426
rect -5756 -4684 589680 -4662
rect -5756 -4686 -5156 -4684
rect 589080 -4686 589680 -4684
rect -6696 -5024 -6096 -5022
rect 590020 -5024 590620 -5022
rect -6696 -5046 590620 -5024
rect -6696 -5282 -6514 -5046
rect -6278 -5282 590202 -5046
rect 590438 -5282 590620 -5046
rect -6696 -5366 590620 -5282
rect -6696 -5602 -6514 -5366
rect -6278 -5602 590202 -5366
rect 590438 -5602 590620 -5366
rect -6696 -5624 590620 -5602
rect -6696 -5626 -6096 -5624
rect 590020 -5626 590620 -5624
rect -7636 -5964 -7036 -5962
rect 590960 -5964 591560 -5962
rect -7636 -5986 591560 -5964
rect -7636 -6222 -7454 -5986
rect -7218 -6222 591142 -5986
rect 591378 -6222 591560 -5986
rect -7636 -6306 591560 -6222
rect -7636 -6542 -7454 -6306
rect -7218 -6542 591142 -6306
rect 591378 -6542 591560 -6306
rect -7636 -6564 591560 -6542
rect -7636 -6566 -7036 -6564
rect 590960 -6566 591560 -6564
rect -8576 -6904 -7976 -6902
rect 591900 -6904 592500 -6902
rect -8576 -6926 592500 -6904
rect -8576 -7162 -8394 -6926
rect -8158 -7162 592082 -6926
rect 592318 -7162 592500 -6926
rect -8576 -7246 592500 -7162
rect -8576 -7482 -8394 -7246
rect -8158 -7482 592082 -7246
rect 592318 -7482 592500 -7246
rect -8576 -7504 592500 -7482
rect -8576 -7506 -7976 -7504
rect 591900 -7506 592500 -7504
use decred_hash_macro  decred_hash_block3
timestamp 1608074288
transform -1 0 558784 0 -1 583916
box 0 0 240000 200000
use decred_hash_macro  decred_hash_block2
timestamp 1608074288
transform -1 0 266656 0 -1 583916
box 0 0 240000 200000
use decred_hash_macro  decred_hash_block1
timestamp 1608074288
transform -1 0 558784 0 -1 273600
box 0 0 240000 200000
use decred_hash_macro  decred_hash_block0
timestamp 1608074288
transform -1 0 266656 0 -1 273600
box 0 0 240000 200000
use decred_controller  decred_controller_block
timestamp 1608074288
transform -1 0 312000 0 -1 355560
box 0 0 40000 40000
<< labels >>
rlabel metal3 s 583520 5796 584960 6036 6 analog_io[0]
port 0 nsew default bidirectional
rlabel metal3 s 583520 474996 584960 475236 6 analog_io[10]
port 1 nsew default bidirectional
rlabel metal3 s 583520 521916 584960 522156 6 analog_io[11]
port 2 nsew default bidirectional
rlabel metal3 s 583520 568836 584960 569076 6 analog_io[12]
port 3 nsew default bidirectional
rlabel metal3 s 583520 615756 584960 615996 6 analog_io[13]
port 4 nsew default bidirectional
rlabel metal3 s 583520 662676 584960 662916 6 analog_io[14]
port 5 nsew default bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[15]
port 6 nsew default bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[16]
port 7 nsew default bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[17]
port 8 nsew default bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[18]
port 9 nsew default bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[19]
port 10 nsew default bidirectional
rlabel metal3 s 583520 52716 584960 52956 6 analog_io[1]
port 11 nsew default bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[20]
port 12 nsew default bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[21]
port 13 nsew default bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[22]
port 14 nsew default bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[23]
port 15 nsew default bidirectional
rlabel metal3 s -960 696540 480 696780 4 analog_io[24]
port 16 nsew default bidirectional
rlabel metal3 s -960 639012 480 639252 4 analog_io[25]
port 17 nsew default bidirectional
rlabel metal3 s -960 581620 480 581860 4 analog_io[26]
port 18 nsew default bidirectional
rlabel metal3 s -960 524092 480 524332 4 analog_io[27]
port 19 nsew default bidirectional
rlabel metal3 s -960 466700 480 466940 4 analog_io[28]
port 20 nsew default bidirectional
rlabel metal3 s -960 409172 480 409412 4 analog_io[29]
port 21 nsew default bidirectional
rlabel metal3 s 583520 99636 584960 99876 6 analog_io[2]
port 22 nsew default bidirectional
rlabel metal3 s -960 351780 480 352020 4 analog_io[30]
port 23 nsew default bidirectional
rlabel metal3 s 583520 146556 584960 146796 6 analog_io[3]
port 24 nsew default bidirectional
rlabel metal3 s 583520 193476 584960 193716 6 analog_io[4]
port 25 nsew default bidirectional
rlabel metal3 s 583520 240396 584960 240636 6 analog_io[5]
port 26 nsew default bidirectional
rlabel metal3 s 583520 287316 584960 287556 6 analog_io[6]
port 27 nsew default bidirectional
rlabel metal3 s 583520 334236 584960 334476 6 analog_io[7]
port 28 nsew default bidirectional
rlabel metal3 s 583520 381156 584960 381396 6 analog_io[8]
port 29 nsew default bidirectional
rlabel metal3 s 583520 428076 584960 428316 6 analog_io[9]
port 30 nsew default bidirectional
rlabel metal3 s 583520 17492 584960 17732 6 io_in[0]
port 31 nsew default input
rlabel metal3 s 583520 486692 584960 486932 6 io_in[10]
port 32 nsew default input
rlabel metal3 s 583520 533748 584960 533988 6 io_in[11]
port 33 nsew default input
rlabel metal3 s 583520 580668 584960 580908 6 io_in[12]
port 34 nsew default input
rlabel metal3 s 583520 627588 584960 627828 6 io_in[13]
port 35 nsew default input
rlabel metal3 s 583520 674508 584960 674748 6 io_in[14]
port 36 nsew default input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 37 nsew default input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 38 nsew default input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 39 nsew default input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 40 nsew default input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 41 nsew default input
rlabel metal3 s 583520 64412 584960 64652 6 io_in[1]
port 42 nsew default input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 43 nsew default input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 44 nsew default input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 45 nsew default input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 46 nsew default input
rlabel metal3 s -960 682124 480 682364 4 io_in[24]
port 47 nsew default input
rlabel metal3 s -960 624732 480 624972 4 io_in[25]
port 48 nsew default input
rlabel metal3 s -960 567204 480 567444 4 io_in[26]
port 49 nsew default input
rlabel metal3 s -960 509812 480 510052 4 io_in[27]
port 50 nsew default input
rlabel metal3 s -960 452284 480 452524 4 io_in[28]
port 51 nsew default input
rlabel metal3 s -960 394892 480 395132 4 io_in[29]
port 52 nsew default input
rlabel metal3 s 583520 111332 584960 111572 6 io_in[2]
port 53 nsew default input
rlabel metal3 s -960 337364 480 337604 4 io_in[30]
port 54 nsew default input
rlabel metal3 s -960 294252 480 294492 4 io_in[31]
port 55 nsew default input
rlabel metal3 s -960 251140 480 251380 4 io_in[32]
port 56 nsew default input
rlabel metal3 s -960 208028 480 208268 4 io_in[33]
port 57 nsew default input
rlabel metal3 s -960 164916 480 165156 4 io_in[34]
port 58 nsew default input
rlabel metal3 s -960 121940 480 122180 4 io_in[35]
port 59 nsew default input
rlabel metal3 s -960 78828 480 79068 4 io_in[36]
port 60 nsew default input
rlabel metal3 s -960 35716 480 35956 4 io_in[37]
port 61 nsew default input
rlabel metal3 s 583520 158252 584960 158492 6 io_in[3]
port 62 nsew default input
rlabel metal3 s 583520 205172 584960 205412 6 io_in[4]
port 63 nsew default input
rlabel metal3 s 583520 252092 584960 252332 6 io_in[5]
port 64 nsew default input
rlabel metal3 s 583520 299012 584960 299252 6 io_in[6]
port 65 nsew default input
rlabel metal3 s 583520 345932 584960 346172 6 io_in[7]
port 66 nsew default input
rlabel metal3 s 583520 392852 584960 393092 6 io_in[8]
port 67 nsew default input
rlabel metal3 s 583520 439772 584960 440012 6 io_in[9]
port 68 nsew default input
rlabel metal3 s 583520 40884 584960 41124 6 io_oeb[0]
port 69 nsew default tristate
rlabel metal3 s 583520 87804 584960 88044 6 io_oeb[1]
port 70 nsew default tristate
rlabel metal3 s -960 366060 480 366300 4 io_oeb[29]
port 71 nsew default tristate
rlabel metal3 s 583520 134724 584960 134964 6 io_oeb[2]
port 72 nsew default tristate
rlabel metal3 s -960 308668 480 308908 4 io_oeb[30]
port 73 nsew default tristate
rlabel metal3 s -960 265556 480 265796 4 io_oeb[31]
port 74 nsew default tristate
rlabel metal3 s -960 222444 480 222684 4 io_oeb[32]
port 75 nsew default tristate
rlabel metal3 s -960 179332 480 179572 4 io_oeb[33]
port 76 nsew default tristate
rlabel metal3 s -960 136220 480 136460 4 io_oeb[34]
port 77 nsew default tristate
rlabel metal3 s -960 93108 480 93348 4 io_oeb[35]
port 78 nsew default tristate
rlabel metal3 s -960 49996 480 50236 4 io_oeb[36]
port 79 nsew default tristate
rlabel metal3 s -960 7020 480 7260 4 io_oeb[37]
port 80 nsew default tristate
rlabel metal3 s 583520 181780 584960 182020 6 io_oeb[3]
port 81 nsew default tristate
rlabel metal3 s 583520 228700 584960 228940 6 io_oeb[4]
port 82 nsew default tristate
rlabel metal3 s 583520 275620 584960 275860 6 io_oeb[5]
port 83 nsew default tristate
rlabel metal3 s 583520 322540 584960 322780 6 io_oeb[6]
port 84 nsew default tristate
rlabel metal3 s 583520 369460 584960 369700 6 io_oeb[7]
port 85 nsew default tristate
rlabel metal3 s 583520 29188 584960 29428 6 io_out[0]
port 86 nsew default tristate
rlabel metal3 s 583520 498524 584960 498764 6 io_out[10]
port 87 nsew default tristate
rlabel metal3 s 583520 545444 584960 545684 6 io_out[11]
port 88 nsew default tristate
rlabel metal3 s 583520 592364 584960 592604 6 io_out[12]
port 89 nsew default tristate
rlabel metal3 s 583520 639284 584960 639524 6 io_out[13]
port 90 nsew default tristate
rlabel metal3 s 583520 686204 584960 686444 6 io_out[14]
port 91 nsew default tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 92 nsew default tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 93 nsew default tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 94 nsew default tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 95 nsew default tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 96 nsew default tristate
rlabel metal3 s 583520 76108 584960 76348 6 io_out[1]
port 97 nsew default tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 98 nsew default tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 99 nsew default tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 100 nsew default tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 101 nsew default tristate
rlabel metal3 s -960 667844 480 668084 4 io_out[24]
port 102 nsew default tristate
rlabel metal3 s -960 610316 480 610556 4 io_out[25]
port 103 nsew default tristate
rlabel metal3 s -960 552924 480 553164 4 io_out[26]
port 104 nsew default tristate
rlabel metal3 s -960 495396 480 495636 4 io_out[27]
port 105 nsew default tristate
rlabel metal3 s -960 437868 480 438108 4 io_out[28]
port 106 nsew default tristate
rlabel metal3 s -960 380476 480 380716 4 io_out[29]
port 107 nsew default tristate
rlabel metal3 s 583520 123028 584960 123268 6 io_out[2]
port 108 nsew default tristate
rlabel metal3 s -960 322948 480 323188 4 io_out[30]
port 109 nsew default tristate
rlabel metal3 s -960 279972 480 280212 4 io_out[31]
port 110 nsew default tristate
rlabel metal3 s -960 236860 480 237100 4 io_out[32]
port 111 nsew default tristate
rlabel metal3 s -960 193748 480 193988 4 io_out[33]
port 112 nsew default tristate
rlabel metal3 s -960 150636 480 150876 4 io_out[34]
port 113 nsew default tristate
rlabel metal3 s -960 107524 480 107764 4 io_out[35]
port 114 nsew default tristate
rlabel metal3 s -960 64412 480 64652 4 io_out[36]
port 115 nsew default tristate
rlabel metal3 s -960 21300 480 21540 4 io_out[37]
port 116 nsew default tristate
rlabel metal3 s 583520 169948 584960 170188 6 io_out[3]
port 117 nsew default tristate
rlabel metal3 s 583520 216868 584960 217108 6 io_out[4]
port 118 nsew default tristate
rlabel metal3 s 583520 263788 584960 264028 6 io_out[5]
port 119 nsew default tristate
rlabel metal3 s 583520 310708 584960 310948 6 io_out[6]
port 120 nsew default tristate
rlabel metal3 s 583520 357764 584960 358004 6 io_out[7]
port 121 nsew default tristate
rlabel metal3 s 583520 404684 584960 404924 6 io_out[8]
port 122 nsew default tristate
rlabel metal3 s 583520 451604 584960 451844 6 io_out[9]
port 123 nsew default tristate
rlabel metal2 s 126582 -960 126694 480 8 la_data_in[0]
port 124 nsew default input
rlabel metal2 s 483450 -960 483562 480 8 la_data_in[100]
port 125 nsew default input
rlabel metal2 s 486946 -960 487058 480 8 la_data_in[101]
port 126 nsew default input
rlabel metal2 s 490534 -960 490646 480 8 la_data_in[102]
port 127 nsew default input
rlabel metal2 s 494122 -960 494234 480 8 la_data_in[103]
port 128 nsew default input
rlabel metal2 s 497710 -960 497822 480 8 la_data_in[104]
port 129 nsew default input
rlabel metal2 s 501206 -960 501318 480 8 la_data_in[105]
port 130 nsew default input
rlabel metal2 s 504794 -960 504906 480 8 la_data_in[106]
port 131 nsew default input
rlabel metal2 s 508382 -960 508494 480 8 la_data_in[107]
port 132 nsew default input
rlabel metal2 s 511970 -960 512082 480 8 la_data_in[108]
port 133 nsew default input
rlabel metal2 s 515558 -960 515670 480 8 la_data_in[109]
port 134 nsew default input
rlabel metal2 s 162278 -960 162390 480 8 la_data_in[10]
port 135 nsew default input
rlabel metal2 s 519054 -960 519166 480 8 la_data_in[110]
port 136 nsew default input
rlabel metal2 s 522642 -960 522754 480 8 la_data_in[111]
port 137 nsew default input
rlabel metal2 s 526230 -960 526342 480 8 la_data_in[112]
port 138 nsew default input
rlabel metal2 s 529818 -960 529930 480 8 la_data_in[113]
port 139 nsew default input
rlabel metal2 s 533406 -960 533518 480 8 la_data_in[114]
port 140 nsew default input
rlabel metal2 s 536902 -960 537014 480 8 la_data_in[115]
port 141 nsew default input
rlabel metal2 s 540490 -960 540602 480 8 la_data_in[116]
port 142 nsew default input
rlabel metal2 s 544078 -960 544190 480 8 la_data_in[117]
port 143 nsew default input
rlabel metal2 s 547666 -960 547778 480 8 la_data_in[118]
port 144 nsew default input
rlabel metal2 s 551162 -960 551274 480 8 la_data_in[119]
port 145 nsew default input
rlabel metal2 s 165866 -960 165978 480 8 la_data_in[11]
port 146 nsew default input
rlabel metal2 s 554750 -960 554862 480 8 la_data_in[120]
port 147 nsew default input
rlabel metal2 s 558338 -960 558450 480 8 la_data_in[121]
port 148 nsew default input
rlabel metal2 s 561926 -960 562038 480 8 la_data_in[122]
port 149 nsew default input
rlabel metal2 s 565514 -960 565626 480 8 la_data_in[123]
port 150 nsew default input
rlabel metal2 s 569010 -960 569122 480 8 la_data_in[124]
port 151 nsew default input
rlabel metal2 s 572598 -960 572710 480 8 la_data_in[125]
port 152 nsew default input
rlabel metal2 s 576186 -960 576298 480 8 la_data_in[126]
port 153 nsew default input
rlabel metal2 s 579774 -960 579886 480 8 la_data_in[127]
port 154 nsew default input
rlabel metal2 s 169362 -960 169474 480 8 la_data_in[12]
port 155 nsew default input
rlabel metal2 s 172950 -960 173062 480 8 la_data_in[13]
port 156 nsew default input
rlabel metal2 s 176538 -960 176650 480 8 la_data_in[14]
port 157 nsew default input
rlabel metal2 s 180126 -960 180238 480 8 la_data_in[15]
port 158 nsew default input
rlabel metal2 s 183714 -960 183826 480 8 la_data_in[16]
port 159 nsew default input
rlabel metal2 s 187210 -960 187322 480 8 la_data_in[17]
port 160 nsew default input
rlabel metal2 s 190798 -960 190910 480 8 la_data_in[18]
port 161 nsew default input
rlabel metal2 s 194386 -960 194498 480 8 la_data_in[19]
port 162 nsew default input
rlabel metal2 s 130170 -960 130282 480 8 la_data_in[1]
port 163 nsew default input
rlabel metal2 s 197974 -960 198086 480 8 la_data_in[20]
port 164 nsew default input
rlabel metal2 s 201470 -960 201582 480 8 la_data_in[21]
port 165 nsew default input
rlabel metal2 s 205058 -960 205170 480 8 la_data_in[22]
port 166 nsew default input
rlabel metal2 s 208646 -960 208758 480 8 la_data_in[23]
port 167 nsew default input
rlabel metal2 s 212234 -960 212346 480 8 la_data_in[24]
port 168 nsew default input
rlabel metal2 s 215822 -960 215934 480 8 la_data_in[25]
port 169 nsew default input
rlabel metal2 s 219318 -960 219430 480 8 la_data_in[26]
port 170 nsew default input
rlabel metal2 s 222906 -960 223018 480 8 la_data_in[27]
port 171 nsew default input
rlabel metal2 s 226494 -960 226606 480 8 la_data_in[28]
port 172 nsew default input
rlabel metal2 s 230082 -960 230194 480 8 la_data_in[29]
port 173 nsew default input
rlabel metal2 s 133758 -960 133870 480 8 la_data_in[2]
port 174 nsew default input
rlabel metal2 s 233670 -960 233782 480 8 la_data_in[30]
port 175 nsew default input
rlabel metal2 s 237166 -960 237278 480 8 la_data_in[31]
port 176 nsew default input
rlabel metal2 s 240754 -960 240866 480 8 la_data_in[32]
port 177 nsew default input
rlabel metal2 s 244342 -960 244454 480 8 la_data_in[33]
port 178 nsew default input
rlabel metal2 s 247930 -960 248042 480 8 la_data_in[34]
port 179 nsew default input
rlabel metal2 s 251426 -960 251538 480 8 la_data_in[35]
port 180 nsew default input
rlabel metal2 s 255014 -960 255126 480 8 la_data_in[36]
port 181 nsew default input
rlabel metal2 s 258602 -960 258714 480 8 la_data_in[37]
port 182 nsew default input
rlabel metal2 s 262190 -960 262302 480 8 la_data_in[38]
port 183 nsew default input
rlabel metal2 s 265778 -960 265890 480 8 la_data_in[39]
port 184 nsew default input
rlabel metal2 s 137254 -960 137366 480 8 la_data_in[3]
port 185 nsew default input
rlabel metal2 s 269274 -960 269386 480 8 la_data_in[40]
port 186 nsew default input
rlabel metal2 s 272862 -960 272974 480 8 la_data_in[41]
port 187 nsew default input
rlabel metal2 s 276450 -960 276562 480 8 la_data_in[42]
port 188 nsew default input
rlabel metal2 s 280038 -960 280150 480 8 la_data_in[43]
port 189 nsew default input
rlabel metal2 s 283626 -960 283738 480 8 la_data_in[44]
port 190 nsew default input
rlabel metal2 s 287122 -960 287234 480 8 la_data_in[45]
port 191 nsew default input
rlabel metal2 s 290710 -960 290822 480 8 la_data_in[46]
port 192 nsew default input
rlabel metal2 s 294298 -960 294410 480 8 la_data_in[47]
port 193 nsew default input
rlabel metal2 s 297886 -960 297998 480 8 la_data_in[48]
port 194 nsew default input
rlabel metal2 s 301382 -960 301494 480 8 la_data_in[49]
port 195 nsew default input
rlabel metal2 s 140842 -960 140954 480 8 la_data_in[4]
port 196 nsew default input
rlabel metal2 s 304970 -960 305082 480 8 la_data_in[50]
port 197 nsew default input
rlabel metal2 s 308558 -960 308670 480 8 la_data_in[51]
port 198 nsew default input
rlabel metal2 s 312146 -960 312258 480 8 la_data_in[52]
port 199 nsew default input
rlabel metal2 s 315734 -960 315846 480 8 la_data_in[53]
port 200 nsew default input
rlabel metal2 s 319230 -960 319342 480 8 la_data_in[54]
port 201 nsew default input
rlabel metal2 s 322818 -960 322930 480 8 la_data_in[55]
port 202 nsew default input
rlabel metal2 s 326406 -960 326518 480 8 la_data_in[56]
port 203 nsew default input
rlabel metal2 s 329994 -960 330106 480 8 la_data_in[57]
port 204 nsew default input
rlabel metal2 s 333582 -960 333694 480 8 la_data_in[58]
port 205 nsew default input
rlabel metal2 s 337078 -960 337190 480 8 la_data_in[59]
port 206 nsew default input
rlabel metal2 s 144430 -960 144542 480 8 la_data_in[5]
port 207 nsew default input
rlabel metal2 s 340666 -960 340778 480 8 la_data_in[60]
port 208 nsew default input
rlabel metal2 s 344254 -960 344366 480 8 la_data_in[61]
port 209 nsew default input
rlabel metal2 s 347842 -960 347954 480 8 la_data_in[62]
port 210 nsew default input
rlabel metal2 s 351338 -960 351450 480 8 la_data_in[63]
port 211 nsew default input
rlabel metal2 s 354926 -960 355038 480 8 la_data_in[64]
port 212 nsew default input
rlabel metal2 s 358514 -960 358626 480 8 la_data_in[65]
port 213 nsew default input
rlabel metal2 s 362102 -960 362214 480 8 la_data_in[66]
port 214 nsew default input
rlabel metal2 s 365690 -960 365802 480 8 la_data_in[67]
port 215 nsew default input
rlabel metal2 s 369186 -960 369298 480 8 la_data_in[68]
port 216 nsew default input
rlabel metal2 s 372774 -960 372886 480 8 la_data_in[69]
port 217 nsew default input
rlabel metal2 s 148018 -960 148130 480 8 la_data_in[6]
port 218 nsew default input
rlabel metal2 s 376362 -960 376474 480 8 la_data_in[70]
port 219 nsew default input
rlabel metal2 s 379950 -960 380062 480 8 la_data_in[71]
port 220 nsew default input
rlabel metal2 s 383538 -960 383650 480 8 la_data_in[72]
port 221 nsew default input
rlabel metal2 s 387034 -960 387146 480 8 la_data_in[73]
port 222 nsew default input
rlabel metal2 s 390622 -960 390734 480 8 la_data_in[74]
port 223 nsew default input
rlabel metal2 s 394210 -960 394322 480 8 la_data_in[75]
port 224 nsew default input
rlabel metal2 s 397798 -960 397910 480 8 la_data_in[76]
port 225 nsew default input
rlabel metal2 s 401294 -960 401406 480 8 la_data_in[77]
port 226 nsew default input
rlabel metal2 s 404882 -960 404994 480 8 la_data_in[78]
port 227 nsew default input
rlabel metal2 s 408470 -960 408582 480 8 la_data_in[79]
port 228 nsew default input
rlabel metal2 s 151514 -960 151626 480 8 la_data_in[7]
port 229 nsew default input
rlabel metal2 s 412058 -960 412170 480 8 la_data_in[80]
port 230 nsew default input
rlabel metal2 s 415646 -960 415758 480 8 la_data_in[81]
port 231 nsew default input
rlabel metal2 s 419142 -960 419254 480 8 la_data_in[82]
port 232 nsew default input
rlabel metal2 s 422730 -960 422842 480 8 la_data_in[83]
port 233 nsew default input
rlabel metal2 s 426318 -960 426430 480 8 la_data_in[84]
port 234 nsew default input
rlabel metal2 s 429906 -960 430018 480 8 la_data_in[85]
port 235 nsew default input
rlabel metal2 s 433494 -960 433606 480 8 la_data_in[86]
port 236 nsew default input
rlabel metal2 s 436990 -960 437102 480 8 la_data_in[87]
port 237 nsew default input
rlabel metal2 s 440578 -960 440690 480 8 la_data_in[88]
port 238 nsew default input
rlabel metal2 s 444166 -960 444278 480 8 la_data_in[89]
port 239 nsew default input
rlabel metal2 s 155102 -960 155214 480 8 la_data_in[8]
port 240 nsew default input
rlabel metal2 s 447754 -960 447866 480 8 la_data_in[90]
port 241 nsew default input
rlabel metal2 s 451250 -960 451362 480 8 la_data_in[91]
port 242 nsew default input
rlabel metal2 s 454838 -960 454950 480 8 la_data_in[92]
port 243 nsew default input
rlabel metal2 s 458426 -960 458538 480 8 la_data_in[93]
port 244 nsew default input
rlabel metal2 s 462014 -960 462126 480 8 la_data_in[94]
port 245 nsew default input
rlabel metal2 s 465602 -960 465714 480 8 la_data_in[95]
port 246 nsew default input
rlabel metal2 s 469098 -960 469210 480 8 la_data_in[96]
port 247 nsew default input
rlabel metal2 s 472686 -960 472798 480 8 la_data_in[97]
port 248 nsew default input
rlabel metal2 s 476274 -960 476386 480 8 la_data_in[98]
port 249 nsew default input
rlabel metal2 s 479862 -960 479974 480 8 la_data_in[99]
port 250 nsew default input
rlabel metal2 s 158690 -960 158802 480 8 la_data_in[9]
port 251 nsew default input
rlabel metal2 s 127778 -960 127890 480 8 la_data_out[0]
port 252 nsew default tristate
rlabel metal2 s 484554 -960 484666 480 8 la_data_out[100]
port 253 nsew default tristate
rlabel metal2 s 488142 -960 488254 480 8 la_data_out[101]
port 254 nsew default tristate
rlabel metal2 s 491730 -960 491842 480 8 la_data_out[102]
port 255 nsew default tristate
rlabel metal2 s 495318 -960 495430 480 8 la_data_out[103]
port 256 nsew default tristate
rlabel metal2 s 498906 -960 499018 480 8 la_data_out[104]
port 257 nsew default tristate
rlabel metal2 s 502402 -960 502514 480 8 la_data_out[105]
port 258 nsew default tristate
rlabel metal2 s 505990 -960 506102 480 8 la_data_out[106]
port 259 nsew default tristate
rlabel metal2 s 509578 -960 509690 480 8 la_data_out[107]
port 260 nsew default tristate
rlabel metal2 s 513166 -960 513278 480 8 la_data_out[108]
port 261 nsew default tristate
rlabel metal2 s 516754 -960 516866 480 8 la_data_out[109]
port 262 nsew default tristate
rlabel metal2 s 163474 -960 163586 480 8 la_data_out[10]
port 263 nsew default tristate
rlabel metal2 s 520250 -960 520362 480 8 la_data_out[110]
port 264 nsew default tristate
rlabel metal2 s 523838 -960 523950 480 8 la_data_out[111]
port 265 nsew default tristate
rlabel metal2 s 527426 -960 527538 480 8 la_data_out[112]
port 266 nsew default tristate
rlabel metal2 s 531014 -960 531126 480 8 la_data_out[113]
port 267 nsew default tristate
rlabel metal2 s 534510 -960 534622 480 8 la_data_out[114]
port 268 nsew default tristate
rlabel metal2 s 538098 -960 538210 480 8 la_data_out[115]
port 269 nsew default tristate
rlabel metal2 s 541686 -960 541798 480 8 la_data_out[116]
port 270 nsew default tristate
rlabel metal2 s 545274 -960 545386 480 8 la_data_out[117]
port 271 nsew default tristate
rlabel metal2 s 548862 -960 548974 480 8 la_data_out[118]
port 272 nsew default tristate
rlabel metal2 s 552358 -960 552470 480 8 la_data_out[119]
port 273 nsew default tristate
rlabel metal2 s 167062 -960 167174 480 8 la_data_out[11]
port 274 nsew default tristate
rlabel metal2 s 555946 -960 556058 480 8 la_data_out[120]
port 275 nsew default tristate
rlabel metal2 s 559534 -960 559646 480 8 la_data_out[121]
port 276 nsew default tristate
rlabel metal2 s 563122 -960 563234 480 8 la_data_out[122]
port 277 nsew default tristate
rlabel metal2 s 566710 -960 566822 480 8 la_data_out[123]
port 278 nsew default tristate
rlabel metal2 s 570206 -960 570318 480 8 la_data_out[124]
port 279 nsew default tristate
rlabel metal2 s 573794 -960 573906 480 8 la_data_out[125]
port 280 nsew default tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[126]
port 281 nsew default tristate
rlabel metal2 s 580970 -960 581082 480 8 la_data_out[127]
port 282 nsew default tristate
rlabel metal2 s 170558 -960 170670 480 8 la_data_out[12]
port 283 nsew default tristate
rlabel metal2 s 174146 -960 174258 480 8 la_data_out[13]
port 284 nsew default tristate
rlabel metal2 s 177734 -960 177846 480 8 la_data_out[14]
port 285 nsew default tristate
rlabel metal2 s 181322 -960 181434 480 8 la_data_out[15]
port 286 nsew default tristate
rlabel metal2 s 184818 -960 184930 480 8 la_data_out[16]
port 287 nsew default tristate
rlabel metal2 s 188406 -960 188518 480 8 la_data_out[17]
port 288 nsew default tristate
rlabel metal2 s 191994 -960 192106 480 8 la_data_out[18]
port 289 nsew default tristate
rlabel metal2 s 195582 -960 195694 480 8 la_data_out[19]
port 290 nsew default tristate
rlabel metal2 s 131366 -960 131478 480 8 la_data_out[1]
port 291 nsew default tristate
rlabel metal2 s 199170 -960 199282 480 8 la_data_out[20]
port 292 nsew default tristate
rlabel metal2 s 202666 -960 202778 480 8 la_data_out[21]
port 293 nsew default tristate
rlabel metal2 s 206254 -960 206366 480 8 la_data_out[22]
port 294 nsew default tristate
rlabel metal2 s 209842 -960 209954 480 8 la_data_out[23]
port 295 nsew default tristate
rlabel metal2 s 213430 -960 213542 480 8 la_data_out[24]
port 296 nsew default tristate
rlabel metal2 s 217018 -960 217130 480 8 la_data_out[25]
port 297 nsew default tristate
rlabel metal2 s 220514 -960 220626 480 8 la_data_out[26]
port 298 nsew default tristate
rlabel metal2 s 224102 -960 224214 480 8 la_data_out[27]
port 299 nsew default tristate
rlabel metal2 s 227690 -960 227802 480 8 la_data_out[28]
port 300 nsew default tristate
rlabel metal2 s 231278 -960 231390 480 8 la_data_out[29]
port 301 nsew default tristate
rlabel metal2 s 134862 -960 134974 480 8 la_data_out[2]
port 302 nsew default tristate
rlabel metal2 s 234774 -960 234886 480 8 la_data_out[30]
port 303 nsew default tristate
rlabel metal2 s 238362 -960 238474 480 8 la_data_out[31]
port 304 nsew default tristate
rlabel metal2 s 241950 -960 242062 480 8 la_data_out[32]
port 305 nsew default tristate
rlabel metal2 s 245538 -960 245650 480 8 la_data_out[33]
port 306 nsew default tristate
rlabel metal2 s 249126 -960 249238 480 8 la_data_out[34]
port 307 nsew default tristate
rlabel metal2 s 252622 -960 252734 480 8 la_data_out[35]
port 308 nsew default tristate
rlabel metal2 s 256210 -960 256322 480 8 la_data_out[36]
port 309 nsew default tristate
rlabel metal2 s 259798 -960 259910 480 8 la_data_out[37]
port 310 nsew default tristate
rlabel metal2 s 263386 -960 263498 480 8 la_data_out[38]
port 311 nsew default tristate
rlabel metal2 s 266974 -960 267086 480 8 la_data_out[39]
port 312 nsew default tristate
rlabel metal2 s 138450 -960 138562 480 8 la_data_out[3]
port 313 nsew default tristate
rlabel metal2 s 270470 -960 270582 480 8 la_data_out[40]
port 314 nsew default tristate
rlabel metal2 s 274058 -960 274170 480 8 la_data_out[41]
port 315 nsew default tristate
rlabel metal2 s 277646 -960 277758 480 8 la_data_out[42]
port 316 nsew default tristate
rlabel metal2 s 281234 -960 281346 480 8 la_data_out[43]
port 317 nsew default tristate
rlabel metal2 s 284730 -960 284842 480 8 la_data_out[44]
port 318 nsew default tristate
rlabel metal2 s 288318 -960 288430 480 8 la_data_out[45]
port 319 nsew default tristate
rlabel metal2 s 291906 -960 292018 480 8 la_data_out[46]
port 320 nsew default tristate
rlabel metal2 s 295494 -960 295606 480 8 la_data_out[47]
port 321 nsew default tristate
rlabel metal2 s 299082 -960 299194 480 8 la_data_out[48]
port 322 nsew default tristate
rlabel metal2 s 302578 -960 302690 480 8 la_data_out[49]
port 323 nsew default tristate
rlabel metal2 s 142038 -960 142150 480 8 la_data_out[4]
port 324 nsew default tristate
rlabel metal2 s 306166 -960 306278 480 8 la_data_out[50]
port 325 nsew default tristate
rlabel metal2 s 309754 -960 309866 480 8 la_data_out[51]
port 326 nsew default tristate
rlabel metal2 s 313342 -960 313454 480 8 la_data_out[52]
port 327 nsew default tristate
rlabel metal2 s 316930 -960 317042 480 8 la_data_out[53]
port 328 nsew default tristate
rlabel metal2 s 320426 -960 320538 480 8 la_data_out[54]
port 329 nsew default tristate
rlabel metal2 s 324014 -960 324126 480 8 la_data_out[55]
port 330 nsew default tristate
rlabel metal2 s 327602 -960 327714 480 8 la_data_out[56]
port 331 nsew default tristate
rlabel metal2 s 331190 -960 331302 480 8 la_data_out[57]
port 332 nsew default tristate
rlabel metal2 s 334686 -960 334798 480 8 la_data_out[58]
port 333 nsew default tristate
rlabel metal2 s 338274 -960 338386 480 8 la_data_out[59]
port 334 nsew default tristate
rlabel metal2 s 145626 -960 145738 480 8 la_data_out[5]
port 335 nsew default tristate
rlabel metal2 s 341862 -960 341974 480 8 la_data_out[60]
port 336 nsew default tristate
rlabel metal2 s 345450 -960 345562 480 8 la_data_out[61]
port 337 nsew default tristate
rlabel metal2 s 349038 -960 349150 480 8 la_data_out[62]
port 338 nsew default tristate
rlabel metal2 s 352534 -960 352646 480 8 la_data_out[63]
port 339 nsew default tristate
rlabel metal2 s 356122 -960 356234 480 8 la_data_out[64]
port 340 nsew default tristate
rlabel metal2 s 359710 -960 359822 480 8 la_data_out[65]
port 341 nsew default tristate
rlabel metal2 s 363298 -960 363410 480 8 la_data_out[66]
port 342 nsew default tristate
rlabel metal2 s 366886 -960 366998 480 8 la_data_out[67]
port 343 nsew default tristate
rlabel metal2 s 370382 -960 370494 480 8 la_data_out[68]
port 344 nsew default tristate
rlabel metal2 s 373970 -960 374082 480 8 la_data_out[69]
port 345 nsew default tristate
rlabel metal2 s 149214 -960 149326 480 8 la_data_out[6]
port 346 nsew default tristate
rlabel metal2 s 377558 -960 377670 480 8 la_data_out[70]
port 347 nsew default tristate
rlabel metal2 s 381146 -960 381258 480 8 la_data_out[71]
port 348 nsew default tristate
rlabel metal2 s 384642 -960 384754 480 8 la_data_out[72]
port 349 nsew default tristate
rlabel metal2 s 388230 -960 388342 480 8 la_data_out[73]
port 350 nsew default tristate
rlabel metal2 s 391818 -960 391930 480 8 la_data_out[74]
port 351 nsew default tristate
rlabel metal2 s 395406 -960 395518 480 8 la_data_out[75]
port 352 nsew default tristate
rlabel metal2 s 398994 -960 399106 480 8 la_data_out[76]
port 353 nsew default tristate
rlabel metal2 s 402490 -960 402602 480 8 la_data_out[77]
port 354 nsew default tristate
rlabel metal2 s 406078 -960 406190 480 8 la_data_out[78]
port 355 nsew default tristate
rlabel metal2 s 409666 -960 409778 480 8 la_data_out[79]
port 356 nsew default tristate
rlabel metal2 s 152710 -960 152822 480 8 la_data_out[7]
port 357 nsew default tristate
rlabel metal2 s 413254 -960 413366 480 8 la_data_out[80]
port 358 nsew default tristate
rlabel metal2 s 416842 -960 416954 480 8 la_data_out[81]
port 359 nsew default tristate
rlabel metal2 s 420338 -960 420450 480 8 la_data_out[82]
port 360 nsew default tristate
rlabel metal2 s 423926 -960 424038 480 8 la_data_out[83]
port 361 nsew default tristate
rlabel metal2 s 427514 -960 427626 480 8 la_data_out[84]
port 362 nsew default tristate
rlabel metal2 s 431102 -960 431214 480 8 la_data_out[85]
port 363 nsew default tristate
rlabel metal2 s 434598 -960 434710 480 8 la_data_out[86]
port 364 nsew default tristate
rlabel metal2 s 438186 -960 438298 480 8 la_data_out[87]
port 365 nsew default tristate
rlabel metal2 s 441774 -960 441886 480 8 la_data_out[88]
port 366 nsew default tristate
rlabel metal2 s 445362 -960 445474 480 8 la_data_out[89]
port 367 nsew default tristate
rlabel metal2 s 156298 -960 156410 480 8 la_data_out[8]
port 368 nsew default tristate
rlabel metal2 s 448950 -960 449062 480 8 la_data_out[90]
port 369 nsew default tristate
rlabel metal2 s 452446 -960 452558 480 8 la_data_out[91]
port 370 nsew default tristate
rlabel metal2 s 456034 -960 456146 480 8 la_data_out[92]
port 371 nsew default tristate
rlabel metal2 s 459622 -960 459734 480 8 la_data_out[93]
port 372 nsew default tristate
rlabel metal2 s 463210 -960 463322 480 8 la_data_out[94]
port 373 nsew default tristate
rlabel metal2 s 466798 -960 466910 480 8 la_data_out[95]
port 374 nsew default tristate
rlabel metal2 s 470294 -960 470406 480 8 la_data_out[96]
port 375 nsew default tristate
rlabel metal2 s 473882 -960 473994 480 8 la_data_out[97]
port 376 nsew default tristate
rlabel metal2 s 477470 -960 477582 480 8 la_data_out[98]
port 377 nsew default tristate
rlabel metal2 s 481058 -960 481170 480 8 la_data_out[99]
port 378 nsew default tristate
rlabel metal2 s 159886 -960 159998 480 8 la_data_out[9]
port 379 nsew default tristate
rlabel metal2 s 128974 -960 129086 480 8 la_oen[0]
port 380 nsew default input
rlabel metal2 s 485750 -960 485862 480 8 la_oen[100]
port 381 nsew default input
rlabel metal2 s 489338 -960 489450 480 8 la_oen[101]
port 382 nsew default input
rlabel metal2 s 492926 -960 493038 480 8 la_oen[102]
port 383 nsew default input
rlabel metal2 s 496514 -960 496626 480 8 la_oen[103]
port 384 nsew default input
rlabel metal2 s 500102 -960 500214 480 8 la_oen[104]
port 385 nsew default input
rlabel metal2 s 503598 -960 503710 480 8 la_oen[105]
port 386 nsew default input
rlabel metal2 s 507186 -960 507298 480 8 la_oen[106]
port 387 nsew default input
rlabel metal2 s 510774 -960 510886 480 8 la_oen[107]
port 388 nsew default input
rlabel metal2 s 514362 -960 514474 480 8 la_oen[108]
port 389 nsew default input
rlabel metal2 s 517858 -960 517970 480 8 la_oen[109]
port 390 nsew default input
rlabel metal2 s 164670 -960 164782 480 8 la_oen[10]
port 391 nsew default input
rlabel metal2 s 521446 -960 521558 480 8 la_oen[110]
port 392 nsew default input
rlabel metal2 s 525034 -960 525146 480 8 la_oen[111]
port 393 nsew default input
rlabel metal2 s 528622 -960 528734 480 8 la_oen[112]
port 394 nsew default input
rlabel metal2 s 532210 -960 532322 480 8 la_oen[113]
port 395 nsew default input
rlabel metal2 s 535706 -960 535818 480 8 la_oen[114]
port 396 nsew default input
rlabel metal2 s 539294 -960 539406 480 8 la_oen[115]
port 397 nsew default input
rlabel metal2 s 542882 -960 542994 480 8 la_oen[116]
port 398 nsew default input
rlabel metal2 s 546470 -960 546582 480 8 la_oen[117]
port 399 nsew default input
rlabel metal2 s 550058 -960 550170 480 8 la_oen[118]
port 400 nsew default input
rlabel metal2 s 553554 -960 553666 480 8 la_oen[119]
port 401 nsew default input
rlabel metal2 s 168166 -960 168278 480 8 la_oen[11]
port 402 nsew default input
rlabel metal2 s 557142 -960 557254 480 8 la_oen[120]
port 403 nsew default input
rlabel metal2 s 560730 -960 560842 480 8 la_oen[121]
port 404 nsew default input
rlabel metal2 s 564318 -960 564430 480 8 la_oen[122]
port 405 nsew default input
rlabel metal2 s 567814 -960 567926 480 8 la_oen[123]
port 406 nsew default input
rlabel metal2 s 571402 -960 571514 480 8 la_oen[124]
port 407 nsew default input
rlabel metal2 s 574990 -960 575102 480 8 la_oen[125]
port 408 nsew default input
rlabel metal2 s 578578 -960 578690 480 8 la_oen[126]
port 409 nsew default input
rlabel metal2 s 582166 -960 582278 480 8 la_oen[127]
port 410 nsew default input
rlabel metal2 s 171754 -960 171866 480 8 la_oen[12]
port 411 nsew default input
rlabel metal2 s 175342 -960 175454 480 8 la_oen[13]
port 412 nsew default input
rlabel metal2 s 178930 -960 179042 480 8 la_oen[14]
port 413 nsew default input
rlabel metal2 s 182518 -960 182630 480 8 la_oen[15]
port 414 nsew default input
rlabel metal2 s 186014 -960 186126 480 8 la_oen[16]
port 415 nsew default input
rlabel metal2 s 189602 -960 189714 480 8 la_oen[17]
port 416 nsew default input
rlabel metal2 s 193190 -960 193302 480 8 la_oen[18]
port 417 nsew default input
rlabel metal2 s 196778 -960 196890 480 8 la_oen[19]
port 418 nsew default input
rlabel metal2 s 132562 -960 132674 480 8 la_oen[1]
port 419 nsew default input
rlabel metal2 s 200366 -960 200478 480 8 la_oen[20]
port 420 nsew default input
rlabel metal2 s 203862 -960 203974 480 8 la_oen[21]
port 421 nsew default input
rlabel metal2 s 207450 -960 207562 480 8 la_oen[22]
port 422 nsew default input
rlabel metal2 s 211038 -960 211150 480 8 la_oen[23]
port 423 nsew default input
rlabel metal2 s 214626 -960 214738 480 8 la_oen[24]
port 424 nsew default input
rlabel metal2 s 218122 -960 218234 480 8 la_oen[25]
port 425 nsew default input
rlabel metal2 s 221710 -960 221822 480 8 la_oen[26]
port 426 nsew default input
rlabel metal2 s 225298 -960 225410 480 8 la_oen[27]
port 427 nsew default input
rlabel metal2 s 228886 -960 228998 480 8 la_oen[28]
port 428 nsew default input
rlabel metal2 s 232474 -960 232586 480 8 la_oen[29]
port 429 nsew default input
rlabel metal2 s 136058 -960 136170 480 8 la_oen[2]
port 430 nsew default input
rlabel metal2 s 235970 -960 236082 480 8 la_oen[30]
port 431 nsew default input
rlabel metal2 s 239558 -960 239670 480 8 la_oen[31]
port 432 nsew default input
rlabel metal2 s 243146 -960 243258 480 8 la_oen[32]
port 433 nsew default input
rlabel metal2 s 246734 -960 246846 480 8 la_oen[33]
port 434 nsew default input
rlabel metal2 s 250322 -960 250434 480 8 la_oen[34]
port 435 nsew default input
rlabel metal2 s 253818 -960 253930 480 8 la_oen[35]
port 436 nsew default input
rlabel metal2 s 257406 -960 257518 480 8 la_oen[36]
port 437 nsew default input
rlabel metal2 s 260994 -960 261106 480 8 la_oen[37]
port 438 nsew default input
rlabel metal2 s 264582 -960 264694 480 8 la_oen[38]
port 439 nsew default input
rlabel metal2 s 268078 -960 268190 480 8 la_oen[39]
port 440 nsew default input
rlabel metal2 s 139646 -960 139758 480 8 la_oen[3]
port 441 nsew default input
rlabel metal2 s 271666 -960 271778 480 8 la_oen[40]
port 442 nsew default input
rlabel metal2 s 275254 -960 275366 480 8 la_oen[41]
port 443 nsew default input
rlabel metal2 s 278842 -960 278954 480 8 la_oen[42]
port 444 nsew default input
rlabel metal2 s 282430 -960 282542 480 8 la_oen[43]
port 445 nsew default input
rlabel metal2 s 285926 -960 286038 480 8 la_oen[44]
port 446 nsew default input
rlabel metal2 s 289514 -960 289626 480 8 la_oen[45]
port 447 nsew default input
rlabel metal2 s 293102 -960 293214 480 8 la_oen[46]
port 448 nsew default input
rlabel metal2 s 296690 -960 296802 480 8 la_oen[47]
port 449 nsew default input
rlabel metal2 s 300278 -960 300390 480 8 la_oen[48]
port 450 nsew default input
rlabel metal2 s 303774 -960 303886 480 8 la_oen[49]
port 451 nsew default input
rlabel metal2 s 143234 -960 143346 480 8 la_oen[4]
port 452 nsew default input
rlabel metal2 s 307362 -960 307474 480 8 la_oen[50]
port 453 nsew default input
rlabel metal2 s 310950 -960 311062 480 8 la_oen[51]
port 454 nsew default input
rlabel metal2 s 314538 -960 314650 480 8 la_oen[52]
port 455 nsew default input
rlabel metal2 s 318034 -960 318146 480 8 la_oen[53]
port 456 nsew default input
rlabel metal2 s 321622 -960 321734 480 8 la_oen[54]
port 457 nsew default input
rlabel metal2 s 325210 -960 325322 480 8 la_oen[55]
port 458 nsew default input
rlabel metal2 s 328798 -960 328910 480 8 la_oen[56]
port 459 nsew default input
rlabel metal2 s 332386 -960 332498 480 8 la_oen[57]
port 460 nsew default input
rlabel metal2 s 335882 -960 335994 480 8 la_oen[58]
port 461 nsew default input
rlabel metal2 s 339470 -960 339582 480 8 la_oen[59]
port 462 nsew default input
rlabel metal2 s 146822 -960 146934 480 8 la_oen[5]
port 463 nsew default input
rlabel metal2 s 343058 -960 343170 480 8 la_oen[60]
port 464 nsew default input
rlabel metal2 s 346646 -960 346758 480 8 la_oen[61]
port 465 nsew default input
rlabel metal2 s 350234 -960 350346 480 8 la_oen[62]
port 466 nsew default input
rlabel metal2 s 353730 -960 353842 480 8 la_oen[63]
port 467 nsew default input
rlabel metal2 s 357318 -960 357430 480 8 la_oen[64]
port 468 nsew default input
rlabel metal2 s 360906 -960 361018 480 8 la_oen[65]
port 469 nsew default input
rlabel metal2 s 364494 -960 364606 480 8 la_oen[66]
port 470 nsew default input
rlabel metal2 s 367990 -960 368102 480 8 la_oen[67]
port 471 nsew default input
rlabel metal2 s 371578 -960 371690 480 8 la_oen[68]
port 472 nsew default input
rlabel metal2 s 375166 -960 375278 480 8 la_oen[69]
port 473 nsew default input
rlabel metal2 s 150410 -960 150522 480 8 la_oen[6]
port 474 nsew default input
rlabel metal2 s 378754 -960 378866 480 8 la_oen[70]
port 475 nsew default input
rlabel metal2 s 382342 -960 382454 480 8 la_oen[71]
port 476 nsew default input
rlabel metal2 s 385838 -960 385950 480 8 la_oen[72]
port 477 nsew default input
rlabel metal2 s 389426 -960 389538 480 8 la_oen[73]
port 478 nsew default input
rlabel metal2 s 393014 -960 393126 480 8 la_oen[74]
port 479 nsew default input
rlabel metal2 s 396602 -960 396714 480 8 la_oen[75]
port 480 nsew default input
rlabel metal2 s 400190 -960 400302 480 8 la_oen[76]
port 481 nsew default input
rlabel metal2 s 403686 -960 403798 480 8 la_oen[77]
port 482 nsew default input
rlabel metal2 s 407274 -960 407386 480 8 la_oen[78]
port 483 nsew default input
rlabel metal2 s 410862 -960 410974 480 8 la_oen[79]
port 484 nsew default input
rlabel metal2 s 153906 -960 154018 480 8 la_oen[7]
port 485 nsew default input
rlabel metal2 s 414450 -960 414562 480 8 la_oen[80]
port 486 nsew default input
rlabel metal2 s 417946 -960 418058 480 8 la_oen[81]
port 487 nsew default input
rlabel metal2 s 421534 -960 421646 480 8 la_oen[82]
port 488 nsew default input
rlabel metal2 s 425122 -960 425234 480 8 la_oen[83]
port 489 nsew default input
rlabel metal2 s 428710 -960 428822 480 8 la_oen[84]
port 490 nsew default input
rlabel metal2 s 432298 -960 432410 480 8 la_oen[85]
port 491 nsew default input
rlabel metal2 s 435794 -960 435906 480 8 la_oen[86]
port 492 nsew default input
rlabel metal2 s 439382 -960 439494 480 8 la_oen[87]
port 493 nsew default input
rlabel metal2 s 442970 -960 443082 480 8 la_oen[88]
port 494 nsew default input
rlabel metal2 s 446558 -960 446670 480 8 la_oen[89]
port 495 nsew default input
rlabel metal2 s 157494 -960 157606 480 8 la_oen[8]
port 496 nsew default input
rlabel metal2 s 450146 -960 450258 480 8 la_oen[90]
port 497 nsew default input
rlabel metal2 s 453642 -960 453754 480 8 la_oen[91]
port 498 nsew default input
rlabel metal2 s 457230 -960 457342 480 8 la_oen[92]
port 499 nsew default input
rlabel metal2 s 460818 -960 460930 480 8 la_oen[93]
port 500 nsew default input
rlabel metal2 s 464406 -960 464518 480 8 la_oen[94]
port 501 nsew default input
rlabel metal2 s 467902 -960 468014 480 8 la_oen[95]
port 502 nsew default input
rlabel metal2 s 471490 -960 471602 480 8 la_oen[96]
port 503 nsew default input
rlabel metal2 s 475078 -960 475190 480 8 la_oen[97]
port 504 nsew default input
rlabel metal2 s 478666 -960 478778 480 8 la_oen[98]
port 505 nsew default input
rlabel metal2 s 482254 -960 482366 480 8 la_oen[99]
port 506 nsew default input
rlabel metal2 s 161082 -960 161194 480 8 la_oen[9]
port 507 nsew default input
rlabel metal3 s 583520 510220 584960 510460 6 io_oeb[10]
port 508 nsew default tristate
rlabel metal3 s 583520 557140 584960 557380 6 io_oeb[11]
port 509 nsew default tristate
rlabel metal3 s 583520 604060 584960 604300 6 io_oeb[12]
port 510 nsew default tristate
rlabel metal3 s 583520 650980 584960 651220 6 io_oeb[13]
port 511 nsew default tristate
rlabel metal3 s 583520 697900 584960 698140 6 io_oeb[14]
port 512 nsew default tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 513 nsew default tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 514 nsew default tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 515 nsew default tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 516 nsew default tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 517 nsew default tristate
rlabel metal3 s 583520 416380 584960 416620 6 io_oeb[8]
port 518 nsew default tristate
rlabel metal3 s 583520 463300 584960 463540 6 io_oeb[9]
port 519 nsew default tristate
rlabel metal2 s 583362 -960 583474 480 8 user_clock2
port 520 nsew default input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 521 nsew default input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 522 nsew default input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 523 nsew default tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 524 nsew default input
rlabel metal2 s 48106 -960 48218 480 8 wbs_adr_i[10]
port 525 nsew default input
rlabel metal2 s 51602 -960 51714 480 8 wbs_adr_i[11]
port 526 nsew default input
rlabel metal2 s 55190 -960 55302 480 8 wbs_adr_i[12]
port 527 nsew default input
rlabel metal2 s 58778 -960 58890 480 8 wbs_adr_i[13]
port 528 nsew default input
rlabel metal2 s 62366 -960 62478 480 8 wbs_adr_i[14]
port 529 nsew default input
rlabel metal2 s 65954 -960 66066 480 8 wbs_adr_i[15]
port 530 nsew default input
rlabel metal2 s 69450 -960 69562 480 8 wbs_adr_i[16]
port 531 nsew default input
rlabel metal2 s 73038 -960 73150 480 8 wbs_adr_i[17]
port 532 nsew default input
rlabel metal2 s 76626 -960 76738 480 8 wbs_adr_i[18]
port 533 nsew default input
rlabel metal2 s 80214 -960 80326 480 8 wbs_adr_i[19]
port 534 nsew default input
rlabel metal2 s 12410 -960 12522 480 8 wbs_adr_i[1]
port 535 nsew default input
rlabel metal2 s 83802 -960 83914 480 8 wbs_adr_i[20]
port 536 nsew default input
rlabel metal2 s 87298 -960 87410 480 8 wbs_adr_i[21]
port 537 nsew default input
rlabel metal2 s 90886 -960 90998 480 8 wbs_adr_i[22]
port 538 nsew default input
rlabel metal2 s 94474 -960 94586 480 8 wbs_adr_i[23]
port 539 nsew default input
rlabel metal2 s 98062 -960 98174 480 8 wbs_adr_i[24]
port 540 nsew default input
rlabel metal2 s 101558 -960 101670 480 8 wbs_adr_i[25]
port 541 nsew default input
rlabel metal2 s 105146 -960 105258 480 8 wbs_adr_i[26]
port 542 nsew default input
rlabel metal2 s 108734 -960 108846 480 8 wbs_adr_i[27]
port 543 nsew default input
rlabel metal2 s 112322 -960 112434 480 8 wbs_adr_i[28]
port 544 nsew default input
rlabel metal2 s 115910 -960 116022 480 8 wbs_adr_i[29]
port 545 nsew default input
rlabel metal2 s 17194 -960 17306 480 8 wbs_adr_i[2]
port 546 nsew default input
rlabel metal2 s 119406 -960 119518 480 8 wbs_adr_i[30]
port 547 nsew default input
rlabel metal2 s 122994 -960 123106 480 8 wbs_adr_i[31]
port 548 nsew default input
rlabel metal2 s 21886 -960 21998 480 8 wbs_adr_i[3]
port 549 nsew default input
rlabel metal2 s 26670 -960 26782 480 8 wbs_adr_i[4]
port 550 nsew default input
rlabel metal2 s 30258 -960 30370 480 8 wbs_adr_i[5]
port 551 nsew default input
rlabel metal2 s 33846 -960 33958 480 8 wbs_adr_i[6]
port 552 nsew default input
rlabel metal2 s 37342 -960 37454 480 8 wbs_adr_i[7]
port 553 nsew default input
rlabel metal2 s 40930 -960 41042 480 8 wbs_adr_i[8]
port 554 nsew default input
rlabel metal2 s 44518 -960 44630 480 8 wbs_adr_i[9]
port 555 nsew default input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 556 nsew default input
rlabel metal2 s 8822 -960 8934 480 8 wbs_dat_i[0]
port 557 nsew default input
rlabel metal2 s 49302 -960 49414 480 8 wbs_dat_i[10]
port 558 nsew default input
rlabel metal2 s 52798 -960 52910 480 8 wbs_dat_i[11]
port 559 nsew default input
rlabel metal2 s 56386 -960 56498 480 8 wbs_dat_i[12]
port 560 nsew default input
rlabel metal2 s 59974 -960 60086 480 8 wbs_dat_i[13]
port 561 nsew default input
rlabel metal2 s 63562 -960 63674 480 8 wbs_dat_i[14]
port 562 nsew default input
rlabel metal2 s 67150 -960 67262 480 8 wbs_dat_i[15]
port 563 nsew default input
rlabel metal2 s 70646 -960 70758 480 8 wbs_dat_i[16]
port 564 nsew default input
rlabel metal2 s 74234 -960 74346 480 8 wbs_dat_i[17]
port 565 nsew default input
rlabel metal2 s 77822 -960 77934 480 8 wbs_dat_i[18]
port 566 nsew default input
rlabel metal2 s 81410 -960 81522 480 8 wbs_dat_i[19]
port 567 nsew default input
rlabel metal2 s 13606 -960 13718 480 8 wbs_dat_i[1]
port 568 nsew default input
rlabel metal2 s 84906 -960 85018 480 8 wbs_dat_i[20]
port 569 nsew default input
rlabel metal2 s 88494 -960 88606 480 8 wbs_dat_i[21]
port 570 nsew default input
rlabel metal2 s 92082 -960 92194 480 8 wbs_dat_i[22]
port 571 nsew default input
rlabel metal2 s 95670 -960 95782 480 8 wbs_dat_i[23]
port 572 nsew default input
rlabel metal2 s 99258 -960 99370 480 8 wbs_dat_i[24]
port 573 nsew default input
rlabel metal2 s 102754 -960 102866 480 8 wbs_dat_i[25]
port 574 nsew default input
rlabel metal2 s 106342 -960 106454 480 8 wbs_dat_i[26]
port 575 nsew default input
rlabel metal2 s 109930 -960 110042 480 8 wbs_dat_i[27]
port 576 nsew default input
rlabel metal2 s 113518 -960 113630 480 8 wbs_dat_i[28]
port 577 nsew default input
rlabel metal2 s 117106 -960 117218 480 8 wbs_dat_i[29]
port 578 nsew default input
rlabel metal2 s 18298 -960 18410 480 8 wbs_dat_i[2]
port 579 nsew default input
rlabel metal2 s 120602 -960 120714 480 8 wbs_dat_i[30]
port 580 nsew default input
rlabel metal2 s 124190 -960 124302 480 8 wbs_dat_i[31]
port 581 nsew default input
rlabel metal2 s 23082 -960 23194 480 8 wbs_dat_i[3]
port 582 nsew default input
rlabel metal2 s 27866 -960 27978 480 8 wbs_dat_i[4]
port 583 nsew default input
rlabel metal2 s 31454 -960 31566 480 8 wbs_dat_i[5]
port 584 nsew default input
rlabel metal2 s 34950 -960 35062 480 8 wbs_dat_i[6]
port 585 nsew default input
rlabel metal2 s 38538 -960 38650 480 8 wbs_dat_i[7]
port 586 nsew default input
rlabel metal2 s 42126 -960 42238 480 8 wbs_dat_i[8]
port 587 nsew default input
rlabel metal2 s 45714 -960 45826 480 8 wbs_dat_i[9]
port 588 nsew default input
rlabel metal2 s 10018 -960 10130 480 8 wbs_dat_o[0]
port 589 nsew default tristate
rlabel metal2 s 50498 -960 50610 480 8 wbs_dat_o[10]
port 590 nsew default tristate
rlabel metal2 s 53994 -960 54106 480 8 wbs_dat_o[11]
port 591 nsew default tristate
rlabel metal2 s 57582 -960 57694 480 8 wbs_dat_o[12]
port 592 nsew default tristate
rlabel metal2 s 61170 -960 61282 480 8 wbs_dat_o[13]
port 593 nsew default tristate
rlabel metal2 s 64758 -960 64870 480 8 wbs_dat_o[14]
port 594 nsew default tristate
rlabel metal2 s 68254 -960 68366 480 8 wbs_dat_o[15]
port 595 nsew default tristate
rlabel metal2 s 71842 -960 71954 480 8 wbs_dat_o[16]
port 596 nsew default tristate
rlabel metal2 s 75430 -960 75542 480 8 wbs_dat_o[17]
port 597 nsew default tristate
rlabel metal2 s 79018 -960 79130 480 8 wbs_dat_o[18]
port 598 nsew default tristate
rlabel metal2 s 82606 -960 82718 480 8 wbs_dat_o[19]
port 599 nsew default tristate
rlabel metal2 s 14802 -960 14914 480 8 wbs_dat_o[1]
port 600 nsew default tristate
rlabel metal2 s 86102 -960 86214 480 8 wbs_dat_o[20]
port 601 nsew default tristate
rlabel metal2 s 89690 -960 89802 480 8 wbs_dat_o[21]
port 602 nsew default tristate
rlabel metal2 s 93278 -960 93390 480 8 wbs_dat_o[22]
port 603 nsew default tristate
rlabel metal2 s 96866 -960 96978 480 8 wbs_dat_o[23]
port 604 nsew default tristate
rlabel metal2 s 100454 -960 100566 480 8 wbs_dat_o[24]
port 605 nsew default tristate
rlabel metal2 s 103950 -960 104062 480 8 wbs_dat_o[25]
port 606 nsew default tristate
rlabel metal2 s 107538 -960 107650 480 8 wbs_dat_o[26]
port 607 nsew default tristate
rlabel metal2 s 111126 -960 111238 480 8 wbs_dat_o[27]
port 608 nsew default tristate
rlabel metal2 s 114714 -960 114826 480 8 wbs_dat_o[28]
port 609 nsew default tristate
rlabel metal2 s 118210 -960 118322 480 8 wbs_dat_o[29]
port 610 nsew default tristate
rlabel metal2 s 19494 -960 19606 480 8 wbs_dat_o[2]
port 611 nsew default tristate
rlabel metal2 s 121798 -960 121910 480 8 wbs_dat_o[30]
port 612 nsew default tristate
rlabel metal2 s 125386 -960 125498 480 8 wbs_dat_o[31]
port 613 nsew default tristate
rlabel metal2 s 24278 -960 24390 480 8 wbs_dat_o[3]
port 614 nsew default tristate
rlabel metal2 s 29062 -960 29174 480 8 wbs_dat_o[4]
port 615 nsew default tristate
rlabel metal2 s 32650 -960 32762 480 8 wbs_dat_o[5]
port 616 nsew default tristate
rlabel metal2 s 36146 -960 36258 480 8 wbs_dat_o[6]
port 617 nsew default tristate
rlabel metal2 s 39734 -960 39846 480 8 wbs_dat_o[7]
port 618 nsew default tristate
rlabel metal2 s 43322 -960 43434 480 8 wbs_dat_o[8]
port 619 nsew default tristate
rlabel metal2 s 46910 -960 47022 480 8 wbs_dat_o[9]
port 620 nsew default tristate
rlabel metal2 s 11214 -960 11326 480 8 wbs_sel_i[0]
port 621 nsew default input
rlabel metal2 s 15998 -960 16110 480 8 wbs_sel_i[1]
port 622 nsew default input
rlabel metal2 s 20690 -960 20802 480 8 wbs_sel_i[2]
port 623 nsew default input
rlabel metal2 s 25474 -960 25586 480 8 wbs_sel_i[3]
port 624 nsew default input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 625 nsew default input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 626 nsew default input
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 627 nsew default tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 628 nsew default tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 629 nsew default tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 630 nsew default tristate
rlabel metal3 s -960 653428 480 653668 4 io_oeb[24]
port 631 nsew default tristate
rlabel metal3 s -960 595900 480 596140 4 io_oeb[25]
port 632 nsew default tristate
rlabel metal3 s -960 538508 480 538748 4 io_oeb[26]
port 633 nsew default tristate
rlabel metal3 s -960 480980 480 481220 4 io_oeb[27]
port 634 nsew default tristate
rlabel metal3 s -960 423588 480 423828 4 io_oeb[28]
port 635 nsew default tristate
rlabel metal5 s -1996 -924 585920 -324 8 vccd1
port 636 nsew default input
rlabel metal5 s -2936 -1864 586860 -1264 8 vssd1
port 637 nsew default input
rlabel metal5 s -3876 -2804 587800 -2204 8 vccd2
port 638 nsew default input
rlabel metal5 s -4816 -3744 588740 -3144 8 vssd2
port 639 nsew default input
rlabel metal5 s -5756 -4684 589680 -4084 8 vdda1
port 640 nsew default input
rlabel metal5 s -6696 -5624 590620 -5024 8 vssa1
port 641 nsew default input
rlabel metal5 s -7636 -6564 591560 -5964 8 vdda2
port 642 nsew default input
rlabel metal5 s -8576 -7504 592500 -6904 8 vssa2
port 643 nsew default input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>

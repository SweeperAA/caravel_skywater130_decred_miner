magic
tech sky130A
magscale 1 2
timestamp 1611787880
<< obsli1 >>
rect 1104 2159 242880 201841
<< obsm1 >>
rect 382 1776 242880 201872
<< metal2 >>
rect 10506 203200 10562 204000
rect 35162 203200 35218 204000
rect 59634 203200 59690 204000
rect 84106 203200 84162 204000
rect 108578 203200 108634 204000
rect 133050 203200 133106 204000
rect 157522 203200 157578 204000
rect 182178 203200 182234 204000
rect 206650 203200 206706 204000
rect 231122 203200 231178 204000
rect 570 0 626 800
rect 25042 0 25098 800
rect 49514 0 49570 800
rect 73986 0 74042 800
rect 98458 0 98514 800
rect 122930 0 122986 800
rect 147402 0 147458 800
rect 172058 0 172114 800
rect 196530 0 196586 800
rect 221002 0 221058 800
<< obsm2 >>
rect 386 203144 10450 203200
rect 10618 203144 35106 203200
rect 35274 203144 59578 203200
rect 59746 203144 84050 203200
rect 84218 203144 108522 203200
rect 108690 203144 132994 203200
rect 133162 203144 157466 203200
rect 157634 203144 182122 203200
rect 182290 203144 206594 203200
rect 206762 203144 231066 203200
rect 231234 203144 242126 203200
rect 386 856 242126 203144
rect 386 800 514 856
rect 682 800 24986 856
rect 25154 800 49458 856
rect 49626 800 73930 856
rect 74098 800 98402 856
rect 98570 800 122874 856
rect 123042 800 147346 856
rect 147514 800 172002 856
rect 172170 800 196474 856
rect 196642 800 220946 856
rect 221114 800 242126 856
<< metal3 >>
rect 243200 184968 244000 185088
rect 0 181704 800 181824
rect 243200 148792 244000 148912
rect 0 145528 800 145648
rect 243200 112616 244000 112736
rect 0 109352 800 109472
rect 243200 76168 244000 76288
rect 0 73176 800 73296
rect 243200 39992 244000 40112
rect 0 37000 800 37120
rect 243200 3816 244000 3936
<< obsm3 >>
rect 381 185168 243200 201857
rect 381 184888 243120 185168
rect 381 181904 243200 184888
rect 880 181624 243200 181904
rect 381 148992 243200 181624
rect 381 148712 243120 148992
rect 381 145728 243200 148712
rect 880 145448 243200 145728
rect 381 112816 243200 145448
rect 381 112536 243120 112816
rect 381 109552 243200 112536
rect 880 109272 243200 109552
rect 381 76368 243200 109272
rect 381 76088 243120 76368
rect 381 73376 243200 76088
rect 880 73096 243200 73376
rect 381 40192 243200 73096
rect 381 39912 243120 40192
rect 381 37200 243200 39912
rect 880 36920 243200 37200
rect 381 4016 243200 36920
rect 381 3736 243120 4016
rect 381 2143 243200 3736
<< metal4 >>
rect 4208 2128 4528 201872
rect 4868 2176 5188 201824
rect 5528 2176 5848 201824
rect 6188 2176 6508 201824
rect 19568 2128 19888 201872
rect 20228 2176 20548 201824
rect 20888 2176 21208 201824
rect 21548 2176 21868 201824
rect 34928 2128 35248 201872
rect 35588 2176 35908 201824
rect 36248 2176 36568 201824
rect 36908 2176 37228 201824
rect 50288 2128 50608 201872
rect 50948 2176 51268 201824
rect 51608 2176 51928 201824
rect 52268 2176 52588 201824
rect 65648 2128 65968 201872
rect 66308 2176 66628 201824
rect 66968 2176 67288 201824
rect 67628 2176 67948 201824
rect 81008 2128 81328 201872
rect 81668 2176 81988 201824
rect 82328 2176 82648 201824
rect 82988 2176 83308 201824
rect 96368 2128 96688 201872
rect 97028 2176 97348 201824
rect 97688 2176 98008 201824
rect 98348 2176 98668 201824
rect 111728 2128 112048 201872
rect 112388 2176 112708 201824
rect 113048 2176 113368 201824
rect 113708 2176 114028 201824
rect 127088 2128 127408 201872
rect 127748 2176 128068 201824
rect 128408 2176 128728 201824
rect 129068 2176 129388 201824
rect 142448 2128 142768 201872
rect 143108 2176 143428 201824
rect 143768 2176 144088 201824
rect 144428 2176 144748 201824
rect 157808 2128 158128 201872
rect 158468 2176 158788 201824
rect 159128 2176 159448 201824
rect 159788 2176 160108 201824
rect 173168 2128 173488 201872
rect 173828 2176 174148 201824
rect 174488 2176 174808 201824
rect 175148 2176 175468 201824
rect 188528 2128 188848 201872
rect 189188 2176 189508 201824
rect 189848 2176 190168 201824
rect 190508 2176 190828 201824
rect 203888 2128 204208 201872
rect 204548 2176 204868 201824
rect 205208 2176 205528 201824
rect 205868 2176 206188 201824
rect 219248 2128 219568 201872
rect 219908 2176 220228 201824
rect 220568 2176 220888 201824
rect 221228 2176 221548 201824
rect 234608 2128 234928 201872
rect 235268 2176 235588 201824
rect 235928 2176 236248 201824
rect 236588 2176 236908 201824
<< obsm4 >>
rect 611 3299 4128 200973
rect 4608 3299 4788 200973
rect 5268 3299 5448 200973
rect 5928 3299 6108 200973
rect 6588 3299 19488 200973
rect 19968 3299 20148 200973
rect 20628 3299 20808 200973
rect 21288 3299 21468 200973
rect 21948 3299 34848 200973
rect 35328 3299 35508 200973
rect 35988 3299 36168 200973
rect 36648 3299 36828 200973
rect 37308 3299 50208 200973
rect 50688 3299 50868 200973
rect 51348 3299 51528 200973
rect 52008 3299 52188 200973
rect 52668 3299 65568 200973
rect 66048 3299 66228 200973
rect 66708 3299 66888 200973
rect 67368 3299 67548 200973
rect 68028 3299 80928 200973
rect 81408 3299 81588 200973
rect 82068 3299 82248 200973
rect 82728 3299 82908 200973
rect 83388 3299 96288 200973
rect 96768 3299 96948 200973
rect 97428 3299 97608 200973
rect 98088 3299 98268 200973
rect 98748 3299 111648 200973
rect 112128 3299 112308 200973
rect 112788 3299 112968 200973
rect 113448 3299 113628 200973
rect 114108 3299 127008 200973
rect 127488 3299 127668 200973
rect 128148 3299 128328 200973
rect 128808 3299 128988 200973
rect 129468 3299 142368 200973
rect 142848 3299 143028 200973
rect 143508 3299 143688 200973
rect 144168 3299 144348 200973
rect 144828 3299 157728 200973
rect 158208 3299 158388 200973
rect 158868 3299 159048 200973
rect 159528 3299 159708 200973
rect 160188 3299 173088 200973
rect 173568 3299 173748 200973
rect 174228 3299 174408 200973
rect 174888 3299 175068 200973
rect 175548 3299 188448 200973
rect 188928 3299 189108 200973
rect 189588 3299 189768 200973
rect 190248 3299 190428 200973
rect 190908 3299 203808 200973
rect 204288 3299 204468 200973
rect 204948 3299 205128 200973
rect 205608 3299 205788 200973
rect 206268 3299 219168 200973
rect 219648 3299 219828 200973
rect 220308 3299 220488 200973
rect 220968 3299 221148 200973
rect 221628 3299 234528 200973
rect 235008 3299 235188 200973
rect 235668 3299 235848 200973
rect 236328 3299 236508 200973
rect 236988 3299 239325 200973
<< obsm5 >>
rect 153020 146380 161620 148060
<< labels >>
rlabel metal2 s 133050 203200 133106 204000 6 CLK
port 1 nsew signal input
rlabel metal2 s 147402 0 147458 800 6 DATA_AVAILABLE
port 2 nsew signal output
rlabel metal2 s 25042 0 25098 800 6 DATA_FROM_HASH[0]
port 3 nsew signal output
rlabel metal2 s 570 0 626 800 6 DATA_FROM_HASH[1]
port 4 nsew signal output
rlabel metal2 s 182178 203200 182234 204000 6 DATA_FROM_HASH[2]
port 5 nsew signal output
rlabel metal2 s 221002 0 221058 800 6 DATA_FROM_HASH[3]
port 6 nsew signal output
rlabel metal3 s 243200 39992 244000 40112 6 DATA_FROM_HASH[4]
port 7 nsew signal output
rlabel metal2 s 73986 0 74042 800 6 DATA_FROM_HASH[5]
port 8 nsew signal output
rlabel metal2 s 35162 203200 35218 204000 6 DATA_FROM_HASH[6]
port 9 nsew signal output
rlabel metal3 s 0 145528 800 145648 6 DATA_FROM_HASH[7]
port 10 nsew signal output
rlabel metal2 s 84106 203200 84162 204000 6 DATA_TO_HASH[0]
port 11 nsew signal input
rlabel metal3 s 0 73176 800 73296 6 DATA_TO_HASH[1]
port 12 nsew signal input
rlabel metal3 s 243200 76168 244000 76288 6 DATA_TO_HASH[2]
port 13 nsew signal input
rlabel metal3 s 243200 3816 244000 3936 6 DATA_TO_HASH[3]
port 14 nsew signal input
rlabel metal3 s 0 181704 800 181824 6 DATA_TO_HASH[4]
port 15 nsew signal input
rlabel metal2 s 49514 0 49570 800 6 DATA_TO_HASH[5]
port 16 nsew signal input
rlabel metal2 s 206650 203200 206706 204000 6 DATA_TO_HASH[6]
port 17 nsew signal input
rlabel metal2 s 59634 203200 59690 204000 6 DATA_TO_HASH[7]
port 18 nsew signal input
rlabel metal2 s 157522 203200 157578 204000 6 HASH_ADDR[0]
port 19 nsew signal input
rlabel metal2 s 10506 203200 10562 204000 6 HASH_ADDR[1]
port 20 nsew signal input
rlabel metal2 s 231122 203200 231178 204000 6 HASH_ADDR[2]
port 21 nsew signal input
rlabel metal2 s 196530 0 196586 800 6 HASH_ADDR[3]
port 22 nsew signal input
rlabel metal3 s 0 37000 800 37120 6 HASH_ADDR[4]
port 23 nsew signal input
rlabel metal3 s 243200 184968 244000 185088 6 HASH_ADDR[5]
port 24 nsew signal input
rlabel metal2 s 98458 0 98514 800 6 HASH_EN
port 25 nsew signal input
rlabel metal2 s 122930 0 122986 800 6 MACRO_RD_SELECT
port 26 nsew signal input
rlabel metal3 s 243200 112616 244000 112736 6 MACRO_WR_SELECT
port 27 nsew signal input
rlabel metal3 s 243200 148792 244000 148912 6 THREAD_COUNT[0]
port 28 nsew signal output
rlabel metal3 s 0 109352 800 109472 6 THREAD_COUNT[1]
port 29 nsew signal output
rlabel metal2 s 108578 203200 108634 204000 6 THREAD_COUNT[2]
port 30 nsew signal output
rlabel metal2 s 172058 0 172114 800 6 THREAD_COUNT[3]
port 31 nsew signal output
rlabel metal4 s 219248 2128 219568 201872 6 vccd1
port 32 nsew power bidirectional
rlabel metal4 s 188528 2128 188848 201872 6 vccd1
port 33 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 201872 6 vccd1
port 34 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 201872 6 vccd1
port 35 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 201872 6 vccd1
port 36 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 201872 6 vccd1
port 37 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 201872 6 vccd1
port 38 nsew power bidirectional
rlabel metal4 s 4208 2128 4528 201872 6 vccd1
port 39 nsew power bidirectional
rlabel metal4 s 234608 2128 234928 201872 6 vssd1
port 40 nsew ground bidirectional
rlabel metal4 s 203888 2128 204208 201872 6 vssd1
port 41 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 201872 6 vssd1
port 42 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 201872 6 vssd1
port 43 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 201872 6 vssd1
port 44 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 201872 6 vssd1
port 45 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 201872 6 vssd1
port 46 nsew ground bidirectional
rlabel metal4 s 19568 2128 19888 201872 6 vssd1
port 47 nsew ground bidirectional
rlabel metal4 s 219908 2176 220228 201824 6 vccd2
port 48 nsew power bidirectional
rlabel metal4 s 189188 2176 189508 201824 6 vccd2
port 49 nsew power bidirectional
rlabel metal4 s 158468 2176 158788 201824 6 vccd2
port 50 nsew power bidirectional
rlabel metal4 s 127748 2176 128068 201824 6 vccd2
port 51 nsew power bidirectional
rlabel metal4 s 97028 2176 97348 201824 6 vccd2
port 52 nsew power bidirectional
rlabel metal4 s 66308 2176 66628 201824 6 vccd2
port 53 nsew power bidirectional
rlabel metal4 s 35588 2176 35908 201824 6 vccd2
port 54 nsew power bidirectional
rlabel metal4 s 4868 2176 5188 201824 6 vccd2
port 55 nsew power bidirectional
rlabel metal4 s 235268 2176 235588 201824 6 vssd2
port 56 nsew ground bidirectional
rlabel metal4 s 204548 2176 204868 201824 6 vssd2
port 57 nsew ground bidirectional
rlabel metal4 s 173828 2176 174148 201824 6 vssd2
port 58 nsew ground bidirectional
rlabel metal4 s 143108 2176 143428 201824 6 vssd2
port 59 nsew ground bidirectional
rlabel metal4 s 112388 2176 112708 201824 6 vssd2
port 60 nsew ground bidirectional
rlabel metal4 s 81668 2176 81988 201824 6 vssd2
port 61 nsew ground bidirectional
rlabel metal4 s 50948 2176 51268 201824 6 vssd2
port 62 nsew ground bidirectional
rlabel metal4 s 20228 2176 20548 201824 6 vssd2
port 63 nsew ground bidirectional
rlabel metal4 s 220568 2176 220888 201824 6 vdda1
port 64 nsew power bidirectional
rlabel metal4 s 189848 2176 190168 201824 6 vdda1
port 65 nsew power bidirectional
rlabel metal4 s 159128 2176 159448 201824 6 vdda1
port 66 nsew power bidirectional
rlabel metal4 s 128408 2176 128728 201824 6 vdda1
port 67 nsew power bidirectional
rlabel metal4 s 97688 2176 98008 201824 6 vdda1
port 68 nsew power bidirectional
rlabel metal4 s 66968 2176 67288 201824 6 vdda1
port 69 nsew power bidirectional
rlabel metal4 s 36248 2176 36568 201824 6 vdda1
port 70 nsew power bidirectional
rlabel metal4 s 5528 2176 5848 201824 6 vdda1
port 71 nsew power bidirectional
rlabel metal4 s 235928 2176 236248 201824 6 vssa1
port 72 nsew ground bidirectional
rlabel metal4 s 205208 2176 205528 201824 6 vssa1
port 73 nsew ground bidirectional
rlabel metal4 s 174488 2176 174808 201824 6 vssa1
port 74 nsew ground bidirectional
rlabel metal4 s 143768 2176 144088 201824 6 vssa1
port 75 nsew ground bidirectional
rlabel metal4 s 113048 2176 113368 201824 6 vssa1
port 76 nsew ground bidirectional
rlabel metal4 s 82328 2176 82648 201824 6 vssa1
port 77 nsew ground bidirectional
rlabel metal4 s 51608 2176 51928 201824 6 vssa1
port 78 nsew ground bidirectional
rlabel metal4 s 20888 2176 21208 201824 6 vssa1
port 79 nsew ground bidirectional
rlabel metal4 s 221228 2176 221548 201824 6 vdda2
port 80 nsew power bidirectional
rlabel metal4 s 190508 2176 190828 201824 6 vdda2
port 81 nsew power bidirectional
rlabel metal4 s 159788 2176 160108 201824 6 vdda2
port 82 nsew power bidirectional
rlabel metal4 s 129068 2176 129388 201824 6 vdda2
port 83 nsew power bidirectional
rlabel metal4 s 98348 2176 98668 201824 6 vdda2
port 84 nsew power bidirectional
rlabel metal4 s 67628 2176 67948 201824 6 vdda2
port 85 nsew power bidirectional
rlabel metal4 s 36908 2176 37228 201824 6 vdda2
port 86 nsew power bidirectional
rlabel metal4 s 6188 2176 6508 201824 6 vdda2
port 87 nsew power bidirectional
rlabel metal4 s 236588 2176 236908 201824 6 vssa2
port 88 nsew ground bidirectional
rlabel metal4 s 205868 2176 206188 201824 6 vssa2
port 89 nsew ground bidirectional
rlabel metal4 s 175148 2176 175468 201824 6 vssa2
port 90 nsew ground bidirectional
rlabel metal4 s 144428 2176 144748 201824 6 vssa2
port 91 nsew ground bidirectional
rlabel metal4 s 113708 2176 114028 201824 6 vssa2
port 92 nsew ground bidirectional
rlabel metal4 s 82988 2176 83308 201824 6 vssa2
port 93 nsew ground bidirectional
rlabel metal4 s 52268 2176 52588 201824 6 vssa2
port 94 nsew ground bidirectional
rlabel metal4 s 21548 2176 21868 201824 6 vssa2
port 95 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 244000 204000
string LEFview TRUE
<< end >>

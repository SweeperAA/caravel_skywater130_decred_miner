magic
tech sky130A
magscale 1 2
timestamp 1608325398
<< locali >>
rect 14105 31195 14139 31433
rect 27261 29495 27295 29733
rect 39957 26435 39991 27217
rect 35633 19907 35667 20009
rect 10425 19159 10459 19261
rect 4445 18071 4479 18173
rect 15669 17527 15703 17765
rect 31217 15419 31251 15521
rect 17969 14263 18003 14569
rect 15393 11543 15427 11645
rect 32229 8891 32263 9129
rect 35265 6239 35299 6409
rect 36737 2975 36771 3077
<< viali >>
rect 11345 38505 11379 38539
rect 8309 38369 8343 38403
rect 8585 38369 8619 38403
rect 12817 38369 12851 38403
rect 14197 38369 14231 38403
rect 14749 38369 14783 38403
rect 15485 38369 15519 38403
rect 18797 38369 18831 38403
rect 19717 38369 19751 38403
rect 19809 38369 19843 38403
rect 20453 38369 20487 38403
rect 21649 38369 21683 38403
rect 22017 38369 22051 38403
rect 22385 38369 22419 38403
rect 26341 38369 26375 38403
rect 26985 38369 27019 38403
rect 27997 38369 28031 38403
rect 29837 38369 29871 38403
rect 30849 38369 30883 38403
rect 8401 38301 8435 38335
rect 9965 38301 9999 38335
rect 10241 38301 10275 38335
rect 14565 38301 14599 38335
rect 19533 38301 19567 38335
rect 24685 38301 24719 38335
rect 24961 38301 24995 38335
rect 26893 38301 26927 38335
rect 27905 38301 27939 38335
rect 29745 38301 29779 38335
rect 30757 38301 30791 38335
rect 12909 38165 12943 38199
rect 15577 38165 15611 38199
rect 18889 38165 18923 38199
rect 21741 38165 21775 38199
rect 27169 38165 27203 38199
rect 28181 38165 28215 38199
rect 30021 38165 30055 38199
rect 31033 38165 31067 38199
rect 4997 37961 5031 37995
rect 10885 37961 10919 37995
rect 16865 37961 16899 37995
rect 28457 37961 28491 37995
rect 31585 37961 31619 37995
rect 38853 37961 38887 37995
rect 10057 37893 10091 37927
rect 3617 37825 3651 37859
rect 6837 37825 6871 37859
rect 7941 37825 7975 37859
rect 8769 37825 8803 37859
rect 12449 37825 12483 37859
rect 12725 37825 12759 37859
rect 15485 37825 15519 37859
rect 20269 37825 20303 37859
rect 22569 37825 22603 37859
rect 23949 37825 23983 37859
rect 26433 37825 26467 37859
rect 33609 37825 33643 37859
rect 3893 37757 3927 37791
rect 7849 37757 7883 37791
rect 8493 37757 8527 37791
rect 10609 37757 10643 37791
rect 10701 37757 10735 37791
rect 14105 37757 14139 37791
rect 14565 37757 14599 37791
rect 15761 37757 15795 37791
rect 18613 37757 18647 37791
rect 18705 37757 18739 37791
rect 18981 37757 19015 37791
rect 19165 37757 19199 37791
rect 19441 37757 19475 37791
rect 20545 37757 20579 37791
rect 22661 37757 22695 37791
rect 23673 37757 23707 37791
rect 26157 37757 26191 37791
rect 28273 37757 28307 37791
rect 30021 37757 30055 37791
rect 30297 37757 30331 37791
rect 32229 37757 32263 37791
rect 32505 37757 32539 37791
rect 38669 37757 38703 37791
rect 23121 37689 23155 37723
rect 14657 37621 14691 37655
rect 18153 37621 18187 37655
rect 21649 37621 21683 37655
rect 25053 37621 25087 37655
rect 27537 37621 27571 37655
rect 29837 37621 29871 37655
rect 38485 37621 38519 37655
rect 9781 37417 9815 37451
rect 11897 37417 11931 37451
rect 18797 37417 18831 37451
rect 21005 37417 21039 37451
rect 21741 37417 21775 37451
rect 33701 37417 33735 37451
rect 35633 37417 35667 37451
rect 4629 37349 4663 37383
rect 17877 37349 17911 37383
rect 22293 37349 22327 37383
rect 4721 37281 4755 37315
rect 5181 37281 5215 37315
rect 5917 37281 5951 37315
rect 8125 37281 8159 37315
rect 8493 37281 8527 37315
rect 8677 37281 8711 37315
rect 9689 37281 9723 37315
rect 10609 37281 10643 37315
rect 12909 37281 12943 37315
rect 13829 37281 13863 37315
rect 14105 37281 14139 37315
rect 14473 37281 14507 37315
rect 15485 37281 15519 37315
rect 15577 37281 15611 37315
rect 16497 37281 16531 37315
rect 18521 37281 18555 37315
rect 19165 37281 19199 37315
rect 19533 37281 19567 37315
rect 19901 37281 19935 37315
rect 20913 37281 20947 37315
rect 21649 37281 21683 37315
rect 22845 37281 22879 37315
rect 22937 37281 22971 37315
rect 23213 37281 23247 37315
rect 23397 37281 23431 37315
rect 23581 37281 23615 37315
rect 24593 37281 24627 37315
rect 25973 37281 26007 37315
rect 27629 37281 27663 37315
rect 29469 37281 29503 37315
rect 29745 37281 29779 37315
rect 31125 37281 31159 37315
rect 32137 37281 32171 37315
rect 34253 37281 34287 37315
rect 34529 37281 34563 37315
rect 5641 37213 5675 37247
rect 8401 37213 8435 37247
rect 10333 37213 10367 37247
rect 14197 37213 14231 37247
rect 16221 37213 16255 37247
rect 24317 37213 24351 37247
rect 27353 37213 27387 37247
rect 32413 37213 32447 37247
rect 4445 37077 4479 37111
rect 7205 37077 7239 37111
rect 13001 37077 13035 37111
rect 28733 37077 28767 37111
rect 2789 36873 2823 36907
rect 21557 36873 21591 36907
rect 24593 36873 24627 36907
rect 28457 36873 28491 36907
rect 32781 36873 32815 36907
rect 16865 36805 16899 36839
rect 1409 36737 1443 36771
rect 4813 36737 4847 36771
rect 8125 36737 8159 36771
rect 11529 36737 11563 36771
rect 12909 36737 12943 36771
rect 14657 36737 14691 36771
rect 14933 36737 14967 36771
rect 18061 36737 18095 36771
rect 18337 36737 18371 36771
rect 25789 36737 25823 36771
rect 29285 36737 29319 36771
rect 29561 36737 29595 36771
rect 1685 36669 1719 36703
rect 5365 36669 5399 36703
rect 5549 36669 5583 36703
rect 5733 36669 5767 36703
rect 5917 36669 5951 36703
rect 6193 36669 6227 36703
rect 7113 36669 7147 36703
rect 7481 36669 7515 36703
rect 7849 36669 7883 36703
rect 8401 36669 8435 36703
rect 9873 36669 9907 36703
rect 10149 36669 10183 36703
rect 11437 36669 11471 36703
rect 11897 36669 11931 36703
rect 12449 36669 12483 36703
rect 12817 36669 12851 36703
rect 13185 36669 13219 36703
rect 16773 36669 16807 36703
rect 17509 36669 17543 36703
rect 20361 36669 20395 36703
rect 21741 36669 21775 36703
rect 21925 36669 21959 36703
rect 22293 36669 22327 36703
rect 22937 36669 22971 36703
rect 24317 36669 24351 36703
rect 24409 36669 24443 36703
rect 26065 36669 26099 36703
rect 28181 36669 28215 36703
rect 28273 36669 28307 36703
rect 32505 36669 32539 36703
rect 32597 36669 32631 36703
rect 16313 36601 16347 36635
rect 9873 36533 9907 36567
rect 19441 36533 19475 36567
rect 20453 36533 20487 36567
rect 27169 36533 27203 36567
rect 30665 36533 30699 36567
rect 8585 36329 8619 36363
rect 11069 36329 11103 36363
rect 13737 36261 13771 36295
rect 18245 36261 18279 36295
rect 27077 36261 27111 36295
rect 33425 36261 33459 36295
rect 4261 36193 4295 36227
rect 4813 36193 4847 36227
rect 6193 36193 6227 36227
rect 6377 36193 6411 36227
rect 6653 36193 6687 36227
rect 7389 36193 7423 36227
rect 7849 36193 7883 36227
rect 8493 36193 8527 36227
rect 9965 36193 9999 36227
rect 12817 36193 12851 36227
rect 13001 36193 13035 36227
rect 14565 36193 14599 36227
rect 15301 36193 15335 36227
rect 16405 36193 16439 36227
rect 16589 36193 16623 36227
rect 16865 36193 16899 36227
rect 18153 36193 18187 36227
rect 19073 36193 19107 36227
rect 19257 36193 19291 36227
rect 19625 36193 19659 36227
rect 19993 36193 20027 36227
rect 20269 36193 20303 36227
rect 21281 36193 21315 36227
rect 21741 36193 21775 36227
rect 22753 36193 22787 36227
rect 22845 36193 22879 36227
rect 23305 36193 23339 36227
rect 24041 36193 24075 36227
rect 26617 36193 26651 36227
rect 27813 36193 27847 36227
rect 30389 36193 30423 36227
rect 32873 36193 32907 36227
rect 32965 36193 32999 36227
rect 33977 36193 34011 36227
rect 34989 36193 35023 36227
rect 35081 36193 35115 36227
rect 5089 36125 5123 36159
rect 9689 36125 9723 36159
rect 13093 36125 13127 36159
rect 14289 36125 14323 36159
rect 14749 36125 14783 36159
rect 17325 36125 17359 36159
rect 21005 36125 21039 36159
rect 23765 36125 23799 36159
rect 26525 36125 26559 36159
rect 27537 36125 27571 36159
rect 30297 36125 30331 36159
rect 30849 36125 30883 36159
rect 33885 36125 33919 36159
rect 4353 36057 4387 36091
rect 6009 36057 6043 36091
rect 21741 36057 21775 36091
rect 7941 35989 7975 36023
rect 15393 35989 15427 36023
rect 22569 35989 22603 36023
rect 25329 35989 25363 36023
rect 28917 35989 28951 36023
rect 34161 35989 34195 36023
rect 35265 35989 35299 36023
rect 9229 35785 9263 35819
rect 16681 35785 16715 35819
rect 23857 35785 23891 35819
rect 27261 35785 27295 35819
rect 33609 35785 33643 35819
rect 36277 35785 36311 35819
rect 4721 35717 4755 35751
rect 11253 35717 11287 35751
rect 28457 35717 28491 35751
rect 4077 35649 4111 35683
rect 6285 35649 6319 35683
rect 7849 35649 7883 35683
rect 13001 35649 13035 35683
rect 16129 35649 16163 35683
rect 18797 35649 18831 35683
rect 29929 35649 29963 35683
rect 32045 35649 32079 35683
rect 32321 35649 32355 35683
rect 35173 35649 35207 35683
rect 4445 35581 4479 35615
rect 4721 35581 4755 35615
rect 5825 35581 5859 35615
rect 6101 35581 6135 35615
rect 6837 35581 6871 35615
rect 8125 35581 8159 35615
rect 10517 35581 10551 35615
rect 11161 35581 11195 35615
rect 11897 35581 11931 35615
rect 12449 35581 12483 35615
rect 13277 35581 13311 35615
rect 13461 35581 13495 35615
rect 14933 35581 14967 35615
rect 15577 35581 15611 35615
rect 15853 35581 15887 35615
rect 16773 35581 16807 35615
rect 17141 35581 17175 35615
rect 18245 35581 18279 35615
rect 18889 35581 18923 35615
rect 19625 35581 19659 35615
rect 20085 35581 20119 35615
rect 21557 35581 21591 35615
rect 21649 35581 21683 35615
rect 21833 35581 21867 35615
rect 22017 35581 22051 35615
rect 22385 35581 22419 35615
rect 23673 35581 23707 35615
rect 24777 35581 24811 35615
rect 25053 35581 25087 35615
rect 27445 35581 27479 35615
rect 27537 35581 27571 35615
rect 28273 35581 28307 35615
rect 29837 35581 29871 35615
rect 30205 35581 30239 35615
rect 34897 35581 34931 35615
rect 20361 35513 20395 35547
rect 21005 35513 21039 35547
rect 7021 35445 7055 35479
rect 10609 35445 10643 35479
rect 18337 35445 18371 35479
rect 26157 35445 26191 35479
rect 27721 35445 27755 35479
rect 29653 35445 29687 35479
rect 31309 35445 31343 35479
rect 10425 35241 10459 35275
rect 22109 35241 22143 35275
rect 27813 35241 27847 35275
rect 35633 35241 35667 35275
rect 9781 35173 9815 35207
rect 20913 35173 20947 35207
rect 21281 35173 21315 35207
rect 4077 35105 4111 35139
rect 4353 35105 4387 35139
rect 6193 35105 6227 35139
rect 7389 35105 7423 35139
rect 7757 35105 7791 35139
rect 8401 35105 8435 35139
rect 9689 35105 9723 35139
rect 10333 35105 10367 35139
rect 11253 35105 11287 35139
rect 13093 35105 13127 35139
rect 13645 35105 13679 35139
rect 15117 35105 15151 35139
rect 15945 35105 15979 35139
rect 16129 35105 16163 35139
rect 18521 35105 18555 35139
rect 18981 35105 19015 35139
rect 19349 35105 19383 35139
rect 19717 35105 19751 35139
rect 21097 35105 21131 35139
rect 21189 35105 21223 35139
rect 22301 35105 22335 35139
rect 22661 35105 22695 35139
rect 22937 35105 22971 35139
rect 23121 35105 23155 35139
rect 23673 35105 23707 35139
rect 24317 35105 24351 35139
rect 25513 35105 25547 35139
rect 26617 35105 26651 35139
rect 27629 35105 27663 35139
rect 28457 35105 28491 35139
rect 28917 35105 28951 35139
rect 29653 35105 29687 35139
rect 31953 35105 31987 35139
rect 32413 35105 32447 35139
rect 34529 35105 34563 35139
rect 38025 35105 38059 35139
rect 38209 35105 38243 35139
rect 8585 35037 8619 35071
rect 10977 35037 11011 35071
rect 16313 35037 16347 35071
rect 16865 35037 16899 35071
rect 17141 35037 17175 35071
rect 21649 35037 21683 35071
rect 22845 35037 22879 35071
rect 25421 35037 25455 35071
rect 25973 35037 26007 35071
rect 26525 35037 26559 35071
rect 28365 35037 28399 35071
rect 29377 35037 29411 35071
rect 32137 35037 32171 35071
rect 34253 35037 34287 35071
rect 6377 34969 6411 35003
rect 24409 34969 24443 35003
rect 31769 34969 31803 35003
rect 5641 34901 5675 34935
rect 12541 34901 12575 34935
rect 13185 34901 13219 34935
rect 14933 34901 14967 34935
rect 26801 34901 26835 34935
rect 30941 34901 30975 34935
rect 33517 34901 33551 34935
rect 38301 34901 38335 34935
rect 14473 34697 14507 34731
rect 17049 34697 17083 34731
rect 27721 34697 27755 34731
rect 30113 34697 30147 34731
rect 23857 34629 23891 34663
rect 28641 34629 28675 34663
rect 31033 34629 31067 34663
rect 6285 34561 6319 34595
rect 9229 34561 9263 34595
rect 15301 34561 15335 34595
rect 19257 34561 19291 34595
rect 24409 34561 24443 34595
rect 24961 34561 24995 34595
rect 26617 34561 26651 34595
rect 29837 34561 29871 34595
rect 31953 34561 31987 34595
rect 37105 34561 37139 34595
rect 38485 34561 38519 34595
rect 3893 34493 3927 34527
rect 5181 34493 5215 34527
rect 5733 34493 5767 34527
rect 6101 34493 6135 34527
rect 6837 34493 6871 34527
rect 7297 34493 7331 34527
rect 7665 34493 7699 34527
rect 8033 34493 8067 34527
rect 9505 34493 9539 34527
rect 10885 34493 10919 34527
rect 11345 34493 11379 34527
rect 12449 34493 12483 34527
rect 13369 34493 13403 34527
rect 13461 34493 13495 34527
rect 13829 34493 13863 34527
rect 14381 34493 14415 34527
rect 15025 34493 15059 34527
rect 15669 34493 15703 34527
rect 15853 34493 15887 34527
rect 16497 34493 16531 34527
rect 16957 34493 16991 34527
rect 18337 34493 18371 34527
rect 19165 34493 19199 34527
rect 20085 34493 20119 34527
rect 20545 34493 20579 34527
rect 20913 34493 20947 34527
rect 21925 34493 21959 34527
rect 22017 34493 22051 34527
rect 22661 34493 22695 34527
rect 22845 34493 22879 34527
rect 23121 34493 23155 34527
rect 23673 34493 23707 34527
rect 24501 34493 24535 34527
rect 26341 34493 26375 34527
rect 28457 34493 28491 34527
rect 29929 34493 29963 34527
rect 30849 34493 30883 34527
rect 31585 34493 31619 34527
rect 32229 34493 32263 34527
rect 32965 34493 32999 34527
rect 33149 34493 33183 34527
rect 33333 34493 33367 34527
rect 35357 34493 35391 34527
rect 36093 34493 36127 34527
rect 36369 34493 36403 34527
rect 37381 34493 37415 34527
rect 12541 34425 12575 34459
rect 4077 34357 4111 34391
rect 6929 34357 6963 34391
rect 11529 34357 11563 34391
rect 18613 34357 18647 34391
rect 19993 34357 20027 34391
rect 35449 34357 35483 34391
rect 7573 34153 7607 34187
rect 9045 34153 9079 34187
rect 17693 34153 17727 34187
rect 24041 34153 24075 34187
rect 37841 34153 37875 34187
rect 8125 34085 8159 34119
rect 25973 34085 26007 34119
rect 1593 34017 1627 34051
rect 4077 34017 4111 34051
rect 6745 34017 6779 34051
rect 7113 34017 7147 34051
rect 7297 34017 7331 34051
rect 8033 34017 8067 34051
rect 8953 34017 8987 34051
rect 9873 34017 9907 34051
rect 10793 34017 10827 34051
rect 11069 34017 11103 34051
rect 11529 34017 11563 34051
rect 11989 34017 12023 34051
rect 12725 34017 12759 34051
rect 12817 34017 12851 34051
rect 13185 34017 13219 34051
rect 13737 34017 13771 34051
rect 16037 34017 16071 34051
rect 16313 34017 16347 34051
rect 16957 34017 16991 34051
rect 17601 34017 17635 34051
rect 18429 34017 18463 34051
rect 18705 34017 18739 34051
rect 21189 34017 21223 34051
rect 21373 34017 21407 34051
rect 21649 34017 21683 34051
rect 22385 34017 22419 34051
rect 22845 34017 22879 34051
rect 23489 34017 23523 34051
rect 24225 34017 24259 34051
rect 24317 34017 24351 34051
rect 26525 34017 26559 34051
rect 26801 34017 26835 34051
rect 30849 34017 30883 34051
rect 32137 34017 32171 34051
rect 34253 34017 34287 34051
rect 34805 34017 34839 34051
rect 35449 34017 35483 34051
rect 35725 34017 35759 34051
rect 37749 34017 37783 34051
rect 38301 34017 38335 34051
rect 1869 33949 1903 33983
rect 4353 33949 4387 33983
rect 11161 33949 11195 33983
rect 15485 33949 15519 33983
rect 16497 33949 16531 33983
rect 23213 33949 23247 33983
rect 24593 33949 24627 33983
rect 28641 33949 28675 33983
rect 28917 33949 28951 33983
rect 30757 33949 30791 33983
rect 32413 33949 32447 33983
rect 38577 33949 38611 33983
rect 3157 33813 3191 33847
rect 5641 33813 5675 33847
rect 9965 33813 9999 33847
rect 12541 33813 12575 33847
rect 17049 33813 17083 33847
rect 19993 33813 20027 33847
rect 22293 33813 22327 33847
rect 27905 33813 27939 33847
rect 30205 33813 30239 33847
rect 31033 33813 31067 33847
rect 33517 33813 33551 33847
rect 34345 33813 34379 33847
rect 36829 33813 36863 33847
rect 5457 33609 5491 33643
rect 7297 33609 7331 33643
rect 10793 33609 10827 33643
rect 13829 33609 13863 33643
rect 14565 33609 14599 33643
rect 17233 33609 17267 33643
rect 21557 33609 21591 33643
rect 26065 33609 26099 33643
rect 28641 33609 28675 33643
rect 29561 33609 29595 33643
rect 30573 33609 30607 33643
rect 34069 33609 34103 33643
rect 1501 33541 1535 33575
rect 9965 33541 9999 33575
rect 22109 33541 22143 33575
rect 35817 33541 35851 33575
rect 38945 33541 38979 33575
rect 9321 33473 9355 33507
rect 12449 33473 12483 33507
rect 13185 33473 13219 33507
rect 15945 33473 15979 33507
rect 25145 33473 25179 33507
rect 25789 33473 25823 33507
rect 30297 33473 30331 33507
rect 31769 33473 31803 33507
rect 32689 33473 32723 33507
rect 32965 33473 32999 33507
rect 38301 33473 38335 33507
rect 1685 33405 1719 33439
rect 2145 33405 2179 33439
rect 2697 33405 2731 33439
rect 3341 33405 3375 33439
rect 3801 33405 3835 33439
rect 3893 33405 3927 33439
rect 4537 33405 4571 33439
rect 4997 33405 5031 33439
rect 5273 33405 5307 33439
rect 7205 33405 7239 33439
rect 8493 33405 8527 33439
rect 9689 33405 9723 33439
rect 10057 33405 10091 33439
rect 10977 33405 11011 33439
rect 11161 33405 11195 33439
rect 11529 33405 11563 33439
rect 12725 33405 12759 33439
rect 13645 33405 13679 33439
rect 14749 33405 14783 33439
rect 15209 33405 15243 33439
rect 15669 33405 15703 33439
rect 18245 33405 18279 33439
rect 18797 33405 18831 33439
rect 18981 33405 19015 33439
rect 19809 33405 19843 33439
rect 19993 33405 20027 33439
rect 20637 33405 20671 33439
rect 21005 33405 21039 33439
rect 21741 33405 21775 33439
rect 21833 33405 21867 33439
rect 22385 33405 22419 33439
rect 22845 33405 22879 33439
rect 23673 33405 23707 33439
rect 23949 33405 23983 33439
rect 25605 33405 25639 33439
rect 25881 33405 25915 33439
rect 27261 33405 27295 33439
rect 27445 33405 27479 33439
rect 27813 33405 27847 33439
rect 27905 33405 27939 33439
rect 28457 33405 28491 33439
rect 29285 33405 29319 33439
rect 29377 33405 29411 33439
rect 30389 33405 30423 33439
rect 31677 33405 31711 33439
rect 31953 33405 31987 33439
rect 34897 33405 34931 33439
rect 35265 33405 35299 33439
rect 35817 33405 35851 33439
rect 36461 33405 36495 33439
rect 37197 33405 37231 33439
rect 37749 33405 37783 33439
rect 38117 33405 38151 33439
rect 38761 33405 38795 33439
rect 2973 33337 3007 33371
rect 5181 33337 5215 33371
rect 12817 33337 12851 33371
rect 26801 33337 26835 33371
rect 8585 33269 8619 33303
rect 12633 33269 12667 33303
rect 18153 33269 18187 33303
rect 19625 33269 19659 33303
rect 20085 33269 20119 33303
rect 29929 33269 29963 33303
rect 36645 33269 36679 33303
rect 4905 33065 4939 33099
rect 16497 33065 16531 33099
rect 20085 33065 20119 33099
rect 21465 33065 21499 33099
rect 31769 33065 31803 33099
rect 2329 32997 2363 33031
rect 5089 32997 5123 33031
rect 10057 32997 10091 33031
rect 12449 32997 12483 33031
rect 15669 32997 15703 33031
rect 16037 32997 16071 33031
rect 35357 32997 35391 33031
rect 38301 32997 38335 33031
rect 2881 32929 2915 32963
rect 3157 32929 3191 32963
rect 3341 32929 3375 32963
rect 4997 32929 5031 32963
rect 6285 32929 6319 32963
rect 6377 32929 6411 32963
rect 6837 32929 6871 32963
rect 7205 32929 7239 32963
rect 7849 32929 7883 32963
rect 8585 32929 8619 32963
rect 9689 32929 9723 32963
rect 10425 32929 10459 32963
rect 10885 32929 10919 32963
rect 11069 32929 11103 32963
rect 11621 32929 11655 32963
rect 12265 32929 12299 32963
rect 12357 32929 12391 32963
rect 12817 32929 12851 32963
rect 14105 32929 14139 32963
rect 15485 32929 15519 32963
rect 15577 32929 15611 32963
rect 16681 32929 16715 32963
rect 16957 32929 16991 32963
rect 17509 32929 17543 32963
rect 17785 32929 17819 32963
rect 18337 32929 18371 32963
rect 19073 32929 19107 32963
rect 19349 32929 19383 32963
rect 19901 32929 19935 32963
rect 21557 32929 21591 32963
rect 22109 32929 22143 32963
rect 22937 32929 22971 32963
rect 23489 32929 23523 32963
rect 24961 32929 24995 32963
rect 25421 32929 25455 32963
rect 26525 32929 26559 32963
rect 29101 32929 29135 32963
rect 29929 32929 29963 32963
rect 31953 32929 31987 32963
rect 32505 32929 32539 32963
rect 32965 32929 32999 32963
rect 34253 32929 34287 32963
rect 34621 32929 34655 32963
rect 35173 32929 35207 32963
rect 36645 32929 36679 32963
rect 36921 32929 36955 32963
rect 38485 32929 38519 32963
rect 4721 32861 4755 32895
rect 5457 32861 5491 32895
rect 12081 32861 12115 32895
rect 13277 32861 13311 32895
rect 13829 32861 13863 32895
rect 14289 32861 14323 32895
rect 15301 32861 15335 32895
rect 22201 32861 22235 32895
rect 25053 32861 25087 32895
rect 27445 32861 27479 32895
rect 27721 32861 27755 32895
rect 29653 32861 29687 32895
rect 36277 32861 36311 32895
rect 38761 32861 38795 32895
rect 5917 32793 5951 32827
rect 16865 32793 16899 32827
rect 18613 32793 18647 32827
rect 32321 32793 32355 32827
rect 36921 32793 36955 32827
rect 8769 32725 8803 32759
rect 23029 32725 23063 32759
rect 26709 32725 26743 32759
rect 31033 32725 31067 32759
rect 6193 32521 6227 32555
rect 8217 32521 8251 32555
rect 17049 32521 17083 32555
rect 24501 32521 24535 32555
rect 39037 32521 39071 32555
rect 12725 32453 12759 32487
rect 13277 32453 13311 32487
rect 18889 32453 18923 32487
rect 35725 32453 35759 32487
rect 2513 32385 2547 32419
rect 3341 32385 3375 32419
rect 9229 32385 9263 32419
rect 10609 32385 10643 32419
rect 13645 32385 13679 32419
rect 15669 32385 15703 32419
rect 15945 32385 15979 32419
rect 20453 32385 20487 32419
rect 22569 32385 22603 32419
rect 30849 32385 30883 32419
rect 31585 32385 31619 32419
rect 36921 32385 36955 32419
rect 1961 32317 1995 32351
rect 2973 32317 3007 32351
rect 3525 32317 3559 32351
rect 4169 32317 4203 32351
rect 4813 32317 4847 32351
rect 5365 32317 5399 32351
rect 5549 32317 5583 32351
rect 6101 32317 6135 32351
rect 6837 32317 6871 32351
rect 7113 32317 7147 32351
rect 8953 32317 8987 32351
rect 11621 32317 11655 32351
rect 12541 32317 12575 32351
rect 14013 32317 14047 32351
rect 14381 32317 14415 32351
rect 14565 32317 14599 32351
rect 14933 32317 14967 32351
rect 18245 32317 18279 32351
rect 18613 32317 18647 32351
rect 18981 32317 19015 32351
rect 19625 32317 19659 32351
rect 20361 32317 20395 32351
rect 21925 32317 21959 32351
rect 22477 32317 22511 32351
rect 23673 32317 23707 32351
rect 24409 32317 24443 32351
rect 25329 32317 25363 32351
rect 25605 32317 25639 32351
rect 27169 32317 27203 32351
rect 27353 32317 27387 32351
rect 27721 32317 27755 32351
rect 27905 32317 27939 32351
rect 28365 32317 28399 32351
rect 29469 32317 29503 32351
rect 29745 32317 29779 32351
rect 31677 32317 31711 32351
rect 32781 32317 32815 32351
rect 32965 32317 32999 32351
rect 33333 32317 33367 32351
rect 34897 32317 34931 32351
rect 35357 32317 35391 32351
rect 35817 32317 35851 32351
rect 36645 32317 36679 32351
rect 37473 32317 37507 32351
rect 37749 32317 37783 32351
rect 1777 32249 1811 32283
rect 2145 32249 2179 32283
rect 4261 32249 4295 32283
rect 32137 32249 32171 32283
rect 36461 32249 36495 32283
rect 2053 32181 2087 32215
rect 11805 32181 11839 32215
rect 19717 32181 19751 32215
rect 21833 32181 21867 32215
rect 23857 32181 23891 32215
rect 25145 32181 25179 32215
rect 26801 32181 26835 32215
rect 28549 32181 28583 32215
rect 3709 31977 3743 32011
rect 7205 31977 7239 32011
rect 9045 31977 9079 32011
rect 22569 31977 22603 32011
rect 33793 31977 33827 32011
rect 36369 31977 36403 32011
rect 4353 31909 4387 31943
rect 18429 31909 18463 31943
rect 30849 31909 30883 31943
rect 1409 31841 1443 31875
rect 3893 31841 3927 31875
rect 4813 31841 4847 31875
rect 4997 31841 5031 31875
rect 5181 31841 5215 31875
rect 5365 31841 5399 31875
rect 5641 31841 5675 31875
rect 6561 31841 6595 31875
rect 6929 31841 6963 31875
rect 7113 31841 7147 31875
rect 8217 31841 8251 31875
rect 8861 31841 8895 31875
rect 9689 31841 9723 31875
rect 10057 31841 10091 31875
rect 10517 31841 10551 31875
rect 12265 31841 12299 31875
rect 12633 31841 12667 31875
rect 13185 31841 13219 31875
rect 13369 31841 13403 31875
rect 14565 31841 14599 31875
rect 15301 31841 15335 31875
rect 16221 31841 16255 31875
rect 16681 31841 16715 31875
rect 17049 31841 17083 31875
rect 17233 31841 17267 31875
rect 17969 31841 18003 31875
rect 18705 31841 18739 31875
rect 18981 31841 19015 31875
rect 19441 31841 19475 31875
rect 19901 31841 19935 31875
rect 20361 31841 20395 31875
rect 21281 31841 21315 31875
rect 21833 31841 21867 31875
rect 22477 31841 22511 31875
rect 23673 31841 23707 31875
rect 24041 31841 24075 31875
rect 25421 31841 25455 31875
rect 25743 31841 25777 31875
rect 25973 31841 26007 31875
rect 26985 31841 27019 31875
rect 27169 31841 27203 31875
rect 27537 31841 27571 31875
rect 27721 31841 27755 31875
rect 28181 31841 28215 31875
rect 28273 31841 28307 31875
rect 29561 31841 29595 31875
rect 30021 31841 30055 31875
rect 30481 31841 30515 31875
rect 30665 31841 30699 31875
rect 30757 31841 30791 31875
rect 38025 31841 38059 31875
rect 38393 31841 38427 31875
rect 38761 31841 38795 31875
rect 1685 31773 1719 31807
rect 8309 31773 8343 31807
rect 11713 31773 11747 31807
rect 12081 31773 12115 31807
rect 14657 31773 14691 31807
rect 16313 31773 16347 31807
rect 21097 31773 21131 31807
rect 23305 31773 23339 31807
rect 24777 31773 24811 31807
rect 25513 31773 25547 31807
rect 26525 31773 26559 31807
rect 29653 31773 29687 31807
rect 31217 31773 31251 31807
rect 32229 31773 32263 31807
rect 32505 31773 32539 31807
rect 34989 31773 35023 31807
rect 35265 31773 35299 31807
rect 38669 31773 38703 31807
rect 9781 31705 9815 31739
rect 21741 31705 21775 31739
rect 23949 31705 23983 31739
rect 2973 31637 3007 31671
rect 15485 31637 15519 31671
rect 28457 31637 28491 31671
rect 1685 31433 1719 31467
rect 14105 31433 14139 31467
rect 14381 31433 14415 31467
rect 17141 31433 17175 31467
rect 35173 31433 35207 31467
rect 2881 31297 2915 31331
rect 7481 31297 7515 31331
rect 10333 31297 10367 31331
rect 13001 31297 13035 31331
rect 13461 31297 13495 31331
rect 1593 31229 1627 31263
rect 2513 31229 2547 31263
rect 2697 31229 2731 31263
rect 3249 31229 3283 31263
rect 3709 31229 3743 31263
rect 4353 31229 4387 31263
rect 4997 31229 5031 31263
rect 5365 31229 5399 31263
rect 6009 31229 6043 31263
rect 6837 31229 6871 31263
rect 7757 31229 7791 31263
rect 9873 31229 9907 31263
rect 10149 31229 10183 31263
rect 10793 31229 10827 31263
rect 11253 31229 11287 31263
rect 11621 31229 11655 31263
rect 13277 31229 13311 31263
rect 22845 31365 22879 31399
rect 23949 31365 23983 31399
rect 25329 31365 25363 31399
rect 32413 31365 32447 31399
rect 15301 31297 15335 31331
rect 19441 31297 19475 31331
rect 22201 31297 22235 31331
rect 24685 31297 24719 31331
rect 29745 31297 29779 31331
rect 31769 31297 31803 31331
rect 36737 31297 36771 31331
rect 14197 31229 14231 31263
rect 15025 31229 15059 31263
rect 17325 31229 17359 31263
rect 19349 31229 19383 31263
rect 19809 31229 19843 31263
rect 19993 31229 20027 31263
rect 20361 31229 20395 31263
rect 21097 31229 21131 31263
rect 22569 31229 22603 31263
rect 22937 31229 22971 31263
rect 23673 31229 23707 31263
rect 24225 31229 24259 31263
rect 25237 31229 25271 31263
rect 25789 31229 25823 31263
rect 26525 31229 26559 31263
rect 26709 31229 26743 31263
rect 27169 31229 27203 31263
rect 27261 31229 27295 31263
rect 28365 31229 28399 31263
rect 29469 31229 29503 31263
rect 31953 31229 31987 31263
rect 32413 31229 32447 31263
rect 33425 31229 33459 31263
rect 33793 31229 33827 31263
rect 34161 31229 34195 31263
rect 34989 31229 35023 31263
rect 36001 31229 36035 31263
rect 36461 31229 36495 31263
rect 36829 31229 36863 31263
rect 37473 31229 37507 31263
rect 37749 31229 37783 31263
rect 9137 31161 9171 31195
rect 12449 31161 12483 31195
rect 14105 31161 14139 31195
rect 34345 31161 34379 31195
rect 4445 31093 4479 31127
rect 6193 31093 6227 31127
rect 6929 31093 6963 31127
rect 11897 31093 11931 31127
rect 16405 31093 16439 31127
rect 27721 31093 27755 31127
rect 28549 31093 28583 31127
rect 30849 31093 30883 31127
rect 38853 31093 38887 31127
rect 7021 30889 7055 30923
rect 10425 30889 10459 30923
rect 12357 30889 12391 30923
rect 23765 30889 23799 30923
rect 34069 30889 34103 30923
rect 35081 30889 35115 30923
rect 36921 30889 36955 30923
rect 37841 30889 37875 30923
rect 2513 30821 2547 30855
rect 9781 30821 9815 30855
rect 29653 30821 29687 30855
rect 3341 30753 3375 30787
rect 3525 30753 3559 30787
rect 4353 30753 4387 30787
rect 4905 30753 4939 30787
rect 5181 30753 5215 30787
rect 5917 30753 5951 30787
rect 8217 30753 8251 30787
rect 8677 30753 8711 30787
rect 9505 30753 9539 30787
rect 9689 30753 9723 30787
rect 10333 30753 10367 30787
rect 10793 30753 10827 30787
rect 11161 30753 11195 30787
rect 11529 30753 11563 30787
rect 12265 30753 12299 30787
rect 13553 30753 13587 30787
rect 13829 30753 13863 30787
rect 14013 30753 14047 30787
rect 14749 30753 14783 30787
rect 16129 30753 16163 30787
rect 17049 30753 17083 30787
rect 17233 30753 17267 30787
rect 17601 30753 17635 30787
rect 17969 30753 18003 30787
rect 18705 30753 18739 30787
rect 19349 30753 19383 30787
rect 19717 30753 19751 30787
rect 20085 30753 20119 30787
rect 21649 30753 21683 30787
rect 22385 30753 22419 30787
rect 23673 30753 23707 30787
rect 24225 30753 24259 30787
rect 25237 30753 25271 30787
rect 25789 30753 25823 30787
rect 26893 30753 26927 30787
rect 27077 30753 27111 30787
rect 30389 30753 30423 30787
rect 30849 30753 30883 30787
rect 31401 30753 31435 30787
rect 31585 30753 31619 30787
rect 32965 30753 32999 30787
rect 35173 30753 35207 30787
rect 35725 30753 35759 30787
rect 36645 30753 36679 30787
rect 36829 30753 36863 30787
rect 37749 30753 37783 30787
rect 38485 30753 38519 30787
rect 3065 30685 3099 30719
rect 4997 30685 5031 30719
rect 5641 30685 5675 30719
rect 8493 30685 8527 30719
rect 15301 30685 15335 30719
rect 15853 30685 15887 30719
rect 16313 30685 16347 30719
rect 22477 30685 22511 30719
rect 24685 30685 24719 30719
rect 26985 30685 27019 30719
rect 27537 30685 27571 30719
rect 27997 30685 28031 30719
rect 28273 30685 28307 30719
rect 30573 30685 30607 30719
rect 32689 30685 32723 30719
rect 35817 30685 35851 30719
rect 38577 30685 38611 30719
rect 17049 30617 17083 30651
rect 19993 30617 20027 30651
rect 21925 30617 21959 30651
rect 25329 30617 25363 30651
rect 9321 30549 9355 30583
rect 14657 30549 14691 30583
rect 30205 30549 30239 30583
rect 7113 30345 7147 30379
rect 8953 30345 8987 30379
rect 28641 30345 28675 30379
rect 32965 30345 32999 30379
rect 34253 30345 34287 30379
rect 17325 30277 17359 30311
rect 22661 30277 22695 30311
rect 31953 30277 31987 30311
rect 35817 30277 35851 30311
rect 4353 30209 4387 30243
rect 10517 30209 10551 30243
rect 12725 30209 12759 30243
rect 14657 30209 14691 30243
rect 15393 30209 15427 30243
rect 16589 30209 16623 30243
rect 19625 30209 19659 30243
rect 24501 30209 24535 30243
rect 25881 30209 25915 30243
rect 26341 30209 26375 30243
rect 30573 30209 30607 30243
rect 37473 30209 37507 30243
rect 39129 30209 39163 30243
rect 2789 30141 2823 30175
rect 2973 30141 3007 30175
rect 3249 30141 3283 30175
rect 3433 30141 3467 30175
rect 3617 30141 3651 30175
rect 4261 30141 4295 30175
rect 4629 30141 4663 30175
rect 4997 30141 5031 30175
rect 5549 30141 5583 30175
rect 6377 30141 6411 30175
rect 7021 30141 7055 30175
rect 7941 30141 7975 30175
rect 8033 30141 8067 30175
rect 8401 30141 8435 30175
rect 9045 30141 9079 30175
rect 9229 30141 9263 30175
rect 9873 30141 9907 30175
rect 10977 30141 11011 30175
rect 11161 30141 11195 30175
rect 11345 30141 11379 30175
rect 12449 30141 12483 30175
rect 16957 30141 16991 30175
rect 17325 30141 17359 30175
rect 19533 30141 19567 30175
rect 19809 30141 19843 30175
rect 20177 30141 20211 30175
rect 20545 30141 20579 30175
rect 21281 30141 21315 30175
rect 21741 30141 21775 30175
rect 22109 30141 22143 30175
rect 22569 30141 22603 30175
rect 23673 30141 23707 30175
rect 24225 30141 24259 30175
rect 25421 30141 25455 30175
rect 26065 30141 26099 30175
rect 26433 30141 26467 30175
rect 27353 30141 27387 30175
rect 27629 30141 27663 30175
rect 28457 30141 28491 30175
rect 29837 30141 29871 30175
rect 31217 30141 31251 30175
rect 31401 30141 31435 30175
rect 31953 30141 31987 30175
rect 32781 30141 32815 30175
rect 33057 30141 33091 30175
rect 33517 30141 33551 30175
rect 34069 30141 34103 30175
rect 34897 30141 34931 30175
rect 35449 30141 35483 30175
rect 35817 30141 35851 30175
rect 36645 30141 36679 30175
rect 37749 30141 37783 30175
rect 2329 30073 2363 30107
rect 14841 30073 14875 30107
rect 15025 30073 15059 30107
rect 27445 30073 27479 30107
rect 30205 30073 30239 30107
rect 36461 30073 36495 30107
rect 37013 30073 37047 30107
rect 6193 30005 6227 30039
rect 14013 30005 14047 30039
rect 14933 30005 14967 30039
rect 23765 30005 23799 30039
rect 27169 30005 27203 30039
rect 27721 30005 27755 30039
rect 30021 30005 30055 30039
rect 30113 30005 30147 30039
rect 32597 30005 32631 30039
rect 2789 29801 2823 29835
rect 6009 29801 6043 29835
rect 9781 29801 9815 29835
rect 30757 29801 30791 29835
rect 32413 29801 32447 29835
rect 8125 29733 8159 29767
rect 27261 29733 27295 29767
rect 30849 29733 30883 29767
rect 31217 29733 31251 29767
rect 1409 29665 1443 29699
rect 4077 29665 4111 29699
rect 4813 29665 4847 29699
rect 5549 29665 5583 29699
rect 5825 29665 5859 29699
rect 6009 29665 6043 29699
rect 6745 29665 6779 29699
rect 7389 29665 7423 29699
rect 8677 29665 8711 29699
rect 8953 29665 8987 29699
rect 9965 29665 9999 29699
rect 10517 29665 10551 29699
rect 10701 29665 10735 29699
rect 11253 29665 11287 29699
rect 11805 29665 11839 29699
rect 12265 29665 12299 29699
rect 12817 29665 12851 29699
rect 13461 29665 13495 29699
rect 14289 29665 14323 29699
rect 14473 29665 14507 29699
rect 15301 29665 15335 29699
rect 15853 29665 15887 29699
rect 16681 29665 16715 29699
rect 17417 29665 17451 29699
rect 18245 29665 18279 29699
rect 18889 29665 18923 29699
rect 19073 29665 19107 29699
rect 19809 29665 19843 29699
rect 20913 29665 20947 29699
rect 21741 29665 21775 29699
rect 22569 29665 22603 29699
rect 22937 29665 22971 29699
rect 23213 29665 23247 29699
rect 24133 29665 24167 29699
rect 24685 29665 24719 29699
rect 25513 29665 25547 29699
rect 26525 29665 26559 29699
rect 1685 29597 1719 29631
rect 6837 29597 6871 29631
rect 9137 29597 9171 29631
rect 14565 29597 14599 29631
rect 15669 29597 15703 29631
rect 17509 29597 17543 29631
rect 24777 29597 24811 29631
rect 11345 29529 11379 29563
rect 12909 29529 12943 29563
rect 16957 29529 16991 29563
rect 18429 29529 18463 29563
rect 19993 29529 20027 29563
rect 21097 29529 21131 29563
rect 23305 29529 23339 29563
rect 24225 29529 24259 29563
rect 25697 29529 25731 29563
rect 27629 29665 27663 29699
rect 29469 29665 29503 29699
rect 29561 29665 29595 29699
rect 30665 29665 30699 29699
rect 32229 29665 32263 29699
rect 32965 29665 32999 29699
rect 35541 29665 35575 29699
rect 37749 29665 37783 29699
rect 38117 29665 38151 29699
rect 38577 29665 38611 29699
rect 27353 29597 27387 29631
rect 30481 29597 30515 29631
rect 33241 29597 33275 29631
rect 35817 29597 35851 29631
rect 38577 29529 38611 29563
rect 4261 29461 4295 29495
rect 7481 29461 7515 29495
rect 21833 29461 21867 29495
rect 26709 29461 26743 29495
rect 27261 29461 27295 29495
rect 28917 29461 28951 29495
rect 29745 29461 29779 29495
rect 34529 29461 34563 29495
rect 36921 29461 36955 29495
rect 1501 29257 1535 29291
rect 1961 29257 1995 29291
rect 7021 29257 7055 29291
rect 11437 29257 11471 29291
rect 21189 29257 21223 29291
rect 25513 29257 25547 29291
rect 27169 29257 27203 29291
rect 38761 29257 38795 29291
rect 17417 29189 17451 29223
rect 18981 29189 19015 29223
rect 24409 29189 24443 29223
rect 27997 29189 28031 29223
rect 30665 29189 30699 29223
rect 33057 29189 33091 29223
rect 35725 29189 35759 29223
rect 37289 29189 37323 29223
rect 2697 29121 2731 29155
rect 3433 29121 3467 29155
rect 4629 29121 4663 29155
rect 5733 29121 5767 29155
rect 7573 29121 7607 29155
rect 9781 29121 9815 29155
rect 15853 29121 15887 29155
rect 19993 29121 20027 29155
rect 36461 29121 36495 29155
rect 1777 29053 1811 29087
rect 2881 29053 2915 29087
rect 2973 29053 3007 29087
rect 4169 29053 4203 29087
rect 4445 29053 4479 29087
rect 5273 29053 5307 29087
rect 5549 29053 5583 29087
rect 6101 29053 6135 29087
rect 6837 29053 6871 29087
rect 7849 29053 7883 29087
rect 9965 29053 9999 29087
rect 10149 29053 10183 29087
rect 10425 29053 10459 29087
rect 11345 29053 11379 29087
rect 13277 29053 13311 29087
rect 13553 29053 13587 29087
rect 13737 29053 13771 29087
rect 14197 29053 14231 29087
rect 14289 29053 14323 29087
rect 14933 29053 14967 29087
rect 15485 29053 15519 29087
rect 16313 29053 16347 29087
rect 16589 29053 16623 29087
rect 17233 29053 17267 29087
rect 18061 29053 18095 29087
rect 18429 29053 18463 29087
rect 18889 29053 18923 29087
rect 19625 29053 19659 29087
rect 20361 29053 20395 29087
rect 21741 29053 21775 29087
rect 21833 29053 21867 29087
rect 22109 29053 22143 29087
rect 22293 29053 22327 29087
rect 22937 29053 22971 29087
rect 23949 29053 23983 29087
rect 24501 29053 24535 29087
rect 24685 29053 24719 29087
rect 25329 29053 25363 29087
rect 26065 29053 26099 29087
rect 26198 29053 26232 29087
rect 26617 29053 26651 29087
rect 27077 29053 27111 29087
rect 28181 29053 28215 29087
rect 28549 29053 28583 29087
rect 28641 29053 28675 29087
rect 29285 29053 29319 29087
rect 29561 29053 29595 29087
rect 31861 29053 31895 29087
rect 32137 29053 32171 29087
rect 32321 29053 32355 29087
rect 32781 29053 32815 29087
rect 33333 29053 33367 29087
rect 33793 29053 33827 29087
rect 35449 29053 35483 29087
rect 36185 29053 36219 29087
rect 37013 29053 37047 29087
rect 37749 29053 37783 29087
rect 37841 29053 37875 29087
rect 38577 29053 38611 29087
rect 1685 28985 1719 29019
rect 3065 28985 3099 29019
rect 9229 28985 9263 29019
rect 12725 28985 12759 29019
rect 23029 28917 23063 28951
rect 3249 28713 3283 28747
rect 4813 28713 4847 28747
rect 7481 28713 7515 28747
rect 8309 28713 8343 28747
rect 9045 28713 9079 28747
rect 29929 28713 29963 28747
rect 12265 28645 12299 28679
rect 17969 28645 18003 28679
rect 24041 28645 24075 28679
rect 31493 28645 31527 28679
rect 36369 28645 36403 28679
rect 4629 28577 4663 28611
rect 5365 28577 5399 28611
rect 6377 28577 6411 28611
rect 8217 28577 8251 28611
rect 8953 28577 8987 28611
rect 9689 28577 9723 28611
rect 10885 28577 10919 28611
rect 15301 28577 15335 28611
rect 15669 28577 15703 28611
rect 16589 28577 16623 28611
rect 16957 28577 16991 28611
rect 17877 28577 17911 28611
rect 18245 28577 18279 28611
rect 18705 28577 18739 28611
rect 19073 28577 19107 28611
rect 19533 28577 19567 28611
rect 19993 28577 20027 28611
rect 20913 28577 20947 28611
rect 21649 28577 21683 28611
rect 22109 28577 22143 28611
rect 22661 28577 22695 28611
rect 22845 28577 22879 28611
rect 23489 28577 23523 28611
rect 24501 28577 24535 28611
rect 24869 28577 24903 28611
rect 24961 28577 24995 28611
rect 25697 28577 25731 28611
rect 26893 28577 26927 28611
rect 27445 28577 27479 28611
rect 28273 28577 28307 28611
rect 28825 28577 28859 28611
rect 29285 28577 29319 28611
rect 30113 28577 30147 28611
rect 30389 28577 30423 28611
rect 30665 28577 30699 28611
rect 31401 28577 31435 28611
rect 32229 28577 32263 28611
rect 33149 28577 33183 28611
rect 35725 28577 35759 28611
rect 36093 28577 36127 28611
rect 36829 28577 36863 28611
rect 38117 28577 38151 28611
rect 38301 28577 38335 28611
rect 38761 28577 38795 28611
rect 1685 28509 1719 28543
rect 1961 28509 1995 28543
rect 5457 28509 5491 28543
rect 6101 28509 6135 28543
rect 10609 28509 10643 28543
rect 13093 28509 13127 28543
rect 13369 28509 13403 28543
rect 26617 28509 26651 28543
rect 27353 28509 27387 28543
rect 32137 28509 32171 28543
rect 33425 28509 33459 28543
rect 35357 28509 35391 28543
rect 16221 28441 16255 28475
rect 21741 28441 21775 28475
rect 28549 28441 28583 28475
rect 38761 28441 38795 28475
rect 9873 28373 9907 28407
rect 14473 28373 14507 28407
rect 20177 28373 20211 28407
rect 21097 28373 21131 28407
rect 25881 28373 25915 28407
rect 32413 28373 32447 28407
rect 34529 28373 34563 28407
rect 37013 28373 37047 28407
rect 1685 28169 1719 28203
rect 8033 28169 8067 28203
rect 9229 28169 9263 28203
rect 11345 28169 11379 28203
rect 12633 28169 12667 28203
rect 15209 28169 15243 28203
rect 25513 28169 25547 28203
rect 29561 28169 29595 28203
rect 34161 28169 34195 28203
rect 36737 28169 36771 28203
rect 2329 28101 2363 28135
rect 5273 28101 5307 28135
rect 6193 28101 6227 28135
rect 6929 28101 6963 28135
rect 13829 28101 13863 28135
rect 24133 28101 24167 28135
rect 28641 28101 28675 28135
rect 10701 28033 10735 28067
rect 14565 28033 14599 28067
rect 16681 28033 16715 28067
rect 18705 28033 18739 28067
rect 20637 28033 20671 28067
rect 27813 28033 27847 28067
rect 29285 28033 29319 28067
rect 30297 28033 30331 28067
rect 30573 28033 30607 28067
rect 33425 28033 33459 28067
rect 35173 28033 35207 28067
rect 37565 28033 37599 28067
rect 1593 27965 1627 27999
rect 2237 27965 2271 27999
rect 3065 27965 3099 27999
rect 3433 27965 3467 27999
rect 3801 27965 3835 27999
rect 4445 27965 4479 27999
rect 4997 27965 5031 27999
rect 5365 27965 5399 27999
rect 6009 27965 6043 27999
rect 7113 27965 7147 27999
rect 7389 27965 7423 27999
rect 8217 27965 8251 27999
rect 8309 27965 8343 27999
rect 9045 27965 9079 27999
rect 9873 27965 9907 27999
rect 10241 27965 10275 27999
rect 10609 27965 10643 27999
rect 11529 27965 11563 27999
rect 11713 27965 11747 27999
rect 12449 27965 12483 27999
rect 13553 27965 13587 27999
rect 14289 27965 14323 27999
rect 15117 27965 15151 27999
rect 15853 27965 15887 27999
rect 16497 27965 16531 27999
rect 18337 27965 18371 27999
rect 18521 27965 18555 27999
rect 19165 27965 19199 27999
rect 19349 27965 19383 27999
rect 19717 27965 19751 27999
rect 20545 27965 20579 27999
rect 21189 27965 21223 27999
rect 21373 27965 21407 27999
rect 21925 27965 21959 27999
rect 22293 27965 22327 27999
rect 22937 27965 22971 27999
rect 23949 27965 23983 27999
rect 24691 27965 24725 27999
rect 25421 27965 25455 27999
rect 25973 27965 26007 27999
rect 26433 27965 26467 27999
rect 27353 27965 27387 27999
rect 28457 27965 28491 27999
rect 29377 27965 29411 27999
rect 32597 27965 32631 27999
rect 32781 27965 32815 27999
rect 33333 27965 33367 27999
rect 33977 27965 34011 27999
rect 35449 27965 35483 27999
rect 37289 27965 37323 27999
rect 3985 27897 4019 27931
rect 23029 27897 23063 27931
rect 27077 27897 27111 27931
rect 27445 27897 27479 27931
rect 8493 27829 8527 27863
rect 11805 27829 11839 27863
rect 15945 27829 15979 27863
rect 24869 27829 24903 27863
rect 27261 27829 27295 27863
rect 31861 27829 31895 27863
rect 38669 27829 38703 27863
rect 4169 27625 4203 27659
rect 1777 27557 1811 27591
rect 7113 27557 7147 27591
rect 10885 27557 10919 27591
rect 15393 27557 15427 27591
rect 16129 27557 16163 27591
rect 27445 27557 27479 27591
rect 27813 27557 27847 27591
rect 28181 27557 28215 27591
rect 36645 27557 36679 27591
rect 37197 27557 37231 27591
rect 1685 27489 1719 27523
rect 2513 27489 2547 27523
rect 2605 27489 2639 27523
rect 3893 27489 3927 27523
rect 4077 27489 4111 27523
rect 4629 27489 4663 27523
rect 4997 27489 5031 27523
rect 5641 27489 5675 27523
rect 6285 27489 6319 27523
rect 7665 27489 7699 27523
rect 7941 27489 7975 27523
rect 8861 27489 8895 27523
rect 10241 27489 10275 27523
rect 10609 27489 10643 27523
rect 11345 27489 11379 27523
rect 12081 27489 12115 27523
rect 12449 27489 12483 27523
rect 13093 27489 13127 27523
rect 13369 27489 13403 27523
rect 14013 27489 14047 27523
rect 14381 27489 14415 27523
rect 14565 27489 14599 27523
rect 15301 27489 15335 27523
rect 16773 27489 16807 27523
rect 17141 27489 17175 27523
rect 17785 27489 17819 27523
rect 18521 27489 18555 27523
rect 19809 27489 19843 27523
rect 20085 27489 20119 27523
rect 21097 27489 21131 27523
rect 21557 27489 21591 27523
rect 22477 27489 22511 27523
rect 23673 27489 23707 27523
rect 24225 27489 24259 27523
rect 25145 27489 25179 27523
rect 25605 27489 25639 27523
rect 26709 27489 26743 27523
rect 27629 27489 27663 27523
rect 27721 27489 27755 27523
rect 28917 27489 28951 27523
rect 29101 27489 29135 27523
rect 29469 27489 29503 27523
rect 30665 27489 30699 27523
rect 32413 27489 32447 27523
rect 33241 27489 33275 27523
rect 33425 27489 33459 27523
rect 33793 27489 33827 27523
rect 34253 27489 34287 27523
rect 35541 27489 35575 27523
rect 35817 27489 35851 27523
rect 36829 27489 36863 27523
rect 38025 27489 38059 27523
rect 38301 27489 38335 27523
rect 38669 27489 38703 27523
rect 8125 27421 8159 27455
rect 9965 27421 9999 27455
rect 13461 27421 13495 27455
rect 16865 27421 16899 27455
rect 17233 27421 17267 27455
rect 19349 27421 19383 27455
rect 20361 27421 20395 27455
rect 21925 27421 21959 27455
rect 23489 27421 23523 27455
rect 30812 27421 30846 27455
rect 31033 27421 31067 27455
rect 35081 27421 35115 27455
rect 3709 27353 3743 27387
rect 17877 27353 17911 27387
rect 21005 27353 21039 27387
rect 22661 27353 22695 27387
rect 24133 27353 24167 27387
rect 24961 27353 24995 27387
rect 29469 27353 29503 27387
rect 30941 27353 30975 27387
rect 32505 27353 32539 27387
rect 35909 27353 35943 27387
rect 38669 27353 38703 27387
rect 2329 27285 2363 27319
rect 2789 27285 2823 27319
rect 5733 27285 5767 27319
rect 6469 27285 6503 27319
rect 9045 27285 9079 27319
rect 11529 27285 11563 27319
rect 26893 27285 26927 27319
rect 31125 27285 31159 27319
rect 34437 27285 34471 27319
rect 39957 27217 39991 27251
rect 5089 27081 5123 27115
rect 6193 27081 6227 27115
rect 9597 27081 9631 27115
rect 25973 27081 26007 27115
rect 29634 27081 29668 27115
rect 32045 27081 32079 27115
rect 35173 27081 35207 27115
rect 27997 27013 28031 27047
rect 29745 27013 29779 27047
rect 36093 27013 36127 27047
rect 1869 26945 1903 26979
rect 7113 26945 7147 26979
rect 11529 26945 11563 26979
rect 20453 26945 20487 26979
rect 22385 26945 22419 26979
rect 24041 26945 24075 26979
rect 29837 26945 29871 26979
rect 34161 26945 34195 26979
rect 36921 26945 36955 26979
rect 38577 26945 38611 26979
rect 1593 26877 1627 26911
rect 3249 26877 3283 26911
rect 3709 26877 3743 26911
rect 4261 26877 4295 26911
rect 4721 26877 4755 26911
rect 5181 26877 5215 26911
rect 6009 26877 6043 26911
rect 6837 26877 6871 26911
rect 9413 26877 9447 26911
rect 10333 26877 10367 26911
rect 10425 26877 10459 26911
rect 11437 26877 11471 26911
rect 11897 26877 11931 26911
rect 12449 26877 12483 26911
rect 13553 26877 13587 26911
rect 13829 26877 13863 26911
rect 15669 26877 15703 26911
rect 16589 26877 16623 26911
rect 16865 26877 16899 26911
rect 17325 26877 17359 26911
rect 18061 26877 18095 26911
rect 18337 26877 18371 26911
rect 18521 26877 18555 26911
rect 18797 26877 18831 26911
rect 18990 26877 19024 26911
rect 19625 26877 19659 26911
rect 20085 26877 20119 26911
rect 20637 26877 20671 26911
rect 21925 26877 21959 26911
rect 22201 26877 22235 26911
rect 22845 26877 22879 26911
rect 23765 26877 23799 26911
rect 25881 26877 25915 26911
rect 26249 26877 26283 26911
rect 26893 26877 26927 26911
rect 28181 26877 28215 26911
rect 28549 26877 28583 26911
rect 28641 26877 28675 26911
rect 30665 26877 30699 26911
rect 30941 26877 30975 26911
rect 33149 26877 33183 26911
rect 33701 26877 33735 26911
rect 34989 26877 35023 26911
rect 35909 26877 35943 26911
rect 36645 26877 36679 26911
rect 38209 26877 38243 26911
rect 8493 26809 8527 26843
rect 15209 26809 15243 26843
rect 17509 26809 17543 26843
rect 25421 26809 25455 26843
rect 29469 26809 29503 26843
rect 30205 26809 30239 26843
rect 38025 26809 38059 26843
rect 10149 26741 10183 26775
rect 10609 26741 10643 26775
rect 12541 26741 12575 26775
rect 15853 26741 15887 26775
rect 23029 26741 23063 26775
rect 33241 26741 33275 26775
rect 5641 26537 5675 26571
rect 6377 26537 6411 26571
rect 18521 26537 18555 26571
rect 19257 26537 19291 26571
rect 21741 26537 21775 26571
rect 29745 26537 29779 26571
rect 31493 26537 31527 26571
rect 37841 26537 37875 26571
rect 38485 26537 38519 26571
rect 2053 26469 2087 26503
rect 33057 26469 33091 26503
rect 2605 26401 2639 26435
rect 2697 26401 2731 26435
rect 2881 26401 2915 26435
rect 3157 26401 3191 26435
rect 3341 26401 3375 26435
rect 4084 26401 4118 26435
rect 6193 26401 6227 26435
rect 7389 26401 7423 26435
rect 7757 26401 7791 26435
rect 8125 26401 8159 26435
rect 8585 26401 8619 26435
rect 12081 26401 12115 26435
rect 12265 26401 12299 26435
rect 12541 26401 12575 26435
rect 13093 26401 13127 26435
rect 13737 26401 13771 26435
rect 14289 26401 14323 26435
rect 15117 26401 15151 26435
rect 15301 26401 15335 26435
rect 16129 26401 16163 26435
rect 16313 26401 16347 26435
rect 17509 26401 17543 26435
rect 18061 26401 18095 26435
rect 18245 26401 18279 26435
rect 19165 26401 19199 26435
rect 19717 26401 19751 26435
rect 20913 26401 20947 26435
rect 21649 26401 21683 26435
rect 22385 26401 22419 26435
rect 22937 26401 22971 26435
rect 23857 26401 23891 26435
rect 24501 26401 24535 26435
rect 25145 26401 25179 26435
rect 25513 26401 25547 26435
rect 25789 26401 25823 26435
rect 26525 26401 26559 26435
rect 29653 26401 29687 26435
rect 30205 26401 30239 26435
rect 31401 26401 31435 26435
rect 32321 26401 32355 26435
rect 32873 26401 32907 26435
rect 33793 26401 33827 26435
rect 36001 26401 36035 26435
rect 36369 26401 36403 26435
rect 37013 26401 37047 26435
rect 37749 26401 37783 26435
rect 38577 26401 38611 26435
rect 38945 26401 38979 26435
rect 39957 26401 39991 26435
rect 4353 26333 4387 26367
rect 7205 26333 7239 26367
rect 9689 26333 9723 26367
rect 9965 26333 9999 26367
rect 11345 26333 11379 26367
rect 12817 26333 12851 26367
rect 14105 26333 14139 26367
rect 17325 26333 17359 26367
rect 23121 26333 23155 26367
rect 24593 26333 24627 26367
rect 27261 26333 27295 26367
rect 27537 26333 27571 26367
rect 30665 26333 30699 26367
rect 33517 26333 33551 26367
rect 35173 26333 35207 26367
rect 16405 26265 16439 26299
rect 22569 26265 22603 26299
rect 23949 26265 23983 26299
rect 26709 26265 26743 26299
rect 14933 26197 14967 26231
rect 21097 26197 21131 26231
rect 28641 26197 28675 26231
rect 36093 26197 36127 26231
rect 14473 25993 14507 26027
rect 16497 25993 16531 26027
rect 18337 25993 18371 26027
rect 23029 25993 23063 26027
rect 33333 25993 33367 26027
rect 36553 25993 36587 26027
rect 38669 25993 38703 26027
rect 3065 25925 3099 25959
rect 20913 25925 20947 25959
rect 25237 25925 25271 25959
rect 29929 25925 29963 25959
rect 2421 25857 2455 25891
rect 5457 25857 5491 25891
rect 8217 25857 8251 25891
rect 8953 25857 8987 25891
rect 15393 25857 15427 25891
rect 20269 25857 20303 25891
rect 31401 25857 31435 25891
rect 32229 25857 32263 25891
rect 35173 25857 35207 25891
rect 37289 25857 37323 25891
rect 1777 25789 1811 25823
rect 2283 25789 2317 25823
rect 3525 25789 3559 25823
rect 3985 25789 4019 25823
rect 4353 25789 4387 25823
rect 4721 25789 4755 25823
rect 5733 25789 5767 25823
rect 6193 25789 6227 25823
rect 7573 25789 7607 25823
rect 8125 25789 8159 25823
rect 9505 25789 9539 25823
rect 9781 25789 9815 25823
rect 9965 25789 9999 25823
rect 10885 25789 10919 25823
rect 11069 25789 11103 25823
rect 11345 25789 11379 25823
rect 11437 25789 11471 25823
rect 11805 25789 11839 25823
rect 13369 25789 13403 25823
rect 13645 25789 13679 25823
rect 13829 25789 13863 25823
rect 14289 25789 14323 25823
rect 15485 25789 15519 25823
rect 16037 25789 16071 25823
rect 16221 25789 16255 25823
rect 17141 25789 17175 25823
rect 18061 25789 18095 25823
rect 18205 25789 18239 25823
rect 19165 25789 19199 25823
rect 19717 25789 19751 25823
rect 19993 25789 20027 25823
rect 20729 25789 20763 25823
rect 22017 25789 22051 25823
rect 22293 25789 22327 25823
rect 22937 25789 22971 25823
rect 23673 25789 23707 25823
rect 24225 25789 24259 25823
rect 25421 25789 25455 25823
rect 25605 25789 25639 25823
rect 25789 25789 25823 25823
rect 26893 25789 26927 25823
rect 27077 25789 27111 25823
rect 27261 25789 27295 25823
rect 28181 25789 28215 25823
rect 28365 25789 28399 25823
rect 29653 25789 29687 25823
rect 30205 25789 30239 25823
rect 30573 25789 30607 25823
rect 31309 25789 31343 25823
rect 31953 25789 31987 25823
rect 34069 25789 34103 25823
rect 35449 25789 35483 25823
rect 37565 25789 37599 25823
rect 3433 25721 3467 25755
rect 5825 25721 5859 25755
rect 10425 25721 10459 25755
rect 12817 25721 12851 25755
rect 22477 25721 22511 25755
rect 26433 25721 26467 25755
rect 1593 25653 1627 25687
rect 5641 25653 5675 25687
rect 7481 25653 7515 25687
rect 17325 25653 17359 25687
rect 23949 25653 23983 25687
rect 27997 25653 28031 25687
rect 34253 25653 34287 25687
rect 5733 25449 5767 25483
rect 9045 25449 9079 25483
rect 9781 25449 9815 25483
rect 11529 25449 11563 25483
rect 35449 25449 35483 25483
rect 4077 25381 4111 25415
rect 11621 25381 11655 25415
rect 11713 25381 11747 25415
rect 12081 25381 12115 25415
rect 18337 25381 18371 25415
rect 20361 25381 20395 25415
rect 22017 25381 22051 25415
rect 28273 25381 28307 25415
rect 31493 25381 31527 25415
rect 1409 25313 1443 25347
rect 1685 25313 1719 25347
rect 4629 25313 4663 25347
rect 4905 25313 4939 25347
rect 5089 25313 5123 25347
rect 5549 25313 5583 25347
rect 6561 25313 6595 25347
rect 8861 25313 8895 25347
rect 9873 25313 9907 25347
rect 10241 25313 10275 25347
rect 10609 25313 10643 25347
rect 13277 25313 13311 25347
rect 13645 25313 13679 25347
rect 14013 25313 14047 25347
rect 15485 25313 15519 25347
rect 16221 25313 16255 25347
rect 17233 25313 17267 25347
rect 17785 25313 17819 25347
rect 17969 25313 18003 25347
rect 19165 25313 19199 25347
rect 19809 25313 19843 25347
rect 20177 25313 20211 25347
rect 20913 25313 20947 25347
rect 21281 25313 21315 25347
rect 21833 25313 21867 25347
rect 23029 25313 23063 25347
rect 23305 25313 23339 25347
rect 23765 25313 23799 25347
rect 24225 25313 24259 25347
rect 25053 25313 25087 25347
rect 25421 25313 25455 25347
rect 26617 25313 26651 25347
rect 29193 25313 29227 25347
rect 29561 25313 29595 25347
rect 30389 25313 30423 25347
rect 30573 25313 30607 25347
rect 30757 25313 30791 25347
rect 31401 25313 31435 25347
rect 32321 25313 32355 25347
rect 32689 25313 32723 25347
rect 34069 25313 34103 25347
rect 34529 25313 34563 25347
rect 35541 25313 35575 25347
rect 36093 25313 36127 25347
rect 36921 25313 36955 25347
rect 38209 25313 38243 25347
rect 38761 25313 38795 25347
rect 6837 25245 6871 25279
rect 8217 25245 8251 25279
rect 11345 25245 11379 25279
rect 13461 25245 13495 25279
rect 17049 25245 17083 25279
rect 25881 25245 25915 25279
rect 26893 25245 26927 25279
rect 28733 25245 28767 25279
rect 29653 25245 29687 25279
rect 32965 25245 32999 25279
rect 33793 25245 33827 25279
rect 36185 25245 36219 25279
rect 38853 25245 38887 25279
rect 23121 25177 23155 25211
rect 24961 25177 24995 25211
rect 32413 25177 32447 25211
rect 34529 25177 34563 25211
rect 38301 25177 38335 25211
rect 2789 25109 2823 25143
rect 15669 25109 15703 25143
rect 16405 25109 16439 25143
rect 24317 25109 24351 25143
rect 37105 25109 37139 25143
rect 19625 24905 19659 24939
rect 23857 24905 23891 24939
rect 2329 24837 2363 24871
rect 6009 24837 6043 24871
rect 20361 24837 20395 24871
rect 21097 24837 21131 24871
rect 22937 24837 22971 24871
rect 7757 24769 7791 24803
rect 11345 24769 11379 24803
rect 13185 24769 13219 24803
rect 15669 24769 15703 24803
rect 24501 24769 24535 24803
rect 24777 24769 24811 24803
rect 25881 24769 25915 24803
rect 27445 24769 27479 24803
rect 29561 24769 29595 24803
rect 30665 24769 30699 24803
rect 33057 24769 33091 24803
rect 35265 24769 35299 24803
rect 36737 24769 36771 24803
rect 2513 24701 2547 24735
rect 2973 24701 3007 24735
rect 3249 24701 3283 24735
rect 3709 24701 3743 24735
rect 4077 24701 4111 24735
rect 5365 24701 5399 24735
rect 5733 24701 5767 24735
rect 6101 24701 6135 24735
rect 7113 24701 7147 24735
rect 7665 24701 7699 24735
rect 8493 24701 8527 24735
rect 8769 24701 8803 24735
rect 10609 24701 10643 24735
rect 12725 24701 12759 24735
rect 14013 24701 14047 24735
rect 14289 24701 14323 24735
rect 16681 24701 16715 24735
rect 18613 24701 18647 24735
rect 19441 24701 19475 24735
rect 20177 24701 20211 24735
rect 20913 24701 20947 24735
rect 22017 24701 22051 24735
rect 22753 24701 22787 24735
rect 23673 24701 23707 24735
rect 26617 24701 26651 24735
rect 27721 24701 27755 24735
rect 28181 24701 28215 24735
rect 29101 24701 29135 24735
rect 29469 24701 29503 24735
rect 30941 24701 30975 24735
rect 31125 24701 31159 24735
rect 31953 24701 31987 24735
rect 32413 24701 32447 24735
rect 32781 24701 32815 24735
rect 34069 24701 34103 24735
rect 35173 24701 35207 24735
rect 35449 24701 35483 24735
rect 36185 24701 36219 24735
rect 36277 24701 36311 24735
rect 37197 24701 37231 24735
rect 37473 24701 37507 24735
rect 10149 24633 10183 24667
rect 10977 24633 11011 24667
rect 12449 24633 12483 24667
rect 12817 24633 12851 24667
rect 28457 24633 28491 24667
rect 30113 24633 30147 24667
rect 6929 24565 6963 24599
rect 10793 24565 10827 24599
rect 10885 24565 10919 24599
rect 12633 24565 12667 24599
rect 16865 24565 16899 24599
rect 18797 24565 18831 24599
rect 22201 24565 22235 24599
rect 26801 24565 26835 24599
rect 28917 24565 28951 24599
rect 34253 24565 34287 24599
rect 38577 24565 38611 24599
rect 1869 24361 1903 24395
rect 8953 24361 8987 24395
rect 9781 24361 9815 24395
rect 15393 24361 15427 24395
rect 21097 24361 21131 24395
rect 24317 24361 24351 24395
rect 27813 24361 27847 24395
rect 12357 24293 12391 24327
rect 15945 24293 15979 24327
rect 1777 24225 1811 24259
rect 2605 24225 2639 24259
rect 3341 24225 3375 24259
rect 4077 24225 4111 24259
rect 7113 24225 7147 24259
rect 8033 24225 8067 24259
rect 8861 24225 8895 24259
rect 9045 24225 9079 24259
rect 9965 24225 9999 24259
rect 10241 24225 10275 24259
rect 11161 24225 11195 24259
rect 11345 24225 11379 24259
rect 11897 24225 11931 24259
rect 12265 24225 12299 24259
rect 13461 24225 13495 24259
rect 13921 24225 13955 24259
rect 14565 24225 14599 24259
rect 15301 24225 15335 24259
rect 16221 24225 16255 24259
rect 16589 24225 16623 24259
rect 16957 24225 16991 24259
rect 17141 24225 17175 24259
rect 17785 24225 17819 24259
rect 18337 24225 18371 24259
rect 18613 24225 18647 24259
rect 18889 24225 18923 24259
rect 19073 24225 19107 24259
rect 19349 24225 19383 24259
rect 19809 24225 19843 24259
rect 20913 24225 20947 24259
rect 21741 24225 21775 24259
rect 22385 24225 22419 24259
rect 22753 24225 22787 24259
rect 23673 24225 23707 24259
rect 23857 24225 23891 24259
rect 24225 24225 24259 24259
rect 25421 24225 25455 24259
rect 25789 24225 25823 24259
rect 27077 24225 27111 24259
rect 27813 24225 27847 24259
rect 28365 24225 28399 24259
rect 28549 24225 28583 24259
rect 30113 24225 30147 24259
rect 32321 24225 32355 24259
rect 33149 24225 33183 24259
rect 33333 24225 33367 24259
rect 36369 24225 36403 24259
rect 36645 24225 36679 24259
rect 38025 24225 38059 24259
rect 38301 24225 38335 24259
rect 38945 24225 38979 24259
rect 2697 24157 2731 24191
rect 4997 24157 5031 24191
rect 5273 24157 5307 24191
rect 7205 24157 7239 24191
rect 13737 24157 13771 24191
rect 25881 24157 25915 24191
rect 27169 24157 27203 24191
rect 29837 24157 29871 24191
rect 33977 24157 34011 24191
rect 34253 24157 34287 24191
rect 35357 24157 35391 24191
rect 36461 24157 36495 24191
rect 39037 24157 39071 24191
rect 14657 24089 14691 24123
rect 25237 24089 25271 24123
rect 33149 24089 33183 24123
rect 37841 24089 37875 24123
rect 3433 24021 3467 24055
rect 4169 24021 4203 24055
rect 6561 24021 6595 24055
rect 21833 24021 21867 24055
rect 31401 24021 31435 24055
rect 7757 23817 7791 23851
rect 17417 23817 17451 23851
rect 19717 23817 19751 23851
rect 28641 23817 28675 23851
rect 32413 23817 32447 23851
rect 39037 23817 39071 23851
rect 2605 23749 2639 23783
rect 4261 23749 4295 23783
rect 5549 23749 5583 23783
rect 12541 23749 12575 23783
rect 15577 23749 15611 23783
rect 20361 23749 20395 23783
rect 22845 23749 22879 23783
rect 3341 23681 3375 23715
rect 9689 23681 9723 23715
rect 14013 23681 14047 23715
rect 14289 23681 14323 23715
rect 16865 23681 16899 23715
rect 18337 23681 18371 23715
rect 22201 23681 22235 23715
rect 23765 23681 23799 23715
rect 25881 23681 25915 23715
rect 30849 23681 30883 23715
rect 31401 23681 31435 23715
rect 31861 23681 31895 23715
rect 33057 23681 33091 23715
rect 35081 23681 35115 23715
rect 37473 23681 37507 23715
rect 2697 23613 2731 23647
rect 3249 23613 3283 23647
rect 4077 23613 4111 23647
rect 5733 23613 5767 23647
rect 6101 23613 6135 23647
rect 6193 23613 6227 23647
rect 7573 23613 7607 23647
rect 8953 23613 8987 23647
rect 9137 23613 9171 23647
rect 9597 23613 9631 23647
rect 11069 23613 11103 23647
rect 11621 23613 11655 23647
rect 11805 23613 11839 23647
rect 12633 23613 12667 23647
rect 13185 23613 13219 23647
rect 16129 23613 16163 23647
rect 16405 23613 16439 23647
rect 17325 23613 17359 23647
rect 18705 23613 18739 23647
rect 18889 23613 18923 23647
rect 19073 23613 19107 23647
rect 19349 23613 19383 23647
rect 20545 23613 20579 23647
rect 20821 23613 20855 23647
rect 21465 23613 21499 23647
rect 21925 23613 21959 23647
rect 22661 23613 22695 23647
rect 23857 23613 23891 23647
rect 24041 23613 24075 23647
rect 24409 23613 24443 23647
rect 25145 23613 25179 23647
rect 26249 23613 26283 23647
rect 26617 23613 26651 23647
rect 27261 23613 27295 23647
rect 27905 23613 27939 23647
rect 27997 23613 28031 23647
rect 28549 23613 28583 23647
rect 29561 23613 29595 23647
rect 30205 23613 30239 23647
rect 31677 23613 31711 23647
rect 32965 23613 32999 23647
rect 33333 23613 33367 23647
rect 33425 23613 33459 23647
rect 33977 23613 34011 23647
rect 35357 23613 35391 23647
rect 37749 23613 37783 23647
rect 16313 23545 16347 23579
rect 26801 23545 26835 23579
rect 29653 23545 29687 23579
rect 11069 23477 11103 23511
rect 30297 23477 30331 23511
rect 34161 23477 34195 23511
rect 36461 23477 36495 23511
rect 5181 23273 5215 23307
rect 8769 23273 8803 23307
rect 9781 23273 9815 23307
rect 17509 23273 17543 23307
rect 22385 23273 22419 23307
rect 24317 23273 24351 23307
rect 26617 23273 26651 23307
rect 28181 23273 28215 23307
rect 30849 23273 30883 23307
rect 32229 23273 32263 23307
rect 33701 23273 33735 23307
rect 35909 23273 35943 23307
rect 3157 23205 3191 23239
rect 19717 23205 19751 23239
rect 34161 23205 34195 23239
rect 1501 23137 1535 23171
rect 1777 23137 1811 23171
rect 4077 23137 4111 23171
rect 4905 23137 4939 23171
rect 5089 23137 5123 23171
rect 6009 23137 6043 23171
rect 6561 23137 6595 23171
rect 7205 23137 7239 23171
rect 7849 23137 7883 23171
rect 8585 23137 8619 23171
rect 9689 23137 9723 23171
rect 10333 23137 10367 23171
rect 10517 23137 10551 23171
rect 11529 23137 11563 23171
rect 12081 23137 12115 23171
rect 12357 23137 12391 23171
rect 13737 23137 13771 23171
rect 13921 23137 13955 23171
rect 14105 23137 14139 23171
rect 14289 23137 14323 23171
rect 14565 23137 14599 23171
rect 15393 23137 15427 23171
rect 16497 23137 16531 23171
rect 16681 23137 16715 23171
rect 16957 23137 16991 23171
rect 17141 23137 17175 23171
rect 18245 23137 18279 23171
rect 18613 23137 18647 23171
rect 18797 23137 18831 23171
rect 18981 23137 19015 23171
rect 19165 23137 19199 23171
rect 20177 23137 20211 23171
rect 21097 23137 21131 23171
rect 21557 23137 21591 23171
rect 22293 23137 22327 23171
rect 22937 23137 22971 23171
rect 25329 23137 25363 23171
rect 25605 23137 25639 23171
rect 25973 23137 26007 23171
rect 26801 23137 26835 23171
rect 27353 23137 27387 23171
rect 28089 23137 28123 23171
rect 28641 23137 28675 23171
rect 30205 23137 30239 23171
rect 30757 23137 30791 23171
rect 30941 23137 30975 23171
rect 31953 23137 31987 23171
rect 32137 23137 32171 23171
rect 32597 23137 32631 23171
rect 32965 23137 32999 23171
rect 33885 23137 33919 23171
rect 34805 23137 34839 23171
rect 35173 23137 35207 23171
rect 35357 23137 35391 23171
rect 35817 23137 35851 23171
rect 36461 23137 36495 23171
rect 38025 23137 38059 23171
rect 38301 23137 38335 23171
rect 38945 23137 38979 23171
rect 5825 23069 5859 23103
rect 6745 23069 6779 23103
rect 12449 23069 12483 23103
rect 13185 23069 13219 23103
rect 16129 23069 16163 23103
rect 21649 23069 21683 23103
rect 23213 23069 23247 23103
rect 27261 23069 27295 23103
rect 28917 23069 28951 23103
rect 34897 23069 34931 23103
rect 36645 23069 36679 23103
rect 8033 23001 8067 23035
rect 20269 23001 20303 23035
rect 37841 23001 37875 23035
rect 7297 22933 7331 22967
rect 15577 22933 15611 22967
rect 31769 22933 31803 22967
rect 39037 22933 39071 22967
rect 6929 22729 6963 22763
rect 11713 22729 11747 22763
rect 18245 22729 18279 22763
rect 18981 22729 19015 22763
rect 22753 22729 22787 22763
rect 25973 22729 26007 22763
rect 28917 22729 28951 22763
rect 31125 22729 31159 22763
rect 38393 22729 38427 22763
rect 4905 22661 4939 22695
rect 19901 22661 19935 22695
rect 33793 22661 33827 22695
rect 2973 22593 3007 22627
rect 6193 22593 6227 22627
rect 8033 22593 8067 22627
rect 9597 22593 9631 22627
rect 13829 22593 13863 22627
rect 17509 22593 17543 22627
rect 25329 22593 25363 22627
rect 32321 22593 32355 22627
rect 35909 22593 35943 22627
rect 37933 22593 37967 22627
rect 2145 22525 2179 22559
rect 2697 22525 2731 22559
rect 3525 22525 3559 22559
rect 4077 22525 4111 22559
rect 4537 22525 4571 22559
rect 4905 22525 4939 22559
rect 5549 22525 5583 22559
rect 6009 22525 6043 22559
rect 6837 22525 6871 22559
rect 7389 22525 7423 22559
rect 8309 22525 8343 22559
rect 10149 22525 10183 22559
rect 10425 22525 10459 22559
rect 12449 22525 12483 22559
rect 13001 22525 13035 22559
rect 14105 22525 14139 22559
rect 16037 22525 16071 22559
rect 16405 22525 16439 22559
rect 16589 22525 16623 22559
rect 16773 22525 16807 22559
rect 17049 22525 17083 22559
rect 18061 22525 18095 22559
rect 18797 22525 18831 22559
rect 19993 22525 20027 22559
rect 20361 22525 20395 22559
rect 20637 22525 20671 22559
rect 21373 22525 21407 22559
rect 21649 22525 21683 22559
rect 23673 22525 23707 22559
rect 24869 22525 24903 22559
rect 25237 22525 25271 22559
rect 26433 22525 26467 22559
rect 26617 22525 26651 22559
rect 26801 22525 26835 22559
rect 27077 22525 27111 22559
rect 27169 22525 27203 22559
rect 27997 22525 28031 22559
rect 29101 22525 29135 22559
rect 29561 22525 29595 22559
rect 29837 22525 29871 22559
rect 31677 22525 31711 22559
rect 32045 22525 32079 22559
rect 32413 22525 32447 22559
rect 32965 22525 32999 22559
rect 33609 22525 33643 22559
rect 34897 22525 34931 22559
rect 36185 22525 36219 22559
rect 37105 22525 37139 22559
rect 38117 22525 38151 22559
rect 38209 22525 38243 22559
rect 15485 22457 15519 22491
rect 24409 22457 24443 22491
rect 36093 22457 36127 22491
rect 36645 22457 36679 22491
rect 2053 22389 2087 22423
rect 12541 22389 12575 22423
rect 23857 22389 23891 22423
rect 28181 22389 28215 22423
rect 35081 22389 35115 22423
rect 37289 22389 37323 22423
rect 1593 22185 1627 22219
rect 4353 22185 4387 22219
rect 7389 22185 7423 22219
rect 8309 22185 8343 22219
rect 9781 22185 9815 22219
rect 11437 22185 11471 22219
rect 25329 22185 25363 22219
rect 26985 22185 27019 22219
rect 29837 22185 29871 22219
rect 33333 22185 33367 22219
rect 37841 22185 37875 22219
rect 14013 22117 14047 22151
rect 15393 22117 15427 22151
rect 1409 22049 1443 22083
rect 2329 22049 2363 22083
rect 2697 22049 2731 22083
rect 2973 22049 3007 22083
rect 4537 22049 4571 22083
rect 4813 22049 4847 22083
rect 5825 22049 5859 22083
rect 8033 22049 8067 22083
rect 8861 22049 8895 22083
rect 9045 22049 9079 22083
rect 9689 22049 9723 22083
rect 10609 22049 10643 22083
rect 10701 22049 10735 22083
rect 11253 22049 11287 22083
rect 12449 22049 12483 22083
rect 12725 22049 12759 22083
rect 13185 22049 13219 22083
rect 14197 22049 14231 22083
rect 14565 22049 14599 22083
rect 15301 22049 15335 22083
rect 16497 22049 16531 22083
rect 16681 22049 16715 22083
rect 16957 22049 16991 22083
rect 17049 22049 17083 22083
rect 18153 22049 18187 22083
rect 18797 22049 18831 22083
rect 19165 22049 19199 22083
rect 19625 22049 19659 22083
rect 20085 22049 20119 22083
rect 20913 22049 20947 22083
rect 22569 22049 22603 22083
rect 23673 22049 23707 22083
rect 24317 22049 24351 22083
rect 25513 22049 25547 22083
rect 25697 22049 25731 22083
rect 26985 22049 27019 22083
rect 27169 22049 27203 22083
rect 27721 22049 27755 22083
rect 28089 22049 28123 22083
rect 29101 22049 29135 22083
rect 29745 22049 29779 22083
rect 29929 22049 29963 22083
rect 30665 22049 30699 22083
rect 31033 22049 31067 22083
rect 31401 22049 31435 22083
rect 32321 22049 32355 22083
rect 33057 22049 33091 22083
rect 33885 22049 33919 22083
rect 36829 22049 36863 22083
rect 37749 22049 37783 22083
rect 38577 22049 38611 22083
rect 6101 21981 6135 22015
rect 13553 21981 13587 22015
rect 16129 21981 16163 22015
rect 17417 21981 17451 22015
rect 21189 21981 21223 22015
rect 24409 21981 24443 22015
rect 33793 21981 33827 22015
rect 35173 21981 35207 22015
rect 35449 21981 35483 22015
rect 38485 21981 38519 22015
rect 2973 21913 3007 21947
rect 20269 21913 20303 21947
rect 23857 21913 23891 21947
rect 31401 21913 31435 21947
rect 19349 21845 19383 21879
rect 32505 21845 32539 21879
rect 2973 21641 3007 21675
rect 18153 21641 18187 21675
rect 25237 21641 25271 21675
rect 38853 21641 38887 21675
rect 6101 21573 6135 21607
rect 6929 21573 6963 21607
rect 31493 21573 31527 21607
rect 33609 21573 33643 21607
rect 5365 21505 5399 21539
rect 7665 21505 7699 21539
rect 13737 21505 13771 21539
rect 14197 21505 14231 21539
rect 17049 21505 17083 21539
rect 23673 21505 23707 21539
rect 23949 21505 23983 21539
rect 29285 21505 29319 21539
rect 29561 21505 29595 21539
rect 32321 21505 32355 21539
rect 35449 21505 35483 21539
rect 37473 21505 37507 21539
rect 37749 21505 37783 21539
rect 1409 21437 1443 21471
rect 1685 21437 1719 21471
rect 4077 21437 4111 21471
rect 4353 21437 4387 21471
rect 4997 21437 5031 21471
rect 5273 21437 5307 21471
rect 5917 21437 5951 21471
rect 6837 21437 6871 21471
rect 7481 21437 7515 21471
rect 10701 21437 10735 21471
rect 11069 21437 11103 21471
rect 11437 21437 11471 21471
rect 12817 21437 12851 21471
rect 13185 21437 13219 21471
rect 13553 21437 13587 21471
rect 14473 21437 14507 21471
rect 16589 21437 16623 21471
rect 16773 21437 16807 21471
rect 18061 21437 18095 21471
rect 18889 21437 18923 21471
rect 19165 21437 19199 21471
rect 21465 21437 21499 21471
rect 21649 21437 21683 21471
rect 21833 21437 21867 21471
rect 22569 21437 22603 21471
rect 22753 21437 22787 21471
rect 22937 21437 22971 21471
rect 23213 21437 23247 21471
rect 26157 21437 26191 21471
rect 26801 21437 26835 21471
rect 26985 21437 27019 21471
rect 27721 21437 27755 21471
rect 28181 21437 28215 21471
rect 31401 21437 31435 21471
rect 31953 21437 31987 21471
rect 33241 21437 33275 21471
rect 33793 21437 33827 21471
rect 34161 21437 34195 21471
rect 34253 21437 34287 21471
rect 34897 21437 34931 21471
rect 35541 21437 35575 21471
rect 35817 21437 35851 21471
rect 36093 21437 36127 21471
rect 36829 21437 36863 21471
rect 11621 21369 11655 21403
rect 15853 21369 15887 21403
rect 21005 21369 21039 21403
rect 22109 21369 22143 21403
rect 20453 21301 20487 21335
rect 23305 21301 23339 21335
rect 26249 21301 26283 21335
rect 27813 21301 27847 21335
rect 30665 21301 30699 21335
rect 33057 21301 33091 21335
rect 1961 21097 1995 21131
rect 7205 21097 7239 21131
rect 15393 21097 15427 21131
rect 21189 21097 21223 21131
rect 23581 21097 23615 21131
rect 26985 21097 27019 21131
rect 29377 21097 29411 21131
rect 31493 21097 31527 21131
rect 32597 21097 32631 21131
rect 4813 21029 4847 21063
rect 10057 21029 10091 21063
rect 16221 21029 16255 21063
rect 18889 21029 18923 21063
rect 19809 21029 19843 21063
rect 19993 21029 20027 21063
rect 29285 21029 29319 21063
rect 29469 21029 29503 21063
rect 34805 21029 34839 21063
rect 1869 20961 1903 20995
rect 2973 20961 3007 20995
rect 3341 20961 3375 20995
rect 4905 20961 4939 20995
rect 8033 20961 8067 20995
rect 8769 20961 8803 20995
rect 9965 20961 9999 20995
rect 10425 20961 10459 20995
rect 10885 20961 10919 20995
rect 11161 20961 11195 20995
rect 11621 20961 11655 20995
rect 12725 20961 12759 20995
rect 12817 20961 12851 20995
rect 13461 20961 13495 20995
rect 13737 20961 13771 20995
rect 14381 20961 14415 20995
rect 15301 20961 15335 20995
rect 16681 20961 16715 20995
rect 16865 20961 16899 20995
rect 17141 20961 17175 20995
rect 17325 20961 17359 20995
rect 17601 20961 17635 20995
rect 18153 20961 18187 20995
rect 18613 20961 18647 20995
rect 19901 20961 19935 20995
rect 21097 20961 21131 20995
rect 21649 20961 21683 20995
rect 22569 20961 22603 20995
rect 23121 20961 23155 20995
rect 23489 20961 23523 20995
rect 23765 20961 23799 20995
rect 24133 20961 24167 20995
rect 24501 20961 24535 20995
rect 25421 20961 25455 20995
rect 25789 20961 25823 20995
rect 26801 20961 26835 20995
rect 27537 20961 27571 20995
rect 28089 20961 28123 20995
rect 29101 20961 29135 20995
rect 30573 20961 30607 20995
rect 31309 20961 31343 20995
rect 32413 20961 32447 20995
rect 33149 20961 33183 20995
rect 35817 20961 35851 20995
rect 37749 20961 37783 20995
rect 38117 20961 38151 20995
rect 38669 20961 38703 20995
rect 2513 20893 2547 20927
rect 3433 20893 3467 20927
rect 5825 20893 5859 20927
rect 6101 20893 6135 20927
rect 9045 20893 9079 20927
rect 19625 20893 19659 20927
rect 20361 20893 20395 20927
rect 21925 20893 21959 20927
rect 22477 20893 22511 20927
rect 25881 20893 25915 20927
rect 28365 20893 28399 20927
rect 29837 20893 29871 20927
rect 33425 20893 33459 20927
rect 35541 20893 35575 20927
rect 37841 20893 37875 20927
rect 8309 20825 8343 20859
rect 23305 20825 23339 20859
rect 25237 20825 25271 20859
rect 27813 20825 27847 20859
rect 4629 20757 4663 20791
rect 5089 20757 5123 20791
rect 12541 20757 12575 20791
rect 14565 20757 14599 20791
rect 22753 20757 22787 20791
rect 30757 20757 30791 20791
rect 36921 20757 36955 20791
rect 2973 20553 3007 20587
rect 3893 20553 3927 20587
rect 9505 20553 9539 20587
rect 16313 20553 16347 20587
rect 20729 20485 20763 20519
rect 23765 20485 23799 20519
rect 31401 20485 31435 20519
rect 4905 20417 4939 20451
rect 7941 20417 7975 20451
rect 10701 20417 10735 20451
rect 12449 20417 12483 20451
rect 14197 20417 14231 20451
rect 26709 20417 26743 20451
rect 30389 20417 30423 20451
rect 32137 20417 32171 20451
rect 36461 20417 36495 20451
rect 1409 20349 1443 20383
rect 1685 20349 1719 20383
rect 3801 20349 3835 20383
rect 4629 20349 4663 20383
rect 8217 20349 8251 20383
rect 10333 20349 10367 20383
rect 10609 20349 10643 20383
rect 10885 20349 10919 20383
rect 11713 20349 11747 20383
rect 12909 20349 12943 20383
rect 13093 20349 13127 20383
rect 13277 20349 13311 20383
rect 13921 20349 13955 20383
rect 16037 20349 16071 20383
rect 16129 20349 16163 20383
rect 17233 20349 17267 20383
rect 23673 20349 23707 20383
rect 24133 20349 24167 20383
rect 24409 20349 24443 20383
rect 24869 20349 24903 20383
rect 25605 20349 25639 20383
rect 26433 20349 26467 20383
rect 28549 20349 28583 20383
rect 29561 20349 29595 20383
rect 30481 20349 30515 20383
rect 30941 20349 30975 20383
rect 31033 20349 31067 20383
rect 32597 20349 32631 20383
rect 32781 20349 32815 20383
rect 32965 20349 32999 20383
rect 33609 20349 33643 20383
rect 34161 20349 34195 20383
rect 35173 20349 35207 20383
rect 35449 20349 35483 20383
rect 36737 20349 36771 20383
rect 38577 20349 38611 20383
rect 3617 20281 3651 20315
rect 19441 20281 19475 20315
rect 21649 20281 21683 20315
rect 23397 20281 23431 20315
rect 6009 20213 6043 20247
rect 11805 20213 11839 20247
rect 15301 20213 15335 20247
rect 17417 20213 17451 20247
rect 27813 20213 27847 20247
rect 28641 20213 28675 20247
rect 29745 20213 29779 20247
rect 33701 20213 33735 20247
rect 34989 20213 35023 20247
rect 37841 20213 37875 20247
rect 38669 20213 38703 20247
rect 10149 20009 10183 20043
rect 20361 20009 20395 20043
rect 25881 20009 25915 20043
rect 35633 20009 35667 20043
rect 8125 19941 8159 19975
rect 13185 19941 13219 19975
rect 16129 19941 16163 19975
rect 32689 19941 32723 19975
rect 37749 19941 37783 19975
rect 2605 19873 2639 19907
rect 2881 19873 2915 19907
rect 3341 19873 3375 19907
rect 4077 19873 4111 19907
rect 4813 19873 4847 19907
rect 4997 19873 5031 19907
rect 5733 19873 5767 19907
rect 8677 19873 8711 19907
rect 8953 19873 8987 19907
rect 9965 19873 9999 19907
rect 10701 19873 10735 19907
rect 11805 19873 11839 19907
rect 14197 19873 14231 19907
rect 15301 19873 15335 19907
rect 16589 19873 16623 19907
rect 16865 19873 16899 19907
rect 16957 19873 16991 19907
rect 17141 19873 17175 19907
rect 17509 19873 17543 19907
rect 17693 19873 17727 19907
rect 18613 19873 18647 19907
rect 18705 19873 18739 19907
rect 18889 19873 18923 19907
rect 19165 19873 19199 19907
rect 19349 19873 19383 19907
rect 20177 19873 20211 19907
rect 20913 19873 20947 19907
rect 22569 19873 22603 19907
rect 22937 19873 22971 19907
rect 23029 19873 23063 19907
rect 24225 19873 24259 19907
rect 24593 19873 24627 19907
rect 25789 19873 25823 19907
rect 27077 19873 27111 19907
rect 27629 19873 27663 19907
rect 27905 19873 27939 19907
rect 29653 19873 29687 19907
rect 29929 19873 29963 19907
rect 30665 19873 30699 19907
rect 31217 19873 31251 19907
rect 32229 19873 32263 19907
rect 33333 19873 33367 19907
rect 33885 19873 33919 19907
rect 33977 19873 34011 19907
rect 34437 19873 34471 19907
rect 35173 19873 35207 19907
rect 35633 19873 35667 19907
rect 35725 19873 35759 19907
rect 36277 19873 36311 19907
rect 36645 19873 36679 19907
rect 36921 19873 36955 19907
rect 38393 19873 38427 19907
rect 38485 19873 38519 19907
rect 38761 19873 38795 19907
rect 3525 19805 3559 19839
rect 6009 19805 6043 19839
rect 9137 19805 9171 19839
rect 11529 19805 11563 19839
rect 14105 19805 14139 19839
rect 18061 19805 18095 19839
rect 21925 19805 21959 19839
rect 22385 19805 22419 19839
rect 24685 19805 24719 19839
rect 27997 19805 28031 19839
rect 29285 19805 29319 19839
rect 31033 19805 31067 19839
rect 32137 19805 32171 19839
rect 33425 19805 33459 19839
rect 36185 19805 36219 19839
rect 38853 19805 38887 19839
rect 4353 19737 4387 19771
rect 15485 19737 15519 19771
rect 24041 19737 24075 19771
rect 29929 19737 29963 19771
rect 7113 19669 7147 19703
rect 10885 19669 10919 19703
rect 14381 19669 14415 19703
rect 17877 19669 17911 19703
rect 21097 19669 21131 19703
rect 2053 19465 2087 19499
rect 4353 19465 4387 19499
rect 9873 19465 9907 19499
rect 14013 19465 14047 19499
rect 31309 19465 31343 19499
rect 34253 19465 34287 19499
rect 35081 19465 35115 19499
rect 25881 19329 25915 19363
rect 30205 19329 30239 19363
rect 1685 19261 1719 19295
rect 1777 19261 1811 19295
rect 1910 19261 1944 19295
rect 2789 19261 2823 19295
rect 3065 19261 3099 19295
rect 5917 19261 5951 19295
rect 7113 19261 7147 19295
rect 7297 19261 7331 19295
rect 8401 19261 8435 19295
rect 9689 19261 9723 19295
rect 10425 19261 10459 19295
rect 10517 19261 10551 19295
rect 10609 19261 10643 19295
rect 11529 19261 11563 19295
rect 12449 19261 12483 19295
rect 12725 19261 12759 19295
rect 15025 19261 15059 19295
rect 15117 19261 15151 19295
rect 15577 19261 15611 19295
rect 16497 19261 16531 19295
rect 16773 19261 16807 19295
rect 16957 19261 16991 19295
rect 17141 19261 17175 19295
rect 17417 19261 17451 19295
rect 18061 19261 18095 19295
rect 18613 19261 18647 19295
rect 19441 19261 19475 19295
rect 19625 19261 19659 19295
rect 19717 19261 19751 19295
rect 19993 19261 20027 19295
rect 20269 19261 20303 19295
rect 20637 19261 20671 19295
rect 21189 19261 21223 19295
rect 21465 19261 21499 19295
rect 21833 19261 21867 19295
rect 22293 19261 22327 19295
rect 22477 19261 22511 19295
rect 22845 19261 22879 19295
rect 22937 19261 22971 19295
rect 23673 19261 23707 19295
rect 24225 19261 24259 19295
rect 24685 19261 24719 19295
rect 26065 19261 26099 19295
rect 26525 19261 26559 19295
rect 26617 19261 26651 19295
rect 27261 19261 27295 19295
rect 28273 19261 28307 19295
rect 28457 19261 28491 19295
rect 29469 19261 29503 19295
rect 29653 19261 29687 19295
rect 30113 19261 30147 19295
rect 31401 19261 31435 19295
rect 31585 19261 31619 19295
rect 32229 19261 32263 19295
rect 33149 19261 33183 19295
rect 33333 19261 33367 19295
rect 33701 19261 33735 19295
rect 34161 19261 34195 19295
rect 34897 19261 34931 19295
rect 35633 19261 35667 19295
rect 36369 19261 36403 19295
rect 36737 19261 36771 19295
rect 37473 19261 37507 19295
rect 37749 19261 37783 19295
rect 11069 19193 11103 19227
rect 16037 19193 16071 19227
rect 18889 19193 18923 19227
rect 28733 19193 28767 19227
rect 37013 19193 37047 19227
rect 6101 19125 6135 19159
rect 6929 19125 6963 19159
rect 8585 19125 8619 19159
rect 10425 19125 10459 19159
rect 11713 19125 11747 19159
rect 18153 19125 18187 19159
rect 20545 19125 20579 19159
rect 23765 19125 23799 19159
rect 35725 19125 35759 19159
rect 38853 19125 38887 19159
rect 2789 18921 2823 18955
rect 4169 18921 4203 18955
rect 9045 18921 9079 18955
rect 19809 18921 19843 18955
rect 19901 18921 19935 18955
rect 21005 18921 21039 18955
rect 37841 18921 37875 18955
rect 19625 18853 19659 18887
rect 19993 18853 20027 18887
rect 30757 18853 30791 18887
rect 32873 18853 32907 18887
rect 34437 18853 34471 18887
rect 39037 18853 39071 18887
rect 1409 18785 1443 18819
rect 4077 18785 4111 18819
rect 5181 18785 5215 18819
rect 6285 18785 6319 18819
rect 6837 18785 6871 18819
rect 7113 18785 7147 18819
rect 8953 18785 8987 18819
rect 9689 18785 9723 18819
rect 14565 18785 14599 18819
rect 15577 18785 15611 18819
rect 17693 18785 17727 18819
rect 18429 18785 18463 18819
rect 18705 18785 18739 18819
rect 19073 18785 19107 18819
rect 19257 18785 19291 18819
rect 21097 18785 21131 18819
rect 21465 18785 21499 18819
rect 21925 18785 21959 18819
rect 22477 18785 22511 18819
rect 23673 18785 23707 18819
rect 24041 18785 24075 18819
rect 25053 18785 25087 18819
rect 25697 18785 25731 18819
rect 26801 18785 26835 18819
rect 27169 18785 27203 18819
rect 27445 18785 27479 18819
rect 27721 18785 27755 18819
rect 28457 18785 28491 18819
rect 29377 18785 29411 18819
rect 31217 18785 31251 18819
rect 32137 18785 32171 18819
rect 32597 18785 32631 18819
rect 33609 18785 33643 18819
rect 33977 18785 34011 18819
rect 34253 18785 34287 18819
rect 35265 18785 35299 18819
rect 35449 18785 35483 18819
rect 35725 18785 35759 18819
rect 36461 18785 36495 18819
rect 36921 18785 36955 18819
rect 37749 18785 37783 18819
rect 38301 18785 38335 18819
rect 38945 18785 38979 18819
rect 1685 18717 1719 18751
rect 5089 18717 5123 18751
rect 10333 18717 10367 18751
rect 10609 18717 10643 18751
rect 12449 18717 12483 18751
rect 12725 18717 12759 18751
rect 15301 18717 15335 18751
rect 20361 18717 20395 18751
rect 24501 18717 24535 18751
rect 26893 18717 26927 18751
rect 29101 18717 29135 18751
rect 6101 18649 6135 18683
rect 14657 18649 14691 18683
rect 16865 18649 16899 18683
rect 19073 18649 19107 18683
rect 23765 18649 23799 18683
rect 31401 18649 31435 18683
rect 33425 18649 33459 18683
rect 5365 18581 5399 18615
rect 8217 18581 8251 18615
rect 9781 18581 9815 18615
rect 11897 18581 11931 18615
rect 13829 18581 13863 18615
rect 19441 18581 19475 18615
rect 22661 18581 22695 18615
rect 25145 18581 25179 18615
rect 25881 18581 25915 18615
rect 28549 18581 28583 18615
rect 36369 18581 36403 18615
rect 37105 18581 37139 18615
rect 5917 18377 5951 18411
rect 11253 18377 11287 18411
rect 28641 18377 28675 18411
rect 37013 18377 37047 18411
rect 16221 18309 16255 18343
rect 16773 18309 16807 18343
rect 21557 18309 21591 18343
rect 32321 18309 32355 18343
rect 32689 18309 32723 18343
rect 2973 18241 3007 18275
rect 3525 18241 3559 18275
rect 9873 18241 9907 18275
rect 14105 18241 14139 18275
rect 19625 18241 19659 18275
rect 22293 18241 22327 18275
rect 26893 18241 26927 18275
rect 31493 18241 31527 18275
rect 33425 18241 33459 18275
rect 36093 18241 36127 18275
rect 37381 18241 37415 18275
rect 3801 18173 3835 18207
rect 3985 18173 4019 18207
rect 4445 18173 4479 18207
rect 4537 18173 4571 18207
rect 4813 18173 4847 18207
rect 7113 18173 7147 18207
rect 7757 18173 7791 18207
rect 8033 18173 8067 18207
rect 10149 18173 10183 18207
rect 12449 18173 12483 18207
rect 12541 18173 12575 18207
rect 13829 18173 13863 18207
rect 16037 18173 16071 18207
rect 16957 18173 16991 18207
rect 17049 18173 17083 18207
rect 18613 18173 18647 18207
rect 19349 18173 19383 18207
rect 21465 18173 21499 18207
rect 22201 18173 22235 18207
rect 24133 18173 24167 18207
rect 24409 18173 24443 18207
rect 24593 18173 24627 18207
rect 24869 18173 24903 18207
rect 25122 18173 25156 18207
rect 26709 18173 26743 18207
rect 27169 18173 27203 18207
rect 27261 18173 27295 18207
rect 27721 18173 27755 18207
rect 28457 18173 28491 18207
rect 29469 18173 29503 18207
rect 29653 18173 29687 18207
rect 29837 18173 29871 18207
rect 30849 18173 30883 18207
rect 31217 18173 31251 18207
rect 32505 18173 32539 18207
rect 32597 18173 32631 18207
rect 33241 18173 33275 18207
rect 34161 18173 34195 18207
rect 35265 18173 35299 18207
rect 35449 18173 35483 18207
rect 35909 18173 35943 18207
rect 36461 18173 36495 18207
rect 37197 18173 37231 18207
rect 37657 18173 37691 18207
rect 13001 18105 13035 18139
rect 17509 18105 17543 18139
rect 25697 18105 25731 18139
rect 34253 18105 34287 18139
rect 4445 18037 4479 18071
rect 7205 18037 7239 18071
rect 9321 18037 9355 18071
rect 15209 18037 15243 18071
rect 18797 18037 18831 18071
rect 20729 18037 20763 18071
rect 30757 18037 30791 18071
rect 38761 18037 38795 18071
rect 25881 17833 25915 17867
rect 33701 17833 33735 17867
rect 36921 17833 36955 17867
rect 37841 17833 37875 17867
rect 39037 17833 39071 17867
rect 3065 17765 3099 17799
rect 7757 17765 7791 17799
rect 10241 17765 10275 17799
rect 14749 17765 14783 17799
rect 15669 17765 15703 17799
rect 26525 17765 26559 17799
rect 1409 17697 1443 17731
rect 5181 17697 5215 17731
rect 5365 17697 5399 17731
rect 8401 17697 8435 17731
rect 9781 17697 9815 17731
rect 11437 17697 11471 17731
rect 11805 17697 11839 17731
rect 11989 17697 12023 17731
rect 12633 17697 12667 17731
rect 13185 17697 13219 17731
rect 14289 17697 14323 17731
rect 1685 17629 1719 17663
rect 5457 17629 5491 17663
rect 6101 17629 6135 17663
rect 6377 17629 6411 17663
rect 9689 17629 9723 17663
rect 12265 17629 12299 17663
rect 14197 17629 14231 17663
rect 8585 17561 8619 17595
rect 15853 17697 15887 17731
rect 17325 17697 17359 17731
rect 17601 17697 17635 17731
rect 18153 17697 18187 17731
rect 18521 17697 18555 17731
rect 19073 17697 19107 17731
rect 19809 17697 19843 17731
rect 20085 17697 20119 17731
rect 23857 17697 23891 17731
rect 25697 17697 25731 17731
rect 26985 17697 27019 17731
rect 27353 17697 27387 17731
rect 27445 17697 27479 17731
rect 28549 17697 28583 17731
rect 28733 17697 28767 17731
rect 29377 17697 29411 17731
rect 29561 17697 29595 17731
rect 29929 17697 29963 17731
rect 30849 17697 30883 17731
rect 31401 17697 31435 17731
rect 32321 17697 32355 17731
rect 32597 17697 32631 17731
rect 35265 17697 35299 17731
rect 35449 17697 35483 17731
rect 36001 17697 36035 17731
rect 36737 17697 36771 17731
rect 37749 17697 37783 17731
rect 38301 17697 38335 17731
rect 38945 17697 38979 17731
rect 15761 17629 15795 17663
rect 21465 17629 21499 17663
rect 21741 17629 21775 17663
rect 23581 17629 23615 17663
rect 28641 17629 28675 17663
rect 31217 17629 31251 17663
rect 34437 17629 34471 17663
rect 34989 17629 35023 17663
rect 17233 17561 17267 17595
rect 19625 17561 19659 17595
rect 36185 17561 36219 17595
rect 15669 17493 15703 17527
rect 16037 17493 16071 17527
rect 23029 17493 23063 17527
rect 24961 17493 24995 17527
rect 2789 17289 2823 17323
rect 5917 17289 5951 17323
rect 8861 17289 8895 17323
rect 16129 17289 16163 17323
rect 26433 17289 26467 17323
rect 33057 17289 33091 17323
rect 34989 17289 35023 17323
rect 9781 17221 9815 17255
rect 17417 17221 17451 17255
rect 19533 17221 19567 17255
rect 38853 17221 38887 17255
rect 1409 17153 1443 17187
rect 1685 17153 1719 17187
rect 5641 17153 5675 17187
rect 7297 17153 7331 17187
rect 12449 17153 12483 17187
rect 12725 17153 12759 17187
rect 14749 17153 14783 17187
rect 18521 17153 18555 17187
rect 26157 17153 26191 17187
rect 27445 17153 27479 17187
rect 3525 17085 3559 17119
rect 3801 17085 3835 17119
rect 5733 17085 5767 17119
rect 7573 17085 7607 17119
rect 9597 17085 9631 17119
rect 10701 17085 10735 17119
rect 10977 17085 11011 17119
rect 11621 17085 11655 17119
rect 15025 17085 15059 17119
rect 17325 17085 17359 17119
rect 18337 17085 18371 17119
rect 18613 17085 18647 17119
rect 19441 17085 19475 17119
rect 19901 17085 19935 17119
rect 20177 17085 20211 17119
rect 20729 17085 20763 17119
rect 21281 17085 21315 17119
rect 22017 17085 22051 17119
rect 22845 17085 22879 17119
rect 24041 17085 24075 17119
rect 24317 17085 24351 17119
rect 26249 17085 26283 17119
rect 27629 17085 27663 17119
rect 27721 17085 27755 17119
rect 29469 17085 29503 17119
rect 30205 17085 30239 17119
rect 30665 17085 30699 17119
rect 31309 17085 31343 17119
rect 31401 17085 31435 17119
rect 31769 17085 31803 17119
rect 32965 17085 32999 17119
rect 33793 17085 33827 17119
rect 34161 17085 34195 17119
rect 34897 17085 34931 17119
rect 35541 17085 35575 17119
rect 36185 17085 36219 17119
rect 36553 17085 36587 17119
rect 36921 17085 36955 17119
rect 37473 17085 37507 17119
rect 37749 17085 37783 17119
rect 5181 17017 5215 17051
rect 25697 17017 25731 17051
rect 27813 17017 27847 17051
rect 28181 17017 28215 17051
rect 30481 17017 30515 17051
rect 34345 17017 34379 17051
rect 10517 16949 10551 16983
rect 11805 16949 11839 16983
rect 13829 16949 13863 16983
rect 22201 16949 22235 16983
rect 23029 16949 23063 16983
rect 29561 16949 29595 16983
rect 36737 16949 36771 16983
rect 1961 16745 1995 16779
rect 2513 16745 2547 16779
rect 5273 16745 5307 16779
rect 6377 16745 6411 16779
rect 11529 16745 11563 16779
rect 14657 16745 14691 16779
rect 15485 16745 15519 16779
rect 16221 16745 16255 16779
rect 20269 16745 20303 16779
rect 31217 16745 31251 16779
rect 32321 16745 32355 16779
rect 33149 16745 33183 16779
rect 36001 16745 36035 16779
rect 38117 16745 38151 16779
rect 7389 16677 7423 16711
rect 38209 16677 38243 16711
rect 38577 16677 38611 16711
rect 1777 16609 1811 16643
rect 2697 16609 2731 16643
rect 4169 16609 4203 16643
rect 5365 16609 5399 16643
rect 5733 16609 5767 16643
rect 6561 16609 6595 16643
rect 6837 16609 6871 16643
rect 7205 16609 7239 16643
rect 8217 16609 8251 16643
rect 8401 16609 8435 16643
rect 8953 16609 8987 16643
rect 9965 16609 9999 16643
rect 10057 16609 10091 16643
rect 10425 16609 10459 16643
rect 11345 16609 11379 16643
rect 12449 16609 12483 16643
rect 12725 16609 12759 16643
rect 14565 16609 14599 16643
rect 15301 16609 15335 16643
rect 16037 16609 16071 16643
rect 17049 16609 17083 16643
rect 19165 16609 19199 16643
rect 20177 16609 20211 16643
rect 21005 16609 21039 16643
rect 21649 16609 21683 16643
rect 21925 16609 21959 16643
rect 22385 16609 22419 16643
rect 22661 16609 22695 16643
rect 23397 16609 23431 16643
rect 24317 16609 24351 16643
rect 25697 16609 25731 16643
rect 26801 16609 26835 16643
rect 27169 16609 27203 16643
rect 27445 16609 27479 16643
rect 27813 16609 27847 16643
rect 28273 16609 28307 16643
rect 29193 16609 29227 16643
rect 31033 16609 31067 16643
rect 32137 16609 32171 16643
rect 32965 16609 32999 16643
rect 33701 16609 33735 16643
rect 33977 16609 34011 16643
rect 35817 16609 35851 16643
rect 36645 16609 36679 16643
rect 36829 16609 36863 16643
rect 38025 16609 38059 16643
rect 4077 16541 4111 16575
rect 9137 16541 9171 16575
rect 9781 16541 9815 16575
rect 16773 16541 16807 16575
rect 21833 16541 21867 16575
rect 24041 16541 24075 16575
rect 26893 16541 26927 16575
rect 28917 16541 28951 16575
rect 37197 16541 37231 16575
rect 37841 16541 37875 16575
rect 4353 16405 4387 16439
rect 14013 16405 14047 16439
rect 18153 16405 18187 16439
rect 19349 16405 19383 16439
rect 23489 16405 23523 16439
rect 30297 16405 30331 16439
rect 35081 16405 35115 16439
rect 4537 16201 4571 16235
rect 10977 16201 11011 16235
rect 16865 16201 16899 16235
rect 34989 16201 35023 16235
rect 38853 16201 38887 16235
rect 7113 16133 7147 16167
rect 11713 16133 11747 16167
rect 14013 16133 14047 16167
rect 18153 16133 18187 16167
rect 2973 16065 3007 16099
rect 3249 16065 3283 16099
rect 5733 16065 5767 16099
rect 9689 16065 9723 16099
rect 19993 16065 20027 16099
rect 23121 16065 23155 16099
rect 24317 16065 24351 16099
rect 26341 16065 26375 16099
rect 27813 16065 27847 16099
rect 30573 16065 30607 16099
rect 37565 16065 37599 16099
rect 5365 15997 5399 16031
rect 5641 15997 5675 16031
rect 6837 15997 6871 16031
rect 7389 15997 7423 16031
rect 7573 15997 7607 16031
rect 8217 15997 8251 16031
rect 8769 15997 8803 16031
rect 9413 15997 9447 16031
rect 11529 15997 11563 16031
rect 12817 15997 12851 16031
rect 13277 15997 13311 16031
rect 13461 15997 13495 16031
rect 14105 15997 14139 16031
rect 14565 15997 14599 16031
rect 14933 15997 14967 16031
rect 15301 15997 15335 16031
rect 15853 15997 15887 16031
rect 16681 15997 16715 16031
rect 18061 15997 18095 16031
rect 18705 15997 18739 16031
rect 19625 15997 19659 16031
rect 20085 15997 20119 16031
rect 20269 15997 20303 16031
rect 20729 15997 20763 16031
rect 21097 15997 21131 16031
rect 22661 15997 22695 16031
rect 22845 15997 22879 16031
rect 23673 15997 23707 16031
rect 24225 15997 24259 16031
rect 26617 15997 26651 16031
rect 26801 15997 26835 16031
rect 28089 15997 28123 16031
rect 28273 15997 28307 16031
rect 30297 15997 30331 16031
rect 32413 15997 32447 16031
rect 33333 15997 33367 16031
rect 33517 15997 33551 16031
rect 34161 15997 34195 16031
rect 34345 15997 34379 16031
rect 34897 15997 34931 16031
rect 35633 15997 35667 16031
rect 36001 15997 36035 16031
rect 36185 15997 36219 16031
rect 36553 15997 36587 16031
rect 37289 15997 37323 16031
rect 25789 15929 25823 15963
rect 27261 15929 27295 15963
rect 18797 15861 18831 15895
rect 31677 15861 31711 15895
rect 32505 15861 32539 15895
rect 7573 15657 7607 15691
rect 14289 15657 14323 15691
rect 16037 15657 16071 15691
rect 33977 15657 34011 15691
rect 36921 15657 36955 15691
rect 18429 15589 18463 15623
rect 27077 15589 27111 15623
rect 1409 15521 1443 15555
rect 1685 15521 1719 15555
rect 4077 15521 4111 15555
rect 5733 15521 5767 15555
rect 6469 15521 6503 15555
rect 8309 15521 8343 15555
rect 10149 15521 10183 15555
rect 10885 15521 10919 15555
rect 11437 15521 11471 15555
rect 11805 15521 11839 15555
rect 12081 15521 12115 15555
rect 12725 15521 12759 15555
rect 13277 15521 13311 15555
rect 13921 15521 13955 15555
rect 14013 15521 14047 15555
rect 14565 15521 14599 15555
rect 15301 15521 15335 15555
rect 15945 15521 15979 15555
rect 16773 15521 16807 15555
rect 19073 15521 19107 15555
rect 19625 15521 19659 15555
rect 19809 15521 19843 15555
rect 21281 15521 21315 15555
rect 21925 15521 21959 15555
rect 22293 15521 22327 15555
rect 22477 15521 22511 15555
rect 22937 15521 22971 15555
rect 23673 15521 23707 15555
rect 24133 15521 24167 15555
rect 26617 15521 26651 15555
rect 28457 15521 28491 15555
rect 28825 15521 28859 15555
rect 30021 15521 30055 15555
rect 30481 15521 30515 15555
rect 31217 15521 31251 15555
rect 31315 15521 31349 15555
rect 32137 15521 32171 15555
rect 32781 15521 32815 15555
rect 33885 15521 33919 15555
rect 34529 15521 34563 15555
rect 34713 15521 34747 15555
rect 35081 15521 35115 15555
rect 35817 15521 35851 15555
rect 37933 15521 37967 15555
rect 38485 15521 38519 15555
rect 4353 15453 4387 15487
rect 6193 15453 6227 15487
rect 10517 15453 10551 15487
rect 15393 15453 15427 15487
rect 17049 15453 17083 15487
rect 18889 15453 18923 15487
rect 22201 15453 22235 15487
rect 24409 15453 24443 15487
rect 26525 15453 26559 15487
rect 28089 15453 28123 15487
rect 29745 15453 29779 15487
rect 32965 15453 32999 15487
rect 35541 15453 35575 15487
rect 38393 15453 38427 15487
rect 11621 15385 11655 15419
rect 19993 15385 20027 15419
rect 28733 15385 28767 15419
rect 30481 15385 30515 15419
rect 31217 15385 31251 15419
rect 32413 15385 32447 15419
rect 2789 15317 2823 15351
rect 8493 15317 8527 15351
rect 13737 15317 13771 15351
rect 31493 15317 31527 15351
rect 38669 15317 38703 15351
rect 5181 15113 5215 15147
rect 8401 15113 8435 15147
rect 11897 15113 11931 15147
rect 21833 15113 21867 15147
rect 31493 15113 31527 15147
rect 34069 15113 34103 15147
rect 38853 15113 38887 15147
rect 3341 14977 3375 15011
rect 4077 14977 4111 15011
rect 7113 14977 7147 15011
rect 9137 14977 9171 15011
rect 13461 14977 13495 15011
rect 14289 14977 14323 15011
rect 16589 14977 16623 15011
rect 19441 14977 19475 15011
rect 24409 14977 24443 15011
rect 26249 14977 26283 15011
rect 26525 14977 26559 15011
rect 29469 14977 29503 15011
rect 30481 14977 30515 15011
rect 33057 14977 33091 15011
rect 37473 14977 37507 15011
rect 1685 14909 1719 14943
rect 1961 14909 1995 14943
rect 3801 14909 3835 14943
rect 6009 14909 6043 14943
rect 6837 14909 6871 14943
rect 9321 14909 9355 14943
rect 9781 14909 9815 14943
rect 10701 14909 10735 14943
rect 11069 14909 11103 14943
rect 11345 14909 11379 14943
rect 12081 14909 12115 14943
rect 12449 14909 12483 14943
rect 13369 14909 13403 14943
rect 13737 14909 13771 14943
rect 14565 14909 14599 14943
rect 16957 14909 16991 14943
rect 17233 14909 17267 14943
rect 18245 14909 18279 14943
rect 18705 14909 18739 14943
rect 19349 14909 19383 14943
rect 19809 14909 19843 14943
rect 20361 14909 20395 14943
rect 20729 14909 20763 14943
rect 21005 14909 21039 14943
rect 21741 14909 21775 14943
rect 22937 14909 22971 14943
rect 24133 14909 24167 14943
rect 30021 14909 30055 14943
rect 30297 14909 30331 14943
rect 31309 14909 31343 14943
rect 32321 14909 32355 14943
rect 32413 14909 32447 14943
rect 32781 14909 32815 14943
rect 33517 14909 33551 14943
rect 33977 14909 34011 14943
rect 35909 14909 35943 14943
rect 36093 14909 36127 14943
rect 36277 14909 36311 14943
rect 37749 14909 37783 14943
rect 10057 14841 10091 14875
rect 17509 14841 17543 14875
rect 27905 14841 27939 14875
rect 35449 14841 35483 14875
rect 6193 14773 6227 14807
rect 12541 14773 12575 14807
rect 15853 14773 15887 14807
rect 18245 14773 18279 14807
rect 23029 14773 23063 14807
rect 25697 14773 25731 14807
rect 2789 14569 2823 14603
rect 13553 14569 13587 14603
rect 16497 14569 16531 14603
rect 17969 14569 18003 14603
rect 23305 14569 23339 14603
rect 34989 14569 35023 14603
rect 37841 14569 37875 14603
rect 17233 14501 17267 14535
rect 1685 14433 1719 14467
rect 3893 14433 3927 14467
rect 6193 14433 6227 14467
rect 8677 14433 8711 14467
rect 9137 14433 9171 14467
rect 9965 14433 9999 14467
rect 10057 14433 10091 14467
rect 10425 14433 10459 14467
rect 11345 14433 11379 14467
rect 11621 14433 11655 14467
rect 13645 14433 13679 14467
rect 14013 14433 14047 14467
rect 15485 14433 15519 14467
rect 15577 14433 15611 14467
rect 15945 14433 15979 14467
rect 16037 14433 16071 14467
rect 17141 14433 17175 14467
rect 1409 14365 1443 14399
rect 4077 14365 4111 14399
rect 4353 14365 4387 14399
rect 6469 14365 6503 14399
rect 8769 14365 8803 14399
rect 9781 14365 9815 14399
rect 13001 14365 13035 14399
rect 14289 14365 14323 14399
rect 5457 14297 5491 14331
rect 18337 14433 18371 14467
rect 20177 14433 20211 14467
rect 22201 14433 22235 14467
rect 24409 14433 24443 14467
rect 26617 14433 26651 14467
rect 27813 14433 27847 14467
rect 28365 14433 28399 14467
rect 28549 14433 28583 14467
rect 29101 14433 29135 14467
rect 30113 14433 30147 14467
rect 30665 14433 30699 14467
rect 31309 14433 31343 14467
rect 32137 14433 32171 14467
rect 32965 14433 32999 14467
rect 33609 14433 33643 14467
rect 35725 14433 35759 14467
rect 36277 14433 36311 14467
rect 36553 14433 36587 14467
rect 37749 14433 37783 14467
rect 38301 14433 38335 14467
rect 18061 14365 18095 14399
rect 21925 14365 21959 14399
rect 24133 14365 24167 14399
rect 26525 14365 26559 14399
rect 29929 14365 29963 14399
rect 33885 14365 33919 14399
rect 38577 14365 38611 14399
rect 30573 14297 30607 14331
rect 31493 14297 31527 14331
rect 35817 14297 35851 14331
rect 3709 14229 3743 14263
rect 7757 14229 7791 14263
rect 17969 14229 18003 14263
rect 19441 14229 19475 14263
rect 20269 14229 20303 14263
rect 25513 14229 25547 14263
rect 26801 14229 26835 14263
rect 27905 14229 27939 14263
rect 32321 14229 32355 14263
rect 33057 14229 33091 14263
rect 10609 14025 10643 14059
rect 11529 14025 11563 14059
rect 12081 14025 12115 14059
rect 6193 13957 6227 13991
rect 6929 13957 6963 13991
rect 22109 13957 22143 13991
rect 9505 13889 9539 13923
rect 14013 13889 14047 13923
rect 17049 13889 17083 13923
rect 19441 13889 19475 13923
rect 21097 13889 21131 13923
rect 21833 13889 21867 13923
rect 22845 13889 22879 13923
rect 24317 13889 24351 13923
rect 24961 13889 24995 13923
rect 28089 13889 28123 13923
rect 29285 13889 29319 13923
rect 30021 13889 30055 13923
rect 30849 13889 30883 13923
rect 34161 13889 34195 13923
rect 35541 13889 35575 13923
rect 35817 13889 35851 13923
rect 38301 13889 38335 13923
rect 2689 13821 2723 13855
rect 3157 13821 3191 13855
rect 3433 13821 3467 13855
rect 6009 13821 6043 13855
rect 6837 13821 6871 13855
rect 7297 13821 7331 13855
rect 7573 13821 7607 13855
rect 8217 13821 8251 13855
rect 8769 13821 8803 13855
rect 9229 13821 9263 13855
rect 11345 13821 11379 13855
rect 12265 13821 12299 13855
rect 12541 13821 12575 13855
rect 12633 13821 12667 13855
rect 13369 13821 13403 13855
rect 13921 13821 13955 13855
rect 14933 13821 14967 13855
rect 15209 13821 15243 13855
rect 15669 13821 15703 13855
rect 15945 13821 15979 13855
rect 16221 13821 16255 13855
rect 16681 13821 16715 13855
rect 17233 13821 17267 13855
rect 18061 13821 18095 13855
rect 18429 13821 18463 13855
rect 18613 13821 18647 13855
rect 19717 13821 19751 13855
rect 22569 13821 22603 13855
rect 23673 13821 23707 13855
rect 24133 13821 24167 13855
rect 25053 13821 25087 13855
rect 26249 13821 26283 13855
rect 26341 13821 26375 13855
rect 26709 13821 26743 13855
rect 27169 13821 27203 13855
rect 27721 13821 27755 13855
rect 27997 13821 28031 13855
rect 29469 13821 29503 13855
rect 31401 13821 31435 13855
rect 31769 13821 31803 13855
rect 32137 13821 32171 13855
rect 32505 13821 32539 13855
rect 33241 13821 33275 13855
rect 33609 13821 33643 13855
rect 34069 13821 34103 13855
rect 38117 13821 38151 13855
rect 38485 13821 38519 13855
rect 25513 13753 25547 13787
rect 29653 13753 29687 13787
rect 31217 13753 31251 13787
rect 2513 13685 2547 13719
rect 4537 13685 4571 13719
rect 13277 13685 13311 13719
rect 14749 13685 14783 13719
rect 29561 13685 29595 13719
rect 36921 13685 36955 13719
rect 5641 13481 5675 13515
rect 6377 13481 6411 13515
rect 9045 13481 9079 13515
rect 21005 13481 21039 13515
rect 29377 13481 29411 13515
rect 32321 13481 32355 13515
rect 33241 13481 33275 13515
rect 25329 13413 25363 13447
rect 29469 13413 29503 13447
rect 29837 13413 29871 13447
rect 37197 13413 37231 13447
rect 4077 13345 4111 13379
rect 4353 13345 4387 13379
rect 6285 13345 6319 13379
rect 7481 13345 7515 13379
rect 7849 13345 7883 13379
rect 8861 13345 8895 13379
rect 10149 13345 10183 13379
rect 10425 13345 10459 13379
rect 10793 13345 10827 13379
rect 11437 13345 11471 13379
rect 11989 13345 12023 13379
rect 12449 13345 12483 13379
rect 13369 13345 13403 13379
rect 13737 13345 13771 13379
rect 14473 13345 14507 13379
rect 15761 13345 15795 13379
rect 16129 13345 16163 13379
rect 16405 13345 16439 13379
rect 16865 13345 16899 13379
rect 18613 13345 18647 13379
rect 19901 13345 19935 13379
rect 20361 13345 20395 13379
rect 21097 13345 21131 13379
rect 21465 13345 21499 13379
rect 23213 13345 23247 13379
rect 23489 13345 23523 13379
rect 24593 13345 24627 13379
rect 25053 13345 25087 13379
rect 27445 13345 27479 13379
rect 27629 13345 27663 13379
rect 27813 13345 27847 13379
rect 28089 13345 28123 13379
rect 28365 13345 28399 13379
rect 29285 13345 29319 13379
rect 30849 13345 30883 13379
rect 31309 13345 31343 13379
rect 32137 13345 32171 13379
rect 33333 13345 33367 13379
rect 33701 13345 33735 13379
rect 34161 13345 34195 13379
rect 34805 13345 34839 13379
rect 36093 13345 36127 13379
rect 36553 13345 36587 13379
rect 36737 13345 36771 13379
rect 37749 13345 37783 13379
rect 38301 13345 38335 13379
rect 1409 13277 1443 13311
rect 1685 13277 1719 13311
rect 7113 13277 7147 13311
rect 12633 13277 12667 13311
rect 15485 13277 15519 13311
rect 17877 13277 17911 13311
rect 19073 13277 19107 13311
rect 19993 13277 20027 13311
rect 21741 13277 21775 13311
rect 22477 13277 22511 13311
rect 24317 13277 24351 13311
rect 26985 13277 27019 13311
rect 29101 13277 29135 13311
rect 30665 13277 30699 13311
rect 38577 13277 38611 13311
rect 7757 13209 7791 13243
rect 13185 13209 13219 13243
rect 18337 13209 18371 13243
rect 22937 13209 22971 13243
rect 31309 13209 31343 13243
rect 37841 13209 37875 13243
rect 2973 13141 3007 13175
rect 14657 13141 14691 13175
rect 17049 13141 17083 13175
rect 34989 13141 35023 13175
rect 2789 12937 2823 12971
rect 4905 12937 4939 12971
rect 6193 12937 6227 12971
rect 14105 12937 14139 12971
rect 24593 12937 24627 12971
rect 36921 12937 36955 12971
rect 12541 12869 12575 12903
rect 18521 12869 18555 12903
rect 22661 12869 22695 12903
rect 1409 12801 1443 12835
rect 3801 12801 3835 12835
rect 7021 12801 7055 12835
rect 7297 12801 7331 12835
rect 9505 12801 9539 12835
rect 14841 12801 14875 12835
rect 15761 12801 15795 12835
rect 17233 12801 17267 12835
rect 19165 12801 19199 12835
rect 20453 12801 20487 12835
rect 22017 12801 22051 12835
rect 27629 12801 27663 12835
rect 30113 12801 30147 12835
rect 30849 12801 30883 12835
rect 32689 12801 32723 12835
rect 37749 12801 37783 12835
rect 39129 12801 39163 12835
rect 1685 12733 1719 12767
rect 3525 12733 3559 12767
rect 6101 12733 6135 12767
rect 9137 12733 9171 12767
rect 9689 12733 9723 12767
rect 10333 12733 10367 12767
rect 10701 12733 10735 12767
rect 10885 12733 10919 12767
rect 11713 12733 11747 12767
rect 12725 12733 12759 12767
rect 13185 12733 13219 12767
rect 13921 12733 13955 12767
rect 15117 12733 15151 12767
rect 15577 12733 15611 12767
rect 16221 12733 16255 12767
rect 16957 12733 16991 12767
rect 18061 12733 18095 12767
rect 18797 12733 18831 12767
rect 19993 12733 20027 12767
rect 20545 12733 20579 12767
rect 20913 12733 20947 12767
rect 21097 12733 21131 12767
rect 22201 12733 22235 12767
rect 22661 12733 22695 12767
rect 24501 12733 24535 12767
rect 25789 12733 25823 12767
rect 26525 12733 26559 12767
rect 27813 12733 27847 12767
rect 29285 12733 29319 12767
rect 30389 12733 30423 12767
rect 31309 12733 31343 12767
rect 31677 12733 31711 12767
rect 32045 12733 32079 12767
rect 32597 12733 32631 12767
rect 33241 12733 33275 12767
rect 33609 12733 33643 12767
rect 34069 12733 34103 12767
rect 34897 12733 34931 12767
rect 35541 12733 35575 12767
rect 36093 12733 36127 12767
rect 36277 12733 36311 12767
rect 36829 12733 36863 12767
rect 37473 12733 37507 12767
rect 8677 12665 8711 12699
rect 27077 12665 27111 12699
rect 27997 12665 28031 12699
rect 28365 12665 28399 12699
rect 30481 12665 30515 12699
rect 34345 12665 34379 12699
rect 34989 12665 35023 12699
rect 11805 12597 11839 12631
rect 16313 12597 16347 12631
rect 27905 12597 27939 12631
rect 29469 12597 29503 12631
rect 30297 12597 30331 12631
rect 3249 12393 3283 12427
rect 29377 12393 29411 12427
rect 30205 12393 30239 12427
rect 16773 12325 16807 12359
rect 18429 12325 18463 12359
rect 25789 12325 25823 12359
rect 30389 12325 30423 12359
rect 1869 12257 1903 12291
rect 4629 12257 4663 12291
rect 5549 12257 5583 12291
rect 6009 12257 6043 12291
rect 6285 12257 6319 12291
rect 6653 12257 6687 12291
rect 7297 12257 7331 12291
rect 8033 12257 8067 12291
rect 8401 12257 8435 12291
rect 8769 12257 8803 12291
rect 9965 12257 9999 12291
rect 10333 12257 10367 12291
rect 10701 12257 10735 12291
rect 11529 12257 11563 12291
rect 11805 12257 11839 12291
rect 12081 12257 12115 12291
rect 13001 12257 13035 12291
rect 13369 12257 13403 12291
rect 14013 12257 14047 12291
rect 14197 12257 14231 12291
rect 15301 12257 15335 12291
rect 15853 12257 15887 12291
rect 17417 12257 17451 12291
rect 17785 12257 17819 12291
rect 19073 12257 19107 12291
rect 19441 12257 19475 12291
rect 20085 12257 20119 12291
rect 20913 12257 20947 12291
rect 21465 12257 21499 12291
rect 22477 12257 22511 12291
rect 22937 12257 22971 12291
rect 23029 12257 23063 12291
rect 24409 12257 24443 12291
rect 26985 12257 27019 12291
rect 27629 12257 27663 12291
rect 28273 12257 28307 12291
rect 29193 12257 29227 12291
rect 30297 12257 30331 12291
rect 31217 12257 31251 12291
rect 32137 12257 32171 12291
rect 32597 12257 32631 12291
rect 32873 12257 32907 12291
rect 33333 12257 33367 12291
rect 34069 12257 34103 12291
rect 37013 12257 37047 12291
rect 38393 12257 38427 12291
rect 38577 12257 38611 12291
rect 38761 12257 38795 12291
rect 2145 12189 2179 12223
rect 6377 12189 6411 12223
rect 8309 12189 8343 12223
rect 10149 12189 10183 12223
rect 12541 12189 12575 12223
rect 17325 12189 17359 12223
rect 17877 12189 17911 12223
rect 18981 12189 19015 12223
rect 19533 12189 19567 12223
rect 22385 12189 22419 12223
rect 23581 12189 23615 12223
rect 24133 12189 24167 12223
rect 27077 12189 27111 12223
rect 28457 12189 28491 12223
rect 30021 12189 30055 12223
rect 30757 12189 30791 12223
rect 33057 12189 33091 12223
rect 34529 12189 34563 12223
rect 34805 12189 34839 12223
rect 35909 12189 35943 12223
rect 37105 12189 37139 12223
rect 15393 12121 15427 12155
rect 21005 12121 21039 12155
rect 27905 12121 27939 12155
rect 4445 12053 4479 12087
rect 20269 12053 20303 12087
rect 31309 12053 31343 12087
rect 4721 11849 4755 11883
rect 8401 11849 8435 11883
rect 9321 11849 9355 11883
rect 12633 11849 12667 11883
rect 18245 11849 18279 11883
rect 28549 11849 28583 11883
rect 32137 11849 32171 11883
rect 15761 11781 15795 11815
rect 19165 11781 19199 11815
rect 20729 11781 20763 11815
rect 22293 11781 22327 11815
rect 31493 11781 31527 11815
rect 33517 11781 33551 11815
rect 35633 11781 35667 11815
rect 3341 11713 3375 11747
rect 7113 11713 7147 11747
rect 10793 11713 10827 11747
rect 13829 11713 13863 11747
rect 29469 11713 29503 11747
rect 34253 11713 34287 11747
rect 37473 11713 37507 11747
rect 37749 11713 37783 11747
rect 2697 11645 2731 11679
rect 3617 11645 3651 11679
rect 6837 11645 6871 11679
rect 9229 11645 9263 11679
rect 9873 11645 9907 11679
rect 10241 11645 10275 11679
rect 10885 11645 10919 11679
rect 11529 11645 11563 11679
rect 12449 11645 12483 11679
rect 13461 11645 13495 11679
rect 13921 11645 13955 11679
rect 14197 11645 14231 11679
rect 15393 11645 15427 11679
rect 15669 11645 15703 11679
rect 16221 11645 16255 11679
rect 16313 11645 16347 11679
rect 17233 11645 17267 11679
rect 18061 11645 18095 11679
rect 19073 11645 19107 11679
rect 19625 11645 19659 11679
rect 19901 11645 19935 11679
rect 20637 11645 20671 11679
rect 21005 11645 21039 11679
rect 21465 11645 21499 11679
rect 22109 11645 22143 11679
rect 22569 11645 22603 11679
rect 22937 11645 22971 11679
rect 25421 11645 25455 11679
rect 26157 11645 26191 11679
rect 26709 11645 26743 11679
rect 27169 11645 27203 11679
rect 27353 11645 27387 11679
rect 27721 11645 27755 11679
rect 27905 11645 27939 11679
rect 28089 11645 28123 11679
rect 29377 11645 29411 11679
rect 30113 11645 30147 11679
rect 30205 11645 30239 11679
rect 30573 11645 30607 11679
rect 31309 11645 31343 11679
rect 32321 11645 32355 11679
rect 32781 11645 32815 11679
rect 33425 11645 33459 11679
rect 33977 11645 34011 11679
rect 35817 11645 35851 11679
rect 36001 11645 36035 11679
rect 36185 11645 36219 11679
rect 2789 11509 2823 11543
rect 11713 11509 11747 11543
rect 15393 11509 15427 11543
rect 17417 11509 17451 11543
rect 38853 11509 38887 11543
rect 7849 11305 7883 11339
rect 11069 11305 11103 11339
rect 14381 11305 14415 11339
rect 16681 11305 16715 11339
rect 19165 11305 19199 11339
rect 21097 11305 21131 11339
rect 25237 11305 25271 11339
rect 36921 11305 36955 11339
rect 38853 11305 38887 11339
rect 10425 11237 10459 11271
rect 25881 11237 25915 11271
rect 27261 11237 27295 11271
rect 38301 11237 38335 11271
rect 1961 11169 1995 11203
rect 2789 11169 2823 11203
rect 2973 11169 3007 11203
rect 5457 11169 5491 11203
rect 5917 11169 5951 11203
rect 6285 11169 6319 11203
rect 6653 11169 6687 11203
rect 7205 11169 7239 11203
rect 7757 11169 7791 11203
rect 8401 11169 8435 11203
rect 8861 11169 8895 11203
rect 9689 11169 9723 11203
rect 10149 11169 10183 11203
rect 11253 11169 11287 11203
rect 11989 11169 12023 11203
rect 12357 11169 12391 11203
rect 12449 11169 12483 11203
rect 13001 11169 13035 11203
rect 13553 11169 13587 11203
rect 14197 11169 14231 11203
rect 15577 11169 15611 11203
rect 17969 11169 18003 11203
rect 18429 11169 18463 11203
rect 19073 11169 19107 11203
rect 19441 11169 19475 11203
rect 20085 11169 20119 11203
rect 21005 11169 21039 11203
rect 21557 11169 21591 11203
rect 22569 11169 22603 11203
rect 23489 11169 23523 11203
rect 24041 11169 24075 11203
rect 24225 11169 24259 11203
rect 25145 11169 25179 11203
rect 25789 11169 25823 11203
rect 26525 11169 26559 11203
rect 26985 11169 27019 11203
rect 28181 11169 28215 11203
rect 28917 11169 28951 11203
rect 29285 11169 29319 11203
rect 29469 11169 29503 11203
rect 30573 11169 30607 11203
rect 30941 11169 30975 11203
rect 31033 11169 31067 11203
rect 32137 11169 32171 11203
rect 32505 11169 32539 11203
rect 33057 11169 33091 11203
rect 33701 11169 33735 11203
rect 34253 11169 34287 11203
rect 35817 11169 35851 11203
rect 37841 11169 37875 11203
rect 38761 11169 38795 11203
rect 9137 11101 9171 11135
rect 11897 11101 11931 11135
rect 13369 11101 13403 11135
rect 15301 11101 15335 11135
rect 22017 11101 22051 11135
rect 22661 11101 22695 11135
rect 23305 11101 23339 11135
rect 28733 11101 28767 11135
rect 30665 11101 30699 11135
rect 32965 11101 32999 11135
rect 34529 11101 34563 11135
rect 35541 11101 35575 11135
rect 37749 11101 37783 11135
rect 2697 11033 2731 11067
rect 5549 11033 5583 11067
rect 11437 11033 11471 11067
rect 17785 11033 17819 11067
rect 20269 11033 20303 11067
rect 27997 11033 28031 11067
rect 28549 11033 28583 11067
rect 33977 11033 34011 11067
rect 24501 10965 24535 10999
rect 30205 10965 30239 10999
rect 2789 10761 2823 10795
rect 4905 10761 4939 10795
rect 6009 10761 6043 10795
rect 16773 10761 16807 10795
rect 27169 10761 27203 10795
rect 34989 10761 35023 10795
rect 37749 10761 37783 10795
rect 11161 10693 11195 10727
rect 12541 10693 12575 10727
rect 19257 10693 19291 10727
rect 23949 10693 23983 10727
rect 6837 10625 6871 10659
rect 9689 10625 9723 10659
rect 13921 10625 13955 10659
rect 22017 10625 22051 10659
rect 23029 10625 23063 10659
rect 28733 10625 28767 10659
rect 29745 10625 29779 10659
rect 32781 10625 32815 10659
rect 36185 10625 36219 10659
rect 1409 10557 1443 10591
rect 1685 10557 1719 10591
rect 3525 10557 3559 10591
rect 3801 10557 3835 10591
rect 5917 10557 5951 10591
rect 7113 10557 7147 10591
rect 9321 10557 9355 10591
rect 9873 10557 9907 10591
rect 11345 10557 11379 10591
rect 11529 10557 11563 10591
rect 11713 10557 11747 10591
rect 12449 10557 12483 10591
rect 13001 10557 13035 10591
rect 14013 10557 14047 10591
rect 14289 10557 14323 10591
rect 14841 10557 14875 10591
rect 15117 10557 15151 10591
rect 15761 10557 15795 10591
rect 16405 10557 16439 10591
rect 16957 10557 16991 10591
rect 17325 10557 17359 10591
rect 18061 10557 18095 10591
rect 18889 10557 18923 10591
rect 19625 10557 19659 10591
rect 19901 10557 19935 10591
rect 20821 10557 20855 10591
rect 21005 10557 21039 10591
rect 21741 10557 21775 10591
rect 22845 10557 22879 10591
rect 22937 10557 22971 10591
rect 23765 10557 23799 10591
rect 24685 10557 24719 10591
rect 24915 10557 24949 10591
rect 25053 10557 25087 10591
rect 25513 10557 25547 10591
rect 25697 10557 25731 10591
rect 26985 10557 27019 10591
rect 28273 10557 28307 10591
rect 28549 10557 28583 10591
rect 29653 10557 29687 10591
rect 30297 10557 30331 10591
rect 30665 10557 30699 10591
rect 30849 10557 30883 10591
rect 32045 10557 32079 10591
rect 32321 10557 32355 10591
rect 32505 10557 32539 10591
rect 33057 10557 33091 10591
rect 33701 10557 33735 10591
rect 34897 10557 34931 10591
rect 35449 10557 35483 10591
rect 36461 10557 36495 10591
rect 8493 10489 8527 10523
rect 27721 10489 27755 10523
rect 16221 10421 16255 10455
rect 18245 10421 18279 10455
rect 20637 10421 20671 10455
rect 21097 10421 21131 10455
rect 22661 10421 22695 10455
rect 24501 10421 24535 10455
rect 25973 10421 26007 10455
rect 33885 10421 33919 10455
rect 2789 10217 2823 10251
rect 6009 10217 6043 10251
rect 9781 10217 9815 10251
rect 23581 10217 23615 10251
rect 25697 10217 25731 10251
rect 28273 10217 28307 10251
rect 29193 10217 29227 10251
rect 29285 10217 29319 10251
rect 33149 10217 33183 10251
rect 34805 10217 34839 10251
rect 11253 10149 11287 10183
rect 14565 10149 14599 10183
rect 18981 10149 19015 10183
rect 29009 10149 29043 10183
rect 29377 10149 29411 10183
rect 29745 10149 29779 10183
rect 1685 10081 1719 10115
rect 3801 10081 3835 10115
rect 4721 10081 4755 10115
rect 6561 10081 6595 10115
rect 7205 10081 7239 10115
rect 7297 10081 7331 10115
rect 7757 10081 7791 10115
rect 8493 10081 8527 10115
rect 8953 10081 8987 10115
rect 9689 10081 9723 10115
rect 10149 10081 10183 10115
rect 11897 10081 11931 10115
rect 12265 10081 12299 10115
rect 13185 10081 13219 10115
rect 15853 10081 15887 10115
rect 16497 10081 16531 10115
rect 16589 10081 16623 10115
rect 17141 10081 17175 10115
rect 17509 10081 17543 10115
rect 18245 10081 18279 10115
rect 19625 10081 19659 10115
rect 19993 10081 20027 10115
rect 20913 10081 20947 10115
rect 21465 10081 21499 10115
rect 22201 10081 22235 10115
rect 30205 10081 30239 10115
rect 30941 10081 30975 10115
rect 31217 10081 31251 10115
rect 32249 10081 32283 10115
rect 33333 10081 33367 10115
rect 33701 10081 33735 10115
rect 35817 10081 35851 10115
rect 37197 10081 37231 10115
rect 37933 10081 37967 10115
rect 38117 10081 38151 10115
rect 38393 10081 38427 10115
rect 38945 10081 38979 10115
rect 1409 10013 1443 10047
rect 4445 10013 4479 10047
rect 7113 10013 7147 10047
rect 9045 10013 9079 10047
rect 11805 10013 11839 10047
rect 12357 10013 12391 10047
rect 12909 10013 12943 10047
rect 19717 10013 19751 10047
rect 20085 10013 20119 10047
rect 21281 10013 21315 10047
rect 22477 10013 22511 10047
rect 24317 10013 24351 10047
rect 24593 10013 24627 10047
rect 26893 10013 26927 10047
rect 27169 10013 27203 10047
rect 32137 10013 32171 10047
rect 33425 10013 33459 10047
rect 35541 10013 35575 10047
rect 16129 9945 16163 9979
rect 30389 9945 30423 9979
rect 3617 9877 3651 9911
rect 18429 9877 18463 9911
rect 32413 9877 32447 9911
rect 39037 9877 39071 9911
rect 3893 9673 3927 9707
rect 9321 9673 9355 9707
rect 18337 9673 18371 9707
rect 12633 9605 12667 9639
rect 20821 9605 20855 9639
rect 24869 9605 24903 9639
rect 26893 9605 26927 9639
rect 28549 9605 28583 9639
rect 30849 9605 30883 9639
rect 35081 9605 35115 9639
rect 2605 9537 2639 9571
rect 7665 9537 7699 9571
rect 15117 9537 15151 9571
rect 21373 9537 21407 9571
rect 25513 9537 25547 9571
rect 25789 9537 25823 9571
rect 29377 9537 29411 9571
rect 30205 9537 30239 9571
rect 32965 9537 32999 9571
rect 37013 9537 37047 9571
rect 2329 9469 2363 9503
rect 4629 9469 4663 9503
rect 4905 9469 4939 9503
rect 7021 9469 7055 9503
rect 7389 9469 7423 9503
rect 7757 9469 7791 9503
rect 8585 9469 8619 9503
rect 9873 9469 9907 9503
rect 9965 9469 9999 9503
rect 10241 9469 10275 9503
rect 10425 9469 10459 9503
rect 11345 9469 11379 9503
rect 11529 9469 11563 9503
rect 11713 9469 11747 9503
rect 12449 9469 12483 9503
rect 13185 9469 13219 9503
rect 14381 9469 14415 9503
rect 14657 9469 14691 9503
rect 14933 9469 14967 9503
rect 15485 9469 15519 9503
rect 15853 9469 15887 9503
rect 16589 9469 16623 9503
rect 16681 9469 16715 9503
rect 17233 9469 17267 9503
rect 18245 9469 18279 9503
rect 18613 9469 18647 9503
rect 18981 9469 19015 9503
rect 19901 9469 19935 9503
rect 20637 9469 20671 9503
rect 21097 9469 21131 9503
rect 22109 9469 22143 9503
rect 22477 9469 22511 9503
rect 22661 9469 22695 9503
rect 23489 9469 23523 9503
rect 23673 9469 23707 9503
rect 23857 9469 23891 9503
rect 24317 9469 24351 9503
rect 24409 9469 24443 9503
rect 27629 9469 27663 9503
rect 27997 9469 28031 9503
rect 28549 9469 28583 9503
rect 29653 9469 29687 9503
rect 30113 9469 30147 9503
rect 31033 9469 31067 9503
rect 31125 9469 31159 9503
rect 31861 9469 31895 9503
rect 32229 9469 32263 9503
rect 32781 9469 32815 9503
rect 33425 9469 33459 9503
rect 33793 9469 33827 9503
rect 33977 9469 34011 9503
rect 34897 9469 34931 9503
rect 36001 9469 36035 9503
rect 36185 9469 36219 9503
rect 36829 9469 36863 9503
rect 37473 9469 37507 9503
rect 37749 9469 37783 9503
rect 10885 9401 10919 9435
rect 19993 9401 20027 9435
rect 6193 9333 6227 9367
rect 8677 9333 8711 9367
rect 13369 9333 13403 9367
rect 17417 9333 17451 9367
rect 23305 9333 23339 9367
rect 31309 9333 31343 9367
rect 37289 9333 37323 9367
rect 38853 9333 38887 9367
rect 2881 9129 2915 9163
rect 7849 9129 7883 9163
rect 17417 9129 17451 9163
rect 19717 9129 19751 9163
rect 22661 9129 22695 9163
rect 23397 9129 23431 9163
rect 26617 9129 26651 9163
rect 28917 9129 28951 9163
rect 29561 9129 29595 9163
rect 32229 9129 32263 9163
rect 9689 9061 9723 9095
rect 11529 9061 11563 9095
rect 27261 9061 27295 9095
rect 1777 8993 1811 9027
rect 2237 8993 2271 9027
rect 3065 8993 3099 9027
rect 3341 8993 3375 9027
rect 4077 8993 4111 9027
rect 4353 8993 4387 9027
rect 5365 8993 5399 9027
rect 6009 8993 6043 9027
rect 6377 8993 6411 9027
rect 6745 8993 6779 9027
rect 7205 8993 7239 9027
rect 7757 8993 7791 9027
rect 9505 8993 9539 9027
rect 10333 8993 10367 9027
rect 10425 8993 10459 9027
rect 10701 8993 10735 9027
rect 12173 8993 12207 9027
rect 12265 8993 12299 9027
rect 12541 8993 12575 9027
rect 12633 8993 12667 9027
rect 13369 8993 13403 9027
rect 13829 8993 13863 9027
rect 14289 8993 14323 9027
rect 16129 8993 16163 9027
rect 17969 8993 18003 9027
rect 18613 8993 18647 9027
rect 18981 8993 19015 9027
rect 19625 8993 19659 9027
rect 20177 8993 20211 9027
rect 21281 8993 21315 9027
rect 21741 8993 21775 9027
rect 22477 8993 22511 9027
rect 23213 8993 23247 9027
rect 24317 8993 24351 9027
rect 24409 8993 24443 9027
rect 24777 8993 24811 9027
rect 24869 8993 24903 9027
rect 26525 8993 26559 9027
rect 27813 8993 27847 9027
rect 28089 8993 28123 9027
rect 28273 8993 28307 9027
rect 28733 8993 28767 9027
rect 29745 8993 29779 9027
rect 30757 8993 30791 9027
rect 31401 8993 31435 9027
rect 31493 8993 31527 9027
rect 1869 8925 1903 8959
rect 4169 8925 4203 8959
rect 4629 8925 4663 8959
rect 5457 8925 5491 8959
rect 10793 8925 10827 8959
rect 15853 8925 15887 8959
rect 21005 8925 21039 8959
rect 29929 8925 29963 8959
rect 30481 8925 30515 8959
rect 30941 8925 30975 8959
rect 32781 8993 32815 9027
rect 32965 8993 32999 9027
rect 33149 8993 33183 9027
rect 34345 8993 34379 9027
rect 36001 8993 36035 9027
rect 36553 8993 36587 9027
rect 38301 8993 38335 9027
rect 38577 8993 38611 9027
rect 34621 8925 34655 8959
rect 36461 8925 36495 8959
rect 37749 8925 37783 8959
rect 38439 8925 38473 8959
rect 18061 8857 18095 8891
rect 21741 8857 21775 8891
rect 25237 8857 25271 8891
rect 32229 8857 32263 8891
rect 32597 8857 32631 8891
rect 9321 8789 9355 8823
rect 13185 8789 13219 8823
rect 13829 8789 13863 8823
rect 36737 8789 36771 8823
rect 10793 8585 10827 8619
rect 17509 8585 17543 8619
rect 21281 8585 21315 8619
rect 27905 8585 27939 8619
rect 37933 8585 37967 8619
rect 3525 8517 3559 8551
rect 24133 8517 24167 8551
rect 28641 8517 28675 8551
rect 7849 8449 7883 8483
rect 9965 8449 9999 8483
rect 11253 8449 11287 8483
rect 13001 8449 13035 8483
rect 13829 8449 13863 8483
rect 18153 8449 18187 8483
rect 19993 8449 20027 8483
rect 22385 8449 22419 8483
rect 24961 8449 24995 8483
rect 27169 8449 27203 8483
rect 29285 8449 29319 8483
rect 30941 8449 30975 8483
rect 32045 8449 32079 8483
rect 32781 8449 32815 8483
rect 36001 8449 36035 8483
rect 36829 8449 36863 8483
rect 38761 8449 38795 8483
rect 3249 8381 3283 8415
rect 3617 8381 3651 8415
rect 6929 8381 6963 8415
rect 7573 8381 7607 8415
rect 7941 8381 7975 8415
rect 8585 8381 8619 8415
rect 8861 8381 8895 8415
rect 11345 8381 11379 8415
rect 11713 8381 11747 8415
rect 11897 8381 11931 8415
rect 12449 8381 12483 8415
rect 12909 8381 12943 8415
rect 13737 8381 13771 8415
rect 14105 8381 14139 8415
rect 14657 8381 14691 8415
rect 15025 8381 15059 8415
rect 15577 8381 15611 8415
rect 16037 8381 16071 8415
rect 16773 8381 16807 8415
rect 17693 8381 17727 8415
rect 18245 8381 18279 8415
rect 18613 8381 18647 8415
rect 19073 8381 19107 8415
rect 19717 8381 19751 8415
rect 22017 8381 22051 8415
rect 22293 8381 22327 8415
rect 22569 8381 22603 8415
rect 24041 8381 24075 8415
rect 24685 8381 24719 8415
rect 26341 8381 26375 8415
rect 27077 8381 27111 8415
rect 27721 8381 27755 8415
rect 28457 8381 28491 8415
rect 29561 8381 29595 8415
rect 31493 8381 31527 8415
rect 31585 8381 31619 8415
rect 32505 8381 32539 8415
rect 35081 8381 35115 8415
rect 35541 8381 35575 8415
rect 35909 8381 35943 8415
rect 36553 8381 36587 8415
rect 38669 8381 38703 8415
rect 16221 8245 16255 8279
rect 16957 8245 16991 8279
rect 33885 8245 33919 8279
rect 3249 8041 3283 8075
rect 6469 8041 6503 8075
rect 11621 8041 11655 8075
rect 21281 8041 21315 8075
rect 24041 8041 24075 8075
rect 27905 8041 27939 8075
rect 32229 8041 32263 8075
rect 25881 7973 25915 8007
rect 29469 7973 29503 8007
rect 33333 7973 33367 8007
rect 2145 7905 2179 7939
rect 4169 7905 4203 7939
rect 5089 7905 5123 7939
rect 5365 7905 5399 7939
rect 7481 7905 7515 7939
rect 8033 7905 8067 7939
rect 8401 7905 8435 7939
rect 9873 7905 9907 7939
rect 10057 7905 10091 7939
rect 10517 7905 10551 7939
rect 11805 7905 11839 7939
rect 12081 7905 12115 7939
rect 13001 7905 13035 7939
rect 15301 7905 15335 7939
rect 16221 7905 16255 7939
rect 16589 7905 16623 7939
rect 17141 7905 17175 7939
rect 17325 7905 17359 7939
rect 18245 7905 18279 7939
rect 18613 7905 18647 7939
rect 19257 7905 19291 7939
rect 19901 7905 19935 7939
rect 21189 7905 21223 7939
rect 23949 7905 23983 7939
rect 24777 7905 24811 7939
rect 25329 7905 25363 7939
rect 25513 7905 25547 7939
rect 26801 7905 26835 7939
rect 28641 7905 28675 7939
rect 30021 7905 30055 7939
rect 30297 7905 30331 7939
rect 30481 7905 30515 7939
rect 31125 7905 31159 7939
rect 32137 7905 32171 7939
rect 32873 7905 32907 7939
rect 36093 7905 36127 7939
rect 36645 7905 36679 7939
rect 37013 7905 37047 7939
rect 37933 7905 37967 7939
rect 38117 7905 38151 7939
rect 38485 7905 38519 7939
rect 1869 7837 1903 7871
rect 7665 7837 7699 7871
rect 12725 7837 12759 7871
rect 16497 7837 16531 7871
rect 21833 7837 21867 7871
rect 22109 7837 22143 7871
rect 24685 7837 24719 7871
rect 26525 7837 26559 7871
rect 31033 7837 31067 7871
rect 32781 7837 32815 7871
rect 33793 7837 33827 7871
rect 34069 7837 34103 7871
rect 38393 7837 38427 7871
rect 10517 7769 10551 7803
rect 17509 7769 17543 7803
rect 36921 7769 36955 7803
rect 4261 7701 4295 7735
rect 14105 7701 14139 7735
rect 15485 7701 15519 7735
rect 16037 7701 16071 7735
rect 18337 7701 18371 7735
rect 20085 7701 20119 7735
rect 23213 7701 23247 7735
rect 28825 7701 28859 7735
rect 31309 7701 31343 7735
rect 35357 7701 35391 7735
rect 3157 7497 3191 7531
rect 5181 7497 5215 7531
rect 25053 7497 25087 7531
rect 26249 7497 26283 7531
rect 31309 7497 31343 7531
rect 36553 7497 36587 7531
rect 7665 7429 7699 7463
rect 22293 7429 22327 7463
rect 29377 7429 29411 7463
rect 2145 7361 2179 7395
rect 2605 7361 2639 7395
rect 4077 7361 4111 7395
rect 7021 7361 7055 7395
rect 9873 7361 9907 7395
rect 13001 7361 13035 7395
rect 14013 7361 14047 7395
rect 18981 7361 19015 7395
rect 20821 7361 20855 7395
rect 23673 7361 23707 7395
rect 27629 7361 27663 7395
rect 28181 7361 28215 7395
rect 28733 7361 28767 7395
rect 30205 7361 30239 7395
rect 32505 7361 32539 7395
rect 35449 7361 35483 7395
rect 37841 7361 37875 7395
rect 2421 7293 2455 7327
rect 3065 7293 3099 7327
rect 3801 7293 3835 7327
rect 7389 7293 7423 7327
rect 7665 7293 7699 7327
rect 8953 7293 8987 7327
rect 9229 7293 9263 7327
rect 9505 7293 9539 7327
rect 10609 7293 10643 7327
rect 10885 7293 10919 7327
rect 11529 7293 11563 7327
rect 12449 7293 12483 7327
rect 12909 7293 12943 7327
rect 13829 7293 13863 7327
rect 13921 7293 13955 7327
rect 14473 7293 14507 7327
rect 14657 7293 14691 7327
rect 15301 7293 15335 7327
rect 15577 7293 15611 7327
rect 16681 7293 16715 7327
rect 16865 7293 16899 7327
rect 17141 7293 17175 7327
rect 18245 7293 18279 7327
rect 18429 7293 18463 7327
rect 18889 7293 18923 7327
rect 19901 7293 19935 7327
rect 19993 7293 20027 7327
rect 20453 7293 20487 7327
rect 21557 7293 21591 7327
rect 22017 7293 22051 7327
rect 22385 7293 22419 7327
rect 23213 7293 23247 7327
rect 23949 7293 23983 7327
rect 26157 7293 26191 7327
rect 26801 7293 26835 7327
rect 27537 7293 27571 7327
rect 28273 7293 28307 7327
rect 29285 7293 29319 7327
rect 29929 7293 29963 7327
rect 32229 7293 32263 7327
rect 35173 7293 35207 7327
rect 37749 7293 37783 7327
rect 37933 7293 37967 7327
rect 38301 7293 38335 7327
rect 38853 7293 38887 7327
rect 1593 7225 1627 7259
rect 33885 7225 33919 7259
rect 10425 7157 10459 7191
rect 11713 7157 11747 7191
rect 13645 7157 13679 7191
rect 23029 7157 23063 7191
rect 26985 7157 27019 7191
rect 7849 6953 7883 6987
rect 9965 6953 9999 6987
rect 29285 6953 29319 6987
rect 15393 6885 15427 6919
rect 24133 6885 24167 6919
rect 2421 6817 2455 6851
rect 2973 6817 3007 6851
rect 3157 6817 3191 6851
rect 5089 6817 5123 6851
rect 5273 6817 5307 6851
rect 5457 6817 5491 6851
rect 6561 6817 6595 6851
rect 8953 6817 8987 6851
rect 9965 6817 9999 6851
rect 10241 6817 10275 6851
rect 11437 6817 11471 6851
rect 11529 6817 11563 6851
rect 11989 6817 12023 6851
rect 12173 6817 12207 6851
rect 13369 6817 13403 6851
rect 14749 6817 14783 6851
rect 15301 6817 15335 6851
rect 16497 6817 16531 6851
rect 16773 6817 16807 6851
rect 18153 6817 18187 6851
rect 19441 6817 19475 6851
rect 19809 6817 19843 6851
rect 20177 6817 20211 6851
rect 21097 6817 21131 6851
rect 21465 6817 21499 6851
rect 22017 6817 22051 6851
rect 22845 6817 22879 6851
rect 23029 6817 23063 6851
rect 23581 6817 23615 6851
rect 23765 6817 23799 6851
rect 24685 6817 24719 6851
rect 25421 6817 25455 6851
rect 26985 6817 27019 6851
rect 30665 6817 30699 6851
rect 31493 6817 31527 6851
rect 32321 6817 32355 6851
rect 33517 6817 33551 6851
rect 33793 6817 33827 6851
rect 35265 6817 35299 6851
rect 36737 6817 36771 6851
rect 38025 6817 38059 6851
rect 38393 6817 38427 6851
rect 38669 6817 38703 6851
rect 4629 6749 4663 6783
rect 6285 6749 6319 6783
rect 13093 6749 13127 6783
rect 19349 6749 19383 6783
rect 21281 6749 21315 6783
rect 27721 6749 27755 6783
rect 27997 6749 28031 6783
rect 29837 6749 29871 6783
rect 30389 6749 30423 6783
rect 30849 6749 30883 6783
rect 32965 6749 32999 6783
rect 33977 6749 34011 6783
rect 34437 6749 34471 6783
rect 34989 6749 35023 6783
rect 35449 6749 35483 6783
rect 35909 6749 35943 6783
rect 36461 6749 36495 6783
rect 36921 6749 36955 6783
rect 2973 6681 3007 6715
rect 9045 6681 9079 6715
rect 32413 6681 32447 6715
rect 37933 6681 37967 6715
rect 12449 6613 12483 6647
rect 24869 6613 24903 6647
rect 25605 6613 25639 6647
rect 27169 6613 27203 6647
rect 31309 6613 31343 6647
rect 6009 6409 6043 6443
rect 9505 6409 9539 6443
rect 13553 6409 13587 6443
rect 20085 6409 20119 6443
rect 20913 6409 20947 6443
rect 23029 6409 23063 6443
rect 26709 6409 26743 6443
rect 31677 6409 31711 6443
rect 35265 6409 35299 6443
rect 38853 6409 38887 6443
rect 3801 6341 3835 6375
rect 16681 6341 16715 6375
rect 27445 6341 27479 6375
rect 30021 6341 30055 6375
rect 2605 6273 2639 6307
rect 3985 6273 4019 6307
rect 7941 6273 7975 6307
rect 10241 6273 10275 6307
rect 14289 6273 14323 6307
rect 18981 6273 19015 6307
rect 25329 6273 25363 6307
rect 27721 6273 27755 6307
rect 32689 6273 32723 6307
rect 37473 6273 37507 6307
rect 37749 6273 37783 6307
rect 2145 6205 2179 6239
rect 2329 6205 2363 6239
rect 3341 6205 3375 6239
rect 3893 6205 3927 6239
rect 4629 6205 4663 6239
rect 4905 6205 4939 6239
rect 8217 6205 8251 6239
rect 10517 6205 10551 6239
rect 11897 6205 11931 6239
rect 12449 6205 12483 6239
rect 13461 6205 13495 6239
rect 14105 6205 14139 6239
rect 14565 6205 14599 6239
rect 14841 6205 14875 6239
rect 15485 6205 15519 6239
rect 15761 6205 15795 6239
rect 16497 6205 16531 6239
rect 17233 6205 17267 6239
rect 18061 6205 18095 6239
rect 18705 6205 18739 6239
rect 20821 6205 20855 6239
rect 21189 6205 21223 6239
rect 21833 6205 21867 6239
rect 22937 6205 22971 6239
rect 24409 6205 24443 6239
rect 24685 6205 24719 6239
rect 24869 6205 24903 6239
rect 25605 6205 25639 6239
rect 27629 6205 27663 6239
rect 28273 6205 28307 6239
rect 28549 6205 28583 6239
rect 28733 6205 28767 6239
rect 29285 6205 29319 6239
rect 30205 6205 30239 6239
rect 30297 6205 30331 6239
rect 30573 6205 30607 6239
rect 32413 6205 32447 6239
rect 34069 6205 34103 6239
rect 35265 6205 35299 6239
rect 35357 6205 35391 6239
rect 35633 6205 35667 6239
rect 23857 6137 23891 6171
rect 12541 6069 12575 6103
rect 17417 6069 17451 6103
rect 18153 6069 18187 6103
rect 29469 6069 29503 6103
rect 36737 6069 36771 6103
rect 2513 5865 2547 5899
rect 4169 5865 4203 5899
rect 10885 5865 10919 5899
rect 13921 5865 13955 5899
rect 15393 5865 15427 5899
rect 19717 5865 19751 5899
rect 24593 5865 24627 5899
rect 37841 5865 37875 5899
rect 39037 5865 39071 5899
rect 28089 5797 28123 5831
rect 30573 5797 30607 5831
rect 36185 5797 36219 5831
rect 2605 5729 2639 5763
rect 3157 5729 3191 5763
rect 3433 5729 3467 5763
rect 4077 5729 4111 5763
rect 4629 5729 4663 5763
rect 5365 5729 5399 5763
rect 8953 5729 8987 5763
rect 9873 5729 9907 5763
rect 9965 5729 9999 5763
rect 10333 5729 10367 5763
rect 10425 5729 10459 5763
rect 11989 5729 12023 5763
rect 13829 5729 13863 5763
rect 15301 5729 15335 5763
rect 16129 5729 16163 5763
rect 16221 5729 16255 5763
rect 16681 5729 16715 5763
rect 16865 5729 16899 5763
rect 17969 5729 18003 5763
rect 18521 5729 18555 5763
rect 18705 5729 18739 5763
rect 19625 5729 19659 5763
rect 20913 5729 20947 5763
rect 21281 5729 21315 5763
rect 21925 5729 21959 5763
rect 25145 5729 25179 5763
rect 27077 5729 27111 5763
rect 27353 5729 27387 5763
rect 28917 5729 28951 5763
rect 29561 5729 29595 5763
rect 31401 5729 31435 5763
rect 31585 5729 31619 5763
rect 32827 5729 32861 5763
rect 32965 5729 32999 5763
rect 34345 5729 34379 5763
rect 36737 5729 36771 5763
rect 37013 5729 37047 5763
rect 37841 5729 37875 5763
rect 38209 5729 38243 5763
rect 38945 5729 38979 5763
rect 5641 5661 5675 5695
rect 11713 5661 11747 5695
rect 13093 5661 13127 5695
rect 17233 5661 17267 5695
rect 17877 5661 17911 5695
rect 21005 5661 21039 5695
rect 23029 5661 23063 5695
rect 23305 5661 23339 5695
rect 26525 5661 26559 5695
rect 27537 5661 27571 5695
rect 28641 5661 28675 5695
rect 29101 5661 29135 5695
rect 31125 5661 31159 5695
rect 32137 5661 32171 5695
rect 32689 5661 32723 5695
rect 34069 5661 34103 5695
rect 37197 5661 37231 5695
rect 18889 5593 18923 5627
rect 25329 5593 25363 5627
rect 35449 5593 35483 5627
rect 6745 5525 6779 5559
rect 9045 5525 9079 5559
rect 29745 5525 29779 5559
rect 3065 5321 3099 5355
rect 9689 5321 9723 5355
rect 19901 5321 19935 5355
rect 23857 5321 23891 5355
rect 27261 5321 27295 5355
rect 28641 5321 28675 5355
rect 29469 5321 29503 5355
rect 31769 5321 31803 5355
rect 35173 5321 35207 5355
rect 37473 5321 37507 5355
rect 38301 5321 38335 5355
rect 11345 5253 11379 5287
rect 13737 5253 13771 5287
rect 1777 5185 1811 5219
rect 4721 5185 4755 5219
rect 8125 5185 8159 5219
rect 8401 5185 8435 5219
rect 18797 5185 18831 5219
rect 22385 5185 22419 5219
rect 24961 5185 24995 5219
rect 30389 5185 30423 5219
rect 33517 5185 33551 5219
rect 36093 5185 36127 5219
rect 36369 5185 36403 5219
rect 1501 5117 1535 5151
rect 4353 5117 4387 5151
rect 4629 5117 4663 5151
rect 5089 5117 5123 5151
rect 5733 5117 5767 5151
rect 5917 5117 5951 5151
rect 10425 5117 10459 5151
rect 10517 5117 10551 5151
rect 10885 5117 10919 5151
rect 10977 5117 11011 5151
rect 12633 5117 12667 5151
rect 12909 5117 12943 5151
rect 13737 5117 13771 5151
rect 14105 5117 14139 5151
rect 14657 5117 14691 5151
rect 15025 5117 15059 5151
rect 15577 5117 15611 5151
rect 16037 5117 16071 5151
rect 16221 5117 16255 5151
rect 16681 5117 16715 5151
rect 16773 5117 16807 5151
rect 18521 5117 18555 5151
rect 20637 5117 20671 5151
rect 22017 5117 22051 5151
rect 22109 5117 22143 5151
rect 22753 5117 22787 5151
rect 23673 5117 23707 5151
rect 25237 5117 25271 5151
rect 25421 5117 25455 5151
rect 25881 5117 25915 5151
rect 26157 5117 26191 5151
rect 28457 5117 28491 5151
rect 29285 5117 29319 5151
rect 30665 5117 30699 5151
rect 33057 5117 33091 5151
rect 33333 5117 33367 5151
rect 34897 5117 34931 5151
rect 34989 5117 35023 5151
rect 38209 5117 38243 5151
rect 38761 5117 38795 5151
rect 20729 5049 20763 5083
rect 24409 5049 24443 5083
rect 32505 5049 32539 5083
rect 6009 4981 6043 5015
rect 12725 4981 12759 5015
rect 17233 4981 17267 5015
rect 22845 4777 22879 4811
rect 29653 4777 29687 4811
rect 37013 4777 37047 4811
rect 11437 4709 11471 4743
rect 14657 4709 14691 4743
rect 20269 4709 20303 4743
rect 32137 4709 32171 4743
rect 4537 4641 4571 4675
rect 5181 4641 5215 4675
rect 10333 4641 10367 4675
rect 10425 4641 10459 4675
rect 10885 4641 10919 4675
rect 11069 4641 11103 4675
rect 12265 4641 12299 4675
rect 14197 4641 14231 4675
rect 15577 4641 15611 4675
rect 16589 4641 16623 4675
rect 18981 4641 19015 4675
rect 19441 4641 19475 4675
rect 20177 4641 20211 4675
rect 24409 4641 24443 4675
rect 24685 4641 24719 4675
rect 24869 4641 24903 4675
rect 27353 4641 27387 4675
rect 28089 4641 28123 4675
rect 30757 4641 30791 4675
rect 31033 4641 31067 4675
rect 32689 4641 32723 4675
rect 32965 4641 32999 4675
rect 34299 4641 34333 4675
rect 34437 4641 34471 4675
rect 35909 4641 35943 4675
rect 36093 4641 36127 4675
rect 36921 4641 36955 4675
rect 4905 4573 4939 4607
rect 6837 4573 6871 4607
rect 7113 4573 7147 4607
rect 11989 4573 12023 4607
rect 14105 4573 14139 4607
rect 16313 4573 16347 4607
rect 19717 4573 19751 4607
rect 21281 4573 21315 4607
rect 21557 4573 21591 4607
rect 23857 4573 23891 4607
rect 26525 4573 26559 4607
rect 27077 4573 27111 4607
rect 27537 4573 27571 4607
rect 28365 4573 28399 4607
rect 30205 4573 30239 4607
rect 31217 4573 31251 4607
rect 32827 4573 32861 4607
rect 33609 4573 33643 4607
rect 34161 4573 34195 4607
rect 35081 4573 35115 4607
rect 35633 4573 35667 4607
rect 15761 4505 15795 4539
rect 8217 4437 8251 4471
rect 13369 4437 13403 4471
rect 17877 4437 17911 4471
rect 18153 4165 18187 4199
rect 34253 4165 34287 4199
rect 4353 4097 4387 4131
rect 5089 4097 5123 4131
rect 6285 4097 6319 4131
rect 7481 4097 7515 4131
rect 14013 4097 14047 4131
rect 14289 4097 14323 4131
rect 15393 4097 15427 4131
rect 20269 4097 20303 4131
rect 23673 4097 23707 4131
rect 24225 4097 24259 4131
rect 25145 4097 25179 4131
rect 25697 4097 25731 4131
rect 26157 4097 26191 4131
rect 27169 4097 27203 4131
rect 27629 4097 27663 4131
rect 29561 4097 29595 4131
rect 30573 4097 30607 4131
rect 30849 4097 30883 4131
rect 34897 4097 34931 4131
rect 38945 4097 38979 4131
rect 4629 4029 4663 4063
rect 5549 4029 5583 4063
rect 5825 4029 5859 4063
rect 7573 4029 7607 4063
rect 8493 4029 8527 4063
rect 8769 4029 8803 4063
rect 11069 4029 11103 4063
rect 11253 4029 11287 4063
rect 12817 4029 12851 4063
rect 13369 4029 13403 4063
rect 16681 4029 16715 4063
rect 17049 4029 17083 4063
rect 18061 4029 18095 4063
rect 18797 4029 18831 4063
rect 19349 4029 19383 4063
rect 19993 4029 20027 4063
rect 22109 4029 22143 4063
rect 22201 4029 22235 4063
rect 24501 4029 24535 4063
rect 24685 4029 24719 4063
rect 25973 4029 26007 4063
rect 26617 4029 26651 4063
rect 27445 4029 27479 4063
rect 29469 4029 29503 4063
rect 33241 4029 33275 4063
rect 33517 4029 33551 4063
rect 33701 4029 33735 4063
rect 34161 4029 34195 4063
rect 35449 4029 35483 4063
rect 35725 4029 35759 4063
rect 35909 4029 35943 4063
rect 37473 4029 37507 4063
rect 37749 4029 37783 4063
rect 4537 3961 4571 3995
rect 5733 3961 5767 3995
rect 8033 3961 8067 3995
rect 10149 3961 10183 3995
rect 13553 3961 13587 3995
rect 19533 3961 19567 3995
rect 22661 3961 22695 3995
rect 32689 3961 32723 3995
rect 10885 3893 10919 3927
rect 16589 3893 16623 3927
rect 21557 3893 21591 3927
rect 32137 3893 32171 3927
rect 19809 3689 19843 3723
rect 29653 3689 29687 3723
rect 34529 3689 34563 3723
rect 10241 3621 10275 3655
rect 24685 3621 24719 3655
rect 7205 3553 7239 3587
rect 7481 3553 7515 3587
rect 8861 3553 8895 3587
rect 9781 3553 9815 3587
rect 10977 3553 11011 3587
rect 11345 3553 11379 3587
rect 15577 3553 15611 3587
rect 17877 3553 17911 3587
rect 19257 3553 19291 3587
rect 19717 3553 19751 3587
rect 23029 3553 23063 3587
rect 25145 3553 25179 3587
rect 27353 3553 27387 3587
rect 28089 3553 28123 3587
rect 28365 3553 28399 3587
rect 31033 3553 31067 3587
rect 32229 3553 32263 3587
rect 35817 3553 35851 3587
rect 9689 3485 9723 3519
rect 11253 3485 11287 3519
rect 12449 3485 12483 3519
rect 12725 3485 12759 3519
rect 15301 3485 15335 3519
rect 17601 3485 17635 3519
rect 20913 3485 20947 3519
rect 21189 3485 21223 3519
rect 23305 3485 23339 3519
rect 26525 3485 26559 3519
rect 27077 3485 27111 3519
rect 27537 3485 27571 3519
rect 30205 3485 30239 3519
rect 30757 3485 30791 3519
rect 31217 3485 31251 3519
rect 32965 3485 32999 3519
rect 33241 3485 33275 3519
rect 35541 3485 35575 3519
rect 25237 3417 25271 3451
rect 14013 3349 14047 3383
rect 16681 3349 16715 3383
rect 22477 3349 22511 3383
rect 32413 3349 32447 3383
rect 37105 3349 37139 3383
rect 14013 3145 14047 3179
rect 18337 3145 18371 3179
rect 25697 3145 25731 3179
rect 11805 3077 11839 3111
rect 36737 3077 36771 3111
rect 3433 3009 3467 3043
rect 9045 3009 9079 3043
rect 9781 3009 9815 3043
rect 12725 3009 12759 3043
rect 14841 3009 14875 3043
rect 15393 3009 15427 3043
rect 16129 3009 16163 3043
rect 18061 3009 18095 3043
rect 19809 3009 19843 3043
rect 24593 3009 24627 3043
rect 26709 3009 26743 3043
rect 29285 3009 29319 3043
rect 29837 3009 29871 3043
rect 31585 3009 31619 3043
rect 34897 3009 34931 3043
rect 37105 3009 37139 3043
rect 3157 2941 3191 2975
rect 7297 2941 7331 2975
rect 7389 2941 7423 2975
rect 8585 2941 8619 2975
rect 8861 2941 8895 2975
rect 9505 2941 9539 2975
rect 11713 2941 11747 2975
rect 12449 2941 12483 2975
rect 14933 2941 14967 2975
rect 15853 2941 15887 2975
rect 18153 2941 18187 2975
rect 19073 2941 19107 2975
rect 19533 2941 19567 2975
rect 20361 2941 20395 2975
rect 20637 2941 20671 2975
rect 22477 2941 22511 2975
rect 22569 2941 22603 2975
rect 24317 2941 24351 2975
rect 26433 2941 26467 2975
rect 29975 2941 30009 2975
rect 30113 2941 30147 2975
rect 31861 2941 31895 2975
rect 33701 2941 33735 2975
rect 35449 2941 35483 2975
rect 35725 2941 35759 2975
rect 35909 2941 35943 2975
rect 36737 2941 36771 2975
rect 36829 2941 36863 2975
rect 7849 2873 7883 2907
rect 17509 2873 17543 2907
rect 23029 2873 23063 2907
rect 33241 2873 33275 2907
rect 38485 2873 38519 2907
rect 4537 2805 4571 2839
rect 10885 2805 10919 2839
rect 21925 2805 21959 2839
rect 27813 2805 27847 2839
rect 33885 2805 33919 2839
rect 18889 2533 18923 2567
rect 22477 2533 22511 2567
rect 25145 2533 25179 2567
rect 32597 2533 32631 2567
rect 7205 2465 7239 2499
rect 7481 2465 7515 2499
rect 10701 2465 10735 2499
rect 12633 2465 12667 2499
rect 13093 2465 13127 2499
rect 14105 2465 14139 2499
rect 14565 2465 14599 2499
rect 15761 2465 15795 2499
rect 19717 2465 19751 2499
rect 21189 2465 21223 2499
rect 21925 2465 21959 2499
rect 23305 2465 23339 2499
rect 23489 2465 23523 2499
rect 24133 2465 24167 2499
rect 25697 2465 25731 2499
rect 25973 2465 26007 2499
rect 27445 2465 27479 2499
rect 27721 2465 27755 2499
rect 27905 2465 27939 2499
rect 28365 2465 28399 2499
rect 29745 2465 29779 2499
rect 30021 2465 30055 2499
rect 31493 2465 31527 2499
rect 33471 2465 33505 2499
rect 35449 2465 35483 2499
rect 35725 2465 35759 2499
rect 10425 2397 10459 2431
rect 13185 2397 13219 2431
rect 14013 2397 14047 2431
rect 15485 2397 15519 2431
rect 19441 2397 19475 2431
rect 19901 2397 19935 2431
rect 23029 2397 23063 2431
rect 24041 2397 24075 2431
rect 24593 2397 24627 2431
rect 26157 2397 26191 2431
rect 26893 2397 26927 2431
rect 33149 2397 33183 2431
rect 33609 2397 33643 2431
rect 21281 2329 21315 2363
rect 8585 2261 8619 2295
rect 11989 2261 12023 2295
rect 16865 2261 16899 2295
rect 28549 2261 28583 2295
rect 31309 2261 31343 2295
rect 37013 2261 37047 2295
<< metal1 >>
rect 1104 38650 39836 38672
rect 1104 38598 19606 38650
rect 19658 38598 19670 38650
rect 19722 38598 19734 38650
rect 19786 38598 19798 38650
rect 19850 38598 39836 38650
rect 1104 38576 39836 38598
rect 10502 38496 10508 38548
rect 10560 38536 10566 38548
rect 11333 38539 11391 38545
rect 11333 38536 11345 38539
rect 10560 38508 11345 38536
rect 10560 38496 10566 38508
rect 11333 38505 11345 38508
rect 11379 38505 11391 38539
rect 11333 38499 11391 38505
rect 14366 38496 14372 38548
rect 14424 38536 14430 38548
rect 17310 38536 17316 38548
rect 14424 38508 17316 38536
rect 14424 38496 14430 38508
rect 17310 38496 17316 38508
rect 17368 38496 17374 38548
rect 35894 38536 35900 38548
rect 29748 38508 35900 38536
rect 5994 38428 6000 38480
rect 6052 38468 6058 38480
rect 6052 38440 8616 38468
rect 6052 38428 6058 38440
rect 8294 38400 8300 38412
rect 8255 38372 8300 38400
rect 8294 38360 8300 38372
rect 8352 38360 8358 38412
rect 8588 38409 8616 38440
rect 8662 38428 8668 38480
rect 8720 38468 8726 38480
rect 9582 38468 9588 38480
rect 8720 38440 9588 38468
rect 8720 38428 8726 38440
rect 9582 38428 9588 38440
rect 9640 38428 9646 38480
rect 16574 38428 16580 38480
rect 16632 38468 16638 38480
rect 16632 38440 22048 38468
rect 16632 38428 16638 38440
rect 8573 38403 8631 38409
rect 8573 38369 8585 38403
rect 8619 38369 8631 38403
rect 8573 38363 8631 38369
rect 12805 38403 12863 38409
rect 12805 38369 12817 38403
rect 12851 38400 12863 38403
rect 12894 38400 12900 38412
rect 12851 38372 12900 38400
rect 12851 38369 12863 38372
rect 12805 38363 12863 38369
rect 12894 38360 12900 38372
rect 12952 38360 12958 38412
rect 14182 38400 14188 38412
rect 14143 38372 14188 38400
rect 14182 38360 14188 38372
rect 14240 38360 14246 38412
rect 14734 38400 14740 38412
rect 14695 38372 14740 38400
rect 14734 38360 14740 38372
rect 14792 38360 14798 38412
rect 19812 38409 19840 38440
rect 15473 38403 15531 38409
rect 15473 38369 15485 38403
rect 15519 38369 15531 38403
rect 15473 38363 15531 38369
rect 18785 38403 18843 38409
rect 18785 38369 18797 38403
rect 18831 38369 18843 38403
rect 18785 38363 18843 38369
rect 19705 38403 19763 38409
rect 19705 38369 19717 38403
rect 19751 38369 19763 38403
rect 19705 38363 19763 38369
rect 19797 38403 19855 38409
rect 19797 38369 19809 38403
rect 19843 38369 19855 38403
rect 19797 38363 19855 38369
rect 20441 38403 20499 38409
rect 20441 38369 20453 38403
rect 20487 38400 20499 38403
rect 20990 38400 20996 38412
rect 20487 38372 20996 38400
rect 20487 38369 20499 38372
rect 20441 38363 20499 38369
rect 8389 38335 8447 38341
rect 8389 38301 8401 38335
rect 8435 38332 8447 38335
rect 8662 38332 8668 38344
rect 8435 38304 8668 38332
rect 8435 38301 8447 38304
rect 8389 38295 8447 38301
rect 8662 38292 8668 38304
rect 8720 38292 8726 38344
rect 9306 38292 9312 38344
rect 9364 38332 9370 38344
rect 9953 38335 10011 38341
rect 9953 38332 9965 38335
rect 9364 38304 9965 38332
rect 9364 38292 9370 38304
rect 9953 38301 9965 38304
rect 9999 38301 10011 38335
rect 9953 38295 10011 38301
rect 10229 38335 10287 38341
rect 10229 38301 10241 38335
rect 10275 38332 10287 38335
rect 10870 38332 10876 38344
rect 10275 38304 10876 38332
rect 10275 38301 10287 38304
rect 10229 38295 10287 38301
rect 10870 38292 10876 38304
rect 10928 38292 10934 38344
rect 14553 38335 14611 38341
rect 14553 38301 14565 38335
rect 14599 38332 14611 38335
rect 15488 38332 15516 38363
rect 14599 38304 15516 38332
rect 18800 38332 18828 38363
rect 19521 38335 19579 38341
rect 19521 38332 19533 38335
rect 18800 38304 19533 38332
rect 14599 38301 14611 38304
rect 14553 38295 14611 38301
rect 19521 38301 19533 38304
rect 19567 38301 19579 38335
rect 19720 38332 19748 38363
rect 20990 38360 20996 38372
rect 21048 38360 21054 38412
rect 21542 38360 21548 38412
rect 21600 38400 21606 38412
rect 22020 38409 22048 38440
rect 26234 38428 26240 38480
rect 26292 38468 26298 38480
rect 26292 38440 28028 38468
rect 26292 38428 26298 38440
rect 21637 38403 21695 38409
rect 21637 38400 21649 38403
rect 21600 38372 21649 38400
rect 21600 38360 21606 38372
rect 21637 38369 21649 38372
rect 21683 38369 21695 38403
rect 21637 38363 21695 38369
rect 22005 38403 22063 38409
rect 22005 38369 22017 38403
rect 22051 38369 22063 38403
rect 22005 38363 22063 38369
rect 22278 38360 22284 38412
rect 22336 38400 22342 38412
rect 28000 38409 28028 38440
rect 22373 38403 22431 38409
rect 22373 38400 22385 38403
rect 22336 38372 22385 38400
rect 22336 38360 22342 38372
rect 22373 38369 22385 38372
rect 22419 38369 22431 38403
rect 22373 38363 22431 38369
rect 26329 38403 26387 38409
rect 26329 38369 26341 38403
rect 26375 38400 26387 38403
rect 26973 38403 27031 38409
rect 26973 38400 26985 38403
rect 26375 38372 26985 38400
rect 26375 38369 26387 38372
rect 26329 38363 26387 38369
rect 26973 38369 26985 38372
rect 27019 38369 27031 38403
rect 26973 38363 27031 38369
rect 27985 38403 28043 38409
rect 27985 38369 27997 38403
rect 28031 38369 28043 38403
rect 29748 38400 29776 38508
rect 35894 38496 35900 38508
rect 35952 38496 35958 38548
rect 29825 38403 29883 38409
rect 29825 38400 29837 38403
rect 29748 38372 29837 38400
rect 27985 38363 28043 38369
rect 29825 38369 29837 38372
rect 29871 38369 29883 38403
rect 29825 38363 29883 38369
rect 29914 38360 29920 38412
rect 29972 38400 29978 38412
rect 30837 38403 30895 38409
rect 30837 38400 30849 38403
rect 29972 38372 30849 38400
rect 29972 38360 29978 38372
rect 30837 38369 30849 38372
rect 30883 38369 30895 38403
rect 30837 38363 30895 38369
rect 20714 38332 20720 38344
rect 19720 38304 20720 38332
rect 19521 38295 19579 38301
rect 20714 38292 20720 38304
rect 20772 38292 20778 38344
rect 24673 38335 24731 38341
rect 24673 38301 24685 38335
rect 24719 38301 24731 38335
rect 24946 38332 24952 38344
rect 24907 38304 24952 38332
rect 24673 38295 24731 38301
rect 14090 38224 14096 38276
rect 14148 38264 14154 38276
rect 21818 38264 21824 38276
rect 14148 38236 21824 38264
rect 14148 38224 14154 38236
rect 21818 38224 21824 38236
rect 21876 38224 21882 38276
rect 12710 38156 12716 38208
rect 12768 38196 12774 38208
rect 12897 38199 12955 38205
rect 12897 38196 12909 38199
rect 12768 38168 12909 38196
rect 12768 38156 12774 38168
rect 12897 38165 12909 38168
rect 12943 38165 12955 38199
rect 15562 38196 15568 38208
rect 15523 38168 15568 38196
rect 12897 38159 12955 38165
rect 15562 38156 15568 38168
rect 15620 38156 15626 38208
rect 18877 38199 18935 38205
rect 18877 38165 18889 38199
rect 18923 38196 18935 38199
rect 20530 38196 20536 38208
rect 18923 38168 20536 38196
rect 18923 38165 18935 38168
rect 18877 38159 18935 38165
rect 20530 38156 20536 38168
rect 20588 38156 20594 38208
rect 21634 38156 21640 38208
rect 21692 38196 21698 38208
rect 21729 38199 21787 38205
rect 21729 38196 21741 38199
rect 21692 38168 21741 38196
rect 21692 38156 21698 38168
rect 21729 38165 21741 38168
rect 21775 38165 21787 38199
rect 24688 38196 24716 38295
rect 24946 38292 24952 38304
rect 25004 38292 25010 38344
rect 26881 38335 26939 38341
rect 26881 38301 26893 38335
rect 26927 38332 26939 38335
rect 27430 38332 27436 38344
rect 26927 38304 27436 38332
rect 26927 38301 26939 38304
rect 26881 38295 26939 38301
rect 27430 38292 27436 38304
rect 27488 38292 27494 38344
rect 27893 38335 27951 38341
rect 27893 38301 27905 38335
rect 27939 38332 27951 38335
rect 28626 38332 28632 38344
rect 27939 38304 28632 38332
rect 27939 38301 27951 38304
rect 27893 38295 27951 38301
rect 28626 38292 28632 38304
rect 28684 38332 28690 38344
rect 29733 38335 29791 38341
rect 29733 38332 29745 38335
rect 28684 38304 29745 38332
rect 28684 38292 28690 38304
rect 29733 38301 29745 38304
rect 29779 38332 29791 38335
rect 30745 38335 30803 38341
rect 30745 38332 30757 38335
rect 29779 38304 30757 38332
rect 29779 38301 29791 38304
rect 29733 38295 29791 38301
rect 30745 38301 30757 38304
rect 30791 38301 30803 38335
rect 30745 38295 30803 38301
rect 24854 38196 24860 38208
rect 24688 38168 24860 38196
rect 21729 38159 21787 38165
rect 24854 38156 24860 38168
rect 24912 38156 24918 38208
rect 26418 38156 26424 38208
rect 26476 38196 26482 38208
rect 27157 38199 27215 38205
rect 27157 38196 27169 38199
rect 26476 38168 27169 38196
rect 26476 38156 26482 38168
rect 27157 38165 27169 38168
rect 27203 38165 27215 38199
rect 27157 38159 27215 38165
rect 27614 38156 27620 38208
rect 27672 38196 27678 38208
rect 28169 38199 28227 38205
rect 28169 38196 28181 38199
rect 27672 38168 28181 38196
rect 27672 38156 27678 38168
rect 28169 38165 28181 38168
rect 28215 38165 28227 38199
rect 30006 38196 30012 38208
rect 29967 38168 30012 38196
rect 28169 38159 28227 38165
rect 30006 38156 30012 38168
rect 30064 38156 30070 38208
rect 31018 38196 31024 38208
rect 30979 38168 31024 38196
rect 31018 38156 31024 38168
rect 31076 38156 31082 38208
rect 1104 38106 39836 38128
rect 1104 38054 4246 38106
rect 4298 38054 4310 38106
rect 4362 38054 4374 38106
rect 4426 38054 4438 38106
rect 4490 38054 34966 38106
rect 35018 38054 35030 38106
rect 35082 38054 35094 38106
rect 35146 38054 35158 38106
rect 35210 38054 39836 38106
rect 1104 38032 39836 38054
rect 4614 37952 4620 38004
rect 4672 37992 4678 38004
rect 4985 37995 5043 38001
rect 4985 37992 4997 37995
rect 4672 37964 4997 37992
rect 4672 37952 4678 37964
rect 4985 37961 4997 37964
rect 5031 37961 5043 37995
rect 10870 37992 10876 38004
rect 10831 37964 10876 37992
rect 4985 37955 5043 37961
rect 10870 37952 10876 37964
rect 10928 37952 10934 38004
rect 12452 37964 15516 37992
rect 9674 37884 9680 37936
rect 9732 37924 9738 37936
rect 10045 37927 10103 37933
rect 10045 37924 10057 37927
rect 9732 37896 10057 37924
rect 9732 37884 9738 37896
rect 10045 37893 10057 37896
rect 10091 37924 10103 37927
rect 12342 37924 12348 37936
rect 10091 37896 12348 37924
rect 10091 37893 10103 37896
rect 10045 37887 10103 37893
rect 12342 37884 12348 37896
rect 12400 37884 12406 37936
rect 12452 37868 12480 37964
rect 3602 37856 3608 37868
rect 3515 37828 3608 37856
rect 3602 37816 3608 37828
rect 3660 37856 3666 37868
rect 5626 37856 5632 37868
rect 3660 37828 5632 37856
rect 3660 37816 3666 37828
rect 5626 37816 5632 37828
rect 5684 37816 5690 37868
rect 6638 37816 6644 37868
rect 6696 37856 6702 37868
rect 6825 37859 6883 37865
rect 6825 37856 6837 37859
rect 6696 37828 6837 37856
rect 6696 37816 6702 37828
rect 6825 37825 6837 37828
rect 6871 37825 6883 37859
rect 6825 37819 6883 37825
rect 7929 37859 7987 37865
rect 7929 37825 7941 37859
rect 7975 37856 7987 37859
rect 8757 37859 8815 37865
rect 8757 37856 8769 37859
rect 7975 37828 8769 37856
rect 7975 37825 7987 37828
rect 7929 37819 7987 37825
rect 8757 37825 8769 37828
rect 8803 37825 8815 37859
rect 12434 37856 12440 37868
rect 12347 37828 12440 37856
rect 8757 37819 8815 37825
rect 12434 37816 12440 37828
rect 12492 37816 12498 37868
rect 12710 37856 12716 37868
rect 12671 37828 12716 37856
rect 12710 37816 12716 37828
rect 12768 37816 12774 37868
rect 15488 37865 15516 37964
rect 16206 37952 16212 38004
rect 16264 37992 16270 38004
rect 16853 37995 16911 38001
rect 16853 37992 16865 37995
rect 16264 37964 16865 37992
rect 16264 37952 16270 37964
rect 16853 37961 16865 37964
rect 16899 37961 16911 37995
rect 16853 37955 16911 37961
rect 17218 37952 17224 38004
rect 17276 37992 17282 38004
rect 22094 37992 22100 38004
rect 17276 37964 22100 37992
rect 17276 37952 17282 37964
rect 22094 37952 22100 37964
rect 22152 37952 22158 38004
rect 24302 37992 24308 38004
rect 22572 37964 24308 37992
rect 15473 37859 15531 37865
rect 15473 37825 15485 37859
rect 15519 37856 15531 37859
rect 16206 37856 16212 37868
rect 15519 37828 16212 37856
rect 15519 37825 15531 37828
rect 15473 37819 15531 37825
rect 16206 37816 16212 37828
rect 16264 37816 16270 37868
rect 20257 37859 20315 37865
rect 20257 37825 20269 37859
rect 20303 37856 20315 37859
rect 22462 37856 22468 37868
rect 20303 37828 22468 37856
rect 20303 37825 20315 37828
rect 20257 37819 20315 37825
rect 22462 37816 22468 37828
rect 22520 37816 22526 37868
rect 22572 37865 22600 37964
rect 24302 37952 24308 37964
rect 24360 37952 24366 38004
rect 27798 37952 27804 38004
rect 27856 37992 27862 38004
rect 28445 37995 28503 38001
rect 28445 37992 28457 37995
rect 27856 37964 28457 37992
rect 27856 37952 27862 37964
rect 28445 37961 28457 37964
rect 28491 37961 28503 37995
rect 28445 37955 28503 37961
rect 31573 37995 31631 38001
rect 31573 37961 31585 37995
rect 31619 37992 31631 37995
rect 31662 37992 31668 38004
rect 31619 37964 31668 37992
rect 31619 37961 31631 37964
rect 31573 37955 31631 37961
rect 31662 37952 31668 37964
rect 31720 37952 31726 38004
rect 38841 37995 38899 38001
rect 38841 37961 38853 37995
rect 38887 37992 38899 37995
rect 39390 37992 39396 38004
rect 38887 37964 39396 37992
rect 38887 37961 38899 37964
rect 38841 37955 38899 37961
rect 39390 37952 39396 37964
rect 39448 37952 39454 38004
rect 22557 37859 22615 37865
rect 22557 37825 22569 37859
rect 22603 37825 22615 37859
rect 23937 37859 23995 37865
rect 23937 37856 23949 37859
rect 22557 37819 22615 37825
rect 23032 37828 23949 37856
rect 3881 37791 3939 37797
rect 3881 37757 3893 37791
rect 3927 37788 3939 37791
rect 3970 37788 3976 37800
rect 3927 37760 3976 37788
rect 3927 37757 3939 37760
rect 3881 37751 3939 37757
rect 3970 37748 3976 37760
rect 4028 37748 4034 37800
rect 7837 37791 7895 37797
rect 7837 37757 7849 37791
rect 7883 37788 7895 37791
rect 8386 37788 8392 37800
rect 7883 37760 8392 37788
rect 7883 37757 7895 37760
rect 7837 37751 7895 37757
rect 8386 37748 8392 37760
rect 8444 37748 8450 37800
rect 8481 37791 8539 37797
rect 8481 37757 8493 37791
rect 8527 37788 8539 37791
rect 9214 37788 9220 37800
rect 8527 37760 9220 37788
rect 8527 37757 8539 37760
rect 8481 37751 8539 37757
rect 9214 37748 9220 37760
rect 9272 37748 9278 37800
rect 10594 37788 10600 37800
rect 10555 37760 10600 37788
rect 10594 37748 10600 37760
rect 10652 37748 10658 37800
rect 10689 37791 10747 37797
rect 10689 37757 10701 37791
rect 10735 37788 10747 37791
rect 11054 37788 11060 37800
rect 10735 37760 11060 37788
rect 10735 37757 10747 37760
rect 10689 37751 10747 37757
rect 11054 37748 11060 37760
rect 11112 37748 11118 37800
rect 13814 37748 13820 37800
rect 13872 37788 13878 37800
rect 14093 37791 14151 37797
rect 14093 37788 14105 37791
rect 13872 37760 14105 37788
rect 13872 37748 13878 37760
rect 14093 37757 14105 37760
rect 14139 37788 14151 37791
rect 14553 37791 14611 37797
rect 14553 37788 14565 37791
rect 14139 37760 14565 37788
rect 14139 37757 14151 37760
rect 14093 37751 14151 37757
rect 14553 37757 14565 37760
rect 14599 37788 14611 37791
rect 15010 37788 15016 37800
rect 14599 37760 15016 37788
rect 14599 37757 14611 37760
rect 14553 37751 14611 37757
rect 15010 37748 15016 37760
rect 15068 37748 15074 37800
rect 15746 37788 15752 37800
rect 15707 37760 15752 37788
rect 15746 37748 15752 37760
rect 15804 37748 15810 37800
rect 18506 37748 18512 37800
rect 18564 37788 18570 37800
rect 18601 37791 18659 37797
rect 18601 37788 18613 37791
rect 18564 37760 18613 37788
rect 18564 37748 18570 37760
rect 18601 37757 18613 37760
rect 18647 37757 18659 37791
rect 18601 37751 18659 37757
rect 18690 37748 18696 37800
rect 18748 37788 18754 37800
rect 18969 37791 19027 37797
rect 18748 37760 18793 37788
rect 18748 37748 18754 37760
rect 18969 37757 18981 37791
rect 19015 37757 19027 37791
rect 19150 37788 19156 37800
rect 19111 37760 19156 37788
rect 18969 37751 19027 37757
rect 18984 37720 19012 37751
rect 19150 37748 19156 37760
rect 19208 37748 19214 37800
rect 19426 37788 19432 37800
rect 19387 37760 19432 37788
rect 19426 37748 19432 37760
rect 19484 37748 19490 37800
rect 20530 37788 20536 37800
rect 20491 37760 20536 37788
rect 20530 37748 20536 37760
rect 20588 37748 20594 37800
rect 22646 37788 22652 37800
rect 22607 37760 22652 37788
rect 22646 37748 22652 37760
rect 22704 37748 22710 37800
rect 19334 37720 19340 37732
rect 18984 37692 19340 37720
rect 19334 37680 19340 37692
rect 19392 37680 19398 37732
rect 21726 37680 21732 37732
rect 21784 37720 21790 37732
rect 23032 37720 23060 37828
rect 23937 37825 23949 37828
rect 23983 37825 23995 37859
rect 26418 37856 26424 37868
rect 23937 37819 23995 37825
rect 24780 37828 26280 37856
rect 26379 37828 26424 37856
rect 23382 37748 23388 37800
rect 23440 37788 23446 37800
rect 23661 37791 23719 37797
rect 23661 37788 23673 37791
rect 23440 37760 23673 37788
rect 23440 37748 23446 37760
rect 23661 37757 23673 37760
rect 23707 37788 23719 37791
rect 24780 37788 24808 37828
rect 23707 37760 24808 37788
rect 23707 37757 23719 37760
rect 23661 37751 23719 37757
rect 24854 37748 24860 37800
rect 24912 37788 24918 37800
rect 25774 37788 25780 37800
rect 24912 37760 25780 37788
rect 24912 37748 24918 37760
rect 25774 37748 25780 37760
rect 25832 37788 25838 37800
rect 26145 37791 26203 37797
rect 26145 37788 26157 37791
rect 25832 37760 26157 37788
rect 25832 37748 25838 37760
rect 26145 37757 26157 37760
rect 26191 37757 26203 37791
rect 26252 37788 26280 37828
rect 26418 37816 26424 37828
rect 26476 37816 26482 37868
rect 28994 37816 29000 37868
rect 29052 37856 29058 37868
rect 33597 37859 33655 37865
rect 33597 37856 33609 37859
rect 29052 37828 33609 37856
rect 29052 37816 29058 37828
rect 33597 37825 33609 37828
rect 33643 37825 33655 37859
rect 33597 37819 33655 37825
rect 26252 37760 27108 37788
rect 26145 37751 26203 37757
rect 21784 37692 23060 37720
rect 23109 37723 23167 37729
rect 21784 37680 21790 37692
rect 23109 37689 23121 37723
rect 23155 37720 23167 37723
rect 23750 37720 23756 37732
rect 23155 37692 23756 37720
rect 23155 37689 23167 37692
rect 23109 37683 23167 37689
rect 23750 37680 23756 37692
rect 23808 37680 23814 37732
rect 27080 37720 27108 37760
rect 28074 37748 28080 37800
rect 28132 37788 28138 37800
rect 28261 37791 28319 37797
rect 28261 37788 28273 37791
rect 28132 37760 28273 37788
rect 28132 37748 28138 37760
rect 28261 37757 28273 37760
rect 28307 37757 28319 37791
rect 28261 37751 28319 37757
rect 30009 37791 30067 37797
rect 30009 37757 30021 37791
rect 30055 37757 30067 37791
rect 30009 37751 30067 37757
rect 30024 37720 30052 37751
rect 30098 37748 30104 37800
rect 30156 37788 30162 37800
rect 30285 37791 30343 37797
rect 30285 37788 30297 37791
rect 30156 37760 30297 37788
rect 30156 37748 30162 37760
rect 30285 37757 30297 37760
rect 30331 37757 30343 37791
rect 30285 37751 30343 37757
rect 32030 37748 32036 37800
rect 32088 37788 32094 37800
rect 32217 37791 32275 37797
rect 32217 37788 32229 37791
rect 32088 37760 32229 37788
rect 32088 37748 32094 37760
rect 32217 37757 32229 37760
rect 32263 37757 32275 37791
rect 32217 37751 32275 37757
rect 32493 37791 32551 37797
rect 32493 37757 32505 37791
rect 32539 37788 32551 37791
rect 32766 37788 32772 37800
rect 32539 37760 32772 37788
rect 32539 37757 32551 37760
rect 32493 37751 32551 37757
rect 32766 37748 32772 37760
rect 32824 37748 32830 37800
rect 38657 37791 38715 37797
rect 38657 37788 38669 37791
rect 38488 37760 38669 37788
rect 27080 37692 30144 37720
rect 14645 37655 14703 37661
rect 14645 37621 14657 37655
rect 14691 37652 14703 37655
rect 14918 37652 14924 37664
rect 14691 37624 14924 37652
rect 14691 37621 14703 37624
rect 14645 37615 14703 37621
rect 14918 37612 14924 37624
rect 14976 37612 14982 37664
rect 18141 37655 18199 37661
rect 18141 37621 18153 37655
rect 18187 37652 18199 37655
rect 18874 37652 18880 37664
rect 18187 37624 18880 37652
rect 18187 37621 18199 37624
rect 18141 37615 18199 37621
rect 18874 37612 18880 37624
rect 18932 37612 18938 37664
rect 21174 37612 21180 37664
rect 21232 37652 21238 37664
rect 21637 37655 21695 37661
rect 21637 37652 21649 37655
rect 21232 37624 21649 37652
rect 21232 37612 21238 37624
rect 21637 37621 21649 37624
rect 21683 37621 21695 37655
rect 21637 37615 21695 37621
rect 22462 37612 22468 37664
rect 22520 37652 22526 37664
rect 23382 37652 23388 37664
rect 22520 37624 23388 37652
rect 22520 37612 22526 37624
rect 23382 37612 23388 37624
rect 23440 37612 23446 37664
rect 23474 37612 23480 37664
rect 23532 37652 23538 37664
rect 25041 37655 25099 37661
rect 25041 37652 25053 37655
rect 23532 37624 25053 37652
rect 23532 37612 23538 37624
rect 25041 37621 25053 37624
rect 25087 37621 25099 37655
rect 27522 37652 27528 37664
rect 27483 37624 27528 37652
rect 25041 37615 25099 37621
rect 27522 37612 27528 37624
rect 27580 37612 27586 37664
rect 29822 37652 29828 37664
rect 29783 37624 29828 37652
rect 29822 37612 29828 37624
rect 29880 37612 29886 37664
rect 30116 37652 30144 37692
rect 32122 37652 32128 37664
rect 30116 37624 32128 37652
rect 32122 37612 32128 37624
rect 32180 37612 32186 37664
rect 38286 37612 38292 37664
rect 38344 37652 38350 37664
rect 38488 37661 38516 37760
rect 38657 37757 38669 37760
rect 38703 37757 38715 37791
rect 38657 37751 38715 37757
rect 38473 37655 38531 37661
rect 38473 37652 38485 37655
rect 38344 37624 38485 37652
rect 38344 37612 38350 37624
rect 38473 37621 38485 37624
rect 38519 37621 38531 37655
rect 38473 37615 38531 37621
rect 1104 37562 39836 37584
rect 1104 37510 19606 37562
rect 19658 37510 19670 37562
rect 19722 37510 19734 37562
rect 19786 37510 19798 37562
rect 19850 37510 39836 37562
rect 1104 37488 39836 37510
rect 7650 37448 7656 37460
rect 4632 37420 7656 37448
rect 4632 37389 4660 37420
rect 7650 37408 7656 37420
rect 7708 37408 7714 37460
rect 8294 37408 8300 37460
rect 8352 37448 8358 37460
rect 9769 37451 9827 37457
rect 9769 37448 9781 37451
rect 8352 37420 9781 37448
rect 8352 37408 8358 37420
rect 9769 37417 9781 37420
rect 9815 37417 9827 37451
rect 11885 37451 11943 37457
rect 9769 37411 9827 37417
rect 10428 37420 11284 37448
rect 4617 37383 4675 37389
rect 4617 37349 4629 37383
rect 4663 37349 4675 37383
rect 10134 37380 10140 37392
rect 4617 37343 4675 37349
rect 8496 37352 10140 37380
rect 4709 37315 4767 37321
rect 4709 37281 4721 37315
rect 4755 37312 4767 37315
rect 5169 37315 5227 37321
rect 4755 37284 5028 37312
rect 4755 37281 4767 37284
rect 4709 37275 4767 37281
rect 5000 37176 5028 37284
rect 5169 37281 5181 37315
rect 5215 37312 5227 37315
rect 5905 37315 5963 37321
rect 5905 37312 5917 37315
rect 5215 37284 5917 37312
rect 5215 37281 5227 37284
rect 5169 37275 5227 37281
rect 5905 37281 5917 37284
rect 5951 37281 5963 37315
rect 8110 37312 8116 37324
rect 8071 37284 8116 37312
rect 5905 37275 5963 37281
rect 8110 37272 8116 37284
rect 8168 37272 8174 37324
rect 8496 37321 8524 37352
rect 10134 37340 10140 37352
rect 10192 37380 10198 37392
rect 10428 37380 10456 37420
rect 10192 37352 10456 37380
rect 11256 37380 11284 37420
rect 11885 37417 11897 37451
rect 11931 37448 11943 37451
rect 17218 37448 17224 37460
rect 11931 37420 17224 37448
rect 11931 37417 11943 37420
rect 11885 37411 11943 37417
rect 17218 37408 17224 37420
rect 17276 37408 17282 37460
rect 18782 37448 18788 37460
rect 18743 37420 18788 37448
rect 18782 37408 18788 37420
rect 18840 37408 18846 37460
rect 20990 37448 20996 37460
rect 20951 37420 20996 37448
rect 20990 37408 20996 37420
rect 21048 37408 21054 37460
rect 21726 37448 21732 37460
rect 21687 37420 21732 37448
rect 21726 37408 21732 37420
rect 21784 37408 21790 37460
rect 21818 37408 21824 37460
rect 21876 37448 21882 37460
rect 29822 37448 29828 37460
rect 21876 37420 29828 37448
rect 21876 37408 21882 37420
rect 29822 37408 29828 37420
rect 29880 37448 29886 37460
rect 30098 37448 30104 37460
rect 29880 37420 30104 37448
rect 29880 37408 29886 37420
rect 30098 37408 30104 37420
rect 30156 37408 30162 37460
rect 33686 37448 33692 37460
rect 33647 37420 33692 37448
rect 33686 37408 33692 37420
rect 33744 37408 33750 37460
rect 35526 37408 35532 37460
rect 35584 37448 35590 37460
rect 35621 37451 35679 37457
rect 35621 37448 35633 37451
rect 35584 37420 35633 37448
rect 35584 37408 35590 37420
rect 35621 37417 35633 37420
rect 35667 37417 35679 37451
rect 35621 37411 35679 37417
rect 12802 37380 12808 37392
rect 11256 37352 12808 37380
rect 10192 37340 10198 37352
rect 12802 37340 12808 37352
rect 12860 37340 12866 37392
rect 12986 37340 12992 37392
rect 13044 37380 13050 37392
rect 17865 37383 17923 37389
rect 13044 37352 14412 37380
rect 13044 37340 13050 37352
rect 8481 37315 8539 37321
rect 8481 37281 8493 37315
rect 8527 37281 8539 37315
rect 8662 37312 8668 37324
rect 8623 37284 8668 37312
rect 8481 37275 8539 37281
rect 8662 37272 8668 37284
rect 8720 37272 8726 37324
rect 9674 37312 9680 37324
rect 9635 37284 9680 37312
rect 9674 37272 9680 37284
rect 9732 37272 9738 37324
rect 10597 37315 10655 37321
rect 10597 37281 10609 37315
rect 10643 37312 10655 37315
rect 10686 37312 10692 37324
rect 10643 37284 10692 37312
rect 10643 37281 10655 37284
rect 10597 37275 10655 37281
rect 10686 37272 10692 37284
rect 10744 37272 10750 37324
rect 12897 37315 12955 37321
rect 12897 37281 12909 37315
rect 12943 37312 12955 37315
rect 13078 37312 13084 37324
rect 12943 37284 13084 37312
rect 12943 37281 12955 37284
rect 12897 37275 12955 37281
rect 13078 37272 13084 37284
rect 13136 37272 13142 37324
rect 13814 37312 13820 37324
rect 13775 37284 13820 37312
rect 13814 37272 13820 37284
rect 13872 37272 13878 37324
rect 14093 37315 14151 37321
rect 14093 37281 14105 37315
rect 14139 37312 14151 37315
rect 14139 37284 14320 37312
rect 14139 37281 14151 37284
rect 14093 37275 14151 37281
rect 5626 37244 5632 37256
rect 5587 37216 5632 37244
rect 5626 37204 5632 37216
rect 5684 37204 5690 37256
rect 8386 37244 8392 37256
rect 8347 37216 8392 37244
rect 8386 37204 8392 37216
rect 8444 37204 8450 37256
rect 10321 37247 10379 37253
rect 10321 37213 10333 37247
rect 10367 37244 10379 37247
rect 12434 37244 12440 37256
rect 10367 37216 12440 37244
rect 10367 37213 10379 37216
rect 10321 37207 10379 37213
rect 12434 37204 12440 37216
rect 12492 37204 12498 37256
rect 14182 37244 14188 37256
rect 14143 37216 14188 37244
rect 14182 37204 14188 37216
rect 14240 37204 14246 37256
rect 5000 37148 5580 37176
rect 4433 37111 4491 37117
rect 4433 37077 4445 37111
rect 4479 37108 4491 37111
rect 4798 37108 4804 37120
rect 4479 37080 4804 37108
rect 4479 37077 4491 37080
rect 4433 37071 4491 37077
rect 4798 37068 4804 37080
rect 4856 37068 4862 37120
rect 5552 37108 5580 37148
rect 9582 37136 9588 37188
rect 9640 37136 9646 37188
rect 14292 37176 14320 37284
rect 14384 37244 14412 37352
rect 14476 37352 15608 37380
rect 14476 37321 14504 37352
rect 15580 37321 15608 37352
rect 17865 37349 17877 37383
rect 17911 37380 17923 37383
rect 18230 37380 18236 37392
rect 17911 37352 18236 37380
rect 17911 37349 17923 37352
rect 17865 37343 17923 37349
rect 18230 37340 18236 37352
rect 18288 37340 18294 37392
rect 19334 37340 19340 37392
rect 19392 37380 19398 37392
rect 22278 37380 22284 37392
rect 19392 37352 19564 37380
rect 22239 37352 22284 37380
rect 19392 37340 19398 37352
rect 14461 37315 14519 37321
rect 14461 37281 14473 37315
rect 14507 37281 14519 37315
rect 14461 37275 14519 37281
rect 15473 37315 15531 37321
rect 15473 37281 15485 37315
rect 15519 37281 15531 37315
rect 15473 37275 15531 37281
rect 15565 37315 15623 37321
rect 15565 37281 15577 37315
rect 15611 37312 15623 37315
rect 15838 37312 15844 37324
rect 15611 37284 15844 37312
rect 15611 37281 15623 37284
rect 15565 37275 15623 37281
rect 15488 37244 15516 37275
rect 15838 37272 15844 37284
rect 15896 37272 15902 37324
rect 16482 37312 16488 37324
rect 15948 37284 16344 37312
rect 16443 37284 16488 37312
rect 15948 37244 15976 37284
rect 16206 37244 16212 37256
rect 14384 37216 15976 37244
rect 16167 37216 16212 37244
rect 16206 37204 16212 37216
rect 16264 37204 16270 37256
rect 16316 37244 16344 37284
rect 16482 37272 16488 37284
rect 16540 37272 16546 37324
rect 18506 37312 18512 37324
rect 18467 37284 18512 37312
rect 18506 37272 18512 37284
rect 18564 37272 18570 37324
rect 19536 37321 19564 37352
rect 22278 37340 22284 37352
rect 22336 37340 22342 37392
rect 19153 37315 19211 37321
rect 19153 37281 19165 37315
rect 19199 37281 19211 37315
rect 19153 37275 19211 37281
rect 19521 37315 19579 37321
rect 19521 37281 19533 37315
rect 19567 37281 19579 37315
rect 19886 37312 19892 37324
rect 19847 37284 19892 37312
rect 19521 37275 19579 37281
rect 18690 37244 18696 37256
rect 16316 37216 18696 37244
rect 18690 37204 18696 37216
rect 18748 37204 18754 37256
rect 19168 37244 19196 37275
rect 19886 37272 19892 37284
rect 19944 37272 19950 37324
rect 20898 37312 20904 37324
rect 20859 37284 20904 37312
rect 20898 37272 20904 37284
rect 20956 37272 20962 37324
rect 21634 37312 21640 37324
rect 21595 37284 21640 37312
rect 21634 37272 21640 37284
rect 21692 37272 21698 37324
rect 22833 37315 22891 37321
rect 22833 37281 22845 37315
rect 22879 37281 22891 37315
rect 22833 37275 22891 37281
rect 19426 37244 19432 37256
rect 19168 37216 19432 37244
rect 19426 37204 19432 37216
rect 19484 37204 19490 37256
rect 21910 37204 21916 37256
rect 21968 37244 21974 37256
rect 22848 37244 22876 37275
rect 22922 37272 22928 37324
rect 22980 37312 22986 37324
rect 23198 37312 23204 37324
rect 22980 37284 23025 37312
rect 23159 37284 23204 37312
rect 22980 37272 22986 37284
rect 23198 37272 23204 37284
rect 23256 37272 23262 37324
rect 23382 37312 23388 37324
rect 23343 37284 23388 37312
rect 23382 37272 23388 37284
rect 23440 37272 23446 37324
rect 23566 37312 23572 37324
rect 23527 37284 23572 37312
rect 23566 37272 23572 37284
rect 23624 37272 23630 37324
rect 23750 37272 23756 37324
rect 23808 37312 23814 37324
rect 24581 37315 24639 37321
rect 24581 37312 24593 37315
rect 23808 37284 24593 37312
rect 23808 37272 23814 37284
rect 24581 37281 24593 37284
rect 24627 37281 24639 37315
rect 24854 37312 24860 37324
rect 24581 37275 24639 37281
rect 24688 37284 24860 37312
rect 23474 37244 23480 37256
rect 21968 37216 22784 37244
rect 22848 37216 23480 37244
rect 21968 37204 21974 37216
rect 15102 37176 15108 37188
rect 12912 37148 13308 37176
rect 14292 37148 15108 37176
rect 5994 37108 6000 37120
rect 5552 37080 6000 37108
rect 5994 37068 6000 37080
rect 6052 37068 6058 37120
rect 7190 37108 7196 37120
rect 7151 37080 7196 37108
rect 7190 37068 7196 37080
rect 7248 37068 7254 37120
rect 9600 37108 9628 37136
rect 12912 37108 12940 37148
rect 9600 37080 12940 37108
rect 12989 37111 13047 37117
rect 12989 37077 13001 37111
rect 13035 37108 13047 37111
rect 13170 37108 13176 37120
rect 13035 37080 13176 37108
rect 13035 37077 13047 37080
rect 12989 37071 13047 37077
rect 13170 37068 13176 37080
rect 13228 37068 13234 37120
rect 13280 37108 13308 37148
rect 15102 37136 15108 37148
rect 15160 37136 15166 37188
rect 17310 37136 17316 37188
rect 17368 37176 17374 37188
rect 22646 37176 22652 37188
rect 17368 37148 22652 37176
rect 17368 37136 17374 37148
rect 22646 37136 22652 37148
rect 22704 37136 22710 37188
rect 22756 37176 22784 37216
rect 23474 37204 23480 37216
rect 23532 37204 23538 37256
rect 24305 37247 24363 37253
rect 24305 37213 24317 37247
rect 24351 37244 24363 37247
rect 24688 37244 24716 37284
rect 24854 37272 24860 37284
rect 24912 37272 24918 37324
rect 25961 37315 26019 37321
rect 25961 37281 25973 37315
rect 26007 37312 26019 37315
rect 26602 37312 26608 37324
rect 26007 37284 26608 37312
rect 26007 37281 26019 37284
rect 25961 37275 26019 37281
rect 26602 37272 26608 37284
rect 26660 37272 26666 37324
rect 27614 37312 27620 37324
rect 27575 37284 27620 37312
rect 27614 37272 27620 37284
rect 27672 37272 27678 37324
rect 29270 37312 29276 37324
rect 27724 37284 29276 37312
rect 24351 37216 24716 37244
rect 24351 37213 24363 37216
rect 24305 37207 24363 37213
rect 25774 37204 25780 37256
rect 25832 37244 25838 37256
rect 27341 37247 27399 37253
rect 27341 37244 27353 37247
rect 25832 37216 27353 37244
rect 25832 37204 25838 37216
rect 27341 37213 27353 37216
rect 27387 37244 27399 37247
rect 27724 37244 27752 37284
rect 29270 37272 29276 37284
rect 29328 37312 29334 37324
rect 29457 37315 29515 37321
rect 29457 37312 29469 37315
rect 29328 37284 29469 37312
rect 29328 37272 29334 37284
rect 29457 37281 29469 37284
rect 29503 37281 29515 37315
rect 29457 37275 29515 37281
rect 29733 37315 29791 37321
rect 29733 37281 29745 37315
rect 29779 37312 29791 37315
rect 31018 37312 31024 37324
rect 29779 37284 31024 37312
rect 29779 37281 29791 37284
rect 29733 37275 29791 37281
rect 31018 37272 31024 37284
rect 31076 37272 31082 37324
rect 31113 37315 31171 37321
rect 31113 37281 31125 37315
rect 31159 37312 31171 37315
rect 31938 37312 31944 37324
rect 31159 37284 31944 37312
rect 31159 37281 31171 37284
rect 31113 37275 31171 37281
rect 31938 37272 31944 37284
rect 31996 37272 32002 37324
rect 32122 37312 32128 37324
rect 32035 37284 32128 37312
rect 32122 37272 32128 37284
rect 32180 37312 32186 37324
rect 34241 37315 34299 37321
rect 34241 37312 34253 37315
rect 32180 37284 34253 37312
rect 32180 37272 32186 37284
rect 34241 37281 34253 37284
rect 34287 37281 34299 37315
rect 34241 37275 34299 37281
rect 34517 37315 34575 37321
rect 34517 37281 34529 37315
rect 34563 37312 34575 37315
rect 35526 37312 35532 37324
rect 34563 37284 35532 37312
rect 34563 37281 34575 37284
rect 34517 37275 34575 37281
rect 35526 37272 35532 37284
rect 35584 37272 35590 37324
rect 27387 37216 27752 37244
rect 27387 37213 27399 37216
rect 27341 37207 27399 37213
rect 31846 37204 31852 37256
rect 31904 37244 31910 37256
rect 32401 37247 32459 37253
rect 32401 37244 32413 37247
rect 31904 37216 32413 37244
rect 31904 37204 31910 37216
rect 32401 37213 32413 37216
rect 32447 37213 32459 37247
rect 32401 37207 32459 37213
rect 23198 37176 23204 37188
rect 22756 37148 23204 37176
rect 23198 37136 23204 37148
rect 23256 37136 23262 37188
rect 27982 37108 27988 37120
rect 13280 37080 27988 37108
rect 27982 37068 27988 37080
rect 28040 37068 28046 37120
rect 28718 37108 28724 37120
rect 28679 37080 28724 37108
rect 28718 37068 28724 37080
rect 28776 37068 28782 37120
rect 1104 37018 39836 37040
rect 1104 36966 4246 37018
rect 4298 36966 4310 37018
rect 4362 36966 4374 37018
rect 4426 36966 4438 37018
rect 4490 36966 34966 37018
rect 35018 36966 35030 37018
rect 35082 36966 35094 37018
rect 35146 36966 35158 37018
rect 35210 36966 39836 37018
rect 1104 36944 39836 36966
rect 2774 36864 2780 36916
rect 2832 36904 2838 36916
rect 2832 36876 2877 36904
rect 2832 36864 2838 36876
rect 2958 36864 2964 36916
rect 3016 36904 3022 36916
rect 11146 36904 11152 36916
rect 3016 36876 11152 36904
rect 3016 36864 3022 36876
rect 11146 36864 11152 36876
rect 11204 36864 11210 36916
rect 16206 36904 16212 36916
rect 14660 36876 16212 36904
rect 9674 36836 9680 36848
rect 5552 36808 7052 36836
rect 1397 36771 1455 36777
rect 1397 36737 1409 36771
rect 1443 36768 1455 36771
rect 3602 36768 3608 36780
rect 1443 36740 3608 36768
rect 1443 36737 1455 36740
rect 1397 36731 1455 36737
rect 3602 36728 3608 36740
rect 3660 36728 3666 36780
rect 4798 36768 4804 36780
rect 4759 36740 4804 36768
rect 4798 36728 4804 36740
rect 4856 36728 4862 36780
rect 1673 36703 1731 36709
rect 1673 36669 1685 36703
rect 1719 36700 1731 36703
rect 1946 36700 1952 36712
rect 1719 36672 1952 36700
rect 1719 36669 1731 36672
rect 1673 36663 1731 36669
rect 1946 36660 1952 36672
rect 2004 36660 2010 36712
rect 5350 36700 5356 36712
rect 5311 36672 5356 36700
rect 5350 36660 5356 36672
rect 5408 36660 5414 36712
rect 5552 36709 5580 36808
rect 6454 36768 6460 36780
rect 5736 36740 6460 36768
rect 5736 36709 5764 36740
rect 6454 36728 6460 36740
rect 6512 36728 6518 36780
rect 5537 36703 5595 36709
rect 5537 36669 5549 36703
rect 5583 36669 5595 36703
rect 5537 36663 5595 36669
rect 5721 36703 5779 36709
rect 5721 36669 5733 36703
rect 5767 36669 5779 36703
rect 5721 36663 5779 36669
rect 5905 36703 5963 36709
rect 5905 36669 5917 36703
rect 5951 36669 5963 36703
rect 5905 36663 5963 36669
rect 6181 36703 6239 36709
rect 6181 36669 6193 36703
rect 6227 36700 6239 36703
rect 6914 36700 6920 36712
rect 6227 36672 6920 36700
rect 6227 36669 6239 36672
rect 6181 36663 6239 36669
rect 5920 36564 5948 36663
rect 6914 36660 6920 36672
rect 6972 36660 6978 36712
rect 7024 36632 7052 36808
rect 7116 36808 9680 36836
rect 7116 36709 7144 36808
rect 9674 36796 9680 36808
rect 9732 36796 9738 36848
rect 7282 36728 7288 36780
rect 7340 36768 7346 36780
rect 8110 36768 8116 36780
rect 7340 36740 7972 36768
rect 8071 36740 8116 36768
rect 7340 36728 7346 36740
rect 7101 36703 7159 36709
rect 7101 36669 7113 36703
rect 7147 36669 7159 36703
rect 7101 36663 7159 36669
rect 7190 36660 7196 36712
rect 7248 36700 7254 36712
rect 7469 36703 7527 36709
rect 7469 36700 7481 36703
rect 7248 36672 7481 36700
rect 7248 36660 7254 36672
rect 7469 36669 7481 36672
rect 7515 36669 7527 36703
rect 7834 36700 7840 36712
rect 7795 36672 7840 36700
rect 7469 36663 7527 36669
rect 7834 36660 7840 36672
rect 7892 36660 7898 36712
rect 7944 36700 7972 36740
rect 8110 36728 8116 36740
rect 8168 36728 8174 36780
rect 11517 36771 11575 36777
rect 11517 36737 11529 36771
rect 11563 36768 11575 36771
rect 11563 36740 12480 36768
rect 11563 36737 11575 36740
rect 11517 36731 11575 36737
rect 8389 36703 8447 36709
rect 8389 36700 8401 36703
rect 7944 36672 8401 36700
rect 8389 36669 8401 36672
rect 8435 36669 8447 36703
rect 8389 36663 8447 36669
rect 9861 36703 9919 36709
rect 9861 36669 9873 36703
rect 9907 36700 9919 36703
rect 10137 36703 10195 36709
rect 9907 36672 10088 36700
rect 9907 36669 9919 36672
rect 9861 36663 9919 36669
rect 8570 36632 8576 36644
rect 7024 36604 8576 36632
rect 8570 36592 8576 36604
rect 8628 36592 8634 36644
rect 7374 36564 7380 36576
rect 5920 36536 7380 36564
rect 7374 36524 7380 36536
rect 7432 36524 7438 36576
rect 9861 36567 9919 36573
rect 9861 36533 9873 36567
rect 9907 36564 9919 36567
rect 9950 36564 9956 36576
rect 9907 36536 9956 36564
rect 9907 36533 9919 36536
rect 9861 36527 9919 36533
rect 9950 36524 9956 36536
rect 10008 36524 10014 36576
rect 10060 36564 10088 36672
rect 10137 36669 10149 36703
rect 10183 36700 10195 36703
rect 10318 36700 10324 36712
rect 10183 36672 10324 36700
rect 10183 36669 10195 36672
rect 10137 36663 10195 36669
rect 10318 36660 10324 36672
rect 10376 36660 10382 36712
rect 11422 36700 11428 36712
rect 11383 36672 11428 36700
rect 11422 36660 11428 36672
rect 11480 36660 11486 36712
rect 12452 36709 12480 36740
rect 12894 36728 12900 36780
rect 12952 36768 12958 36780
rect 14660 36777 14688 36876
rect 16206 36864 16212 36876
rect 16264 36864 16270 36916
rect 18782 36864 18788 36916
rect 18840 36904 18846 36916
rect 21542 36904 21548 36916
rect 18840 36876 21404 36904
rect 21503 36876 21548 36904
rect 18840 36864 18846 36876
rect 16298 36796 16304 36848
rect 16356 36836 16362 36848
rect 16853 36839 16911 36845
rect 16853 36836 16865 36839
rect 16356 36808 16865 36836
rect 16356 36796 16362 36808
rect 16853 36805 16865 36808
rect 16899 36805 16911 36839
rect 16853 36799 16911 36805
rect 19886 36796 19892 36848
rect 19944 36836 19950 36848
rect 21266 36836 21272 36848
rect 19944 36808 21272 36836
rect 19944 36796 19950 36808
rect 21266 36796 21272 36808
rect 21324 36796 21330 36848
rect 21376 36836 21404 36876
rect 21542 36864 21548 36876
rect 21600 36864 21606 36916
rect 24581 36907 24639 36913
rect 24581 36873 24593 36907
rect 24627 36904 24639 36907
rect 24946 36904 24952 36916
rect 24627 36876 24952 36904
rect 24627 36873 24639 36876
rect 24581 36867 24639 36873
rect 24946 36864 24952 36876
rect 25004 36864 25010 36916
rect 27798 36864 27804 36916
rect 27856 36904 27862 36916
rect 28445 36907 28503 36913
rect 28445 36904 28457 36907
rect 27856 36876 28457 36904
rect 27856 36864 27862 36876
rect 28445 36873 28457 36876
rect 28491 36873 28503 36907
rect 32766 36904 32772 36916
rect 32727 36876 32772 36904
rect 28445 36867 28503 36873
rect 32766 36864 32772 36876
rect 32824 36864 32830 36916
rect 21376 36808 22324 36836
rect 14645 36771 14703 36777
rect 12952 36740 12997 36768
rect 12952 36728 12958 36740
rect 14645 36737 14657 36771
rect 14691 36737 14703 36771
rect 14645 36731 14703 36737
rect 14921 36771 14979 36777
rect 14921 36737 14933 36771
rect 14967 36768 14979 36771
rect 15562 36768 15568 36780
rect 14967 36740 15568 36768
rect 14967 36737 14979 36740
rect 14921 36731 14979 36737
rect 15562 36728 15568 36740
rect 15620 36728 15626 36780
rect 16206 36728 16212 36780
rect 16264 36768 16270 36780
rect 18049 36771 18107 36777
rect 18049 36768 18061 36771
rect 16264 36740 18061 36768
rect 16264 36728 16270 36740
rect 18049 36737 18061 36740
rect 18095 36768 18107 36771
rect 18230 36768 18236 36780
rect 18095 36740 18236 36768
rect 18095 36737 18107 36740
rect 18049 36731 18107 36737
rect 18230 36728 18236 36740
rect 18288 36728 18294 36780
rect 18325 36771 18383 36777
rect 18325 36737 18337 36771
rect 18371 36768 18383 36771
rect 18414 36768 18420 36780
rect 18371 36740 18420 36768
rect 18371 36737 18383 36740
rect 18325 36731 18383 36737
rect 18414 36728 18420 36740
rect 18472 36728 18478 36780
rect 11885 36703 11943 36709
rect 11885 36669 11897 36703
rect 11931 36669 11943 36703
rect 11885 36663 11943 36669
rect 12437 36703 12495 36709
rect 12437 36669 12449 36703
rect 12483 36669 12495 36703
rect 12802 36700 12808 36712
rect 12763 36672 12808 36700
rect 12437 36663 12495 36669
rect 11900 36632 11928 36663
rect 12802 36660 12808 36672
rect 12860 36660 12866 36712
rect 13170 36700 13176 36712
rect 13131 36672 13176 36700
rect 13170 36660 13176 36672
rect 13228 36660 13234 36712
rect 15010 36660 15016 36712
rect 15068 36700 15074 36712
rect 16761 36703 16819 36709
rect 16761 36700 16773 36703
rect 15068 36672 16773 36700
rect 15068 36660 15074 36672
rect 16761 36669 16773 36672
rect 16807 36669 16819 36703
rect 16761 36663 16819 36669
rect 17497 36703 17555 36709
rect 17497 36669 17509 36703
rect 17543 36700 17555 36703
rect 19794 36700 19800 36712
rect 17543 36672 19800 36700
rect 17543 36669 17555 36672
rect 17497 36663 17555 36669
rect 12986 36632 12992 36644
rect 11900 36604 12992 36632
rect 12986 36592 12992 36604
rect 13044 36592 13050 36644
rect 16301 36635 16359 36641
rect 16301 36601 16313 36635
rect 16347 36632 16359 36635
rect 17512 36632 17540 36663
rect 19794 36660 19800 36672
rect 19852 36660 19858 36712
rect 20349 36703 20407 36709
rect 20349 36669 20361 36703
rect 20395 36700 20407 36703
rect 21174 36700 21180 36712
rect 20395 36672 21180 36700
rect 20395 36669 20407 36672
rect 20349 36663 20407 36669
rect 21174 36660 21180 36672
rect 21232 36660 21238 36712
rect 21729 36703 21787 36709
rect 21729 36669 21741 36703
rect 21775 36669 21787 36703
rect 21910 36700 21916 36712
rect 21871 36672 21916 36700
rect 21729 36663 21787 36669
rect 16347 36604 17540 36632
rect 16347 36601 16359 36604
rect 16301 36595 16359 36601
rect 12158 36564 12164 36576
rect 10060 36536 12164 36564
rect 12158 36524 12164 36536
rect 12216 36524 12222 36576
rect 12802 36524 12808 36576
rect 12860 36564 12866 36576
rect 14918 36564 14924 36576
rect 12860 36536 14924 36564
rect 12860 36524 12866 36536
rect 14918 36524 14924 36536
rect 14976 36524 14982 36576
rect 15010 36524 15016 36576
rect 15068 36564 15074 36576
rect 16316 36564 16344 36595
rect 20070 36592 20076 36644
rect 20128 36632 20134 36644
rect 21744 36632 21772 36663
rect 21910 36660 21916 36672
rect 21968 36660 21974 36712
rect 22296 36709 22324 36808
rect 23934 36728 23940 36780
rect 23992 36768 23998 36780
rect 25774 36768 25780 36780
rect 23992 36740 24440 36768
rect 25735 36740 25780 36768
rect 23992 36728 23998 36740
rect 22281 36703 22339 36709
rect 22281 36669 22293 36703
rect 22327 36669 22339 36703
rect 22281 36663 22339 36669
rect 22925 36703 22983 36709
rect 22925 36669 22937 36703
rect 22971 36700 22983 36703
rect 23474 36700 23480 36712
rect 22971 36672 23480 36700
rect 22971 36669 22983 36672
rect 22925 36663 22983 36669
rect 23474 36660 23480 36672
rect 23532 36700 23538 36712
rect 24118 36700 24124 36712
rect 23532 36672 24124 36700
rect 23532 36660 23538 36672
rect 24118 36660 24124 36672
rect 24176 36660 24182 36712
rect 24302 36700 24308 36712
rect 24263 36672 24308 36700
rect 24302 36660 24308 36672
rect 24360 36660 24366 36712
rect 24412 36709 24440 36740
rect 25774 36728 25780 36740
rect 25832 36728 25838 36780
rect 29270 36768 29276 36780
rect 29231 36740 29276 36768
rect 29270 36728 29276 36740
rect 29328 36728 29334 36780
rect 29549 36771 29607 36777
rect 29549 36737 29561 36771
rect 29595 36768 29607 36771
rect 30006 36768 30012 36780
rect 29595 36740 30012 36768
rect 29595 36737 29607 36740
rect 29549 36731 29607 36737
rect 30006 36728 30012 36740
rect 30064 36728 30070 36780
rect 24397 36703 24455 36709
rect 24397 36669 24409 36703
rect 24443 36669 24455 36703
rect 26050 36700 26056 36712
rect 26011 36672 26056 36700
rect 24397 36663 24455 36669
rect 26050 36660 26056 36672
rect 26108 36660 26114 36712
rect 28166 36700 28172 36712
rect 28127 36672 28172 36700
rect 28166 36660 28172 36672
rect 28224 36660 28230 36712
rect 28261 36703 28319 36709
rect 28261 36669 28273 36703
rect 28307 36700 28319 36703
rect 28994 36700 29000 36712
rect 28307 36672 29000 36700
rect 28307 36669 28319 36672
rect 28261 36663 28319 36669
rect 28994 36660 29000 36672
rect 29052 36660 29058 36712
rect 32490 36700 32496 36712
rect 29380 36672 32496 36700
rect 23566 36632 23572 36644
rect 20128 36604 21128 36632
rect 21744 36604 23572 36632
rect 20128 36592 20134 36604
rect 15068 36536 16344 36564
rect 15068 36524 15074 36536
rect 18138 36524 18144 36576
rect 18196 36564 18202 36576
rect 19429 36567 19487 36573
rect 19429 36564 19441 36567
rect 18196 36536 19441 36564
rect 18196 36524 18202 36536
rect 19429 36533 19441 36536
rect 19475 36564 19487 36567
rect 20254 36564 20260 36576
rect 19475 36536 20260 36564
rect 19475 36533 19487 36536
rect 19429 36527 19487 36533
rect 20254 36524 20260 36536
rect 20312 36524 20318 36576
rect 20438 36564 20444 36576
rect 20399 36536 20444 36564
rect 20438 36524 20444 36536
rect 20496 36524 20502 36576
rect 21100 36564 21128 36604
rect 23566 36592 23572 36604
rect 23624 36592 23630 36644
rect 27430 36592 27436 36644
rect 27488 36632 27494 36644
rect 29380 36632 29408 36672
rect 32490 36660 32496 36672
rect 32548 36660 32554 36712
rect 32585 36703 32643 36709
rect 32585 36669 32597 36703
rect 32631 36700 32643 36703
rect 37550 36700 37556 36712
rect 32631 36672 37556 36700
rect 32631 36669 32643 36672
rect 32585 36663 32643 36669
rect 37550 36660 37556 36672
rect 37608 36660 37614 36712
rect 27488 36604 29408 36632
rect 27488 36592 27494 36604
rect 25130 36564 25136 36576
rect 21100 36536 25136 36564
rect 25130 36524 25136 36536
rect 25188 36524 25194 36576
rect 26418 36524 26424 36576
rect 26476 36564 26482 36576
rect 27157 36567 27215 36573
rect 27157 36564 27169 36567
rect 26476 36536 27169 36564
rect 26476 36524 26482 36536
rect 27157 36533 27169 36536
rect 27203 36533 27215 36567
rect 30650 36564 30656 36576
rect 30611 36536 30656 36564
rect 27157 36527 27215 36533
rect 30650 36524 30656 36536
rect 30708 36524 30714 36576
rect 1104 36474 39836 36496
rect 1104 36422 19606 36474
rect 19658 36422 19670 36474
rect 19722 36422 19734 36474
rect 19786 36422 19798 36474
rect 19850 36422 39836 36474
rect 1104 36400 39836 36422
rect 7190 36320 7196 36372
rect 7248 36320 7254 36372
rect 8570 36360 8576 36372
rect 8531 36332 8576 36360
rect 8570 36320 8576 36332
rect 8628 36320 8634 36372
rect 11054 36360 11060 36372
rect 11015 36332 11060 36360
rect 11054 36320 11060 36332
rect 11112 36320 11118 36372
rect 11146 36320 11152 36372
rect 11204 36360 11210 36372
rect 11204 36332 30420 36360
rect 11204 36320 11210 36332
rect 5350 36252 5356 36304
rect 5408 36292 5414 36304
rect 7208 36292 7236 36320
rect 5408 36264 7236 36292
rect 5408 36252 5414 36264
rect 4249 36227 4307 36233
rect 4249 36193 4261 36227
rect 4295 36193 4307 36227
rect 4798 36224 4804 36236
rect 4759 36196 4804 36224
rect 4249 36187 4307 36193
rect 4264 36156 4292 36187
rect 4798 36184 4804 36196
rect 4856 36184 4862 36236
rect 6196 36233 6224 36264
rect 7650 36252 7656 36304
rect 7708 36292 7714 36304
rect 9674 36292 9680 36304
rect 7708 36264 9680 36292
rect 7708 36252 7714 36264
rect 9674 36252 9680 36264
rect 9732 36252 9738 36304
rect 13725 36295 13783 36301
rect 13725 36261 13737 36295
rect 13771 36292 13783 36295
rect 14734 36292 14740 36304
rect 13771 36264 14740 36292
rect 13771 36261 13783 36264
rect 13725 36255 13783 36261
rect 14734 36252 14740 36264
rect 14792 36252 14798 36304
rect 14918 36252 14924 36304
rect 14976 36292 14982 36304
rect 17034 36292 17040 36304
rect 14976 36264 17040 36292
rect 14976 36252 14982 36264
rect 17034 36252 17040 36264
rect 17092 36252 17098 36304
rect 18233 36295 18291 36301
rect 18233 36261 18245 36295
rect 18279 36292 18291 36295
rect 18506 36292 18512 36304
rect 18279 36264 18512 36292
rect 18279 36261 18291 36264
rect 18233 36255 18291 36261
rect 18506 36252 18512 36264
rect 18564 36252 18570 36304
rect 19426 36292 19432 36304
rect 19076 36264 19432 36292
rect 6181 36227 6239 36233
rect 6181 36193 6193 36227
rect 6227 36193 6239 36227
rect 6181 36187 6239 36193
rect 6365 36227 6423 36233
rect 6365 36193 6377 36227
rect 6411 36193 6423 36227
rect 6638 36224 6644 36236
rect 6599 36196 6644 36224
rect 6365 36187 6423 36193
rect 4706 36156 4712 36168
rect 4264 36128 4712 36156
rect 4706 36116 4712 36128
rect 4764 36116 4770 36168
rect 5074 36156 5080 36168
rect 5035 36128 5080 36156
rect 5074 36116 5080 36128
rect 5132 36116 5138 36168
rect 4341 36091 4399 36097
rect 4341 36057 4353 36091
rect 4387 36088 4399 36091
rect 4614 36088 4620 36100
rect 4387 36060 4620 36088
rect 4387 36057 4399 36060
rect 4341 36051 4399 36057
rect 4614 36048 4620 36060
rect 4672 36048 4678 36100
rect 5994 36088 6000 36100
rect 5955 36060 6000 36088
rect 5994 36048 6000 36060
rect 6052 36048 6058 36100
rect 14 35980 20 36032
rect 72 36020 78 36032
rect 750 36020 756 36032
rect 72 35992 756 36020
rect 72 35980 78 35992
rect 750 35980 756 35992
rect 808 35980 814 36032
rect 6380 36020 6408 36187
rect 6638 36184 6644 36196
rect 6696 36184 6702 36236
rect 7374 36224 7380 36236
rect 7335 36196 7380 36224
rect 7374 36184 7380 36196
rect 7432 36184 7438 36236
rect 7837 36227 7895 36233
rect 7837 36193 7849 36227
rect 7883 36193 7895 36227
rect 7837 36187 7895 36193
rect 8481 36227 8539 36233
rect 8481 36193 8493 36227
rect 8527 36193 8539 36227
rect 9950 36224 9956 36236
rect 9911 36196 9956 36224
rect 8481 36187 8539 36193
rect 6454 36116 6460 36168
rect 6512 36156 6518 36168
rect 7852 36156 7880 36187
rect 6512 36128 7880 36156
rect 6512 36116 6518 36128
rect 6730 36048 6736 36100
rect 6788 36088 6794 36100
rect 8496 36088 8524 36187
rect 9950 36184 9956 36196
rect 10008 36184 10014 36236
rect 11422 36184 11428 36236
rect 11480 36224 11486 36236
rect 12802 36224 12808 36236
rect 11480 36196 12808 36224
rect 11480 36184 11486 36196
rect 12802 36184 12808 36196
rect 12860 36184 12866 36236
rect 12986 36224 12992 36236
rect 12947 36196 12992 36224
rect 12986 36184 12992 36196
rect 13044 36184 13050 36236
rect 14553 36227 14611 36233
rect 14553 36224 14565 36227
rect 13096 36196 14565 36224
rect 13096 36168 13124 36196
rect 14553 36193 14565 36196
rect 14599 36193 14611 36227
rect 15102 36224 15108 36236
rect 14553 36187 14611 36193
rect 14660 36196 15108 36224
rect 9306 36116 9312 36168
rect 9364 36156 9370 36168
rect 9677 36159 9735 36165
rect 9677 36156 9689 36159
rect 9364 36128 9689 36156
rect 9364 36116 9370 36128
rect 9677 36125 9689 36128
rect 9723 36125 9735 36159
rect 13078 36156 13084 36168
rect 13039 36128 13084 36156
rect 9677 36119 9735 36125
rect 13078 36116 13084 36128
rect 13136 36116 13142 36168
rect 14277 36159 14335 36165
rect 14277 36125 14289 36159
rect 14323 36156 14335 36159
rect 14660 36156 14688 36196
rect 15102 36184 15108 36196
rect 15160 36184 15166 36236
rect 15289 36227 15347 36233
rect 15289 36193 15301 36227
rect 15335 36224 15347 36227
rect 16298 36224 16304 36236
rect 15335 36196 16304 36224
rect 15335 36193 15347 36196
rect 15289 36187 15347 36193
rect 16298 36184 16304 36196
rect 16356 36184 16362 36236
rect 16393 36227 16451 36233
rect 16393 36193 16405 36227
rect 16439 36193 16451 36227
rect 16574 36224 16580 36236
rect 16535 36196 16580 36224
rect 16393 36187 16451 36193
rect 14323 36128 14688 36156
rect 14737 36159 14795 36165
rect 14323 36125 14335 36128
rect 14277 36119 14335 36125
rect 14737 36125 14749 36159
rect 14783 36156 14795 36159
rect 15010 36156 15016 36168
rect 14783 36128 15016 36156
rect 14783 36125 14795 36128
rect 14737 36119 14795 36125
rect 15010 36116 15016 36128
rect 15068 36116 15074 36168
rect 16316 36088 16344 36184
rect 16408 36156 16436 36187
rect 16574 36184 16580 36196
rect 16632 36184 16638 36236
rect 16850 36224 16856 36236
rect 16811 36196 16856 36224
rect 16850 36184 16856 36196
rect 16908 36184 16914 36236
rect 18138 36224 18144 36236
rect 18099 36196 18144 36224
rect 18138 36184 18144 36196
rect 18196 36184 18202 36236
rect 19076 36233 19104 36264
rect 19426 36252 19432 36264
rect 19484 36292 19490 36304
rect 20438 36292 20444 36304
rect 19484 36264 20444 36292
rect 19484 36252 19490 36264
rect 20438 36252 20444 36264
rect 20496 36292 20502 36304
rect 20496 36264 21772 36292
rect 20496 36252 20502 36264
rect 19061 36227 19119 36233
rect 19061 36193 19073 36227
rect 19107 36193 19119 36227
rect 19061 36187 19119 36193
rect 19150 36184 19156 36236
rect 19208 36224 19214 36236
rect 19245 36227 19303 36233
rect 19245 36224 19257 36227
rect 19208 36196 19257 36224
rect 19208 36184 19214 36196
rect 19245 36193 19257 36196
rect 19291 36193 19303 36227
rect 19245 36187 19303 36193
rect 19334 36184 19340 36236
rect 19392 36224 19398 36236
rect 19613 36227 19671 36233
rect 19613 36224 19625 36227
rect 19392 36196 19625 36224
rect 19392 36184 19398 36196
rect 19613 36193 19625 36196
rect 19659 36193 19671 36227
rect 19613 36187 19671 36193
rect 19981 36227 20039 36233
rect 19981 36193 19993 36227
rect 20027 36193 20039 36227
rect 19981 36187 20039 36193
rect 20257 36227 20315 36233
rect 20257 36193 20269 36227
rect 20303 36224 20315 36227
rect 20530 36224 20536 36236
rect 20303 36196 20536 36224
rect 20303 36193 20315 36196
rect 20257 36187 20315 36193
rect 16666 36156 16672 36168
rect 16408 36128 16672 36156
rect 16666 36116 16672 36128
rect 16724 36116 16730 36168
rect 17310 36156 17316 36168
rect 17271 36128 17316 36156
rect 17310 36116 17316 36128
rect 17368 36116 17374 36168
rect 18690 36116 18696 36168
rect 18748 36156 18754 36168
rect 19996 36156 20024 36187
rect 20530 36184 20536 36196
rect 20588 36224 20594 36236
rect 20898 36224 20904 36236
rect 20588 36196 20904 36224
rect 20588 36184 20594 36196
rect 20898 36184 20904 36196
rect 20956 36184 20962 36236
rect 21266 36224 21272 36236
rect 21227 36196 21272 36224
rect 21266 36184 21272 36196
rect 21324 36184 21330 36236
rect 21744 36233 21772 36264
rect 26050 36252 26056 36304
rect 26108 36292 26114 36304
rect 27065 36295 27123 36301
rect 27065 36292 27077 36295
rect 26108 36264 27077 36292
rect 26108 36252 26114 36264
rect 27065 36261 27077 36264
rect 27111 36261 27123 36295
rect 27065 36255 27123 36261
rect 21729 36227 21787 36233
rect 21729 36193 21741 36227
rect 21775 36193 21787 36227
rect 21729 36187 21787 36193
rect 22741 36227 22799 36233
rect 22741 36193 22753 36227
rect 22787 36193 22799 36227
rect 22741 36187 22799 36193
rect 18748 36128 20024 36156
rect 18748 36116 18754 36128
rect 20622 36116 20628 36168
rect 20680 36156 20686 36168
rect 20993 36159 21051 36165
rect 20993 36156 21005 36159
rect 20680 36128 21005 36156
rect 20680 36116 20686 36128
rect 20993 36125 21005 36128
rect 21039 36125 21051 36159
rect 22756 36156 22784 36187
rect 22830 36184 22836 36236
rect 22888 36224 22894 36236
rect 23293 36227 23351 36233
rect 22888 36196 22933 36224
rect 22888 36184 22894 36196
rect 23293 36193 23305 36227
rect 23339 36224 23351 36227
rect 24029 36227 24087 36233
rect 24029 36224 24041 36227
rect 23339 36196 24041 36224
rect 23339 36193 23351 36196
rect 23293 36187 23351 36193
rect 24029 36193 24041 36196
rect 24075 36193 24087 36227
rect 26602 36224 26608 36236
rect 26563 36196 26608 36224
rect 24029 36187 24087 36193
rect 26602 36184 26608 36196
rect 26660 36184 26666 36236
rect 27798 36224 27804 36236
rect 27448 36196 27660 36224
rect 27759 36196 27804 36224
rect 23750 36156 23756 36168
rect 20993 36119 21051 36125
rect 21836 36128 22784 36156
rect 23711 36128 23756 36156
rect 19150 36088 19156 36100
rect 6788 36060 8524 36088
rect 12452 36060 15608 36088
rect 16316 36060 19156 36088
rect 6788 36048 6794 36060
rect 6914 36020 6920 36032
rect 6380 35992 6920 36020
rect 6914 35980 6920 35992
rect 6972 36020 6978 36032
rect 7190 36020 7196 36032
rect 6972 35992 7196 36020
rect 6972 35980 6978 35992
rect 7190 35980 7196 35992
rect 7248 35980 7254 36032
rect 7926 36020 7932 36032
rect 7887 35992 7932 36020
rect 7926 35980 7932 35992
rect 7984 35980 7990 36032
rect 9674 35980 9680 36032
rect 9732 36020 9738 36032
rect 12452 36020 12480 36060
rect 9732 35992 12480 36020
rect 9732 35980 9738 35992
rect 14918 35980 14924 36032
rect 14976 36020 14982 36032
rect 15381 36023 15439 36029
rect 15381 36020 15393 36023
rect 14976 35992 15393 36020
rect 14976 35980 14982 35992
rect 15381 35989 15393 35992
rect 15427 35989 15439 36023
rect 15580 36020 15608 36060
rect 19150 36048 19156 36060
rect 19208 36048 19214 36100
rect 20714 36048 20720 36100
rect 20772 36088 20778 36100
rect 21729 36091 21787 36097
rect 21729 36088 21741 36091
rect 20772 36060 21741 36088
rect 20772 36048 20778 36060
rect 21729 36057 21741 36060
rect 21775 36057 21787 36091
rect 21729 36051 21787 36057
rect 21836 36020 21864 36128
rect 23750 36116 23756 36128
rect 23808 36116 23814 36168
rect 25406 36116 25412 36168
rect 25464 36156 25470 36168
rect 26513 36159 26571 36165
rect 26513 36156 26525 36159
rect 25464 36128 26525 36156
rect 25464 36116 25470 36128
rect 26513 36125 26525 36128
rect 26559 36156 26571 36159
rect 27448 36156 27476 36196
rect 26559 36128 27476 36156
rect 27525 36159 27583 36165
rect 26559 36125 26571 36128
rect 26513 36119 26571 36125
rect 27525 36125 27537 36159
rect 27571 36125 27583 36159
rect 27632 36156 27660 36196
rect 27798 36184 27804 36196
rect 27856 36184 27862 36236
rect 30392 36233 30420 36332
rect 31202 36320 31208 36372
rect 31260 36360 31266 36372
rect 31260 36332 35020 36360
rect 31260 36320 31266 36332
rect 33413 36295 33471 36301
rect 33413 36261 33425 36295
rect 33459 36292 33471 36295
rect 34514 36292 34520 36304
rect 33459 36264 34520 36292
rect 33459 36261 33471 36264
rect 33413 36255 33471 36261
rect 34514 36252 34520 36264
rect 34572 36252 34578 36304
rect 30377 36227 30435 36233
rect 30377 36193 30389 36227
rect 30423 36193 30435 36227
rect 30377 36187 30435 36193
rect 32490 36184 32496 36236
rect 32548 36224 32554 36236
rect 32861 36227 32919 36233
rect 32861 36224 32873 36227
rect 32548 36196 32873 36224
rect 32548 36184 32554 36196
rect 32861 36193 32873 36196
rect 32907 36193 32919 36227
rect 32861 36187 32919 36193
rect 32953 36227 33011 36233
rect 32953 36193 32965 36227
rect 32999 36224 33011 36227
rect 33134 36224 33140 36236
rect 32999 36196 33140 36224
rect 32999 36193 33011 36196
rect 32953 36187 33011 36193
rect 28166 36156 28172 36168
rect 27632 36128 28172 36156
rect 27525 36119 27583 36125
rect 27246 36048 27252 36100
rect 27304 36088 27310 36100
rect 27540 36088 27568 36119
rect 28166 36116 28172 36128
rect 28224 36116 28230 36168
rect 30285 36159 30343 36165
rect 30285 36125 30297 36159
rect 30331 36125 30343 36159
rect 30285 36119 30343 36125
rect 30837 36159 30895 36165
rect 30837 36125 30849 36159
rect 30883 36156 30895 36159
rect 32306 36156 32312 36168
rect 30883 36128 32312 36156
rect 30883 36125 30895 36128
rect 30837 36119 30895 36125
rect 27304 36060 27568 36088
rect 30300 36088 30328 36119
rect 32306 36116 32312 36128
rect 32364 36116 32370 36168
rect 32876 36156 32904 36187
rect 33134 36184 33140 36196
rect 33192 36184 33198 36236
rect 33962 36224 33968 36236
rect 33923 36196 33968 36224
rect 33962 36184 33968 36196
rect 34020 36184 34026 36236
rect 34992 36233 35020 36332
rect 34977 36227 35035 36233
rect 34977 36193 34989 36227
rect 35023 36193 35035 36227
rect 34977 36187 35035 36193
rect 35069 36227 35127 36233
rect 35069 36193 35081 36227
rect 35115 36224 35127 36227
rect 35894 36224 35900 36236
rect 35115 36196 35900 36224
rect 35115 36193 35127 36196
rect 35069 36187 35127 36193
rect 35894 36184 35900 36196
rect 35952 36184 35958 36236
rect 33873 36159 33931 36165
rect 33873 36156 33885 36159
rect 32876 36128 33885 36156
rect 33873 36125 33885 36128
rect 33919 36125 33931 36159
rect 33873 36119 33931 36125
rect 31202 36088 31208 36100
rect 30300 36060 31208 36088
rect 27304 36048 27310 36060
rect 31202 36048 31208 36060
rect 31260 36048 31266 36100
rect 22554 36020 22560 36032
rect 15580 35992 21864 36020
rect 22515 35992 22560 36020
rect 15381 35983 15439 35989
rect 22554 35980 22560 35992
rect 22612 35980 22618 36032
rect 25317 36023 25375 36029
rect 25317 35989 25329 36023
rect 25363 36020 25375 36023
rect 25866 36020 25872 36032
rect 25363 35992 25872 36020
rect 25363 35989 25375 35992
rect 25317 35983 25375 35989
rect 25866 35980 25872 35992
rect 25924 35980 25930 36032
rect 27798 35980 27804 36032
rect 27856 36020 27862 36032
rect 28905 36023 28963 36029
rect 28905 36020 28917 36023
rect 27856 35992 28917 36020
rect 27856 35980 27862 35992
rect 28905 35989 28917 35992
rect 28951 35989 28963 36023
rect 34146 36020 34152 36032
rect 34107 35992 34152 36020
rect 28905 35983 28963 35989
rect 34146 35980 34152 35992
rect 34204 35980 34210 36032
rect 35250 36020 35256 36032
rect 35211 35992 35256 36020
rect 35250 35980 35256 35992
rect 35308 35980 35314 36032
rect 1104 35930 39836 35952
rect 1104 35878 4246 35930
rect 4298 35878 4310 35930
rect 4362 35878 4374 35930
rect 4426 35878 4438 35930
rect 4490 35878 34966 35930
rect 35018 35878 35030 35930
rect 35082 35878 35094 35930
rect 35146 35878 35158 35930
rect 35210 35878 39836 35930
rect 1104 35856 39836 35878
rect 7374 35776 7380 35828
rect 7432 35816 7438 35828
rect 8018 35816 8024 35828
rect 7432 35788 8024 35816
rect 7432 35776 7438 35788
rect 8018 35776 8024 35788
rect 8076 35816 8082 35828
rect 9217 35819 9275 35825
rect 9217 35816 9229 35819
rect 8076 35788 9229 35816
rect 8076 35776 8082 35788
rect 9217 35785 9229 35788
rect 9263 35785 9275 35819
rect 16666 35816 16672 35828
rect 16627 35788 16672 35816
rect 9217 35779 9275 35785
rect 16666 35776 16672 35788
rect 16724 35776 16730 35828
rect 23382 35776 23388 35828
rect 23440 35816 23446 35828
rect 23845 35819 23903 35825
rect 23845 35816 23857 35819
rect 23440 35788 23857 35816
rect 23440 35776 23446 35788
rect 23845 35785 23857 35788
rect 23891 35785 23903 35819
rect 23845 35779 23903 35785
rect 25774 35776 25780 35828
rect 25832 35816 25838 35828
rect 26326 35816 26332 35828
rect 25832 35788 26332 35816
rect 25832 35776 25838 35788
rect 26326 35776 26332 35788
rect 26384 35816 26390 35828
rect 27246 35816 27252 35828
rect 26384 35788 27252 35816
rect 26384 35776 26390 35788
rect 27246 35776 27252 35788
rect 27304 35776 27310 35828
rect 33597 35819 33655 35825
rect 33597 35785 33609 35819
rect 33643 35816 33655 35819
rect 33962 35816 33968 35828
rect 33643 35788 33968 35816
rect 33643 35785 33655 35788
rect 33597 35779 33655 35785
rect 33962 35776 33968 35788
rect 34020 35776 34026 35828
rect 36265 35819 36323 35825
rect 36265 35816 36277 35819
rect 34072 35788 36277 35816
rect 4706 35748 4712 35760
rect 4667 35720 4712 35748
rect 4706 35708 4712 35720
rect 4764 35708 4770 35760
rect 11241 35751 11299 35757
rect 11241 35717 11253 35751
rect 11287 35717 11299 35751
rect 11241 35711 11299 35717
rect 4065 35683 4123 35689
rect 4065 35649 4077 35683
rect 4111 35680 4123 35683
rect 4798 35680 4804 35692
rect 4111 35652 4804 35680
rect 4111 35649 4123 35652
rect 4065 35643 4123 35649
rect 4798 35640 4804 35652
rect 4856 35640 4862 35692
rect 6273 35683 6331 35689
rect 6273 35649 6285 35683
rect 6319 35680 6331 35683
rect 6638 35680 6644 35692
rect 6319 35652 6644 35680
rect 6319 35649 6331 35652
rect 6273 35643 6331 35649
rect 6638 35640 6644 35652
rect 6696 35640 6702 35692
rect 7837 35683 7895 35689
rect 7837 35649 7849 35683
rect 7883 35680 7895 35683
rect 9306 35680 9312 35692
rect 7883 35652 9312 35680
rect 7883 35649 7895 35652
rect 7837 35643 7895 35649
rect 9306 35640 9312 35652
rect 9364 35640 9370 35692
rect 11256 35680 11284 35711
rect 12158 35708 12164 35760
rect 12216 35748 12222 35760
rect 12216 35720 18276 35748
rect 12216 35708 12222 35720
rect 10520 35652 11284 35680
rect 12989 35683 13047 35689
rect 4433 35615 4491 35621
rect 4433 35581 4445 35615
rect 4479 35581 4491 35615
rect 4433 35575 4491 35581
rect 4709 35615 4767 35621
rect 4709 35581 4721 35615
rect 4755 35612 4767 35615
rect 5813 35615 5871 35621
rect 4755 35584 5764 35612
rect 4755 35581 4767 35584
rect 4709 35575 4767 35581
rect 4448 35544 4476 35575
rect 5074 35544 5080 35556
rect 4448 35516 5080 35544
rect 5074 35504 5080 35516
rect 5132 35504 5138 35556
rect 5736 35476 5764 35584
rect 5813 35581 5825 35615
rect 5859 35581 5871 35615
rect 6086 35612 6092 35624
rect 6047 35584 6092 35612
rect 5813 35575 5871 35581
rect 5828 35544 5856 35575
rect 6086 35572 6092 35584
rect 6144 35612 6150 35624
rect 6730 35612 6736 35624
rect 6144 35584 6736 35612
rect 6144 35572 6150 35584
rect 6730 35572 6736 35584
rect 6788 35612 6794 35624
rect 6825 35615 6883 35621
rect 6825 35612 6837 35615
rect 6788 35584 6837 35612
rect 6788 35572 6794 35584
rect 6825 35581 6837 35584
rect 6871 35581 6883 35615
rect 6825 35575 6883 35581
rect 8113 35615 8171 35621
rect 8113 35581 8125 35615
rect 8159 35612 8171 35615
rect 10410 35612 10416 35624
rect 8159 35584 10416 35612
rect 8159 35581 8171 35584
rect 8113 35575 8171 35581
rect 10410 35572 10416 35584
rect 10468 35572 10474 35624
rect 10520 35621 10548 35652
rect 12989 35649 13001 35683
rect 13035 35680 13047 35683
rect 15102 35680 15108 35692
rect 13035 35652 15108 35680
rect 13035 35649 13047 35652
rect 12989 35643 13047 35649
rect 15102 35640 15108 35652
rect 15160 35640 15166 35692
rect 16117 35683 16175 35689
rect 16117 35649 16129 35683
rect 16163 35680 16175 35683
rect 16850 35680 16856 35692
rect 16163 35652 16856 35680
rect 16163 35649 16175 35652
rect 16117 35643 16175 35649
rect 16850 35640 16856 35652
rect 16908 35640 16914 35692
rect 17144 35652 18184 35680
rect 10505 35615 10563 35621
rect 10505 35581 10517 35615
rect 10551 35581 10563 35615
rect 11146 35612 11152 35624
rect 11107 35584 11152 35612
rect 10505 35575 10563 35581
rect 11146 35572 11152 35584
rect 11204 35572 11210 35624
rect 11885 35615 11943 35621
rect 11885 35581 11897 35615
rect 11931 35612 11943 35615
rect 12437 35615 12495 35621
rect 12437 35612 12449 35615
rect 11931 35584 12449 35612
rect 11931 35581 11943 35584
rect 11885 35575 11943 35581
rect 12437 35581 12449 35584
rect 12483 35581 12495 35615
rect 13262 35612 13268 35624
rect 13223 35584 13268 35612
rect 12437 35575 12495 35581
rect 13262 35572 13268 35584
rect 13320 35572 13326 35624
rect 13449 35615 13507 35621
rect 13449 35581 13461 35615
rect 13495 35612 13507 35615
rect 13630 35612 13636 35624
rect 13495 35584 13636 35612
rect 13495 35581 13507 35584
rect 13449 35575 13507 35581
rect 13630 35572 13636 35584
rect 13688 35572 13694 35624
rect 14918 35612 14924 35624
rect 14879 35584 14924 35612
rect 14918 35572 14924 35584
rect 14976 35572 14982 35624
rect 15562 35612 15568 35624
rect 15523 35584 15568 35612
rect 15562 35572 15568 35584
rect 15620 35572 15626 35624
rect 15838 35612 15844 35624
rect 15799 35584 15844 35612
rect 15838 35572 15844 35584
rect 15896 35572 15902 35624
rect 16758 35612 16764 35624
rect 16719 35584 16764 35612
rect 16758 35572 16764 35584
rect 16816 35572 16822 35624
rect 16942 35572 16948 35624
rect 17000 35612 17006 35624
rect 17144 35621 17172 35652
rect 17129 35615 17187 35621
rect 17129 35612 17141 35615
rect 17000 35584 17141 35612
rect 17000 35572 17006 35584
rect 17129 35581 17141 35584
rect 17175 35581 17187 35615
rect 17129 35575 17187 35581
rect 6178 35544 6184 35556
rect 5828 35516 6184 35544
rect 6178 35504 6184 35516
rect 6236 35544 6242 35556
rect 7926 35544 7932 35556
rect 6236 35516 7932 35544
rect 6236 35504 6242 35516
rect 7926 35504 7932 35516
rect 7984 35504 7990 35556
rect 18156 35544 18184 35652
rect 18248 35621 18276 35720
rect 20254 35708 20260 35760
rect 20312 35748 20318 35760
rect 21358 35748 21364 35760
rect 20312 35720 21364 35748
rect 20312 35708 20318 35720
rect 21358 35708 21364 35720
rect 21416 35748 21422 35760
rect 21818 35748 21824 35760
rect 21416 35720 21824 35748
rect 21416 35708 21422 35720
rect 21818 35708 21824 35720
rect 21876 35748 21882 35760
rect 21876 35720 23704 35748
rect 21876 35708 21882 35720
rect 18782 35680 18788 35692
rect 18743 35652 18788 35680
rect 18782 35640 18788 35652
rect 18840 35640 18846 35692
rect 20622 35680 20628 35692
rect 19628 35652 20628 35680
rect 18233 35615 18291 35621
rect 18233 35581 18245 35615
rect 18279 35612 18291 35615
rect 18322 35612 18328 35624
rect 18279 35584 18328 35612
rect 18279 35581 18291 35584
rect 18233 35575 18291 35581
rect 18322 35572 18328 35584
rect 18380 35572 18386 35624
rect 18874 35612 18880 35624
rect 18835 35584 18880 35612
rect 18874 35572 18880 35584
rect 18932 35572 18938 35624
rect 19334 35572 19340 35624
rect 19392 35612 19398 35624
rect 19628 35621 19656 35652
rect 20622 35640 20628 35652
rect 20680 35640 20686 35692
rect 21910 35680 21916 35692
rect 21560 35652 21916 35680
rect 21560 35621 21588 35652
rect 21910 35640 21916 35652
rect 21968 35640 21974 35692
rect 19613 35615 19671 35621
rect 19613 35612 19625 35615
rect 19392 35584 19625 35612
rect 19392 35572 19398 35584
rect 19613 35581 19625 35584
rect 19659 35581 19671 35615
rect 19613 35575 19671 35581
rect 20073 35615 20131 35621
rect 20073 35581 20085 35615
rect 20119 35581 20131 35615
rect 20073 35575 20131 35581
rect 21545 35615 21603 35621
rect 21545 35581 21557 35615
rect 21591 35581 21603 35615
rect 21545 35575 21603 35581
rect 19886 35544 19892 35556
rect 18156 35516 19892 35544
rect 19886 35504 19892 35516
rect 19944 35544 19950 35556
rect 20088 35544 20116 35575
rect 21634 35572 21640 35624
rect 21692 35612 21698 35624
rect 21818 35612 21824 35624
rect 21692 35584 21737 35612
rect 21779 35584 21824 35612
rect 21692 35572 21698 35584
rect 21818 35572 21824 35584
rect 21876 35572 21882 35624
rect 22002 35612 22008 35624
rect 21963 35584 22008 35612
rect 22002 35572 22008 35584
rect 22060 35572 22066 35624
rect 22373 35615 22431 35621
rect 22373 35581 22385 35615
rect 22419 35612 22431 35615
rect 22646 35612 22652 35624
rect 22419 35584 22652 35612
rect 22419 35581 22431 35584
rect 22373 35575 22431 35581
rect 22646 35572 22652 35584
rect 22704 35572 22710 35624
rect 23676 35621 23704 35720
rect 26234 35708 26240 35760
rect 26292 35748 26298 35760
rect 28445 35751 28503 35757
rect 28445 35748 28457 35751
rect 26292 35720 28457 35748
rect 26292 35708 26298 35720
rect 28445 35717 28457 35720
rect 28491 35717 28503 35751
rect 28445 35711 28503 35717
rect 33134 35708 33140 35760
rect 33192 35748 33198 35760
rect 34072 35748 34100 35788
rect 36265 35785 36277 35788
rect 36311 35785 36323 35819
rect 36265 35779 36323 35785
rect 33192 35720 34100 35748
rect 33192 35708 33198 35720
rect 29362 35640 29368 35692
rect 29420 35680 29426 35692
rect 29917 35683 29975 35689
rect 29917 35680 29929 35683
rect 29420 35652 29929 35680
rect 29420 35640 29426 35652
rect 29917 35649 29929 35652
rect 29963 35649 29975 35683
rect 32030 35680 32036 35692
rect 31943 35652 32036 35680
rect 29917 35643 29975 35649
rect 32030 35640 32036 35652
rect 32088 35680 32094 35692
rect 32306 35680 32312 35692
rect 32088 35652 32168 35680
rect 32267 35652 32312 35680
rect 32088 35640 32094 35652
rect 23661 35615 23719 35621
rect 23661 35581 23673 35615
rect 23707 35581 23719 35615
rect 23661 35575 23719 35581
rect 24765 35615 24823 35621
rect 24765 35581 24777 35615
rect 24811 35612 24823 35615
rect 24854 35612 24860 35624
rect 24811 35584 24860 35612
rect 24811 35581 24823 35584
rect 24765 35575 24823 35581
rect 24854 35572 24860 35584
rect 24912 35572 24918 35624
rect 25038 35612 25044 35624
rect 24999 35584 25044 35612
rect 25038 35572 25044 35584
rect 25096 35572 25102 35624
rect 27433 35615 27491 35621
rect 27433 35581 27445 35615
rect 27479 35581 27491 35615
rect 27433 35575 27491 35581
rect 27525 35615 27583 35621
rect 27525 35581 27537 35615
rect 27571 35612 27583 35615
rect 27614 35612 27620 35624
rect 27571 35584 27620 35612
rect 27571 35581 27583 35584
rect 27525 35575 27583 35581
rect 19944 35516 20116 35544
rect 20349 35547 20407 35553
rect 19944 35504 19950 35516
rect 20349 35513 20361 35547
rect 20395 35544 20407 35547
rect 20898 35544 20904 35556
rect 20395 35516 20904 35544
rect 20395 35513 20407 35516
rect 20349 35507 20407 35513
rect 20898 35504 20904 35516
rect 20956 35504 20962 35556
rect 20993 35547 21051 35553
rect 20993 35513 21005 35547
rect 21039 35544 21051 35547
rect 22554 35544 22560 35556
rect 21039 35516 22560 35544
rect 21039 35513 21051 35516
rect 20993 35507 21051 35513
rect 22554 35504 22560 35516
rect 22612 35504 22618 35556
rect 27448 35544 27476 35575
rect 27614 35572 27620 35584
rect 27672 35612 27678 35624
rect 28261 35615 28319 35621
rect 28261 35612 28273 35615
rect 27672 35584 28273 35612
rect 27672 35572 27678 35584
rect 28261 35581 28273 35584
rect 28307 35612 28319 35615
rect 28442 35612 28448 35624
rect 28307 35584 28448 35612
rect 28307 35581 28319 35584
rect 28261 35575 28319 35581
rect 28442 35572 28448 35584
rect 28500 35572 28506 35624
rect 29825 35615 29883 35621
rect 29825 35581 29837 35615
rect 29871 35581 29883 35615
rect 30190 35612 30196 35624
rect 30151 35584 30196 35612
rect 29825 35575 29883 35581
rect 27448 35516 29684 35544
rect 6638 35476 6644 35488
rect 5736 35448 6644 35476
rect 6638 35436 6644 35448
rect 6696 35436 6702 35488
rect 7009 35479 7067 35485
rect 7009 35445 7021 35479
rect 7055 35476 7067 35479
rect 7742 35476 7748 35488
rect 7055 35448 7748 35476
rect 7055 35445 7067 35448
rect 7009 35439 7067 35445
rect 7742 35436 7748 35448
rect 7800 35436 7806 35488
rect 10597 35479 10655 35485
rect 10597 35445 10609 35479
rect 10643 35476 10655 35479
rect 11238 35476 11244 35488
rect 10643 35448 11244 35476
rect 10643 35445 10655 35448
rect 10597 35439 10655 35445
rect 11238 35436 11244 35448
rect 11296 35436 11302 35488
rect 18325 35479 18383 35485
rect 18325 35445 18337 35479
rect 18371 35476 18383 35479
rect 18414 35476 18420 35488
rect 18371 35448 18420 35476
rect 18371 35445 18383 35448
rect 18325 35439 18383 35445
rect 18414 35436 18420 35448
rect 18472 35436 18478 35488
rect 25498 35436 25504 35488
rect 25556 35476 25562 35488
rect 26145 35479 26203 35485
rect 26145 35476 26157 35479
rect 25556 35448 26157 35476
rect 25556 35436 25562 35448
rect 26145 35445 26157 35448
rect 26191 35445 26203 35479
rect 26145 35439 26203 35445
rect 27709 35479 27767 35485
rect 27709 35445 27721 35479
rect 27755 35476 27767 35479
rect 28166 35476 28172 35488
rect 27755 35448 28172 35476
rect 27755 35445 27767 35448
rect 27709 35439 27767 35445
rect 28166 35436 28172 35448
rect 28224 35436 28230 35488
rect 29656 35485 29684 35516
rect 29641 35479 29699 35485
rect 29641 35445 29653 35479
rect 29687 35476 29699 35479
rect 29730 35476 29736 35488
rect 29687 35448 29736 35476
rect 29687 35445 29699 35448
rect 29641 35439 29699 35445
rect 29730 35436 29736 35448
rect 29788 35436 29794 35488
rect 29840 35476 29868 35575
rect 30190 35572 30196 35584
rect 30248 35572 30254 35624
rect 32140 35544 32168 35652
rect 32306 35640 32312 35652
rect 32364 35640 32370 35692
rect 35161 35683 35219 35689
rect 35161 35649 35173 35683
rect 35207 35680 35219 35683
rect 35250 35680 35256 35692
rect 35207 35652 35256 35680
rect 35207 35649 35219 35652
rect 35161 35643 35219 35649
rect 35250 35640 35256 35652
rect 35308 35640 35314 35692
rect 34885 35615 34943 35621
rect 34885 35581 34897 35615
rect 34931 35612 34943 35615
rect 35434 35612 35440 35624
rect 34931 35584 35440 35612
rect 34931 35581 34943 35584
rect 34885 35575 34943 35581
rect 35434 35572 35440 35584
rect 35492 35572 35498 35624
rect 32048 35516 32168 35544
rect 32048 35488 32076 35516
rect 30834 35476 30840 35488
rect 29840 35448 30840 35476
rect 30834 35436 30840 35448
rect 30892 35436 30898 35488
rect 31294 35476 31300 35488
rect 31255 35448 31300 35476
rect 31294 35436 31300 35448
rect 31352 35436 31358 35488
rect 32030 35436 32036 35488
rect 32088 35436 32094 35488
rect 1104 35386 39836 35408
rect 1104 35334 19606 35386
rect 19658 35334 19670 35386
rect 19722 35334 19734 35386
rect 19786 35334 19798 35386
rect 19850 35334 39836 35386
rect 1104 35312 39836 35334
rect 4062 35232 4068 35284
rect 4120 35272 4126 35284
rect 10410 35272 10416 35284
rect 4120 35244 9904 35272
rect 10371 35244 10416 35272
rect 4120 35232 4126 35244
rect 9769 35207 9827 35213
rect 9769 35204 9781 35207
rect 8404 35176 9781 35204
rect 3602 35096 3608 35148
rect 3660 35136 3666 35148
rect 4065 35139 4123 35145
rect 4065 35136 4077 35139
rect 3660 35108 4077 35136
rect 3660 35096 3666 35108
rect 4065 35105 4077 35108
rect 4111 35105 4123 35139
rect 4065 35099 4123 35105
rect 4341 35139 4399 35145
rect 4341 35105 4353 35139
rect 4387 35136 4399 35139
rect 4614 35136 4620 35148
rect 4387 35108 4620 35136
rect 4387 35105 4399 35108
rect 4341 35099 4399 35105
rect 4614 35096 4620 35108
rect 4672 35096 4678 35148
rect 6178 35136 6184 35148
rect 6139 35108 6184 35136
rect 6178 35096 6184 35108
rect 6236 35096 6242 35148
rect 6270 35096 6276 35148
rect 6328 35136 6334 35148
rect 7377 35139 7435 35145
rect 7377 35136 7389 35139
rect 6328 35108 7389 35136
rect 6328 35096 6334 35108
rect 7377 35105 7389 35108
rect 7423 35105 7435 35139
rect 7377 35099 7435 35105
rect 7650 35096 7656 35148
rect 7708 35136 7714 35148
rect 8404 35145 8432 35176
rect 9769 35173 9781 35176
rect 9815 35173 9827 35207
rect 9876 35204 9904 35244
rect 10410 35232 10416 35244
rect 10468 35232 10474 35284
rect 19426 35272 19432 35284
rect 10520 35244 19432 35272
rect 10520 35204 10548 35244
rect 19426 35232 19432 35244
rect 19484 35232 19490 35284
rect 21634 35272 21640 35284
rect 21008 35244 21640 35272
rect 16758 35204 16764 35216
rect 9876 35176 10548 35204
rect 15948 35176 16764 35204
rect 9769 35167 9827 35173
rect 7745 35139 7803 35145
rect 7745 35136 7757 35139
rect 7708 35108 7757 35136
rect 7708 35096 7714 35108
rect 7745 35105 7757 35108
rect 7791 35105 7803 35139
rect 7745 35099 7803 35105
rect 8389 35139 8447 35145
rect 8389 35105 8401 35139
rect 8435 35105 8447 35139
rect 9677 35139 9735 35145
rect 9677 35136 9689 35139
rect 8389 35099 8447 35105
rect 8496 35108 9689 35136
rect 4798 35028 4804 35080
rect 4856 35068 4862 35080
rect 4856 35040 6408 35068
rect 4856 35028 4862 35040
rect 6380 35009 6408 35040
rect 7834 35028 7840 35080
rect 7892 35068 7898 35080
rect 8496 35068 8524 35108
rect 9677 35105 9689 35108
rect 9723 35105 9735 35139
rect 9677 35099 9735 35105
rect 10321 35139 10379 35145
rect 10321 35105 10333 35139
rect 10367 35105 10379 35139
rect 11238 35136 11244 35148
rect 11199 35108 11244 35136
rect 10321 35099 10379 35105
rect 7892 35040 8524 35068
rect 8573 35071 8631 35077
rect 7892 35028 7898 35040
rect 8573 35037 8585 35071
rect 8619 35068 8631 35071
rect 10336 35068 10364 35099
rect 11238 35096 11244 35108
rect 11296 35096 11302 35148
rect 11330 35096 11336 35148
rect 11388 35136 11394 35148
rect 13081 35139 13139 35145
rect 13081 35136 13093 35139
rect 11388 35108 13093 35136
rect 11388 35096 11394 35108
rect 13081 35105 13093 35108
rect 13127 35105 13139 35139
rect 13630 35136 13636 35148
rect 13591 35108 13636 35136
rect 13081 35099 13139 35105
rect 13630 35096 13636 35108
rect 13688 35096 13694 35148
rect 15948 35145 15976 35176
rect 16758 35164 16764 35176
rect 16816 35164 16822 35216
rect 20898 35204 20904 35216
rect 20811 35176 20904 35204
rect 20898 35164 20904 35176
rect 20956 35204 20962 35216
rect 21008 35204 21036 35244
rect 21634 35232 21640 35244
rect 21692 35232 21698 35284
rect 22097 35275 22155 35281
rect 22097 35241 22109 35275
rect 22143 35272 22155 35275
rect 22462 35272 22468 35284
rect 22143 35244 22468 35272
rect 22143 35241 22155 35244
rect 22097 35235 22155 35241
rect 22462 35232 22468 35244
rect 22520 35232 22526 35284
rect 27430 35232 27436 35284
rect 27488 35272 27494 35284
rect 27801 35275 27859 35281
rect 27801 35272 27813 35275
rect 27488 35244 27813 35272
rect 27488 35232 27494 35244
rect 27801 35241 27813 35244
rect 27847 35241 27859 35275
rect 27801 35235 27859 35241
rect 30282 35232 30288 35284
rect 30340 35272 30346 35284
rect 35621 35275 35679 35281
rect 35621 35272 35633 35275
rect 30340 35244 35633 35272
rect 30340 35232 30346 35244
rect 35621 35241 35633 35244
rect 35667 35241 35679 35275
rect 35621 35235 35679 35241
rect 21266 35204 21272 35216
rect 20956 35176 21036 35204
rect 21227 35176 21272 35204
rect 20956 35164 20962 35176
rect 21266 35164 21272 35176
rect 21324 35204 21330 35216
rect 22002 35204 22008 35216
rect 21324 35176 22008 35204
rect 21324 35164 21330 35176
rect 22002 35164 22008 35176
rect 22060 35164 22066 35216
rect 25866 35204 25872 35216
rect 23676 35176 25872 35204
rect 15105 35139 15163 35145
rect 15105 35105 15117 35139
rect 15151 35105 15163 35139
rect 15105 35099 15163 35105
rect 15933 35139 15991 35145
rect 15933 35105 15945 35139
rect 15979 35105 15991 35139
rect 16114 35136 16120 35148
rect 16075 35108 16120 35136
rect 15933 35099 15991 35105
rect 10962 35068 10968 35080
rect 8619 35040 10364 35068
rect 10875 35040 10968 35068
rect 8619 35037 8631 35040
rect 8573 35031 8631 35037
rect 10962 35028 10968 35040
rect 11020 35068 11026 35080
rect 11020 35040 14964 35068
rect 11020 35028 11026 35040
rect 6365 35003 6423 35009
rect 6365 34969 6377 35003
rect 6411 35000 6423 35003
rect 6822 35000 6828 35012
rect 6411 34972 6828 35000
rect 6411 34969 6423 34972
rect 6365 34963 6423 34969
rect 6822 34960 6828 34972
rect 6880 34960 6886 35012
rect 5629 34935 5687 34941
rect 5629 34901 5641 34935
rect 5675 34932 5687 34935
rect 6454 34932 6460 34944
rect 5675 34904 6460 34932
rect 5675 34901 5687 34904
rect 5629 34895 5687 34901
rect 6454 34892 6460 34904
rect 6512 34892 6518 34944
rect 12526 34932 12532 34944
rect 12487 34904 12532 34932
rect 12526 34892 12532 34904
rect 12584 34892 12590 34944
rect 12618 34892 12624 34944
rect 12676 34932 12682 34944
rect 14936 34941 14964 35040
rect 15120 35000 15148 35099
rect 16114 35096 16120 35108
rect 16172 35136 16178 35148
rect 16942 35136 16948 35148
rect 16172 35108 16948 35136
rect 16172 35096 16178 35108
rect 16942 35096 16948 35108
rect 17000 35096 17006 35148
rect 18509 35139 18567 35145
rect 18509 35105 18521 35139
rect 18555 35136 18567 35139
rect 18966 35136 18972 35148
rect 18555 35108 18972 35136
rect 18555 35105 18567 35108
rect 18509 35099 18567 35105
rect 18966 35096 18972 35108
rect 19024 35096 19030 35148
rect 19334 35136 19340 35148
rect 19295 35108 19340 35136
rect 19334 35096 19340 35108
rect 19392 35096 19398 35148
rect 19705 35139 19763 35145
rect 19705 35105 19717 35139
rect 19751 35136 19763 35139
rect 20254 35136 20260 35148
rect 19751 35108 20260 35136
rect 19751 35105 19763 35108
rect 19705 35099 19763 35105
rect 20254 35096 20260 35108
rect 20312 35096 20318 35148
rect 20714 35096 20720 35148
rect 20772 35136 20778 35148
rect 21085 35139 21143 35145
rect 21085 35136 21097 35139
rect 20772 35108 21097 35136
rect 20772 35096 20778 35108
rect 21085 35105 21097 35108
rect 21131 35105 21143 35139
rect 21085 35099 21143 35105
rect 21177 35139 21235 35145
rect 21177 35105 21189 35139
rect 21223 35136 21235 35139
rect 21450 35136 21456 35148
rect 21223 35108 21456 35136
rect 21223 35105 21235 35108
rect 21177 35099 21235 35105
rect 21450 35096 21456 35108
rect 21508 35096 21514 35148
rect 22289 35139 22347 35145
rect 22289 35105 22301 35139
rect 22335 35136 22347 35139
rect 22554 35136 22560 35148
rect 22335 35108 22560 35136
rect 22335 35105 22347 35108
rect 22289 35099 22347 35105
rect 22554 35096 22560 35108
rect 22612 35096 22618 35148
rect 22646 35096 22652 35148
rect 22704 35136 22710 35148
rect 22925 35139 22983 35145
rect 22704 35108 22797 35136
rect 22704 35096 22710 35108
rect 22925 35105 22937 35139
rect 22971 35105 22983 35139
rect 23106 35136 23112 35148
rect 23067 35108 23112 35136
rect 22925 35099 22983 35105
rect 16298 35068 16304 35080
rect 16259 35040 16304 35068
rect 16298 35028 16304 35040
rect 16356 35028 16362 35080
rect 16390 35028 16396 35080
rect 16448 35068 16454 35080
rect 16853 35071 16911 35077
rect 16853 35068 16865 35071
rect 16448 35040 16865 35068
rect 16448 35028 16454 35040
rect 16853 35037 16865 35040
rect 16899 35037 16911 35071
rect 17126 35068 17132 35080
rect 17087 35040 17132 35068
rect 16853 35031 16911 35037
rect 17126 35028 17132 35040
rect 17184 35028 17190 35080
rect 20990 35028 20996 35080
rect 21048 35068 21054 35080
rect 21637 35071 21695 35077
rect 21637 35068 21649 35071
rect 21048 35040 21649 35068
rect 21048 35028 21054 35040
rect 21637 35037 21649 35040
rect 21683 35037 21695 35071
rect 21637 35031 21695 35037
rect 16574 35000 16580 35012
rect 15120 34972 16580 35000
rect 16574 34960 16580 34972
rect 16632 34960 16638 35012
rect 22664 35000 22692 35096
rect 22830 35068 22836 35080
rect 22791 35040 22836 35068
rect 22830 35028 22836 35040
rect 22888 35028 22894 35080
rect 22940 35068 22968 35099
rect 23106 35096 23112 35108
rect 23164 35096 23170 35148
rect 23198 35096 23204 35148
rect 23256 35136 23262 35148
rect 23676 35145 23704 35176
rect 25866 35164 25872 35176
rect 25924 35164 25930 35216
rect 23661 35139 23719 35145
rect 23661 35136 23673 35139
rect 23256 35108 23673 35136
rect 23256 35096 23262 35108
rect 23661 35105 23673 35108
rect 23707 35105 23719 35139
rect 23661 35099 23719 35105
rect 23750 35096 23756 35148
rect 23808 35136 23814 35148
rect 24305 35139 24363 35145
rect 24305 35136 24317 35139
rect 23808 35108 24317 35136
rect 23808 35096 23814 35108
rect 24305 35105 24317 35108
rect 24351 35105 24363 35139
rect 25498 35136 25504 35148
rect 25459 35108 25504 35136
rect 24305 35099 24363 35105
rect 25498 35096 25504 35108
rect 25556 35096 25562 35148
rect 26602 35136 26608 35148
rect 26563 35108 26608 35136
rect 26602 35096 26608 35108
rect 26660 35096 26666 35148
rect 27614 35136 27620 35148
rect 27575 35108 27620 35136
rect 27614 35096 27620 35108
rect 27672 35096 27678 35148
rect 28445 35139 28503 35145
rect 28445 35105 28457 35139
rect 28491 35136 28503 35139
rect 28718 35136 28724 35148
rect 28491 35108 28724 35136
rect 28491 35105 28503 35108
rect 28445 35099 28503 35105
rect 28718 35096 28724 35108
rect 28776 35096 28782 35148
rect 28905 35139 28963 35145
rect 28905 35105 28917 35139
rect 28951 35136 28963 35139
rect 29641 35139 29699 35145
rect 29641 35136 29653 35139
rect 28951 35108 29653 35136
rect 28951 35105 28963 35108
rect 28905 35099 28963 35105
rect 29641 35105 29653 35108
rect 29687 35105 29699 35139
rect 29641 35099 29699 35105
rect 29730 35096 29736 35148
rect 29788 35136 29794 35148
rect 31941 35139 31999 35145
rect 31941 35136 31953 35139
rect 29788 35108 31953 35136
rect 29788 35096 29794 35108
rect 31941 35105 31953 35108
rect 31987 35105 31999 35139
rect 31941 35099 31999 35105
rect 32401 35139 32459 35145
rect 32401 35105 32413 35139
rect 32447 35136 32459 35139
rect 34146 35136 34152 35148
rect 32447 35108 34152 35136
rect 32447 35105 32459 35108
rect 32401 35099 32459 35105
rect 34146 35096 34152 35108
rect 34204 35096 34210 35148
rect 34514 35136 34520 35148
rect 34475 35108 34520 35136
rect 34514 35096 34520 35108
rect 34572 35096 34578 35148
rect 37918 35096 37924 35148
rect 37976 35136 37982 35148
rect 38013 35139 38071 35145
rect 38013 35136 38025 35139
rect 37976 35108 38025 35136
rect 37976 35096 37982 35108
rect 38013 35105 38025 35108
rect 38059 35105 38071 35139
rect 38194 35136 38200 35148
rect 38155 35108 38200 35136
rect 38013 35099 38071 35105
rect 38194 35096 38200 35108
rect 38252 35096 38258 35148
rect 23382 35068 23388 35080
rect 22940 35040 23388 35068
rect 23382 35028 23388 35040
rect 23440 35028 23446 35080
rect 25406 35068 25412 35080
rect 25367 35040 25412 35068
rect 25406 35028 25412 35040
rect 25464 35028 25470 35080
rect 25958 35068 25964 35080
rect 25919 35040 25964 35068
rect 25958 35028 25964 35040
rect 26016 35028 26022 35080
rect 26513 35071 26571 35077
rect 26513 35037 26525 35071
rect 26559 35068 26571 35071
rect 27430 35068 27436 35080
rect 26559 35040 27436 35068
rect 26559 35037 26571 35040
rect 26513 35031 26571 35037
rect 27430 35028 27436 35040
rect 27488 35028 27494 35080
rect 28353 35071 28411 35077
rect 28353 35037 28365 35071
rect 28399 35068 28411 35071
rect 29270 35068 29276 35080
rect 28399 35040 29276 35068
rect 28399 35037 28411 35040
rect 28353 35031 28411 35037
rect 29270 35028 29276 35040
rect 29328 35028 29334 35080
rect 29362 35028 29368 35080
rect 29420 35068 29426 35080
rect 32030 35068 32036 35080
rect 29420 35040 29465 35068
rect 31772 35040 32036 35068
rect 29420 35028 29426 35040
rect 23566 35000 23572 35012
rect 22664 34972 23572 35000
rect 23566 34960 23572 34972
rect 23624 35000 23630 35012
rect 31772 35009 31800 35040
rect 32030 35028 32036 35040
rect 32088 35068 32094 35080
rect 32125 35071 32183 35077
rect 32125 35068 32137 35071
rect 32088 35040 32137 35068
rect 32088 35028 32094 35040
rect 32125 35037 32137 35040
rect 32171 35068 32183 35071
rect 32858 35068 32864 35080
rect 32171 35040 32864 35068
rect 32171 35037 32183 35040
rect 32125 35031 32183 35037
rect 32858 35028 32864 35040
rect 32916 35068 32922 35080
rect 34241 35071 34299 35077
rect 34241 35068 34253 35071
rect 32916 35040 34253 35068
rect 32916 35028 32922 35040
rect 34241 35037 34253 35040
rect 34287 35068 34299 35071
rect 35434 35068 35440 35080
rect 34287 35040 35440 35068
rect 34287 35037 34299 35040
rect 34241 35031 34299 35037
rect 35434 35028 35440 35040
rect 35492 35028 35498 35080
rect 24397 35003 24455 35009
rect 24397 35000 24409 35003
rect 23624 34972 24409 35000
rect 23624 34960 23630 34972
rect 24397 34969 24409 34972
rect 24443 34969 24455 35003
rect 24397 34963 24455 34969
rect 31757 35003 31815 35009
rect 31757 34969 31769 35003
rect 31803 34969 31815 35003
rect 31757 34963 31815 34969
rect 13173 34935 13231 34941
rect 13173 34932 13185 34935
rect 12676 34904 13185 34932
rect 12676 34892 12682 34904
rect 13173 34901 13185 34904
rect 13219 34901 13231 34935
rect 13173 34895 13231 34901
rect 14921 34935 14979 34941
rect 14921 34901 14933 34935
rect 14967 34932 14979 34935
rect 16206 34932 16212 34944
rect 14967 34904 16212 34932
rect 14967 34901 14979 34904
rect 14921 34895 14979 34901
rect 16206 34892 16212 34904
rect 16264 34892 16270 34944
rect 26786 34932 26792 34944
rect 26747 34904 26792 34932
rect 26786 34892 26792 34904
rect 26844 34892 26850 34944
rect 30926 34932 30932 34944
rect 30887 34904 30932 34932
rect 30926 34892 30932 34904
rect 30984 34892 30990 34944
rect 33226 34892 33232 34944
rect 33284 34932 33290 34944
rect 33505 34935 33563 34941
rect 33505 34932 33517 34935
rect 33284 34904 33517 34932
rect 33284 34892 33290 34904
rect 33505 34901 33517 34904
rect 33551 34901 33563 34935
rect 33505 34895 33563 34901
rect 38102 34892 38108 34944
rect 38160 34932 38166 34944
rect 38289 34935 38347 34941
rect 38289 34932 38301 34935
rect 38160 34904 38301 34932
rect 38160 34892 38166 34904
rect 38289 34901 38301 34904
rect 38335 34901 38347 34935
rect 38289 34895 38347 34901
rect 1104 34842 39836 34864
rect 1104 34790 4246 34842
rect 4298 34790 4310 34842
rect 4362 34790 4374 34842
rect 4426 34790 4438 34842
rect 4490 34790 34966 34842
rect 35018 34790 35030 34842
rect 35082 34790 35094 34842
rect 35146 34790 35158 34842
rect 35210 34790 39836 34842
rect 1104 34768 39836 34790
rect 14461 34731 14519 34737
rect 14461 34697 14473 34731
rect 14507 34728 14519 34731
rect 16114 34728 16120 34740
rect 14507 34700 16120 34728
rect 14507 34697 14519 34700
rect 14461 34691 14519 34697
rect 16114 34688 16120 34700
rect 16172 34688 16178 34740
rect 16758 34688 16764 34740
rect 16816 34728 16822 34740
rect 17037 34731 17095 34737
rect 17037 34728 17049 34731
rect 16816 34700 17049 34728
rect 16816 34688 16822 34700
rect 17037 34697 17049 34700
rect 17083 34697 17095 34731
rect 17037 34691 17095 34697
rect 19426 34688 19432 34740
rect 19484 34728 19490 34740
rect 19484 34700 24532 34728
rect 19484 34688 19490 34700
rect 5074 34620 5080 34672
rect 5132 34660 5138 34672
rect 5258 34660 5264 34672
rect 5132 34632 5264 34660
rect 5132 34620 5138 34632
rect 5258 34620 5264 34632
rect 5316 34660 5322 34672
rect 7742 34660 7748 34672
rect 5316 34632 7748 34660
rect 5316 34620 5322 34632
rect 3881 34527 3939 34533
rect 3881 34493 3893 34527
rect 3927 34524 3939 34527
rect 4706 34524 4712 34536
rect 3927 34496 4712 34524
rect 3927 34493 3939 34496
rect 3881 34487 3939 34493
rect 4706 34484 4712 34496
rect 4764 34484 4770 34536
rect 4798 34484 4804 34536
rect 4856 34524 4862 34536
rect 5736 34533 5764 34632
rect 7742 34620 7748 34632
rect 7800 34620 7806 34672
rect 16022 34620 16028 34672
rect 16080 34660 16086 34672
rect 16482 34660 16488 34672
rect 16080 34632 16488 34660
rect 16080 34620 16086 34632
rect 16482 34620 16488 34632
rect 16540 34620 16546 34672
rect 23382 34660 23388 34672
rect 21928 34632 23388 34660
rect 6270 34592 6276 34604
rect 6231 34564 6276 34592
rect 6270 34552 6276 34564
rect 6328 34552 6334 34604
rect 7098 34592 7104 34604
rect 6656 34564 7104 34592
rect 5169 34527 5227 34533
rect 5169 34524 5181 34527
rect 4856 34496 5181 34524
rect 4856 34484 4862 34496
rect 5169 34493 5181 34496
rect 5215 34493 5227 34527
rect 5169 34487 5227 34493
rect 5721 34527 5779 34533
rect 5721 34493 5733 34527
rect 5767 34493 5779 34527
rect 5721 34487 5779 34493
rect 6089 34527 6147 34533
rect 6089 34493 6101 34527
rect 6135 34524 6147 34527
rect 6656 34524 6684 34564
rect 7098 34552 7104 34564
rect 7156 34592 7162 34604
rect 9217 34595 9275 34601
rect 7156 34564 7328 34592
rect 7156 34552 7162 34564
rect 6822 34524 6828 34536
rect 6135 34496 6684 34524
rect 6783 34496 6828 34524
rect 6135 34493 6147 34496
rect 6089 34487 6147 34493
rect 6822 34484 6828 34496
rect 6880 34484 6886 34536
rect 7300 34533 7328 34564
rect 9217 34561 9229 34595
rect 9263 34592 9275 34595
rect 10962 34592 10968 34604
rect 9263 34564 10968 34592
rect 9263 34561 9275 34564
rect 9217 34555 9275 34561
rect 10962 34552 10968 34564
rect 11020 34552 11026 34604
rect 14918 34592 14924 34604
rect 13372 34564 14924 34592
rect 7285 34527 7343 34533
rect 7285 34493 7297 34527
rect 7331 34493 7343 34527
rect 7650 34524 7656 34536
rect 7611 34496 7656 34524
rect 7285 34487 7343 34493
rect 7650 34484 7656 34496
rect 7708 34484 7714 34536
rect 7742 34484 7748 34536
rect 7800 34524 7806 34536
rect 8021 34527 8079 34533
rect 8021 34524 8033 34527
rect 7800 34496 8033 34524
rect 7800 34484 7806 34496
rect 8021 34493 8033 34496
rect 8067 34493 8079 34527
rect 9490 34524 9496 34536
rect 9451 34496 9496 34524
rect 8021 34487 8079 34493
rect 9490 34484 9496 34496
rect 9548 34484 9554 34536
rect 10873 34527 10931 34533
rect 10873 34493 10885 34527
rect 10919 34524 10931 34527
rect 11330 34524 11336 34536
rect 10919 34496 11336 34524
rect 10919 34493 10931 34496
rect 10873 34487 10931 34493
rect 11330 34484 11336 34496
rect 11388 34484 11394 34536
rect 12437 34527 12495 34533
rect 12437 34493 12449 34527
rect 12483 34524 12495 34527
rect 12618 34524 12624 34536
rect 12483 34496 12624 34524
rect 12483 34493 12495 34496
rect 12437 34487 12495 34493
rect 12618 34484 12624 34496
rect 12676 34484 12682 34536
rect 13372 34533 13400 34564
rect 14918 34552 14924 34564
rect 14976 34592 14982 34604
rect 15286 34592 15292 34604
rect 14976 34564 15056 34592
rect 15247 34564 15292 34592
rect 14976 34552 14982 34564
rect 13357 34527 13415 34533
rect 13357 34493 13369 34527
rect 13403 34493 13415 34527
rect 13357 34487 13415 34493
rect 13449 34527 13507 34533
rect 13449 34493 13461 34527
rect 13495 34493 13507 34527
rect 13814 34524 13820 34536
rect 13775 34496 13820 34524
rect 13449 34487 13507 34493
rect 12529 34459 12587 34465
rect 12529 34425 12541 34459
rect 12575 34456 12587 34459
rect 12710 34456 12716 34468
rect 12575 34428 12716 34456
rect 12575 34425 12587 34428
rect 12529 34419 12587 34425
rect 12710 34416 12716 34428
rect 12768 34456 12774 34468
rect 13464 34456 13492 34487
rect 13814 34484 13820 34496
rect 13872 34484 13878 34536
rect 14366 34524 14372 34536
rect 14327 34496 14372 34524
rect 14366 34484 14372 34496
rect 14424 34484 14430 34536
rect 15028 34533 15056 34564
rect 15286 34552 15292 34564
rect 15344 34552 15350 34604
rect 15562 34552 15568 34604
rect 15620 34592 15626 34604
rect 18966 34592 18972 34604
rect 15620 34564 18972 34592
rect 15620 34552 15626 34564
rect 15672 34533 15700 34564
rect 15013 34527 15071 34533
rect 15013 34493 15025 34527
rect 15059 34493 15071 34527
rect 15013 34487 15071 34493
rect 15657 34527 15715 34533
rect 15657 34493 15669 34527
rect 15703 34493 15715 34527
rect 15838 34524 15844 34536
rect 15799 34496 15844 34524
rect 15657 34487 15715 34493
rect 15838 34484 15844 34496
rect 15896 34484 15902 34536
rect 16482 34524 16488 34536
rect 16443 34496 16488 34524
rect 16482 34484 16488 34496
rect 16540 34484 16546 34536
rect 16960 34533 16988 34564
rect 18966 34552 18972 34564
rect 19024 34552 19030 34604
rect 19245 34595 19303 34601
rect 19245 34561 19257 34595
rect 19291 34592 19303 34595
rect 20990 34592 20996 34604
rect 19291 34564 20996 34592
rect 19291 34561 19303 34564
rect 19245 34555 19303 34561
rect 20990 34552 20996 34564
rect 21048 34552 21054 34604
rect 16945 34527 17003 34533
rect 16945 34493 16957 34527
rect 16991 34493 17003 34527
rect 18322 34524 18328 34536
rect 18283 34496 18328 34524
rect 16945 34487 17003 34493
rect 18322 34484 18328 34496
rect 18380 34484 18386 34536
rect 19153 34527 19211 34533
rect 19153 34493 19165 34527
rect 19199 34524 19211 34527
rect 20073 34527 20131 34533
rect 19199 34496 19380 34524
rect 19199 34493 19211 34496
rect 19153 34487 19211 34493
rect 12768 34428 13492 34456
rect 12768 34416 12774 34428
rect 3326 34348 3332 34400
rect 3384 34388 3390 34400
rect 4065 34391 4123 34397
rect 4065 34388 4077 34391
rect 3384 34360 4077 34388
rect 3384 34348 3390 34360
rect 4065 34357 4077 34360
rect 4111 34357 4123 34391
rect 6914 34388 6920 34400
rect 6875 34360 6920 34388
rect 4065 34351 4123 34357
rect 6914 34348 6920 34360
rect 6972 34348 6978 34400
rect 11517 34391 11575 34397
rect 11517 34357 11529 34391
rect 11563 34388 11575 34391
rect 11698 34388 11704 34400
rect 11563 34360 11704 34388
rect 11563 34357 11575 34360
rect 11517 34351 11575 34357
rect 11698 34348 11704 34360
rect 11756 34348 11762 34400
rect 18601 34391 18659 34397
rect 18601 34357 18613 34391
rect 18647 34388 18659 34391
rect 18690 34388 18696 34400
rect 18647 34360 18696 34388
rect 18647 34357 18659 34360
rect 18601 34351 18659 34357
rect 18690 34348 18696 34360
rect 18748 34348 18754 34400
rect 19352 34388 19380 34496
rect 20073 34493 20085 34527
rect 20119 34493 20131 34527
rect 20530 34524 20536 34536
rect 20491 34496 20536 34524
rect 20073 34487 20131 34493
rect 20088 34456 20116 34487
rect 20530 34484 20536 34496
rect 20588 34484 20594 34536
rect 20901 34527 20959 34533
rect 20901 34493 20913 34527
rect 20947 34524 20959 34527
rect 21450 34524 21456 34536
rect 20947 34496 21456 34524
rect 20947 34493 20959 34496
rect 20901 34487 20959 34493
rect 21450 34484 21456 34496
rect 21508 34524 21514 34536
rect 21928 34533 21956 34632
rect 23382 34620 23388 34632
rect 23440 34620 23446 34672
rect 23845 34663 23903 34669
rect 23845 34629 23857 34663
rect 23891 34629 23903 34663
rect 23845 34623 23903 34629
rect 23860 34592 23888 34623
rect 22204 34564 23888 34592
rect 21913 34527 21971 34533
rect 21913 34524 21925 34527
rect 21508 34496 21925 34524
rect 21508 34484 21514 34496
rect 21913 34493 21925 34496
rect 21959 34493 21971 34527
rect 21913 34487 21971 34493
rect 22005 34527 22063 34533
rect 22005 34493 22017 34527
rect 22051 34524 22063 34527
rect 22051 34496 22085 34524
rect 22051 34493 22063 34496
rect 22005 34487 22063 34493
rect 20162 34456 20168 34468
rect 20088 34428 20168 34456
rect 20162 34416 20168 34428
rect 20220 34456 20226 34468
rect 20622 34456 20628 34468
rect 20220 34428 20628 34456
rect 20220 34416 20226 34428
rect 20622 34416 20628 34428
rect 20680 34456 20686 34468
rect 22020 34456 22048 34487
rect 22094 34456 22100 34468
rect 20680 34428 22100 34456
rect 20680 34416 20686 34428
rect 22094 34416 22100 34428
rect 22152 34416 22158 34468
rect 19981 34391 20039 34397
rect 19981 34388 19993 34391
rect 19352 34360 19993 34388
rect 19981 34357 19993 34360
rect 20027 34357 20039 34391
rect 19981 34351 20039 34357
rect 21542 34348 21548 34400
rect 21600 34388 21606 34400
rect 22204 34388 22232 34564
rect 24302 34552 24308 34604
rect 24360 34592 24366 34604
rect 24397 34595 24455 34601
rect 24397 34592 24409 34595
rect 24360 34564 24409 34592
rect 24360 34552 24366 34564
rect 24397 34561 24409 34564
rect 24443 34561 24455 34595
rect 24397 34555 24455 34561
rect 22649 34527 22707 34533
rect 22649 34493 22661 34527
rect 22695 34493 22707 34527
rect 22830 34524 22836 34536
rect 22791 34496 22836 34524
rect 22649 34487 22707 34493
rect 22664 34456 22692 34487
rect 22830 34484 22836 34496
rect 22888 34484 22894 34536
rect 23109 34527 23167 34533
rect 23109 34493 23121 34527
rect 23155 34524 23167 34527
rect 23474 34524 23480 34536
rect 23155 34496 23480 34524
rect 23155 34493 23167 34496
rect 23109 34487 23167 34493
rect 23474 34484 23480 34496
rect 23532 34484 23538 34536
rect 23658 34524 23664 34536
rect 23619 34496 23664 34524
rect 23658 34484 23664 34496
rect 23716 34484 23722 34536
rect 23014 34456 23020 34468
rect 22664 34428 23020 34456
rect 23014 34416 23020 34428
rect 23072 34416 23078 34468
rect 24412 34456 24440 34555
rect 24504 34533 24532 34700
rect 25682 34688 25688 34740
rect 25740 34728 25746 34740
rect 27709 34731 27767 34737
rect 27709 34728 27721 34731
rect 25740 34700 27721 34728
rect 25740 34688 25746 34700
rect 27709 34697 27721 34700
rect 27755 34697 27767 34731
rect 27709 34691 27767 34697
rect 30101 34731 30159 34737
rect 30101 34697 30113 34731
rect 30147 34728 30159 34731
rect 30190 34728 30196 34740
rect 30147 34700 30196 34728
rect 30147 34697 30159 34700
rect 30101 34691 30159 34697
rect 30190 34688 30196 34700
rect 30248 34688 30254 34740
rect 28442 34620 28448 34672
rect 28500 34660 28506 34672
rect 28629 34663 28687 34669
rect 28629 34660 28641 34663
rect 28500 34632 28641 34660
rect 28500 34620 28506 34632
rect 28629 34629 28641 34632
rect 28675 34660 28687 34663
rect 31021 34663 31079 34669
rect 28675 34632 30880 34660
rect 28675 34629 28687 34632
rect 28629 34623 28687 34629
rect 24949 34595 25007 34601
rect 24949 34561 24961 34595
rect 24995 34592 25007 34595
rect 25038 34592 25044 34604
rect 24995 34564 25044 34592
rect 24995 34561 25007 34564
rect 24949 34555 25007 34561
rect 25038 34552 25044 34564
rect 25096 34552 25102 34604
rect 25958 34552 25964 34604
rect 26016 34592 26022 34604
rect 26605 34595 26663 34601
rect 26605 34592 26617 34595
rect 26016 34564 26617 34592
rect 26016 34552 26022 34564
rect 26605 34561 26617 34564
rect 26651 34561 26663 34595
rect 26605 34555 26663 34561
rect 29270 34552 29276 34604
rect 29328 34592 29334 34604
rect 29822 34592 29828 34604
rect 29328 34564 29828 34592
rect 29328 34552 29334 34564
rect 29822 34552 29828 34564
rect 29880 34552 29886 34604
rect 24489 34527 24547 34533
rect 24489 34493 24501 34527
rect 24535 34493 24547 34527
rect 26326 34524 26332 34536
rect 26287 34496 26332 34524
rect 24489 34487 24547 34493
rect 26326 34484 26332 34496
rect 26384 34484 26390 34536
rect 28445 34527 28503 34533
rect 28445 34493 28457 34527
rect 28491 34524 28503 34527
rect 28718 34524 28724 34536
rect 28491 34496 28724 34524
rect 28491 34493 28503 34496
rect 28445 34487 28503 34493
rect 28718 34484 28724 34496
rect 28776 34484 28782 34536
rect 29917 34527 29975 34533
rect 29917 34493 29929 34527
rect 29963 34524 29975 34527
rect 30650 34524 30656 34536
rect 29963 34496 30656 34524
rect 29963 34493 29975 34496
rect 29917 34487 29975 34493
rect 30650 34484 30656 34496
rect 30708 34484 30714 34536
rect 30852 34533 30880 34632
rect 31021 34629 31033 34663
rect 31067 34660 31079 34663
rect 31202 34660 31208 34672
rect 31067 34632 31208 34660
rect 31067 34629 31079 34632
rect 31021 34623 31079 34629
rect 31202 34620 31208 34632
rect 31260 34620 31266 34672
rect 31941 34595 31999 34601
rect 31941 34561 31953 34595
rect 31987 34592 31999 34595
rect 32490 34592 32496 34604
rect 31987 34564 32496 34592
rect 31987 34561 31999 34564
rect 31941 34555 31999 34561
rect 32490 34552 32496 34564
rect 32548 34552 32554 34604
rect 34054 34592 34060 34604
rect 32968 34564 34060 34592
rect 30837 34527 30895 34533
rect 30837 34493 30849 34527
rect 30883 34493 30895 34527
rect 31573 34527 31631 34533
rect 31573 34524 31585 34527
rect 30837 34487 30895 34493
rect 30944 34496 31585 34524
rect 26234 34456 26240 34468
rect 24412 34428 26240 34456
rect 26234 34416 26240 34428
rect 26292 34416 26298 34468
rect 30190 34416 30196 34468
rect 30248 34456 30254 34468
rect 30944 34456 30972 34496
rect 31573 34493 31585 34496
rect 31619 34493 31631 34527
rect 32214 34524 32220 34536
rect 32175 34496 32220 34524
rect 31573 34487 31631 34493
rect 32214 34484 32220 34496
rect 32272 34484 32278 34536
rect 32968 34533 32996 34564
rect 34054 34552 34060 34564
rect 34112 34552 34118 34604
rect 35434 34552 35440 34604
rect 35492 34592 35498 34604
rect 37093 34595 37151 34601
rect 37093 34592 37105 34595
rect 35492 34564 37105 34592
rect 35492 34552 35498 34564
rect 37093 34561 37105 34564
rect 37139 34561 37151 34595
rect 37093 34555 37151 34561
rect 38010 34552 38016 34604
rect 38068 34592 38074 34604
rect 38194 34592 38200 34604
rect 38068 34564 38200 34592
rect 38068 34552 38074 34564
rect 38194 34552 38200 34564
rect 38252 34592 38258 34604
rect 38473 34595 38531 34601
rect 38473 34592 38485 34595
rect 38252 34564 38485 34592
rect 38252 34552 38258 34564
rect 38473 34561 38485 34564
rect 38519 34561 38531 34595
rect 38473 34555 38531 34561
rect 32953 34527 33011 34533
rect 32953 34493 32965 34527
rect 32999 34493 33011 34527
rect 33134 34524 33140 34536
rect 33095 34496 33140 34524
rect 32953 34487 33011 34493
rect 33134 34484 33140 34496
rect 33192 34484 33198 34536
rect 33318 34524 33324 34536
rect 33279 34496 33324 34524
rect 33318 34484 33324 34496
rect 33376 34484 33382 34536
rect 35345 34527 35403 34533
rect 35345 34493 35357 34527
rect 35391 34493 35403 34527
rect 36078 34524 36084 34536
rect 36039 34496 36084 34524
rect 35345 34487 35403 34493
rect 30248 34428 30972 34456
rect 30248 34416 30254 34428
rect 35360 34400 35388 34487
rect 36078 34484 36084 34496
rect 36136 34484 36142 34536
rect 36354 34524 36360 34536
rect 36315 34496 36360 34524
rect 36354 34484 36360 34496
rect 36412 34484 36418 34536
rect 37366 34524 37372 34536
rect 37327 34496 37372 34524
rect 37366 34484 37372 34496
rect 37424 34484 37430 34536
rect 21600 34360 22232 34388
rect 21600 34348 21606 34360
rect 35342 34348 35348 34400
rect 35400 34348 35406 34400
rect 35437 34391 35495 34397
rect 35437 34357 35449 34391
rect 35483 34388 35495 34391
rect 35710 34388 35716 34400
rect 35483 34360 35716 34388
rect 35483 34357 35495 34360
rect 35437 34351 35495 34357
rect 35710 34348 35716 34360
rect 35768 34348 35774 34400
rect 1104 34298 39836 34320
rect 1104 34246 19606 34298
rect 19658 34246 19670 34298
rect 19722 34246 19734 34298
rect 19786 34246 19798 34298
rect 19850 34246 39836 34298
rect 1104 34224 39836 34246
rect 7561 34187 7619 34193
rect 7561 34153 7573 34187
rect 7607 34184 7619 34187
rect 7834 34184 7840 34196
rect 7607 34156 7840 34184
rect 7607 34153 7619 34156
rect 7561 34147 7619 34153
rect 7834 34144 7840 34156
rect 7892 34144 7898 34196
rect 9033 34187 9091 34193
rect 9033 34153 9045 34187
rect 9079 34184 9091 34187
rect 9490 34184 9496 34196
rect 9079 34156 9496 34184
rect 9079 34153 9091 34156
rect 9033 34147 9091 34153
rect 9490 34144 9496 34156
rect 9548 34144 9554 34196
rect 17126 34144 17132 34196
rect 17184 34184 17190 34196
rect 17681 34187 17739 34193
rect 17681 34184 17693 34187
rect 17184 34156 17693 34184
rect 17184 34144 17190 34156
rect 17681 34153 17693 34156
rect 17727 34153 17739 34187
rect 17681 34147 17739 34153
rect 23842 34144 23848 34196
rect 23900 34184 23906 34196
rect 24029 34187 24087 34193
rect 24029 34184 24041 34187
rect 23900 34156 24041 34184
rect 23900 34144 23906 34156
rect 24029 34153 24041 34156
rect 24075 34184 24087 34187
rect 28902 34184 28908 34196
rect 24075 34156 28908 34184
rect 24075 34153 24087 34156
rect 24029 34147 24087 34153
rect 28902 34144 28908 34156
rect 28960 34144 28966 34196
rect 37366 34144 37372 34196
rect 37424 34184 37430 34196
rect 37829 34187 37887 34193
rect 37829 34184 37841 34187
rect 37424 34156 37841 34184
rect 37424 34144 37430 34156
rect 37829 34153 37841 34156
rect 37875 34153 37887 34187
rect 37829 34147 37887 34153
rect 8113 34119 8171 34125
rect 8113 34116 8125 34119
rect 7116 34088 8125 34116
rect 7116 34060 7144 34088
rect 8113 34085 8125 34088
rect 8159 34085 8171 34119
rect 13906 34116 13912 34128
rect 8113 34079 8171 34085
rect 12820 34088 13912 34116
rect 1581 34051 1639 34057
rect 1581 34017 1593 34051
rect 1627 34048 1639 34051
rect 2682 34048 2688 34060
rect 1627 34020 2688 34048
rect 1627 34017 1639 34020
rect 1581 34011 1639 34017
rect 2682 34008 2688 34020
rect 2740 34048 2746 34060
rect 3602 34048 3608 34060
rect 2740 34020 3608 34048
rect 2740 34008 2746 34020
rect 3602 34008 3608 34020
rect 3660 34048 3666 34060
rect 4065 34051 4123 34057
rect 4065 34048 4077 34051
rect 3660 34020 4077 34048
rect 3660 34008 3666 34020
rect 4065 34017 4077 34020
rect 4111 34017 4123 34051
rect 4065 34011 4123 34017
rect 6733 34051 6791 34057
rect 6733 34017 6745 34051
rect 6779 34048 6791 34051
rect 6822 34048 6828 34060
rect 6779 34020 6828 34048
rect 6779 34017 6791 34020
rect 6733 34011 6791 34017
rect 6822 34008 6828 34020
rect 6880 34008 6886 34060
rect 7098 34048 7104 34060
rect 7059 34020 7104 34048
rect 7098 34008 7104 34020
rect 7156 34008 7162 34060
rect 7285 34051 7343 34057
rect 7285 34017 7297 34051
rect 7331 34017 7343 34051
rect 8018 34048 8024 34060
rect 7979 34020 8024 34048
rect 7285 34011 7343 34017
rect 1854 33980 1860 33992
rect 1815 33952 1860 33980
rect 1854 33940 1860 33952
rect 1912 33940 1918 33992
rect 4341 33983 4399 33989
rect 4341 33949 4353 33983
rect 4387 33980 4399 33983
rect 5442 33980 5448 33992
rect 4387 33952 5448 33980
rect 4387 33949 4399 33952
rect 4341 33943 4399 33949
rect 5442 33940 5448 33952
rect 5500 33940 5506 33992
rect 6178 33940 6184 33992
rect 6236 33980 6242 33992
rect 7300 33980 7328 34011
rect 8018 34008 8024 34020
rect 8076 34008 8082 34060
rect 8938 34048 8944 34060
rect 8899 34020 8944 34048
rect 8938 34008 8944 34020
rect 8996 34008 9002 34060
rect 9858 34048 9864 34060
rect 9819 34020 9864 34048
rect 9858 34008 9864 34020
rect 9916 34008 9922 34060
rect 10781 34051 10839 34057
rect 10781 34017 10793 34051
rect 10827 34017 10839 34051
rect 10781 34011 10839 34017
rect 11057 34051 11115 34057
rect 11057 34017 11069 34051
rect 11103 34048 11115 34051
rect 11517 34051 11575 34057
rect 11103 34020 11284 34048
rect 11103 34017 11115 34020
rect 11057 34011 11115 34017
rect 6236 33952 7328 33980
rect 6236 33940 6242 33952
rect 10796 33912 10824 34011
rect 11146 33980 11152 33992
rect 11107 33952 11152 33980
rect 11146 33940 11152 33952
rect 11204 33940 11210 33992
rect 11256 33980 11284 34020
rect 11517 34017 11529 34051
rect 11563 34048 11575 34051
rect 11882 34048 11888 34060
rect 11563 34020 11888 34048
rect 11563 34017 11575 34020
rect 11517 34011 11575 34017
rect 11882 34008 11888 34020
rect 11940 34008 11946 34060
rect 11977 34051 12035 34057
rect 11977 34017 11989 34051
rect 12023 34017 12035 34051
rect 12710 34048 12716 34060
rect 12671 34020 12716 34048
rect 11977 34011 12035 34017
rect 11698 33980 11704 33992
rect 11256 33952 11704 33980
rect 11698 33940 11704 33952
rect 11756 33940 11762 33992
rect 11992 33980 12020 34011
rect 12710 34008 12716 34020
rect 12768 34008 12774 34060
rect 12820 34057 12848 34088
rect 13906 34076 13912 34088
rect 13964 34076 13970 34128
rect 22646 34076 22652 34128
rect 22704 34116 22710 34128
rect 25961 34119 26019 34125
rect 22704 34088 24256 34116
rect 22704 34076 22710 34088
rect 12805 34051 12863 34057
rect 12805 34017 12817 34051
rect 12851 34017 12863 34051
rect 12805 34011 12863 34017
rect 12894 34008 12900 34060
rect 12952 34048 12958 34060
rect 13173 34051 13231 34057
rect 13173 34048 13185 34051
rect 12952 34020 13185 34048
rect 12952 34008 12958 34020
rect 13173 34017 13185 34020
rect 13219 34017 13231 34051
rect 13173 34011 13231 34017
rect 13725 34051 13783 34057
rect 13725 34017 13737 34051
rect 13771 34017 13783 34051
rect 13725 34011 13783 34017
rect 12526 33980 12532 33992
rect 11992 33952 12532 33980
rect 12526 33940 12532 33952
rect 12584 33980 12590 33992
rect 13630 33980 13636 33992
rect 12584 33952 13636 33980
rect 12584 33940 12590 33952
rect 13630 33940 13636 33952
rect 13688 33940 13694 33992
rect 11054 33912 11060 33924
rect 10796 33884 11060 33912
rect 11054 33872 11060 33884
rect 11112 33872 11118 33924
rect 12342 33872 12348 33924
rect 12400 33912 12406 33924
rect 13740 33912 13768 34011
rect 15102 34008 15108 34060
rect 15160 34048 15166 34060
rect 16025 34051 16083 34057
rect 16025 34048 16037 34051
rect 15160 34020 16037 34048
rect 15160 34008 15166 34020
rect 16025 34017 16037 34020
rect 16071 34017 16083 34051
rect 16298 34048 16304 34060
rect 16259 34020 16304 34048
rect 16025 34011 16083 34017
rect 16298 34008 16304 34020
rect 16356 34008 16362 34060
rect 16942 34048 16948 34060
rect 16903 34020 16948 34048
rect 16942 34008 16948 34020
rect 17000 34008 17006 34060
rect 17310 34008 17316 34060
rect 17368 34048 17374 34060
rect 17589 34051 17647 34057
rect 17589 34048 17601 34051
rect 17368 34020 17601 34048
rect 17368 34008 17374 34020
rect 17589 34017 17601 34020
rect 17635 34017 17647 34051
rect 17589 34011 17647 34017
rect 18230 34008 18236 34060
rect 18288 34048 18294 34060
rect 18417 34051 18475 34057
rect 18417 34048 18429 34051
rect 18288 34020 18429 34048
rect 18288 34008 18294 34020
rect 18417 34017 18429 34020
rect 18463 34017 18475 34051
rect 18690 34048 18696 34060
rect 18651 34020 18696 34048
rect 18417 34011 18475 34017
rect 18690 34008 18696 34020
rect 18748 34008 18754 34060
rect 21174 34048 21180 34060
rect 21135 34020 21180 34048
rect 21174 34008 21180 34020
rect 21232 34008 21238 34060
rect 21358 34048 21364 34060
rect 21319 34020 21364 34048
rect 21358 34008 21364 34020
rect 21416 34008 21422 34060
rect 21634 34048 21640 34060
rect 21595 34020 21640 34048
rect 21634 34008 21640 34020
rect 21692 34008 21698 34060
rect 22094 34008 22100 34060
rect 22152 34048 22158 34060
rect 22373 34051 22431 34057
rect 22373 34048 22385 34051
rect 22152 34020 22385 34048
rect 22152 34008 22158 34020
rect 22373 34017 22385 34020
rect 22419 34048 22431 34051
rect 22833 34051 22891 34057
rect 22833 34048 22845 34051
rect 22419 34020 22845 34048
rect 22419 34017 22431 34020
rect 22373 34011 22431 34017
rect 22833 34017 22845 34020
rect 22879 34017 22891 34051
rect 23474 34048 23480 34060
rect 23435 34020 23480 34048
rect 22833 34011 22891 34017
rect 23474 34008 23480 34020
rect 23532 34008 23538 34060
rect 24228 34057 24256 34088
rect 25961 34085 25973 34119
rect 26007 34116 26019 34119
rect 26602 34116 26608 34128
rect 26007 34088 26608 34116
rect 26007 34085 26019 34088
rect 25961 34079 26019 34085
rect 26602 34076 26608 34088
rect 26660 34076 26666 34128
rect 24213 34051 24271 34057
rect 24213 34017 24225 34051
rect 24259 34017 24271 34051
rect 24213 34011 24271 34017
rect 24305 34051 24363 34057
rect 24305 34017 24317 34051
rect 24351 34048 24363 34051
rect 26326 34048 26332 34060
rect 24351 34020 26332 34048
rect 24351 34017 24363 34020
rect 24305 34011 24363 34017
rect 26326 34008 26332 34020
rect 26384 34048 26390 34060
rect 26513 34051 26571 34057
rect 26513 34048 26525 34051
rect 26384 34020 26525 34048
rect 26384 34008 26390 34020
rect 26513 34017 26525 34020
rect 26559 34017 26571 34051
rect 26786 34048 26792 34060
rect 26747 34020 26792 34048
rect 26513 34011 26571 34017
rect 15194 33940 15200 33992
rect 15252 33980 15258 33992
rect 15473 33983 15531 33989
rect 15473 33980 15485 33983
rect 15252 33952 15485 33980
rect 15252 33940 15258 33952
rect 15473 33949 15485 33952
rect 15519 33949 15531 33983
rect 16482 33980 16488 33992
rect 16395 33952 16488 33980
rect 15473 33943 15531 33949
rect 16482 33940 16488 33952
rect 16540 33980 16546 33992
rect 17218 33980 17224 33992
rect 16540 33952 17224 33980
rect 16540 33940 16546 33952
rect 17218 33940 17224 33952
rect 17276 33940 17282 33992
rect 23201 33983 23259 33989
rect 23201 33949 23213 33983
rect 23247 33980 23259 33983
rect 23750 33980 23756 33992
rect 23247 33952 23756 33980
rect 23247 33949 23259 33952
rect 23201 33943 23259 33949
rect 23750 33940 23756 33952
rect 23808 33940 23814 33992
rect 24578 33980 24584 33992
rect 24539 33952 24584 33980
rect 24578 33940 24584 33952
rect 24636 33940 24642 33992
rect 26528 33980 26556 34011
rect 26786 34008 26792 34020
rect 26844 34008 26850 34060
rect 29638 34008 29644 34060
rect 29696 34048 29702 34060
rect 30837 34051 30895 34057
rect 30837 34048 30849 34051
rect 29696 34020 30849 34048
rect 29696 34008 29702 34020
rect 30837 34017 30849 34020
rect 30883 34017 30895 34051
rect 30837 34011 30895 34017
rect 32125 34051 32183 34057
rect 32125 34017 32137 34051
rect 32171 34048 32183 34051
rect 32858 34048 32864 34060
rect 32171 34020 32864 34048
rect 32171 34017 32183 34020
rect 32125 34011 32183 34017
rect 32858 34008 32864 34020
rect 32916 34008 32922 34060
rect 33134 34008 33140 34060
rect 33192 34048 33198 34060
rect 34241 34051 34299 34057
rect 34241 34048 34253 34051
rect 33192 34020 34253 34048
rect 33192 34008 33198 34020
rect 34241 34017 34253 34020
rect 34287 34017 34299 34051
rect 34790 34048 34796 34060
rect 34751 34020 34796 34048
rect 34241 34011 34299 34017
rect 34790 34008 34796 34020
rect 34848 34008 34854 34060
rect 35434 34048 35440 34060
rect 35395 34020 35440 34048
rect 35434 34008 35440 34020
rect 35492 34008 35498 34060
rect 35710 34048 35716 34060
rect 35671 34020 35716 34048
rect 35710 34008 35716 34020
rect 35768 34008 35774 34060
rect 35802 34008 35808 34060
rect 35860 34048 35866 34060
rect 37737 34051 37795 34057
rect 37737 34048 37749 34051
rect 35860 34020 37749 34048
rect 35860 34008 35866 34020
rect 37737 34017 37749 34020
rect 37783 34017 37795 34051
rect 38286 34048 38292 34060
rect 38247 34020 38292 34048
rect 37737 34011 37795 34017
rect 38286 34008 38292 34020
rect 38344 34008 38350 34060
rect 28629 33983 28687 33989
rect 28629 33980 28641 33983
rect 26528 33952 28641 33980
rect 28629 33949 28641 33952
rect 28675 33949 28687 33983
rect 28629 33943 28687 33949
rect 28905 33983 28963 33989
rect 28905 33949 28917 33983
rect 28951 33980 28963 33983
rect 29546 33980 29552 33992
rect 28951 33952 29552 33980
rect 28951 33949 28963 33952
rect 28905 33943 28963 33949
rect 29546 33940 29552 33952
rect 29604 33940 29610 33992
rect 29822 33940 29828 33992
rect 29880 33980 29886 33992
rect 30745 33983 30803 33989
rect 30745 33980 30757 33983
rect 29880 33952 30757 33980
rect 29880 33940 29886 33952
rect 30745 33949 30757 33952
rect 30791 33949 30803 33983
rect 32398 33980 32404 33992
rect 32359 33952 32404 33980
rect 30745 33943 30803 33949
rect 32398 33940 32404 33952
rect 32456 33940 32462 33992
rect 37642 33940 37648 33992
rect 37700 33980 37706 33992
rect 38565 33983 38623 33989
rect 38565 33980 38577 33983
rect 37700 33952 38577 33980
rect 37700 33940 37706 33952
rect 38565 33949 38577 33952
rect 38611 33949 38623 33983
rect 38565 33943 38623 33949
rect 12400 33884 13768 33912
rect 12400 33872 12406 33884
rect 29730 33872 29736 33924
rect 29788 33912 29794 33924
rect 29788 33884 31064 33912
rect 29788 33872 29794 33884
rect 3145 33847 3203 33853
rect 3145 33813 3157 33847
rect 3191 33844 3203 33847
rect 3234 33844 3240 33856
rect 3191 33816 3240 33844
rect 3191 33813 3203 33816
rect 3145 33807 3203 33813
rect 3234 33804 3240 33816
rect 3292 33804 3298 33856
rect 5626 33844 5632 33856
rect 5587 33816 5632 33844
rect 5626 33804 5632 33816
rect 5684 33804 5690 33856
rect 9674 33804 9680 33856
rect 9732 33844 9738 33856
rect 9953 33847 10011 33853
rect 9953 33844 9965 33847
rect 9732 33816 9965 33844
rect 9732 33804 9738 33816
rect 9953 33813 9965 33816
rect 9999 33813 10011 33847
rect 9953 33807 10011 33813
rect 12529 33847 12587 33853
rect 12529 33813 12541 33847
rect 12575 33844 12587 33847
rect 12986 33844 12992 33856
rect 12575 33816 12992 33844
rect 12575 33813 12587 33816
rect 12529 33807 12587 33813
rect 12986 33804 12992 33816
rect 13044 33804 13050 33856
rect 15930 33804 15936 33856
rect 15988 33844 15994 33856
rect 17037 33847 17095 33853
rect 17037 33844 17049 33847
rect 15988 33816 17049 33844
rect 15988 33804 15994 33816
rect 17037 33813 17049 33816
rect 17083 33813 17095 33847
rect 19978 33844 19984 33856
rect 19939 33816 19984 33844
rect 17037 33807 17095 33813
rect 19978 33804 19984 33816
rect 20036 33804 20042 33856
rect 22281 33847 22339 33853
rect 22281 33813 22293 33847
rect 22327 33844 22339 33847
rect 22370 33844 22376 33856
rect 22327 33816 22376 33844
rect 22327 33813 22339 33816
rect 22281 33807 22339 33813
rect 22370 33804 22376 33816
rect 22428 33804 22434 33856
rect 26694 33804 26700 33856
rect 26752 33844 26758 33856
rect 27893 33847 27951 33853
rect 27893 33844 27905 33847
rect 26752 33816 27905 33844
rect 26752 33804 26758 33816
rect 27893 33813 27905 33816
rect 27939 33813 27951 33847
rect 27893 33807 27951 33813
rect 30193 33847 30251 33853
rect 30193 33813 30205 33847
rect 30239 33844 30251 33847
rect 30374 33844 30380 33856
rect 30239 33816 30380 33844
rect 30239 33813 30251 33816
rect 30193 33807 30251 33813
rect 30374 33804 30380 33816
rect 30432 33804 30438 33856
rect 31036 33853 31064 33884
rect 31021 33847 31079 33853
rect 31021 33813 31033 33847
rect 31067 33813 31079 33847
rect 33502 33844 33508 33856
rect 33463 33816 33508 33844
rect 31021 33807 31079 33813
rect 33502 33804 33508 33816
rect 33560 33804 33566 33856
rect 34330 33844 34336 33856
rect 34291 33816 34336 33844
rect 34330 33804 34336 33816
rect 34388 33804 34394 33856
rect 36630 33804 36636 33856
rect 36688 33844 36694 33856
rect 36817 33847 36875 33853
rect 36817 33844 36829 33847
rect 36688 33816 36829 33844
rect 36688 33804 36694 33816
rect 36817 33813 36829 33816
rect 36863 33813 36875 33847
rect 36817 33807 36875 33813
rect 1104 33754 39836 33776
rect 1104 33702 4246 33754
rect 4298 33702 4310 33754
rect 4362 33702 4374 33754
rect 4426 33702 4438 33754
rect 4490 33702 34966 33754
rect 35018 33702 35030 33754
rect 35082 33702 35094 33754
rect 35146 33702 35158 33754
rect 35210 33702 39836 33754
rect 1104 33680 39836 33702
rect 5442 33640 5448 33652
rect 5403 33612 5448 33640
rect 5442 33600 5448 33612
rect 5500 33600 5506 33652
rect 7285 33643 7343 33649
rect 7285 33609 7297 33643
rect 7331 33640 7343 33643
rect 7650 33640 7656 33652
rect 7331 33612 7656 33640
rect 7331 33609 7343 33612
rect 7285 33603 7343 33609
rect 7650 33600 7656 33612
rect 7708 33600 7714 33652
rect 9858 33600 9864 33652
rect 9916 33640 9922 33652
rect 10781 33643 10839 33649
rect 10781 33640 10793 33643
rect 9916 33612 10793 33640
rect 9916 33600 9922 33612
rect 10781 33609 10793 33612
rect 10827 33609 10839 33643
rect 13814 33640 13820 33652
rect 13775 33612 13820 33640
rect 10781 33603 10839 33609
rect 13814 33600 13820 33612
rect 13872 33600 13878 33652
rect 14553 33643 14611 33649
rect 14553 33609 14565 33643
rect 14599 33640 14611 33643
rect 16942 33640 16948 33652
rect 14599 33612 16948 33640
rect 14599 33609 14611 33612
rect 14553 33603 14611 33609
rect 16942 33600 16948 33612
rect 17000 33600 17006 33652
rect 17218 33640 17224 33652
rect 17131 33612 17224 33640
rect 17218 33600 17224 33612
rect 17276 33640 17282 33652
rect 20254 33640 20260 33652
rect 17276 33612 20260 33640
rect 17276 33600 17282 33612
rect 20254 33600 20260 33612
rect 20312 33600 20318 33652
rect 21545 33643 21603 33649
rect 21545 33609 21557 33643
rect 21591 33640 21603 33643
rect 22646 33640 22652 33652
rect 21591 33612 22652 33640
rect 21591 33609 21603 33612
rect 21545 33603 21603 33609
rect 22646 33600 22652 33612
rect 22704 33600 22710 33652
rect 24578 33600 24584 33652
rect 24636 33640 24642 33652
rect 26053 33643 26111 33649
rect 26053 33640 26065 33643
rect 24636 33612 26065 33640
rect 24636 33600 24642 33612
rect 26053 33609 26065 33612
rect 26099 33609 26111 33643
rect 28626 33640 28632 33652
rect 28587 33612 28632 33640
rect 26053 33603 26111 33609
rect 28626 33600 28632 33612
rect 28684 33600 28690 33652
rect 28902 33600 28908 33652
rect 28960 33640 28966 33652
rect 29178 33640 29184 33652
rect 28960 33612 29184 33640
rect 28960 33600 28966 33612
rect 29178 33600 29184 33612
rect 29236 33600 29242 33652
rect 29546 33640 29552 33652
rect 29507 33612 29552 33640
rect 29546 33600 29552 33612
rect 29604 33600 29610 33652
rect 30558 33640 30564 33652
rect 30519 33612 30564 33640
rect 30558 33600 30564 33612
rect 30616 33600 30622 33652
rect 34054 33640 34060 33652
rect 34015 33612 34060 33640
rect 34054 33600 34060 33612
rect 34112 33600 34118 33652
rect 1489 33575 1547 33581
rect 1489 33541 1501 33575
rect 1535 33572 1547 33575
rect 1578 33572 1584 33584
rect 1535 33544 1584 33572
rect 1535 33541 1547 33544
rect 1489 33535 1547 33541
rect 1578 33532 1584 33544
rect 1636 33532 1642 33584
rect 8938 33532 8944 33584
rect 8996 33572 9002 33584
rect 9953 33575 10011 33581
rect 9953 33572 9965 33575
rect 8996 33544 9965 33572
rect 8996 33532 9002 33544
rect 9953 33541 9965 33544
rect 9999 33541 10011 33575
rect 9953 33535 10011 33541
rect 11514 33532 11520 33584
rect 11572 33532 11578 33584
rect 19058 33532 19064 33584
rect 19116 33572 19122 33584
rect 22097 33575 22155 33581
rect 19116 33544 20668 33572
rect 19116 33532 19122 33544
rect 3234 33464 3240 33516
rect 3292 33504 3298 33516
rect 5074 33504 5080 33516
rect 3292 33476 3924 33504
rect 3292 33464 3298 33476
rect 1673 33439 1731 33445
rect 1673 33405 1685 33439
rect 1719 33405 1731 33439
rect 2130 33436 2136 33448
rect 2091 33408 2136 33436
rect 1673 33399 1731 33405
rect 1688 33368 1716 33399
rect 2130 33396 2136 33408
rect 2188 33396 2194 33448
rect 2685 33439 2743 33445
rect 2685 33405 2697 33439
rect 2731 33436 2743 33439
rect 3326 33436 3332 33448
rect 2731 33408 3188 33436
rect 3287 33408 3332 33436
rect 2731 33405 2743 33408
rect 2685 33399 2743 33405
rect 2774 33368 2780 33380
rect 1688 33340 2780 33368
rect 2774 33328 2780 33340
rect 2832 33328 2838 33380
rect 2866 33328 2872 33380
rect 2924 33368 2930 33380
rect 2961 33371 3019 33377
rect 2961 33368 2973 33371
rect 2924 33340 2973 33368
rect 2924 33328 2930 33340
rect 2961 33337 2973 33340
rect 3007 33337 3019 33371
rect 3160 33368 3188 33408
rect 3326 33396 3332 33408
rect 3384 33396 3390 33448
rect 3896 33445 3924 33476
rect 4540 33476 5080 33504
rect 4540 33445 4568 33476
rect 5074 33464 5080 33476
rect 5132 33464 5138 33516
rect 9309 33507 9367 33513
rect 9309 33473 9321 33507
rect 9355 33504 9367 33507
rect 10410 33504 10416 33516
rect 9355 33476 10416 33504
rect 9355 33473 9367 33476
rect 9309 33467 9367 33473
rect 10410 33464 10416 33476
rect 10468 33464 10474 33516
rect 11532 33504 11560 33532
rect 12342 33504 12348 33516
rect 11532 33476 12348 33504
rect 3789 33439 3847 33445
rect 3789 33405 3801 33439
rect 3835 33405 3847 33439
rect 3789 33399 3847 33405
rect 3881 33439 3939 33445
rect 3881 33405 3893 33439
rect 3927 33405 3939 33439
rect 3881 33399 3939 33405
rect 4525 33439 4583 33445
rect 4525 33405 4537 33439
rect 4571 33405 4583 33439
rect 4525 33399 4583 33405
rect 3602 33368 3608 33380
rect 3160 33340 3608 33368
rect 2961 33331 3019 33337
rect 3602 33328 3608 33340
rect 3660 33328 3666 33380
rect 3804 33368 3832 33399
rect 4614 33396 4620 33448
rect 4672 33436 4678 33448
rect 4985 33439 5043 33445
rect 4985 33436 4997 33439
rect 4672 33408 4997 33436
rect 4672 33396 4678 33408
rect 4985 33405 4997 33408
rect 5031 33405 5043 33439
rect 5258 33436 5264 33448
rect 5219 33408 5264 33436
rect 4985 33399 5043 33405
rect 5258 33396 5264 33408
rect 5316 33396 5322 33448
rect 7190 33436 7196 33448
rect 7103 33408 7196 33436
rect 7190 33396 7196 33408
rect 7248 33436 7254 33448
rect 8202 33436 8208 33448
rect 7248 33408 8208 33436
rect 7248 33396 7254 33408
rect 8202 33396 8208 33408
rect 8260 33396 8266 33448
rect 8481 33439 8539 33445
rect 8481 33405 8493 33439
rect 8527 33405 8539 33439
rect 9674 33436 9680 33448
rect 9635 33408 9680 33436
rect 8481 33399 8539 33405
rect 4890 33368 4896 33380
rect 3804 33340 4896 33368
rect 4890 33328 4896 33340
rect 4948 33328 4954 33380
rect 5169 33371 5227 33377
rect 5169 33337 5181 33371
rect 5215 33337 5227 33371
rect 8496 33368 8524 33399
rect 9674 33396 9680 33408
rect 9732 33396 9738 33448
rect 10042 33436 10048 33448
rect 10003 33408 10048 33436
rect 10042 33396 10048 33408
rect 10100 33396 10106 33448
rect 10965 33439 11023 33445
rect 10965 33405 10977 33439
rect 11011 33405 11023 33439
rect 11146 33436 11152 33448
rect 11107 33408 11152 33436
rect 10965 33399 11023 33405
rect 9766 33368 9772 33380
rect 8496 33340 9772 33368
rect 5169 33331 5227 33337
rect 2038 33260 2044 33312
rect 2096 33300 2102 33312
rect 5184 33300 5212 33331
rect 9766 33328 9772 33340
rect 9824 33328 9830 33380
rect 10980 33368 11008 33399
rect 11146 33396 11152 33408
rect 11204 33396 11210 33448
rect 11532 33445 11560 33476
rect 12342 33464 12348 33476
rect 12400 33504 12406 33516
rect 12437 33507 12495 33513
rect 12437 33504 12449 33507
rect 12400 33476 12449 33504
rect 12400 33464 12406 33476
rect 12437 33473 12449 33476
rect 12483 33473 12495 33507
rect 12437 33467 12495 33473
rect 13173 33507 13231 33513
rect 13173 33473 13185 33507
rect 13219 33504 13231 33507
rect 13262 33504 13268 33516
rect 13219 33476 13268 33504
rect 13219 33473 13231 33476
rect 13173 33467 13231 33473
rect 13262 33464 13268 33476
rect 13320 33464 13326 33516
rect 15286 33504 15292 33516
rect 14752 33476 15292 33504
rect 11517 33439 11575 33445
rect 11517 33405 11529 33439
rect 11563 33405 11575 33439
rect 11517 33399 11575 33405
rect 12713 33439 12771 33445
rect 12713 33405 12725 33439
rect 12759 33436 12771 33439
rect 12894 33436 12900 33448
rect 12759 33408 12900 33436
rect 12759 33405 12771 33408
rect 12713 33399 12771 33405
rect 12894 33396 12900 33408
rect 12952 33396 12958 33448
rect 13633 33439 13691 33445
rect 13633 33405 13645 33439
rect 13679 33436 13691 33439
rect 13906 33436 13912 33448
rect 13679 33408 13912 33436
rect 13679 33405 13691 33408
rect 13633 33399 13691 33405
rect 13906 33396 13912 33408
rect 13964 33396 13970 33448
rect 14752 33445 14780 33476
rect 15286 33464 15292 33476
rect 15344 33464 15350 33516
rect 15930 33504 15936 33516
rect 15891 33476 15936 33504
rect 15930 33464 15936 33476
rect 15988 33464 15994 33516
rect 20640 33504 20668 33544
rect 22097 33541 22109 33575
rect 22143 33572 22155 33575
rect 23474 33572 23480 33584
rect 22143 33544 23480 33572
rect 22143 33541 22155 33544
rect 22097 33535 22155 33541
rect 23474 33532 23480 33544
rect 23532 33532 23538 33584
rect 23566 33532 23572 33584
rect 23624 33532 23630 33584
rect 35802 33572 35808 33584
rect 35763 33544 35808 33572
rect 35802 33532 35808 33544
rect 35860 33532 35866 33584
rect 38470 33572 38476 33584
rect 37752 33544 38476 33572
rect 21542 33504 21548 33516
rect 18340 33476 20024 33504
rect 18340 33448 18368 33476
rect 14737 33439 14795 33445
rect 14737 33405 14749 33439
rect 14783 33405 14795 33439
rect 15194 33436 15200 33448
rect 15155 33408 15200 33436
rect 14737 33399 14795 33405
rect 15194 33396 15200 33408
rect 15252 33396 15258 33448
rect 15654 33436 15660 33448
rect 15567 33408 15660 33436
rect 15654 33396 15660 33408
rect 15712 33436 15718 33448
rect 16390 33436 16396 33448
rect 15712 33408 16396 33436
rect 15712 33396 15718 33408
rect 16390 33396 16396 33408
rect 16448 33396 16454 33448
rect 18233 33439 18291 33445
rect 18233 33405 18245 33439
rect 18279 33436 18291 33439
rect 18322 33436 18328 33448
rect 18279 33408 18328 33436
rect 18279 33405 18291 33408
rect 18233 33399 18291 33405
rect 18322 33396 18328 33408
rect 18380 33396 18386 33448
rect 18785 33439 18843 33445
rect 18785 33405 18797 33439
rect 18831 33405 18843 33439
rect 18966 33436 18972 33448
rect 18927 33408 18972 33436
rect 18785 33399 18843 33405
rect 11054 33368 11060 33380
rect 10967 33340 11060 33368
rect 11054 33328 11060 33340
rect 11112 33368 11118 33380
rect 11606 33368 11612 33380
rect 11112 33340 11612 33368
rect 11112 33328 11118 33340
rect 11606 33328 11612 33340
rect 11664 33368 11670 33380
rect 12805 33371 12863 33377
rect 12805 33368 12817 33371
rect 11664 33340 12817 33368
rect 11664 33328 11670 33340
rect 12805 33337 12817 33340
rect 12851 33368 12863 33371
rect 13814 33368 13820 33380
rect 12851 33340 13820 33368
rect 12851 33337 12863 33340
rect 12805 33331 12863 33337
rect 13814 33328 13820 33340
rect 13872 33328 13878 33380
rect 18800 33368 18828 33399
rect 18966 33396 18972 33408
rect 19024 33396 19030 33448
rect 19797 33439 19855 33445
rect 19797 33405 19809 33439
rect 19843 33436 19855 33439
rect 19886 33436 19892 33448
rect 19843 33408 19892 33436
rect 19843 33405 19855 33408
rect 19797 33399 19855 33405
rect 19886 33396 19892 33408
rect 19944 33396 19950 33448
rect 19996 33445 20024 33476
rect 20640 33476 21548 33504
rect 20640 33445 20668 33476
rect 21542 33464 21548 33476
rect 21600 33464 21606 33516
rect 23584 33504 23612 33532
rect 24394 33504 24400 33516
rect 23584 33476 24400 33504
rect 24394 33464 24400 33476
rect 24452 33504 24458 33516
rect 25133 33507 25191 33513
rect 25133 33504 25145 33507
rect 24452 33476 25145 33504
rect 24452 33464 24458 33476
rect 25133 33473 25145 33476
rect 25179 33473 25191 33507
rect 25133 33467 25191 33473
rect 25777 33507 25835 33513
rect 25777 33473 25789 33507
rect 25823 33504 25835 33507
rect 26234 33504 26240 33516
rect 25823 33476 26240 33504
rect 25823 33473 25835 33476
rect 25777 33467 25835 33473
rect 26234 33464 26240 33476
rect 26292 33504 26298 33516
rect 26292 33476 28120 33504
rect 26292 33464 26298 33476
rect 19981 33439 20039 33445
rect 19981 33405 19993 33439
rect 20027 33405 20039 33439
rect 19981 33399 20039 33405
rect 20625 33439 20683 33445
rect 20625 33405 20637 33439
rect 20671 33405 20683 33439
rect 20625 33399 20683 33405
rect 20993 33439 21051 33445
rect 20993 33405 21005 33439
rect 21039 33436 21051 33439
rect 21358 33436 21364 33448
rect 21039 33408 21364 33436
rect 21039 33405 21051 33408
rect 20993 33399 21051 33405
rect 21358 33396 21364 33408
rect 21416 33396 21422 33448
rect 21729 33439 21787 33445
rect 21729 33405 21741 33439
rect 21775 33405 21787 33439
rect 21729 33399 21787 33405
rect 19058 33368 19064 33380
rect 18800 33340 19064 33368
rect 19058 33328 19064 33340
rect 19116 33328 19122 33380
rect 21744 33368 21772 33399
rect 21818 33396 21824 33448
rect 21876 33436 21882 33448
rect 22370 33436 22376 33448
rect 21876 33408 21921 33436
rect 22331 33408 22376 33436
rect 21876 33396 21882 33408
rect 22370 33396 22376 33408
rect 22428 33396 22434 33448
rect 22833 33439 22891 33445
rect 22833 33405 22845 33439
rect 22879 33436 22891 33439
rect 23566 33436 23572 33448
rect 22879 33408 23572 33436
rect 22879 33405 22891 33408
rect 22833 33399 22891 33405
rect 23566 33396 23572 33408
rect 23624 33396 23630 33448
rect 23661 33439 23719 33445
rect 23661 33405 23673 33439
rect 23707 33436 23719 33439
rect 23750 33436 23756 33448
rect 23707 33408 23756 33436
rect 23707 33405 23719 33408
rect 23661 33399 23719 33405
rect 23750 33396 23756 33408
rect 23808 33396 23814 33448
rect 23934 33436 23940 33448
rect 23895 33408 23940 33436
rect 23934 33396 23940 33408
rect 23992 33396 23998 33448
rect 25038 33396 25044 33448
rect 25096 33436 25102 33448
rect 25593 33439 25651 33445
rect 25593 33436 25605 33439
rect 25096 33408 25605 33436
rect 25096 33396 25102 33408
rect 25593 33405 25605 33408
rect 25639 33405 25651 33439
rect 25593 33399 25651 33405
rect 25869 33439 25927 33445
rect 25869 33405 25881 33439
rect 25915 33405 25927 33439
rect 25869 33399 25927 33405
rect 19628 33340 21772 33368
rect 25608 33368 25636 33399
rect 25884 33368 25912 33399
rect 27154 33396 27160 33448
rect 27212 33436 27218 33448
rect 27249 33439 27307 33445
rect 27249 33436 27261 33439
rect 27212 33408 27261 33436
rect 27212 33396 27218 33408
rect 27249 33405 27261 33408
rect 27295 33405 27307 33439
rect 27249 33399 27307 33405
rect 27338 33396 27344 33448
rect 27396 33436 27402 33448
rect 27433 33439 27491 33445
rect 27433 33436 27445 33439
rect 27396 33408 27445 33436
rect 27396 33396 27402 33408
rect 27433 33405 27445 33408
rect 27479 33405 27491 33439
rect 27798 33436 27804 33448
rect 27759 33408 27804 33436
rect 27433 33399 27491 33405
rect 27798 33396 27804 33408
rect 27856 33396 27862 33448
rect 27890 33396 27896 33448
rect 27948 33436 27954 33448
rect 27948 33408 27993 33436
rect 27948 33396 27954 33408
rect 26786 33368 26792 33380
rect 25608 33340 25912 33368
rect 26747 33340 26792 33368
rect 8570 33300 8576 33312
rect 2096 33272 5212 33300
rect 8531 33272 8576 33300
rect 2096 33260 2102 33272
rect 8570 33260 8576 33272
rect 8628 33260 8634 33312
rect 10410 33260 10416 33312
rect 10468 33300 10474 33312
rect 11698 33300 11704 33312
rect 10468 33272 11704 33300
rect 10468 33260 10474 33272
rect 11698 33260 11704 33272
rect 11756 33300 11762 33312
rect 12621 33303 12679 33309
rect 12621 33300 12633 33303
rect 11756 33272 12633 33300
rect 11756 33260 11762 33272
rect 12621 33269 12633 33272
rect 12667 33300 12679 33303
rect 17678 33300 17684 33312
rect 12667 33272 17684 33300
rect 12667 33269 12679 33272
rect 12621 33263 12679 33269
rect 17678 33260 17684 33272
rect 17736 33260 17742 33312
rect 18138 33300 18144 33312
rect 18099 33272 18144 33300
rect 18138 33260 18144 33272
rect 18196 33260 18202 33312
rect 19242 33260 19248 33312
rect 19300 33300 19306 33312
rect 19628 33309 19656 33340
rect 26786 33328 26792 33340
rect 26844 33328 26850 33380
rect 28092 33368 28120 33476
rect 28166 33464 28172 33516
rect 28224 33504 28230 33516
rect 30285 33507 30343 33513
rect 30285 33504 30297 33507
rect 28224 33476 30297 33504
rect 28224 33464 28230 33476
rect 30285 33473 30297 33476
rect 30331 33473 30343 33507
rect 30285 33467 30343 33473
rect 31757 33507 31815 33513
rect 31757 33473 31769 33507
rect 31803 33504 31815 33507
rect 32398 33504 32404 33516
rect 31803 33476 32404 33504
rect 31803 33473 31815 33476
rect 31757 33467 31815 33473
rect 32398 33464 32404 33476
rect 32456 33464 32462 33516
rect 32677 33507 32735 33513
rect 32677 33473 32689 33507
rect 32723 33504 32735 33507
rect 32858 33504 32864 33516
rect 32723 33476 32864 33504
rect 32723 33473 32735 33476
rect 32677 33467 32735 33473
rect 32858 33464 32864 33476
rect 32916 33464 32922 33516
rect 32953 33507 33011 33513
rect 32953 33473 32965 33507
rect 32999 33504 33011 33507
rect 34330 33504 34336 33516
rect 32999 33476 34336 33504
rect 32999 33473 33011 33476
rect 32953 33467 33011 33473
rect 34330 33464 34336 33476
rect 34388 33464 34394 33516
rect 28442 33436 28448 33448
rect 28403 33408 28448 33436
rect 28442 33396 28448 33408
rect 28500 33396 28506 33448
rect 29273 33439 29331 33445
rect 29273 33405 29285 33439
rect 29319 33405 29331 33439
rect 29273 33399 29331 33405
rect 29365 33439 29423 33445
rect 29365 33405 29377 33439
rect 29411 33405 29423 33439
rect 30374 33436 30380 33448
rect 30335 33408 30380 33436
rect 29365 33399 29423 33405
rect 29288 33368 29316 33399
rect 28092 33340 29316 33368
rect 19613 33303 19671 33309
rect 19613 33300 19625 33303
rect 19300 33272 19625 33300
rect 19300 33260 19306 33272
rect 19613 33269 19625 33272
rect 19659 33269 19671 33303
rect 20070 33300 20076 33312
rect 20031 33272 20076 33300
rect 19613 33263 19671 33269
rect 20070 33260 20076 33272
rect 20128 33260 20134 33312
rect 29380 33300 29408 33399
rect 30374 33396 30380 33408
rect 30432 33396 30438 33448
rect 31665 33439 31723 33445
rect 31665 33405 31677 33439
rect 31711 33405 31723 33439
rect 31938 33436 31944 33448
rect 31899 33408 31944 33436
rect 31665 33399 31723 33405
rect 31680 33368 31708 33399
rect 31938 33396 31944 33408
rect 31996 33396 32002 33448
rect 33594 33396 33600 33448
rect 33652 33436 33658 33448
rect 34885 33439 34943 33445
rect 34885 33436 34897 33439
rect 33652 33408 34897 33436
rect 33652 33396 33658 33408
rect 34885 33405 34897 33408
rect 34931 33405 34943 33439
rect 34885 33399 34943 33405
rect 35253 33439 35311 33445
rect 35253 33405 35265 33439
rect 35299 33405 35311 33439
rect 35802 33436 35808 33448
rect 35763 33408 35808 33436
rect 35253 33399 35311 33405
rect 32306 33368 32312 33380
rect 31680 33340 32312 33368
rect 32306 33328 32312 33340
rect 32364 33328 32370 33380
rect 35268 33368 35296 33399
rect 35802 33396 35808 33408
rect 35860 33396 35866 33448
rect 36449 33439 36507 33445
rect 36449 33405 36461 33439
rect 36495 33405 36507 33439
rect 36449 33399 36507 33405
rect 36464 33368 36492 33399
rect 36630 33396 36636 33448
rect 36688 33436 36694 33448
rect 37752 33445 37780 33544
rect 38470 33532 38476 33544
rect 38528 33572 38534 33584
rect 38933 33575 38991 33581
rect 38933 33572 38945 33575
rect 38528 33544 38945 33572
rect 38528 33532 38534 33544
rect 38933 33541 38945 33544
rect 38979 33541 38991 33575
rect 38933 33535 38991 33541
rect 38286 33504 38292 33516
rect 38247 33476 38292 33504
rect 38286 33464 38292 33476
rect 38344 33464 38350 33516
rect 37185 33439 37243 33445
rect 37185 33436 37197 33439
rect 36688 33408 37197 33436
rect 36688 33396 36694 33408
rect 37185 33405 37197 33408
rect 37231 33405 37243 33439
rect 37185 33399 37243 33405
rect 37737 33439 37795 33445
rect 37737 33405 37749 33439
rect 37783 33405 37795 33439
rect 38102 33436 38108 33448
rect 38063 33408 38108 33436
rect 37737 33399 37795 33405
rect 38102 33396 38108 33408
rect 38160 33396 38166 33448
rect 38749 33439 38807 33445
rect 38749 33405 38761 33439
rect 38795 33405 38807 33439
rect 38749 33399 38807 33405
rect 35268 33340 36492 33368
rect 29914 33300 29920 33312
rect 29380 33272 29920 33300
rect 29914 33260 29920 33272
rect 29972 33260 29978 33312
rect 34514 33260 34520 33312
rect 34572 33300 34578 33312
rect 35268 33300 35296 33340
rect 36722 33328 36728 33380
rect 36780 33368 36786 33380
rect 38764 33368 38792 33399
rect 36780 33340 38792 33368
rect 36780 33328 36786 33340
rect 34572 33272 35296 33300
rect 34572 33260 34578 33272
rect 36354 33260 36360 33312
rect 36412 33300 36418 33312
rect 36633 33303 36691 33309
rect 36633 33300 36645 33303
rect 36412 33272 36645 33300
rect 36412 33260 36418 33272
rect 36633 33269 36645 33272
rect 36679 33300 36691 33303
rect 37642 33300 37648 33312
rect 36679 33272 37648 33300
rect 36679 33269 36691 33272
rect 36633 33263 36691 33269
rect 37642 33260 37648 33272
rect 37700 33260 37706 33312
rect 1104 33210 39836 33232
rect 1104 33158 19606 33210
rect 19658 33158 19670 33210
rect 19722 33158 19734 33210
rect 19786 33158 19798 33210
rect 19850 33158 39836 33210
rect 1104 33136 39836 33158
rect 4798 33056 4804 33108
rect 4856 33096 4862 33108
rect 4893 33099 4951 33105
rect 4893 33096 4905 33099
rect 4856 33068 4905 33096
rect 4856 33056 4862 33068
rect 4893 33065 4905 33068
rect 4939 33096 4951 33099
rect 5166 33096 5172 33108
rect 4939 33068 5172 33096
rect 4939 33065 4951 33068
rect 4893 33059 4951 33065
rect 5166 33056 5172 33068
rect 5224 33056 5230 33108
rect 13906 33056 13912 33108
rect 13964 33096 13970 33108
rect 16485 33099 16543 33105
rect 13964 33068 16068 33096
rect 13964 33056 13970 33068
rect 1854 32988 1860 33040
rect 1912 33028 1918 33040
rect 2317 33031 2375 33037
rect 2317 33028 2329 33031
rect 1912 33000 2329 33028
rect 1912 32988 1918 33000
rect 2317 32997 2329 33000
rect 2363 32997 2375 33031
rect 5074 33028 5080 33040
rect 5035 33000 5080 33028
rect 2317 32991 2375 32997
rect 5074 32988 5080 33000
rect 5132 32988 5138 33040
rect 5626 32988 5632 33040
rect 5684 33028 5690 33040
rect 5684 33000 6408 33028
rect 5684 32988 5690 33000
rect 2866 32960 2872 32972
rect 2827 32932 2872 32960
rect 2866 32920 2872 32932
rect 2924 32920 2930 32972
rect 3142 32960 3148 32972
rect 3103 32932 3148 32960
rect 3142 32920 3148 32932
rect 3200 32920 3206 32972
rect 3234 32920 3240 32972
rect 3292 32960 3298 32972
rect 3329 32963 3387 32969
rect 3329 32960 3341 32963
rect 3292 32932 3341 32960
rect 3292 32920 3298 32932
rect 3329 32929 3341 32932
rect 3375 32960 3387 32963
rect 4985 32963 5043 32969
rect 4985 32960 4997 32963
rect 3375 32932 4997 32960
rect 3375 32929 3387 32932
rect 3329 32923 3387 32929
rect 4985 32929 4997 32932
rect 5031 32960 5043 32963
rect 5258 32960 5264 32972
rect 5031 32932 5264 32960
rect 5031 32929 5043 32932
rect 4985 32923 5043 32929
rect 5258 32920 5264 32932
rect 5316 32920 5322 32972
rect 6270 32960 6276 32972
rect 6231 32932 6276 32960
rect 6270 32920 6276 32932
rect 6328 32920 6334 32972
rect 6380 32969 6408 33000
rect 6454 32988 6460 33040
rect 6512 33028 6518 33040
rect 10042 33028 10048 33040
rect 6512 33000 7236 33028
rect 10003 33000 10048 33028
rect 6512 32988 6518 33000
rect 7208 32969 7236 33000
rect 10042 32988 10048 33000
rect 10100 32988 10106 33040
rect 12434 32988 12440 33040
rect 12492 33028 12498 33040
rect 12492 33000 12537 33028
rect 12492 32988 12498 33000
rect 12618 32988 12624 33040
rect 12676 33028 12682 33040
rect 16040 33037 16068 33068
rect 16485 33065 16497 33099
rect 16531 33096 16543 33099
rect 16574 33096 16580 33108
rect 16531 33068 16580 33096
rect 16531 33065 16543 33068
rect 16485 33059 16543 33065
rect 16574 33056 16580 33068
rect 16632 33096 16638 33108
rect 17310 33096 17316 33108
rect 16632 33068 17316 33096
rect 16632 33056 16638 33068
rect 17310 33056 17316 33068
rect 17368 33056 17374 33108
rect 20073 33099 20131 33105
rect 20073 33065 20085 33099
rect 20119 33096 20131 33099
rect 20162 33096 20168 33108
rect 20119 33068 20168 33096
rect 20119 33065 20131 33068
rect 20073 33059 20131 33065
rect 20162 33056 20168 33068
rect 20220 33056 20226 33108
rect 21453 33099 21511 33105
rect 21453 33065 21465 33099
rect 21499 33096 21511 33099
rect 24486 33096 24492 33108
rect 21499 33068 24492 33096
rect 21499 33065 21511 33068
rect 21453 33059 21511 33065
rect 24486 33056 24492 33068
rect 24544 33056 24550 33108
rect 24964 33068 30604 33096
rect 15657 33031 15715 33037
rect 15657 33028 15669 33031
rect 12676 33000 15669 33028
rect 12676 32988 12682 33000
rect 15657 32997 15669 33000
rect 15703 33028 15715 33031
rect 16025 33031 16083 33037
rect 15703 33000 15792 33028
rect 15703 32997 15715 33000
rect 15657 32991 15715 32997
rect 6365 32963 6423 32969
rect 6365 32929 6377 32963
rect 6411 32929 6423 32963
rect 6365 32923 6423 32929
rect 6825 32963 6883 32969
rect 6825 32929 6837 32963
rect 6871 32929 6883 32963
rect 6825 32923 6883 32929
rect 7193 32963 7251 32969
rect 7193 32929 7205 32963
rect 7239 32929 7251 32963
rect 7193 32923 7251 32929
rect 7837 32963 7895 32969
rect 7837 32929 7849 32963
rect 7883 32960 7895 32963
rect 8018 32960 8024 32972
rect 7883 32932 8024 32960
rect 7883 32929 7895 32932
rect 7837 32923 7895 32929
rect 4709 32895 4767 32901
rect 4709 32861 4721 32895
rect 4755 32892 4767 32895
rect 4890 32892 4896 32904
rect 4755 32864 4896 32892
rect 4755 32861 4767 32864
rect 4709 32855 4767 32861
rect 4890 32852 4896 32864
rect 4948 32852 4954 32904
rect 5445 32895 5503 32901
rect 5445 32861 5457 32895
rect 5491 32892 5503 32895
rect 6840 32892 6868 32923
rect 8018 32920 8024 32932
rect 8076 32920 8082 32972
rect 8573 32963 8631 32969
rect 8573 32929 8585 32963
rect 8619 32960 8631 32963
rect 8662 32960 8668 32972
rect 8619 32932 8668 32960
rect 8619 32929 8631 32932
rect 8573 32923 8631 32929
rect 8662 32920 8668 32932
rect 8720 32960 8726 32972
rect 9677 32963 9735 32969
rect 9677 32960 9689 32963
rect 8720 32932 9689 32960
rect 8720 32920 8726 32932
rect 9677 32929 9689 32932
rect 9723 32929 9735 32963
rect 10410 32960 10416 32972
rect 10371 32932 10416 32960
rect 9677 32923 9735 32929
rect 10410 32920 10416 32932
rect 10468 32920 10474 32972
rect 10873 32963 10931 32969
rect 10873 32929 10885 32963
rect 10919 32929 10931 32963
rect 11054 32960 11060 32972
rect 11015 32932 11060 32960
rect 10873 32923 10931 32929
rect 5491 32864 6868 32892
rect 10888 32892 10916 32923
rect 11054 32920 11060 32932
rect 11112 32920 11118 32972
rect 11606 32960 11612 32972
rect 11567 32932 11612 32960
rect 11606 32920 11612 32932
rect 11664 32920 11670 32972
rect 12250 32960 12256 32972
rect 12211 32932 12256 32960
rect 12250 32920 12256 32932
rect 12308 32920 12314 32972
rect 12345 32963 12403 32969
rect 12345 32929 12357 32963
rect 12391 32929 12403 32963
rect 12345 32923 12403 32929
rect 12805 32963 12863 32969
rect 12805 32929 12817 32963
rect 12851 32960 12863 32963
rect 14093 32963 14151 32969
rect 14093 32960 14105 32963
rect 12851 32932 14105 32960
rect 12851 32929 12863 32932
rect 12805 32923 12863 32929
rect 14093 32929 14105 32932
rect 14139 32929 14151 32963
rect 15470 32960 15476 32972
rect 15431 32932 15476 32960
rect 14093 32923 14151 32929
rect 11790 32892 11796 32904
rect 10888 32864 11796 32892
rect 5491 32861 5503 32864
rect 5445 32855 5503 32861
rect 11790 32852 11796 32864
rect 11848 32892 11854 32904
rect 12069 32895 12127 32901
rect 12069 32892 12081 32895
rect 11848 32864 12081 32892
rect 11848 32852 11854 32864
rect 12069 32861 12081 32864
rect 12115 32861 12127 32895
rect 12360 32892 12388 32923
rect 15470 32920 15476 32932
rect 15528 32920 15534 32972
rect 15562 32920 15568 32972
rect 15620 32960 15626 32972
rect 15764 32960 15792 33000
rect 16025 32997 16037 33031
rect 16071 32997 16083 33031
rect 17218 33028 17224 33040
rect 16025 32991 16083 32997
rect 16132 33000 17224 33028
rect 16132 32960 16160 33000
rect 17218 32988 17224 33000
rect 17276 32988 17282 33040
rect 22186 33028 22192 33040
rect 21560 33000 22192 33028
rect 15620 32932 15665 32960
rect 15764 32932 16160 32960
rect 16669 32963 16727 32969
rect 15620 32920 15626 32932
rect 16669 32929 16681 32963
rect 16715 32929 16727 32963
rect 16942 32960 16948 32972
rect 16903 32932 16948 32960
rect 16669 32923 16727 32929
rect 12069 32855 12127 32861
rect 12176 32864 12388 32892
rect 13265 32895 13323 32901
rect 5905 32827 5963 32833
rect 5905 32793 5917 32827
rect 5951 32824 5963 32827
rect 7190 32824 7196 32836
rect 5951 32796 7196 32824
rect 5951 32793 5963 32796
rect 5905 32787 5963 32793
rect 7190 32784 7196 32796
rect 7248 32784 7254 32836
rect 11974 32784 11980 32836
rect 12032 32824 12038 32836
rect 12176 32824 12204 32864
rect 13265 32861 13277 32895
rect 13311 32861 13323 32895
rect 13814 32892 13820 32904
rect 13775 32864 13820 32892
rect 13265 32855 13323 32861
rect 12032 32796 12204 32824
rect 13280 32824 13308 32855
rect 13814 32852 13820 32864
rect 13872 32852 13878 32904
rect 14274 32892 14280 32904
rect 14235 32864 14280 32892
rect 14274 32852 14280 32864
rect 14332 32852 14338 32904
rect 15286 32892 15292 32904
rect 15247 32864 15292 32892
rect 15286 32852 15292 32864
rect 15344 32852 15350 32904
rect 16684 32892 16712 32923
rect 16942 32920 16948 32932
rect 17000 32920 17006 32972
rect 17494 32960 17500 32972
rect 17455 32932 17500 32960
rect 17494 32920 17500 32932
rect 17552 32920 17558 32972
rect 17773 32963 17831 32969
rect 17773 32929 17785 32963
rect 17819 32960 17831 32963
rect 18138 32960 18144 32972
rect 17819 32932 18144 32960
rect 17819 32929 17831 32932
rect 17773 32923 17831 32929
rect 18138 32920 18144 32932
rect 18196 32920 18202 32972
rect 18322 32960 18328 32972
rect 18283 32932 18328 32960
rect 18322 32920 18328 32932
rect 18380 32920 18386 32972
rect 19058 32960 19064 32972
rect 19019 32932 19064 32960
rect 19058 32920 19064 32932
rect 19116 32920 19122 32972
rect 19337 32963 19395 32969
rect 19337 32929 19349 32963
rect 19383 32960 19395 32963
rect 19889 32963 19947 32969
rect 19889 32960 19901 32963
rect 19383 32932 19901 32960
rect 19383 32929 19395 32932
rect 19337 32923 19395 32929
rect 19889 32929 19901 32932
rect 19935 32960 19947 32963
rect 19978 32960 19984 32972
rect 19935 32932 19984 32960
rect 19935 32929 19947 32932
rect 19889 32923 19947 32929
rect 19978 32920 19984 32932
rect 20036 32920 20042 32972
rect 21560 32969 21588 33000
rect 22186 32988 22192 33000
rect 22244 32988 22250 33040
rect 21545 32963 21603 32969
rect 21545 32929 21557 32963
rect 21591 32929 21603 32963
rect 21545 32923 21603 32929
rect 22094 32920 22100 32972
rect 22152 32960 22158 32972
rect 22152 32932 22197 32960
rect 22152 32920 22158 32932
rect 22830 32920 22836 32972
rect 22888 32960 22894 32972
rect 22925 32963 22983 32969
rect 22925 32960 22937 32963
rect 22888 32932 22937 32960
rect 22888 32920 22894 32932
rect 22925 32929 22937 32932
rect 22971 32929 22983 32963
rect 23474 32960 23480 32972
rect 23435 32932 23480 32960
rect 22925 32923 22983 32929
rect 23474 32920 23480 32932
rect 23532 32920 23538 32972
rect 24964 32969 24992 33068
rect 30576 33028 30604 33068
rect 30834 33056 30840 33108
rect 30892 33096 30898 33108
rect 31110 33096 31116 33108
rect 30892 33068 31116 33096
rect 30892 33056 30898 33068
rect 31110 33056 31116 33068
rect 31168 33096 31174 33108
rect 31757 33099 31815 33105
rect 31757 33096 31769 33099
rect 31168 33068 31769 33096
rect 31168 33056 31174 33068
rect 31757 33065 31769 33068
rect 31803 33065 31815 33099
rect 33226 33096 33232 33108
rect 31757 33059 31815 33065
rect 32416 33068 33232 33096
rect 32416 33028 32444 33068
rect 33226 33056 33232 33068
rect 33284 33056 33290 33108
rect 33502 33028 33508 33040
rect 30576 33000 32444 33028
rect 32508 33000 33508 33028
rect 24949 32963 25007 32969
rect 24949 32929 24961 32963
rect 24995 32929 25007 32963
rect 24949 32923 25007 32929
rect 25409 32963 25467 32969
rect 25409 32929 25421 32963
rect 25455 32960 25467 32963
rect 25498 32960 25504 32972
rect 25455 32932 25504 32960
rect 25455 32929 25467 32932
rect 25409 32923 25467 32929
rect 25498 32920 25504 32932
rect 25556 32920 25562 32972
rect 26513 32963 26571 32969
rect 26513 32929 26525 32963
rect 26559 32960 26571 32963
rect 27154 32960 27160 32972
rect 26559 32932 27160 32960
rect 26559 32929 26571 32932
rect 26513 32923 26571 32929
rect 27154 32920 27160 32932
rect 27212 32920 27218 32972
rect 29089 32963 29147 32969
rect 29089 32929 29101 32963
rect 29135 32960 29147 32963
rect 29917 32963 29975 32969
rect 29135 32932 29868 32960
rect 29135 32929 29147 32932
rect 29089 32923 29147 32929
rect 19242 32892 19248 32904
rect 16684 32864 19248 32892
rect 19242 32852 19248 32864
rect 19300 32852 19306 32904
rect 20254 32852 20260 32904
rect 20312 32892 20318 32904
rect 22189 32895 22247 32901
rect 22189 32892 22201 32895
rect 20312 32864 22201 32892
rect 20312 32852 20318 32864
rect 22189 32861 22201 32864
rect 22235 32861 22247 32895
rect 22189 32855 22247 32861
rect 24854 32852 24860 32904
rect 24912 32892 24918 32904
rect 25041 32895 25099 32901
rect 25041 32892 25053 32895
rect 24912 32864 25053 32892
rect 24912 32852 24918 32864
rect 25041 32861 25053 32864
rect 25087 32861 25099 32895
rect 25041 32855 25099 32861
rect 26326 32852 26332 32904
rect 26384 32892 26390 32904
rect 27433 32895 27491 32901
rect 27433 32892 27445 32895
rect 26384 32864 27445 32892
rect 26384 32852 26390 32864
rect 27433 32861 27445 32864
rect 27479 32861 27491 32895
rect 27706 32892 27712 32904
rect 27667 32864 27712 32892
rect 27433 32855 27491 32861
rect 27706 32852 27712 32864
rect 27764 32852 27770 32904
rect 29546 32852 29552 32904
rect 29604 32892 29610 32904
rect 29641 32895 29699 32901
rect 29641 32892 29653 32895
rect 29604 32864 29653 32892
rect 29604 32852 29610 32864
rect 29641 32861 29653 32864
rect 29687 32861 29699 32895
rect 29840 32892 29868 32932
rect 29917 32929 29929 32963
rect 29963 32960 29975 32963
rect 30558 32960 30564 32972
rect 29963 32932 30564 32960
rect 29963 32929 29975 32932
rect 29917 32923 29975 32929
rect 30558 32920 30564 32932
rect 30616 32920 30622 32972
rect 32508 32969 32536 33000
rect 33502 32988 33508 33000
rect 33560 32988 33566 33040
rect 35342 33028 35348 33040
rect 35303 33000 35348 33028
rect 35342 32988 35348 33000
rect 35400 32988 35406 33040
rect 37918 32988 37924 33040
rect 37976 33028 37982 33040
rect 38289 33031 38347 33037
rect 38289 33028 38301 33031
rect 37976 33000 38301 33028
rect 37976 32988 37982 33000
rect 38289 32997 38301 33000
rect 38335 32997 38347 33031
rect 38289 32991 38347 32997
rect 31941 32963 31999 32969
rect 31941 32929 31953 32963
rect 31987 32929 31999 32963
rect 31941 32923 31999 32929
rect 32493 32963 32551 32969
rect 32493 32929 32505 32963
rect 32539 32929 32551 32963
rect 32493 32923 32551 32929
rect 32953 32963 33011 32969
rect 32953 32929 32965 32963
rect 32999 32960 33011 32963
rect 33318 32960 33324 32972
rect 32999 32932 33324 32960
rect 32999 32929 33011 32932
rect 32953 32923 33011 32929
rect 31662 32892 31668 32904
rect 29840 32864 31668 32892
rect 29641 32855 29699 32861
rect 31662 32852 31668 32864
rect 31720 32852 31726 32904
rect 31956 32892 31984 32923
rect 33318 32920 33324 32932
rect 33376 32920 33382 32972
rect 34054 32920 34060 32972
rect 34112 32960 34118 32972
rect 34241 32963 34299 32969
rect 34241 32960 34253 32963
rect 34112 32932 34253 32960
rect 34112 32920 34118 32932
rect 34241 32929 34253 32932
rect 34287 32929 34299 32963
rect 34241 32923 34299 32929
rect 34514 32920 34520 32972
rect 34572 32960 34578 32972
rect 34609 32963 34667 32969
rect 34609 32960 34621 32963
rect 34572 32932 34621 32960
rect 34572 32920 34578 32932
rect 34609 32929 34621 32932
rect 34655 32929 34667 32963
rect 34609 32923 34667 32929
rect 35161 32963 35219 32969
rect 35161 32929 35173 32963
rect 35207 32960 35219 32963
rect 35802 32960 35808 32972
rect 35207 32932 35808 32960
rect 35207 32929 35219 32932
rect 35161 32923 35219 32929
rect 35802 32920 35808 32932
rect 35860 32920 35866 32972
rect 36446 32920 36452 32972
rect 36504 32960 36510 32972
rect 36633 32963 36691 32969
rect 36633 32960 36645 32963
rect 36504 32932 36645 32960
rect 36504 32920 36510 32932
rect 36633 32929 36645 32932
rect 36679 32960 36691 32963
rect 36722 32960 36728 32972
rect 36679 32932 36728 32960
rect 36679 32929 36691 32932
rect 36633 32923 36691 32929
rect 36722 32920 36728 32932
rect 36780 32920 36786 32972
rect 36906 32960 36912 32972
rect 36867 32932 36912 32960
rect 36906 32920 36912 32932
rect 36964 32920 36970 32972
rect 38473 32963 38531 32969
rect 38473 32929 38485 32963
rect 38519 32960 38531 32963
rect 38562 32960 38568 32972
rect 38519 32932 38568 32960
rect 38519 32929 38531 32932
rect 38473 32923 38531 32929
rect 38562 32920 38568 32932
rect 38620 32920 38626 32972
rect 36262 32892 36268 32904
rect 31956 32864 32812 32892
rect 36223 32864 36268 32892
rect 32784 32836 32812 32864
rect 36262 32852 36268 32864
rect 36320 32852 36326 32904
rect 38746 32892 38752 32904
rect 38707 32864 38752 32892
rect 38746 32852 38752 32864
rect 38804 32852 38810 32904
rect 15930 32824 15936 32836
rect 13280 32796 15936 32824
rect 12032 32784 12038 32796
rect 15930 32784 15936 32796
rect 15988 32784 15994 32836
rect 16850 32824 16856 32836
rect 16811 32796 16856 32824
rect 16850 32784 16856 32796
rect 16908 32784 16914 32836
rect 18601 32827 18659 32833
rect 18601 32793 18613 32827
rect 18647 32824 18659 32827
rect 19058 32824 19064 32836
rect 18647 32796 19064 32824
rect 18647 32793 18659 32796
rect 18601 32787 18659 32793
rect 19058 32784 19064 32796
rect 19116 32784 19122 32836
rect 19150 32784 19156 32836
rect 19208 32824 19214 32836
rect 21818 32824 21824 32836
rect 19208 32796 21824 32824
rect 19208 32784 19214 32796
rect 21818 32784 21824 32796
rect 21876 32784 21882 32836
rect 32306 32824 32312 32836
rect 32267 32796 32312 32824
rect 32306 32784 32312 32796
rect 32364 32784 32370 32836
rect 32766 32784 32772 32836
rect 32824 32784 32830 32836
rect 36078 32784 36084 32836
rect 36136 32824 36142 32836
rect 36909 32827 36967 32833
rect 36909 32824 36921 32827
rect 36136 32796 36921 32824
rect 36136 32784 36142 32796
rect 36909 32793 36921 32796
rect 36955 32793 36967 32827
rect 36909 32787 36967 32793
rect 3602 32716 3608 32768
rect 3660 32756 3666 32768
rect 8757 32759 8815 32765
rect 8757 32756 8769 32759
rect 3660 32728 8769 32756
rect 3660 32716 3666 32728
rect 8757 32725 8769 32728
rect 8803 32756 8815 32759
rect 10410 32756 10416 32768
rect 8803 32728 10416 32756
rect 8803 32725 8815 32728
rect 8757 32719 8815 32725
rect 10410 32716 10416 32728
rect 10468 32716 10474 32768
rect 17862 32716 17868 32768
rect 17920 32756 17926 32768
rect 21726 32756 21732 32768
rect 17920 32728 21732 32756
rect 17920 32716 17926 32728
rect 21726 32716 21732 32728
rect 21784 32716 21790 32768
rect 22462 32716 22468 32768
rect 22520 32756 22526 32768
rect 23017 32759 23075 32765
rect 23017 32756 23029 32759
rect 22520 32728 23029 32756
rect 22520 32716 22526 32728
rect 23017 32725 23029 32728
rect 23063 32725 23075 32759
rect 23017 32719 23075 32725
rect 23474 32716 23480 32768
rect 23532 32756 23538 32768
rect 24578 32756 24584 32768
rect 23532 32728 24584 32756
rect 23532 32716 23538 32728
rect 24578 32716 24584 32728
rect 24636 32756 24642 32768
rect 26697 32759 26755 32765
rect 26697 32756 26709 32759
rect 24636 32728 26709 32756
rect 24636 32716 24642 32728
rect 26697 32725 26709 32728
rect 26743 32725 26755 32759
rect 26697 32719 26755 32725
rect 29086 32716 29092 32768
rect 29144 32756 29150 32768
rect 31021 32759 31079 32765
rect 31021 32756 31033 32759
rect 29144 32728 31033 32756
rect 29144 32716 29150 32728
rect 31021 32725 31033 32728
rect 31067 32725 31079 32759
rect 31021 32719 31079 32725
rect 1104 32666 39836 32688
rect 1104 32614 4246 32666
rect 4298 32614 4310 32666
rect 4362 32614 4374 32666
rect 4426 32614 4438 32666
rect 4490 32614 34966 32666
rect 35018 32614 35030 32666
rect 35082 32614 35094 32666
rect 35146 32614 35158 32666
rect 35210 32614 39836 32666
rect 1104 32592 39836 32614
rect 6178 32552 6184 32564
rect 6139 32524 6184 32552
rect 6178 32512 6184 32524
rect 6236 32512 6242 32564
rect 8202 32552 8208 32564
rect 8163 32524 8208 32552
rect 8202 32512 8208 32524
rect 8260 32512 8266 32564
rect 15470 32512 15476 32564
rect 15528 32552 15534 32564
rect 17037 32555 17095 32561
rect 17037 32552 17049 32555
rect 15528 32524 17049 32552
rect 15528 32512 15534 32524
rect 17037 32521 17049 32524
rect 17083 32521 17095 32555
rect 19978 32552 19984 32564
rect 17037 32515 17095 32521
rect 17144 32524 19984 32552
rect 3418 32484 3424 32496
rect 1964 32456 3424 32484
rect 1964 32357 1992 32456
rect 3418 32444 3424 32456
rect 3476 32444 3482 32496
rect 11054 32444 11060 32496
rect 11112 32484 11118 32496
rect 12434 32484 12440 32496
rect 11112 32456 12440 32484
rect 11112 32444 11118 32456
rect 12434 32444 12440 32456
rect 12492 32484 12498 32496
rect 12710 32484 12716 32496
rect 12492 32456 12716 32484
rect 12492 32444 12498 32456
rect 12710 32444 12716 32456
rect 12768 32444 12774 32496
rect 13265 32487 13323 32493
rect 13265 32453 13277 32487
rect 13311 32484 13323 32487
rect 13311 32456 15332 32484
rect 13311 32453 13323 32456
rect 13265 32447 13323 32453
rect 2501 32419 2559 32425
rect 2501 32385 2513 32419
rect 2547 32416 2559 32419
rect 3142 32416 3148 32428
rect 2547 32388 3148 32416
rect 2547 32385 2559 32388
rect 2501 32379 2559 32385
rect 3142 32376 3148 32388
rect 3200 32376 3206 32428
rect 3329 32419 3387 32425
rect 3329 32385 3341 32419
rect 3375 32416 3387 32419
rect 5626 32416 5632 32428
rect 3375 32388 4200 32416
rect 3375 32385 3387 32388
rect 3329 32379 3387 32385
rect 1949 32351 2007 32357
rect 1949 32317 1961 32351
rect 1995 32317 2007 32351
rect 1949 32311 2007 32317
rect 2148 32320 2636 32348
rect 1765 32283 1823 32289
rect 1765 32249 1777 32283
rect 1811 32280 1823 32283
rect 1854 32280 1860 32292
rect 1811 32252 1860 32280
rect 1811 32249 1823 32252
rect 1765 32243 1823 32249
rect 1854 32240 1860 32252
rect 1912 32240 1918 32292
rect 2148 32289 2176 32320
rect 2133 32283 2191 32289
rect 2133 32249 2145 32283
rect 2179 32249 2191 32283
rect 2608 32280 2636 32320
rect 2774 32308 2780 32360
rect 2832 32348 2838 32360
rect 2961 32351 3019 32357
rect 2961 32348 2973 32351
rect 2832 32320 2973 32348
rect 2832 32308 2838 32320
rect 2961 32317 2973 32320
rect 3007 32317 3019 32351
rect 2961 32311 3019 32317
rect 3050 32308 3056 32360
rect 3108 32348 3114 32360
rect 4172 32357 4200 32388
rect 5368 32388 5632 32416
rect 3513 32351 3571 32357
rect 3513 32348 3525 32351
rect 3108 32320 3525 32348
rect 3108 32308 3114 32320
rect 3513 32317 3525 32320
rect 3559 32317 3571 32351
rect 3513 32311 3571 32317
rect 4157 32351 4215 32357
rect 4157 32317 4169 32351
rect 4203 32317 4215 32351
rect 4157 32311 4215 32317
rect 4801 32351 4859 32357
rect 4801 32317 4813 32351
rect 4847 32348 4859 32351
rect 5074 32348 5080 32360
rect 4847 32320 5080 32348
rect 4847 32317 4859 32320
rect 4801 32311 4859 32317
rect 4249 32283 4307 32289
rect 4249 32280 4261 32283
rect 2608 32252 4261 32280
rect 2133 32243 2191 32249
rect 4249 32249 4261 32252
rect 4295 32280 4307 32283
rect 4816 32280 4844 32311
rect 5074 32308 5080 32320
rect 5132 32308 5138 32360
rect 5368 32357 5396 32388
rect 5626 32376 5632 32388
rect 5684 32376 5690 32428
rect 8570 32376 8576 32428
rect 8628 32416 8634 32428
rect 9217 32419 9275 32425
rect 9217 32416 9229 32419
rect 8628 32388 9229 32416
rect 8628 32376 8634 32388
rect 9217 32385 9229 32388
rect 9263 32385 9275 32419
rect 9217 32379 9275 32385
rect 9674 32376 9680 32428
rect 9732 32416 9738 32428
rect 10597 32419 10655 32425
rect 10597 32416 10609 32419
rect 9732 32388 10609 32416
rect 9732 32376 9738 32388
rect 10597 32385 10609 32388
rect 10643 32416 10655 32419
rect 12618 32416 12624 32428
rect 10643 32388 12624 32416
rect 10643 32385 10655 32388
rect 10597 32379 10655 32385
rect 12618 32376 12624 32388
rect 12676 32376 12682 32428
rect 5353 32351 5411 32357
rect 5353 32348 5365 32351
rect 5184 32320 5365 32348
rect 4295 32252 4844 32280
rect 4295 32249 4307 32252
rect 4249 32243 4307 32249
rect 2041 32215 2099 32221
rect 2041 32181 2053 32215
rect 2087 32212 2099 32215
rect 3326 32212 3332 32224
rect 2087 32184 3332 32212
rect 2087 32181 2099 32184
rect 2041 32175 2099 32181
rect 3326 32172 3332 32184
rect 3384 32172 3390 32224
rect 4706 32172 4712 32224
rect 4764 32212 4770 32224
rect 5184 32212 5212 32320
rect 5353 32317 5365 32320
rect 5399 32317 5411 32351
rect 5534 32348 5540 32360
rect 5495 32320 5540 32348
rect 5353 32311 5411 32317
rect 5534 32308 5540 32320
rect 5592 32308 5598 32360
rect 6089 32351 6147 32357
rect 6089 32317 6101 32351
rect 6135 32317 6147 32351
rect 6089 32311 6147 32317
rect 5258 32240 5264 32292
rect 5316 32280 5322 32292
rect 6104 32280 6132 32311
rect 6730 32308 6736 32360
rect 6788 32348 6794 32360
rect 6825 32351 6883 32357
rect 6825 32348 6837 32351
rect 6788 32320 6837 32348
rect 6788 32308 6794 32320
rect 6825 32317 6837 32320
rect 6871 32317 6883 32351
rect 7098 32348 7104 32360
rect 7059 32320 7104 32348
rect 6825 32311 6883 32317
rect 7098 32308 7104 32320
rect 7156 32308 7162 32360
rect 8941 32351 8999 32357
rect 8941 32317 8953 32351
rect 8987 32348 8999 32351
rect 9306 32348 9312 32360
rect 8987 32320 9312 32348
rect 8987 32317 8999 32320
rect 8941 32311 8999 32317
rect 9306 32308 9312 32320
rect 9364 32308 9370 32360
rect 11514 32308 11520 32360
rect 11572 32348 11578 32360
rect 11609 32351 11667 32357
rect 11609 32348 11621 32351
rect 11572 32320 11621 32348
rect 11572 32308 11578 32320
rect 11609 32317 11621 32320
rect 11655 32317 11667 32351
rect 12526 32348 12532 32360
rect 12439 32320 12532 32348
rect 11609 32311 11667 32317
rect 12526 32308 12532 32320
rect 12584 32348 12590 32360
rect 12894 32348 12900 32360
rect 12584 32320 12900 32348
rect 12584 32308 12590 32320
rect 12894 32308 12900 32320
rect 12952 32308 12958 32360
rect 5316 32252 6132 32280
rect 5316 32240 5322 32252
rect 10410 32240 10416 32292
rect 10468 32280 10474 32292
rect 13280 32280 13308 32447
rect 13633 32419 13691 32425
rect 13633 32385 13645 32419
rect 13679 32416 13691 32419
rect 13814 32416 13820 32428
rect 13679 32388 13820 32416
rect 13679 32385 13691 32388
rect 13633 32379 13691 32385
rect 13814 32376 13820 32388
rect 13872 32376 13878 32428
rect 14274 32416 14280 32428
rect 14016 32388 14280 32416
rect 14016 32357 14044 32388
rect 14274 32376 14280 32388
rect 14332 32416 14338 32428
rect 14826 32416 14832 32428
rect 14332 32388 14832 32416
rect 14332 32376 14338 32388
rect 14826 32376 14832 32388
rect 14884 32376 14890 32428
rect 14001 32351 14059 32357
rect 14001 32317 14013 32351
rect 14047 32317 14059 32351
rect 14366 32348 14372 32360
rect 14327 32320 14372 32348
rect 14001 32311 14059 32317
rect 14366 32308 14372 32320
rect 14424 32308 14430 32360
rect 14550 32348 14556 32360
rect 14511 32320 14556 32348
rect 14550 32308 14556 32320
rect 14608 32308 14614 32360
rect 14921 32351 14979 32357
rect 14921 32317 14933 32351
rect 14967 32317 14979 32351
rect 15304 32348 15332 32456
rect 15378 32376 15384 32428
rect 15436 32416 15442 32428
rect 15654 32416 15660 32428
rect 15436 32388 15660 32416
rect 15436 32376 15442 32388
rect 15654 32376 15660 32388
rect 15712 32376 15718 32428
rect 15930 32416 15936 32428
rect 15891 32388 15936 32416
rect 15930 32376 15936 32388
rect 15988 32376 15994 32428
rect 16390 32376 16396 32428
rect 16448 32416 16454 32428
rect 17144 32416 17172 32524
rect 19978 32512 19984 32524
rect 20036 32512 20042 32564
rect 21726 32512 21732 32564
rect 21784 32552 21790 32564
rect 23474 32552 23480 32564
rect 21784 32524 23480 32552
rect 21784 32512 21790 32524
rect 23474 32512 23480 32524
rect 23532 32512 23538 32564
rect 23566 32512 23572 32564
rect 23624 32552 23630 32564
rect 24489 32555 24547 32561
rect 24489 32552 24501 32555
rect 23624 32524 24501 32552
rect 23624 32512 23630 32524
rect 24489 32521 24501 32524
rect 24535 32521 24547 32555
rect 24489 32515 24547 32521
rect 29362 32512 29368 32564
rect 29420 32552 29426 32564
rect 39022 32552 39028 32564
rect 29420 32524 31616 32552
rect 38983 32524 39028 32552
rect 29420 32512 29426 32524
rect 17494 32444 17500 32496
rect 17552 32484 17558 32496
rect 18877 32487 18935 32493
rect 18877 32484 18889 32487
rect 17552 32456 18889 32484
rect 17552 32444 17558 32456
rect 18877 32453 18889 32456
rect 18923 32453 18935 32487
rect 19150 32484 19156 32496
rect 18877 32447 18935 32453
rect 18984 32456 19156 32484
rect 18984 32416 19012 32456
rect 19150 32444 19156 32456
rect 19208 32444 19214 32496
rect 26786 32484 26792 32496
rect 19260 32456 26792 32484
rect 16448 32388 17172 32416
rect 17236 32388 19012 32416
rect 16448 32376 16454 32388
rect 17236 32348 17264 32388
rect 15304 32320 17264 32348
rect 18233 32351 18291 32357
rect 14921 32311 14979 32317
rect 18233 32317 18245 32351
rect 18279 32317 18291 32351
rect 18598 32348 18604 32360
rect 18559 32320 18604 32348
rect 18233 32311 18291 32317
rect 10468 32252 13308 32280
rect 10468 32240 10474 32252
rect 14458 32240 14464 32292
rect 14516 32280 14522 32292
rect 14936 32280 14964 32311
rect 14516 32252 14964 32280
rect 14516 32240 14522 32252
rect 4764 32184 5212 32212
rect 4764 32172 4770 32184
rect 6638 32172 6644 32224
rect 6696 32212 6702 32224
rect 9490 32212 9496 32224
rect 6696 32184 9496 32212
rect 6696 32172 6702 32184
rect 9490 32172 9496 32184
rect 9548 32172 9554 32224
rect 11790 32212 11796 32224
rect 11751 32184 11796 32212
rect 11790 32172 11796 32184
rect 11848 32172 11854 32224
rect 18248 32212 18276 32311
rect 18598 32308 18604 32320
rect 18656 32308 18662 32360
rect 18969 32351 19027 32357
rect 18969 32317 18981 32351
rect 19015 32348 19027 32351
rect 19260 32348 19288 32456
rect 26786 32444 26792 32456
rect 26844 32444 26850 32496
rect 29086 32484 29092 32496
rect 27816 32456 29092 32484
rect 20070 32376 20076 32428
rect 20128 32416 20134 32428
rect 20441 32419 20499 32425
rect 20441 32416 20453 32419
rect 20128 32388 20453 32416
rect 20128 32376 20134 32388
rect 20441 32385 20453 32388
rect 20487 32385 20499 32419
rect 20441 32379 20499 32385
rect 21174 32376 21180 32428
rect 21232 32416 21238 32428
rect 22557 32419 22615 32425
rect 22557 32416 22569 32419
rect 21232 32388 22569 32416
rect 21232 32376 21238 32388
rect 22557 32385 22569 32388
rect 22603 32385 22615 32419
rect 27816 32416 27844 32456
rect 29086 32444 29092 32456
rect 29144 32444 29150 32496
rect 22557 32379 22615 32385
rect 27724 32388 27844 32416
rect 19015 32320 19288 32348
rect 19015 32317 19027 32320
rect 18969 32311 19027 32317
rect 19334 32308 19340 32360
rect 19392 32348 19398 32360
rect 19613 32351 19671 32357
rect 19613 32348 19625 32351
rect 19392 32320 19625 32348
rect 19392 32308 19398 32320
rect 19613 32317 19625 32320
rect 19659 32317 19671 32351
rect 19613 32311 19671 32317
rect 20349 32351 20407 32357
rect 20349 32317 20361 32351
rect 20395 32348 20407 32351
rect 21818 32348 21824 32360
rect 20395 32320 21824 32348
rect 20395 32317 20407 32320
rect 20349 32311 20407 32317
rect 21818 32308 21824 32320
rect 21876 32308 21882 32360
rect 21913 32351 21971 32357
rect 21913 32317 21925 32351
rect 21959 32317 21971 32351
rect 21913 32311 21971 32317
rect 20254 32280 20260 32292
rect 19628 32252 20260 32280
rect 19628 32212 19656 32252
rect 20254 32240 20260 32252
rect 20312 32240 20318 32292
rect 21928 32280 21956 32311
rect 22094 32308 22100 32360
rect 22152 32348 22158 32360
rect 22465 32351 22523 32357
rect 22465 32348 22477 32351
rect 22152 32320 22477 32348
rect 22152 32308 22158 32320
rect 22465 32317 22477 32320
rect 22511 32348 22523 32351
rect 23566 32348 23572 32360
rect 22511 32320 23572 32348
rect 22511 32317 22523 32320
rect 22465 32311 22523 32317
rect 23566 32308 23572 32320
rect 23624 32308 23630 32360
rect 23661 32351 23719 32357
rect 23661 32317 23673 32351
rect 23707 32317 23719 32351
rect 23661 32311 23719 32317
rect 22186 32280 22192 32292
rect 21928 32252 22192 32280
rect 22186 32240 22192 32252
rect 22244 32280 22250 32292
rect 23676 32280 23704 32311
rect 23842 32308 23848 32360
rect 23900 32348 23906 32360
rect 24394 32348 24400 32360
rect 23900 32320 24400 32348
rect 23900 32308 23906 32320
rect 24394 32308 24400 32320
rect 24452 32308 24458 32360
rect 25314 32348 25320 32360
rect 25275 32320 25320 32348
rect 25314 32308 25320 32320
rect 25372 32308 25378 32360
rect 25593 32351 25651 32357
rect 25593 32317 25605 32351
rect 25639 32317 25651 32351
rect 27154 32348 27160 32360
rect 27115 32320 27160 32348
rect 25593 32311 25651 32317
rect 22244 32252 23704 32280
rect 22244 32240 22250 32252
rect 23750 32240 23756 32292
rect 23808 32280 23814 32292
rect 25608 32280 25636 32311
rect 27154 32308 27160 32320
rect 27212 32308 27218 32360
rect 27338 32348 27344 32360
rect 27299 32320 27344 32348
rect 27338 32308 27344 32320
rect 27396 32308 27402 32360
rect 27724 32357 27752 32388
rect 30374 32376 30380 32428
rect 30432 32416 30438 32428
rect 31588 32425 31616 32524
rect 39022 32512 39028 32524
rect 39080 32512 39086 32564
rect 35342 32444 35348 32496
rect 35400 32484 35406 32496
rect 35713 32487 35771 32493
rect 35713 32484 35725 32487
rect 35400 32456 35725 32484
rect 35400 32444 35406 32456
rect 35713 32453 35725 32456
rect 35759 32453 35771 32487
rect 35713 32447 35771 32453
rect 30837 32419 30895 32425
rect 30837 32416 30849 32419
rect 30432 32388 30849 32416
rect 30432 32376 30438 32388
rect 30837 32385 30849 32388
rect 30883 32385 30895 32419
rect 30837 32379 30895 32385
rect 31573 32419 31631 32425
rect 31573 32385 31585 32419
rect 31619 32385 31631 32419
rect 36906 32416 36912 32428
rect 36867 32388 36912 32416
rect 31573 32379 31631 32385
rect 36906 32376 36912 32388
rect 36964 32376 36970 32428
rect 37918 32416 37924 32428
rect 37292 32388 37924 32416
rect 27709 32351 27767 32357
rect 27709 32317 27721 32351
rect 27755 32317 27767 32351
rect 27890 32348 27896 32360
rect 27851 32320 27896 32348
rect 27709 32311 27767 32317
rect 27890 32308 27896 32320
rect 27948 32308 27954 32360
rect 28353 32351 28411 32357
rect 28353 32317 28365 32351
rect 28399 32317 28411 32351
rect 28353 32311 28411 32317
rect 29457 32351 29515 32357
rect 29457 32317 29469 32351
rect 29503 32348 29515 32351
rect 29546 32348 29552 32360
rect 29503 32320 29552 32348
rect 29503 32317 29515 32320
rect 29457 32311 29515 32317
rect 26050 32280 26056 32292
rect 23808 32252 25176 32280
rect 25608 32252 26056 32280
rect 23808 32240 23814 32252
rect 18248 32184 19656 32212
rect 19705 32215 19763 32221
rect 19705 32181 19717 32215
rect 19751 32212 19763 32215
rect 20070 32212 20076 32224
rect 19751 32184 20076 32212
rect 19751 32181 19763 32184
rect 19705 32175 19763 32181
rect 20070 32172 20076 32184
rect 20128 32172 20134 32224
rect 21821 32215 21879 32221
rect 21821 32181 21833 32215
rect 21867 32212 21879 32215
rect 22278 32212 22284 32224
rect 21867 32184 22284 32212
rect 21867 32181 21879 32184
rect 21821 32175 21879 32181
rect 22278 32172 22284 32184
rect 22336 32172 22342 32224
rect 22554 32172 22560 32224
rect 22612 32212 22618 32224
rect 25148 32221 25176 32252
rect 26050 32240 26056 32252
rect 26108 32280 26114 32292
rect 28368 32280 28396 32311
rect 26108 32252 28396 32280
rect 26108 32240 26114 32252
rect 28994 32240 29000 32292
rect 29052 32280 29058 32292
rect 29472 32280 29500 32311
rect 29546 32308 29552 32320
rect 29604 32308 29610 32360
rect 29733 32351 29791 32357
rect 29733 32317 29745 32351
rect 29779 32348 29791 32351
rect 31662 32348 31668 32360
rect 29779 32320 30788 32348
rect 31623 32320 31668 32348
rect 29779 32317 29791 32320
rect 29733 32311 29791 32317
rect 29052 32252 29500 32280
rect 30760 32280 30788 32320
rect 31662 32308 31668 32320
rect 31720 32308 31726 32360
rect 32769 32351 32827 32357
rect 32769 32317 32781 32351
rect 32815 32317 32827 32351
rect 32950 32348 32956 32360
rect 32911 32320 32956 32348
rect 32769 32311 32827 32317
rect 32125 32283 32183 32289
rect 32125 32280 32137 32283
rect 30760 32252 32137 32280
rect 29052 32240 29058 32252
rect 32125 32249 32137 32252
rect 32171 32249 32183 32283
rect 32784 32280 32812 32311
rect 32950 32308 32956 32320
rect 33008 32308 33014 32360
rect 33318 32348 33324 32360
rect 33279 32320 33324 32348
rect 33318 32308 33324 32320
rect 33376 32308 33382 32360
rect 33778 32308 33784 32360
rect 33836 32348 33842 32360
rect 34885 32351 34943 32357
rect 34885 32348 34897 32351
rect 33836 32320 34897 32348
rect 33836 32308 33842 32320
rect 34885 32317 34897 32320
rect 34931 32317 34943 32351
rect 34885 32311 34943 32317
rect 35345 32351 35403 32357
rect 35345 32317 35357 32351
rect 35391 32317 35403 32351
rect 35802 32348 35808 32360
rect 35763 32320 35808 32348
rect 35345 32311 35403 32317
rect 33226 32280 33232 32292
rect 32784 32252 33232 32280
rect 32125 32243 32183 32249
rect 33226 32240 33232 32252
rect 33284 32240 33290 32292
rect 34514 32240 34520 32292
rect 34572 32280 34578 32292
rect 35360 32280 35388 32311
rect 35802 32308 35808 32320
rect 35860 32308 35866 32360
rect 36630 32348 36636 32360
rect 36591 32320 36636 32348
rect 36630 32308 36636 32320
rect 36688 32308 36694 32360
rect 34572 32252 35388 32280
rect 36449 32283 36507 32289
rect 34572 32240 34578 32252
rect 36449 32249 36461 32283
rect 36495 32280 36507 32283
rect 36538 32280 36544 32292
rect 36495 32252 36544 32280
rect 36495 32249 36507 32252
rect 36449 32243 36507 32249
rect 36538 32240 36544 32252
rect 36596 32280 36602 32292
rect 37292 32280 37320 32388
rect 37918 32376 37924 32388
rect 37976 32376 37982 32428
rect 37458 32348 37464 32360
rect 37419 32320 37464 32348
rect 37458 32308 37464 32320
rect 37516 32308 37522 32360
rect 37734 32348 37740 32360
rect 37695 32320 37740 32348
rect 37734 32308 37740 32320
rect 37792 32308 37798 32360
rect 36596 32252 37320 32280
rect 36596 32240 36602 32252
rect 23845 32215 23903 32221
rect 23845 32212 23857 32215
rect 22612 32184 23857 32212
rect 22612 32172 22618 32184
rect 23845 32181 23857 32184
rect 23891 32181 23903 32215
rect 23845 32175 23903 32181
rect 25133 32215 25191 32221
rect 25133 32181 25145 32215
rect 25179 32181 25191 32215
rect 25133 32175 25191 32181
rect 25222 32172 25228 32224
rect 25280 32212 25286 32224
rect 26789 32215 26847 32221
rect 26789 32212 26801 32215
rect 25280 32184 26801 32212
rect 25280 32172 25286 32184
rect 26789 32181 26801 32184
rect 26835 32181 26847 32215
rect 26789 32175 26847 32181
rect 27338 32172 27344 32224
rect 27396 32212 27402 32224
rect 28537 32215 28595 32221
rect 28537 32212 28549 32215
rect 27396 32184 28549 32212
rect 27396 32172 27402 32184
rect 28537 32181 28549 32184
rect 28583 32181 28595 32215
rect 28537 32175 28595 32181
rect 30006 32172 30012 32224
rect 30064 32212 30070 32224
rect 33502 32212 33508 32224
rect 30064 32184 33508 32212
rect 30064 32172 30070 32184
rect 33502 32172 33508 32184
rect 33560 32172 33566 32224
rect 1104 32122 39836 32144
rect 1104 32070 19606 32122
rect 19658 32070 19670 32122
rect 19722 32070 19734 32122
rect 19786 32070 19798 32122
rect 19850 32070 39836 32122
rect 1104 32048 39836 32070
rect 2682 32008 2688 32020
rect 1412 31980 2688 32008
rect 1412 31884 1440 31980
rect 2682 31968 2688 31980
rect 2740 32008 2746 32020
rect 3697 32011 3755 32017
rect 3697 32008 3709 32011
rect 2740 31980 3709 32008
rect 2740 31968 2746 31980
rect 3697 31977 3709 31980
rect 3743 31977 3755 32011
rect 3697 31971 3755 31977
rect 1394 31872 1400 31884
rect 1307 31844 1400 31872
rect 1394 31832 1400 31844
rect 1452 31832 1458 31884
rect 1670 31804 1676 31816
rect 1631 31776 1676 31804
rect 1670 31764 1676 31776
rect 1728 31764 1734 31816
rect 3712 31804 3740 31971
rect 5074 31968 5080 32020
rect 5132 32008 5138 32020
rect 5132 31980 5488 32008
rect 5132 31968 5138 31980
rect 4341 31943 4399 31949
rect 4341 31909 4353 31943
rect 4387 31940 4399 31943
rect 4614 31940 4620 31952
rect 4387 31912 4620 31940
rect 4387 31909 4399 31912
rect 4341 31903 4399 31909
rect 4614 31900 4620 31912
rect 4672 31900 4678 31952
rect 3878 31872 3884 31884
rect 3839 31844 3884 31872
rect 3878 31832 3884 31844
rect 3936 31832 3942 31884
rect 4706 31832 4712 31884
rect 4764 31872 4770 31884
rect 4801 31875 4859 31881
rect 4801 31872 4813 31875
rect 4764 31844 4813 31872
rect 4764 31832 4770 31844
rect 4801 31841 4813 31844
rect 4847 31841 4859 31875
rect 4982 31872 4988 31884
rect 4943 31844 4988 31872
rect 4801 31835 4859 31841
rect 4982 31832 4988 31844
rect 5040 31832 5046 31884
rect 5166 31872 5172 31884
rect 5127 31844 5172 31872
rect 5166 31832 5172 31844
rect 5224 31832 5230 31884
rect 5258 31832 5264 31884
rect 5316 31872 5322 31884
rect 5353 31875 5411 31881
rect 5353 31872 5365 31875
rect 5316 31844 5365 31872
rect 5316 31832 5322 31844
rect 5353 31841 5365 31844
rect 5399 31841 5411 31875
rect 5460 31872 5488 31980
rect 7098 31968 7104 32020
rect 7156 32008 7162 32020
rect 7193 32011 7251 32017
rect 7193 32008 7205 32011
rect 7156 31980 7205 32008
rect 7156 31968 7162 31980
rect 7193 31977 7205 31980
rect 7239 31977 7251 32011
rect 7193 31971 7251 31977
rect 9033 32011 9091 32017
rect 9033 31977 9045 32011
rect 9079 32008 9091 32011
rect 9079 31980 10916 32008
rect 9079 31977 9091 31980
rect 9033 31971 9091 31977
rect 6270 31900 6276 31952
rect 6328 31940 6334 31952
rect 6328 31912 7144 31940
rect 6328 31900 6334 31912
rect 5629 31875 5687 31881
rect 5629 31872 5641 31875
rect 5460 31844 5641 31872
rect 5353 31835 5411 31841
rect 5629 31841 5641 31844
rect 5675 31841 5687 31875
rect 5629 31835 5687 31841
rect 6549 31875 6607 31881
rect 6549 31841 6561 31875
rect 6595 31841 6607 31875
rect 6914 31872 6920 31884
rect 6875 31844 6920 31872
rect 6549 31835 6607 31841
rect 5184 31804 5212 31832
rect 5442 31804 5448 31816
rect 3712 31776 4844 31804
rect 5184 31776 5448 31804
rect 4816 31748 4844 31776
rect 5442 31764 5448 31776
rect 5500 31764 5506 31816
rect 6564 31804 6592 31835
rect 6914 31832 6920 31844
rect 6972 31832 6978 31884
rect 7116 31881 7144 31912
rect 9490 31900 9496 31952
rect 9548 31940 9554 31952
rect 9548 31912 9720 31940
rect 9548 31900 9554 31912
rect 7101 31875 7159 31881
rect 7101 31841 7113 31875
rect 7147 31841 7159 31875
rect 7101 31835 7159 31841
rect 8205 31875 8263 31881
rect 8205 31841 8217 31875
rect 8251 31872 8263 31875
rect 8754 31872 8760 31884
rect 8251 31844 8760 31872
rect 8251 31841 8263 31844
rect 8205 31835 8263 31841
rect 8754 31832 8760 31844
rect 8812 31832 8818 31884
rect 8849 31875 8907 31881
rect 8849 31841 8861 31875
rect 8895 31872 8907 31875
rect 9582 31872 9588 31884
rect 8895 31844 9588 31872
rect 8895 31841 8907 31844
rect 8849 31835 8907 31841
rect 9582 31832 9588 31844
rect 9640 31832 9646 31884
rect 9692 31881 9720 31912
rect 10888 31884 10916 31980
rect 11790 31968 11796 32020
rect 11848 32008 11854 32020
rect 17862 32008 17868 32020
rect 11848 31980 12664 32008
rect 11848 31968 11854 31980
rect 9677 31875 9735 31881
rect 9677 31841 9689 31875
rect 9723 31841 9735 31875
rect 9677 31835 9735 31841
rect 10045 31875 10103 31881
rect 10045 31841 10057 31875
rect 10091 31841 10103 31875
rect 10502 31872 10508 31884
rect 10463 31844 10508 31872
rect 10045 31835 10103 31841
rect 7006 31804 7012 31816
rect 6564 31776 7012 31804
rect 7006 31764 7012 31776
rect 7064 31764 7070 31816
rect 8297 31807 8355 31813
rect 8297 31773 8309 31807
rect 8343 31804 8355 31807
rect 10060 31804 10088 31835
rect 10502 31832 10508 31844
rect 10560 31832 10566 31884
rect 10870 31832 10876 31884
rect 10928 31872 10934 31884
rect 12250 31872 12256 31884
rect 10928 31844 12020 31872
rect 12211 31844 12256 31872
rect 10928 31832 10934 31844
rect 11992 31816 12020 31844
rect 12250 31832 12256 31844
rect 12308 31832 12314 31884
rect 12636 31881 12664 31980
rect 16224 31980 17868 32008
rect 12710 31900 12716 31952
rect 12768 31940 12774 31952
rect 15654 31940 15660 31952
rect 12768 31912 13400 31940
rect 12768 31900 12774 31912
rect 13372 31881 13400 31912
rect 14568 31912 15660 31940
rect 14568 31881 14596 31912
rect 15654 31900 15660 31912
rect 15712 31900 15718 31952
rect 12621 31875 12679 31881
rect 12621 31841 12633 31875
rect 12667 31841 12679 31875
rect 12621 31835 12679 31841
rect 13173 31875 13231 31881
rect 13173 31841 13185 31875
rect 13219 31841 13231 31875
rect 13173 31835 13231 31841
rect 13357 31875 13415 31881
rect 13357 31841 13369 31875
rect 13403 31841 13415 31875
rect 13357 31835 13415 31841
rect 14553 31875 14611 31881
rect 14553 31841 14565 31875
rect 14599 31841 14611 31875
rect 14553 31835 14611 31841
rect 15289 31875 15347 31881
rect 15289 31841 15301 31875
rect 15335 31872 15347 31875
rect 15470 31872 15476 31884
rect 15335 31844 15476 31872
rect 15335 31841 15347 31844
rect 15289 31835 15347 31841
rect 8343 31776 10088 31804
rect 8343 31773 8355 31776
rect 8297 31767 8355 31773
rect 10410 31764 10416 31816
rect 10468 31804 10474 31816
rect 11701 31807 11759 31813
rect 11701 31804 11713 31807
rect 10468 31776 11713 31804
rect 10468 31764 10474 31776
rect 11701 31773 11713 31776
rect 11747 31773 11759 31807
rect 11701 31767 11759 31773
rect 11974 31764 11980 31816
rect 12032 31764 12038 31816
rect 12069 31807 12127 31813
rect 12069 31773 12081 31807
rect 12115 31804 12127 31807
rect 12434 31804 12440 31816
rect 12115 31776 12440 31804
rect 12115 31773 12127 31776
rect 12069 31767 12127 31773
rect 12434 31764 12440 31776
rect 12492 31764 12498 31816
rect 13188 31804 13216 31835
rect 15470 31832 15476 31844
rect 15528 31832 15534 31884
rect 16224 31881 16252 31980
rect 17862 31968 17868 31980
rect 17920 31968 17926 32020
rect 18782 32008 18788 32020
rect 18524 31980 18788 32008
rect 17126 31940 17132 31952
rect 16684 31912 17132 31940
rect 16684 31881 16712 31912
rect 17126 31900 17132 31912
rect 17184 31900 17190 31952
rect 18414 31940 18420 31952
rect 17604 31912 18276 31940
rect 18375 31912 18420 31940
rect 16209 31875 16267 31881
rect 16209 31841 16221 31875
rect 16255 31841 16267 31875
rect 16209 31835 16267 31841
rect 16669 31875 16727 31881
rect 16669 31841 16681 31875
rect 16715 31841 16727 31875
rect 16669 31835 16727 31841
rect 17037 31875 17095 31881
rect 17037 31841 17049 31875
rect 17083 31841 17095 31875
rect 17218 31872 17224 31884
rect 17179 31844 17224 31872
rect 17037 31835 17095 31841
rect 14458 31804 14464 31816
rect 12544 31776 14464 31804
rect 4798 31696 4804 31748
rect 4856 31696 4862 31748
rect 9766 31736 9772 31748
rect 9727 31708 9772 31736
rect 9766 31696 9772 31708
rect 9824 31696 9830 31748
rect 11992 31736 12020 31764
rect 12544 31736 12572 31776
rect 14458 31764 14464 31776
rect 14516 31764 14522 31816
rect 14645 31807 14703 31813
rect 14645 31773 14657 31807
rect 14691 31804 14703 31807
rect 15194 31804 15200 31816
rect 14691 31776 15200 31804
rect 14691 31773 14703 31776
rect 14645 31767 14703 31773
rect 15194 31764 15200 31776
rect 15252 31764 15258 31816
rect 16301 31807 16359 31813
rect 16301 31773 16313 31807
rect 16347 31804 16359 31807
rect 16942 31804 16948 31816
rect 16347 31776 16948 31804
rect 16347 31773 16359 31776
rect 16301 31767 16359 31773
rect 16942 31764 16948 31776
rect 17000 31764 17006 31816
rect 17052 31804 17080 31835
rect 17218 31832 17224 31844
rect 17276 31832 17282 31884
rect 17604 31816 17632 31912
rect 17957 31875 18015 31881
rect 17957 31841 17969 31875
rect 18003 31841 18015 31875
rect 18248 31872 18276 31912
rect 18414 31900 18420 31912
rect 18472 31900 18478 31952
rect 18524 31872 18552 31980
rect 18782 31968 18788 31980
rect 18840 32008 18846 32020
rect 19426 32008 19432 32020
rect 18840 31980 19432 32008
rect 18840 31968 18846 31980
rect 19426 31968 19432 31980
rect 19484 31968 19490 32020
rect 22557 32011 22615 32017
rect 22557 31977 22569 32011
rect 22603 32008 22615 32011
rect 23934 32008 23940 32020
rect 22603 31980 23940 32008
rect 22603 31977 22615 31980
rect 22557 31971 22615 31977
rect 23934 31968 23940 31980
rect 23992 31968 23998 32020
rect 33778 32008 33784 32020
rect 29564 31980 33784 32008
rect 18598 31900 18604 31952
rect 18656 31940 18662 31952
rect 19242 31940 19248 31952
rect 18656 31912 19248 31940
rect 18656 31900 18662 31912
rect 19242 31900 19248 31912
rect 19300 31900 19306 31952
rect 24302 31940 24308 31952
rect 21836 31912 24308 31940
rect 18248 31844 18552 31872
rect 18693 31875 18751 31881
rect 17957 31835 18015 31841
rect 18693 31841 18705 31875
rect 18739 31872 18751 31875
rect 18874 31872 18880 31884
rect 18739 31844 18880 31872
rect 18739 31841 18751 31844
rect 18693 31835 18751 31841
rect 17586 31804 17592 31816
rect 17052 31776 17592 31804
rect 17586 31764 17592 31776
rect 17644 31764 17650 31816
rect 17972 31804 18000 31835
rect 18874 31832 18880 31844
rect 18932 31832 18938 31884
rect 18966 31832 18972 31884
rect 19024 31872 19030 31884
rect 19334 31872 19340 31884
rect 19024 31844 19069 31872
rect 19168 31844 19340 31872
rect 19024 31832 19030 31844
rect 19168 31804 19196 31844
rect 19334 31832 19340 31844
rect 19392 31832 19398 31884
rect 19426 31832 19432 31884
rect 19484 31872 19490 31884
rect 19889 31875 19947 31881
rect 19484 31844 19529 31872
rect 19484 31832 19490 31844
rect 19889 31841 19901 31875
rect 19935 31872 19947 31875
rect 19978 31872 19984 31884
rect 19935 31844 19984 31872
rect 19935 31841 19947 31844
rect 19889 31835 19947 31841
rect 19978 31832 19984 31844
rect 20036 31832 20042 31884
rect 20346 31872 20352 31884
rect 20259 31844 20352 31872
rect 20346 31832 20352 31844
rect 20404 31872 20410 31884
rect 20990 31872 20996 31884
rect 20404 31844 20996 31872
rect 20404 31832 20410 31844
rect 20990 31832 20996 31844
rect 21048 31832 21054 31884
rect 21266 31872 21272 31884
rect 21227 31844 21272 31872
rect 21266 31832 21272 31844
rect 21324 31832 21330 31884
rect 21836 31881 21864 31912
rect 24302 31900 24308 31912
rect 24360 31900 24366 31952
rect 24762 31900 24768 31952
rect 24820 31940 24826 31952
rect 24820 31912 27016 31940
rect 24820 31900 24826 31912
rect 21821 31875 21879 31881
rect 21821 31841 21833 31875
rect 21867 31841 21879 31875
rect 22462 31872 22468 31884
rect 22423 31844 22468 31872
rect 21821 31835 21879 31841
rect 22462 31832 22468 31844
rect 22520 31832 22526 31884
rect 23658 31872 23664 31884
rect 23619 31844 23664 31872
rect 23658 31832 23664 31844
rect 23716 31832 23722 31884
rect 24029 31875 24087 31881
rect 24029 31841 24041 31875
rect 24075 31872 24087 31875
rect 25222 31872 25228 31884
rect 24075 31844 25228 31872
rect 24075 31841 24087 31844
rect 24029 31835 24087 31841
rect 25222 31832 25228 31844
rect 25280 31832 25286 31884
rect 25409 31875 25467 31881
rect 25409 31841 25421 31875
rect 25455 31841 25467 31875
rect 25409 31835 25467 31841
rect 17972 31776 19196 31804
rect 21085 31807 21143 31813
rect 21085 31773 21097 31807
rect 21131 31804 21143 31807
rect 22002 31804 22008 31816
rect 21131 31776 22008 31804
rect 21131 31773 21143 31776
rect 21085 31767 21143 31773
rect 22002 31764 22008 31776
rect 22060 31764 22066 31816
rect 23290 31804 23296 31816
rect 23251 31776 23296 31804
rect 23290 31764 23296 31776
rect 23348 31764 23354 31816
rect 23566 31764 23572 31816
rect 23624 31804 23630 31816
rect 24765 31807 24823 31813
rect 24765 31804 24777 31807
rect 23624 31776 24777 31804
rect 23624 31764 23630 31776
rect 24765 31773 24777 31776
rect 24811 31773 24823 31807
rect 24765 31767 24823 31773
rect 11992 31708 12572 31736
rect 17218 31696 17224 31748
rect 17276 31736 17282 31748
rect 18966 31736 18972 31748
rect 17276 31708 18972 31736
rect 17276 31696 17282 31708
rect 18966 31696 18972 31708
rect 19024 31736 19030 31748
rect 19794 31736 19800 31748
rect 19024 31708 19800 31736
rect 19024 31696 19030 31708
rect 19794 31696 19800 31708
rect 19852 31696 19858 31748
rect 21729 31739 21787 31745
rect 21729 31705 21741 31739
rect 21775 31705 21787 31739
rect 21729 31699 21787 31705
rect 2498 31628 2504 31680
rect 2556 31668 2562 31680
rect 2774 31668 2780 31680
rect 2556 31640 2780 31668
rect 2556 31628 2562 31640
rect 2774 31628 2780 31640
rect 2832 31668 2838 31680
rect 2961 31671 3019 31677
rect 2961 31668 2973 31671
rect 2832 31640 2973 31668
rect 2832 31628 2838 31640
rect 2961 31637 2973 31640
rect 3007 31668 3019 31671
rect 3510 31668 3516 31680
rect 3007 31640 3516 31668
rect 3007 31637 3019 31640
rect 2961 31631 3019 31637
rect 3510 31628 3516 31640
rect 3568 31628 3574 31680
rect 14826 31628 14832 31680
rect 14884 31668 14890 31680
rect 15473 31671 15531 31677
rect 15473 31668 15485 31671
rect 14884 31640 15485 31668
rect 14884 31628 14890 31640
rect 15473 31637 15485 31640
rect 15519 31668 15531 31671
rect 20346 31668 20352 31680
rect 15519 31640 20352 31668
rect 15519 31637 15531 31640
rect 15473 31631 15531 31637
rect 20346 31628 20352 31640
rect 20404 31628 20410 31680
rect 21744 31668 21772 31699
rect 21818 31696 21824 31748
rect 21876 31736 21882 31748
rect 23937 31739 23995 31745
rect 23937 31736 23949 31739
rect 21876 31708 23949 31736
rect 21876 31696 21882 31708
rect 23937 31705 23949 31708
rect 23983 31705 23995 31739
rect 23937 31699 23995 31705
rect 23842 31668 23848 31680
rect 21744 31640 23848 31668
rect 23842 31628 23848 31640
rect 23900 31628 23906 31680
rect 25424 31668 25452 31835
rect 25682 31832 25688 31884
rect 25740 31881 25746 31884
rect 25740 31875 25789 31881
rect 25740 31841 25743 31875
rect 25777 31841 25789 31875
rect 25740 31835 25789 31841
rect 25961 31875 26019 31881
rect 25961 31841 25973 31875
rect 26007 31872 26019 31875
rect 26326 31872 26332 31884
rect 26007 31844 26332 31872
rect 26007 31841 26019 31844
rect 25961 31835 26019 31841
rect 25740 31832 25746 31835
rect 26326 31832 26332 31844
rect 26384 31832 26390 31884
rect 26988 31881 27016 31912
rect 26973 31875 27031 31881
rect 26973 31841 26985 31875
rect 27019 31841 27031 31875
rect 27157 31875 27215 31881
rect 27157 31872 27169 31875
rect 26973 31835 27031 31841
rect 27080 31844 27169 31872
rect 25501 31807 25559 31813
rect 25501 31773 25513 31807
rect 25547 31773 25559 31807
rect 25501 31767 25559 31773
rect 25516 31736 25544 31767
rect 26142 31764 26148 31816
rect 26200 31804 26206 31816
rect 26513 31807 26571 31813
rect 26513 31804 26525 31807
rect 26200 31776 26525 31804
rect 26200 31764 26206 31776
rect 26513 31773 26525 31776
rect 26559 31773 26571 31807
rect 26513 31767 26571 31773
rect 25682 31736 25688 31748
rect 25516 31708 25688 31736
rect 25682 31696 25688 31708
rect 25740 31696 25746 31748
rect 27080 31668 27108 31844
rect 27157 31841 27169 31844
rect 27203 31841 27215 31875
rect 27522 31872 27528 31884
rect 27483 31844 27528 31872
rect 27157 31835 27215 31841
rect 27522 31832 27528 31844
rect 27580 31832 27586 31884
rect 27709 31875 27767 31881
rect 27709 31841 27721 31875
rect 27755 31841 27767 31875
rect 28166 31872 28172 31884
rect 28127 31844 28172 31872
rect 27709 31835 27767 31841
rect 27724 31804 27752 31835
rect 28166 31832 28172 31844
rect 28224 31832 28230 31884
rect 28261 31875 28319 31881
rect 28261 31841 28273 31875
rect 28307 31872 28319 31875
rect 28810 31872 28816 31884
rect 28307 31844 28816 31872
rect 28307 31841 28319 31844
rect 28261 31835 28319 31841
rect 28810 31832 28816 31844
rect 28868 31832 28874 31884
rect 29564 31881 29592 31980
rect 33778 31968 33784 31980
rect 33836 31968 33842 32020
rect 36262 31968 36268 32020
rect 36320 32008 36326 32020
rect 36357 32011 36415 32017
rect 36357 32008 36369 32011
rect 36320 31980 36369 32008
rect 36320 31968 36326 31980
rect 36357 31977 36369 31980
rect 36403 31977 36415 32011
rect 36357 31971 36415 31977
rect 30834 31940 30840 31952
rect 30795 31912 30840 31940
rect 30834 31900 30840 31912
rect 30892 31900 30898 31952
rect 38470 31940 38476 31952
rect 38396 31912 38476 31940
rect 29549 31875 29607 31881
rect 29549 31841 29561 31875
rect 29595 31841 29607 31875
rect 30006 31872 30012 31884
rect 29967 31844 30012 31872
rect 29549 31835 29607 31841
rect 30006 31832 30012 31844
rect 30064 31832 30070 31884
rect 30098 31832 30104 31884
rect 30156 31872 30162 31884
rect 30469 31875 30527 31881
rect 30469 31872 30481 31875
rect 30156 31844 30481 31872
rect 30156 31832 30162 31844
rect 30469 31841 30481 31844
rect 30515 31841 30527 31875
rect 30469 31835 30527 31841
rect 30653 31875 30711 31881
rect 30653 31841 30665 31875
rect 30699 31841 30711 31875
rect 30653 31835 30711 31841
rect 30745 31875 30803 31881
rect 30745 31841 30757 31875
rect 30791 31872 30803 31875
rect 30926 31872 30932 31884
rect 30791 31844 30932 31872
rect 30791 31841 30803 31844
rect 30745 31835 30803 31841
rect 27890 31804 27896 31816
rect 27724 31776 27896 31804
rect 27890 31764 27896 31776
rect 27948 31804 27954 31816
rect 28442 31804 28448 31816
rect 27948 31776 28448 31804
rect 27948 31764 27954 31776
rect 28442 31764 28448 31776
rect 28500 31764 28506 31816
rect 28626 31764 28632 31816
rect 28684 31804 28690 31816
rect 28902 31804 28908 31816
rect 28684 31776 28908 31804
rect 28684 31764 28690 31776
rect 28902 31764 28908 31776
rect 28960 31764 28966 31816
rect 29641 31807 29699 31813
rect 29641 31773 29653 31807
rect 29687 31804 29699 31807
rect 30190 31804 30196 31816
rect 29687 31776 30196 31804
rect 29687 31773 29699 31776
rect 29641 31767 29699 31773
rect 30190 31764 30196 31776
rect 30248 31764 30254 31816
rect 30668 31804 30696 31835
rect 30926 31832 30932 31844
rect 30984 31832 30990 31884
rect 35526 31872 35532 31884
rect 32232 31844 32628 31872
rect 31018 31804 31024 31816
rect 30668 31776 31024 31804
rect 31018 31764 31024 31776
rect 31076 31764 31082 31816
rect 31205 31807 31263 31813
rect 31205 31773 31217 31807
rect 31251 31804 31263 31807
rect 31754 31804 31760 31816
rect 31251 31776 31760 31804
rect 31251 31773 31263 31776
rect 31205 31767 31263 31773
rect 31754 31764 31760 31776
rect 31812 31764 31818 31816
rect 32232 31813 32260 31844
rect 32217 31807 32275 31813
rect 32217 31804 32229 31807
rect 32127 31776 32229 31804
rect 32217 31773 32229 31776
rect 32263 31773 32275 31807
rect 32490 31804 32496 31816
rect 32451 31776 32496 31804
rect 32217 31767 32275 31773
rect 27246 31668 27252 31680
rect 25424 31640 27252 31668
rect 27246 31628 27252 31640
rect 27304 31628 27310 31680
rect 27706 31628 27712 31680
rect 27764 31668 27770 31680
rect 28445 31671 28503 31677
rect 28445 31668 28457 31671
rect 27764 31640 28457 31668
rect 27764 31628 27770 31640
rect 28445 31637 28457 31640
rect 28491 31637 28503 31671
rect 32232 31668 32260 31767
rect 32490 31764 32496 31776
rect 32548 31764 32554 31816
rect 32600 31804 32628 31844
rect 34716 31844 35532 31872
rect 34716 31816 34744 31844
rect 35526 31832 35532 31844
rect 35584 31832 35590 31884
rect 38010 31872 38016 31884
rect 37971 31844 38016 31872
rect 38010 31832 38016 31844
rect 38068 31832 38074 31884
rect 38286 31832 38292 31884
rect 38344 31872 38350 31884
rect 38396 31881 38424 31912
rect 38470 31900 38476 31912
rect 38528 31900 38534 31952
rect 38381 31875 38439 31881
rect 38381 31872 38393 31875
rect 38344 31844 38393 31872
rect 38344 31832 38350 31844
rect 38381 31841 38393 31844
rect 38427 31841 38439 31875
rect 38746 31872 38752 31884
rect 38707 31844 38752 31872
rect 38381 31835 38439 31841
rect 38746 31832 38752 31844
rect 38804 31832 38810 31884
rect 32600 31776 33180 31804
rect 33152 31736 33180 31776
rect 34698 31764 34704 31816
rect 34756 31764 34762 31816
rect 34977 31807 35035 31813
rect 34977 31773 34989 31807
rect 35023 31804 35035 31807
rect 35250 31804 35256 31816
rect 35023 31776 35057 31804
rect 35211 31776 35256 31804
rect 35023 31773 35035 31776
rect 34977 31767 35035 31773
rect 34992 31736 35020 31767
rect 35250 31764 35256 31776
rect 35308 31764 35314 31816
rect 38470 31764 38476 31816
rect 38528 31804 38534 31816
rect 38657 31807 38715 31813
rect 38657 31804 38669 31807
rect 38528 31776 38669 31804
rect 38528 31764 38534 31776
rect 38657 31773 38669 31776
rect 38703 31773 38715 31807
rect 38657 31767 38715 31773
rect 33152 31708 35020 31736
rect 32674 31668 32680 31680
rect 32232 31640 32680 31668
rect 28445 31631 28503 31637
rect 32674 31628 32680 31640
rect 32732 31628 32738 31680
rect 34992 31668 35020 31708
rect 35434 31668 35440 31680
rect 34992 31640 35440 31668
rect 35434 31628 35440 31640
rect 35492 31628 35498 31680
rect 1104 31578 39836 31600
rect 1104 31526 4246 31578
rect 4298 31526 4310 31578
rect 4362 31526 4374 31578
rect 4426 31526 4438 31578
rect 4490 31526 34966 31578
rect 35018 31526 35030 31578
rect 35082 31526 35094 31578
rect 35146 31526 35158 31578
rect 35210 31526 39836 31578
rect 1104 31504 39836 31526
rect 1670 31464 1676 31476
rect 1631 31436 1676 31464
rect 1670 31424 1676 31436
rect 1728 31424 1734 31476
rect 4798 31424 4804 31476
rect 4856 31464 4862 31476
rect 5626 31464 5632 31476
rect 4856 31436 5632 31464
rect 4856 31424 4862 31436
rect 5626 31424 5632 31436
rect 5684 31464 5690 31476
rect 6730 31464 6736 31476
rect 5684 31436 6736 31464
rect 5684 31424 5690 31436
rect 6730 31424 6736 31436
rect 6788 31424 6794 31476
rect 13078 31424 13084 31476
rect 13136 31464 13142 31476
rect 14093 31467 14151 31473
rect 14093 31464 14105 31467
rect 13136 31436 14105 31464
rect 13136 31424 13142 31436
rect 14093 31433 14105 31436
rect 14139 31433 14151 31467
rect 14093 31427 14151 31433
rect 14369 31467 14427 31473
rect 14369 31433 14381 31467
rect 14415 31464 14427 31467
rect 14550 31464 14556 31476
rect 14415 31436 14556 31464
rect 14415 31433 14427 31436
rect 14369 31427 14427 31433
rect 2866 31328 2872 31340
rect 2827 31300 2872 31328
rect 2866 31288 2872 31300
rect 2924 31288 2930 31340
rect 6748 31328 6776 31424
rect 12250 31356 12256 31408
rect 12308 31396 12314 31408
rect 12308 31368 13492 31396
rect 12308 31356 12314 31368
rect 7469 31331 7527 31337
rect 7469 31328 7481 31331
rect 6748 31300 7481 31328
rect 7469 31297 7481 31300
rect 7515 31297 7527 31331
rect 10321 31331 10379 31337
rect 7469 31291 7527 31297
rect 9876 31300 10272 31328
rect 1578 31260 1584 31272
rect 1539 31232 1584 31260
rect 1578 31220 1584 31232
rect 1636 31220 1642 31272
rect 2498 31260 2504 31272
rect 2459 31232 2504 31260
rect 2498 31220 2504 31232
rect 2556 31220 2562 31272
rect 2685 31263 2743 31269
rect 2685 31229 2697 31263
rect 2731 31260 2743 31263
rect 2774 31260 2780 31272
rect 2731 31232 2780 31260
rect 2731 31229 2743 31232
rect 2685 31223 2743 31229
rect 2774 31220 2780 31232
rect 2832 31260 2838 31272
rect 3050 31260 3056 31272
rect 2832 31232 3056 31260
rect 2832 31220 2838 31232
rect 3050 31220 3056 31232
rect 3108 31220 3114 31272
rect 3237 31263 3295 31269
rect 3237 31229 3249 31263
rect 3283 31229 3295 31263
rect 3237 31223 3295 31229
rect 3252 31192 3280 31223
rect 3326 31220 3332 31272
rect 3384 31260 3390 31272
rect 3697 31263 3755 31269
rect 3697 31260 3709 31263
rect 3384 31232 3709 31260
rect 3384 31220 3390 31232
rect 3697 31229 3709 31232
rect 3743 31260 3755 31263
rect 4062 31260 4068 31272
rect 3743 31232 4068 31260
rect 3743 31229 3755 31232
rect 3697 31223 3755 31229
rect 4062 31220 4068 31232
rect 4120 31260 4126 31272
rect 4341 31263 4399 31269
rect 4341 31260 4353 31263
rect 4120 31232 4353 31260
rect 4120 31220 4126 31232
rect 4341 31229 4353 31232
rect 4387 31229 4399 31263
rect 4982 31260 4988 31272
rect 4943 31232 4988 31260
rect 4341 31223 4399 31229
rect 4982 31220 4988 31232
rect 5040 31220 5046 31272
rect 5350 31260 5356 31272
rect 5311 31232 5356 31260
rect 5350 31220 5356 31232
rect 5408 31220 5414 31272
rect 5997 31263 6055 31269
rect 5997 31229 6009 31263
rect 6043 31260 6055 31263
rect 6822 31260 6828 31272
rect 6043 31232 6828 31260
rect 6043 31229 6055 31232
rect 5997 31223 6055 31229
rect 6822 31220 6828 31232
rect 6880 31220 6886 31272
rect 7742 31260 7748 31272
rect 7703 31232 7748 31260
rect 7742 31220 7748 31232
rect 7800 31220 7806 31272
rect 9876 31269 9904 31300
rect 9861 31263 9919 31269
rect 9861 31229 9873 31263
rect 9907 31229 9919 31263
rect 9861 31223 9919 31229
rect 10137 31263 10195 31269
rect 10137 31229 10149 31263
rect 10183 31229 10195 31263
rect 10244 31260 10272 31300
rect 10321 31297 10333 31331
rect 10367 31328 10379 31331
rect 11514 31328 11520 31340
rect 10367 31300 11520 31328
rect 10367 31297 10379 31300
rect 10321 31291 10379 31297
rect 11514 31288 11520 31300
rect 11572 31288 11578 31340
rect 12434 31288 12440 31340
rect 12492 31328 12498 31340
rect 13464 31337 13492 31368
rect 12989 31331 13047 31337
rect 12989 31328 13001 31331
rect 12492 31300 13001 31328
rect 12492 31288 12498 31300
rect 12989 31297 13001 31300
rect 13035 31297 13047 31331
rect 12989 31291 13047 31297
rect 13449 31331 13507 31337
rect 13449 31297 13461 31331
rect 13495 31328 13507 31331
rect 13814 31328 13820 31340
rect 13495 31300 13820 31328
rect 13495 31297 13507 31300
rect 13449 31291 13507 31297
rect 13814 31288 13820 31300
rect 13872 31328 13878 31340
rect 14384 31328 14412 31427
rect 14550 31424 14556 31436
rect 14608 31424 14614 31476
rect 15378 31424 15384 31476
rect 15436 31464 15442 31476
rect 17129 31467 17187 31473
rect 17129 31464 17141 31467
rect 15436 31436 17141 31464
rect 15436 31424 15442 31436
rect 17129 31433 17141 31436
rect 17175 31433 17187 31467
rect 17129 31427 17187 31433
rect 19886 31424 19892 31476
rect 19944 31464 19950 31476
rect 20622 31464 20628 31476
rect 19944 31436 20628 31464
rect 19944 31424 19950 31436
rect 20622 31424 20628 31436
rect 20680 31424 20686 31476
rect 35161 31467 35219 31473
rect 23952 31436 31984 31464
rect 22370 31356 22376 31408
rect 22428 31396 22434 31408
rect 23952 31405 23980 31436
rect 22833 31399 22891 31405
rect 22833 31396 22845 31399
rect 22428 31368 22845 31396
rect 22428 31356 22434 31368
rect 22833 31365 22845 31368
rect 22879 31365 22891 31399
rect 22833 31359 22891 31365
rect 23937 31399 23995 31405
rect 23937 31365 23949 31399
rect 23983 31365 23995 31399
rect 23937 31359 23995 31365
rect 25317 31399 25375 31405
rect 25317 31365 25329 31399
rect 25363 31365 25375 31399
rect 25317 31359 25375 31365
rect 13872 31300 14412 31328
rect 13872 31288 13878 31300
rect 15194 31288 15200 31340
rect 15252 31328 15258 31340
rect 15289 31331 15347 31337
rect 15289 31328 15301 31331
rect 15252 31300 15301 31328
rect 15252 31288 15258 31300
rect 15289 31297 15301 31300
rect 15335 31297 15347 31331
rect 15289 31291 15347 31297
rect 19429 31331 19487 31337
rect 19429 31297 19441 31331
rect 19475 31328 19487 31331
rect 21634 31328 21640 31340
rect 19475 31300 21640 31328
rect 19475 31297 19487 31300
rect 19429 31291 19487 31297
rect 21634 31288 21640 31300
rect 21692 31288 21698 31340
rect 21726 31288 21732 31340
rect 21784 31328 21790 31340
rect 22189 31331 22247 31337
rect 22189 31328 22201 31331
rect 21784 31300 22201 31328
rect 21784 31288 21790 31300
rect 22189 31297 22201 31300
rect 22235 31328 22247 31331
rect 23290 31328 23296 31340
rect 22235 31300 23296 31328
rect 22235 31297 22247 31300
rect 22189 31291 22247 31297
rect 23290 31288 23296 31300
rect 23348 31288 23354 31340
rect 24673 31331 24731 31337
rect 24673 31297 24685 31331
rect 24719 31328 24731 31331
rect 25332 31328 25360 31359
rect 26326 31356 26332 31408
rect 26384 31396 26390 31408
rect 26384 31368 28396 31396
rect 26384 31356 26390 31368
rect 24719 31300 25360 31328
rect 24719 31297 24731 31300
rect 24673 31291 24731 31297
rect 10686 31260 10692 31272
rect 10244 31232 10692 31260
rect 10137 31223 10195 31229
rect 4798 31192 4804 31204
rect 3252 31164 4804 31192
rect 4798 31152 4804 31164
rect 4856 31152 4862 31204
rect 9125 31195 9183 31201
rect 9125 31161 9137 31195
rect 9171 31192 9183 31195
rect 9214 31192 9220 31204
rect 9171 31164 9220 31192
rect 9171 31161 9183 31164
rect 9125 31155 9183 31161
rect 9214 31152 9220 31164
rect 9272 31152 9278 31204
rect 10152 31192 10180 31223
rect 10686 31220 10692 31232
rect 10744 31260 10750 31272
rect 10781 31263 10839 31269
rect 10781 31260 10793 31263
rect 10744 31232 10793 31260
rect 10744 31220 10750 31232
rect 10781 31229 10793 31232
rect 10827 31229 10839 31263
rect 10781 31223 10839 31229
rect 11146 31220 11152 31272
rect 11204 31260 11210 31272
rect 11241 31263 11299 31269
rect 11241 31260 11253 31263
rect 11204 31232 11253 31260
rect 11204 31220 11210 31232
rect 11241 31229 11253 31232
rect 11287 31229 11299 31263
rect 11241 31223 11299 31229
rect 11609 31263 11667 31269
rect 11609 31229 11621 31263
rect 11655 31229 11667 31263
rect 11609 31223 11667 31229
rect 11514 31192 11520 31204
rect 10152 31164 11520 31192
rect 11514 31152 11520 31164
rect 11572 31192 11578 31204
rect 11624 31192 11652 31223
rect 11698 31220 11704 31272
rect 11756 31260 11762 31272
rect 13265 31263 13323 31269
rect 13265 31260 13277 31263
rect 11756 31232 13277 31260
rect 11756 31220 11762 31232
rect 13265 31229 13277 31232
rect 13311 31229 13323 31263
rect 14182 31260 14188 31272
rect 14143 31232 14188 31260
rect 13265 31223 13323 31229
rect 11572 31164 11652 31192
rect 12437 31195 12495 31201
rect 11572 31152 11578 31164
rect 12437 31161 12449 31195
rect 12483 31192 12495 31195
rect 12710 31192 12716 31204
rect 12483 31164 12716 31192
rect 12483 31161 12495 31164
rect 12437 31155 12495 31161
rect 12710 31152 12716 31164
rect 12768 31152 12774 31204
rect 13280 31192 13308 31223
rect 14182 31220 14188 31232
rect 14240 31220 14246 31272
rect 15013 31263 15071 31269
rect 15013 31229 15025 31263
rect 15059 31260 15071 31263
rect 15378 31260 15384 31272
rect 15059 31232 15384 31260
rect 15059 31229 15071 31232
rect 15013 31223 15071 31229
rect 13998 31192 14004 31204
rect 13280 31164 14004 31192
rect 13998 31152 14004 31164
rect 14056 31152 14062 31204
rect 14093 31195 14151 31201
rect 14093 31161 14105 31195
rect 14139 31192 14151 31195
rect 15028 31192 15056 31223
rect 15378 31220 15384 31232
rect 15436 31220 15442 31272
rect 17310 31260 17316 31272
rect 17271 31232 17316 31260
rect 17310 31220 17316 31232
rect 17368 31220 17374 31272
rect 18874 31220 18880 31272
rect 18932 31260 18938 31272
rect 19334 31260 19340 31272
rect 18932 31232 19340 31260
rect 18932 31220 18938 31232
rect 19334 31220 19340 31232
rect 19392 31260 19398 31272
rect 19794 31260 19800 31272
rect 19392 31232 19437 31260
rect 19707 31232 19800 31260
rect 19392 31220 19398 31232
rect 19794 31220 19800 31232
rect 19852 31220 19858 31272
rect 19886 31220 19892 31272
rect 19944 31260 19950 31272
rect 19981 31263 20039 31269
rect 19981 31260 19993 31263
rect 19944 31232 19993 31260
rect 19944 31220 19950 31232
rect 19981 31229 19993 31232
rect 20027 31229 20039 31263
rect 20346 31260 20352 31272
rect 20307 31232 20352 31260
rect 19981 31223 20039 31229
rect 20346 31220 20352 31232
rect 20404 31220 20410 31272
rect 21082 31260 21088 31272
rect 21043 31232 21088 31260
rect 21082 31220 21088 31232
rect 21140 31220 21146 31272
rect 22557 31263 22615 31269
rect 22557 31229 22569 31263
rect 22603 31229 22615 31263
rect 22557 31223 22615 31229
rect 22925 31263 22983 31269
rect 22925 31229 22937 31263
rect 22971 31260 22983 31263
rect 23566 31260 23572 31272
rect 22971 31232 23572 31260
rect 22971 31229 22983 31232
rect 22925 31223 22983 31229
rect 14139 31164 15056 31192
rect 19812 31192 19840 31220
rect 20162 31192 20168 31204
rect 19812 31164 20168 31192
rect 14139 31161 14151 31164
rect 14093 31155 14151 31161
rect 20162 31152 20168 31164
rect 20220 31152 20226 31204
rect 22572 31192 22600 31223
rect 23566 31220 23572 31232
rect 23624 31220 23630 31272
rect 23661 31263 23719 31269
rect 23661 31229 23673 31263
rect 23707 31229 23719 31263
rect 23661 31223 23719 31229
rect 23106 31192 23112 31204
rect 22572 31164 23112 31192
rect 23106 31152 23112 31164
rect 23164 31152 23170 31204
rect 4433 31127 4491 31133
rect 4433 31093 4445 31127
rect 4479 31124 4491 31127
rect 4890 31124 4896 31136
rect 4479 31096 4896 31124
rect 4479 31093 4491 31096
rect 4433 31087 4491 31093
rect 4890 31084 4896 31096
rect 4948 31084 4954 31136
rect 5442 31084 5448 31136
rect 5500 31124 5506 31136
rect 6181 31127 6239 31133
rect 6181 31124 6193 31127
rect 5500 31096 6193 31124
rect 5500 31084 5506 31096
rect 6181 31093 6193 31096
rect 6227 31093 6239 31127
rect 6914 31124 6920 31136
rect 6875 31096 6920 31124
rect 6181 31087 6239 31093
rect 6914 31084 6920 31096
rect 6972 31084 6978 31136
rect 11882 31124 11888 31136
rect 11795 31096 11888 31124
rect 11882 31084 11888 31096
rect 11940 31124 11946 31136
rect 14366 31124 14372 31136
rect 11940 31096 14372 31124
rect 11940 31084 11946 31096
rect 14366 31084 14372 31096
rect 14424 31084 14430 31136
rect 16390 31124 16396 31136
rect 16351 31096 16396 31124
rect 16390 31084 16396 31096
rect 16448 31084 16454 31136
rect 22002 31084 22008 31136
rect 22060 31124 22066 31136
rect 22462 31124 22468 31136
rect 22060 31096 22468 31124
rect 22060 31084 22066 31096
rect 22462 31084 22468 31096
rect 22520 31084 22526 31136
rect 23566 31084 23572 31136
rect 23624 31124 23630 31136
rect 23676 31124 23704 31223
rect 23750 31220 23756 31272
rect 23808 31260 23814 31272
rect 24213 31263 24271 31269
rect 24213 31260 24225 31263
rect 23808 31232 24225 31260
rect 23808 31220 23814 31232
rect 24213 31229 24225 31232
rect 24259 31229 24271 31263
rect 24213 31223 24271 31229
rect 25130 31220 25136 31272
rect 25188 31260 25194 31272
rect 25225 31263 25283 31269
rect 25225 31260 25237 31263
rect 25188 31232 25237 31260
rect 25188 31220 25194 31232
rect 25225 31229 25237 31232
rect 25271 31229 25283 31263
rect 25774 31260 25780 31272
rect 25735 31232 25780 31260
rect 25225 31223 25283 31229
rect 25774 31220 25780 31232
rect 25832 31220 25838 31272
rect 26510 31260 26516 31272
rect 26471 31232 26516 31260
rect 26510 31220 26516 31232
rect 26568 31220 26574 31272
rect 26694 31260 26700 31272
rect 26655 31232 26700 31260
rect 26694 31220 26700 31232
rect 26752 31220 26758 31272
rect 27154 31260 27160 31272
rect 27067 31232 27160 31260
rect 27154 31220 27160 31232
rect 27212 31220 27218 31272
rect 27246 31220 27252 31272
rect 27304 31260 27310 31272
rect 28368 31269 28396 31368
rect 29730 31328 29736 31340
rect 29691 31300 29736 31328
rect 29730 31288 29736 31300
rect 29788 31288 29794 31340
rect 31754 31288 31760 31340
rect 31812 31328 31818 31340
rect 31812 31300 31857 31328
rect 31812 31288 31818 31300
rect 31956 31269 31984 31436
rect 35161 31433 35173 31467
rect 35207 31464 35219 31467
rect 35802 31464 35808 31476
rect 35207 31436 35808 31464
rect 35207 31433 35219 31436
rect 35161 31427 35219 31433
rect 32214 31356 32220 31408
rect 32272 31396 32278 31408
rect 32401 31399 32459 31405
rect 32401 31396 32413 31399
rect 32272 31368 32413 31396
rect 32272 31356 32278 31368
rect 32401 31365 32413 31368
rect 32447 31365 32459 31399
rect 32401 31359 32459 31365
rect 34514 31328 34520 31340
rect 33796 31300 34520 31328
rect 28353 31263 28411 31269
rect 27304 31232 27349 31260
rect 27304 31220 27310 31232
rect 28353 31229 28365 31263
rect 28399 31229 28411 31263
rect 28353 31223 28411 31229
rect 29457 31263 29515 31269
rect 29457 31229 29469 31263
rect 29503 31260 29515 31263
rect 31941 31263 31999 31269
rect 29503 31232 31892 31260
rect 29503 31229 29515 31232
rect 29457 31223 29515 31229
rect 25682 31152 25688 31204
rect 25740 31192 25746 31204
rect 27172 31192 27200 31220
rect 31864 31192 31892 31232
rect 31941 31229 31953 31263
rect 31987 31229 31999 31263
rect 31941 31223 31999 31229
rect 32030 31220 32036 31272
rect 32088 31260 32094 31272
rect 32401 31263 32459 31269
rect 32401 31260 32413 31263
rect 32088 31232 32413 31260
rect 32088 31220 32094 31232
rect 32401 31229 32413 31232
rect 32447 31229 32459 31263
rect 33410 31260 33416 31272
rect 33371 31232 33416 31260
rect 32401 31223 32459 31229
rect 33410 31220 33416 31232
rect 33468 31220 33474 31272
rect 33796 31269 33824 31300
rect 34514 31288 34520 31300
rect 34572 31288 34578 31340
rect 35176 31328 35204 31427
rect 35802 31424 35808 31436
rect 35860 31424 35866 31476
rect 34808 31300 35204 31328
rect 33781 31263 33839 31269
rect 33781 31229 33793 31263
rect 33827 31229 33839 31263
rect 33781 31223 33839 31229
rect 34149 31263 34207 31269
rect 34149 31229 34161 31263
rect 34195 31260 34207 31263
rect 34808 31260 34836 31300
rect 35710 31288 35716 31340
rect 35768 31328 35774 31340
rect 36725 31331 36783 31337
rect 36725 31328 36737 31331
rect 35768 31300 36737 31328
rect 35768 31288 35774 31300
rect 36725 31297 36737 31300
rect 36771 31297 36783 31331
rect 36725 31291 36783 31297
rect 34195 31232 34836 31260
rect 34977 31263 35035 31269
rect 34195 31229 34207 31232
rect 34149 31223 34207 31229
rect 34977 31229 34989 31263
rect 35023 31260 35035 31263
rect 35158 31260 35164 31272
rect 35023 31232 35164 31260
rect 35023 31229 35035 31232
rect 34977 31223 35035 31229
rect 35158 31220 35164 31232
rect 35216 31220 35222 31272
rect 35986 31260 35992 31272
rect 35947 31232 35992 31260
rect 35986 31220 35992 31232
rect 36044 31220 36050 31272
rect 36446 31260 36452 31272
rect 36359 31232 36452 31260
rect 36446 31220 36452 31232
rect 36504 31260 36510 31272
rect 36630 31260 36636 31272
rect 36504 31232 36636 31260
rect 36504 31220 36510 31232
rect 36630 31220 36636 31232
rect 36688 31220 36694 31272
rect 36814 31260 36820 31272
rect 36775 31232 36820 31260
rect 36814 31220 36820 31232
rect 36872 31220 36878 31272
rect 37461 31263 37519 31269
rect 37461 31229 37473 31263
rect 37507 31229 37519 31263
rect 37734 31260 37740 31272
rect 37695 31232 37740 31260
rect 37461 31223 37519 31229
rect 32674 31192 32680 31204
rect 25740 31164 27200 31192
rect 27632 31164 29500 31192
rect 31864 31164 32680 31192
rect 25740 31152 25746 31164
rect 27632 31124 27660 31164
rect 29472 31136 29500 31164
rect 32674 31152 32680 31164
rect 32732 31152 32738 31204
rect 34333 31195 34391 31201
rect 34333 31161 34345 31195
rect 34379 31192 34391 31195
rect 35434 31192 35440 31204
rect 34379 31164 35440 31192
rect 34379 31161 34391 31164
rect 34333 31155 34391 31161
rect 35434 31152 35440 31164
rect 35492 31152 35498 31204
rect 35526 31152 35532 31204
rect 35584 31192 35590 31204
rect 37476 31192 37504 31223
rect 37734 31220 37740 31232
rect 37792 31220 37798 31272
rect 35584 31164 37504 31192
rect 35584 31152 35590 31164
rect 23624 31096 27660 31124
rect 27709 31127 27767 31133
rect 23624 31084 23630 31096
rect 27709 31093 27721 31127
rect 27755 31124 27767 31127
rect 27982 31124 27988 31136
rect 27755 31096 27988 31124
rect 27755 31093 27767 31096
rect 27709 31087 27767 31093
rect 27982 31084 27988 31096
rect 28040 31084 28046 31136
rect 28442 31084 28448 31136
rect 28500 31124 28506 31136
rect 28537 31127 28595 31133
rect 28537 31124 28549 31127
rect 28500 31096 28549 31124
rect 28500 31084 28506 31096
rect 28537 31093 28549 31096
rect 28583 31093 28595 31127
rect 28537 31087 28595 31093
rect 29454 31084 29460 31136
rect 29512 31084 29518 31136
rect 30374 31084 30380 31136
rect 30432 31124 30438 31136
rect 30837 31127 30895 31133
rect 30837 31124 30849 31127
rect 30432 31096 30849 31124
rect 30432 31084 30438 31096
rect 30837 31093 30849 31096
rect 30883 31093 30895 31127
rect 30837 31087 30895 31093
rect 38102 31084 38108 31136
rect 38160 31124 38166 31136
rect 38562 31124 38568 31136
rect 38160 31096 38568 31124
rect 38160 31084 38166 31096
rect 38562 31084 38568 31096
rect 38620 31124 38626 31136
rect 38841 31127 38899 31133
rect 38841 31124 38853 31127
rect 38620 31096 38853 31124
rect 38620 31084 38626 31096
rect 38841 31093 38853 31096
rect 38887 31093 38899 31127
rect 38841 31087 38899 31093
rect 1104 31034 39836 31056
rect 1104 30982 19606 31034
rect 19658 30982 19670 31034
rect 19722 30982 19734 31034
rect 19786 30982 19798 31034
rect 19850 30982 39836 31034
rect 1104 30960 39836 30982
rect 4356 30892 6776 30920
rect 2130 30812 2136 30864
rect 2188 30852 2194 30864
rect 2501 30855 2559 30861
rect 2501 30852 2513 30855
rect 2188 30824 2513 30852
rect 2188 30812 2194 30824
rect 2501 30821 2513 30824
rect 2547 30821 2559 30855
rect 2501 30815 2559 30821
rect 3326 30784 3332 30796
rect 3287 30756 3332 30784
rect 3326 30744 3332 30756
rect 3384 30744 3390 30796
rect 3510 30784 3516 30796
rect 3471 30756 3516 30784
rect 3510 30744 3516 30756
rect 3568 30744 3574 30796
rect 4356 30793 4384 30892
rect 4341 30787 4399 30793
rect 4341 30753 4353 30787
rect 4387 30753 4399 30787
rect 4890 30784 4896 30796
rect 4851 30756 4896 30784
rect 4341 30747 4399 30753
rect 4890 30744 4896 30756
rect 4948 30744 4954 30796
rect 5169 30787 5227 30793
rect 5169 30753 5181 30787
rect 5215 30784 5227 30787
rect 5905 30787 5963 30793
rect 5905 30784 5917 30787
rect 5215 30756 5917 30784
rect 5215 30753 5227 30756
rect 5169 30747 5227 30753
rect 5905 30753 5917 30756
rect 5951 30753 5963 30787
rect 6748 30784 6776 30892
rect 6822 30880 6828 30932
rect 6880 30920 6886 30932
rect 7009 30923 7067 30929
rect 7009 30920 7021 30923
rect 6880 30892 7021 30920
rect 6880 30880 6886 30892
rect 7009 30889 7021 30892
rect 7055 30889 7067 30923
rect 7009 30883 7067 30889
rect 8754 30880 8760 30932
rect 8812 30920 8818 30932
rect 10413 30923 10471 30929
rect 10413 30920 10425 30923
rect 8812 30892 10425 30920
rect 8812 30880 8818 30892
rect 10413 30889 10425 30892
rect 10459 30920 10471 30923
rect 11698 30920 11704 30932
rect 10459 30892 11704 30920
rect 10459 30889 10471 30892
rect 10413 30883 10471 30889
rect 11698 30880 11704 30892
rect 11756 30880 11762 30932
rect 12345 30923 12403 30929
rect 12345 30889 12357 30923
rect 12391 30920 12403 30923
rect 12526 30920 12532 30932
rect 12391 30892 12532 30920
rect 12391 30889 12403 30892
rect 12345 30883 12403 30889
rect 12526 30880 12532 30892
rect 12584 30880 12590 30932
rect 20254 30920 20260 30932
rect 19352 30892 20260 30920
rect 8938 30852 8944 30864
rect 8220 30824 8944 30852
rect 7006 30784 7012 30796
rect 6748 30756 7012 30784
rect 5905 30747 5963 30753
rect 7006 30744 7012 30756
rect 7064 30744 7070 30796
rect 8220 30793 8248 30824
rect 8938 30812 8944 30824
rect 8996 30812 9002 30864
rect 9769 30855 9827 30861
rect 9769 30821 9781 30855
rect 9815 30852 9827 30855
rect 14826 30852 14832 30864
rect 9815 30824 10364 30852
rect 9815 30821 9827 30824
rect 9769 30815 9827 30821
rect 8205 30787 8263 30793
rect 8205 30753 8217 30787
rect 8251 30753 8263 30787
rect 8205 30747 8263 30753
rect 8294 30744 8300 30796
rect 8352 30784 8358 30796
rect 8665 30787 8723 30793
rect 8665 30784 8677 30787
rect 8352 30756 8677 30784
rect 8352 30744 8358 30756
rect 8665 30753 8677 30756
rect 8711 30753 8723 30787
rect 8665 30747 8723 30753
rect 9493 30787 9551 30793
rect 9493 30753 9505 30787
rect 9539 30753 9551 30787
rect 9493 30747 9551 30753
rect 3053 30719 3111 30725
rect 3053 30685 3065 30719
rect 3099 30716 3111 30719
rect 4706 30716 4712 30728
rect 3099 30688 4712 30716
rect 3099 30685 3111 30688
rect 3053 30679 3111 30685
rect 4706 30676 4712 30688
rect 4764 30676 4770 30728
rect 4985 30719 5043 30725
rect 4985 30685 4997 30719
rect 5031 30716 5043 30719
rect 5626 30716 5632 30728
rect 5031 30688 5488 30716
rect 5587 30688 5632 30716
rect 5031 30685 5043 30688
rect 4985 30679 5043 30685
rect 5460 30648 5488 30688
rect 5626 30676 5632 30688
rect 5684 30676 5690 30728
rect 8478 30716 8484 30728
rect 8439 30688 8484 30716
rect 8478 30676 8484 30688
rect 8536 30676 8542 30728
rect 9508 30716 9536 30747
rect 9674 30744 9680 30796
rect 9732 30784 9738 30796
rect 10336 30793 10364 30824
rect 11164 30824 12296 30852
rect 11164 30796 11192 30824
rect 10321 30787 10379 30793
rect 9732 30756 9777 30784
rect 9732 30744 9738 30756
rect 10321 30753 10333 30787
rect 10367 30753 10379 30787
rect 10321 30747 10379 30753
rect 10686 30744 10692 30796
rect 10744 30784 10750 30796
rect 10781 30787 10839 30793
rect 10781 30784 10793 30787
rect 10744 30756 10793 30784
rect 10744 30744 10750 30756
rect 10781 30753 10793 30756
rect 10827 30753 10839 30787
rect 11146 30784 11152 30796
rect 11107 30756 11152 30784
rect 10781 30747 10839 30753
rect 11146 30744 11152 30756
rect 11204 30744 11210 30796
rect 11514 30784 11520 30796
rect 11475 30756 11520 30784
rect 11514 30744 11520 30756
rect 11572 30744 11578 30796
rect 12268 30793 12296 30824
rect 13832 30824 14832 30852
rect 12253 30787 12311 30793
rect 12253 30753 12265 30787
rect 12299 30753 12311 30787
rect 12253 30747 12311 30753
rect 13541 30787 13599 30793
rect 13541 30753 13553 30787
rect 13587 30784 13599 30787
rect 13722 30784 13728 30796
rect 13587 30756 13728 30784
rect 13587 30753 13599 30756
rect 13541 30747 13599 30753
rect 13722 30744 13728 30756
rect 13780 30744 13786 30796
rect 13832 30793 13860 30824
rect 14826 30812 14832 30824
rect 14884 30812 14890 30864
rect 15286 30812 15292 30864
rect 15344 30812 15350 30864
rect 17862 30852 17868 30864
rect 17144 30824 17868 30852
rect 13817 30787 13875 30793
rect 13817 30753 13829 30787
rect 13863 30753 13875 30787
rect 13998 30784 14004 30796
rect 13959 30756 14004 30784
rect 13817 30747 13875 30753
rect 13998 30744 14004 30756
rect 14056 30744 14062 30796
rect 14737 30787 14795 30793
rect 14737 30753 14749 30787
rect 14783 30784 14795 30787
rect 15304 30784 15332 30812
rect 17144 30796 17172 30824
rect 17862 30812 17868 30824
rect 17920 30812 17926 30864
rect 16114 30784 16120 30796
rect 14783 30756 15976 30784
rect 16075 30756 16120 30784
rect 14783 30753 14795 30756
rect 14737 30747 14795 30753
rect 10962 30716 10968 30728
rect 9508 30688 10968 30716
rect 10962 30676 10968 30688
rect 11020 30676 11026 30728
rect 11532 30716 11560 30744
rect 12802 30716 12808 30728
rect 11532 30688 12808 30716
rect 12802 30676 12808 30688
rect 12860 30676 12866 30728
rect 15289 30719 15347 30725
rect 15289 30685 15301 30719
rect 15335 30716 15347 30719
rect 15378 30716 15384 30728
rect 15335 30688 15384 30716
rect 15335 30685 15347 30688
rect 15289 30679 15347 30685
rect 15378 30676 15384 30688
rect 15436 30676 15442 30728
rect 15841 30719 15899 30725
rect 15841 30685 15853 30719
rect 15887 30685 15899 30719
rect 15948 30716 15976 30756
rect 16114 30744 16120 30756
rect 16172 30744 16178 30796
rect 17037 30787 17095 30793
rect 17037 30753 17049 30787
rect 17083 30784 17095 30787
rect 17126 30784 17132 30796
rect 17083 30756 17132 30784
rect 17083 30753 17095 30756
rect 17037 30747 17095 30753
rect 17126 30744 17132 30756
rect 17184 30744 17190 30796
rect 17218 30744 17224 30796
rect 17276 30784 17282 30796
rect 17586 30784 17592 30796
rect 17276 30756 17321 30784
rect 17547 30756 17592 30784
rect 17276 30744 17282 30756
rect 17586 30744 17592 30756
rect 17644 30744 17650 30796
rect 17678 30744 17684 30796
rect 17736 30784 17742 30796
rect 17957 30787 18015 30793
rect 17957 30784 17969 30787
rect 17736 30756 17969 30784
rect 17736 30744 17742 30756
rect 17957 30753 17969 30756
rect 18003 30753 18015 30787
rect 17957 30747 18015 30753
rect 18693 30787 18751 30793
rect 18693 30753 18705 30787
rect 18739 30784 18751 30787
rect 18874 30784 18880 30796
rect 18739 30756 18880 30784
rect 18739 30753 18751 30756
rect 18693 30747 18751 30753
rect 18874 30744 18880 30756
rect 18932 30744 18938 30796
rect 19352 30793 19380 30892
rect 20254 30880 20260 30892
rect 20312 30920 20318 30932
rect 21726 30920 21732 30932
rect 20312 30892 21732 30920
rect 20312 30880 20318 30892
rect 21726 30880 21732 30892
rect 21784 30880 21790 30932
rect 23753 30923 23811 30929
rect 23753 30889 23765 30923
rect 23799 30920 23811 30923
rect 23799 30892 30880 30920
rect 23799 30889 23811 30892
rect 23753 30883 23811 30889
rect 26142 30852 26148 30864
rect 20088 30824 26148 30852
rect 20088 30793 20116 30824
rect 26142 30812 26148 30824
rect 26200 30812 26206 30864
rect 29638 30852 29644 30864
rect 29599 30824 29644 30852
rect 29638 30812 29644 30824
rect 29696 30812 29702 30864
rect 19337 30787 19395 30793
rect 19337 30753 19349 30787
rect 19383 30753 19395 30787
rect 19337 30747 19395 30753
rect 19705 30787 19763 30793
rect 19705 30753 19717 30787
rect 19751 30753 19763 30787
rect 19705 30747 19763 30753
rect 20073 30787 20131 30793
rect 20073 30753 20085 30787
rect 20119 30753 20131 30787
rect 21634 30784 21640 30796
rect 21595 30756 21640 30784
rect 20073 30747 20131 30753
rect 16301 30719 16359 30725
rect 16301 30716 16313 30719
rect 15948 30688 16313 30716
rect 15841 30679 15899 30685
rect 16301 30685 16313 30688
rect 16347 30716 16359 30719
rect 16390 30716 16396 30728
rect 16347 30688 16396 30716
rect 16347 30685 16359 30688
rect 16301 30679 16359 30685
rect 5534 30648 5540 30660
rect 5460 30620 5540 30648
rect 5534 30608 5540 30620
rect 5592 30608 5598 30660
rect 8754 30608 8760 30660
rect 8812 30648 8818 30660
rect 15102 30648 15108 30660
rect 8812 30620 15108 30648
rect 8812 30608 8818 30620
rect 15102 30608 15108 30620
rect 15160 30648 15166 30660
rect 15856 30648 15884 30679
rect 16390 30676 16396 30688
rect 16448 30676 16454 30728
rect 19720 30716 19748 30747
rect 21634 30744 21640 30756
rect 21692 30744 21698 30796
rect 22370 30784 22376 30796
rect 22331 30756 22376 30784
rect 22370 30744 22376 30756
rect 22428 30744 22434 30796
rect 23566 30744 23572 30796
rect 23624 30784 23630 30796
rect 23661 30787 23719 30793
rect 23661 30784 23673 30787
rect 23624 30756 23673 30784
rect 23624 30744 23630 30756
rect 23661 30753 23673 30756
rect 23707 30753 23719 30787
rect 24210 30784 24216 30796
rect 24171 30756 24216 30784
rect 23661 30747 23719 30753
rect 24210 30744 24216 30756
rect 24268 30744 24274 30796
rect 25222 30784 25228 30796
rect 25183 30756 25228 30784
rect 25222 30744 25228 30756
rect 25280 30744 25286 30796
rect 25406 30744 25412 30796
rect 25464 30784 25470 30796
rect 25774 30784 25780 30796
rect 25464 30756 25780 30784
rect 25464 30744 25470 30756
rect 25774 30744 25780 30756
rect 25832 30744 25838 30796
rect 26881 30787 26939 30793
rect 26881 30753 26893 30787
rect 26927 30784 26939 30787
rect 27062 30784 27068 30796
rect 26927 30756 27068 30784
rect 26927 30753 26939 30756
rect 26881 30747 26939 30753
rect 27062 30744 27068 30756
rect 27120 30744 27126 30796
rect 28626 30784 28632 30796
rect 27448 30756 28632 30784
rect 20346 30716 20352 30728
rect 19720 30688 20352 30716
rect 20346 30676 20352 30688
rect 20404 30676 20410 30728
rect 22278 30676 22284 30728
rect 22336 30716 22342 30728
rect 22465 30719 22523 30725
rect 22465 30716 22477 30719
rect 22336 30688 22477 30716
rect 22336 30676 22342 30688
rect 22465 30685 22477 30688
rect 22511 30685 22523 30719
rect 22465 30679 22523 30685
rect 24673 30719 24731 30725
rect 24673 30685 24685 30719
rect 24719 30685 24731 30719
rect 24673 30679 24731 30685
rect 26973 30719 27031 30725
rect 26973 30685 26985 30719
rect 27019 30716 27031 30719
rect 27448 30716 27476 30756
rect 28626 30744 28632 30756
rect 28684 30744 28690 30796
rect 30852 30793 30880 30892
rect 33410 30880 33416 30932
rect 33468 30920 33474 30932
rect 34057 30923 34115 30929
rect 34057 30920 34069 30923
rect 33468 30892 34069 30920
rect 33468 30880 33474 30892
rect 34057 30889 34069 30892
rect 34103 30889 34115 30923
rect 34057 30883 34115 30889
rect 35069 30923 35127 30929
rect 35069 30889 35081 30923
rect 35115 30920 35127 30923
rect 35250 30920 35256 30932
rect 35115 30892 35256 30920
rect 35115 30889 35127 30892
rect 35069 30883 35127 30889
rect 35250 30880 35256 30892
rect 35308 30880 35314 30932
rect 36814 30880 36820 30932
rect 36872 30920 36878 30932
rect 36909 30923 36967 30929
rect 36909 30920 36921 30923
rect 36872 30892 36921 30920
rect 36872 30880 36878 30892
rect 36909 30889 36921 30892
rect 36955 30889 36967 30923
rect 36909 30883 36967 30889
rect 37734 30880 37740 30932
rect 37792 30920 37798 30932
rect 37829 30923 37887 30929
rect 37829 30920 37841 30923
rect 37792 30892 37841 30920
rect 37792 30880 37798 30892
rect 37829 30889 37841 30892
rect 37875 30889 37887 30923
rect 37829 30883 37887 30889
rect 36262 30812 36268 30864
rect 36320 30852 36326 30864
rect 36320 30824 36860 30852
rect 36320 30812 36326 30824
rect 30377 30787 30435 30793
rect 30377 30753 30389 30787
rect 30423 30784 30435 30787
rect 30837 30787 30895 30793
rect 30423 30756 30788 30784
rect 30423 30753 30435 30756
rect 30377 30747 30435 30753
rect 27019 30688 27476 30716
rect 27525 30719 27583 30725
rect 27019 30685 27031 30688
rect 26973 30679 27031 30685
rect 27525 30685 27537 30719
rect 27571 30716 27583 30719
rect 27614 30716 27620 30728
rect 27571 30688 27620 30716
rect 27571 30685 27583 30688
rect 27525 30679 27583 30685
rect 15160 30620 15884 30648
rect 17037 30651 17095 30657
rect 15160 30608 15166 30620
rect 17037 30617 17049 30651
rect 17083 30648 17095 30651
rect 18230 30648 18236 30660
rect 17083 30620 18236 30648
rect 17083 30617 17095 30620
rect 17037 30611 17095 30617
rect 18230 30608 18236 30620
rect 18288 30608 18294 30660
rect 19978 30648 19984 30660
rect 19939 30620 19984 30648
rect 19978 30608 19984 30620
rect 20036 30608 20042 30660
rect 21913 30651 21971 30657
rect 21913 30617 21925 30651
rect 21959 30648 21971 30651
rect 22094 30648 22100 30660
rect 21959 30620 22100 30648
rect 21959 30617 21971 30620
rect 21913 30611 21971 30617
rect 22094 30608 22100 30620
rect 22152 30608 22158 30660
rect 24688 30648 24716 30679
rect 27614 30676 27620 30688
rect 27672 30676 27678 30728
rect 27985 30719 28043 30725
rect 27985 30685 27997 30719
rect 28031 30685 28043 30719
rect 27985 30679 28043 30685
rect 28261 30719 28319 30725
rect 28261 30685 28273 30719
rect 28307 30716 28319 30719
rect 29730 30716 29736 30728
rect 28307 30688 29736 30716
rect 28307 30685 28319 30688
rect 28261 30679 28319 30685
rect 25317 30651 25375 30657
rect 25317 30648 25329 30651
rect 24688 30620 25329 30648
rect 25317 30617 25329 30620
rect 25363 30617 25375 30651
rect 25317 30611 25375 30617
rect 27246 30608 27252 30660
rect 27304 30648 27310 30660
rect 28000 30648 28028 30679
rect 29730 30676 29736 30688
rect 29788 30676 29794 30728
rect 30558 30716 30564 30728
rect 30519 30688 30564 30716
rect 30558 30676 30564 30688
rect 30616 30676 30622 30728
rect 30760 30716 30788 30756
rect 30837 30753 30849 30787
rect 30883 30753 30895 30787
rect 30837 30747 30895 30753
rect 31389 30787 31447 30793
rect 31389 30753 31401 30787
rect 31435 30753 31447 30787
rect 31389 30747 31447 30753
rect 31573 30787 31631 30793
rect 31573 30753 31585 30787
rect 31619 30784 31631 30787
rect 32950 30784 32956 30796
rect 31619 30756 32812 30784
rect 32911 30756 32956 30784
rect 31619 30753 31631 30756
rect 31573 30747 31631 30753
rect 31110 30716 31116 30728
rect 30760 30688 31116 30716
rect 31110 30676 31116 30688
rect 31168 30676 31174 30728
rect 27304 30620 28028 30648
rect 27304 30608 27310 30620
rect 9306 30580 9312 30592
rect 9267 30552 9312 30580
rect 9306 30540 9312 30552
rect 9364 30540 9370 30592
rect 14645 30583 14703 30589
rect 14645 30549 14657 30583
rect 14691 30580 14703 30583
rect 15286 30580 15292 30592
rect 14691 30552 15292 30580
rect 14691 30549 14703 30552
rect 14645 30543 14703 30549
rect 15286 30540 15292 30552
rect 15344 30540 15350 30592
rect 28000 30580 28028 30620
rect 28994 30580 29000 30592
rect 28000 30552 29000 30580
rect 28994 30540 29000 30552
rect 29052 30580 29058 30592
rect 29178 30580 29184 30592
rect 29052 30552 29184 30580
rect 29052 30540 29058 30552
rect 29178 30540 29184 30552
rect 29236 30540 29242 30592
rect 30193 30583 30251 30589
rect 30193 30549 30205 30583
rect 30239 30580 30251 30583
rect 30742 30580 30748 30592
rect 30239 30552 30748 30580
rect 30239 30549 30251 30552
rect 30193 30543 30251 30549
rect 30742 30540 30748 30552
rect 30800 30540 30806 30592
rect 31404 30580 31432 30747
rect 32674 30716 32680 30728
rect 32635 30688 32680 30716
rect 32674 30676 32680 30688
rect 32732 30676 32738 30728
rect 32784 30716 32812 30756
rect 32950 30744 32956 30756
rect 33008 30744 33014 30796
rect 35161 30787 35219 30793
rect 35161 30753 35173 30787
rect 35207 30784 35219 30787
rect 35342 30784 35348 30796
rect 35207 30756 35348 30784
rect 35207 30753 35219 30756
rect 35161 30747 35219 30753
rect 35342 30744 35348 30756
rect 35400 30744 35406 30796
rect 35710 30784 35716 30796
rect 35671 30756 35716 30784
rect 35710 30744 35716 30756
rect 35768 30744 35774 30796
rect 36446 30744 36452 30796
rect 36504 30784 36510 30796
rect 36832 30793 36860 30824
rect 36633 30787 36691 30793
rect 36633 30784 36645 30787
rect 36504 30756 36645 30784
rect 36504 30744 36510 30756
rect 36633 30753 36645 30756
rect 36679 30753 36691 30787
rect 36633 30747 36691 30753
rect 36817 30787 36875 30793
rect 36817 30753 36829 30787
rect 36863 30753 36875 30787
rect 36817 30747 36875 30753
rect 36906 30744 36912 30796
rect 36964 30784 36970 30796
rect 37737 30787 37795 30793
rect 37737 30784 37749 30787
rect 36964 30756 37749 30784
rect 36964 30744 36970 30756
rect 37737 30753 37749 30756
rect 37783 30753 37795 30787
rect 38470 30784 38476 30796
rect 38431 30756 38476 30784
rect 37737 30747 37795 30753
rect 38470 30744 38476 30756
rect 38528 30744 38534 30796
rect 34790 30716 34796 30728
rect 32784 30688 34796 30716
rect 34790 30676 34796 30688
rect 34848 30676 34854 30728
rect 35805 30719 35863 30725
rect 35805 30685 35817 30719
rect 35851 30716 35863 30719
rect 36354 30716 36360 30728
rect 35851 30688 36360 30716
rect 35851 30685 35863 30688
rect 35805 30679 35863 30685
rect 36354 30676 36360 30688
rect 36412 30676 36418 30728
rect 37642 30676 37648 30728
rect 37700 30716 37706 30728
rect 37826 30716 37832 30728
rect 37700 30688 37832 30716
rect 37700 30676 37706 30688
rect 37826 30676 37832 30688
rect 37884 30716 37890 30728
rect 38565 30719 38623 30725
rect 38565 30716 38577 30719
rect 37884 30688 38577 30716
rect 37884 30676 37890 30688
rect 38565 30685 38577 30688
rect 38611 30685 38623 30719
rect 38565 30679 38623 30685
rect 32030 30580 32036 30592
rect 31404 30552 32036 30580
rect 32030 30540 32036 30552
rect 32088 30540 32094 30592
rect 1104 30490 39836 30512
rect 1104 30438 4246 30490
rect 4298 30438 4310 30490
rect 4362 30438 4374 30490
rect 4426 30438 4438 30490
rect 4490 30438 34966 30490
rect 35018 30438 35030 30490
rect 35082 30438 35094 30490
rect 35146 30438 35158 30490
rect 35210 30438 39836 30490
rect 1104 30416 39836 30438
rect 7101 30379 7159 30385
rect 3252 30348 3556 30376
rect 1762 30200 1768 30252
rect 1820 30240 1826 30252
rect 3252 30240 3280 30348
rect 1820 30212 3280 30240
rect 3528 30240 3556 30348
rect 7101 30345 7113 30379
rect 7147 30376 7159 30379
rect 7742 30376 7748 30388
rect 7147 30348 7748 30376
rect 7147 30345 7159 30348
rect 7101 30339 7159 30345
rect 7742 30336 7748 30348
rect 7800 30336 7806 30388
rect 8478 30376 8484 30388
rect 7944 30348 8484 30376
rect 4062 30268 4068 30320
rect 4120 30308 4126 30320
rect 4120 30280 4660 30308
rect 4120 30268 4126 30280
rect 4341 30243 4399 30249
rect 4341 30240 4353 30243
rect 3528 30212 4353 30240
rect 1820 30200 1826 30212
rect 4341 30209 4353 30212
rect 4387 30209 4399 30243
rect 4341 30203 4399 30209
rect 2774 30132 2780 30184
rect 2832 30172 2838 30184
rect 2958 30172 2964 30184
rect 2832 30144 2877 30172
rect 2919 30144 2964 30172
rect 2832 30132 2838 30144
rect 2958 30132 2964 30144
rect 3016 30132 3022 30184
rect 3234 30172 3240 30184
rect 3195 30144 3240 30172
rect 3234 30132 3240 30144
rect 3292 30132 3298 30184
rect 3418 30172 3424 30184
rect 3379 30144 3424 30172
rect 3418 30132 3424 30144
rect 3476 30132 3482 30184
rect 3510 30132 3516 30184
rect 3568 30172 3574 30184
rect 4632 30181 4660 30280
rect 5810 30268 5816 30320
rect 5868 30308 5874 30320
rect 7558 30308 7564 30320
rect 5868 30280 7564 30308
rect 5868 30268 5874 30280
rect 7558 30268 7564 30280
rect 7616 30268 7622 30320
rect 7944 30240 7972 30348
rect 8478 30336 8484 30348
rect 8536 30336 8542 30388
rect 8938 30376 8944 30388
rect 8899 30348 8944 30376
rect 8938 30336 8944 30348
rect 8996 30336 9002 30388
rect 19518 30336 19524 30388
rect 19576 30376 19582 30388
rect 20254 30376 20260 30388
rect 19576 30348 20260 30376
rect 19576 30336 19582 30348
rect 20254 30336 20260 30348
rect 20312 30336 20318 30388
rect 23750 30376 23756 30388
rect 22572 30348 23756 30376
rect 11146 30308 11152 30320
rect 7024 30212 7972 30240
rect 8036 30280 11152 30308
rect 3605 30175 3663 30181
rect 3605 30172 3617 30175
rect 3568 30144 3617 30172
rect 3568 30132 3574 30144
rect 3605 30141 3617 30144
rect 3651 30141 3663 30175
rect 3605 30135 3663 30141
rect 4249 30175 4307 30181
rect 4249 30141 4261 30175
rect 4295 30141 4307 30175
rect 4249 30135 4307 30141
rect 4617 30175 4675 30181
rect 4617 30141 4629 30175
rect 4663 30141 4675 30175
rect 4982 30172 4988 30184
rect 4943 30144 4988 30172
rect 4617 30135 4675 30141
rect 1486 30064 1492 30116
rect 1544 30104 1550 30116
rect 2317 30107 2375 30113
rect 2317 30104 2329 30107
rect 1544 30076 2329 30104
rect 1544 30064 1550 30076
rect 2317 30073 2329 30076
rect 2363 30073 2375 30107
rect 2792 30104 2820 30132
rect 4264 30104 4292 30135
rect 4982 30132 4988 30144
rect 5040 30132 5046 30184
rect 5350 30132 5356 30184
rect 5408 30172 5414 30184
rect 7024 30181 7052 30212
rect 8036 30181 8064 30280
rect 11146 30268 11152 30280
rect 11204 30268 11210 30320
rect 17313 30311 17371 30317
rect 17313 30277 17325 30311
rect 17359 30308 17371 30311
rect 22572 30308 22600 30348
rect 23750 30336 23756 30348
rect 23808 30336 23814 30388
rect 25498 30336 25504 30388
rect 25556 30376 25562 30388
rect 28629 30379 28687 30385
rect 28629 30376 28641 30379
rect 25556 30348 28641 30376
rect 25556 30336 25562 30348
rect 28629 30345 28641 30348
rect 28675 30345 28687 30379
rect 28629 30339 28687 30345
rect 32953 30379 33011 30385
rect 32953 30345 32965 30379
rect 32999 30376 33011 30379
rect 33042 30376 33048 30388
rect 32999 30348 33048 30376
rect 32999 30345 33011 30348
rect 32953 30339 33011 30345
rect 33042 30336 33048 30348
rect 33100 30336 33106 30388
rect 34241 30379 34299 30385
rect 34241 30345 34253 30379
rect 34287 30376 34299 30379
rect 34514 30376 34520 30388
rect 34287 30348 34520 30376
rect 34287 30345 34299 30348
rect 34241 30339 34299 30345
rect 34514 30336 34520 30348
rect 34572 30336 34578 30388
rect 17359 30280 22600 30308
rect 22649 30311 22707 30317
rect 17359 30277 17371 30280
rect 17313 30271 17371 30277
rect 22649 30277 22661 30311
rect 22695 30308 22707 30311
rect 24210 30308 24216 30320
rect 22695 30280 24216 30308
rect 22695 30277 22707 30280
rect 22649 30271 22707 30277
rect 24210 30268 24216 30280
rect 24268 30268 24274 30320
rect 31938 30308 31944 30320
rect 27356 30280 30788 30308
rect 31899 30280 31944 30308
rect 10502 30240 10508 30252
rect 8956 30212 9260 30240
rect 10463 30212 10508 30240
rect 5537 30175 5595 30181
rect 5537 30172 5549 30175
rect 5408 30144 5549 30172
rect 5408 30132 5414 30144
rect 5537 30141 5549 30144
rect 5583 30141 5595 30175
rect 5537 30135 5595 30141
rect 6365 30175 6423 30181
rect 6365 30141 6377 30175
rect 6411 30141 6423 30175
rect 6365 30135 6423 30141
rect 7009 30175 7067 30181
rect 7009 30141 7021 30175
rect 7055 30141 7067 30175
rect 7009 30135 7067 30141
rect 7929 30175 7987 30181
rect 7929 30141 7941 30175
rect 7975 30141 7987 30175
rect 7929 30135 7987 30141
rect 8021 30175 8079 30181
rect 8021 30141 8033 30175
rect 8067 30141 8079 30175
rect 8021 30135 8079 30141
rect 8389 30175 8447 30181
rect 8389 30141 8401 30175
rect 8435 30172 8447 30175
rect 8956 30172 8984 30212
rect 9232 30184 9260 30212
rect 10502 30200 10508 30212
rect 10560 30200 10566 30252
rect 12710 30240 12716 30252
rect 12671 30212 12716 30240
rect 12710 30200 12716 30212
rect 12768 30200 12774 30252
rect 14366 30200 14372 30252
rect 14424 30240 14430 30252
rect 14645 30243 14703 30249
rect 14645 30240 14657 30243
rect 14424 30212 14657 30240
rect 14424 30200 14430 30212
rect 14645 30209 14657 30212
rect 14691 30209 14703 30243
rect 14645 30203 14703 30209
rect 15381 30243 15439 30249
rect 15381 30209 15393 30243
rect 15427 30240 15439 30243
rect 16114 30240 16120 30252
rect 15427 30212 16120 30240
rect 15427 30209 15439 30212
rect 15381 30203 15439 30209
rect 16114 30200 16120 30212
rect 16172 30200 16178 30252
rect 16577 30243 16635 30249
rect 16577 30209 16589 30243
rect 16623 30240 16635 30243
rect 18506 30240 18512 30252
rect 16623 30212 18512 30240
rect 16623 30209 16635 30212
rect 16577 30203 16635 30209
rect 18506 30200 18512 30212
rect 18564 30200 18570 30252
rect 19613 30243 19671 30249
rect 19613 30209 19625 30243
rect 19659 30240 19671 30243
rect 24486 30240 24492 30252
rect 19659 30212 23704 30240
rect 24447 30212 24492 30240
rect 19659 30209 19671 30212
rect 19613 30203 19671 30209
rect 8435 30144 8984 30172
rect 8435 30141 8447 30144
rect 8389 30135 8447 30141
rect 2792 30076 4292 30104
rect 2317 30067 2375 30073
rect 4706 30064 4712 30116
rect 4764 30104 4770 30116
rect 6380 30104 6408 30135
rect 7834 30104 7840 30116
rect 4764 30076 6316 30104
rect 6380 30076 7840 30104
rect 4764 30064 4770 30076
rect 3878 29996 3884 30048
rect 3936 30036 3942 30048
rect 6181 30039 6239 30045
rect 6181 30036 6193 30039
rect 3936 30008 6193 30036
rect 3936 29996 3942 30008
rect 6181 30005 6193 30008
rect 6227 30005 6239 30039
rect 6288 30036 6316 30076
rect 7834 30064 7840 30076
rect 7892 30064 7898 30116
rect 7944 30104 7972 30135
rect 9030 30132 9036 30184
rect 9088 30172 9094 30184
rect 9214 30172 9220 30184
rect 9088 30144 9133 30172
rect 9175 30144 9220 30172
rect 9088 30132 9094 30144
rect 9214 30132 9220 30144
rect 9272 30132 9278 30184
rect 9861 30175 9919 30181
rect 9861 30141 9873 30175
rect 9907 30141 9919 30175
rect 9861 30135 9919 30141
rect 9048 30104 9076 30132
rect 7944 30076 9076 30104
rect 9876 30104 9904 30135
rect 10870 30132 10876 30184
rect 10928 30172 10934 30184
rect 10965 30175 11023 30181
rect 10965 30172 10977 30175
rect 10928 30144 10977 30172
rect 10928 30132 10934 30144
rect 10965 30141 10977 30144
rect 11011 30141 11023 30175
rect 10965 30135 11023 30141
rect 11054 30132 11060 30184
rect 11112 30172 11118 30184
rect 11149 30175 11207 30181
rect 11149 30172 11161 30175
rect 11112 30144 11161 30172
rect 11112 30132 11118 30144
rect 11149 30141 11161 30144
rect 11195 30141 11207 30175
rect 11149 30135 11207 30141
rect 11333 30175 11391 30181
rect 11333 30141 11345 30175
rect 11379 30172 11391 30175
rect 11790 30172 11796 30184
rect 11379 30144 11796 30172
rect 11379 30141 11391 30144
rect 11333 30135 11391 30141
rect 11348 30104 11376 30135
rect 11790 30132 11796 30144
rect 11848 30132 11854 30184
rect 12437 30175 12495 30181
rect 12437 30141 12449 30175
rect 12483 30172 12495 30175
rect 13078 30172 13084 30184
rect 12483 30144 13084 30172
rect 12483 30141 12495 30144
rect 12437 30135 12495 30141
rect 13078 30132 13084 30144
rect 13136 30132 13142 30184
rect 14458 30132 14464 30184
rect 14516 30172 14522 30184
rect 16945 30175 17003 30181
rect 14516 30144 15056 30172
rect 14516 30132 14522 30144
rect 14826 30104 14832 30116
rect 9876 30076 11376 30104
rect 14787 30076 14832 30104
rect 14826 30064 14832 30076
rect 14884 30064 14890 30116
rect 15028 30113 15056 30144
rect 16945 30141 16957 30175
rect 16991 30172 17003 30175
rect 17313 30175 17371 30181
rect 16991 30144 17172 30172
rect 16991 30141 17003 30144
rect 16945 30135 17003 30141
rect 15013 30107 15071 30113
rect 15013 30073 15025 30107
rect 15059 30073 15071 30107
rect 15013 30067 15071 30073
rect 7650 30036 7656 30048
rect 6288 30008 7656 30036
rect 6181 29999 6239 30005
rect 7650 29996 7656 30008
rect 7708 29996 7714 30048
rect 14001 30039 14059 30045
rect 14001 30005 14013 30039
rect 14047 30036 14059 30039
rect 14182 30036 14188 30048
rect 14047 30008 14188 30036
rect 14047 30005 14059 30008
rect 14001 29999 14059 30005
rect 14182 29996 14188 30008
rect 14240 30036 14246 30048
rect 14921 30039 14979 30045
rect 14921 30036 14933 30039
rect 14240 30008 14933 30036
rect 14240 29996 14246 30008
rect 14921 30005 14933 30008
rect 14967 30036 14979 30039
rect 15194 30036 15200 30048
rect 14967 30008 15200 30036
rect 14967 30005 14979 30008
rect 14921 29999 14979 30005
rect 15194 29996 15200 30008
rect 15252 30036 15258 30048
rect 15562 30036 15568 30048
rect 15252 30008 15568 30036
rect 15252 29996 15258 30008
rect 15562 29996 15568 30008
rect 15620 29996 15626 30048
rect 17144 30036 17172 30144
rect 17313 30141 17325 30175
rect 17359 30172 17371 30175
rect 19150 30172 19156 30184
rect 17359 30144 19156 30172
rect 17359 30141 17371 30144
rect 17313 30135 17371 30141
rect 19150 30132 19156 30144
rect 19208 30132 19214 30184
rect 19518 30172 19524 30184
rect 19479 30144 19524 30172
rect 19518 30132 19524 30144
rect 19576 30132 19582 30184
rect 19794 30172 19800 30184
rect 19755 30144 19800 30172
rect 19794 30132 19800 30144
rect 19852 30132 19858 30184
rect 19886 30132 19892 30184
rect 19944 30172 19950 30184
rect 20165 30175 20223 30181
rect 20165 30172 20177 30175
rect 19944 30144 20177 30172
rect 19944 30132 19950 30144
rect 20165 30141 20177 30144
rect 20211 30141 20223 30175
rect 20530 30172 20536 30184
rect 20491 30144 20536 30172
rect 20165 30135 20223 30141
rect 20530 30132 20536 30144
rect 20588 30132 20594 30184
rect 21082 30132 21088 30184
rect 21140 30172 21146 30184
rect 21269 30175 21327 30181
rect 21269 30172 21281 30175
rect 21140 30144 21281 30172
rect 21140 30132 21146 30144
rect 21269 30141 21281 30144
rect 21315 30172 21327 30175
rect 21634 30172 21640 30184
rect 21315 30144 21640 30172
rect 21315 30141 21327 30144
rect 21269 30135 21327 30141
rect 21634 30132 21640 30144
rect 21692 30132 21698 30184
rect 21729 30175 21787 30181
rect 21729 30141 21741 30175
rect 21775 30141 21787 30175
rect 21729 30135 21787 30141
rect 19334 30064 19340 30116
rect 19392 30104 19398 30116
rect 21744 30104 21772 30135
rect 22094 30132 22100 30184
rect 22152 30172 22158 30184
rect 23676 30181 23704 30212
rect 24486 30200 24492 30212
rect 24544 30200 24550 30252
rect 25314 30200 25320 30252
rect 25372 30240 25378 30252
rect 25498 30240 25504 30252
rect 25372 30212 25504 30240
rect 25372 30200 25378 30212
rect 25498 30200 25504 30212
rect 25556 30240 25562 30252
rect 25869 30243 25927 30249
rect 25869 30240 25881 30243
rect 25556 30212 25881 30240
rect 25556 30200 25562 30212
rect 25869 30209 25881 30212
rect 25915 30209 25927 30243
rect 26326 30240 26332 30252
rect 26287 30212 26332 30240
rect 25869 30203 25927 30209
rect 26326 30200 26332 30212
rect 26384 30200 26390 30252
rect 22557 30175 22615 30181
rect 22152 30144 22197 30172
rect 22152 30132 22158 30144
rect 22557 30141 22569 30175
rect 22603 30141 22615 30175
rect 22557 30135 22615 30141
rect 23661 30175 23719 30181
rect 23661 30141 23673 30175
rect 23707 30141 23719 30175
rect 23661 30135 23719 30141
rect 19392 30076 21772 30104
rect 19392 30064 19398 30076
rect 21818 30064 21824 30116
rect 21876 30104 21882 30116
rect 22572 30104 22600 30135
rect 23842 30132 23848 30184
rect 23900 30172 23906 30184
rect 24213 30175 24271 30181
rect 24213 30172 24225 30175
rect 23900 30144 24225 30172
rect 23900 30132 23906 30144
rect 24213 30141 24225 30144
rect 24259 30141 24271 30175
rect 24213 30135 24271 30141
rect 24302 30132 24308 30184
rect 24360 30172 24366 30184
rect 25409 30175 25467 30181
rect 25409 30172 25421 30175
rect 24360 30144 25421 30172
rect 24360 30132 24366 30144
rect 25409 30141 25421 30144
rect 25455 30141 25467 30175
rect 26050 30172 26056 30184
rect 26011 30144 26056 30172
rect 25409 30135 25467 30141
rect 26050 30132 26056 30144
rect 26108 30132 26114 30184
rect 26418 30172 26424 30184
rect 26379 30144 26424 30172
rect 26418 30132 26424 30144
rect 26476 30132 26482 30184
rect 27356 30181 27384 30280
rect 30760 30252 30788 30280
rect 31938 30268 31944 30280
rect 31996 30268 32002 30320
rect 32030 30268 32036 30320
rect 32088 30308 32094 30320
rect 34146 30308 34152 30320
rect 32088 30280 34152 30308
rect 32088 30268 32094 30280
rect 34146 30268 34152 30280
rect 34204 30268 34210 30320
rect 35805 30311 35863 30317
rect 35805 30277 35817 30311
rect 35851 30308 35863 30311
rect 36906 30308 36912 30320
rect 35851 30280 36912 30308
rect 35851 30277 35863 30280
rect 35805 30271 35863 30277
rect 36906 30268 36912 30280
rect 36964 30268 36970 30320
rect 30282 30240 30288 30252
rect 27632 30212 30288 30240
rect 27632 30181 27660 30212
rect 30282 30200 30288 30212
rect 30340 30200 30346 30252
rect 30558 30240 30564 30252
rect 30519 30212 30564 30240
rect 30558 30200 30564 30212
rect 30616 30200 30622 30252
rect 30742 30200 30748 30252
rect 30800 30240 30806 30252
rect 32048 30240 32076 30268
rect 37458 30240 37464 30252
rect 30800 30212 31800 30240
rect 30800 30200 30806 30212
rect 27341 30175 27399 30181
rect 27341 30141 27353 30175
rect 27387 30141 27399 30175
rect 27341 30135 27399 30141
rect 27617 30175 27675 30181
rect 27617 30141 27629 30175
rect 27663 30141 27675 30175
rect 27617 30135 27675 30141
rect 28445 30175 28503 30181
rect 28445 30141 28457 30175
rect 28491 30172 28503 30175
rect 28534 30172 28540 30184
rect 28491 30144 28540 30172
rect 28491 30141 28503 30144
rect 28445 30135 28503 30141
rect 28534 30132 28540 30144
rect 28592 30132 28598 30184
rect 29822 30172 29828 30184
rect 29735 30144 29828 30172
rect 29822 30132 29828 30144
rect 29880 30172 29886 30184
rect 30098 30172 30104 30184
rect 29880 30144 30104 30172
rect 29880 30132 29886 30144
rect 30098 30132 30104 30144
rect 30156 30132 30162 30184
rect 31202 30172 31208 30184
rect 31163 30144 31208 30172
rect 31202 30132 31208 30144
rect 31260 30132 31266 30184
rect 31389 30175 31447 30181
rect 31389 30141 31401 30175
rect 31435 30141 31447 30175
rect 31389 30135 31447 30141
rect 21876 30076 22600 30104
rect 27433 30107 27491 30113
rect 21876 30064 21882 30076
rect 27433 30073 27445 30107
rect 27479 30104 27491 30107
rect 27479 30076 28488 30104
rect 27479 30073 27491 30076
rect 27433 30067 27491 30073
rect 28460 30048 28488 30076
rect 29638 30064 29644 30116
rect 29696 30104 29702 30116
rect 30193 30107 30251 30113
rect 30193 30104 30205 30107
rect 29696 30076 30205 30104
rect 29696 30064 29702 30076
rect 30193 30073 30205 30076
rect 30239 30073 30251 30107
rect 30193 30067 30251 30073
rect 30466 30064 30472 30116
rect 30524 30104 30530 30116
rect 31404 30104 31432 30135
rect 30524 30076 31432 30104
rect 31772 30104 31800 30212
rect 31956 30212 32076 30240
rect 37419 30212 37464 30240
rect 31956 30181 31984 30212
rect 37458 30200 37464 30212
rect 37516 30200 37522 30252
rect 39114 30240 39120 30252
rect 39075 30212 39120 30240
rect 39114 30200 39120 30212
rect 39172 30200 39178 30252
rect 31941 30175 31999 30181
rect 31941 30141 31953 30175
rect 31987 30141 31999 30175
rect 31941 30135 31999 30141
rect 32769 30175 32827 30181
rect 32769 30141 32781 30175
rect 32815 30141 32827 30175
rect 32769 30135 32827 30141
rect 33045 30175 33103 30181
rect 33045 30141 33057 30175
rect 33091 30172 33103 30175
rect 33318 30172 33324 30184
rect 33091 30144 33324 30172
rect 33091 30141 33103 30144
rect 33045 30135 33103 30141
rect 32784 30104 32812 30135
rect 33318 30132 33324 30144
rect 33376 30132 33382 30184
rect 33502 30172 33508 30184
rect 33463 30144 33508 30172
rect 33502 30132 33508 30144
rect 33560 30132 33566 30184
rect 34057 30175 34115 30181
rect 34057 30141 34069 30175
rect 34103 30172 34115 30175
rect 34422 30172 34428 30184
rect 34103 30144 34428 30172
rect 34103 30141 34115 30144
rect 34057 30135 34115 30141
rect 34422 30132 34428 30144
rect 34480 30132 34486 30184
rect 34514 30132 34520 30184
rect 34572 30172 34578 30184
rect 34885 30175 34943 30181
rect 34885 30172 34897 30175
rect 34572 30144 34897 30172
rect 34572 30132 34578 30144
rect 34885 30141 34897 30144
rect 34931 30141 34943 30175
rect 34885 30135 34943 30141
rect 35437 30175 35495 30181
rect 35437 30141 35449 30175
rect 35483 30172 35495 30175
rect 35618 30172 35624 30184
rect 35483 30144 35624 30172
rect 35483 30141 35495 30144
rect 35437 30135 35495 30141
rect 35618 30132 35624 30144
rect 35676 30132 35682 30184
rect 35802 30172 35808 30184
rect 35763 30144 35808 30172
rect 35802 30132 35808 30144
rect 35860 30132 35866 30184
rect 36633 30175 36691 30181
rect 36633 30141 36645 30175
rect 36679 30172 36691 30175
rect 36906 30172 36912 30184
rect 36679 30144 36912 30172
rect 36679 30141 36691 30144
rect 36633 30135 36691 30141
rect 36906 30132 36912 30144
rect 36964 30132 36970 30184
rect 37366 30132 37372 30184
rect 37424 30172 37430 30184
rect 37737 30175 37795 30181
rect 37737 30172 37749 30175
rect 37424 30144 37749 30172
rect 37424 30132 37430 30144
rect 37737 30141 37749 30144
rect 37783 30141 37795 30175
rect 37737 30135 37795 30141
rect 36446 30104 36452 30116
rect 31772 30076 32812 30104
rect 36407 30076 36452 30104
rect 30524 30064 30530 30076
rect 36446 30064 36452 30076
rect 36504 30064 36510 30116
rect 37001 30107 37059 30113
rect 37001 30073 37013 30107
rect 37047 30073 37059 30107
rect 37001 30067 37059 30073
rect 23753 30039 23811 30045
rect 23753 30036 23765 30039
rect 17144 30008 23765 30036
rect 23753 30005 23765 30008
rect 23799 30005 23811 30039
rect 27154 30036 27160 30048
rect 27115 30008 27160 30036
rect 23753 29999 23811 30005
rect 27154 29996 27160 30008
rect 27212 29996 27218 30048
rect 27706 30036 27712 30048
rect 27667 30008 27712 30036
rect 27706 29996 27712 30008
rect 27764 29996 27770 30048
rect 28442 29996 28448 30048
rect 28500 29996 28506 30048
rect 30006 30036 30012 30048
rect 29967 30008 30012 30036
rect 30006 29996 30012 30008
rect 30064 29996 30070 30048
rect 30098 29996 30104 30048
rect 30156 30036 30162 30048
rect 32585 30039 32643 30045
rect 30156 30008 30201 30036
rect 30156 29996 30162 30008
rect 32585 30005 32597 30039
rect 32631 30036 32643 30039
rect 32674 30036 32680 30048
rect 32631 30008 32680 30036
rect 32631 30005 32643 30008
rect 32585 29999 32643 30005
rect 32674 29996 32680 30008
rect 32732 30036 32738 30048
rect 33042 30036 33048 30048
rect 32732 30008 33048 30036
rect 32732 29996 32738 30008
rect 33042 29996 33048 30008
rect 33100 29996 33106 30048
rect 37016 30036 37044 30067
rect 38562 30036 38568 30048
rect 37016 30008 38568 30036
rect 38562 29996 38568 30008
rect 38620 29996 38626 30048
rect 1104 29946 39836 29968
rect 1104 29894 19606 29946
rect 19658 29894 19670 29946
rect 19722 29894 19734 29946
rect 19786 29894 19798 29946
rect 19850 29894 39836 29946
rect 1104 29872 39836 29894
rect 2774 29792 2780 29844
rect 2832 29832 2838 29844
rect 2832 29804 2877 29832
rect 2832 29792 2838 29804
rect 3510 29792 3516 29844
rect 3568 29832 3574 29844
rect 5442 29832 5448 29844
rect 3568 29804 5448 29832
rect 3568 29792 3574 29804
rect 5442 29792 5448 29804
rect 5500 29792 5506 29844
rect 5534 29792 5540 29844
rect 5592 29832 5598 29844
rect 5997 29835 6055 29841
rect 5997 29832 6009 29835
rect 5592 29804 6009 29832
rect 5592 29792 5598 29804
rect 5997 29801 6009 29804
rect 6043 29801 6055 29835
rect 5997 29795 6055 29801
rect 9769 29835 9827 29841
rect 9769 29801 9781 29835
rect 9815 29801 9827 29835
rect 9769 29795 9827 29801
rect 9876 29804 23980 29832
rect 3142 29724 3148 29776
rect 3200 29764 3206 29776
rect 3418 29764 3424 29776
rect 3200 29736 3424 29764
rect 3200 29724 3206 29736
rect 3418 29724 3424 29736
rect 3476 29764 3482 29776
rect 5350 29764 5356 29776
rect 3476 29736 5356 29764
rect 3476 29724 3482 29736
rect 5350 29724 5356 29736
rect 5408 29724 5414 29776
rect 6914 29764 6920 29776
rect 5828 29736 6920 29764
rect 1394 29696 1400 29708
rect 1355 29668 1400 29696
rect 1394 29656 1400 29668
rect 1452 29656 1458 29708
rect 2866 29656 2872 29708
rect 2924 29696 2930 29708
rect 5828 29705 5856 29736
rect 6914 29724 6920 29736
rect 6972 29724 6978 29776
rect 8113 29767 8171 29773
rect 8113 29733 8125 29767
rect 8159 29764 8171 29767
rect 8294 29764 8300 29776
rect 8159 29736 8300 29764
rect 8159 29733 8171 29736
rect 8113 29727 8171 29733
rect 8294 29724 8300 29736
rect 8352 29724 8358 29776
rect 9784 29764 9812 29795
rect 8956 29736 9812 29764
rect 8956 29708 8984 29736
rect 4065 29699 4123 29705
rect 4065 29696 4077 29699
rect 2924 29668 4077 29696
rect 2924 29656 2930 29668
rect 4065 29665 4077 29668
rect 4111 29696 4123 29699
rect 4801 29699 4859 29705
rect 4801 29696 4813 29699
rect 4111 29668 4813 29696
rect 4111 29665 4123 29668
rect 4065 29659 4123 29665
rect 4801 29665 4813 29668
rect 4847 29665 4859 29699
rect 4801 29659 4859 29665
rect 5537 29699 5595 29705
rect 5537 29665 5549 29699
rect 5583 29665 5595 29699
rect 5537 29659 5595 29665
rect 5813 29699 5871 29705
rect 5813 29665 5825 29699
rect 5859 29665 5871 29699
rect 5994 29696 6000 29708
rect 5955 29668 6000 29696
rect 5813 29659 5871 29665
rect 1670 29628 1676 29640
rect 1631 29600 1676 29628
rect 1670 29588 1676 29600
rect 1728 29588 1734 29640
rect 5442 29588 5448 29640
rect 5500 29628 5506 29640
rect 5552 29628 5580 29659
rect 5994 29656 6000 29668
rect 6052 29656 6058 29708
rect 6733 29699 6791 29705
rect 6733 29665 6745 29699
rect 6779 29696 6791 29699
rect 7006 29696 7012 29708
rect 6779 29668 7012 29696
rect 6779 29665 6791 29668
rect 6733 29659 6791 29665
rect 7006 29656 7012 29668
rect 7064 29656 7070 29708
rect 7377 29699 7435 29705
rect 7377 29665 7389 29699
rect 7423 29665 7435 29699
rect 7377 29659 7435 29665
rect 8665 29699 8723 29705
rect 8665 29665 8677 29699
rect 8711 29696 8723 29699
rect 8754 29696 8760 29708
rect 8711 29668 8760 29696
rect 8711 29665 8723 29668
rect 8665 29659 8723 29665
rect 6825 29631 6883 29637
rect 6825 29628 6837 29631
rect 5500 29600 6837 29628
rect 5500 29588 5506 29600
rect 6825 29597 6837 29600
rect 6871 29597 6883 29631
rect 6825 29591 6883 29597
rect 4798 29520 4804 29572
rect 4856 29560 4862 29572
rect 7392 29560 7420 29659
rect 8754 29656 8760 29668
rect 8812 29656 8818 29708
rect 8938 29696 8944 29708
rect 8851 29668 8944 29696
rect 8938 29656 8944 29668
rect 8996 29656 9002 29708
rect 9398 29656 9404 29708
rect 9456 29696 9462 29708
rect 9876 29696 9904 29804
rect 11422 29764 11428 29776
rect 9968 29736 11428 29764
rect 9968 29705 9996 29736
rect 11422 29724 11428 29736
rect 11480 29724 11486 29776
rect 12618 29764 12624 29776
rect 12268 29736 12624 29764
rect 9456 29668 9904 29696
rect 9953 29699 10011 29705
rect 9456 29656 9462 29668
rect 9953 29665 9965 29699
rect 9999 29665 10011 29699
rect 9953 29659 10011 29665
rect 10226 29656 10232 29708
rect 10284 29696 10290 29708
rect 10502 29696 10508 29708
rect 10284 29668 10508 29696
rect 10284 29656 10290 29668
rect 10502 29656 10508 29668
rect 10560 29656 10566 29708
rect 10686 29696 10692 29708
rect 10647 29668 10692 29696
rect 10686 29656 10692 29668
rect 10744 29656 10750 29708
rect 11238 29696 11244 29708
rect 11199 29668 11244 29696
rect 11238 29656 11244 29668
rect 11296 29656 11302 29708
rect 11790 29696 11796 29708
rect 11751 29668 11796 29696
rect 11790 29656 11796 29668
rect 11848 29656 11854 29708
rect 12268 29705 12296 29736
rect 12618 29724 12624 29736
rect 12676 29764 12682 29776
rect 19978 29764 19984 29776
rect 12676 29736 14504 29764
rect 12676 29724 12682 29736
rect 12253 29699 12311 29705
rect 12253 29665 12265 29699
rect 12299 29665 12311 29699
rect 12253 29659 12311 29665
rect 12434 29656 12440 29708
rect 12492 29696 12498 29708
rect 12805 29699 12863 29705
rect 12805 29696 12817 29699
rect 12492 29668 12817 29696
rect 12492 29656 12498 29668
rect 12805 29665 12817 29668
rect 12851 29665 12863 29699
rect 12805 29659 12863 29665
rect 13449 29699 13507 29705
rect 13449 29665 13461 29699
rect 13495 29696 13507 29699
rect 13722 29696 13728 29708
rect 13495 29668 13728 29696
rect 13495 29665 13507 29668
rect 13449 29659 13507 29665
rect 13722 29656 13728 29668
rect 13780 29656 13786 29708
rect 14274 29696 14280 29708
rect 14235 29668 14280 29696
rect 14274 29656 14280 29668
rect 14332 29656 14338 29708
rect 14476 29705 14504 29736
rect 18892 29736 19984 29764
rect 14461 29699 14519 29705
rect 14461 29665 14473 29699
rect 14507 29665 14519 29699
rect 15286 29696 15292 29708
rect 15247 29668 15292 29696
rect 14461 29659 14519 29665
rect 15286 29656 15292 29668
rect 15344 29656 15350 29708
rect 15378 29656 15384 29708
rect 15436 29696 15442 29708
rect 15841 29699 15899 29705
rect 15841 29696 15853 29699
rect 15436 29668 15853 29696
rect 15436 29656 15442 29668
rect 15841 29665 15853 29668
rect 15887 29665 15899 29699
rect 15841 29659 15899 29665
rect 15930 29656 15936 29708
rect 15988 29696 15994 29708
rect 16669 29699 16727 29705
rect 16669 29696 16681 29699
rect 15988 29668 16681 29696
rect 15988 29656 15994 29668
rect 16669 29665 16681 29668
rect 16715 29665 16727 29699
rect 16669 29659 16727 29665
rect 17405 29699 17463 29705
rect 17405 29665 17417 29699
rect 17451 29696 17463 29699
rect 17586 29696 17592 29708
rect 17451 29668 17592 29696
rect 17451 29665 17463 29668
rect 17405 29659 17463 29665
rect 17586 29656 17592 29668
rect 17644 29656 17650 29708
rect 18230 29696 18236 29708
rect 18191 29668 18236 29696
rect 18230 29656 18236 29668
rect 18288 29656 18294 29708
rect 18892 29705 18920 29736
rect 19978 29724 19984 29736
rect 20036 29724 20042 29776
rect 20530 29764 20536 29776
rect 20180 29736 20536 29764
rect 18877 29699 18935 29705
rect 18877 29665 18889 29699
rect 18923 29665 18935 29699
rect 19058 29696 19064 29708
rect 19019 29668 19064 29696
rect 18877 29659 18935 29665
rect 19058 29656 19064 29668
rect 19116 29656 19122 29708
rect 19794 29656 19800 29708
rect 19852 29696 19858 29708
rect 19852 29668 19897 29696
rect 19852 29656 19858 29668
rect 9125 29631 9183 29637
rect 9125 29597 9137 29631
rect 9171 29628 9183 29631
rect 9214 29628 9220 29640
rect 9171 29600 9220 29628
rect 9171 29597 9183 29600
rect 9125 29591 9183 29597
rect 9214 29588 9220 29600
rect 9272 29588 9278 29640
rect 13538 29588 13544 29640
rect 13596 29628 13602 29640
rect 14553 29631 14611 29637
rect 14553 29628 14565 29631
rect 13596 29600 14565 29628
rect 13596 29588 13602 29600
rect 14553 29597 14565 29600
rect 14599 29597 14611 29631
rect 15654 29628 15660 29640
rect 15615 29600 15660 29628
rect 14553 29591 14611 29597
rect 15654 29588 15660 29600
rect 15712 29588 15718 29640
rect 17497 29631 17555 29637
rect 17497 29628 17509 29631
rect 15764 29600 17509 29628
rect 11330 29560 11336 29572
rect 4856 29532 7420 29560
rect 11291 29532 11336 29560
rect 4856 29520 4862 29532
rect 11330 29520 11336 29532
rect 11388 29520 11394 29572
rect 12894 29560 12900 29572
rect 12855 29532 12900 29560
rect 12894 29520 12900 29532
rect 12952 29520 12958 29572
rect 13630 29520 13636 29572
rect 13688 29560 13694 29572
rect 15764 29560 15792 29600
rect 17497 29597 17509 29600
rect 17543 29597 17555 29631
rect 19610 29628 19616 29640
rect 17497 29591 17555 29597
rect 18248 29600 19616 29628
rect 13688 29532 15792 29560
rect 16945 29563 17003 29569
rect 13688 29520 13694 29532
rect 16945 29529 16957 29563
rect 16991 29560 17003 29563
rect 18248 29560 18276 29600
rect 19610 29588 19616 29600
rect 19668 29588 19674 29640
rect 20180 29628 20208 29736
rect 20530 29724 20536 29736
rect 20588 29724 20594 29776
rect 21174 29724 21180 29776
rect 21232 29764 21238 29776
rect 21818 29764 21824 29776
rect 21232 29736 21824 29764
rect 21232 29724 21238 29736
rect 21818 29724 21824 29736
rect 21876 29724 21882 29776
rect 23952 29764 23980 29804
rect 24228 29804 29592 29832
rect 24228 29764 24256 29804
rect 23952 29736 24256 29764
rect 24486 29724 24492 29776
rect 24544 29764 24550 29776
rect 25314 29764 25320 29776
rect 24544 29736 25320 29764
rect 24544 29724 24550 29736
rect 25314 29724 25320 29736
rect 25372 29724 25378 29776
rect 27249 29767 27307 29773
rect 27249 29764 27261 29767
rect 26528 29736 27261 29764
rect 20714 29656 20720 29708
rect 20772 29696 20778 29708
rect 20898 29696 20904 29708
rect 20772 29668 20904 29696
rect 20772 29656 20778 29668
rect 20898 29656 20904 29668
rect 20956 29656 20962 29708
rect 21082 29656 21088 29708
rect 21140 29696 21146 29708
rect 21542 29696 21548 29708
rect 21140 29668 21548 29696
rect 21140 29656 21146 29668
rect 21542 29656 21548 29668
rect 21600 29696 21606 29708
rect 21729 29699 21787 29705
rect 21729 29696 21741 29699
rect 21600 29668 21741 29696
rect 21600 29656 21606 29668
rect 21729 29665 21741 29668
rect 21775 29665 21787 29699
rect 22554 29696 22560 29708
rect 22515 29668 22560 29696
rect 21729 29659 21787 29665
rect 22554 29656 22560 29668
rect 22612 29656 22618 29708
rect 22922 29696 22928 29708
rect 22883 29668 22928 29696
rect 22922 29656 22928 29668
rect 22980 29656 22986 29708
rect 23198 29696 23204 29708
rect 23159 29668 23204 29696
rect 23198 29656 23204 29668
rect 23256 29656 23262 29708
rect 24121 29699 24179 29705
rect 24121 29665 24133 29699
rect 24167 29696 24179 29699
rect 24394 29696 24400 29708
rect 24167 29668 24400 29696
rect 24167 29665 24179 29668
rect 24121 29659 24179 29665
rect 24394 29656 24400 29668
rect 24452 29656 24458 29708
rect 24673 29699 24731 29705
rect 24673 29665 24685 29699
rect 24719 29696 24731 29699
rect 24719 29668 25452 29696
rect 24719 29665 24731 29668
rect 24673 29659 24731 29665
rect 20088 29600 20208 29628
rect 18414 29560 18420 29572
rect 16991 29532 18276 29560
rect 18375 29532 18420 29560
rect 16991 29529 17003 29532
rect 16945 29523 17003 29529
rect 18414 29520 18420 29532
rect 18472 29520 18478 29572
rect 18782 29520 18788 29572
rect 18840 29560 18846 29572
rect 19981 29563 20039 29569
rect 19981 29560 19993 29563
rect 18840 29532 19993 29560
rect 18840 29520 18846 29532
rect 19981 29529 19993 29532
rect 20027 29529 20039 29563
rect 19981 29523 20039 29529
rect 4249 29495 4307 29501
rect 4249 29461 4261 29495
rect 4295 29492 4307 29495
rect 4614 29492 4620 29504
rect 4295 29464 4620 29492
rect 4295 29461 4307 29464
rect 4249 29455 4307 29461
rect 4614 29452 4620 29464
rect 4672 29452 4678 29504
rect 7466 29492 7472 29504
rect 7427 29464 7472 29492
rect 7466 29452 7472 29464
rect 7524 29452 7530 29504
rect 15194 29452 15200 29504
rect 15252 29492 15258 29504
rect 20088 29492 20116 29600
rect 20990 29588 20996 29640
rect 21048 29628 21054 29640
rect 22572 29628 22600 29656
rect 21048 29600 22600 29628
rect 24765 29631 24823 29637
rect 21048 29588 21054 29600
rect 24765 29597 24777 29631
rect 24811 29597 24823 29631
rect 25424 29628 25452 29668
rect 25498 29656 25504 29708
rect 25556 29696 25562 29708
rect 26528 29705 26556 29736
rect 27249 29733 27261 29736
rect 27295 29733 27307 29767
rect 27249 29727 27307 29733
rect 26513 29699 26571 29705
rect 25556 29668 25601 29696
rect 25556 29656 25562 29668
rect 26513 29665 26525 29699
rect 26559 29665 26571 29699
rect 26513 29659 26571 29665
rect 26602 29656 26608 29708
rect 26660 29696 26666 29708
rect 27614 29696 27620 29708
rect 26660 29668 27476 29696
rect 27575 29668 27620 29696
rect 26660 29656 26666 29668
rect 26694 29628 26700 29640
rect 25424 29600 26700 29628
rect 24765 29591 24823 29597
rect 20162 29520 20168 29572
rect 20220 29560 20226 29572
rect 21085 29563 21143 29569
rect 21085 29560 21097 29563
rect 20220 29532 21097 29560
rect 20220 29520 20226 29532
rect 21085 29529 21097 29532
rect 21131 29529 21143 29563
rect 23290 29560 23296 29572
rect 23251 29532 23296 29560
rect 21085 29523 21143 29529
rect 23290 29520 23296 29532
rect 23348 29520 23354 29572
rect 24210 29560 24216 29572
rect 24171 29532 24216 29560
rect 24210 29520 24216 29532
rect 24268 29520 24274 29572
rect 15252 29464 20116 29492
rect 21821 29495 21879 29501
rect 15252 29452 15258 29464
rect 21821 29461 21833 29495
rect 21867 29492 21879 29495
rect 24780 29492 24808 29591
rect 26694 29588 26700 29600
rect 26752 29588 26758 29640
rect 27246 29588 27252 29640
rect 27304 29628 27310 29640
rect 27341 29631 27399 29637
rect 27341 29628 27353 29631
rect 27304 29600 27353 29628
rect 27304 29588 27310 29600
rect 27341 29597 27353 29600
rect 27387 29597 27399 29631
rect 27448 29628 27476 29668
rect 27614 29656 27620 29668
rect 27672 29656 27678 29708
rect 28902 29656 28908 29708
rect 28960 29696 28966 29708
rect 29564 29705 29592 29804
rect 30098 29792 30104 29844
rect 30156 29832 30162 29844
rect 30466 29832 30472 29844
rect 30156 29804 30472 29832
rect 30156 29792 30162 29804
rect 30466 29792 30472 29804
rect 30524 29792 30530 29844
rect 30650 29792 30656 29844
rect 30708 29832 30714 29844
rect 30745 29835 30803 29841
rect 30745 29832 30757 29835
rect 30708 29804 30757 29832
rect 30708 29792 30714 29804
rect 30745 29801 30757 29804
rect 30791 29832 30803 29835
rect 31294 29832 31300 29844
rect 30791 29804 31300 29832
rect 30791 29801 30803 29804
rect 30745 29795 30803 29801
rect 31294 29792 31300 29804
rect 31352 29792 31358 29844
rect 32401 29835 32459 29841
rect 32401 29801 32413 29835
rect 32447 29832 32459 29835
rect 36262 29832 36268 29844
rect 32447 29804 36268 29832
rect 32447 29801 32459 29804
rect 32401 29795 32459 29801
rect 36262 29792 36268 29804
rect 36320 29792 36326 29844
rect 29638 29724 29644 29776
rect 29696 29764 29702 29776
rect 30834 29764 30840 29776
rect 29696 29736 30840 29764
rect 29696 29724 29702 29736
rect 30834 29724 30840 29736
rect 30892 29724 30898 29776
rect 31202 29764 31208 29776
rect 31163 29736 31208 29764
rect 31202 29724 31208 29736
rect 31260 29724 31266 29776
rect 36630 29724 36636 29776
rect 36688 29764 36694 29776
rect 36688 29736 37964 29764
rect 36688 29724 36694 29736
rect 37936 29708 37964 29736
rect 29457 29699 29515 29705
rect 29457 29696 29469 29699
rect 28960 29668 29469 29696
rect 28960 29656 28966 29668
rect 29457 29665 29469 29668
rect 29503 29665 29515 29699
rect 29457 29659 29515 29665
rect 29549 29699 29607 29705
rect 29549 29665 29561 29699
rect 29595 29665 29607 29699
rect 29549 29659 29607 29665
rect 30006 29656 30012 29708
rect 30064 29696 30070 29708
rect 30653 29699 30711 29705
rect 30653 29696 30665 29699
rect 30064 29668 30665 29696
rect 30064 29656 30070 29668
rect 30653 29665 30665 29668
rect 30699 29696 30711 29699
rect 31018 29696 31024 29708
rect 30699 29668 31024 29696
rect 30699 29665 30711 29668
rect 30653 29659 30711 29665
rect 31018 29656 31024 29668
rect 31076 29656 31082 29708
rect 32217 29699 32275 29705
rect 32217 29665 32229 29699
rect 32263 29696 32275 29699
rect 32953 29699 33011 29705
rect 32263 29668 32536 29696
rect 32263 29665 32275 29668
rect 32217 29659 32275 29665
rect 29822 29628 29828 29640
rect 27448 29600 29828 29628
rect 27341 29591 27399 29597
rect 29822 29588 29828 29600
rect 29880 29628 29886 29640
rect 30469 29631 30527 29637
rect 30469 29628 30481 29631
rect 29880 29600 30481 29628
rect 29880 29588 29886 29600
rect 30469 29597 30481 29600
rect 30515 29597 30527 29631
rect 30469 29591 30527 29597
rect 25682 29560 25688 29572
rect 25643 29532 25688 29560
rect 25682 29520 25688 29532
rect 25740 29520 25746 29572
rect 21867 29464 24808 29492
rect 21867 29461 21879 29464
rect 21821 29455 21879 29461
rect 26510 29452 26516 29504
rect 26568 29492 26574 29504
rect 26697 29495 26755 29501
rect 26697 29492 26709 29495
rect 26568 29464 26709 29492
rect 26568 29452 26574 29464
rect 26697 29461 26709 29464
rect 26743 29461 26755 29495
rect 26697 29455 26755 29461
rect 27249 29495 27307 29501
rect 27249 29461 27261 29495
rect 27295 29492 27307 29495
rect 27798 29492 27804 29504
rect 27295 29464 27804 29492
rect 27295 29461 27307 29464
rect 27249 29455 27307 29461
rect 27798 29452 27804 29464
rect 27856 29492 27862 29504
rect 28534 29492 28540 29504
rect 27856 29464 28540 29492
rect 27856 29452 27862 29464
rect 28534 29452 28540 29464
rect 28592 29452 28598 29504
rect 28905 29495 28963 29501
rect 28905 29461 28917 29495
rect 28951 29492 28963 29495
rect 29362 29492 29368 29504
rect 28951 29464 29368 29492
rect 28951 29461 28963 29464
rect 28905 29455 28963 29461
rect 29362 29452 29368 29464
rect 29420 29452 29426 29504
rect 29730 29492 29736 29504
rect 29691 29464 29736 29492
rect 29730 29452 29736 29464
rect 29788 29452 29794 29504
rect 32508 29492 32536 29668
rect 32953 29665 32965 29699
rect 32999 29696 33011 29699
rect 33042 29696 33048 29708
rect 32999 29668 33048 29696
rect 32999 29665 33011 29668
rect 32953 29659 33011 29665
rect 33042 29656 33048 29668
rect 33100 29656 33106 29708
rect 35526 29696 35532 29708
rect 35487 29668 35532 29696
rect 35526 29656 35532 29668
rect 35584 29656 35590 29708
rect 37734 29696 37740 29708
rect 37695 29668 37740 29696
rect 37734 29656 37740 29668
rect 37792 29656 37798 29708
rect 37918 29656 37924 29708
rect 37976 29696 37982 29708
rect 38105 29699 38163 29705
rect 38105 29696 38117 29699
rect 37976 29668 38117 29696
rect 37976 29656 37982 29668
rect 38105 29665 38117 29668
rect 38151 29665 38163 29699
rect 38562 29696 38568 29708
rect 38523 29668 38568 29696
rect 38105 29659 38163 29665
rect 38562 29656 38568 29668
rect 38620 29656 38626 29708
rect 33226 29628 33232 29640
rect 33187 29600 33232 29628
rect 33226 29588 33232 29600
rect 33284 29588 33290 29640
rect 35710 29588 35716 29640
rect 35768 29628 35774 29640
rect 35805 29631 35863 29637
rect 35805 29628 35817 29631
rect 35768 29600 35817 29628
rect 35768 29588 35774 29600
rect 35805 29597 35817 29600
rect 35851 29597 35863 29631
rect 35805 29591 35863 29597
rect 34422 29560 34428 29572
rect 33888 29532 34428 29560
rect 33888 29492 33916 29532
rect 34422 29520 34428 29532
rect 34480 29520 34486 29572
rect 38565 29563 38623 29569
rect 38565 29560 38577 29563
rect 36464 29532 38577 29560
rect 34514 29492 34520 29504
rect 32508 29464 33916 29492
rect 34475 29464 34520 29492
rect 34514 29452 34520 29464
rect 34572 29452 34578 29504
rect 36170 29452 36176 29504
rect 36228 29492 36234 29504
rect 36464 29492 36492 29532
rect 38565 29529 38577 29532
rect 38611 29529 38623 29563
rect 38565 29523 38623 29529
rect 36906 29492 36912 29504
rect 36228 29464 36492 29492
rect 36867 29464 36912 29492
rect 36228 29452 36234 29464
rect 36906 29452 36912 29464
rect 36964 29452 36970 29504
rect 1104 29402 39836 29424
rect 1104 29350 4246 29402
rect 4298 29350 4310 29402
rect 4362 29350 4374 29402
rect 4426 29350 4438 29402
rect 4490 29350 34966 29402
rect 35018 29350 35030 29402
rect 35082 29350 35094 29402
rect 35146 29350 35158 29402
rect 35210 29350 39836 29402
rect 1104 29328 39836 29350
rect 1486 29288 1492 29300
rect 1447 29260 1492 29288
rect 1486 29248 1492 29260
rect 1544 29248 1550 29300
rect 1670 29248 1676 29300
rect 1728 29288 1734 29300
rect 1949 29291 2007 29297
rect 1949 29288 1961 29291
rect 1728 29260 1961 29288
rect 1728 29248 1734 29260
rect 1949 29257 1961 29260
rect 1995 29257 2007 29291
rect 1949 29251 2007 29257
rect 5350 29248 5356 29300
rect 5408 29288 5414 29300
rect 7009 29291 7067 29297
rect 7009 29288 7021 29291
rect 5408 29260 7021 29288
rect 5408 29248 5414 29260
rect 7009 29257 7021 29260
rect 7055 29257 7067 29291
rect 7009 29251 7067 29257
rect 10870 29248 10876 29300
rect 10928 29288 10934 29300
rect 11238 29288 11244 29300
rect 10928 29260 11244 29288
rect 10928 29248 10934 29260
rect 11238 29248 11244 29260
rect 11296 29248 11302 29300
rect 11422 29288 11428 29300
rect 11383 29260 11428 29288
rect 11422 29248 11428 29260
rect 11480 29248 11486 29300
rect 11790 29248 11796 29300
rect 11848 29288 11854 29300
rect 14274 29288 14280 29300
rect 11848 29260 14280 29288
rect 11848 29248 11854 29260
rect 14274 29248 14280 29260
rect 14332 29248 14338 29300
rect 17586 29248 17592 29300
rect 17644 29288 17650 29300
rect 18322 29288 18328 29300
rect 17644 29260 18328 29288
rect 17644 29248 17650 29260
rect 18322 29248 18328 29260
rect 18380 29288 18386 29300
rect 20990 29288 20996 29300
rect 18380 29260 20996 29288
rect 18380 29248 18386 29260
rect 20990 29248 20996 29260
rect 21048 29248 21054 29300
rect 21177 29291 21235 29297
rect 21177 29257 21189 29291
rect 21223 29288 21235 29291
rect 23198 29288 23204 29300
rect 21223 29260 23204 29288
rect 21223 29257 21235 29260
rect 21177 29251 21235 29257
rect 23198 29248 23204 29260
rect 23256 29248 23262 29300
rect 25314 29248 25320 29300
rect 25372 29288 25378 29300
rect 25501 29291 25559 29297
rect 25501 29288 25513 29291
rect 25372 29260 25513 29288
rect 25372 29248 25378 29260
rect 25501 29257 25513 29260
rect 25547 29257 25559 29291
rect 25501 29251 25559 29257
rect 26326 29248 26332 29300
rect 26384 29288 26390 29300
rect 27157 29291 27215 29297
rect 27157 29288 27169 29291
rect 26384 29260 27169 29288
rect 26384 29248 26390 29260
rect 27157 29257 27169 29260
rect 27203 29257 27215 29291
rect 30006 29288 30012 29300
rect 27157 29251 27215 29257
rect 27908 29260 30012 29288
rect 2700 29192 4660 29220
rect 1854 29112 1860 29164
rect 1912 29152 1918 29164
rect 2700 29161 2728 29192
rect 2685 29155 2743 29161
rect 2685 29152 2697 29155
rect 1912 29124 2697 29152
rect 1912 29112 1918 29124
rect 2685 29121 2697 29124
rect 2731 29121 2743 29155
rect 3142 29152 3148 29164
rect 2685 29115 2743 29121
rect 2884 29124 3148 29152
rect 1762 29084 1768 29096
rect 1723 29056 1768 29084
rect 1762 29044 1768 29056
rect 1820 29044 1826 29096
rect 2884 29093 2912 29124
rect 3142 29112 3148 29124
rect 3200 29112 3206 29164
rect 3326 29112 3332 29164
rect 3384 29152 3390 29164
rect 4632 29161 4660 29192
rect 9214 29180 9220 29232
rect 9272 29220 9278 29232
rect 9272 29192 14964 29220
rect 9272 29180 9278 29192
rect 3421 29155 3479 29161
rect 3421 29152 3433 29155
rect 3384 29124 3433 29152
rect 3384 29112 3390 29124
rect 3421 29121 3433 29124
rect 3467 29121 3479 29155
rect 3421 29115 3479 29121
rect 4617 29155 4675 29161
rect 4617 29121 4629 29155
rect 4663 29152 4675 29155
rect 4982 29152 4988 29164
rect 4663 29124 4988 29152
rect 4663 29121 4675 29124
rect 4617 29115 4675 29121
rect 4982 29112 4988 29124
rect 5040 29112 5046 29164
rect 5718 29152 5724 29164
rect 5679 29124 5724 29152
rect 5718 29112 5724 29124
rect 5776 29112 5782 29164
rect 7466 29152 7472 29164
rect 6104 29124 7472 29152
rect 2869 29087 2927 29093
rect 2869 29053 2881 29087
rect 2915 29053 2927 29087
rect 2869 29047 2927 29053
rect 2961 29087 3019 29093
rect 2961 29053 2973 29087
rect 3007 29084 3019 29087
rect 3510 29084 3516 29096
rect 3007 29056 3516 29084
rect 3007 29053 3019 29056
rect 2961 29047 3019 29053
rect 3510 29044 3516 29056
rect 3568 29044 3574 29096
rect 4157 29087 4215 29093
rect 4157 29053 4169 29087
rect 4203 29053 4215 29087
rect 4157 29047 4215 29053
rect 4433 29087 4491 29093
rect 4433 29053 4445 29087
rect 4479 29084 4491 29087
rect 5258 29084 5264 29096
rect 4479 29056 5120 29084
rect 5219 29056 5264 29084
rect 4479 29053 4491 29056
rect 4433 29047 4491 29053
rect 1673 29019 1731 29025
rect 1673 28985 1685 29019
rect 1719 29016 1731 29019
rect 2038 29016 2044 29028
rect 1719 28988 2044 29016
rect 1719 28985 1731 28988
rect 1673 28979 1731 28985
rect 2038 28976 2044 28988
rect 2096 28976 2102 29028
rect 2774 28976 2780 29028
rect 2832 29016 2838 29028
rect 3053 29019 3111 29025
rect 3053 29016 3065 29019
rect 2832 28988 3065 29016
rect 2832 28976 2838 28988
rect 3053 28985 3065 28988
rect 3099 28985 3111 29019
rect 4172 29016 4200 29047
rect 4614 29016 4620 29028
rect 4172 28988 4620 29016
rect 3053 28979 3111 28985
rect 4614 28976 4620 28988
rect 4672 28976 4678 29028
rect 5092 29016 5120 29056
rect 5258 29044 5264 29056
rect 5316 29044 5322 29096
rect 5537 29087 5595 29093
rect 5537 29053 5549 29087
rect 5583 29084 5595 29087
rect 5810 29084 5816 29096
rect 5583 29056 5816 29084
rect 5583 29053 5595 29056
rect 5537 29047 5595 29053
rect 5810 29044 5816 29056
rect 5868 29044 5874 29096
rect 6104 29093 6132 29124
rect 7466 29112 7472 29124
rect 7524 29112 7530 29164
rect 7561 29155 7619 29161
rect 7561 29121 7573 29155
rect 7607 29152 7619 29155
rect 7607 29124 8432 29152
rect 7607 29121 7619 29124
rect 7561 29115 7619 29121
rect 6089 29087 6147 29093
rect 6089 29053 6101 29087
rect 6135 29053 6147 29087
rect 6089 29047 6147 29053
rect 6825 29087 6883 29093
rect 6825 29053 6837 29087
rect 6871 29084 6883 29087
rect 7006 29084 7012 29096
rect 6871 29056 7012 29084
rect 6871 29053 6883 29056
rect 6825 29047 6883 29053
rect 7006 29044 7012 29056
rect 7064 29044 7070 29096
rect 7837 29087 7895 29093
rect 7837 29053 7849 29087
rect 7883 29084 7895 29087
rect 8294 29084 8300 29096
rect 7883 29056 8300 29084
rect 7883 29053 7895 29056
rect 7837 29047 7895 29053
rect 8294 29044 8300 29056
rect 8352 29044 8358 29096
rect 8404 29084 8432 29124
rect 8478 29112 8484 29164
rect 8536 29152 8542 29164
rect 9769 29155 9827 29161
rect 9769 29152 9781 29155
rect 8536 29124 9781 29152
rect 8536 29112 8542 29124
rect 9769 29121 9781 29124
rect 9815 29121 9827 29155
rect 9769 29115 9827 29121
rect 12434 29112 12440 29164
rect 12492 29152 12498 29164
rect 12492 29124 14228 29152
rect 12492 29112 12498 29124
rect 9306 29084 9312 29096
rect 8404 29056 9312 29084
rect 9306 29044 9312 29056
rect 9364 29044 9370 29096
rect 9950 29084 9956 29096
rect 9911 29056 9956 29084
rect 9950 29044 9956 29056
rect 10008 29044 10014 29096
rect 10134 29084 10140 29096
rect 10095 29056 10140 29084
rect 10134 29044 10140 29056
rect 10192 29044 10198 29096
rect 10410 29084 10416 29096
rect 10371 29056 10416 29084
rect 10410 29044 10416 29056
rect 10468 29044 10474 29096
rect 11333 29087 11391 29093
rect 11333 29053 11345 29087
rect 11379 29053 11391 29087
rect 11333 29047 11391 29053
rect 13265 29087 13323 29093
rect 13265 29053 13277 29087
rect 13311 29084 13323 29087
rect 13354 29084 13360 29096
rect 13311 29056 13360 29084
rect 13311 29053 13323 29056
rect 13265 29047 13323 29053
rect 5626 29016 5632 29028
rect 5092 28988 5632 29016
rect 5626 28976 5632 28988
rect 5684 29016 5690 29028
rect 5994 29016 6000 29028
rect 5684 28988 6000 29016
rect 5684 28976 5690 28988
rect 5994 28976 6000 28988
rect 6052 28976 6058 29028
rect 9030 28976 9036 29028
rect 9088 29016 9094 29028
rect 9217 29019 9275 29025
rect 9217 29016 9229 29019
rect 9088 28988 9229 29016
rect 9088 28976 9094 28988
rect 9217 28985 9229 28988
rect 9263 29016 9275 29019
rect 11348 29016 11376 29047
rect 13354 29044 13360 29056
rect 13412 29044 13418 29096
rect 13538 29084 13544 29096
rect 13499 29056 13544 29084
rect 13538 29044 13544 29056
rect 13596 29044 13602 29096
rect 13722 29084 13728 29096
rect 13683 29056 13728 29084
rect 13722 29044 13728 29056
rect 13780 29044 13786 29096
rect 14200 29093 14228 29124
rect 14185 29087 14243 29093
rect 14185 29053 14197 29087
rect 14231 29053 14243 29087
rect 14185 29047 14243 29053
rect 14274 29044 14280 29096
rect 14332 29084 14338 29096
rect 14642 29084 14648 29096
rect 14332 29056 14648 29084
rect 14332 29044 14338 29056
rect 14642 29044 14648 29056
rect 14700 29044 14706 29096
rect 14936 29093 14964 29192
rect 17310 29180 17316 29232
rect 17368 29220 17374 29232
rect 17405 29223 17463 29229
rect 17405 29220 17417 29223
rect 17368 29192 17417 29220
rect 17368 29180 17374 29192
rect 17405 29189 17417 29192
rect 17451 29220 17463 29223
rect 18782 29220 18788 29232
rect 17451 29192 18788 29220
rect 17451 29189 17463 29192
rect 17405 29183 17463 29189
rect 18782 29180 18788 29192
rect 18840 29180 18846 29232
rect 18969 29223 19027 29229
rect 18969 29189 18981 29223
rect 19015 29220 19027 29223
rect 23934 29220 23940 29232
rect 19015 29192 19932 29220
rect 19015 29189 19027 29192
rect 18969 29183 19027 29189
rect 15841 29155 15899 29161
rect 15841 29121 15853 29155
rect 15887 29152 15899 29155
rect 15887 29124 19288 29152
rect 15887 29121 15899 29124
rect 15841 29115 15899 29121
rect 14921 29087 14979 29093
rect 14921 29053 14933 29087
rect 14967 29053 14979 29087
rect 14921 29047 14979 29053
rect 15473 29087 15531 29093
rect 15473 29053 15485 29087
rect 15519 29084 15531 29087
rect 15654 29084 15660 29096
rect 15519 29056 15660 29084
rect 15519 29053 15531 29056
rect 15473 29047 15531 29053
rect 15654 29044 15660 29056
rect 15712 29084 15718 29096
rect 15930 29084 15936 29096
rect 15712 29056 15936 29084
rect 15712 29044 15718 29056
rect 15930 29044 15936 29056
rect 15988 29044 15994 29096
rect 16301 29087 16359 29093
rect 16301 29053 16313 29087
rect 16347 29084 16359 29087
rect 16390 29084 16396 29096
rect 16347 29056 16396 29084
rect 16347 29053 16359 29056
rect 16301 29047 16359 29053
rect 16390 29044 16396 29056
rect 16448 29044 16454 29096
rect 16577 29087 16635 29093
rect 16577 29053 16589 29087
rect 16623 29084 16635 29087
rect 16942 29084 16948 29096
rect 16623 29056 16948 29084
rect 16623 29053 16635 29056
rect 16577 29047 16635 29053
rect 16942 29044 16948 29056
rect 17000 29044 17006 29096
rect 17218 29084 17224 29096
rect 17179 29056 17224 29084
rect 17218 29044 17224 29056
rect 17276 29044 17282 29096
rect 17954 29044 17960 29096
rect 18012 29084 18018 29096
rect 18049 29087 18107 29093
rect 18049 29084 18061 29087
rect 18012 29056 18061 29084
rect 18012 29044 18018 29056
rect 18049 29053 18061 29056
rect 18095 29053 18107 29087
rect 18414 29084 18420 29096
rect 18375 29056 18420 29084
rect 18049 29047 18107 29053
rect 18414 29044 18420 29056
rect 18472 29044 18478 29096
rect 18877 29087 18935 29093
rect 18877 29053 18889 29087
rect 18923 29053 18935 29087
rect 18877 29047 18935 29053
rect 9263 28988 11376 29016
rect 12713 29019 12771 29025
rect 9263 28985 9275 28988
rect 9217 28979 9275 28985
rect 12713 28985 12725 29019
rect 12759 29016 12771 29019
rect 14550 29016 14556 29028
rect 12759 28988 14556 29016
rect 12759 28985 12771 28988
rect 12713 28979 12771 28985
rect 14550 28976 14556 28988
rect 14608 28976 14614 29028
rect 17494 28976 17500 29028
rect 17552 29016 17558 29028
rect 18892 29016 18920 29047
rect 17552 28988 18920 29016
rect 19260 29016 19288 29124
rect 19426 29044 19432 29096
rect 19484 29084 19490 29096
rect 19613 29087 19671 29093
rect 19613 29084 19625 29087
rect 19484 29056 19625 29084
rect 19484 29044 19490 29056
rect 19613 29053 19625 29056
rect 19659 29053 19671 29087
rect 19904 29084 19932 29192
rect 19996 29192 23940 29220
rect 19996 29161 20024 29192
rect 23934 29180 23940 29192
rect 23992 29180 23998 29232
rect 24394 29220 24400 29232
rect 24355 29192 24400 29220
rect 24394 29180 24400 29192
rect 24452 29180 24458 29232
rect 19981 29155 20039 29161
rect 19981 29121 19993 29155
rect 20027 29121 20039 29155
rect 19981 29115 20039 29121
rect 20088 29124 26740 29152
rect 20088 29084 20116 29124
rect 19904 29056 20116 29084
rect 20349 29087 20407 29093
rect 19613 29047 19671 29053
rect 20349 29053 20361 29087
rect 20395 29084 20407 29087
rect 20530 29084 20536 29096
rect 20395 29056 20536 29084
rect 20395 29053 20407 29056
rect 20349 29047 20407 29053
rect 20530 29044 20536 29056
rect 20588 29044 20594 29096
rect 21008 29056 21220 29084
rect 21008 29016 21036 29056
rect 19260 28988 21036 29016
rect 21192 29016 21220 29056
rect 21358 29044 21364 29096
rect 21416 29084 21422 29096
rect 21729 29087 21787 29093
rect 21729 29084 21741 29087
rect 21416 29056 21741 29084
rect 21416 29044 21422 29056
rect 21729 29053 21741 29056
rect 21775 29053 21787 29087
rect 21729 29047 21787 29053
rect 21818 29044 21824 29096
rect 21876 29084 21882 29096
rect 21876 29056 21921 29084
rect 21876 29044 21882 29056
rect 22002 29044 22008 29096
rect 22060 29084 22066 29096
rect 22097 29087 22155 29093
rect 22097 29084 22109 29087
rect 22060 29056 22109 29084
rect 22060 29044 22066 29056
rect 22097 29053 22109 29056
rect 22143 29053 22155 29087
rect 22097 29047 22155 29053
rect 22281 29087 22339 29093
rect 22281 29053 22293 29087
rect 22327 29084 22339 29087
rect 22830 29084 22836 29096
rect 22327 29056 22836 29084
rect 22327 29053 22339 29056
rect 22281 29047 22339 29053
rect 22830 29044 22836 29056
rect 22888 29044 22894 29096
rect 22925 29087 22983 29093
rect 22925 29053 22937 29087
rect 22971 29084 22983 29087
rect 23842 29084 23848 29096
rect 22971 29056 23848 29084
rect 22971 29053 22983 29056
rect 22925 29047 22983 29053
rect 23842 29044 23848 29056
rect 23900 29044 23906 29096
rect 23937 29087 23995 29093
rect 23937 29053 23949 29087
rect 23983 29084 23995 29087
rect 24026 29084 24032 29096
rect 23983 29056 24032 29084
rect 23983 29053 23995 29056
rect 23937 29047 23995 29053
rect 24026 29044 24032 29056
rect 24084 29044 24090 29096
rect 24486 29084 24492 29096
rect 24447 29056 24492 29084
rect 24486 29044 24492 29056
rect 24544 29044 24550 29096
rect 24578 29044 24584 29096
rect 24636 29084 24642 29096
rect 24673 29087 24731 29093
rect 24673 29084 24685 29087
rect 24636 29056 24685 29084
rect 24636 29044 24642 29056
rect 24673 29053 24685 29056
rect 24719 29053 24731 29087
rect 25317 29087 25375 29093
rect 25317 29084 25329 29087
rect 24673 29047 24731 29053
rect 25056 29056 25329 29084
rect 24946 29016 24952 29028
rect 21192 28988 24952 29016
rect 17552 28976 17558 28988
rect 24946 28976 24952 28988
rect 25004 28976 25010 29028
rect 9858 28908 9864 28960
rect 9916 28948 9922 28960
rect 10134 28948 10140 28960
rect 9916 28920 10140 28948
rect 9916 28908 9922 28920
rect 10134 28908 10140 28920
rect 10192 28908 10198 28960
rect 20254 28908 20260 28960
rect 20312 28948 20318 28960
rect 22830 28948 22836 28960
rect 20312 28920 22836 28948
rect 20312 28908 20318 28920
rect 22830 28908 22836 28920
rect 22888 28908 22894 28960
rect 23017 28951 23075 28957
rect 23017 28917 23029 28951
rect 23063 28948 23075 28951
rect 25056 28948 25084 29056
rect 25317 29053 25329 29056
rect 25363 29084 25375 29087
rect 25958 29084 25964 29096
rect 25363 29056 25964 29084
rect 25363 29053 25375 29056
rect 25317 29047 25375 29053
rect 25958 29044 25964 29056
rect 26016 29044 26022 29096
rect 26050 29044 26056 29096
rect 26108 29084 26114 29096
rect 26186 29087 26244 29093
rect 26108 29056 26153 29084
rect 26108 29044 26114 29056
rect 26186 29053 26198 29087
rect 26232 29053 26244 29087
rect 26602 29084 26608 29096
rect 26563 29056 26608 29084
rect 26186 29047 26244 29053
rect 26201 29016 26229 29047
rect 26602 29044 26608 29056
rect 26660 29044 26666 29096
rect 25976 28988 26229 29016
rect 26712 29016 26740 29124
rect 26970 29112 26976 29164
rect 27028 29152 27034 29164
rect 27908 29152 27936 29260
rect 30006 29248 30012 29260
rect 30064 29248 30070 29300
rect 36446 29248 36452 29300
rect 36504 29288 36510 29300
rect 38749 29291 38807 29297
rect 38749 29288 38761 29291
rect 36504 29260 38761 29288
rect 36504 29248 36510 29260
rect 38749 29257 38761 29260
rect 38795 29257 38807 29291
rect 38749 29251 38807 29257
rect 27985 29223 28043 29229
rect 27985 29189 27997 29223
rect 28031 29189 28043 29223
rect 27985 29183 28043 29189
rect 27028 29124 27936 29152
rect 28000 29152 28028 29183
rect 28166 29180 28172 29232
rect 28224 29220 28230 29232
rect 28994 29220 29000 29232
rect 28224 29192 29000 29220
rect 28224 29180 28230 29192
rect 28994 29180 29000 29192
rect 29052 29180 29058 29232
rect 30282 29180 30288 29232
rect 30340 29220 30346 29232
rect 30653 29223 30711 29229
rect 30653 29220 30665 29223
rect 30340 29192 30665 29220
rect 30340 29180 30346 29192
rect 30653 29189 30665 29192
rect 30699 29189 30711 29223
rect 30653 29183 30711 29189
rect 33045 29223 33103 29229
rect 33045 29189 33057 29223
rect 33091 29220 33103 29223
rect 33226 29220 33232 29232
rect 33091 29192 33232 29220
rect 33091 29189 33103 29192
rect 33045 29183 33103 29189
rect 33226 29180 33232 29192
rect 33284 29180 33290 29232
rect 35710 29220 35716 29232
rect 35671 29192 35716 29220
rect 35710 29180 35716 29192
rect 35768 29180 35774 29232
rect 37277 29223 37335 29229
rect 37277 29189 37289 29223
rect 37323 29220 37335 29223
rect 37550 29220 37556 29232
rect 37323 29192 37556 29220
rect 37323 29189 37335 29192
rect 37277 29183 37335 29189
rect 37550 29180 37556 29192
rect 37608 29180 37614 29232
rect 36446 29152 36452 29164
rect 28000 29124 33364 29152
rect 36407 29124 36452 29152
rect 27028 29112 27034 29124
rect 27065 29087 27123 29093
rect 27065 29053 27077 29087
rect 27111 29084 27123 29087
rect 27798 29084 27804 29096
rect 27111 29056 27804 29084
rect 27111 29053 27123 29056
rect 27065 29047 27123 29053
rect 27798 29044 27804 29056
rect 27856 29044 27862 29096
rect 28166 29084 28172 29096
rect 28127 29056 28172 29084
rect 28166 29044 28172 29056
rect 28224 29044 28230 29096
rect 28537 29087 28595 29093
rect 28537 29053 28549 29087
rect 28583 29053 28595 29087
rect 28537 29047 28595 29053
rect 28629 29087 28687 29093
rect 28629 29053 28641 29087
rect 28675 29084 28687 29087
rect 29086 29084 29092 29096
rect 28675 29056 29092 29084
rect 28675 29053 28687 29056
rect 28629 29047 28687 29053
rect 28552 29016 28580 29047
rect 29086 29044 29092 29056
rect 29144 29044 29150 29096
rect 29178 29044 29184 29096
rect 29236 29084 29242 29096
rect 29273 29087 29331 29093
rect 29273 29084 29285 29087
rect 29236 29056 29285 29084
rect 29236 29044 29242 29056
rect 29273 29053 29285 29056
rect 29319 29053 29331 29087
rect 29546 29084 29552 29096
rect 29507 29056 29552 29084
rect 29273 29047 29331 29053
rect 29546 29044 29552 29056
rect 29604 29044 29610 29096
rect 31849 29087 31907 29093
rect 31849 29053 31861 29087
rect 31895 29084 31907 29087
rect 32030 29084 32036 29096
rect 31895 29056 32036 29084
rect 31895 29053 31907 29056
rect 31849 29047 31907 29053
rect 32030 29044 32036 29056
rect 32088 29044 32094 29096
rect 33336 29093 33364 29124
rect 36446 29112 36452 29124
rect 36504 29112 36510 29164
rect 32125 29087 32183 29093
rect 32125 29053 32137 29087
rect 32171 29053 32183 29087
rect 32125 29047 32183 29053
rect 32309 29087 32367 29093
rect 32309 29053 32321 29087
rect 32355 29084 32367 29087
rect 32769 29087 32827 29093
rect 32769 29084 32781 29087
rect 32355 29056 32781 29084
rect 32355 29053 32367 29056
rect 32309 29047 32367 29053
rect 32769 29053 32781 29056
rect 32815 29053 32827 29087
rect 32769 29047 32827 29053
rect 33321 29087 33379 29093
rect 33321 29053 33333 29087
rect 33367 29053 33379 29087
rect 33321 29047 33379 29053
rect 33781 29087 33839 29093
rect 33781 29053 33793 29087
rect 33827 29084 33839 29087
rect 34146 29084 34152 29096
rect 33827 29056 34152 29084
rect 33827 29053 33839 29056
rect 33781 29047 33839 29053
rect 26712 28988 28580 29016
rect 32140 29016 32168 29047
rect 34146 29044 34152 29056
rect 34204 29044 34210 29096
rect 35434 29084 35440 29096
rect 35395 29056 35440 29084
rect 35434 29044 35440 29056
rect 35492 29044 35498 29096
rect 36170 29084 36176 29096
rect 36131 29056 36176 29084
rect 36170 29044 36176 29056
rect 36228 29044 36234 29096
rect 36354 29044 36360 29096
rect 36412 29084 36418 29096
rect 37001 29087 37059 29093
rect 37001 29084 37013 29087
rect 36412 29056 37013 29084
rect 36412 29044 36418 29056
rect 37001 29053 37013 29056
rect 37047 29053 37059 29087
rect 37001 29047 37059 29053
rect 37737 29087 37795 29093
rect 37737 29053 37749 29087
rect 37783 29053 37795 29087
rect 37737 29047 37795 29053
rect 34514 29016 34520 29028
rect 32140 28988 34520 29016
rect 25976 28960 26004 28988
rect 34514 28976 34520 28988
rect 34572 28976 34578 29028
rect 37752 29016 37780 29047
rect 37826 29044 37832 29096
rect 37884 29084 37890 29096
rect 37884 29056 37929 29084
rect 37884 29044 37890 29056
rect 38470 29044 38476 29096
rect 38528 29084 38534 29096
rect 38565 29087 38623 29093
rect 38565 29084 38577 29087
rect 38528 29056 38577 29084
rect 38528 29044 38534 29056
rect 38565 29053 38577 29056
rect 38611 29053 38623 29087
rect 38565 29047 38623 29053
rect 38654 29016 38660 29028
rect 37752 28988 38660 29016
rect 38654 28976 38660 28988
rect 38712 28976 38718 29028
rect 23063 28920 25084 28948
rect 23063 28917 23075 28920
rect 23017 28911 23075 28917
rect 25958 28908 25964 28960
rect 26016 28908 26022 28960
rect 26234 28908 26240 28960
rect 26292 28948 26298 28960
rect 33134 28948 33140 28960
rect 26292 28920 33140 28948
rect 26292 28908 26298 28920
rect 33134 28908 33140 28920
rect 33192 28908 33198 28960
rect 1104 28858 39836 28880
rect 1104 28806 19606 28858
rect 19658 28806 19670 28858
rect 19722 28806 19734 28858
rect 19786 28806 19798 28858
rect 19850 28806 39836 28858
rect 1104 28784 39836 28806
rect 2866 28704 2872 28756
rect 2924 28744 2930 28756
rect 3234 28744 3240 28756
rect 2924 28716 3240 28744
rect 2924 28704 2930 28716
rect 3234 28704 3240 28716
rect 3292 28704 3298 28756
rect 4798 28744 4804 28756
rect 4759 28716 4804 28744
rect 4798 28704 4804 28716
rect 4856 28704 4862 28756
rect 7006 28704 7012 28756
rect 7064 28744 7070 28756
rect 7469 28747 7527 28753
rect 7469 28744 7481 28747
rect 7064 28716 7481 28744
rect 7064 28704 7070 28716
rect 7469 28713 7481 28716
rect 7515 28713 7527 28747
rect 8294 28744 8300 28756
rect 8255 28716 8300 28744
rect 7469 28707 7527 28713
rect 8294 28704 8300 28716
rect 8352 28704 8358 28756
rect 9033 28747 9091 28753
rect 9033 28713 9045 28747
rect 9079 28744 9091 28747
rect 10410 28744 10416 28756
rect 9079 28716 10416 28744
rect 9079 28713 9091 28716
rect 9033 28707 9091 28713
rect 10410 28704 10416 28716
rect 10468 28704 10474 28756
rect 13446 28704 13452 28756
rect 13504 28744 13510 28756
rect 16666 28744 16672 28756
rect 13504 28716 16672 28744
rect 13504 28704 13510 28716
rect 16666 28704 16672 28716
rect 16724 28704 16730 28756
rect 17126 28704 17132 28756
rect 17184 28744 17190 28756
rect 17184 28716 18276 28744
rect 17184 28704 17190 28716
rect 5626 28676 5632 28688
rect 5368 28648 5632 28676
rect 4614 28608 4620 28620
rect 4575 28580 4620 28608
rect 4614 28568 4620 28580
rect 4672 28568 4678 28620
rect 5368 28617 5396 28648
rect 5626 28636 5632 28648
rect 5684 28636 5690 28688
rect 12253 28679 12311 28685
rect 12253 28645 12265 28679
rect 12299 28676 12311 28679
rect 12434 28676 12440 28688
rect 12299 28648 12440 28676
rect 12299 28645 12311 28648
rect 12253 28639 12311 28645
rect 12434 28636 12440 28648
rect 12492 28636 12498 28688
rect 16684 28676 16712 28704
rect 17402 28676 17408 28688
rect 16684 28648 17408 28676
rect 17402 28636 17408 28648
rect 17460 28636 17466 28688
rect 17954 28676 17960 28688
rect 17915 28648 17960 28676
rect 17954 28636 17960 28648
rect 18012 28636 18018 28688
rect 18248 28620 18276 28716
rect 19150 28704 19156 28756
rect 19208 28744 19214 28756
rect 20254 28744 20260 28756
rect 19208 28716 20260 28744
rect 19208 28704 19214 28716
rect 20254 28704 20260 28716
rect 20312 28704 20318 28756
rect 21450 28704 21456 28756
rect 21508 28744 21514 28756
rect 22462 28744 22468 28756
rect 21508 28716 22468 28744
rect 21508 28704 21514 28716
rect 22462 28704 22468 28716
rect 22520 28744 22526 28756
rect 26510 28744 26516 28756
rect 22520 28716 26516 28744
rect 22520 28704 22526 28716
rect 24029 28679 24087 28685
rect 19076 28648 19472 28676
rect 5353 28611 5411 28617
rect 5353 28577 5365 28611
rect 5399 28577 5411 28611
rect 5353 28571 5411 28577
rect 5534 28568 5540 28620
rect 5592 28608 5598 28620
rect 6365 28611 6423 28617
rect 6365 28608 6377 28611
rect 5592 28580 6377 28608
rect 5592 28568 5598 28580
rect 6365 28577 6377 28580
rect 6411 28577 6423 28611
rect 6365 28571 6423 28577
rect 8205 28611 8263 28617
rect 8205 28577 8217 28611
rect 8251 28608 8263 28611
rect 8478 28608 8484 28620
rect 8251 28580 8484 28608
rect 8251 28577 8263 28580
rect 8205 28571 8263 28577
rect 8478 28568 8484 28580
rect 8536 28568 8542 28620
rect 8938 28608 8944 28620
rect 8899 28580 8944 28608
rect 8938 28568 8944 28580
rect 8996 28568 9002 28620
rect 9122 28568 9128 28620
rect 9180 28608 9186 28620
rect 9677 28611 9735 28617
rect 9677 28608 9689 28611
rect 9180 28580 9689 28608
rect 9180 28568 9186 28580
rect 9677 28577 9689 28580
rect 9723 28577 9735 28611
rect 9677 28571 9735 28577
rect 10873 28611 10931 28617
rect 10873 28577 10885 28611
rect 10919 28608 10931 28611
rect 11330 28608 11336 28620
rect 10919 28580 11336 28608
rect 10919 28577 10931 28580
rect 10873 28571 10931 28577
rect 11330 28568 11336 28580
rect 11388 28568 11394 28620
rect 11514 28568 11520 28620
rect 11572 28608 11578 28620
rect 15289 28611 15347 28617
rect 15289 28608 15301 28611
rect 11572 28580 15301 28608
rect 11572 28568 11578 28580
rect 15289 28577 15301 28580
rect 15335 28577 15347 28611
rect 15654 28608 15660 28620
rect 15615 28580 15660 28608
rect 15289 28571 15347 28577
rect 15654 28568 15660 28580
rect 15712 28568 15718 28620
rect 16390 28568 16396 28620
rect 16448 28608 16454 28620
rect 16577 28611 16635 28617
rect 16577 28608 16589 28611
rect 16448 28580 16589 28608
rect 16448 28568 16454 28580
rect 16577 28577 16589 28580
rect 16623 28577 16635 28611
rect 16942 28608 16948 28620
rect 16855 28580 16948 28608
rect 16577 28571 16635 28577
rect 16942 28568 16948 28580
rect 17000 28608 17006 28620
rect 17865 28611 17923 28617
rect 17000 28580 17632 28608
rect 17000 28568 17006 28580
rect 1394 28500 1400 28552
rect 1452 28540 1458 28552
rect 1673 28543 1731 28549
rect 1673 28540 1685 28543
rect 1452 28512 1685 28540
rect 1452 28500 1458 28512
rect 1673 28509 1685 28512
rect 1719 28509 1731 28543
rect 1673 28503 1731 28509
rect 1949 28543 2007 28549
rect 1949 28509 1961 28543
rect 1995 28540 2007 28543
rect 4062 28540 4068 28552
rect 1995 28512 4068 28540
rect 1995 28509 2007 28512
rect 1949 28503 2007 28509
rect 4062 28500 4068 28512
rect 4120 28500 4126 28552
rect 5442 28540 5448 28552
rect 5403 28512 5448 28540
rect 5442 28500 5448 28512
rect 5500 28500 5506 28552
rect 6089 28543 6147 28549
rect 6089 28509 6101 28543
rect 6135 28540 6147 28543
rect 6546 28540 6552 28552
rect 6135 28512 6552 28540
rect 6135 28509 6147 28512
rect 6089 28503 6147 28509
rect 6546 28500 6552 28512
rect 6604 28500 6610 28552
rect 9306 28500 9312 28552
rect 9364 28540 9370 28552
rect 10597 28543 10655 28549
rect 10597 28540 10609 28543
rect 9364 28512 10609 28540
rect 9364 28500 9370 28512
rect 10597 28509 10609 28512
rect 10643 28509 10655 28543
rect 13078 28540 13084 28552
rect 13039 28512 13084 28540
rect 10597 28503 10655 28509
rect 13078 28500 13084 28512
rect 13136 28500 13142 28552
rect 13357 28543 13415 28549
rect 13357 28509 13369 28543
rect 13403 28540 13415 28543
rect 15194 28540 15200 28552
rect 13403 28512 15200 28540
rect 13403 28509 13415 28512
rect 13357 28503 13415 28509
rect 15194 28500 15200 28512
rect 15252 28500 15258 28552
rect 16209 28475 16267 28481
rect 16209 28441 16221 28475
rect 16255 28472 16267 28475
rect 16666 28472 16672 28484
rect 16255 28444 16672 28472
rect 16255 28441 16267 28444
rect 16209 28435 16267 28441
rect 16666 28432 16672 28444
rect 16724 28432 16730 28484
rect 17604 28472 17632 28580
rect 17865 28577 17877 28611
rect 17911 28577 17923 28611
rect 18230 28608 18236 28620
rect 18191 28580 18236 28608
rect 17865 28571 17923 28577
rect 17880 28540 17908 28571
rect 18230 28568 18236 28580
rect 18288 28568 18294 28620
rect 18693 28611 18751 28617
rect 18693 28577 18705 28611
rect 18739 28608 18751 28611
rect 18966 28608 18972 28620
rect 18739 28580 18972 28608
rect 18739 28577 18751 28580
rect 18693 28571 18751 28577
rect 18966 28568 18972 28580
rect 19024 28568 19030 28620
rect 19076 28617 19104 28648
rect 19444 28620 19472 28648
rect 24029 28645 24041 28679
rect 24075 28676 24087 28679
rect 24075 28648 25636 28676
rect 24075 28645 24087 28648
rect 24029 28639 24087 28645
rect 19061 28611 19119 28617
rect 19061 28577 19073 28611
rect 19107 28577 19119 28611
rect 19334 28608 19340 28620
rect 19061 28571 19119 28577
rect 19168 28580 19340 28608
rect 18322 28540 18328 28552
rect 17880 28512 18328 28540
rect 18322 28500 18328 28512
rect 18380 28500 18386 28552
rect 19168 28472 19196 28580
rect 19334 28568 19340 28580
rect 19392 28568 19398 28620
rect 19426 28568 19432 28620
rect 19484 28568 19490 28620
rect 19521 28611 19579 28617
rect 19521 28577 19533 28611
rect 19567 28577 19579 28611
rect 19521 28571 19579 28577
rect 19981 28611 20039 28617
rect 19981 28577 19993 28611
rect 20027 28577 20039 28611
rect 19981 28571 20039 28577
rect 20901 28611 20959 28617
rect 20901 28577 20913 28611
rect 20947 28608 20959 28611
rect 20947 28580 21128 28608
rect 20947 28577 20959 28580
rect 20901 28571 20959 28577
rect 17604 28444 19196 28472
rect 7650 28364 7656 28416
rect 7708 28404 7714 28416
rect 9861 28407 9919 28413
rect 9861 28404 9873 28407
rect 7708 28376 9873 28404
rect 7708 28364 7714 28376
rect 9861 28373 9873 28376
rect 9907 28404 9919 28407
rect 13354 28404 13360 28416
rect 9907 28376 13360 28404
rect 9907 28373 9919 28376
rect 9861 28367 9919 28373
rect 13354 28364 13360 28376
rect 13412 28364 13418 28416
rect 13722 28364 13728 28416
rect 13780 28404 13786 28416
rect 14461 28407 14519 28413
rect 14461 28404 14473 28407
rect 13780 28376 14473 28404
rect 13780 28364 13786 28376
rect 14461 28373 14473 28376
rect 14507 28373 14519 28407
rect 14461 28367 14519 28373
rect 14642 28364 14648 28416
rect 14700 28404 14706 28416
rect 19536 28404 19564 28571
rect 19996 28540 20024 28571
rect 20162 28540 20168 28552
rect 19996 28512 20168 28540
rect 20162 28500 20168 28512
rect 20220 28540 20226 28552
rect 20990 28540 20996 28552
rect 20220 28512 20996 28540
rect 20220 28500 20226 28512
rect 20990 28500 20996 28512
rect 21048 28500 21054 28552
rect 21100 28540 21128 28580
rect 21358 28568 21364 28620
rect 21416 28608 21422 28620
rect 21637 28611 21695 28617
rect 21637 28608 21649 28611
rect 21416 28580 21649 28608
rect 21416 28568 21422 28580
rect 21637 28577 21649 28580
rect 21683 28577 21695 28611
rect 21637 28571 21695 28577
rect 22094 28568 22100 28620
rect 22152 28608 22158 28620
rect 22649 28611 22707 28617
rect 22152 28580 22197 28608
rect 22152 28568 22158 28580
rect 22649 28577 22661 28611
rect 22695 28577 22707 28611
rect 22830 28608 22836 28620
rect 22791 28580 22836 28608
rect 22649 28571 22707 28577
rect 21818 28540 21824 28552
rect 21100 28512 21824 28540
rect 21818 28500 21824 28512
rect 21876 28500 21882 28552
rect 22664 28540 22692 28571
rect 22830 28568 22836 28580
rect 22888 28568 22894 28620
rect 23474 28608 23480 28620
rect 23435 28580 23480 28608
rect 23474 28568 23480 28580
rect 23532 28568 23538 28620
rect 23750 28568 23756 28620
rect 23808 28608 23814 28620
rect 24489 28611 24547 28617
rect 24489 28608 24501 28611
rect 23808 28580 24501 28608
rect 23808 28568 23814 28580
rect 24489 28577 24501 28580
rect 24535 28577 24547 28611
rect 24489 28571 24547 28577
rect 24578 28568 24584 28620
rect 24636 28608 24642 28620
rect 24857 28611 24915 28617
rect 24857 28608 24869 28611
rect 24636 28580 24869 28608
rect 24636 28568 24642 28580
rect 24857 28577 24869 28580
rect 24903 28577 24915 28611
rect 24857 28571 24915 28577
rect 24946 28568 24952 28620
rect 25004 28608 25010 28620
rect 25004 28580 25049 28608
rect 25004 28568 25010 28580
rect 22922 28540 22928 28552
rect 22664 28512 22928 28540
rect 22922 28500 22928 28512
rect 22980 28540 22986 28552
rect 24394 28540 24400 28552
rect 22980 28512 23428 28540
rect 22980 28500 22986 28512
rect 20714 28432 20720 28484
rect 20772 28472 20778 28484
rect 21729 28475 21787 28481
rect 21729 28472 21741 28475
rect 20772 28444 21741 28472
rect 20772 28432 20778 28444
rect 21729 28441 21741 28444
rect 21775 28441 21787 28475
rect 23400 28472 23428 28512
rect 23676 28512 24400 28540
rect 23676 28472 23704 28512
rect 24394 28500 24400 28512
rect 24452 28500 24458 28552
rect 25608 28540 25636 28648
rect 25700 28617 25728 28716
rect 26510 28704 26516 28716
rect 26568 28704 26574 28756
rect 28994 28704 29000 28756
rect 29052 28744 29058 28756
rect 29917 28747 29975 28753
rect 29917 28744 29929 28747
rect 29052 28716 29929 28744
rect 29052 28704 29058 28716
rect 29917 28713 29929 28716
rect 29963 28713 29975 28747
rect 29917 28707 29975 28713
rect 27614 28636 27620 28688
rect 27672 28676 27678 28688
rect 27672 28648 28856 28676
rect 27672 28636 27678 28648
rect 25685 28611 25743 28617
rect 25685 28577 25697 28611
rect 25731 28577 25743 28611
rect 25685 28571 25743 28577
rect 26326 28568 26332 28620
rect 26384 28608 26390 28620
rect 26881 28611 26939 28617
rect 26881 28608 26893 28611
rect 26384 28580 26893 28608
rect 26384 28568 26390 28580
rect 26881 28577 26893 28580
rect 26927 28577 26939 28611
rect 26881 28571 26939 28577
rect 27433 28611 27491 28617
rect 27433 28577 27445 28611
rect 27479 28608 27491 28611
rect 27706 28608 27712 28620
rect 27479 28580 27712 28608
rect 27479 28577 27491 28580
rect 27433 28571 27491 28577
rect 27706 28568 27712 28580
rect 27764 28568 27770 28620
rect 28258 28608 28264 28620
rect 28219 28580 28264 28608
rect 28258 28568 28264 28580
rect 28316 28568 28322 28620
rect 28828 28617 28856 28648
rect 29086 28636 29092 28688
rect 29144 28676 29150 28688
rect 31481 28679 31539 28685
rect 31481 28676 31493 28679
rect 29144 28648 31493 28676
rect 29144 28636 29150 28648
rect 29288 28617 29316 28648
rect 31481 28645 31493 28648
rect 31527 28645 31539 28679
rect 31481 28639 31539 28645
rect 32122 28636 32128 28688
rect 32180 28636 32186 28688
rect 34422 28636 34428 28688
rect 34480 28676 34486 28688
rect 36354 28676 36360 28688
rect 34480 28648 36216 28676
rect 36315 28648 36360 28676
rect 34480 28636 34486 28648
rect 28813 28611 28871 28617
rect 28813 28577 28825 28611
rect 28859 28577 28871 28611
rect 28813 28571 28871 28577
rect 29273 28611 29331 28617
rect 29273 28577 29285 28611
rect 29319 28577 29331 28611
rect 29273 28571 29331 28577
rect 30101 28611 30159 28617
rect 30101 28577 30113 28611
rect 30147 28608 30159 28611
rect 30282 28608 30288 28620
rect 30147 28580 30288 28608
rect 30147 28577 30159 28580
rect 30101 28571 30159 28577
rect 30282 28568 30288 28580
rect 30340 28568 30346 28620
rect 30377 28611 30435 28617
rect 30377 28577 30389 28611
rect 30423 28577 30435 28611
rect 30377 28571 30435 28577
rect 26234 28540 26240 28552
rect 25608 28512 26240 28540
rect 26234 28500 26240 28512
rect 26292 28500 26298 28552
rect 26602 28540 26608 28552
rect 26563 28512 26608 28540
rect 26602 28500 26608 28512
rect 26660 28500 26666 28552
rect 26694 28500 26700 28552
rect 26752 28540 26758 28552
rect 27341 28543 27399 28549
rect 27341 28540 27353 28543
rect 26752 28512 27353 28540
rect 26752 28500 26758 28512
rect 27341 28509 27353 28512
rect 27387 28509 27399 28543
rect 30392 28540 30420 28571
rect 30466 28568 30472 28620
rect 30524 28608 30530 28620
rect 30653 28611 30711 28617
rect 30653 28608 30665 28611
rect 30524 28580 30665 28608
rect 30524 28568 30530 28580
rect 30653 28577 30665 28580
rect 30699 28577 30711 28611
rect 31386 28608 31392 28620
rect 31347 28580 31392 28608
rect 30653 28571 30711 28577
rect 31386 28568 31392 28580
rect 31444 28568 31450 28620
rect 32140 28608 32168 28636
rect 32217 28611 32275 28617
rect 32217 28608 32229 28611
rect 32140 28580 32229 28608
rect 32217 28577 32229 28580
rect 32263 28577 32275 28611
rect 32217 28571 32275 28577
rect 33042 28568 33048 28620
rect 33100 28608 33106 28620
rect 33137 28611 33195 28617
rect 33137 28608 33149 28611
rect 33100 28580 33149 28608
rect 33100 28568 33106 28580
rect 33137 28577 33149 28580
rect 33183 28577 33195 28611
rect 34790 28608 34796 28620
rect 33137 28571 33195 28577
rect 33244 28580 34796 28608
rect 27341 28503 27399 28509
rect 30116 28512 30420 28540
rect 32125 28543 32183 28549
rect 23400 28444 23704 28472
rect 28537 28475 28595 28481
rect 21729 28435 21787 28441
rect 28537 28441 28549 28475
rect 28583 28472 28595 28475
rect 30006 28472 30012 28484
rect 28583 28444 30012 28472
rect 28583 28441 28595 28444
rect 28537 28435 28595 28441
rect 30006 28432 30012 28444
rect 30064 28432 30070 28484
rect 14700 28376 19564 28404
rect 14700 28364 14706 28376
rect 19610 28364 19616 28416
rect 19668 28404 19674 28416
rect 20165 28407 20223 28413
rect 20165 28404 20177 28407
rect 19668 28376 20177 28404
rect 19668 28364 19674 28376
rect 20165 28373 20177 28376
rect 20211 28373 20223 28407
rect 20165 28367 20223 28373
rect 21085 28407 21143 28413
rect 21085 28373 21097 28407
rect 21131 28404 21143 28407
rect 22370 28404 22376 28416
rect 21131 28376 22376 28404
rect 21131 28373 21143 28376
rect 21085 28367 21143 28373
rect 22370 28364 22376 28376
rect 22428 28364 22434 28416
rect 22830 28364 22836 28416
rect 22888 28404 22894 28416
rect 24118 28404 24124 28416
rect 22888 28376 24124 28404
rect 22888 28364 22894 28376
rect 24118 28364 24124 28376
rect 24176 28404 24182 28416
rect 24762 28404 24768 28416
rect 24176 28376 24768 28404
rect 24176 28364 24182 28376
rect 24762 28364 24768 28376
rect 24820 28364 24826 28416
rect 25869 28407 25927 28413
rect 25869 28373 25881 28407
rect 25915 28404 25927 28407
rect 26602 28404 26608 28416
rect 25915 28376 26608 28404
rect 25915 28373 25927 28376
rect 25869 28367 25927 28373
rect 26602 28364 26608 28376
rect 26660 28404 26666 28416
rect 27430 28404 27436 28416
rect 26660 28376 27436 28404
rect 26660 28364 26666 28376
rect 27430 28364 27436 28376
rect 27488 28364 27494 28416
rect 27522 28364 27528 28416
rect 27580 28404 27586 28416
rect 29086 28404 29092 28416
rect 27580 28376 29092 28404
rect 27580 28364 27586 28376
rect 29086 28364 29092 28376
rect 29144 28404 29150 28416
rect 30116 28404 30144 28512
rect 32125 28509 32137 28543
rect 32171 28540 32183 28543
rect 33244 28540 33272 28580
rect 34790 28568 34796 28580
rect 34848 28568 34854 28620
rect 35710 28608 35716 28620
rect 35671 28580 35716 28608
rect 35710 28568 35716 28580
rect 35768 28568 35774 28620
rect 35802 28568 35808 28620
rect 35860 28608 35866 28620
rect 36081 28611 36139 28617
rect 36081 28608 36093 28611
rect 35860 28580 36093 28608
rect 35860 28568 35866 28580
rect 36081 28577 36093 28580
rect 36127 28577 36139 28611
rect 36188 28608 36216 28648
rect 36354 28636 36360 28648
rect 36412 28636 36418 28688
rect 36817 28611 36875 28617
rect 36817 28608 36829 28611
rect 36188 28580 36829 28608
rect 36081 28571 36139 28577
rect 36817 28577 36829 28580
rect 36863 28577 36875 28611
rect 38102 28608 38108 28620
rect 38063 28580 38108 28608
rect 36817 28571 36875 28577
rect 38102 28568 38108 28580
rect 38160 28568 38166 28620
rect 38286 28608 38292 28620
rect 38247 28580 38292 28608
rect 38286 28568 38292 28580
rect 38344 28568 38350 28620
rect 38378 28568 38384 28620
rect 38436 28608 38442 28620
rect 38749 28611 38807 28617
rect 38749 28608 38761 28611
rect 38436 28580 38761 28608
rect 38436 28568 38442 28580
rect 38749 28577 38761 28580
rect 38795 28577 38807 28611
rect 38749 28571 38807 28577
rect 33410 28540 33416 28552
rect 32171 28512 33272 28540
rect 33371 28512 33416 28540
rect 32171 28509 32183 28512
rect 32125 28503 32183 28509
rect 33410 28500 33416 28512
rect 33468 28500 33474 28552
rect 35345 28543 35403 28549
rect 35345 28540 35357 28543
rect 34532 28512 35357 28540
rect 34532 28416 34560 28512
rect 35345 28509 35357 28512
rect 35391 28509 35403 28543
rect 35345 28503 35403 28509
rect 38654 28432 38660 28484
rect 38712 28472 38718 28484
rect 38749 28475 38807 28481
rect 38749 28472 38761 28475
rect 38712 28444 38761 28472
rect 38712 28432 38718 28444
rect 38749 28441 38761 28444
rect 38795 28441 38807 28475
rect 38749 28435 38807 28441
rect 32398 28404 32404 28416
rect 29144 28376 30144 28404
rect 32359 28376 32404 28404
rect 29144 28364 29150 28376
rect 32398 28364 32404 28376
rect 32456 28364 32462 28416
rect 34514 28404 34520 28416
rect 34475 28376 34520 28404
rect 34514 28364 34520 28376
rect 34572 28364 34578 28416
rect 35710 28364 35716 28416
rect 35768 28404 35774 28416
rect 37001 28407 37059 28413
rect 37001 28404 37013 28407
rect 35768 28376 37013 28404
rect 35768 28364 35774 28376
rect 37001 28373 37013 28376
rect 37047 28373 37059 28407
rect 37001 28367 37059 28373
rect 1104 28314 39836 28336
rect 1104 28262 4246 28314
rect 4298 28262 4310 28314
rect 4362 28262 4374 28314
rect 4426 28262 4438 28314
rect 4490 28262 34966 28314
rect 35018 28262 35030 28314
rect 35082 28262 35094 28314
rect 35146 28262 35158 28314
rect 35210 28262 39836 28314
rect 1104 28240 39836 28262
rect 1673 28203 1731 28209
rect 1673 28169 1685 28203
rect 1719 28200 1731 28203
rect 2958 28200 2964 28212
rect 1719 28172 2964 28200
rect 1719 28169 1731 28172
rect 1673 28163 1731 28169
rect 2958 28160 2964 28172
rect 3016 28160 3022 28212
rect 3068 28172 4384 28200
rect 2317 28135 2375 28141
rect 2317 28101 2329 28135
rect 2363 28132 2375 28135
rect 2774 28132 2780 28144
rect 2363 28104 2780 28132
rect 2363 28101 2375 28104
rect 2317 28095 2375 28101
rect 2774 28092 2780 28104
rect 2832 28092 2838 28144
rect 2866 28064 2872 28076
rect 2240 28036 2872 28064
rect 2240 28005 2268 28036
rect 2866 28024 2872 28036
rect 2924 28024 2930 28076
rect 3068 28005 3096 28172
rect 4356 28132 4384 28172
rect 7834 28160 7840 28212
rect 7892 28200 7898 28212
rect 8021 28203 8079 28209
rect 8021 28200 8033 28203
rect 7892 28172 8033 28200
rect 7892 28160 7898 28172
rect 8021 28169 8033 28172
rect 8067 28169 8079 28203
rect 8021 28163 8079 28169
rect 4430 28132 4436 28144
rect 4356 28104 4436 28132
rect 4430 28092 4436 28104
rect 4488 28132 4494 28144
rect 4614 28132 4620 28144
rect 4488 28104 4620 28132
rect 4488 28092 4494 28104
rect 4614 28092 4620 28104
rect 4672 28092 4678 28144
rect 5258 28132 5264 28144
rect 5219 28104 5264 28132
rect 5258 28092 5264 28104
rect 5316 28092 5322 28144
rect 6181 28135 6239 28141
rect 6181 28101 6193 28135
rect 6227 28101 6239 28135
rect 6914 28132 6920 28144
rect 6875 28104 6920 28132
rect 6181 28095 6239 28101
rect 6196 28064 6224 28095
rect 6914 28092 6920 28104
rect 6972 28092 6978 28144
rect 3436 28036 6224 28064
rect 3436 28008 3464 28036
rect 5000 28008 5028 28036
rect 1581 27999 1639 28005
rect 1581 27996 1593 27999
rect 1504 27968 1593 27996
rect 1504 27860 1532 27968
rect 1581 27965 1593 27968
rect 1627 27965 1639 27999
rect 1581 27959 1639 27965
rect 2225 27999 2283 28005
rect 2225 27965 2237 27999
rect 2271 27965 2283 27999
rect 2225 27959 2283 27965
rect 3053 27999 3111 28005
rect 3053 27965 3065 27999
rect 3099 27965 3111 27999
rect 3418 27996 3424 28008
rect 3331 27968 3424 27996
rect 3053 27959 3111 27965
rect 3418 27956 3424 27968
rect 3476 27956 3482 28008
rect 3789 27999 3847 28005
rect 3789 27965 3801 27999
rect 3835 27996 3847 27999
rect 4430 27996 4436 28008
rect 3835 27968 4292 27996
rect 4391 27968 4436 27996
rect 3835 27965 3847 27968
rect 3789 27959 3847 27965
rect 3973 27931 4031 27937
rect 3973 27897 3985 27931
rect 4019 27928 4031 27931
rect 4062 27928 4068 27940
rect 4019 27900 4068 27928
rect 4019 27897 4031 27900
rect 3973 27891 4031 27897
rect 4062 27888 4068 27900
rect 4120 27888 4126 27940
rect 4264 27928 4292 27968
rect 4430 27956 4436 27968
rect 4488 27956 4494 28008
rect 4982 27996 4988 28008
rect 4895 27968 4988 27996
rect 4982 27956 4988 27968
rect 5040 27956 5046 28008
rect 5353 27999 5411 28005
rect 5353 27965 5365 27999
rect 5399 27996 5411 27999
rect 5442 27996 5448 28008
rect 5399 27968 5448 27996
rect 5399 27965 5411 27968
rect 5353 27959 5411 27965
rect 5442 27956 5448 27968
rect 5500 27956 5506 28008
rect 5626 27956 5632 28008
rect 5684 27996 5690 28008
rect 5997 27999 6055 28005
rect 5997 27996 6009 27999
rect 5684 27968 6009 27996
rect 5684 27956 5690 27968
rect 5997 27965 6009 27968
rect 6043 27965 6055 27999
rect 5997 27959 6055 27965
rect 7101 27999 7159 28005
rect 7101 27965 7113 27999
rect 7147 27996 7159 27999
rect 7190 27996 7196 28008
rect 7147 27968 7196 27996
rect 7147 27965 7159 27968
rect 7101 27959 7159 27965
rect 7190 27956 7196 27968
rect 7248 27956 7254 28008
rect 7374 27996 7380 28008
rect 7335 27968 7380 27996
rect 7374 27956 7380 27968
rect 7432 27956 7438 28008
rect 6638 27928 6644 27940
rect 4264 27900 6644 27928
rect 6638 27888 6644 27900
rect 6696 27888 6702 27940
rect 8036 27928 8064 28163
rect 8754 28160 8760 28212
rect 8812 28200 8818 28212
rect 9217 28203 9275 28209
rect 9217 28200 9229 28203
rect 8812 28172 9229 28200
rect 8812 28160 8818 28172
rect 9217 28169 9229 28172
rect 9263 28169 9275 28203
rect 9217 28163 9275 28169
rect 10502 28160 10508 28212
rect 10560 28200 10566 28212
rect 10962 28200 10968 28212
rect 10560 28172 10968 28200
rect 10560 28160 10566 28172
rect 10962 28160 10968 28172
rect 11020 28200 11026 28212
rect 11333 28203 11391 28209
rect 11333 28200 11345 28203
rect 11020 28172 11345 28200
rect 11020 28160 11026 28172
rect 11333 28169 11345 28172
rect 11379 28169 11391 28203
rect 12618 28200 12624 28212
rect 12579 28172 12624 28200
rect 11333 28163 11391 28169
rect 12618 28160 12624 28172
rect 12676 28160 12682 28212
rect 15194 28200 15200 28212
rect 13648 28172 14964 28200
rect 15155 28172 15200 28200
rect 13648 28132 13676 28172
rect 14936 28144 14964 28172
rect 15194 28160 15200 28172
rect 15252 28160 15258 28212
rect 20622 28200 20628 28212
rect 15304 28172 20628 28200
rect 13814 28132 13820 28144
rect 8220 28104 13676 28132
rect 13775 28104 13820 28132
rect 8220 28005 8248 28104
rect 13814 28092 13820 28104
rect 13872 28092 13878 28144
rect 14918 28092 14924 28144
rect 14976 28132 14982 28144
rect 15304 28132 15332 28172
rect 20622 28160 20628 28172
rect 20680 28160 20686 28212
rect 21726 28160 21732 28212
rect 21784 28200 21790 28212
rect 22278 28200 22284 28212
rect 21784 28172 22284 28200
rect 21784 28160 21790 28172
rect 22278 28160 22284 28172
rect 22336 28160 22342 28212
rect 25498 28200 25504 28212
rect 23952 28172 25504 28200
rect 19702 28132 19708 28144
rect 14976 28104 15332 28132
rect 18708 28104 19708 28132
rect 14976 28092 14982 28104
rect 9950 28024 9956 28076
rect 10008 28064 10014 28076
rect 10689 28067 10747 28073
rect 10689 28064 10701 28067
rect 10008 28036 10701 28064
rect 10008 28024 10014 28036
rect 10689 28033 10701 28036
rect 10735 28033 10747 28067
rect 10689 28027 10747 28033
rect 10962 28024 10968 28076
rect 11020 28064 11026 28076
rect 14553 28067 14611 28073
rect 11020 28036 13584 28064
rect 11020 28024 11026 28036
rect 8205 27999 8263 28005
rect 8205 27965 8217 27999
rect 8251 27965 8263 27999
rect 8205 27959 8263 27965
rect 8294 27956 8300 28008
rect 8352 27996 8358 28008
rect 9033 27999 9091 28005
rect 8352 27968 8397 27996
rect 8352 27956 8358 27968
rect 9033 27965 9045 27999
rect 9079 27996 9091 27999
rect 9122 27996 9128 28008
rect 9079 27968 9128 27996
rect 9079 27965 9091 27968
rect 9033 27959 9091 27965
rect 9122 27956 9128 27968
rect 9180 27956 9186 28008
rect 9861 27999 9919 28005
rect 9861 27965 9873 27999
rect 9907 27996 9919 27999
rect 10042 27996 10048 28008
rect 9907 27968 10048 27996
rect 9907 27965 9919 27968
rect 9861 27959 9919 27965
rect 10042 27956 10048 27968
rect 10100 27956 10106 28008
rect 10226 27996 10232 28008
rect 10187 27968 10232 27996
rect 10226 27956 10232 27968
rect 10284 27956 10290 28008
rect 10597 27999 10655 28005
rect 10597 27965 10609 27999
rect 10643 27996 10655 27999
rect 11422 27996 11428 28008
rect 10643 27968 11428 27996
rect 10643 27965 10655 27968
rect 10597 27959 10655 27965
rect 11422 27956 11428 27968
rect 11480 27956 11486 28008
rect 11517 27999 11575 28005
rect 11517 27965 11529 27999
rect 11563 27965 11575 27999
rect 11517 27959 11575 27965
rect 11701 27999 11759 28005
rect 11701 27965 11713 27999
rect 11747 27965 11759 27999
rect 11701 27959 11759 27965
rect 12437 27999 12495 28005
rect 12437 27965 12449 27999
rect 12483 27996 12495 27999
rect 12802 27996 12808 28008
rect 12483 27968 12808 27996
rect 12483 27965 12495 27968
rect 12437 27959 12495 27965
rect 11532 27928 11560 27959
rect 8036 27900 11560 27928
rect 11716 27928 11744 27959
rect 12802 27956 12808 27968
rect 12860 27956 12866 28008
rect 13556 28005 13584 28036
rect 14553 28033 14565 28067
rect 14599 28064 14611 28067
rect 16666 28064 16672 28076
rect 14599 28036 16436 28064
rect 16627 28036 16672 28064
rect 14599 28033 14611 28036
rect 14553 28027 14611 28033
rect 13541 27999 13599 28005
rect 13541 27965 13553 27999
rect 13587 27965 13599 27999
rect 13541 27959 13599 27965
rect 14277 27999 14335 28005
rect 14277 27965 14289 27999
rect 14323 27965 14335 27999
rect 14277 27959 14335 27965
rect 13170 27928 13176 27940
rect 11716 27900 13176 27928
rect 13170 27888 13176 27900
rect 13228 27888 13234 27940
rect 14292 27928 14320 27959
rect 14458 27956 14464 28008
rect 14516 27996 14522 28008
rect 15105 27999 15163 28005
rect 15105 27996 15117 27999
rect 14516 27968 15117 27996
rect 14516 27956 14522 27968
rect 15105 27965 15117 27968
rect 15151 27965 15163 27999
rect 15838 27996 15844 28008
rect 15799 27968 15844 27996
rect 15105 27959 15163 27965
rect 15838 27956 15844 27968
rect 15896 27956 15902 28008
rect 15378 27928 15384 27940
rect 14292 27900 15384 27928
rect 15378 27888 15384 27900
rect 15436 27888 15442 27940
rect 16408 27928 16436 28036
rect 16666 28024 16672 28036
rect 16724 28024 16730 28076
rect 18230 28024 18236 28076
rect 18288 28064 18294 28076
rect 18708 28073 18736 28104
rect 19702 28092 19708 28104
rect 19760 28092 19766 28144
rect 18693 28067 18751 28073
rect 18288 28036 18552 28064
rect 18288 28024 18294 28036
rect 16485 27999 16543 28005
rect 16485 27965 16497 27999
rect 16531 27996 16543 27999
rect 17862 27996 17868 28008
rect 16531 27968 17868 27996
rect 16531 27965 16543 27968
rect 16485 27959 16543 27965
rect 17862 27956 17868 27968
rect 17920 27956 17926 28008
rect 18322 27996 18328 28008
rect 18283 27968 18328 27996
rect 18322 27956 18328 27968
rect 18380 27956 18386 28008
rect 18524 28005 18552 28036
rect 18693 28033 18705 28067
rect 18739 28033 18751 28067
rect 18693 28027 18751 28033
rect 19426 28024 19432 28076
rect 19484 28064 19490 28076
rect 20625 28067 20683 28073
rect 20625 28064 20637 28067
rect 19484 28036 20637 28064
rect 19484 28024 19490 28036
rect 20625 28033 20637 28036
rect 20671 28033 20683 28067
rect 21542 28064 21548 28076
rect 20625 28027 20683 28033
rect 21192 28036 21548 28064
rect 18509 27999 18567 28005
rect 18509 27965 18521 27999
rect 18555 27965 18567 27999
rect 19150 27996 19156 28008
rect 19111 27968 19156 27996
rect 18509 27959 18567 27965
rect 19150 27956 19156 27968
rect 19208 27956 19214 28008
rect 19334 27956 19340 28008
rect 19392 27996 19398 28008
rect 19610 27996 19616 28008
rect 19392 27968 19616 27996
rect 19392 27956 19398 27968
rect 19610 27956 19616 27968
rect 19668 27956 19674 28008
rect 19705 27999 19763 28005
rect 19705 27965 19717 27999
rect 19751 27965 19763 27999
rect 19705 27959 19763 27965
rect 20533 27999 20591 28005
rect 20533 27965 20545 27999
rect 20579 27996 20591 27999
rect 20806 27996 20812 28008
rect 20579 27968 20812 27996
rect 20579 27965 20591 27968
rect 20533 27959 20591 27965
rect 17586 27928 17592 27940
rect 16408 27900 17592 27928
rect 17586 27888 17592 27900
rect 17644 27928 17650 27940
rect 19720 27928 19748 27959
rect 20806 27956 20812 27968
rect 20864 27956 20870 28008
rect 21192 28005 21220 28036
rect 21542 28024 21548 28036
rect 21600 28024 21606 28076
rect 21177 27999 21235 28005
rect 21177 27965 21189 27999
rect 21223 27965 21235 27999
rect 21358 27996 21364 28008
rect 21319 27968 21364 27996
rect 21177 27959 21235 27965
rect 21358 27956 21364 27968
rect 21416 27956 21422 28008
rect 21910 27996 21916 28008
rect 21871 27968 21916 27996
rect 21910 27956 21916 27968
rect 21968 27956 21974 28008
rect 22278 27996 22284 28008
rect 22239 27968 22284 27996
rect 22278 27956 22284 27968
rect 22336 27956 22342 28008
rect 23952 28005 23980 28172
rect 25498 28160 25504 28172
rect 25556 28160 25562 28212
rect 29546 28200 29552 28212
rect 29507 28172 29552 28200
rect 29546 28160 29552 28172
rect 29604 28160 29610 28212
rect 30006 28160 30012 28212
rect 30064 28200 30070 28212
rect 30064 28172 32812 28200
rect 30064 28160 30070 28172
rect 24118 28132 24124 28144
rect 24079 28104 24124 28132
rect 24118 28092 24124 28104
rect 24176 28092 24182 28144
rect 28629 28135 28687 28141
rect 28629 28101 28641 28135
rect 28675 28101 28687 28135
rect 28629 28095 28687 28101
rect 24026 28024 24032 28076
rect 24084 28064 24090 28076
rect 24302 28064 24308 28076
rect 24084 28036 24308 28064
rect 24084 28024 24090 28036
rect 24302 28024 24308 28036
rect 24360 28064 24366 28076
rect 27798 28064 27804 28076
rect 24360 28036 24716 28064
rect 24360 28024 24366 28036
rect 24688 28005 24716 28036
rect 25792 28036 27384 28064
rect 27759 28036 27804 28064
rect 25792 28008 25820 28036
rect 22925 27999 22983 28005
rect 22925 27965 22937 27999
rect 22971 27965 22983 27999
rect 22925 27959 22983 27965
rect 23937 27999 23995 28005
rect 23937 27965 23949 27999
rect 23983 27965 23995 27999
rect 23937 27959 23995 27965
rect 24679 27999 24737 28005
rect 24679 27965 24691 27999
rect 24725 27965 24737 27999
rect 25406 27996 25412 28008
rect 25367 27968 25412 27996
rect 24679 27959 24737 27965
rect 17644 27900 19748 27928
rect 21376 27928 21404 27956
rect 21726 27928 21732 27940
rect 21376 27900 21732 27928
rect 17644 27888 17650 27900
rect 21726 27888 21732 27900
rect 21784 27888 21790 27940
rect 2590 27860 2596 27872
rect 1504 27832 2596 27860
rect 2590 27820 2596 27832
rect 2648 27820 2654 27872
rect 8481 27863 8539 27869
rect 8481 27829 8493 27863
rect 8527 27860 8539 27863
rect 9858 27860 9864 27872
rect 8527 27832 9864 27860
rect 8527 27829 8539 27832
rect 8481 27823 8539 27829
rect 9858 27820 9864 27832
rect 9916 27860 9922 27872
rect 10778 27860 10784 27872
rect 9916 27832 10784 27860
rect 9916 27820 9922 27832
rect 10778 27820 10784 27832
rect 10836 27820 10842 27872
rect 11793 27863 11851 27869
rect 11793 27829 11805 27863
rect 11839 27860 11851 27863
rect 12066 27860 12072 27872
rect 11839 27832 12072 27860
rect 11839 27829 11851 27832
rect 11793 27823 11851 27829
rect 12066 27820 12072 27832
rect 12124 27820 12130 27872
rect 15930 27860 15936 27872
rect 15891 27832 15936 27860
rect 15930 27820 15936 27832
rect 15988 27820 15994 27872
rect 21634 27820 21640 27872
rect 21692 27860 21698 27872
rect 22738 27860 22744 27872
rect 21692 27832 22744 27860
rect 21692 27820 21698 27832
rect 22738 27820 22744 27832
rect 22796 27820 22802 27872
rect 22940 27860 22968 27959
rect 25406 27956 25412 27968
rect 25464 27996 25470 28008
rect 25774 27996 25780 28008
rect 25464 27968 25780 27996
rect 25464 27956 25470 27968
rect 25774 27956 25780 27968
rect 25832 27956 25838 28008
rect 25958 27996 25964 28008
rect 25919 27968 25964 27996
rect 25958 27956 25964 27968
rect 26016 27956 26022 28008
rect 26418 27996 26424 28008
rect 26331 27968 26424 27996
rect 26418 27956 26424 27968
rect 26476 27996 26482 28008
rect 26878 27996 26884 28008
rect 26476 27968 26884 27996
rect 26476 27956 26482 27968
rect 26878 27956 26884 27968
rect 26936 27956 26942 28008
rect 27356 28005 27384 28036
rect 27798 28024 27804 28036
rect 27856 28024 27862 28076
rect 28644 28064 28672 28095
rect 29178 28092 29184 28144
rect 29236 28132 29242 28144
rect 29236 28104 30328 28132
rect 29236 28092 29242 28104
rect 30024 28076 30052 28104
rect 29270 28064 29276 28076
rect 28644 28036 29276 28064
rect 29270 28024 29276 28036
rect 29328 28024 29334 28076
rect 30006 28024 30012 28076
rect 30064 28024 30070 28076
rect 30300 28073 30328 28104
rect 30285 28067 30343 28073
rect 30285 28033 30297 28067
rect 30331 28033 30343 28067
rect 30285 28027 30343 28033
rect 30561 28067 30619 28073
rect 30561 28033 30573 28067
rect 30607 28064 30619 28067
rect 32398 28064 32404 28076
rect 30607 28036 32404 28064
rect 30607 28033 30619 28036
rect 30561 28027 30619 28033
rect 32398 28024 32404 28036
rect 32456 28024 32462 28076
rect 27341 27999 27399 28005
rect 27341 27965 27353 27999
rect 27387 27965 27399 27999
rect 27341 27959 27399 27965
rect 28445 27999 28503 28005
rect 28445 27965 28457 27999
rect 28491 27965 28503 27999
rect 28445 27959 28503 27965
rect 23017 27931 23075 27937
rect 23017 27897 23029 27931
rect 23063 27928 23075 27931
rect 24762 27928 24768 27940
rect 23063 27900 24768 27928
rect 23063 27897 23075 27900
rect 23017 27891 23075 27897
rect 24762 27888 24768 27900
rect 24820 27888 24826 27940
rect 26510 27888 26516 27940
rect 26568 27928 26574 27940
rect 27062 27928 27068 27940
rect 26568 27900 27068 27928
rect 26568 27888 26574 27900
rect 27062 27888 27068 27900
rect 27120 27888 27126 27940
rect 27433 27931 27491 27937
rect 27433 27897 27445 27931
rect 27479 27928 27491 27931
rect 27522 27928 27528 27940
rect 27479 27900 27528 27928
rect 27479 27897 27491 27900
rect 27433 27891 27491 27897
rect 27522 27888 27528 27900
rect 27580 27888 27586 27940
rect 28460 27928 28488 27959
rect 29362 27956 29368 28008
rect 29420 27996 29426 28008
rect 32784 28005 32812 28172
rect 33502 28160 33508 28212
rect 33560 28200 33566 28212
rect 34149 28203 34207 28209
rect 34149 28200 34161 28203
rect 33560 28172 34161 28200
rect 33560 28160 33566 28172
rect 34149 28169 34161 28172
rect 34195 28169 34207 28203
rect 34149 28163 34207 28169
rect 36725 28203 36783 28209
rect 36725 28169 36737 28203
rect 36771 28200 36783 28203
rect 37734 28200 37740 28212
rect 36771 28172 37740 28200
rect 36771 28169 36783 28172
rect 36725 28163 36783 28169
rect 37734 28160 37740 28172
rect 37792 28160 37798 28212
rect 33410 28064 33416 28076
rect 33371 28036 33416 28064
rect 33410 28024 33416 28036
rect 33468 28024 33474 28076
rect 35161 28067 35219 28073
rect 35161 28033 35173 28067
rect 35207 28064 35219 28067
rect 37550 28064 37556 28076
rect 35207 28036 37320 28064
rect 37511 28036 37556 28064
rect 35207 28033 35219 28036
rect 35161 28027 35219 28033
rect 37292 28008 37320 28036
rect 37550 28024 37556 28036
rect 37608 28024 37614 28076
rect 32585 27999 32643 28005
rect 29420 27968 29465 27996
rect 30392 27968 32536 27996
rect 29420 27956 29426 27968
rect 30392 27928 30420 27968
rect 28460 27900 30420 27928
rect 24026 27860 24032 27872
rect 22940 27832 24032 27860
rect 24026 27820 24032 27832
rect 24084 27820 24090 27872
rect 24857 27863 24915 27869
rect 24857 27829 24869 27863
rect 24903 27860 24915 27863
rect 25682 27860 25688 27872
rect 24903 27832 25688 27860
rect 24903 27829 24915 27832
rect 24857 27823 24915 27829
rect 25682 27820 25688 27832
rect 25740 27820 25746 27872
rect 25866 27820 25872 27872
rect 25924 27860 25930 27872
rect 27249 27863 27307 27869
rect 27249 27860 27261 27863
rect 25924 27832 27261 27860
rect 25924 27820 25930 27832
rect 27249 27829 27261 27832
rect 27295 27829 27307 27863
rect 27249 27823 27307 27829
rect 29454 27820 29460 27872
rect 29512 27860 29518 27872
rect 31386 27860 31392 27872
rect 29512 27832 31392 27860
rect 29512 27820 29518 27832
rect 31386 27820 31392 27832
rect 31444 27820 31450 27872
rect 31846 27860 31852 27872
rect 31807 27832 31852 27860
rect 31846 27820 31852 27832
rect 31904 27820 31910 27872
rect 32508 27860 32536 27968
rect 32585 27965 32597 27999
rect 32631 27965 32643 27999
rect 32585 27959 32643 27965
rect 32769 27999 32827 28005
rect 32769 27965 32781 27999
rect 32815 27965 32827 27999
rect 33318 27996 33324 28008
rect 33279 27968 33324 27996
rect 32769 27959 32827 27965
rect 32600 27928 32628 27959
rect 33318 27956 33324 27968
rect 33376 27956 33382 28008
rect 33962 27996 33968 28008
rect 33923 27968 33968 27996
rect 33962 27956 33968 27968
rect 34020 27956 34026 28008
rect 35437 27999 35495 28005
rect 35437 27965 35449 27999
rect 35483 27996 35495 27999
rect 36078 27996 36084 28008
rect 35483 27968 36084 27996
rect 35483 27965 35495 27968
rect 35437 27959 35495 27965
rect 36078 27956 36084 27968
rect 36136 27956 36142 28008
rect 37274 27996 37280 28008
rect 37235 27968 37280 27996
rect 37274 27956 37280 27968
rect 37332 27956 37338 28008
rect 33502 27928 33508 27940
rect 32600 27900 33508 27928
rect 33502 27888 33508 27900
rect 33560 27888 33566 27940
rect 34054 27860 34060 27872
rect 32508 27832 34060 27860
rect 34054 27820 34060 27832
rect 34112 27820 34118 27872
rect 38010 27820 38016 27872
rect 38068 27860 38074 27872
rect 38657 27863 38715 27869
rect 38657 27860 38669 27863
rect 38068 27832 38669 27860
rect 38068 27820 38074 27832
rect 38657 27829 38669 27832
rect 38703 27829 38715 27863
rect 38657 27823 38715 27829
rect 1104 27770 39836 27792
rect 1104 27718 19606 27770
rect 19658 27718 19670 27770
rect 19722 27718 19734 27770
rect 19786 27718 19798 27770
rect 19850 27718 39836 27770
rect 1104 27696 39836 27718
rect 4154 27656 4160 27668
rect 4115 27628 4160 27656
rect 4154 27616 4160 27628
rect 4212 27616 4218 27668
rect 15930 27616 15936 27668
rect 15988 27656 15994 27668
rect 15988 27628 23704 27656
rect 15988 27616 15994 27628
rect 1765 27591 1823 27597
rect 1765 27557 1777 27591
rect 1811 27588 1823 27591
rect 5534 27588 5540 27600
rect 1811 27560 5540 27588
rect 1811 27557 1823 27560
rect 1765 27551 1823 27557
rect 5534 27548 5540 27560
rect 5592 27548 5598 27600
rect 6914 27588 6920 27600
rect 5644 27560 6920 27588
rect 1673 27523 1731 27529
rect 1673 27489 1685 27523
rect 1719 27489 1731 27523
rect 1673 27483 1731 27489
rect 1688 27452 1716 27483
rect 2038 27480 2044 27532
rect 2096 27520 2102 27532
rect 2498 27520 2504 27532
rect 2096 27492 2504 27520
rect 2096 27480 2102 27492
rect 2498 27480 2504 27492
rect 2556 27480 2562 27532
rect 2590 27480 2596 27532
rect 2648 27520 2654 27532
rect 3418 27520 3424 27532
rect 2648 27492 3424 27520
rect 2648 27480 2654 27492
rect 3418 27480 3424 27492
rect 3476 27480 3482 27532
rect 3878 27520 3884 27532
rect 3839 27492 3884 27520
rect 3878 27480 3884 27492
rect 3936 27480 3942 27532
rect 4062 27520 4068 27532
rect 4023 27492 4068 27520
rect 4062 27480 4068 27492
rect 4120 27480 4126 27532
rect 4614 27520 4620 27532
rect 4575 27492 4620 27520
rect 4614 27480 4620 27492
rect 4672 27480 4678 27532
rect 4982 27520 4988 27532
rect 4943 27492 4988 27520
rect 4982 27480 4988 27492
rect 5040 27480 5046 27532
rect 5644 27529 5672 27560
rect 6914 27548 6920 27560
rect 6972 27548 6978 27600
rect 7101 27591 7159 27597
rect 7101 27557 7113 27591
rect 7147 27588 7159 27591
rect 7374 27588 7380 27600
rect 7147 27560 7380 27588
rect 7147 27557 7159 27560
rect 7101 27551 7159 27557
rect 7374 27548 7380 27560
rect 7432 27548 7438 27600
rect 8294 27588 8300 27600
rect 7576 27560 8300 27588
rect 5629 27523 5687 27529
rect 5629 27489 5641 27523
rect 5675 27489 5687 27523
rect 5629 27483 5687 27489
rect 5994 27480 6000 27532
rect 6052 27520 6058 27532
rect 6273 27523 6331 27529
rect 6273 27520 6285 27523
rect 6052 27492 6285 27520
rect 6052 27480 6058 27492
rect 6273 27489 6285 27492
rect 6319 27520 6331 27523
rect 7576 27520 7604 27560
rect 8294 27548 8300 27560
rect 8352 27548 8358 27600
rect 10870 27588 10876 27600
rect 8772 27560 10640 27588
rect 10831 27560 10876 27588
rect 6319 27492 7604 27520
rect 6319 27489 6331 27492
rect 6273 27483 6331 27489
rect 7650 27480 7656 27532
rect 7708 27520 7714 27532
rect 7926 27520 7932 27532
rect 7708 27492 7753 27520
rect 7887 27492 7932 27520
rect 7708 27480 7714 27492
rect 7926 27480 7932 27492
rect 7984 27480 7990 27532
rect 8772 27520 8800 27560
rect 8036 27492 8800 27520
rect 8849 27523 8907 27529
rect 5718 27452 5724 27464
rect 1688 27424 5724 27452
rect 5718 27412 5724 27424
rect 5776 27412 5782 27464
rect 6638 27412 6644 27464
rect 6696 27452 6702 27464
rect 8036 27452 8064 27492
rect 8849 27489 8861 27523
rect 8895 27520 8907 27523
rect 9122 27520 9128 27532
rect 8895 27492 9128 27520
rect 8895 27489 8907 27492
rect 8849 27483 8907 27489
rect 9122 27480 9128 27492
rect 9180 27480 9186 27532
rect 10226 27520 10232 27532
rect 10187 27492 10232 27520
rect 10226 27480 10232 27492
rect 10284 27480 10290 27532
rect 10612 27529 10640 27560
rect 10870 27548 10876 27560
rect 10928 27548 10934 27600
rect 14274 27588 14280 27600
rect 13096 27560 14280 27588
rect 10597 27523 10655 27529
rect 10597 27489 10609 27523
rect 10643 27489 10655 27523
rect 11330 27520 11336 27532
rect 11291 27492 11336 27520
rect 10597 27483 10655 27489
rect 11330 27480 11336 27492
rect 11388 27480 11394 27532
rect 12066 27520 12072 27532
rect 12027 27492 12072 27520
rect 12066 27480 12072 27492
rect 12124 27480 12130 27532
rect 12434 27480 12440 27532
rect 12492 27520 12498 27532
rect 13096 27529 13124 27560
rect 14274 27548 14280 27560
rect 14332 27588 14338 27600
rect 15378 27588 15384 27600
rect 14332 27560 15240 27588
rect 15339 27560 15384 27588
rect 14332 27548 14338 27560
rect 13081 27523 13139 27529
rect 12492 27492 12537 27520
rect 12492 27480 12498 27492
rect 13081 27489 13093 27523
rect 13127 27489 13139 27523
rect 13081 27483 13139 27489
rect 13357 27523 13415 27529
rect 13357 27489 13369 27523
rect 13403 27489 13415 27523
rect 14001 27523 14059 27529
rect 14001 27520 14013 27523
rect 13357 27483 13415 27489
rect 13464 27492 14013 27520
rect 6696 27424 8064 27452
rect 8113 27455 8171 27461
rect 6696 27412 6702 27424
rect 8113 27421 8125 27455
rect 8159 27452 8171 27455
rect 8570 27452 8576 27464
rect 8159 27424 8576 27452
rect 8159 27421 8171 27424
rect 8113 27415 8171 27421
rect 8570 27412 8576 27424
rect 8628 27412 8634 27464
rect 9953 27455 10011 27461
rect 9953 27421 9965 27455
rect 9999 27452 10011 27455
rect 11790 27452 11796 27464
rect 9999 27424 11796 27452
rect 9999 27421 10011 27424
rect 9953 27415 10011 27421
rect 11790 27412 11796 27424
rect 11848 27412 11854 27464
rect 1394 27344 1400 27396
rect 1452 27384 1458 27396
rect 3697 27387 3755 27393
rect 3697 27384 3709 27387
rect 1452 27356 3709 27384
rect 1452 27344 1458 27356
rect 3697 27353 3709 27356
rect 3743 27384 3755 27387
rect 3970 27384 3976 27396
rect 3743 27356 3976 27384
rect 3743 27353 3755 27356
rect 3697 27347 3755 27353
rect 3970 27344 3976 27356
rect 4028 27384 4034 27396
rect 6546 27384 6552 27396
rect 4028 27356 6552 27384
rect 4028 27344 4034 27356
rect 6546 27344 6552 27356
rect 6604 27344 6610 27396
rect 11974 27384 11980 27396
rect 7944 27356 11980 27384
rect 2038 27276 2044 27328
rect 2096 27316 2102 27328
rect 2317 27319 2375 27325
rect 2317 27316 2329 27319
rect 2096 27288 2329 27316
rect 2096 27276 2102 27288
rect 2317 27285 2329 27288
rect 2363 27285 2375 27319
rect 2317 27279 2375 27285
rect 2774 27276 2780 27328
rect 2832 27316 2838 27328
rect 5718 27316 5724 27328
rect 2832 27288 2877 27316
rect 5679 27288 5724 27316
rect 2832 27276 2838 27288
rect 5718 27276 5724 27288
rect 5776 27276 5782 27328
rect 5810 27276 5816 27328
rect 5868 27316 5874 27328
rect 6457 27319 6515 27325
rect 6457 27316 6469 27319
rect 5868 27288 6469 27316
rect 5868 27276 5874 27288
rect 6457 27285 6469 27288
rect 6503 27316 6515 27319
rect 7944 27316 7972 27356
rect 11974 27344 11980 27356
rect 12032 27344 12038 27396
rect 13372 27384 13400 27483
rect 13464 27461 13492 27492
rect 14001 27489 14013 27492
rect 14047 27489 14059 27523
rect 14001 27483 14059 27489
rect 14369 27523 14427 27529
rect 14369 27489 14381 27523
rect 14415 27520 14427 27523
rect 14458 27520 14464 27532
rect 14415 27492 14464 27520
rect 14415 27489 14427 27492
rect 14369 27483 14427 27489
rect 14458 27480 14464 27492
rect 14516 27480 14522 27532
rect 14550 27480 14556 27532
rect 14608 27520 14614 27532
rect 15212 27520 15240 27560
rect 15378 27548 15384 27560
rect 15436 27548 15442 27600
rect 16117 27591 16175 27597
rect 16117 27557 16129 27591
rect 16163 27588 16175 27591
rect 16163 27560 17816 27588
rect 16163 27557 16175 27560
rect 16117 27551 16175 27557
rect 15289 27523 15347 27529
rect 15289 27520 15301 27523
rect 14608 27492 14653 27520
rect 15212 27492 15301 27520
rect 14608 27480 14614 27492
rect 15289 27489 15301 27492
rect 15335 27489 15347 27523
rect 15289 27483 15347 27489
rect 16761 27523 16819 27529
rect 16761 27489 16773 27523
rect 16807 27489 16819 27523
rect 16761 27483 16819 27489
rect 13449 27455 13507 27461
rect 13449 27421 13461 27455
rect 13495 27421 13507 27455
rect 13449 27415 13507 27421
rect 13722 27384 13728 27396
rect 13372 27356 13728 27384
rect 13722 27344 13728 27356
rect 13780 27344 13786 27396
rect 6503 27288 7972 27316
rect 6503 27285 6515 27288
rect 6457 27279 6515 27285
rect 8294 27276 8300 27328
rect 8352 27316 8358 27328
rect 9030 27316 9036 27328
rect 8352 27288 9036 27316
rect 8352 27276 8358 27288
rect 9030 27276 9036 27288
rect 9088 27276 9094 27328
rect 11054 27276 11060 27328
rect 11112 27316 11118 27328
rect 11517 27319 11575 27325
rect 11517 27316 11529 27319
rect 11112 27288 11529 27316
rect 11112 27276 11118 27288
rect 11517 27285 11529 27288
rect 11563 27285 11575 27319
rect 16776 27316 16804 27483
rect 17034 27480 17040 27532
rect 17092 27520 17098 27532
rect 17788 27529 17816 27560
rect 17954 27548 17960 27600
rect 18012 27588 18018 27600
rect 21818 27588 21824 27600
rect 18012 27560 21824 27588
rect 18012 27548 18018 27560
rect 21818 27548 21824 27560
rect 21876 27588 21882 27600
rect 23566 27588 23572 27600
rect 21876 27560 23572 27588
rect 21876 27548 21882 27560
rect 23566 27548 23572 27560
rect 23624 27548 23630 27600
rect 17129 27523 17187 27529
rect 17129 27520 17141 27523
rect 17092 27492 17141 27520
rect 17092 27480 17098 27492
rect 17129 27489 17141 27492
rect 17175 27489 17187 27523
rect 17129 27483 17187 27489
rect 17773 27523 17831 27529
rect 17773 27489 17785 27523
rect 17819 27489 17831 27523
rect 17773 27483 17831 27489
rect 18509 27523 18567 27529
rect 18509 27489 18521 27523
rect 18555 27520 18567 27523
rect 19426 27520 19432 27532
rect 18555 27492 19432 27520
rect 18555 27489 18567 27492
rect 18509 27483 18567 27489
rect 19426 27480 19432 27492
rect 19484 27480 19490 27532
rect 19797 27523 19855 27529
rect 19797 27489 19809 27523
rect 19843 27520 19855 27523
rect 19886 27520 19892 27532
rect 19843 27492 19892 27520
rect 19843 27489 19855 27492
rect 19797 27483 19855 27489
rect 19886 27480 19892 27492
rect 19944 27480 19950 27532
rect 19978 27480 19984 27532
rect 20036 27520 20042 27532
rect 20073 27523 20131 27529
rect 20073 27520 20085 27523
rect 20036 27492 20085 27520
rect 20036 27480 20042 27492
rect 20073 27489 20085 27492
rect 20119 27489 20131 27523
rect 20714 27520 20720 27532
rect 20073 27483 20131 27489
rect 20180 27492 20720 27520
rect 16853 27455 16911 27461
rect 16853 27421 16865 27455
rect 16899 27421 16911 27455
rect 17218 27452 17224 27464
rect 17179 27424 17224 27452
rect 16853 27415 16911 27421
rect 16868 27384 16896 27415
rect 17218 27412 17224 27424
rect 17276 27412 17282 27464
rect 17402 27412 17408 27464
rect 17460 27452 17466 27464
rect 19337 27455 19395 27461
rect 17460 27424 18000 27452
rect 17460 27412 17466 27424
rect 17034 27384 17040 27396
rect 16868 27356 17040 27384
rect 17034 27344 17040 27356
rect 17092 27384 17098 27396
rect 17310 27384 17316 27396
rect 17092 27356 17316 27384
rect 17092 27344 17098 27356
rect 17310 27344 17316 27356
rect 17368 27344 17374 27396
rect 17862 27384 17868 27396
rect 17823 27356 17868 27384
rect 17862 27344 17868 27356
rect 17920 27344 17926 27396
rect 17972 27384 18000 27424
rect 19337 27421 19349 27455
rect 19383 27452 19395 27455
rect 20180 27452 20208 27492
rect 20714 27480 20720 27492
rect 20772 27480 20778 27532
rect 21082 27520 21088 27532
rect 21043 27492 21088 27520
rect 21082 27480 21088 27492
rect 21140 27480 21146 27532
rect 21542 27520 21548 27532
rect 21503 27492 21548 27520
rect 21542 27480 21548 27492
rect 21600 27480 21606 27532
rect 22278 27480 22284 27532
rect 22336 27520 22342 27532
rect 23676 27529 23704 27628
rect 24026 27616 24032 27668
rect 24084 27656 24090 27668
rect 25406 27656 25412 27668
rect 24084 27628 25412 27656
rect 24084 27616 24090 27628
rect 25406 27616 25412 27628
rect 25464 27616 25470 27668
rect 25682 27616 25688 27668
rect 25740 27656 25746 27668
rect 27522 27656 27528 27668
rect 25740 27628 27528 27656
rect 25740 27616 25746 27628
rect 27522 27616 27528 27628
rect 27580 27656 27586 27668
rect 29638 27656 29644 27668
rect 27580 27628 29644 27656
rect 27580 27616 27586 27628
rect 24762 27548 24768 27600
rect 24820 27588 24826 27600
rect 24820 27560 26740 27588
rect 24820 27548 24826 27560
rect 22465 27523 22523 27529
rect 22465 27520 22477 27523
rect 22336 27492 22477 27520
rect 22336 27480 22342 27492
rect 22465 27489 22477 27492
rect 22511 27489 22523 27523
rect 22465 27483 22523 27489
rect 23661 27523 23719 27529
rect 23661 27489 23673 27523
rect 23707 27489 23719 27523
rect 23661 27483 23719 27489
rect 24213 27523 24271 27529
rect 24213 27489 24225 27523
rect 24259 27489 24271 27523
rect 24213 27483 24271 27489
rect 20346 27452 20352 27464
rect 19383 27424 20208 27452
rect 20307 27424 20352 27452
rect 19383 27421 19395 27424
rect 19337 27415 19395 27421
rect 20346 27412 20352 27424
rect 20404 27412 20410 27464
rect 21913 27455 21971 27461
rect 20456 27424 21588 27452
rect 20456 27384 20484 27424
rect 17972 27356 20484 27384
rect 20806 27344 20812 27396
rect 20864 27384 20870 27396
rect 20993 27387 21051 27393
rect 20993 27384 21005 27387
rect 20864 27356 21005 27384
rect 20864 27344 20870 27356
rect 20993 27353 21005 27356
rect 21039 27353 21051 27387
rect 20993 27347 21051 27353
rect 18598 27316 18604 27328
rect 16776 27288 18604 27316
rect 11517 27279 11575 27285
rect 18598 27276 18604 27288
rect 18656 27316 18662 27328
rect 21358 27316 21364 27328
rect 18656 27288 21364 27316
rect 18656 27276 18662 27288
rect 21358 27276 21364 27288
rect 21416 27276 21422 27328
rect 21560 27316 21588 27424
rect 21913 27421 21925 27455
rect 21959 27452 21971 27455
rect 23477 27455 23535 27461
rect 21959 27424 23428 27452
rect 21959 27421 21971 27424
rect 21913 27415 21971 27421
rect 21726 27344 21732 27396
rect 21784 27384 21790 27396
rect 22649 27387 22707 27393
rect 22649 27384 22661 27387
rect 21784 27356 22661 27384
rect 21784 27344 21790 27356
rect 22649 27353 22661 27356
rect 22695 27353 22707 27387
rect 22649 27347 22707 27353
rect 22462 27316 22468 27328
rect 21560 27288 22468 27316
rect 22462 27276 22468 27288
rect 22520 27276 22526 27328
rect 23400 27316 23428 27424
rect 23477 27421 23489 27455
rect 23523 27452 23535 27455
rect 23934 27452 23940 27464
rect 23523 27424 23940 27452
rect 23523 27421 23535 27424
rect 23477 27415 23535 27421
rect 23934 27412 23940 27424
rect 23992 27412 23998 27464
rect 24228 27452 24256 27483
rect 24486 27480 24492 27532
rect 24544 27520 24550 27532
rect 25133 27523 25191 27529
rect 24544 27492 25084 27520
rect 24544 27480 24550 27492
rect 24228 27424 24992 27452
rect 24026 27344 24032 27396
rect 24084 27384 24090 27396
rect 24964 27393 24992 27424
rect 24121 27387 24179 27393
rect 24121 27384 24133 27387
rect 24084 27356 24133 27384
rect 24084 27344 24090 27356
rect 24121 27353 24133 27356
rect 24167 27353 24179 27387
rect 24121 27347 24179 27353
rect 24949 27387 25007 27393
rect 24949 27353 24961 27387
rect 24995 27353 25007 27387
rect 25056 27384 25084 27492
rect 25133 27489 25145 27523
rect 25179 27520 25191 27523
rect 25406 27520 25412 27532
rect 25179 27492 25412 27520
rect 25179 27489 25191 27492
rect 25133 27483 25191 27489
rect 25406 27480 25412 27492
rect 25464 27480 25470 27532
rect 25590 27520 25596 27532
rect 25551 27492 25596 27520
rect 25590 27480 25596 27492
rect 25648 27480 25654 27532
rect 26712 27529 26740 27560
rect 27062 27548 27068 27600
rect 27120 27588 27126 27600
rect 27816 27597 27844 27628
rect 29638 27616 29644 27628
rect 29696 27616 29702 27668
rect 27433 27591 27491 27597
rect 27433 27588 27445 27591
rect 27120 27560 27445 27588
rect 27120 27548 27126 27560
rect 27433 27557 27445 27560
rect 27479 27557 27491 27591
rect 27433 27551 27491 27557
rect 27801 27591 27859 27597
rect 27801 27557 27813 27591
rect 27847 27557 27859 27591
rect 27801 27551 27859 27557
rect 28169 27591 28227 27597
rect 28169 27557 28181 27591
rect 28215 27588 28227 27591
rect 28258 27588 28264 27600
rect 28215 27560 28264 27588
rect 28215 27557 28227 27560
rect 28169 27551 28227 27557
rect 28258 27548 28264 27560
rect 28316 27548 28322 27600
rect 34514 27588 34520 27600
rect 28920 27560 31064 27588
rect 28920 27529 28948 27560
rect 26697 27523 26755 27529
rect 26697 27489 26709 27523
rect 26743 27520 26755 27523
rect 27617 27523 27675 27529
rect 27617 27520 27629 27523
rect 26743 27492 27629 27520
rect 26743 27489 26755 27492
rect 26697 27483 26755 27489
rect 27617 27489 27629 27492
rect 27663 27489 27675 27523
rect 27617 27483 27675 27489
rect 27709 27523 27767 27529
rect 27709 27489 27721 27523
rect 27755 27489 27767 27523
rect 27709 27483 27767 27489
rect 28905 27523 28963 27529
rect 28905 27489 28917 27523
rect 28951 27489 28963 27523
rect 29086 27520 29092 27532
rect 29047 27492 29092 27520
rect 28905 27483 28963 27489
rect 27724 27452 27752 27483
rect 29086 27480 29092 27492
rect 29144 27480 29150 27532
rect 29178 27480 29184 27532
rect 29236 27520 29242 27532
rect 29457 27523 29515 27529
rect 29457 27520 29469 27523
rect 29236 27492 29469 27520
rect 29236 27480 29242 27492
rect 29457 27489 29469 27492
rect 29503 27520 29515 27523
rect 30466 27520 30472 27532
rect 29503 27492 30472 27520
rect 29503 27489 29515 27492
rect 29457 27483 29515 27489
rect 30466 27480 30472 27492
rect 30524 27480 30530 27532
rect 30650 27520 30656 27532
rect 30611 27492 30656 27520
rect 30650 27480 30656 27492
rect 30708 27480 30714 27532
rect 27724 27424 29776 27452
rect 28994 27384 29000 27396
rect 25056 27356 29000 27384
rect 24949 27347 25007 27353
rect 28994 27344 29000 27356
rect 29052 27344 29058 27396
rect 29454 27384 29460 27396
rect 29415 27356 29460 27384
rect 29454 27344 29460 27356
rect 29512 27344 29518 27396
rect 29748 27328 29776 27424
rect 30374 27412 30380 27464
rect 30432 27452 30438 27464
rect 31036 27461 31064 27560
rect 33244 27560 34520 27588
rect 32030 27480 32036 27532
rect 32088 27520 32094 27532
rect 33244 27529 33272 27560
rect 34514 27548 34520 27560
rect 34572 27548 34578 27600
rect 36633 27591 36691 27597
rect 36633 27557 36645 27591
rect 36679 27588 36691 27591
rect 37090 27588 37096 27600
rect 36679 27560 37096 27588
rect 36679 27557 36691 27560
rect 36633 27551 36691 27557
rect 37090 27548 37096 27560
rect 37148 27548 37154 27600
rect 37185 27591 37243 27597
rect 37185 27557 37197 27591
rect 37231 27588 37243 27591
rect 38378 27588 38384 27600
rect 37231 27560 38384 27588
rect 37231 27557 37243 27560
rect 37185 27551 37243 27557
rect 38378 27548 38384 27560
rect 38436 27548 38442 27600
rect 32401 27523 32459 27529
rect 32401 27520 32413 27523
rect 32088 27492 32413 27520
rect 32088 27480 32094 27492
rect 32401 27489 32413 27492
rect 32447 27489 32459 27523
rect 32401 27483 32459 27489
rect 33229 27523 33287 27529
rect 33229 27489 33241 27523
rect 33275 27489 33287 27523
rect 33229 27483 33287 27489
rect 33318 27480 33324 27532
rect 33376 27520 33382 27532
rect 33413 27523 33471 27529
rect 33413 27520 33425 27523
rect 33376 27492 33425 27520
rect 33376 27480 33382 27492
rect 33413 27489 33425 27492
rect 33459 27489 33471 27523
rect 33413 27483 33471 27489
rect 33781 27523 33839 27529
rect 33781 27489 33793 27523
rect 33827 27520 33839 27523
rect 33962 27520 33968 27532
rect 33827 27492 33968 27520
rect 33827 27489 33839 27492
rect 33781 27483 33839 27489
rect 33962 27480 33968 27492
rect 34020 27480 34026 27532
rect 34238 27520 34244 27532
rect 34199 27492 34244 27520
rect 34238 27480 34244 27492
rect 34296 27480 34302 27532
rect 35529 27523 35587 27529
rect 35529 27489 35541 27523
rect 35575 27520 35587 27523
rect 35710 27520 35716 27532
rect 35575 27492 35716 27520
rect 35575 27489 35587 27492
rect 35529 27483 35587 27489
rect 35710 27480 35716 27492
rect 35768 27480 35774 27532
rect 35802 27480 35808 27532
rect 35860 27520 35866 27532
rect 36817 27523 36875 27529
rect 35860 27492 35905 27520
rect 35860 27480 35866 27492
rect 36817 27489 36829 27523
rect 36863 27520 36875 27523
rect 38010 27520 38016 27532
rect 36863 27492 38016 27520
rect 36863 27489 36875 27492
rect 36817 27483 36875 27489
rect 38010 27480 38016 27492
rect 38068 27480 38074 27532
rect 38286 27520 38292 27532
rect 38247 27492 38292 27520
rect 38286 27480 38292 27492
rect 38344 27480 38350 27532
rect 38562 27480 38568 27532
rect 38620 27520 38626 27532
rect 38657 27523 38715 27529
rect 38657 27520 38669 27523
rect 38620 27492 38669 27520
rect 38620 27480 38626 27492
rect 38657 27489 38669 27492
rect 38703 27489 38715 27523
rect 38657 27483 38715 27489
rect 30800 27455 30858 27461
rect 30800 27452 30812 27455
rect 30432 27424 30812 27452
rect 30432 27412 30438 27424
rect 30800 27421 30812 27424
rect 30846 27421 30858 27455
rect 30800 27415 30858 27421
rect 31021 27455 31079 27461
rect 31021 27421 31033 27455
rect 31067 27452 31079 27455
rect 31846 27452 31852 27464
rect 31067 27424 31852 27452
rect 31067 27421 31079 27424
rect 31021 27415 31079 27421
rect 31846 27412 31852 27424
rect 31904 27412 31910 27464
rect 33042 27412 33048 27464
rect 33100 27452 33106 27464
rect 35069 27455 35127 27461
rect 35069 27452 35081 27455
rect 33100 27424 35081 27452
rect 33100 27412 33106 27424
rect 35069 27421 35081 27424
rect 35115 27421 35127 27455
rect 35069 27415 35127 27421
rect 30926 27384 30932 27396
rect 30887 27356 30932 27384
rect 30926 27344 30932 27356
rect 30984 27344 30990 27396
rect 31478 27344 31484 27396
rect 31536 27384 31542 27396
rect 32490 27384 32496 27396
rect 31536 27356 32352 27384
rect 32403 27356 32496 27384
rect 31536 27344 31542 27356
rect 24854 27316 24860 27328
rect 23400 27288 24860 27316
rect 24854 27276 24860 27288
rect 24912 27276 24918 27328
rect 26881 27319 26939 27325
rect 26881 27285 26893 27319
rect 26927 27316 26939 27319
rect 26970 27316 26976 27328
rect 26927 27288 26976 27316
rect 26927 27285 26939 27288
rect 26881 27279 26939 27285
rect 26970 27276 26976 27288
rect 27028 27276 27034 27328
rect 29730 27276 29736 27328
rect 29788 27316 29794 27328
rect 30558 27316 30564 27328
rect 29788 27288 30564 27316
rect 29788 27276 29794 27288
rect 30558 27276 30564 27288
rect 30616 27276 30622 27328
rect 31018 27276 31024 27328
rect 31076 27316 31082 27328
rect 31113 27319 31171 27325
rect 31113 27316 31125 27319
rect 31076 27288 31125 27316
rect 31076 27276 31082 27288
rect 31113 27285 31125 27288
rect 31159 27285 31171 27319
rect 32324 27316 32352 27356
rect 32490 27344 32496 27356
rect 32548 27384 32554 27396
rect 33962 27384 33968 27396
rect 32548 27356 33968 27384
rect 32548 27344 32554 27356
rect 33962 27344 33968 27356
rect 34020 27344 34026 27396
rect 35894 27384 35900 27396
rect 34072 27356 35296 27384
rect 35855 27356 35900 27384
rect 34072 27316 34100 27356
rect 32324 27288 34100 27316
rect 31113 27279 31171 27285
rect 34146 27276 34152 27328
rect 34204 27316 34210 27328
rect 34425 27319 34483 27325
rect 34425 27316 34437 27319
rect 34204 27288 34437 27316
rect 34204 27276 34210 27288
rect 34425 27285 34437 27288
rect 34471 27285 34483 27319
rect 35268 27316 35296 27356
rect 35894 27344 35900 27356
rect 35952 27344 35958 27396
rect 36630 27344 36636 27396
rect 36688 27384 36694 27396
rect 38657 27387 38715 27393
rect 38657 27384 38669 27387
rect 36688 27356 38669 27384
rect 36688 27344 36694 27356
rect 38657 27353 38669 27356
rect 38703 27353 38715 27387
rect 38657 27347 38715 27353
rect 38838 27316 38844 27328
rect 35268 27288 38844 27316
rect 34425 27279 34483 27285
rect 38838 27276 38844 27288
rect 38896 27276 38902 27328
rect 39942 27248 39948 27260
rect 1104 27226 39836 27248
rect 1104 27174 4246 27226
rect 4298 27174 4310 27226
rect 4362 27174 4374 27226
rect 4426 27174 4438 27226
rect 4490 27174 34966 27226
rect 35018 27174 35030 27226
rect 35082 27174 35094 27226
rect 35146 27174 35158 27226
rect 35210 27174 39836 27226
rect 39903 27220 39948 27248
rect 39942 27208 39948 27220
rect 40000 27208 40006 27260
rect 1104 27152 39836 27174
rect 5077 27115 5135 27121
rect 5077 27081 5089 27115
rect 5123 27112 5135 27115
rect 5626 27112 5632 27124
rect 5123 27084 5632 27112
rect 5123 27081 5135 27084
rect 5077 27075 5135 27081
rect 5626 27072 5632 27084
rect 5684 27072 5690 27124
rect 6181 27115 6239 27121
rect 6181 27081 6193 27115
rect 6227 27112 6239 27115
rect 6638 27112 6644 27124
rect 6227 27084 6644 27112
rect 6227 27081 6239 27084
rect 6181 27075 6239 27081
rect 6638 27072 6644 27084
rect 6696 27072 6702 27124
rect 9585 27115 9643 27121
rect 9585 27081 9597 27115
rect 9631 27112 9643 27115
rect 13446 27112 13452 27124
rect 9631 27084 13452 27112
rect 9631 27081 9643 27084
rect 9585 27075 9643 27081
rect 13446 27072 13452 27084
rect 13504 27072 13510 27124
rect 13722 27072 13728 27124
rect 13780 27112 13786 27124
rect 13780 27084 18092 27112
rect 13780 27072 13786 27084
rect 1857 26979 1915 26985
rect 1857 26945 1869 26979
rect 1903 26976 1915 26979
rect 2774 26976 2780 26988
rect 1903 26948 2780 26976
rect 1903 26945 1915 26948
rect 1857 26939 1915 26945
rect 2774 26936 2780 26948
rect 2832 26936 2838 26988
rect 5718 26936 5724 26988
rect 5776 26976 5782 26988
rect 7101 26979 7159 26985
rect 7101 26976 7113 26979
rect 5776 26948 7113 26976
rect 5776 26936 5782 26948
rect 7101 26945 7113 26948
rect 7147 26945 7159 26979
rect 10502 26976 10508 26988
rect 7101 26939 7159 26945
rect 10336 26948 10508 26976
rect 1394 26868 1400 26920
rect 1452 26908 1458 26920
rect 1581 26911 1639 26917
rect 1581 26908 1593 26911
rect 1452 26880 1593 26908
rect 1452 26868 1458 26880
rect 1581 26877 1593 26880
rect 1627 26877 1639 26911
rect 1581 26871 1639 26877
rect 2590 26868 2596 26920
rect 2648 26908 2654 26920
rect 3237 26911 3295 26917
rect 3237 26908 3249 26911
rect 2648 26880 3249 26908
rect 2648 26868 2654 26880
rect 3237 26877 3249 26880
rect 3283 26908 3295 26911
rect 3697 26911 3755 26917
rect 3697 26908 3709 26911
rect 3283 26880 3709 26908
rect 3283 26877 3295 26880
rect 3237 26871 3295 26877
rect 3697 26877 3709 26880
rect 3743 26877 3755 26911
rect 4246 26908 4252 26920
rect 4207 26880 4252 26908
rect 3697 26871 3755 26877
rect 4246 26868 4252 26880
rect 4304 26868 4310 26920
rect 4709 26911 4767 26917
rect 4709 26877 4721 26911
rect 4755 26908 4767 26911
rect 4798 26908 4804 26920
rect 4755 26880 4804 26908
rect 4755 26877 4767 26880
rect 4709 26871 4767 26877
rect 4798 26868 4804 26880
rect 4856 26868 4862 26920
rect 5169 26911 5227 26917
rect 5169 26877 5181 26911
rect 5215 26908 5227 26911
rect 5626 26908 5632 26920
rect 5215 26880 5632 26908
rect 5215 26877 5227 26880
rect 5169 26871 5227 26877
rect 5626 26868 5632 26880
rect 5684 26868 5690 26920
rect 5994 26908 6000 26920
rect 5955 26880 6000 26908
rect 5994 26868 6000 26880
rect 6052 26868 6058 26920
rect 6546 26868 6552 26920
rect 6604 26908 6610 26920
rect 6825 26911 6883 26917
rect 6825 26908 6837 26911
rect 6604 26880 6837 26908
rect 6604 26868 6610 26880
rect 6825 26877 6837 26880
rect 6871 26877 6883 26911
rect 6825 26871 6883 26877
rect 9030 26868 9036 26920
rect 9088 26908 9094 26920
rect 10336 26917 10364 26948
rect 10502 26936 10508 26948
rect 10560 26936 10566 26988
rect 10594 26936 10600 26988
rect 10652 26976 10658 26988
rect 10870 26976 10876 26988
rect 10652 26948 10876 26976
rect 10652 26936 10658 26948
rect 10870 26936 10876 26948
rect 10928 26936 10934 26988
rect 11517 26979 11575 26985
rect 11517 26945 11529 26979
rect 11563 26976 11575 26979
rect 17954 26976 17960 26988
rect 11563 26948 12480 26976
rect 11563 26945 11575 26948
rect 11517 26939 11575 26945
rect 9401 26911 9459 26917
rect 9401 26908 9413 26911
rect 9088 26880 9413 26908
rect 9088 26868 9094 26880
rect 9401 26877 9413 26880
rect 9447 26877 9459 26911
rect 9401 26871 9459 26877
rect 10321 26911 10379 26917
rect 10321 26877 10333 26911
rect 10367 26877 10379 26911
rect 10321 26871 10379 26877
rect 10413 26911 10471 26917
rect 10413 26877 10425 26911
rect 10459 26908 10471 26911
rect 11054 26908 11060 26920
rect 10459 26880 11060 26908
rect 10459 26877 10471 26880
rect 10413 26871 10471 26877
rect 11054 26868 11060 26880
rect 11112 26868 11118 26920
rect 11422 26908 11428 26920
rect 11383 26880 11428 26908
rect 11422 26868 11428 26880
rect 11480 26868 11486 26920
rect 11882 26908 11888 26920
rect 11843 26880 11888 26908
rect 11882 26868 11888 26880
rect 11940 26868 11946 26920
rect 12452 26917 12480 26948
rect 15672 26948 17960 26976
rect 12437 26911 12495 26917
rect 12437 26877 12449 26911
rect 12483 26877 12495 26911
rect 13538 26908 13544 26920
rect 13499 26880 13544 26908
rect 12437 26871 12495 26877
rect 13538 26868 13544 26880
rect 13596 26868 13602 26920
rect 13814 26868 13820 26920
rect 13872 26908 13878 26920
rect 15672 26917 15700 26948
rect 17954 26936 17960 26948
rect 18012 26936 18018 26988
rect 15657 26911 15715 26917
rect 13872 26880 13917 26908
rect 13872 26868 13878 26880
rect 15657 26877 15669 26911
rect 15703 26877 15715 26911
rect 16574 26908 16580 26920
rect 16535 26880 16580 26908
rect 15657 26871 15715 26877
rect 16574 26868 16580 26880
rect 16632 26868 16638 26920
rect 16850 26908 16856 26920
rect 16811 26880 16856 26908
rect 16850 26868 16856 26880
rect 16908 26868 16914 26920
rect 17313 26911 17371 26917
rect 17313 26877 17325 26911
rect 17359 26908 17371 26911
rect 17402 26908 17408 26920
rect 17359 26880 17408 26908
rect 17359 26877 17371 26880
rect 17313 26871 17371 26877
rect 17402 26868 17408 26880
rect 17460 26868 17466 26920
rect 18064 26917 18092 27084
rect 23566 27072 23572 27124
rect 23624 27112 23630 27124
rect 25961 27115 26019 27121
rect 25961 27112 25973 27115
rect 23624 27084 25973 27112
rect 23624 27072 23630 27084
rect 25961 27081 25973 27084
rect 26007 27081 26019 27115
rect 25961 27075 26019 27081
rect 29622 27115 29680 27121
rect 29622 27081 29634 27115
rect 29668 27112 29680 27115
rect 32033 27115 32091 27121
rect 32033 27112 32045 27115
rect 29668 27084 32045 27112
rect 29668 27081 29680 27084
rect 29622 27075 29680 27081
rect 32033 27081 32045 27084
rect 32079 27081 32091 27115
rect 32033 27075 32091 27081
rect 34790 27072 34796 27124
rect 34848 27112 34854 27124
rect 35161 27115 35219 27121
rect 35161 27112 35173 27115
rect 34848 27084 35173 27112
rect 34848 27072 34854 27084
rect 35161 27081 35173 27084
rect 35207 27112 35219 27115
rect 35618 27112 35624 27124
rect 35207 27084 35624 27112
rect 35207 27081 35219 27084
rect 35161 27075 35219 27081
rect 35618 27072 35624 27084
rect 35676 27072 35682 27124
rect 18156 27016 19564 27044
rect 18049 26911 18107 26917
rect 18049 26877 18061 26911
rect 18095 26877 18107 26911
rect 18049 26871 18107 26877
rect 8481 26843 8539 26849
rect 8481 26809 8493 26843
rect 8527 26840 8539 26843
rect 8570 26840 8576 26852
rect 8527 26812 8576 26840
rect 8527 26809 8539 26812
rect 8481 26803 8539 26809
rect 8570 26800 8576 26812
rect 8628 26840 8634 26852
rect 11900 26840 11928 26868
rect 8628 26812 11928 26840
rect 8628 26800 8634 26812
rect 11974 26800 11980 26852
rect 12032 26840 12038 26852
rect 13630 26840 13636 26852
rect 12032 26812 13636 26840
rect 12032 26800 12038 26812
rect 13630 26800 13636 26812
rect 13688 26800 13694 26852
rect 15197 26843 15255 26849
rect 15197 26809 15209 26843
rect 15243 26840 15255 26843
rect 15470 26840 15476 26852
rect 15243 26812 15476 26840
rect 15243 26809 15255 26812
rect 15197 26803 15255 26809
rect 2498 26732 2504 26784
rect 2556 26772 2562 26784
rect 5718 26772 5724 26784
rect 2556 26744 5724 26772
rect 2556 26732 2562 26744
rect 5718 26732 5724 26744
rect 5776 26732 5782 26784
rect 9674 26732 9680 26784
rect 9732 26772 9738 26784
rect 10137 26775 10195 26781
rect 10137 26772 10149 26775
rect 9732 26744 10149 26772
rect 9732 26732 9738 26744
rect 10137 26741 10149 26744
rect 10183 26741 10195 26775
rect 10594 26772 10600 26784
rect 10555 26744 10600 26772
rect 10137 26735 10195 26741
rect 10594 26732 10600 26744
rect 10652 26732 10658 26784
rect 12434 26732 12440 26784
rect 12492 26772 12498 26784
rect 12529 26775 12587 26781
rect 12529 26772 12541 26775
rect 12492 26744 12541 26772
rect 12492 26732 12498 26744
rect 12529 26741 12541 26744
rect 12575 26741 12587 26775
rect 12529 26735 12587 26741
rect 13814 26732 13820 26784
rect 13872 26772 13878 26784
rect 15212 26772 15240 26803
rect 15470 26800 15476 26812
rect 15528 26800 15534 26852
rect 17497 26843 17555 26849
rect 17497 26809 17509 26843
rect 17543 26840 17555 26843
rect 18156 26840 18184 27016
rect 19150 26976 19156 26988
rect 18340 26948 19156 26976
rect 18340 26917 18368 26948
rect 19150 26936 19156 26948
rect 19208 26936 19214 26988
rect 18325 26911 18383 26917
rect 18325 26877 18337 26911
rect 18371 26877 18383 26911
rect 18325 26871 18383 26877
rect 18509 26911 18567 26917
rect 18509 26877 18521 26911
rect 18555 26908 18567 26911
rect 18598 26908 18604 26920
rect 18555 26880 18604 26908
rect 18555 26877 18567 26880
rect 18509 26871 18567 26877
rect 18598 26868 18604 26880
rect 18656 26868 18662 26920
rect 18782 26908 18788 26920
rect 18743 26880 18788 26908
rect 18782 26868 18788 26880
rect 18840 26868 18846 26920
rect 18978 26911 19036 26917
rect 18978 26908 18990 26911
rect 18892 26880 18990 26908
rect 18892 26840 18920 26880
rect 18978 26877 18990 26880
rect 19024 26877 19036 26911
rect 18978 26871 19036 26877
rect 17543 26812 18184 26840
rect 18708 26812 18920 26840
rect 19536 26840 19564 27016
rect 22186 27004 22192 27056
rect 22244 27044 22250 27056
rect 22244 27016 22416 27044
rect 22244 27004 22250 27016
rect 20441 26979 20499 26985
rect 20441 26945 20453 26979
rect 20487 26976 20499 26979
rect 20530 26976 20536 26988
rect 20487 26948 20536 26976
rect 20487 26945 20499 26948
rect 20441 26939 20499 26945
rect 20530 26936 20536 26948
rect 20588 26936 20594 26988
rect 22094 26976 22100 26988
rect 21928 26948 22100 26976
rect 19613 26911 19671 26917
rect 19613 26877 19625 26911
rect 19659 26908 19671 26911
rect 20073 26911 20131 26917
rect 20073 26908 20085 26911
rect 19659 26880 20085 26908
rect 19659 26877 19671 26880
rect 19613 26871 19671 26877
rect 20073 26877 20085 26880
rect 20119 26877 20131 26911
rect 20073 26871 20131 26877
rect 20346 26868 20352 26920
rect 20404 26908 20410 26920
rect 21928 26917 21956 26948
rect 22094 26936 22100 26948
rect 22152 26936 22158 26988
rect 22388 26985 22416 27016
rect 25314 27004 25320 27056
rect 25372 27044 25378 27056
rect 27985 27047 28043 27053
rect 25372 27016 26004 27044
rect 25372 27004 25378 27016
rect 25976 26988 26004 27016
rect 27985 27013 27997 27047
rect 28031 27044 28043 27047
rect 29730 27044 29736 27056
rect 28031 27016 29592 27044
rect 29691 27016 29736 27044
rect 28031 27013 28043 27016
rect 27985 27007 28043 27013
rect 22373 26979 22431 26985
rect 22373 26945 22385 26979
rect 22419 26945 22431 26979
rect 24026 26976 24032 26988
rect 23987 26948 24032 26976
rect 22373 26939 22431 26945
rect 24026 26936 24032 26948
rect 24084 26936 24090 26988
rect 24762 26936 24768 26988
rect 24820 26976 24826 26988
rect 24820 26948 25912 26976
rect 24820 26936 24826 26948
rect 20625 26911 20683 26917
rect 20625 26908 20637 26911
rect 20404 26880 20637 26908
rect 20404 26868 20410 26880
rect 20625 26877 20637 26880
rect 20671 26877 20683 26911
rect 20625 26871 20683 26877
rect 21913 26911 21971 26917
rect 21913 26877 21925 26911
rect 21959 26877 21971 26911
rect 22186 26908 22192 26920
rect 22147 26880 22192 26908
rect 21913 26871 21971 26877
rect 22186 26868 22192 26880
rect 22244 26868 22250 26920
rect 22738 26868 22744 26920
rect 22796 26908 22802 26920
rect 22833 26911 22891 26917
rect 22833 26908 22845 26911
rect 22796 26880 22845 26908
rect 22796 26868 22802 26880
rect 22833 26877 22845 26880
rect 22879 26877 22891 26911
rect 22833 26871 22891 26877
rect 23566 26868 23572 26920
rect 23624 26908 23630 26920
rect 25884 26917 25912 26948
rect 25958 26936 25964 26988
rect 26016 26976 26022 26988
rect 29454 26976 29460 26988
rect 26016 26948 26109 26976
rect 28184 26948 29460 26976
rect 26016 26936 26022 26948
rect 23753 26911 23811 26917
rect 23753 26908 23765 26911
rect 23624 26880 23765 26908
rect 23624 26868 23630 26880
rect 23753 26877 23765 26880
rect 23799 26877 23811 26911
rect 25869 26911 25927 26917
rect 23753 26871 23811 26877
rect 23860 26880 25360 26908
rect 23860 26840 23888 26880
rect 19536 26812 23888 26840
rect 17543 26809 17555 26812
rect 17497 26803 17555 26809
rect 13872 26744 15240 26772
rect 15841 26775 15899 26781
rect 13872 26732 13878 26744
rect 15841 26741 15853 26775
rect 15887 26772 15899 26775
rect 17862 26772 17868 26784
rect 15887 26744 17868 26772
rect 15887 26741 15899 26744
rect 15841 26735 15899 26741
rect 17862 26732 17868 26744
rect 17920 26772 17926 26784
rect 18708 26772 18736 26812
rect 17920 26744 18736 26772
rect 17920 26732 17926 26744
rect 19150 26732 19156 26784
rect 19208 26772 19214 26784
rect 22554 26772 22560 26784
rect 19208 26744 22560 26772
rect 19208 26732 19214 26744
rect 22554 26732 22560 26744
rect 22612 26732 22618 26784
rect 23014 26772 23020 26784
rect 22975 26744 23020 26772
rect 23014 26732 23020 26744
rect 23072 26732 23078 26784
rect 25332 26772 25360 26880
rect 25869 26877 25881 26911
rect 25915 26877 25927 26911
rect 25976 26908 26004 26936
rect 26237 26911 26295 26917
rect 26237 26908 26249 26911
rect 25976 26880 26249 26908
rect 25869 26871 25927 26877
rect 26237 26877 26249 26880
rect 26283 26877 26295 26911
rect 26878 26908 26884 26920
rect 26839 26880 26884 26908
rect 26237 26871 26295 26877
rect 26878 26868 26884 26880
rect 26936 26868 26942 26920
rect 28184 26917 28212 26948
rect 29454 26936 29460 26948
rect 29512 26936 29518 26988
rect 29564 26976 29592 27016
rect 29730 27004 29736 27016
rect 29788 27004 29794 27056
rect 30282 27044 30288 27056
rect 29840 27016 30288 27044
rect 29840 26985 29868 27016
rect 30282 27004 30288 27016
rect 30340 27004 30346 27056
rect 36078 27044 36084 27056
rect 36039 27016 36084 27044
rect 36078 27004 36084 27016
rect 36136 27004 36142 27056
rect 29825 26979 29883 26985
rect 29564 26948 29776 26976
rect 28169 26911 28227 26917
rect 28169 26877 28181 26911
rect 28215 26877 28227 26911
rect 28169 26871 28227 26877
rect 28537 26911 28595 26917
rect 28537 26877 28549 26911
rect 28583 26877 28595 26911
rect 28537 26871 28595 26877
rect 25406 26800 25412 26852
rect 25464 26840 25470 26852
rect 28350 26840 28356 26852
rect 25464 26812 28356 26840
rect 25464 26800 25470 26812
rect 28350 26800 28356 26812
rect 28408 26800 28414 26852
rect 28552 26772 28580 26871
rect 28626 26868 28632 26920
rect 28684 26908 28690 26920
rect 29748 26908 29776 26948
rect 29825 26945 29837 26979
rect 29871 26945 29883 26979
rect 34146 26976 34152 26988
rect 29825 26939 29883 26945
rect 29932 26948 33732 26976
rect 34107 26948 34152 26976
rect 29932 26908 29960 26948
rect 28684 26880 28729 26908
rect 29748 26880 29960 26908
rect 28684 26868 28690 26880
rect 30006 26868 30012 26920
rect 30064 26908 30070 26920
rect 30653 26911 30711 26917
rect 30653 26908 30665 26911
rect 30064 26880 30665 26908
rect 30064 26868 30070 26880
rect 30653 26877 30665 26880
rect 30699 26877 30711 26911
rect 30926 26908 30932 26920
rect 30887 26880 30932 26908
rect 30653 26871 30711 26877
rect 30926 26868 30932 26880
rect 30984 26868 30990 26920
rect 33134 26908 33140 26920
rect 33095 26880 33140 26908
rect 33134 26868 33140 26880
rect 33192 26868 33198 26920
rect 33704 26917 33732 26948
rect 34146 26936 34152 26948
rect 34204 26936 34210 26988
rect 36909 26979 36967 26985
rect 36909 26945 36921 26979
rect 36955 26976 36967 26979
rect 37826 26976 37832 26988
rect 36955 26948 37832 26976
rect 36955 26945 36967 26948
rect 36909 26939 36967 26945
rect 37826 26936 37832 26948
rect 37884 26936 37890 26988
rect 38562 26976 38568 26988
rect 38523 26948 38568 26976
rect 38562 26936 38568 26948
rect 38620 26936 38626 26988
rect 33689 26911 33747 26917
rect 33689 26877 33701 26911
rect 33735 26877 33747 26911
rect 33689 26871 33747 26877
rect 34054 26868 34060 26920
rect 34112 26908 34118 26920
rect 34977 26911 35035 26917
rect 34977 26908 34989 26911
rect 34112 26880 34989 26908
rect 34112 26868 34118 26880
rect 34977 26877 34989 26880
rect 35023 26908 35035 26911
rect 35250 26908 35256 26920
rect 35023 26880 35256 26908
rect 35023 26877 35035 26880
rect 34977 26871 35035 26877
rect 35250 26868 35256 26880
rect 35308 26868 35314 26920
rect 35894 26908 35900 26920
rect 35855 26880 35900 26908
rect 35894 26868 35900 26880
rect 35952 26868 35958 26920
rect 36630 26908 36636 26920
rect 36591 26880 36636 26908
rect 36630 26868 36636 26880
rect 36688 26868 36694 26920
rect 37734 26868 37740 26920
rect 37792 26908 37798 26920
rect 38197 26911 38255 26917
rect 38197 26908 38209 26911
rect 37792 26880 38209 26908
rect 37792 26868 37798 26880
rect 38197 26877 38209 26880
rect 38243 26877 38255 26911
rect 38197 26871 38255 26877
rect 29457 26843 29515 26849
rect 29457 26809 29469 26843
rect 29503 26809 29515 26843
rect 29457 26803 29515 26809
rect 30193 26843 30251 26849
rect 30193 26809 30205 26843
rect 30239 26840 30251 26843
rect 30558 26840 30564 26852
rect 30239 26812 30564 26840
rect 30239 26809 30251 26812
rect 30193 26803 30251 26809
rect 25332 26744 28580 26772
rect 29472 26772 29500 26803
rect 30558 26800 30564 26812
rect 30616 26800 30622 26852
rect 37090 26800 37096 26852
rect 37148 26840 37154 26852
rect 38013 26843 38071 26849
rect 38013 26840 38025 26843
rect 37148 26812 38025 26840
rect 37148 26800 37154 26812
rect 38013 26809 38025 26812
rect 38059 26809 38071 26843
rect 38013 26803 38071 26809
rect 31018 26772 31024 26784
rect 29472 26744 31024 26772
rect 31018 26732 31024 26744
rect 31076 26732 31082 26784
rect 31202 26732 31208 26784
rect 31260 26772 31266 26784
rect 33042 26772 33048 26784
rect 31260 26744 33048 26772
rect 31260 26732 31266 26744
rect 33042 26732 33048 26744
rect 33100 26732 33106 26784
rect 33229 26775 33287 26781
rect 33229 26741 33241 26775
rect 33275 26772 33287 26775
rect 33778 26772 33784 26784
rect 33275 26744 33784 26772
rect 33275 26741 33287 26744
rect 33229 26735 33287 26741
rect 33778 26732 33784 26744
rect 33836 26732 33842 26784
rect 1104 26682 39836 26704
rect 1104 26630 19606 26682
rect 19658 26630 19670 26682
rect 19722 26630 19734 26682
rect 19786 26630 19798 26682
rect 19850 26630 39836 26682
rect 1104 26608 39836 26630
rect 4062 26568 4068 26580
rect 2884 26540 4068 26568
rect 2038 26500 2044 26512
rect 1999 26472 2044 26500
rect 2038 26460 2044 26472
rect 2096 26460 2102 26512
rect 2590 26432 2596 26444
rect 2551 26404 2596 26432
rect 2590 26392 2596 26404
rect 2648 26392 2654 26444
rect 2682 26392 2688 26444
rect 2740 26432 2746 26444
rect 2884 26441 2912 26540
rect 4062 26528 4068 26540
rect 4120 26528 4126 26580
rect 5626 26568 5632 26580
rect 5587 26540 5632 26568
rect 5626 26528 5632 26540
rect 5684 26528 5690 26580
rect 5718 26528 5724 26580
rect 5776 26568 5782 26580
rect 6365 26571 6423 26577
rect 6365 26568 6377 26571
rect 5776 26540 6377 26568
rect 5776 26528 5782 26540
rect 6365 26537 6377 26540
rect 6411 26537 6423 26571
rect 6365 26531 6423 26537
rect 11882 26528 11888 26580
rect 11940 26568 11946 26580
rect 18506 26568 18512 26580
rect 11940 26540 16252 26568
rect 18467 26540 18512 26568
rect 11940 26528 11946 26540
rect 12434 26500 12440 26512
rect 12268 26472 12440 26500
rect 2869 26435 2927 26441
rect 2740 26404 2785 26432
rect 2740 26392 2746 26404
rect 2869 26401 2881 26435
rect 2915 26401 2927 26435
rect 3142 26432 3148 26444
rect 3103 26404 3148 26432
rect 2869 26395 2927 26401
rect 3142 26392 3148 26404
rect 3200 26392 3206 26444
rect 3329 26435 3387 26441
rect 3329 26401 3341 26435
rect 3375 26401 3387 26435
rect 3329 26395 3387 26401
rect 3344 26364 3372 26395
rect 3970 26392 3976 26444
rect 4028 26432 4034 26444
rect 4072 26435 4130 26441
rect 4072 26432 4084 26435
rect 4028 26404 4084 26432
rect 4028 26392 4034 26404
rect 4072 26401 4084 26404
rect 4118 26401 4130 26435
rect 4072 26395 4130 26401
rect 5994 26392 6000 26444
rect 6052 26432 6058 26444
rect 6181 26435 6239 26441
rect 6181 26432 6193 26435
rect 6052 26404 6193 26432
rect 6052 26392 6058 26404
rect 6181 26401 6193 26404
rect 6227 26401 6239 26435
rect 7374 26432 7380 26444
rect 7335 26404 7380 26432
rect 6181 26395 6239 26401
rect 7374 26392 7380 26404
rect 7432 26392 7438 26444
rect 7742 26432 7748 26444
rect 7703 26404 7748 26432
rect 7742 26392 7748 26404
rect 7800 26392 7806 26444
rect 8110 26432 8116 26444
rect 8071 26404 8116 26432
rect 8110 26392 8116 26404
rect 8168 26392 8174 26444
rect 8570 26432 8576 26444
rect 8531 26404 8576 26432
rect 8570 26392 8576 26404
rect 8628 26392 8634 26444
rect 12066 26432 12072 26444
rect 12027 26404 12072 26432
rect 12066 26392 12072 26404
rect 12124 26392 12130 26444
rect 12268 26441 12296 26472
rect 12434 26460 12440 26472
rect 12492 26460 12498 26512
rect 12618 26460 12624 26512
rect 12676 26500 12682 26512
rect 12676 26472 15332 26500
rect 12676 26460 12682 26472
rect 12253 26435 12311 26441
rect 12253 26401 12265 26435
rect 12299 26401 12311 26435
rect 12253 26395 12311 26401
rect 12342 26392 12348 26444
rect 12400 26432 12406 26444
rect 12529 26435 12587 26441
rect 12529 26432 12541 26435
rect 12400 26404 12541 26432
rect 12400 26392 12406 26404
rect 12529 26401 12541 26404
rect 12575 26401 12587 26435
rect 13081 26435 13139 26441
rect 13081 26432 13093 26435
rect 12529 26395 12587 26401
rect 12728 26404 13093 26432
rect 4246 26364 4252 26376
rect 2792 26336 4252 26364
rect 2792 26308 2820 26336
rect 2774 26256 2780 26308
rect 2832 26256 2838 26308
rect 4080 26228 4108 26336
rect 4246 26324 4252 26336
rect 4304 26324 4310 26376
rect 4341 26367 4399 26373
rect 4341 26333 4353 26367
rect 4387 26364 4399 26367
rect 4706 26364 4712 26376
rect 4387 26336 4712 26364
rect 4387 26333 4399 26336
rect 4341 26327 4399 26333
rect 4706 26324 4712 26336
rect 4764 26324 4770 26376
rect 7190 26364 7196 26376
rect 7151 26336 7196 26364
rect 7190 26324 7196 26336
rect 7248 26324 7254 26376
rect 9674 26364 9680 26376
rect 9635 26336 9680 26364
rect 9674 26324 9680 26336
rect 9732 26324 9738 26376
rect 9858 26324 9864 26376
rect 9916 26364 9922 26376
rect 9953 26367 10011 26373
rect 9953 26364 9965 26367
rect 9916 26336 9965 26364
rect 9916 26324 9922 26336
rect 9953 26333 9965 26336
rect 9999 26333 10011 26367
rect 11330 26364 11336 26376
rect 11243 26336 11336 26364
rect 9953 26327 10011 26333
rect 11330 26324 11336 26336
rect 11388 26364 11394 26376
rect 12728 26364 12756 26404
rect 13081 26401 13093 26404
rect 13127 26401 13139 26435
rect 13081 26395 13139 26401
rect 13262 26392 13268 26444
rect 13320 26432 13326 26444
rect 13722 26432 13728 26444
rect 13320 26404 13728 26432
rect 13320 26392 13326 26404
rect 13722 26392 13728 26404
rect 13780 26392 13786 26444
rect 13814 26392 13820 26444
rect 13872 26432 13878 26444
rect 14277 26435 14335 26441
rect 14277 26432 14289 26435
rect 13872 26404 14289 26432
rect 13872 26392 13878 26404
rect 14277 26401 14289 26404
rect 14323 26401 14335 26435
rect 15102 26432 15108 26444
rect 15063 26404 15108 26432
rect 14277 26395 14335 26401
rect 15102 26392 15108 26404
rect 15160 26392 15166 26444
rect 15304 26441 15332 26472
rect 15289 26435 15347 26441
rect 15289 26401 15301 26435
rect 15335 26401 15347 26435
rect 16114 26432 16120 26444
rect 16075 26404 16120 26432
rect 15289 26395 15347 26401
rect 16114 26392 16120 26404
rect 16172 26392 16178 26444
rect 11388 26336 12756 26364
rect 11388 26324 11394 26336
rect 12802 26324 12808 26376
rect 12860 26364 12866 26376
rect 12860 26336 12905 26364
rect 12860 26324 12866 26336
rect 13170 26324 13176 26376
rect 13228 26364 13234 26376
rect 14093 26367 14151 26373
rect 14093 26364 14105 26367
rect 13228 26336 14105 26364
rect 13228 26324 13234 26336
rect 14093 26333 14105 26336
rect 14139 26333 14151 26367
rect 16224 26364 16252 26540
rect 18506 26528 18512 26540
rect 18564 26528 18570 26580
rect 19245 26571 19303 26577
rect 19245 26537 19257 26571
rect 19291 26537 19303 26571
rect 19245 26531 19303 26537
rect 21729 26571 21787 26577
rect 21729 26537 21741 26571
rect 21775 26568 21787 26571
rect 22094 26568 22100 26580
rect 21775 26540 22100 26568
rect 21775 26537 21787 26540
rect 21729 26531 21787 26537
rect 19260 26500 19288 26531
rect 22094 26528 22100 26540
rect 22152 26528 22158 26580
rect 25590 26528 25596 26580
rect 25648 26568 25654 26580
rect 25648 26540 28304 26568
rect 25648 26528 25654 26540
rect 22186 26500 22192 26512
rect 17512 26472 19288 26500
rect 19720 26472 22192 26500
rect 16301 26435 16359 26441
rect 16301 26401 16313 26435
rect 16347 26432 16359 26435
rect 16390 26432 16396 26444
rect 16347 26404 16396 26432
rect 16347 26401 16359 26404
rect 16301 26395 16359 26401
rect 16390 26392 16396 26404
rect 16448 26392 16454 26444
rect 17126 26392 17132 26444
rect 17184 26432 17190 26444
rect 17512 26441 17540 26472
rect 17497 26435 17555 26441
rect 17497 26432 17509 26435
rect 17184 26404 17509 26432
rect 17184 26392 17190 26404
rect 17497 26401 17509 26404
rect 17543 26401 17555 26435
rect 17497 26395 17555 26401
rect 17862 26392 17868 26444
rect 17920 26432 17926 26444
rect 18049 26435 18107 26441
rect 18049 26432 18061 26435
rect 17920 26404 18061 26432
rect 17920 26392 17926 26404
rect 18049 26401 18061 26404
rect 18095 26401 18107 26435
rect 18049 26395 18107 26401
rect 18138 26392 18144 26444
rect 18196 26432 18202 26444
rect 18233 26435 18291 26441
rect 18233 26432 18245 26435
rect 18196 26404 18245 26432
rect 18196 26392 18202 26404
rect 18233 26401 18245 26404
rect 18279 26432 18291 26435
rect 18782 26432 18788 26444
rect 18279 26404 18788 26432
rect 18279 26401 18291 26404
rect 18233 26395 18291 26401
rect 18782 26392 18788 26404
rect 18840 26392 18846 26444
rect 19150 26432 19156 26444
rect 19111 26404 19156 26432
rect 19150 26392 19156 26404
rect 19208 26392 19214 26444
rect 19720 26441 19748 26472
rect 22186 26460 22192 26472
rect 22244 26500 22250 26512
rect 26878 26500 26884 26512
rect 22244 26472 24624 26500
rect 22244 26460 22250 26472
rect 19705 26435 19763 26441
rect 19705 26401 19717 26435
rect 19751 26401 19763 26435
rect 19705 26395 19763 26401
rect 20806 26392 20812 26444
rect 20864 26432 20870 26444
rect 20901 26435 20959 26441
rect 20901 26432 20913 26435
rect 20864 26404 20913 26432
rect 20864 26392 20870 26404
rect 20901 26401 20913 26404
rect 20947 26401 20959 26435
rect 21634 26432 21640 26444
rect 21595 26404 21640 26432
rect 20901 26395 20959 26401
rect 21634 26392 21640 26404
rect 21692 26392 21698 26444
rect 22370 26432 22376 26444
rect 22331 26404 22376 26432
rect 22370 26392 22376 26404
rect 22428 26392 22434 26444
rect 22922 26432 22928 26444
rect 22883 26404 22928 26432
rect 22922 26392 22928 26404
rect 22980 26392 22986 26444
rect 23842 26432 23848 26444
rect 23803 26404 23848 26432
rect 23842 26392 23848 26404
rect 23900 26392 23906 26444
rect 24486 26432 24492 26444
rect 24447 26404 24492 26432
rect 24486 26392 24492 26404
rect 24544 26392 24550 26444
rect 17313 26367 17371 26373
rect 17313 26364 17325 26367
rect 16224 26336 17325 26364
rect 14093 26327 14151 26333
rect 17313 26333 17325 26336
rect 17359 26333 17371 26367
rect 23106 26364 23112 26376
rect 23067 26336 23112 26364
rect 17313 26327 17371 26333
rect 23106 26324 23112 26336
rect 23164 26324 23170 26376
rect 23566 26324 23572 26376
rect 23624 26364 23630 26376
rect 24596 26373 24624 26472
rect 25516 26472 26884 26500
rect 25133 26435 25191 26441
rect 25133 26401 25145 26435
rect 25179 26432 25191 26435
rect 25314 26432 25320 26444
rect 25179 26404 25320 26432
rect 25179 26401 25191 26404
rect 25133 26395 25191 26401
rect 25314 26392 25320 26404
rect 25372 26392 25378 26444
rect 25516 26441 25544 26472
rect 26878 26460 26884 26472
rect 26936 26460 26942 26512
rect 25501 26435 25559 26441
rect 25501 26401 25513 26435
rect 25547 26401 25559 26435
rect 25774 26432 25780 26444
rect 25735 26404 25780 26432
rect 25501 26395 25559 26401
rect 25774 26392 25780 26404
rect 25832 26392 25838 26444
rect 26513 26435 26571 26441
rect 26513 26401 26525 26435
rect 26559 26432 26571 26435
rect 28166 26432 28172 26444
rect 26559 26404 28172 26432
rect 26559 26401 26571 26404
rect 26513 26395 26571 26401
rect 28166 26392 28172 26404
rect 28224 26392 28230 26444
rect 24581 26367 24639 26373
rect 23624 26336 24532 26364
rect 23624 26324 23630 26336
rect 12618 26256 12624 26308
rect 12676 26256 12682 26308
rect 13630 26256 13636 26308
rect 13688 26296 13694 26308
rect 15194 26296 15200 26308
rect 13688 26268 15200 26296
rect 13688 26256 13694 26268
rect 15194 26256 15200 26268
rect 15252 26256 15258 26308
rect 16393 26299 16451 26305
rect 16393 26265 16405 26299
rect 16439 26296 16451 26299
rect 22557 26299 22615 26305
rect 16439 26268 21312 26296
rect 16439 26265 16451 26268
rect 16393 26259 16451 26265
rect 5350 26228 5356 26240
rect 4080 26200 5356 26228
rect 5350 26188 5356 26200
rect 5408 26188 5414 26240
rect 11054 26188 11060 26240
rect 11112 26228 11118 26240
rect 12636 26228 12664 26256
rect 14918 26228 14924 26240
rect 11112 26200 12664 26228
rect 14879 26200 14924 26228
rect 11112 26188 11118 26200
rect 14918 26188 14924 26200
rect 14976 26188 14982 26240
rect 21082 26228 21088 26240
rect 21043 26200 21088 26228
rect 21082 26188 21088 26200
rect 21140 26188 21146 26240
rect 21284 26228 21312 26268
rect 22557 26265 22569 26299
rect 22603 26296 22615 26299
rect 23934 26296 23940 26308
rect 22603 26268 23796 26296
rect 23895 26268 23940 26296
rect 22603 26265 22615 26268
rect 22557 26259 22615 26265
rect 23290 26228 23296 26240
rect 21284 26200 23296 26228
rect 23290 26188 23296 26200
rect 23348 26188 23354 26240
rect 23768 26228 23796 26268
rect 23934 26256 23940 26268
rect 23992 26256 23998 26308
rect 24504 26296 24532 26336
rect 24581 26333 24593 26367
rect 24627 26333 24639 26367
rect 27246 26364 27252 26376
rect 24581 26327 24639 26333
rect 26620 26336 27252 26364
rect 26620 26308 26648 26336
rect 27246 26324 27252 26336
rect 27304 26324 27310 26376
rect 27525 26367 27583 26373
rect 27525 26333 27537 26367
rect 27571 26364 27583 26367
rect 27614 26364 27620 26376
rect 27571 26336 27620 26364
rect 27571 26333 27583 26336
rect 27525 26327 27583 26333
rect 27614 26324 27620 26336
rect 27672 26324 27678 26376
rect 26602 26296 26608 26308
rect 24504 26268 26608 26296
rect 26602 26256 26608 26268
rect 26660 26256 26666 26308
rect 26697 26299 26755 26305
rect 26697 26265 26709 26299
rect 26743 26296 26755 26299
rect 28276 26296 28304 26540
rect 28626 26528 28632 26580
rect 28684 26568 28690 26580
rect 29733 26571 29791 26577
rect 29733 26568 29745 26571
rect 28684 26540 29745 26568
rect 28684 26528 28690 26540
rect 29733 26537 29745 26540
rect 29779 26537 29791 26571
rect 31478 26568 31484 26580
rect 31439 26540 31484 26568
rect 29733 26531 29791 26537
rect 31478 26528 31484 26540
rect 31536 26528 31542 26580
rect 37829 26571 37887 26577
rect 32968 26540 35020 26568
rect 28350 26460 28356 26512
rect 28408 26500 28414 26512
rect 31202 26500 31208 26512
rect 28408 26472 31208 26500
rect 28408 26460 28414 26472
rect 31202 26460 31208 26472
rect 31260 26460 31266 26512
rect 32968 26500 32996 26540
rect 31404 26472 32996 26500
rect 33045 26503 33103 26509
rect 29546 26392 29552 26444
rect 29604 26432 29610 26444
rect 31404 26441 31432 26472
rect 33045 26469 33057 26503
rect 33091 26500 33103 26503
rect 33134 26500 33140 26512
rect 33091 26472 33140 26500
rect 33091 26469 33103 26472
rect 33045 26463 33103 26469
rect 33134 26460 33140 26472
rect 33192 26460 33198 26512
rect 34992 26500 35020 26540
rect 37829 26537 37841 26571
rect 37875 26568 37887 26571
rect 37918 26568 37924 26580
rect 37875 26540 37924 26568
rect 37875 26537 37887 26540
rect 37829 26531 37887 26537
rect 37918 26528 37924 26540
rect 37976 26528 37982 26580
rect 38470 26568 38476 26580
rect 38431 26540 38476 26568
rect 38470 26528 38476 26540
rect 38528 26528 38534 26580
rect 38654 26500 38660 26512
rect 34992 26472 38660 26500
rect 38654 26460 38660 26472
rect 38712 26460 38718 26512
rect 29641 26435 29699 26441
rect 29641 26432 29653 26435
rect 29604 26404 29653 26432
rect 29604 26392 29610 26404
rect 29641 26401 29653 26404
rect 29687 26401 29699 26435
rect 29641 26395 29699 26401
rect 30193 26435 30251 26441
rect 30193 26401 30205 26435
rect 30239 26401 30251 26435
rect 30193 26395 30251 26401
rect 31389 26435 31447 26441
rect 31389 26401 31401 26435
rect 31435 26401 31447 26435
rect 31389 26395 31447 26401
rect 29362 26324 29368 26376
rect 29420 26364 29426 26376
rect 30208 26364 30236 26395
rect 32030 26392 32036 26444
rect 32088 26432 32094 26444
rect 32309 26435 32367 26441
rect 32309 26432 32321 26435
rect 32088 26404 32321 26432
rect 32088 26392 32094 26404
rect 32309 26401 32321 26404
rect 32355 26401 32367 26435
rect 32309 26395 32367 26401
rect 32861 26435 32919 26441
rect 32861 26401 32873 26435
rect 32907 26432 32919 26435
rect 33778 26432 33784 26444
rect 32907 26404 33640 26432
rect 33739 26404 33784 26432
rect 32907 26401 32919 26404
rect 32861 26395 32919 26401
rect 29420 26336 30236 26364
rect 30653 26367 30711 26373
rect 29420 26324 29426 26336
rect 30653 26333 30665 26367
rect 30699 26364 30711 26367
rect 30742 26364 30748 26376
rect 30699 26336 30748 26364
rect 30699 26333 30711 26336
rect 30653 26327 30711 26333
rect 30742 26324 30748 26336
rect 30800 26324 30806 26376
rect 32324 26364 32352 26395
rect 33318 26364 33324 26376
rect 32324 26336 33324 26364
rect 33318 26324 33324 26336
rect 33376 26324 33382 26376
rect 33502 26364 33508 26376
rect 33463 26336 33508 26364
rect 33502 26324 33508 26336
rect 33560 26324 33566 26376
rect 33612 26364 33640 26404
rect 33778 26392 33784 26404
rect 33836 26392 33842 26444
rect 35986 26432 35992 26444
rect 35947 26404 35992 26432
rect 35986 26392 35992 26404
rect 36044 26432 36050 26444
rect 36262 26432 36268 26444
rect 36044 26404 36268 26432
rect 36044 26392 36050 26404
rect 36262 26392 36268 26404
rect 36320 26392 36326 26444
rect 36357 26435 36415 26441
rect 36357 26401 36369 26435
rect 36403 26401 36415 26435
rect 36357 26395 36415 26401
rect 37001 26435 37059 26441
rect 37001 26401 37013 26435
rect 37047 26401 37059 26435
rect 37734 26432 37740 26444
rect 37695 26404 37740 26432
rect 37001 26395 37059 26401
rect 35161 26367 35219 26373
rect 35161 26364 35173 26367
rect 33612 26336 35173 26364
rect 35161 26333 35173 26336
rect 35207 26364 35219 26367
rect 35342 26364 35348 26376
rect 35207 26336 35348 26364
rect 35207 26333 35219 26336
rect 35161 26327 35219 26333
rect 35342 26324 35348 26336
rect 35400 26324 35406 26376
rect 35710 26324 35716 26376
rect 35768 26364 35774 26376
rect 36372 26364 36400 26395
rect 35768 26336 36400 26364
rect 37016 26364 37044 26395
rect 37734 26392 37740 26404
rect 37792 26432 37798 26444
rect 38378 26432 38384 26444
rect 37792 26404 38384 26432
rect 37792 26392 37798 26404
rect 38378 26392 38384 26404
rect 38436 26392 38442 26444
rect 38565 26435 38623 26441
rect 38565 26401 38577 26435
rect 38611 26432 38623 26435
rect 38746 26432 38752 26444
rect 38611 26404 38752 26432
rect 38611 26401 38623 26404
rect 38565 26395 38623 26401
rect 38746 26392 38752 26404
rect 38804 26392 38810 26444
rect 38933 26435 38991 26441
rect 38933 26401 38945 26435
rect 38979 26432 38991 26435
rect 39945 26435 40003 26441
rect 39945 26432 39957 26435
rect 38979 26404 39957 26432
rect 38979 26401 38991 26404
rect 38933 26395 38991 26401
rect 39945 26401 39957 26404
rect 39991 26401 40003 26435
rect 39945 26395 40003 26401
rect 38286 26364 38292 26376
rect 37016 26336 38292 26364
rect 35768 26324 35774 26336
rect 38286 26324 38292 26336
rect 38344 26324 38350 26376
rect 32490 26296 32496 26308
rect 26743 26268 27292 26296
rect 28276 26268 32496 26296
rect 26743 26265 26755 26268
rect 26697 26259 26755 26265
rect 24578 26228 24584 26240
rect 23768 26200 24584 26228
rect 24578 26188 24584 26200
rect 24636 26188 24642 26240
rect 27264 26228 27292 26268
rect 32490 26256 32496 26268
rect 32548 26256 32554 26308
rect 27706 26228 27712 26240
rect 27264 26200 27712 26228
rect 27706 26188 27712 26200
rect 27764 26188 27770 26240
rect 28166 26188 28172 26240
rect 28224 26228 28230 26240
rect 28629 26231 28687 26237
rect 28629 26228 28641 26231
rect 28224 26200 28641 26228
rect 28224 26188 28230 26200
rect 28629 26197 28641 26200
rect 28675 26197 28687 26231
rect 36078 26228 36084 26240
rect 36039 26200 36084 26228
rect 28629 26191 28687 26197
rect 36078 26188 36084 26200
rect 36136 26188 36142 26240
rect 1104 26138 39836 26160
rect 1104 26086 4246 26138
rect 4298 26086 4310 26138
rect 4362 26086 4374 26138
rect 4426 26086 4438 26138
rect 4490 26086 34966 26138
rect 35018 26086 35030 26138
rect 35082 26086 35094 26138
rect 35146 26086 35158 26138
rect 35210 26086 39836 26138
rect 1104 26064 39836 26086
rect 2682 25984 2688 26036
rect 2740 26024 2746 26036
rect 5442 26024 5448 26036
rect 2740 25996 5448 26024
rect 2740 25984 2746 25996
rect 5442 25984 5448 25996
rect 5500 25984 5506 26036
rect 9398 25984 9404 26036
rect 9456 26024 9462 26036
rect 9456 25996 10088 26024
rect 9456 25984 9462 25996
rect 3053 25959 3111 25965
rect 3053 25925 3065 25959
rect 3099 25956 3111 25959
rect 3602 25956 3608 25968
rect 3099 25928 3608 25956
rect 3099 25925 3111 25928
rect 3053 25919 3111 25925
rect 3602 25916 3608 25928
rect 3660 25916 3666 25968
rect 4062 25916 4068 25968
rect 4120 25956 4126 25968
rect 5902 25956 5908 25968
rect 4120 25928 5908 25956
rect 4120 25916 4126 25928
rect 5902 25916 5908 25928
rect 5960 25916 5966 25968
rect 9950 25956 9956 25968
rect 8220 25928 9956 25956
rect 2406 25888 2412 25900
rect 2367 25860 2412 25888
rect 2406 25848 2412 25860
rect 2464 25848 2470 25900
rect 5442 25848 5448 25900
rect 5500 25888 5506 25900
rect 5500 25860 5545 25888
rect 5500 25848 5506 25860
rect 7374 25848 7380 25900
rect 7432 25888 7438 25900
rect 8220 25897 8248 25928
rect 9950 25916 9956 25928
rect 10008 25916 10014 25968
rect 8205 25891 8263 25897
rect 8205 25888 8217 25891
rect 7432 25860 8217 25888
rect 7432 25848 7438 25860
rect 8205 25857 8217 25860
rect 8251 25857 8263 25891
rect 8205 25851 8263 25857
rect 8941 25891 8999 25897
rect 8941 25857 8953 25891
rect 8987 25888 8999 25891
rect 9858 25888 9864 25900
rect 8987 25860 9864 25888
rect 8987 25857 8999 25860
rect 8941 25851 8999 25857
rect 9858 25848 9864 25860
rect 9916 25848 9922 25900
rect 1762 25820 1768 25832
rect 1723 25792 1768 25820
rect 1762 25780 1768 25792
rect 1820 25780 1826 25832
rect 2314 25829 2320 25832
rect 2271 25823 2320 25829
rect 2271 25789 2283 25823
rect 2317 25789 2320 25823
rect 2271 25783 2320 25789
rect 2314 25780 2320 25783
rect 2372 25780 2378 25832
rect 2958 25780 2964 25832
rect 3016 25820 3022 25832
rect 3513 25823 3571 25829
rect 3513 25820 3525 25823
rect 3016 25792 3525 25820
rect 3016 25780 3022 25792
rect 3513 25789 3525 25792
rect 3559 25789 3571 25823
rect 3513 25783 3571 25789
rect 3602 25780 3608 25832
rect 3660 25820 3666 25832
rect 3973 25823 4031 25829
rect 3973 25820 3985 25823
rect 3660 25792 3985 25820
rect 3660 25780 3666 25792
rect 3973 25789 3985 25792
rect 4019 25789 4031 25823
rect 3973 25783 4031 25789
rect 4062 25780 4068 25832
rect 4120 25820 4126 25832
rect 4341 25823 4399 25829
rect 4341 25820 4353 25823
rect 4120 25792 4353 25820
rect 4120 25780 4126 25792
rect 4341 25789 4353 25792
rect 4387 25789 4399 25823
rect 4341 25783 4399 25789
rect 4709 25823 4767 25829
rect 4709 25789 4721 25823
rect 4755 25820 4767 25823
rect 5718 25820 5724 25832
rect 4755 25792 5724 25820
rect 4755 25789 4767 25792
rect 4709 25783 4767 25789
rect 3421 25755 3479 25761
rect 3421 25721 3433 25755
rect 3467 25752 3479 25755
rect 4614 25752 4620 25764
rect 3467 25724 4620 25752
rect 3467 25721 3479 25724
rect 3421 25715 3479 25721
rect 4614 25712 4620 25724
rect 4672 25712 4678 25764
rect 1581 25687 1639 25693
rect 1581 25653 1593 25687
rect 1627 25684 1639 25687
rect 1670 25684 1676 25696
rect 1627 25656 1676 25684
rect 1627 25653 1639 25656
rect 1581 25647 1639 25653
rect 1670 25644 1676 25656
rect 1728 25644 1734 25696
rect 3142 25644 3148 25696
rect 3200 25684 3206 25696
rect 4062 25684 4068 25696
rect 3200 25656 4068 25684
rect 3200 25644 3206 25656
rect 4062 25644 4068 25656
rect 4120 25684 4126 25696
rect 4724 25684 4752 25783
rect 5718 25780 5724 25792
rect 5776 25780 5782 25832
rect 6178 25820 6184 25832
rect 6139 25792 6184 25820
rect 6178 25780 6184 25792
rect 6236 25780 6242 25832
rect 7561 25823 7619 25829
rect 7561 25789 7573 25823
rect 7607 25820 7619 25823
rect 7742 25820 7748 25832
rect 7607 25792 7748 25820
rect 7607 25789 7619 25792
rect 7561 25783 7619 25789
rect 7742 25780 7748 25792
rect 7800 25780 7806 25832
rect 8110 25820 8116 25832
rect 8071 25792 8116 25820
rect 8110 25780 8116 25792
rect 8168 25780 8174 25832
rect 9490 25820 9496 25832
rect 9451 25792 9496 25820
rect 9490 25780 9496 25792
rect 9548 25780 9554 25832
rect 9769 25823 9827 25829
rect 9769 25789 9781 25823
rect 9815 25789 9827 25823
rect 9950 25820 9956 25832
rect 9911 25792 9956 25820
rect 9769 25783 9827 25789
rect 5813 25755 5871 25761
rect 5813 25752 5825 25755
rect 5552 25724 5825 25752
rect 4120 25656 4752 25684
rect 4120 25644 4126 25656
rect 5350 25644 5356 25696
rect 5408 25684 5414 25696
rect 5552 25684 5580 25724
rect 5813 25721 5825 25724
rect 5859 25721 5871 25755
rect 5813 25715 5871 25721
rect 9030 25712 9036 25764
rect 9088 25752 9094 25764
rect 9784 25752 9812 25783
rect 9950 25780 9956 25792
rect 10008 25780 10014 25832
rect 10060 25820 10088 25996
rect 10686 25984 10692 26036
rect 10744 26024 10750 26036
rect 11422 26024 11428 26036
rect 10744 25996 11428 26024
rect 10744 25984 10750 25996
rect 11422 25984 11428 25996
rect 11480 26024 11486 26036
rect 11480 25996 12480 26024
rect 11480 25984 11486 25996
rect 12452 25956 12480 25996
rect 14274 25984 14280 26036
rect 14332 26024 14338 26036
rect 14461 26027 14519 26033
rect 14461 26024 14473 26027
rect 14332 25996 14473 26024
rect 14332 25984 14338 25996
rect 14461 25993 14473 25996
rect 14507 25993 14519 26027
rect 14461 25987 14519 25993
rect 16485 26027 16543 26033
rect 16485 25993 16497 26027
rect 16531 26024 16543 26027
rect 16574 26024 16580 26036
rect 16531 25996 16580 26024
rect 16531 25993 16543 25996
rect 16485 25987 16543 25993
rect 16574 25984 16580 25996
rect 16632 25984 16638 26036
rect 18322 26024 18328 26036
rect 18283 25996 18328 26024
rect 18322 25984 18328 25996
rect 18380 25984 18386 26036
rect 22554 25984 22560 26036
rect 22612 26024 22618 26036
rect 23017 26027 23075 26033
rect 23017 26024 23029 26027
rect 22612 25996 23029 26024
rect 22612 25984 22618 25996
rect 23017 25993 23029 25996
rect 23063 25993 23075 26027
rect 23017 25987 23075 25993
rect 23566 25984 23572 26036
rect 23624 26024 23630 26036
rect 25590 26024 25596 26036
rect 23624 25996 25596 26024
rect 23624 25984 23630 25996
rect 25590 25984 25596 25996
rect 25648 25984 25654 26036
rect 33318 26024 33324 26036
rect 33279 25996 33324 26024
rect 33318 25984 33324 25996
rect 33376 26024 33382 26036
rect 34238 26024 34244 26036
rect 33376 25996 34244 26024
rect 33376 25984 33382 25996
rect 34238 25984 34244 25996
rect 34296 25984 34302 26036
rect 36262 25984 36268 26036
rect 36320 26024 36326 26036
rect 36541 26027 36599 26033
rect 36541 26024 36553 26027
rect 36320 25996 36553 26024
rect 36320 25984 36326 25996
rect 36541 25993 36553 25996
rect 36587 25993 36599 26027
rect 38654 26024 38660 26036
rect 38615 25996 38660 26024
rect 36541 25987 36599 25993
rect 38654 25984 38660 25996
rect 38712 25984 38718 26036
rect 20901 25959 20959 25965
rect 20901 25956 20913 25959
rect 12452 25928 15424 25956
rect 10594 25848 10600 25900
rect 10652 25888 10658 25900
rect 15396 25897 15424 25928
rect 16960 25928 20913 25956
rect 15381 25891 15439 25897
rect 10652 25860 11468 25888
rect 10652 25848 10658 25860
rect 10873 25823 10931 25829
rect 10873 25820 10885 25823
rect 10060 25792 10885 25820
rect 10873 25789 10885 25792
rect 10919 25789 10931 25823
rect 10873 25783 10931 25789
rect 11057 25823 11115 25829
rect 11057 25789 11069 25823
rect 11103 25789 11115 25823
rect 11330 25820 11336 25832
rect 11291 25792 11336 25820
rect 11057 25783 11115 25789
rect 9088 25724 9812 25752
rect 10413 25755 10471 25761
rect 9088 25712 9094 25724
rect 10413 25721 10425 25755
rect 10459 25752 10471 25755
rect 10962 25752 10968 25764
rect 10459 25724 10968 25752
rect 10459 25721 10471 25724
rect 10413 25715 10471 25721
rect 10962 25712 10968 25724
rect 11020 25712 11026 25764
rect 5408 25656 5580 25684
rect 5629 25687 5687 25693
rect 5408 25644 5414 25656
rect 5629 25653 5641 25687
rect 5675 25684 5687 25687
rect 5902 25684 5908 25696
rect 5675 25656 5908 25684
rect 5675 25653 5687 25656
rect 5629 25647 5687 25653
rect 5902 25644 5908 25656
rect 5960 25644 5966 25696
rect 7469 25687 7527 25693
rect 7469 25653 7481 25687
rect 7515 25684 7527 25687
rect 7650 25684 7656 25696
rect 7515 25656 7656 25684
rect 7515 25653 7527 25656
rect 7469 25647 7527 25653
rect 7650 25644 7656 25656
rect 7708 25644 7714 25696
rect 8846 25644 8852 25696
rect 8904 25684 8910 25696
rect 11072 25684 11100 25783
rect 11330 25780 11336 25792
rect 11388 25780 11394 25832
rect 11440 25829 11468 25860
rect 15381 25857 15393 25891
rect 15427 25857 15439 25891
rect 15381 25851 15439 25857
rect 11425 25823 11483 25829
rect 11425 25789 11437 25823
rect 11471 25789 11483 25823
rect 11425 25783 11483 25789
rect 11793 25823 11851 25829
rect 11793 25789 11805 25823
rect 11839 25820 11851 25823
rect 12434 25820 12440 25832
rect 11839 25792 12440 25820
rect 11839 25789 11851 25792
rect 11793 25783 11851 25789
rect 12434 25780 12440 25792
rect 12492 25780 12498 25832
rect 13354 25820 13360 25832
rect 13315 25792 13360 25820
rect 13354 25780 13360 25792
rect 13412 25780 13418 25832
rect 13630 25820 13636 25832
rect 13591 25792 13636 25820
rect 13630 25780 13636 25792
rect 13688 25780 13694 25832
rect 13814 25820 13820 25832
rect 13775 25792 13820 25820
rect 13814 25780 13820 25792
rect 13872 25780 13878 25832
rect 14274 25820 14280 25832
rect 14235 25792 14280 25820
rect 14274 25780 14280 25792
rect 14332 25780 14338 25832
rect 15473 25823 15531 25829
rect 15473 25789 15485 25823
rect 15519 25789 15531 25823
rect 15473 25783 15531 25789
rect 16025 25823 16083 25829
rect 16025 25789 16037 25823
rect 16071 25820 16083 25823
rect 16114 25820 16120 25832
rect 16071 25792 16120 25820
rect 16071 25789 16083 25792
rect 16025 25783 16083 25789
rect 12805 25755 12863 25761
rect 12805 25721 12817 25755
rect 12851 25752 12863 25755
rect 13906 25752 13912 25764
rect 12851 25724 13912 25752
rect 12851 25721 12863 25724
rect 12805 25715 12863 25721
rect 13906 25712 13912 25724
rect 13964 25712 13970 25764
rect 15488 25752 15516 25783
rect 16114 25780 16120 25792
rect 16172 25780 16178 25832
rect 16209 25823 16267 25829
rect 16209 25789 16221 25823
rect 16255 25820 16267 25823
rect 16390 25820 16396 25832
rect 16255 25792 16396 25820
rect 16255 25789 16267 25792
rect 16209 25783 16267 25789
rect 16390 25780 16396 25792
rect 16448 25820 16454 25832
rect 16960 25820 16988 25928
rect 20901 25925 20913 25928
rect 20947 25956 20959 25959
rect 25222 25956 25228 25968
rect 20947 25928 23888 25956
rect 25183 25928 25228 25956
rect 20947 25925 20959 25928
rect 20901 25919 20959 25925
rect 20070 25888 20076 25900
rect 19720 25860 20076 25888
rect 17126 25820 17132 25832
rect 16448 25792 16988 25820
rect 17087 25792 17132 25820
rect 16448 25780 16454 25792
rect 17126 25780 17132 25792
rect 17184 25780 17190 25832
rect 17954 25780 17960 25832
rect 18012 25820 18018 25832
rect 18049 25823 18107 25829
rect 18049 25820 18061 25823
rect 18012 25792 18061 25820
rect 18012 25780 18018 25792
rect 18049 25789 18061 25792
rect 18095 25789 18107 25823
rect 18049 25783 18107 25789
rect 18138 25780 18144 25832
rect 18196 25829 18202 25832
rect 18196 25823 18251 25829
rect 18196 25789 18205 25823
rect 18239 25789 18251 25823
rect 18196 25783 18251 25789
rect 18196 25780 18202 25783
rect 18322 25780 18328 25832
rect 18380 25820 18386 25832
rect 19720 25829 19748 25860
rect 20070 25848 20076 25860
rect 20128 25848 20134 25900
rect 20257 25891 20315 25897
rect 20257 25857 20269 25891
rect 20303 25888 20315 25891
rect 23860 25888 23888 25928
rect 25222 25916 25228 25928
rect 25280 25916 25286 25968
rect 29917 25959 29975 25965
rect 29917 25925 29929 25959
rect 29963 25956 29975 25959
rect 30098 25956 30104 25968
rect 29963 25928 30104 25956
rect 29963 25925 29975 25928
rect 29917 25919 29975 25925
rect 30098 25916 30104 25928
rect 30156 25916 30162 25968
rect 26970 25888 26976 25900
rect 20303 25860 23796 25888
rect 23860 25860 25636 25888
rect 20303 25857 20315 25860
rect 20257 25851 20315 25857
rect 19153 25823 19211 25829
rect 19153 25820 19165 25823
rect 18380 25792 19165 25820
rect 18380 25780 18386 25792
rect 19153 25789 19165 25792
rect 19199 25789 19211 25823
rect 19153 25783 19211 25789
rect 19705 25823 19763 25829
rect 19705 25789 19717 25823
rect 19751 25789 19763 25823
rect 19978 25820 19984 25832
rect 19939 25792 19984 25820
rect 19705 25783 19763 25789
rect 19978 25780 19984 25792
rect 20036 25780 20042 25832
rect 20714 25820 20720 25832
rect 20675 25792 20720 25820
rect 20714 25780 20720 25792
rect 20772 25780 20778 25832
rect 22002 25820 22008 25832
rect 21963 25792 22008 25820
rect 22002 25780 22008 25792
rect 22060 25780 22066 25832
rect 22278 25820 22284 25832
rect 22239 25792 22284 25820
rect 22278 25780 22284 25792
rect 22336 25780 22342 25832
rect 22646 25780 22652 25832
rect 22704 25820 22710 25832
rect 22925 25823 22983 25829
rect 22925 25820 22937 25823
rect 22704 25792 22937 25820
rect 22704 25780 22710 25792
rect 22925 25789 22937 25792
rect 22971 25789 22983 25823
rect 22925 25783 22983 25789
rect 23566 25780 23572 25832
rect 23624 25820 23630 25832
rect 23661 25823 23719 25829
rect 23661 25820 23673 25823
rect 23624 25792 23673 25820
rect 23624 25780 23630 25792
rect 23661 25789 23673 25792
rect 23707 25789 23719 25823
rect 23768 25820 23796 25860
rect 24213 25823 24271 25829
rect 23768 25792 24072 25820
rect 23661 25783 23719 25789
rect 15654 25752 15660 25764
rect 15488 25724 15660 25752
rect 15654 25712 15660 25724
rect 15712 25752 15718 25764
rect 18156 25752 18184 25780
rect 20732 25752 20760 25780
rect 15712 25724 17356 25752
rect 18156 25724 20760 25752
rect 22465 25755 22523 25761
rect 15712 25712 15718 25724
rect 17328 25696 17356 25724
rect 22465 25721 22477 25755
rect 22511 25752 22523 25755
rect 22554 25752 22560 25764
rect 22511 25724 22560 25752
rect 22511 25721 22523 25724
rect 22465 25715 22523 25721
rect 22554 25712 22560 25724
rect 22612 25712 22618 25764
rect 11974 25684 11980 25696
rect 8904 25656 11980 25684
rect 8904 25644 8910 25656
rect 11974 25644 11980 25656
rect 12032 25684 12038 25696
rect 12250 25684 12256 25696
rect 12032 25656 12256 25684
rect 12032 25644 12038 25656
rect 12250 25644 12256 25656
rect 12308 25644 12314 25696
rect 17310 25684 17316 25696
rect 17271 25656 17316 25684
rect 17310 25644 17316 25656
rect 17368 25644 17374 25696
rect 23842 25644 23848 25696
rect 23900 25684 23906 25696
rect 23937 25687 23995 25693
rect 23937 25684 23949 25687
rect 23900 25656 23949 25684
rect 23900 25644 23906 25656
rect 23937 25653 23949 25656
rect 23983 25653 23995 25687
rect 24044 25684 24072 25792
rect 24213 25789 24225 25823
rect 24259 25820 24271 25823
rect 24578 25820 24584 25832
rect 24259 25792 24584 25820
rect 24259 25789 24271 25792
rect 24213 25783 24271 25789
rect 24578 25780 24584 25792
rect 24636 25780 24642 25832
rect 25406 25820 25412 25832
rect 25367 25792 25412 25820
rect 25406 25780 25412 25792
rect 25464 25780 25470 25832
rect 25608 25829 25636 25860
rect 25792 25860 26976 25888
rect 25792 25829 25820 25860
rect 26970 25848 26976 25860
rect 27028 25888 27034 25900
rect 31389 25891 31447 25897
rect 27028 25860 27108 25888
rect 27028 25848 27034 25860
rect 25593 25823 25651 25829
rect 25593 25789 25605 25823
rect 25639 25789 25651 25823
rect 25593 25783 25651 25789
rect 25777 25823 25835 25829
rect 25777 25789 25789 25823
rect 25823 25789 25835 25823
rect 25777 25783 25835 25789
rect 25958 25780 25964 25832
rect 26016 25820 26022 25832
rect 27080 25829 27108 25860
rect 31389 25857 31401 25891
rect 31435 25888 31447 25891
rect 32217 25891 32275 25897
rect 32217 25888 32229 25891
rect 31435 25860 32229 25888
rect 31435 25857 31447 25860
rect 31389 25851 31447 25857
rect 32217 25857 32229 25860
rect 32263 25857 32275 25891
rect 32217 25851 32275 25857
rect 33502 25848 33508 25900
rect 33560 25888 33566 25900
rect 35161 25891 35219 25897
rect 35161 25888 35173 25891
rect 33560 25860 35173 25888
rect 33560 25848 33566 25860
rect 35161 25857 35173 25860
rect 35207 25888 35219 25891
rect 37274 25888 37280 25900
rect 35207 25860 37280 25888
rect 35207 25857 35219 25860
rect 35161 25851 35219 25857
rect 37274 25848 37280 25860
rect 37332 25848 37338 25900
rect 26881 25823 26939 25829
rect 26881 25820 26893 25823
rect 26016 25792 26893 25820
rect 26016 25780 26022 25792
rect 26881 25789 26893 25792
rect 26927 25789 26939 25823
rect 26881 25783 26939 25789
rect 27065 25823 27123 25829
rect 27065 25789 27077 25823
rect 27111 25789 27123 25823
rect 27246 25820 27252 25832
rect 27207 25792 27252 25820
rect 27065 25783 27123 25789
rect 27246 25780 27252 25792
rect 27304 25780 27310 25832
rect 28166 25820 28172 25832
rect 28127 25792 28172 25820
rect 28166 25780 28172 25792
rect 28224 25780 28230 25832
rect 28258 25780 28264 25832
rect 28316 25820 28322 25832
rect 28353 25823 28411 25829
rect 28353 25820 28365 25823
rect 28316 25792 28365 25820
rect 28316 25780 28322 25792
rect 28353 25789 28365 25792
rect 28399 25789 28411 25823
rect 28353 25783 28411 25789
rect 29546 25780 29552 25832
rect 29604 25820 29610 25832
rect 29641 25823 29699 25829
rect 29641 25820 29653 25823
rect 29604 25792 29653 25820
rect 29604 25780 29610 25792
rect 29641 25789 29653 25792
rect 29687 25789 29699 25823
rect 29641 25783 29699 25789
rect 30193 25823 30251 25829
rect 30193 25789 30205 25823
rect 30239 25789 30251 25823
rect 30558 25820 30564 25832
rect 30519 25792 30564 25820
rect 30193 25783 30251 25789
rect 25038 25712 25044 25764
rect 25096 25752 25102 25764
rect 26421 25755 26479 25761
rect 26421 25752 26433 25755
rect 25096 25724 26433 25752
rect 25096 25712 25102 25724
rect 26421 25721 26433 25724
rect 26467 25721 26479 25755
rect 30208 25752 30236 25783
rect 30558 25780 30564 25792
rect 30616 25780 30622 25832
rect 31297 25823 31355 25829
rect 31297 25789 31309 25823
rect 31343 25789 31355 25823
rect 31297 25783 31355 25789
rect 31941 25823 31999 25829
rect 31941 25789 31953 25823
rect 31987 25820 31999 25823
rect 33520 25820 33548 25848
rect 31987 25792 33548 25820
rect 31987 25789 31999 25792
rect 31941 25783 31999 25789
rect 26421 25715 26479 25721
rect 26528 25724 30236 25752
rect 31312 25752 31340 25783
rect 33870 25780 33876 25832
rect 33928 25820 33934 25832
rect 34054 25820 34060 25832
rect 33928 25792 34060 25820
rect 33928 25780 33934 25792
rect 34054 25780 34060 25792
rect 34112 25780 34118 25832
rect 35434 25820 35440 25832
rect 35395 25792 35440 25820
rect 35434 25780 35440 25792
rect 35492 25780 35498 25832
rect 37550 25820 37556 25832
rect 37511 25792 37556 25820
rect 37550 25780 37556 25792
rect 37608 25780 37614 25832
rect 31312 25724 31800 25752
rect 26528 25684 26556 25724
rect 24044 25656 26556 25684
rect 23937 25647 23995 25653
rect 26878 25644 26884 25696
rect 26936 25684 26942 25696
rect 27985 25687 28043 25693
rect 27985 25684 27997 25687
rect 26936 25656 27997 25684
rect 26936 25644 26942 25656
rect 27985 25653 27997 25656
rect 28031 25653 28043 25687
rect 31772 25684 31800 25724
rect 33962 25684 33968 25696
rect 31772 25656 33968 25684
rect 27985 25647 28043 25653
rect 33962 25644 33968 25656
rect 34020 25644 34026 25696
rect 34241 25687 34299 25693
rect 34241 25653 34253 25687
rect 34287 25684 34299 25687
rect 35802 25684 35808 25696
rect 34287 25656 35808 25684
rect 34287 25653 34299 25656
rect 34241 25647 34299 25653
rect 35802 25644 35808 25656
rect 35860 25684 35866 25696
rect 37918 25684 37924 25696
rect 35860 25656 37924 25684
rect 35860 25644 35866 25656
rect 37918 25644 37924 25656
rect 37976 25644 37982 25696
rect 1104 25594 39836 25616
rect 1104 25542 19606 25594
rect 19658 25542 19670 25594
rect 19722 25542 19734 25594
rect 19786 25542 19798 25594
rect 19850 25542 39836 25594
rect 1104 25520 39836 25542
rect 5718 25480 5724 25492
rect 5679 25452 5724 25480
rect 5718 25440 5724 25452
rect 5776 25440 5782 25492
rect 8110 25440 8116 25492
rect 8168 25480 8174 25492
rect 9030 25480 9036 25492
rect 8168 25452 9036 25480
rect 8168 25440 8174 25452
rect 9030 25440 9036 25452
rect 9088 25440 9094 25492
rect 9490 25440 9496 25492
rect 9548 25480 9554 25492
rect 9769 25483 9827 25489
rect 9769 25480 9781 25483
rect 9548 25452 9781 25480
rect 9548 25440 9554 25452
rect 9769 25449 9781 25452
rect 9815 25449 9827 25483
rect 9769 25443 9827 25449
rect 9950 25440 9956 25492
rect 10008 25480 10014 25492
rect 10594 25480 10600 25492
rect 10008 25452 10600 25480
rect 10008 25440 10014 25452
rect 10594 25440 10600 25452
rect 10652 25440 10658 25492
rect 11054 25440 11060 25492
rect 11112 25480 11118 25492
rect 11238 25480 11244 25492
rect 11112 25452 11244 25480
rect 11112 25440 11118 25452
rect 11238 25440 11244 25452
rect 11296 25480 11302 25492
rect 11517 25483 11575 25489
rect 11517 25480 11529 25483
rect 11296 25452 11529 25480
rect 11296 25440 11302 25452
rect 11517 25449 11529 25452
rect 11563 25449 11575 25483
rect 18046 25480 18052 25492
rect 11517 25443 11575 25449
rect 15488 25452 18052 25480
rect 4065 25415 4123 25421
rect 4065 25381 4077 25415
rect 4111 25412 4123 25415
rect 4706 25412 4712 25424
rect 4111 25384 4712 25412
rect 4111 25381 4123 25384
rect 4065 25375 4123 25381
rect 4706 25372 4712 25384
rect 4764 25372 4770 25424
rect 5736 25412 5764 25440
rect 5092 25384 5764 25412
rect 9048 25412 9076 25440
rect 9048 25384 10272 25412
rect 1397 25347 1455 25353
rect 1397 25313 1409 25347
rect 1443 25344 1455 25347
rect 1486 25344 1492 25356
rect 1443 25316 1492 25344
rect 1443 25313 1455 25316
rect 1397 25307 1455 25313
rect 1486 25304 1492 25316
rect 1544 25304 1550 25356
rect 1670 25344 1676 25356
rect 1631 25316 1676 25344
rect 1670 25304 1676 25316
rect 1728 25304 1734 25356
rect 4614 25344 4620 25356
rect 4575 25316 4620 25344
rect 4614 25304 4620 25316
rect 4672 25304 4678 25356
rect 4798 25304 4804 25356
rect 4856 25344 4862 25356
rect 5092 25353 5120 25384
rect 4893 25347 4951 25353
rect 4893 25344 4905 25347
rect 4856 25316 4905 25344
rect 4856 25304 4862 25316
rect 4893 25313 4905 25316
rect 4939 25313 4951 25347
rect 4893 25307 4951 25313
rect 5077 25347 5135 25353
rect 5077 25313 5089 25347
rect 5123 25313 5135 25347
rect 5077 25307 5135 25313
rect 5537 25347 5595 25353
rect 5537 25313 5549 25347
rect 5583 25344 5595 25347
rect 5626 25344 5632 25356
rect 5583 25316 5632 25344
rect 5583 25313 5595 25316
rect 5537 25307 5595 25313
rect 5626 25304 5632 25316
rect 5684 25304 5690 25356
rect 6546 25344 6552 25356
rect 6507 25316 6552 25344
rect 6546 25304 6552 25316
rect 6604 25304 6610 25356
rect 8846 25344 8852 25356
rect 8807 25316 8852 25344
rect 8846 25304 8852 25316
rect 8904 25304 8910 25356
rect 9858 25344 9864 25356
rect 9819 25316 9864 25344
rect 9858 25304 9864 25316
rect 9916 25304 9922 25356
rect 10244 25353 10272 25384
rect 11146 25372 11152 25424
rect 11204 25412 11210 25424
rect 11609 25415 11667 25421
rect 11609 25412 11621 25415
rect 11204 25384 11621 25412
rect 11204 25372 11210 25384
rect 11609 25381 11621 25384
rect 11655 25381 11667 25415
rect 11609 25375 11667 25381
rect 11701 25415 11759 25421
rect 11701 25381 11713 25415
rect 11747 25381 11759 25415
rect 11701 25375 11759 25381
rect 12069 25415 12127 25421
rect 12069 25381 12081 25415
rect 12115 25412 12127 25415
rect 14274 25412 14280 25424
rect 12115 25384 14280 25412
rect 12115 25381 12127 25384
rect 12069 25375 12127 25381
rect 10229 25347 10287 25353
rect 10229 25313 10241 25347
rect 10275 25313 10287 25347
rect 10594 25344 10600 25356
rect 10555 25316 10600 25344
rect 10229 25307 10287 25313
rect 10594 25304 10600 25316
rect 10652 25304 10658 25356
rect 11716 25344 11744 25375
rect 14274 25372 14280 25384
rect 14332 25372 14338 25424
rect 12434 25344 12440 25356
rect 11716 25316 12440 25344
rect 12434 25304 12440 25316
rect 12492 25344 12498 25356
rect 12802 25344 12808 25356
rect 12492 25316 12808 25344
rect 12492 25304 12498 25316
rect 12802 25304 12808 25316
rect 12860 25304 12866 25356
rect 13262 25344 13268 25356
rect 13223 25316 13268 25344
rect 13262 25304 13268 25316
rect 13320 25304 13326 25356
rect 13633 25347 13691 25353
rect 13633 25313 13645 25347
rect 13679 25313 13691 25347
rect 13633 25307 13691 25313
rect 14001 25347 14059 25353
rect 14001 25313 14013 25347
rect 14047 25344 14059 25347
rect 14182 25344 14188 25356
rect 14047 25316 14188 25344
rect 14047 25313 14059 25316
rect 14001 25307 14059 25313
rect 6825 25279 6883 25285
rect 6825 25245 6837 25279
rect 6871 25276 6883 25279
rect 6914 25276 6920 25288
rect 6871 25248 6920 25276
rect 6871 25245 6883 25248
rect 6825 25239 6883 25245
rect 6914 25236 6920 25248
rect 6972 25236 6978 25288
rect 7742 25236 7748 25288
rect 7800 25276 7806 25288
rect 8205 25279 8263 25285
rect 8205 25276 8217 25279
rect 7800 25248 8217 25276
rect 7800 25236 7806 25248
rect 8205 25245 8217 25248
rect 8251 25276 8263 25279
rect 10686 25276 10692 25288
rect 8251 25248 10692 25276
rect 8251 25245 8263 25248
rect 8205 25239 8263 25245
rect 10686 25236 10692 25248
rect 10744 25236 10750 25288
rect 11054 25236 11060 25288
rect 11112 25276 11118 25288
rect 11333 25279 11391 25285
rect 11333 25276 11345 25279
rect 11112 25248 11345 25276
rect 11112 25236 11118 25248
rect 11333 25245 11345 25248
rect 11379 25245 11391 25279
rect 13446 25276 13452 25288
rect 13407 25248 13452 25276
rect 11333 25239 11391 25245
rect 13446 25236 13452 25248
rect 13504 25236 13510 25288
rect 13648 25276 13676 25307
rect 14182 25304 14188 25316
rect 14240 25304 14246 25356
rect 15488 25353 15516 25452
rect 18046 25440 18052 25452
rect 18104 25480 18110 25492
rect 34054 25480 34060 25492
rect 18104 25452 19196 25480
rect 18104 25440 18110 25452
rect 18322 25412 18328 25424
rect 18283 25384 18328 25412
rect 18322 25372 18328 25384
rect 18380 25372 18386 25424
rect 19168 25356 19196 25452
rect 32508 25452 34060 25480
rect 20349 25415 20407 25421
rect 19812 25384 20300 25412
rect 15473 25347 15531 25353
rect 15473 25313 15485 25347
rect 15519 25313 15531 25347
rect 15473 25307 15531 25313
rect 16114 25304 16120 25356
rect 16172 25344 16178 25356
rect 16209 25347 16267 25353
rect 16209 25344 16221 25347
rect 16172 25316 16221 25344
rect 16172 25304 16178 25316
rect 16209 25313 16221 25316
rect 16255 25313 16267 25347
rect 16209 25307 16267 25313
rect 17221 25347 17279 25353
rect 17221 25313 17233 25347
rect 17267 25344 17279 25347
rect 17310 25344 17316 25356
rect 17267 25316 17316 25344
rect 17267 25313 17279 25316
rect 17221 25307 17279 25313
rect 17310 25304 17316 25316
rect 17368 25304 17374 25356
rect 17773 25347 17831 25353
rect 17773 25313 17785 25347
rect 17819 25344 17831 25347
rect 17862 25344 17868 25356
rect 17819 25316 17868 25344
rect 17819 25313 17831 25316
rect 17773 25307 17831 25313
rect 17862 25304 17868 25316
rect 17920 25304 17926 25356
rect 17957 25347 18015 25353
rect 17957 25313 17969 25347
rect 18003 25344 18015 25347
rect 18138 25344 18144 25356
rect 18003 25316 18144 25344
rect 18003 25313 18015 25316
rect 17957 25307 18015 25313
rect 18138 25304 18144 25316
rect 18196 25304 18202 25356
rect 19150 25344 19156 25356
rect 19063 25316 19156 25344
rect 19150 25304 19156 25316
rect 19208 25304 19214 25356
rect 19812 25353 19840 25384
rect 19797 25347 19855 25353
rect 19797 25313 19809 25347
rect 19843 25313 19855 25347
rect 19797 25307 19855 25313
rect 20165 25347 20223 25353
rect 20165 25313 20177 25347
rect 20211 25313 20223 25347
rect 20272 25344 20300 25384
rect 20349 25381 20361 25415
rect 20395 25412 20407 25415
rect 20714 25412 20720 25424
rect 20395 25384 20720 25412
rect 20395 25381 20407 25384
rect 20349 25375 20407 25381
rect 20714 25372 20720 25384
rect 20772 25372 20778 25424
rect 22002 25412 22008 25424
rect 21963 25384 22008 25412
rect 22002 25372 22008 25384
rect 22060 25372 22066 25424
rect 23934 25412 23940 25424
rect 23032 25384 23940 25412
rect 20898 25344 20904 25356
rect 20272 25316 20904 25344
rect 20165 25307 20223 25313
rect 13814 25276 13820 25288
rect 13648 25248 13820 25276
rect 13814 25236 13820 25248
rect 13872 25276 13878 25288
rect 15654 25276 15660 25288
rect 13872 25248 15660 25276
rect 13872 25236 13878 25248
rect 15654 25236 15660 25248
rect 15712 25276 15718 25288
rect 17037 25279 17095 25285
rect 17037 25276 17049 25279
rect 15712 25248 17049 25276
rect 15712 25236 15718 25248
rect 17037 25245 17049 25248
rect 17083 25245 17095 25279
rect 20180 25276 20208 25307
rect 20898 25304 20904 25316
rect 20956 25304 20962 25356
rect 21082 25304 21088 25356
rect 21140 25344 21146 25356
rect 21269 25347 21327 25353
rect 21269 25344 21281 25347
rect 21140 25316 21281 25344
rect 21140 25304 21146 25316
rect 21269 25313 21281 25316
rect 21315 25313 21327 25347
rect 21818 25344 21824 25356
rect 21779 25316 21824 25344
rect 21269 25307 21327 25313
rect 21818 25304 21824 25316
rect 21876 25304 21882 25356
rect 23032 25353 23060 25384
rect 23934 25372 23940 25384
rect 23992 25372 23998 25424
rect 28258 25412 28264 25424
rect 28219 25384 28264 25412
rect 28258 25372 28264 25384
rect 28316 25372 28322 25424
rect 31481 25415 31539 25421
rect 31481 25381 31493 25415
rect 31527 25412 31539 25415
rect 32398 25412 32404 25424
rect 31527 25384 32404 25412
rect 31527 25381 31539 25384
rect 31481 25375 31539 25381
rect 32398 25372 32404 25384
rect 32456 25372 32462 25424
rect 23017 25347 23075 25353
rect 23017 25313 23029 25347
rect 23063 25313 23075 25347
rect 23290 25344 23296 25356
rect 23251 25316 23296 25344
rect 23017 25307 23075 25313
rect 23290 25304 23296 25316
rect 23348 25304 23354 25356
rect 23750 25344 23756 25356
rect 23711 25316 23756 25344
rect 23750 25304 23756 25316
rect 23808 25304 23814 25356
rect 23842 25304 23848 25356
rect 23900 25344 23906 25356
rect 24213 25347 24271 25353
rect 24213 25344 24225 25347
rect 23900 25316 24225 25344
rect 23900 25304 23906 25316
rect 24213 25313 24225 25316
rect 24259 25313 24271 25347
rect 25038 25344 25044 25356
rect 24999 25316 25044 25344
rect 24213 25307 24271 25313
rect 25038 25304 25044 25316
rect 25096 25304 25102 25356
rect 25222 25304 25228 25356
rect 25280 25344 25286 25356
rect 25409 25347 25467 25353
rect 25409 25344 25421 25347
rect 25280 25316 25421 25344
rect 25280 25304 25286 25316
rect 25409 25313 25421 25316
rect 25455 25313 25467 25347
rect 26602 25344 26608 25356
rect 26563 25316 26608 25344
rect 25409 25307 25467 25313
rect 26602 25304 26608 25316
rect 26660 25304 26666 25356
rect 27246 25304 27252 25356
rect 27304 25344 27310 25356
rect 29181 25347 29239 25353
rect 29181 25344 29193 25347
rect 27304 25316 29193 25344
rect 27304 25304 27310 25316
rect 29181 25313 29193 25316
rect 29227 25313 29239 25347
rect 29546 25344 29552 25356
rect 29507 25316 29552 25344
rect 29181 25307 29239 25313
rect 29546 25304 29552 25316
rect 29604 25304 29610 25356
rect 30377 25347 30435 25353
rect 30377 25313 30389 25347
rect 30423 25313 30435 25347
rect 30558 25344 30564 25356
rect 30519 25316 30564 25344
rect 30377 25307 30435 25313
rect 20806 25276 20812 25288
rect 20180 25248 20812 25276
rect 17037 25239 17095 25245
rect 20806 25236 20812 25248
rect 20864 25276 20870 25288
rect 22002 25276 22008 25288
rect 20864 25248 22008 25276
rect 20864 25236 20870 25248
rect 22002 25236 22008 25248
rect 22060 25236 22066 25288
rect 25866 25276 25872 25288
rect 25827 25248 25872 25276
rect 25866 25236 25872 25248
rect 25924 25236 25930 25288
rect 26881 25279 26939 25285
rect 26881 25245 26893 25279
rect 26927 25276 26939 25279
rect 28166 25276 28172 25288
rect 26927 25248 28172 25276
rect 26927 25245 26939 25248
rect 26881 25239 26939 25245
rect 28166 25236 28172 25248
rect 28224 25236 28230 25288
rect 28350 25236 28356 25288
rect 28408 25276 28414 25288
rect 28721 25279 28779 25285
rect 28721 25276 28733 25279
rect 28408 25248 28733 25276
rect 28408 25236 28414 25248
rect 28721 25245 28733 25248
rect 28767 25245 28779 25279
rect 29638 25276 29644 25288
rect 29599 25248 29644 25276
rect 28721 25239 28779 25245
rect 29638 25236 29644 25248
rect 29696 25236 29702 25288
rect 18874 25208 18880 25220
rect 15672 25180 18880 25208
rect 2774 25100 2780 25152
rect 2832 25140 2838 25152
rect 15672 25149 15700 25180
rect 18874 25168 18880 25180
rect 18932 25168 18938 25220
rect 22554 25168 22560 25220
rect 22612 25208 22618 25220
rect 23109 25211 23167 25217
rect 23109 25208 23121 25211
rect 22612 25180 23121 25208
rect 22612 25168 22618 25180
rect 23109 25177 23121 25180
rect 23155 25208 23167 25211
rect 24946 25208 24952 25220
rect 23155 25180 24808 25208
rect 24907 25180 24952 25208
rect 23155 25177 23167 25180
rect 23109 25171 23167 25177
rect 15657 25143 15715 25149
rect 2832 25112 2877 25140
rect 2832 25100 2838 25112
rect 15657 25109 15669 25143
rect 15703 25109 15715 25143
rect 15657 25103 15715 25109
rect 16393 25143 16451 25149
rect 16393 25109 16405 25143
rect 16439 25140 16451 25143
rect 16666 25140 16672 25152
rect 16439 25112 16672 25140
rect 16439 25109 16451 25112
rect 16393 25103 16451 25109
rect 16666 25100 16672 25112
rect 16724 25140 16730 25152
rect 16942 25140 16948 25152
rect 16724 25112 16948 25140
rect 16724 25100 16730 25112
rect 16942 25100 16948 25112
rect 17000 25100 17006 25152
rect 17034 25100 17040 25152
rect 17092 25140 17098 25152
rect 17310 25140 17316 25152
rect 17092 25112 17316 25140
rect 17092 25100 17098 25112
rect 17310 25100 17316 25112
rect 17368 25100 17374 25152
rect 22186 25100 22192 25152
rect 22244 25140 22250 25152
rect 24305 25143 24363 25149
rect 24305 25140 24317 25143
rect 22244 25112 24317 25140
rect 22244 25100 22250 25112
rect 24305 25109 24317 25112
rect 24351 25140 24363 25143
rect 24486 25140 24492 25152
rect 24351 25112 24492 25140
rect 24351 25109 24363 25112
rect 24305 25103 24363 25109
rect 24486 25100 24492 25112
rect 24544 25100 24550 25152
rect 24780 25140 24808 25180
rect 24946 25168 24952 25180
rect 25004 25168 25010 25220
rect 30392 25208 30420 25307
rect 30558 25304 30564 25316
rect 30616 25304 30622 25356
rect 30742 25344 30748 25356
rect 30703 25316 30748 25344
rect 30742 25304 30748 25316
rect 30800 25304 30806 25356
rect 31389 25347 31447 25353
rect 31389 25313 31401 25347
rect 31435 25344 31447 25347
rect 31846 25344 31852 25356
rect 31435 25316 31852 25344
rect 31435 25313 31447 25316
rect 31389 25307 31447 25313
rect 31846 25304 31852 25316
rect 31904 25304 31910 25356
rect 32309 25347 32367 25353
rect 32309 25313 32321 25347
rect 32355 25344 32367 25347
rect 32508 25344 32536 25452
rect 34054 25440 34060 25452
rect 34112 25440 34118 25492
rect 35434 25480 35440 25492
rect 35395 25452 35440 25480
rect 35434 25440 35440 25452
rect 35492 25440 35498 25492
rect 32674 25344 32680 25356
rect 32355 25316 32536 25344
rect 32635 25316 32680 25344
rect 32355 25313 32367 25316
rect 32309 25307 32367 25313
rect 32674 25304 32680 25316
rect 32732 25344 32738 25356
rect 32732 25316 33088 25344
rect 32732 25304 32738 25316
rect 32490 25236 32496 25288
rect 32548 25276 32554 25288
rect 32953 25279 33011 25285
rect 32953 25276 32965 25279
rect 32548 25248 32965 25276
rect 32548 25236 32554 25248
rect 32953 25245 32965 25248
rect 32999 25245 33011 25279
rect 33060 25276 33088 25316
rect 33134 25304 33140 25356
rect 33192 25344 33198 25356
rect 34057 25347 34115 25353
rect 34057 25344 34069 25347
rect 33192 25316 34069 25344
rect 33192 25304 33198 25316
rect 34057 25313 34069 25316
rect 34103 25313 34115 25347
rect 34057 25307 34115 25313
rect 34517 25347 34575 25353
rect 34517 25313 34529 25347
rect 34563 25313 34575 25347
rect 35526 25344 35532 25356
rect 35487 25316 35532 25344
rect 34517 25307 34575 25313
rect 33781 25279 33839 25285
rect 33781 25276 33793 25279
rect 33060 25248 33793 25276
rect 32953 25239 33011 25245
rect 33781 25245 33793 25248
rect 33827 25245 33839 25279
rect 34532 25276 34560 25307
rect 35526 25304 35532 25316
rect 35584 25304 35590 25356
rect 36078 25344 36084 25356
rect 36039 25316 36084 25344
rect 36078 25304 36084 25316
rect 36136 25304 36142 25356
rect 36909 25347 36967 25353
rect 36909 25313 36921 25347
rect 36955 25313 36967 25347
rect 36909 25307 36967 25313
rect 38197 25347 38255 25353
rect 38197 25313 38209 25347
rect 38243 25344 38255 25347
rect 38470 25344 38476 25356
rect 38243 25316 38476 25344
rect 38243 25313 38255 25316
rect 38197 25307 38255 25313
rect 33781 25239 33839 25245
rect 33888 25248 34560 25276
rect 32401 25211 32459 25217
rect 30392 25180 32352 25208
rect 25498 25140 25504 25152
rect 24780 25112 25504 25140
rect 25498 25100 25504 25112
rect 25556 25140 25562 25152
rect 30742 25140 30748 25152
rect 25556 25112 30748 25140
rect 25556 25100 25562 25112
rect 30742 25100 30748 25112
rect 30800 25100 30806 25152
rect 32324 25140 32352 25180
rect 32401 25177 32413 25211
rect 32447 25208 32459 25211
rect 33888 25208 33916 25248
rect 35894 25236 35900 25288
rect 35952 25276 35958 25288
rect 36173 25279 36231 25285
rect 36173 25276 36185 25279
rect 35952 25248 36185 25276
rect 35952 25236 35958 25248
rect 36173 25245 36185 25248
rect 36219 25245 36231 25279
rect 36924 25276 36952 25307
rect 38470 25304 38476 25316
rect 38528 25304 38534 25356
rect 38746 25344 38752 25356
rect 38659 25316 38752 25344
rect 38746 25304 38752 25316
rect 38804 25344 38810 25356
rect 39114 25344 39120 25356
rect 38804 25316 39120 25344
rect 38804 25304 38810 25316
rect 39114 25304 39120 25316
rect 39172 25304 39178 25356
rect 37734 25276 37740 25288
rect 36924 25248 37740 25276
rect 36173 25239 36231 25245
rect 37734 25236 37740 25248
rect 37792 25276 37798 25288
rect 38378 25276 38384 25288
rect 37792 25248 38384 25276
rect 37792 25236 37798 25248
rect 38378 25236 38384 25248
rect 38436 25236 38442 25288
rect 38838 25276 38844 25288
rect 38799 25248 38844 25276
rect 38838 25236 38844 25248
rect 38896 25236 38902 25288
rect 32447 25180 33916 25208
rect 32447 25177 32459 25180
rect 32401 25171 32459 25177
rect 33962 25168 33968 25220
rect 34020 25208 34026 25220
rect 34517 25211 34575 25217
rect 34517 25208 34529 25211
rect 34020 25180 34529 25208
rect 34020 25168 34026 25180
rect 34517 25177 34529 25180
rect 34563 25177 34575 25211
rect 38286 25208 38292 25220
rect 38247 25180 38292 25208
rect 34517 25171 34575 25177
rect 38286 25168 38292 25180
rect 38344 25168 38350 25220
rect 36078 25140 36084 25152
rect 32324 25112 36084 25140
rect 36078 25100 36084 25112
rect 36136 25100 36142 25152
rect 37090 25140 37096 25152
rect 37051 25112 37096 25140
rect 37090 25100 37096 25112
rect 37148 25100 37154 25152
rect 1104 25050 39836 25072
rect 1104 24998 4246 25050
rect 4298 24998 4310 25050
rect 4362 24998 4374 25050
rect 4426 24998 4438 25050
rect 4490 24998 34966 25050
rect 35018 24998 35030 25050
rect 35082 24998 35094 25050
rect 35146 24998 35158 25050
rect 35210 24998 39836 25050
rect 1104 24976 39836 24998
rect 19613 24939 19671 24945
rect 19613 24905 19625 24939
rect 19659 24936 19671 24939
rect 22738 24936 22744 24948
rect 19659 24908 22744 24936
rect 19659 24905 19671 24908
rect 19613 24899 19671 24905
rect 22738 24896 22744 24908
rect 22796 24896 22802 24948
rect 23842 24936 23848 24948
rect 23803 24908 23848 24936
rect 23842 24896 23848 24908
rect 23900 24896 23906 24948
rect 23934 24896 23940 24948
rect 23992 24936 23998 24948
rect 27982 24936 27988 24948
rect 23992 24908 27988 24936
rect 23992 24896 23998 24908
rect 27982 24896 27988 24908
rect 28040 24896 28046 24948
rect 2317 24871 2375 24877
rect 2317 24837 2329 24871
rect 2363 24868 2375 24871
rect 2406 24868 2412 24880
rect 2363 24840 2412 24868
rect 2363 24837 2375 24840
rect 2317 24831 2375 24837
rect 2406 24828 2412 24840
rect 2464 24828 2470 24880
rect 5718 24828 5724 24880
rect 5776 24868 5782 24880
rect 5997 24871 6055 24877
rect 5997 24868 6009 24871
rect 5776 24840 6009 24868
rect 5776 24828 5782 24840
rect 5997 24837 6009 24840
rect 6043 24837 6055 24871
rect 20346 24868 20352 24880
rect 20307 24840 20352 24868
rect 5997 24831 6055 24837
rect 20346 24828 20352 24840
rect 20404 24828 20410 24880
rect 21085 24871 21143 24877
rect 21085 24837 21097 24871
rect 21131 24837 21143 24871
rect 21085 24831 21143 24837
rect 3970 24800 3976 24812
rect 3712 24772 3976 24800
rect 3712 24744 3740 24772
rect 3970 24760 3976 24772
rect 4028 24760 4034 24812
rect 7558 24800 7564 24812
rect 6104 24772 7564 24800
rect 2501 24735 2559 24741
rect 2501 24701 2513 24735
rect 2547 24732 2559 24735
rect 2774 24732 2780 24744
rect 2547 24704 2780 24732
rect 2547 24701 2559 24704
rect 2501 24695 2559 24701
rect 2774 24692 2780 24704
rect 2832 24692 2838 24744
rect 2958 24732 2964 24744
rect 2919 24704 2964 24732
rect 2958 24692 2964 24704
rect 3016 24692 3022 24744
rect 3234 24732 3240 24744
rect 3195 24704 3240 24732
rect 3234 24692 3240 24704
rect 3292 24732 3298 24744
rect 3602 24732 3608 24744
rect 3292 24704 3608 24732
rect 3292 24692 3298 24704
rect 3602 24692 3608 24704
rect 3660 24692 3666 24744
rect 3694 24692 3700 24744
rect 3752 24732 3758 24744
rect 4062 24732 4068 24744
rect 3752 24704 3797 24732
rect 4023 24704 4068 24732
rect 3752 24692 3758 24704
rect 4062 24692 4068 24704
rect 4120 24692 4126 24744
rect 5353 24735 5411 24741
rect 5353 24701 5365 24735
rect 5399 24732 5411 24735
rect 5626 24732 5632 24744
rect 5399 24704 5632 24732
rect 5399 24701 5411 24704
rect 5353 24695 5411 24701
rect 5626 24692 5632 24704
rect 5684 24692 5690 24744
rect 6104 24741 6132 24772
rect 7558 24760 7564 24772
rect 7616 24760 7622 24812
rect 7745 24803 7803 24809
rect 7745 24769 7757 24803
rect 7791 24800 7803 24803
rect 7926 24800 7932 24812
rect 7791 24772 7932 24800
rect 7791 24769 7803 24772
rect 7745 24763 7803 24769
rect 7926 24760 7932 24772
rect 7984 24800 7990 24812
rect 11333 24803 11391 24809
rect 11333 24800 11345 24803
rect 7984 24772 11345 24800
rect 7984 24760 7990 24772
rect 11333 24769 11345 24772
rect 11379 24769 11391 24803
rect 11333 24763 11391 24769
rect 13173 24803 13231 24809
rect 13173 24769 13185 24803
rect 13219 24800 13231 24803
rect 13630 24800 13636 24812
rect 13219 24772 13636 24800
rect 13219 24769 13231 24772
rect 13173 24763 13231 24769
rect 13630 24760 13636 24772
rect 13688 24760 13694 24812
rect 15654 24800 15660 24812
rect 15615 24772 15660 24800
rect 15654 24760 15660 24772
rect 15712 24760 15718 24812
rect 19150 24760 19156 24812
rect 19208 24800 19214 24812
rect 20530 24800 20536 24812
rect 19208 24772 20536 24800
rect 19208 24760 19214 24772
rect 5721 24735 5779 24741
rect 5721 24701 5733 24735
rect 5767 24701 5779 24735
rect 5721 24695 5779 24701
rect 6089 24735 6147 24741
rect 6089 24701 6101 24735
rect 6135 24701 6147 24735
rect 7098 24732 7104 24744
rect 7059 24704 7104 24732
rect 6089 24695 6147 24701
rect 5736 24664 5764 24695
rect 7098 24692 7104 24704
rect 7156 24692 7162 24744
rect 7650 24732 7656 24744
rect 7611 24704 7656 24732
rect 7650 24692 7656 24704
rect 7708 24692 7714 24744
rect 8481 24735 8539 24741
rect 8481 24701 8493 24735
rect 8527 24701 8539 24735
rect 8754 24732 8760 24744
rect 8715 24704 8760 24732
rect 8481 24695 8539 24701
rect 6178 24664 6184 24676
rect 5736 24636 6184 24664
rect 6178 24624 6184 24636
rect 6236 24624 6242 24676
rect 6914 24596 6920 24608
rect 6875 24568 6920 24596
rect 6914 24556 6920 24568
rect 6972 24556 6978 24608
rect 8496 24596 8524 24695
rect 8754 24692 8760 24704
rect 8812 24692 8818 24744
rect 10597 24735 10655 24741
rect 10597 24701 10609 24735
rect 10643 24732 10655 24735
rect 11054 24732 11060 24744
rect 10643 24704 11060 24732
rect 10643 24701 10655 24704
rect 10597 24695 10655 24701
rect 11054 24692 11060 24704
rect 11112 24692 11118 24744
rect 11238 24692 11244 24744
rect 11296 24732 11302 24744
rect 12713 24735 12771 24741
rect 12713 24732 12725 24735
rect 11296 24704 12725 24732
rect 11296 24692 11302 24704
rect 12713 24701 12725 24704
rect 12759 24701 12771 24735
rect 12713 24695 12771 24701
rect 13538 24692 13544 24744
rect 13596 24732 13602 24744
rect 13998 24732 14004 24744
rect 13596 24704 14004 24732
rect 13596 24692 13602 24704
rect 13998 24692 14004 24704
rect 14056 24692 14062 24744
rect 14277 24735 14335 24741
rect 14277 24701 14289 24735
rect 14323 24732 14335 24735
rect 15378 24732 15384 24744
rect 14323 24704 15384 24732
rect 14323 24701 14335 24704
rect 14277 24695 14335 24701
rect 15378 24692 15384 24704
rect 15436 24692 15442 24744
rect 16669 24735 16727 24741
rect 16669 24701 16681 24735
rect 16715 24732 16727 24735
rect 18322 24732 18328 24744
rect 16715 24704 18328 24732
rect 16715 24701 16727 24704
rect 16669 24695 16727 24701
rect 18322 24692 18328 24704
rect 18380 24692 18386 24744
rect 19444 24741 19472 24772
rect 20530 24760 20536 24772
rect 20588 24800 20594 24812
rect 21100 24800 21128 24831
rect 21910 24828 21916 24880
rect 21968 24868 21974 24880
rect 22830 24868 22836 24880
rect 21968 24840 22836 24868
rect 21968 24828 21974 24840
rect 22830 24828 22836 24840
rect 22888 24868 22894 24880
rect 22925 24871 22983 24877
rect 22925 24868 22937 24871
rect 22888 24840 22937 24868
rect 22888 24828 22894 24840
rect 22925 24837 22937 24840
rect 22971 24837 22983 24871
rect 22925 24831 22983 24837
rect 29454 24828 29460 24880
rect 29512 24828 29518 24880
rect 20588 24772 21128 24800
rect 20588 24760 20594 24772
rect 21818 24760 21824 24812
rect 21876 24800 21882 24812
rect 21876 24772 22784 24800
rect 21876 24760 21882 24772
rect 18601 24735 18659 24741
rect 18601 24701 18613 24735
rect 18647 24701 18659 24735
rect 18601 24695 18659 24701
rect 19429 24735 19487 24741
rect 19429 24701 19441 24735
rect 19475 24701 19487 24735
rect 20162 24732 20168 24744
rect 20075 24704 20168 24732
rect 19429 24695 19487 24701
rect 10137 24667 10195 24673
rect 10137 24633 10149 24667
rect 10183 24664 10195 24667
rect 10965 24667 11023 24673
rect 10965 24664 10977 24667
rect 10183 24636 10977 24664
rect 10183 24633 10195 24636
rect 10137 24627 10195 24633
rect 10965 24633 10977 24636
rect 11011 24664 11023 24667
rect 11146 24664 11152 24676
rect 11011 24636 11152 24664
rect 11011 24633 11023 24636
rect 10965 24627 11023 24633
rect 11146 24624 11152 24636
rect 11204 24624 11210 24676
rect 11974 24624 11980 24676
rect 12032 24664 12038 24676
rect 12437 24667 12495 24673
rect 12437 24664 12449 24667
rect 12032 24636 12449 24664
rect 12032 24624 12038 24636
rect 12437 24633 12449 24636
rect 12483 24633 12495 24667
rect 12802 24664 12808 24676
rect 12763 24636 12808 24664
rect 12437 24627 12495 24633
rect 12802 24624 12808 24636
rect 12860 24624 12866 24676
rect 16574 24624 16580 24676
rect 16632 24664 16638 24676
rect 18616 24664 18644 24695
rect 20162 24692 20168 24704
rect 20220 24732 20226 24744
rect 20901 24735 20959 24741
rect 20220 24704 20300 24732
rect 20220 24692 20226 24704
rect 19150 24664 19156 24676
rect 16632 24636 19156 24664
rect 16632 24624 16638 24636
rect 19150 24624 19156 24636
rect 19208 24624 19214 24676
rect 20272 24664 20300 24704
rect 20901 24701 20913 24735
rect 20947 24732 20959 24735
rect 21726 24732 21732 24744
rect 20947 24704 21732 24732
rect 20947 24701 20959 24704
rect 20901 24695 20959 24701
rect 21726 24692 21732 24704
rect 21784 24692 21790 24744
rect 22005 24735 22063 24741
rect 22005 24701 22017 24735
rect 22051 24732 22063 24735
rect 22646 24732 22652 24744
rect 22051 24704 22652 24732
rect 22051 24701 22063 24704
rect 22005 24695 22063 24701
rect 22646 24692 22652 24704
rect 22704 24692 22710 24744
rect 22756 24741 22784 24772
rect 23474 24760 23480 24812
rect 23532 24800 23538 24812
rect 24489 24803 24547 24809
rect 24489 24800 24501 24803
rect 23532 24772 24501 24800
rect 23532 24760 23538 24772
rect 24489 24769 24501 24772
rect 24535 24769 24547 24803
rect 24489 24763 24547 24769
rect 24765 24803 24823 24809
rect 24765 24769 24777 24803
rect 24811 24800 24823 24803
rect 24946 24800 24952 24812
rect 24811 24772 24952 24800
rect 24811 24769 24823 24772
rect 24765 24763 24823 24769
rect 24946 24760 24952 24772
rect 25004 24760 25010 24812
rect 25774 24760 25780 24812
rect 25832 24800 25838 24812
rect 25869 24803 25927 24809
rect 25869 24800 25881 24803
rect 25832 24772 25881 24800
rect 25832 24760 25838 24772
rect 25869 24769 25881 24772
rect 25915 24769 25927 24803
rect 25869 24763 25927 24769
rect 26510 24760 26516 24812
rect 26568 24800 26574 24812
rect 27246 24800 27252 24812
rect 26568 24772 27252 24800
rect 26568 24760 26574 24772
rect 27246 24760 27252 24772
rect 27304 24800 27310 24812
rect 27433 24803 27491 24809
rect 27433 24800 27445 24803
rect 27304 24772 27445 24800
rect 27304 24760 27310 24772
rect 27433 24769 27445 24772
rect 27479 24769 27491 24803
rect 29472 24800 29500 24828
rect 27433 24763 27491 24769
rect 27540 24772 29500 24800
rect 29549 24803 29607 24809
rect 22741 24735 22799 24741
rect 22741 24701 22753 24735
rect 22787 24701 22799 24735
rect 22741 24695 22799 24701
rect 23661 24735 23719 24741
rect 23661 24701 23673 24735
rect 23707 24732 23719 24735
rect 24394 24732 24400 24744
rect 23707 24704 24400 24732
rect 23707 24701 23719 24704
rect 23661 24695 23719 24701
rect 24394 24692 24400 24704
rect 24452 24692 24458 24744
rect 24578 24692 24584 24744
rect 24636 24732 24642 24744
rect 26605 24735 26663 24741
rect 26605 24732 26617 24735
rect 24636 24704 26617 24732
rect 24636 24692 24642 24704
rect 26605 24701 26617 24704
rect 26651 24701 26663 24735
rect 27540 24732 27568 24772
rect 29549 24769 29561 24803
rect 29595 24800 29607 24803
rect 30558 24800 30564 24812
rect 29595 24772 30564 24800
rect 29595 24769 29607 24772
rect 29549 24763 29607 24769
rect 30558 24760 30564 24772
rect 30616 24760 30622 24812
rect 30653 24803 30711 24809
rect 30653 24769 30665 24803
rect 30699 24800 30711 24803
rect 31018 24800 31024 24812
rect 30699 24772 31024 24800
rect 30699 24769 30711 24772
rect 30653 24763 30711 24769
rect 31018 24760 31024 24772
rect 31076 24760 31082 24812
rect 33045 24803 33103 24809
rect 33045 24769 33057 24803
rect 33091 24800 33103 24803
rect 33134 24800 33140 24812
rect 33091 24772 33140 24800
rect 33091 24769 33103 24772
rect 33045 24763 33103 24769
rect 33134 24760 33140 24772
rect 33192 24760 33198 24812
rect 35253 24803 35311 24809
rect 35253 24769 35265 24803
rect 35299 24800 35311 24803
rect 35894 24800 35900 24812
rect 35299 24772 35900 24800
rect 35299 24769 35311 24772
rect 35253 24763 35311 24769
rect 35894 24760 35900 24772
rect 35952 24760 35958 24812
rect 36725 24803 36783 24809
rect 36725 24769 36737 24803
rect 36771 24800 36783 24803
rect 37550 24800 37556 24812
rect 36771 24772 37556 24800
rect 36771 24769 36783 24772
rect 36725 24763 36783 24769
rect 37550 24760 37556 24772
rect 37608 24760 37614 24812
rect 26605 24695 26663 24701
rect 26804 24704 27568 24732
rect 27709 24735 27767 24741
rect 20272 24636 22232 24664
rect 9674 24596 9680 24608
rect 8496 24568 9680 24596
rect 9674 24556 9680 24568
rect 9732 24596 9738 24608
rect 9950 24596 9956 24608
rect 9732 24568 9956 24596
rect 9732 24556 9738 24568
rect 9950 24556 9956 24568
rect 10008 24556 10014 24608
rect 10686 24556 10692 24608
rect 10744 24596 10750 24608
rect 10781 24599 10839 24605
rect 10781 24596 10793 24599
rect 10744 24568 10793 24596
rect 10744 24556 10750 24568
rect 10781 24565 10793 24568
rect 10827 24565 10839 24599
rect 10781 24559 10839 24565
rect 10873 24599 10931 24605
rect 10873 24565 10885 24599
rect 10919 24596 10931 24599
rect 11238 24596 11244 24608
rect 10919 24568 11244 24596
rect 10919 24565 10931 24568
rect 10873 24559 10931 24565
rect 11238 24556 11244 24568
rect 11296 24556 11302 24608
rect 11330 24556 11336 24608
rect 11388 24596 11394 24608
rect 12621 24599 12679 24605
rect 12621 24596 12633 24599
rect 11388 24568 12633 24596
rect 11388 24556 11394 24568
rect 12621 24565 12633 24568
rect 12667 24596 12679 24599
rect 13262 24596 13268 24608
rect 12667 24568 13268 24596
rect 12667 24565 12679 24568
rect 12621 24559 12679 24565
rect 13262 24556 13268 24568
rect 13320 24556 13326 24608
rect 16114 24556 16120 24608
rect 16172 24596 16178 24608
rect 16853 24599 16911 24605
rect 16853 24596 16865 24599
rect 16172 24568 16865 24596
rect 16172 24556 16178 24568
rect 16853 24565 16865 24568
rect 16899 24565 16911 24599
rect 18782 24596 18788 24608
rect 18743 24568 18788 24596
rect 16853 24559 16911 24565
rect 18782 24556 18788 24568
rect 18840 24556 18846 24608
rect 22204 24605 22232 24636
rect 26804 24605 26832 24704
rect 27709 24701 27721 24735
rect 27755 24701 27767 24735
rect 28169 24735 28227 24741
rect 28169 24732 28181 24735
rect 27709 24695 27767 24701
rect 27816 24704 28181 24732
rect 26878 24624 26884 24676
rect 26936 24664 26942 24676
rect 27724 24664 27752 24695
rect 26936 24636 27752 24664
rect 26936 24624 26942 24636
rect 22189 24599 22247 24605
rect 22189 24565 22201 24599
rect 22235 24565 22247 24599
rect 22189 24559 22247 24565
rect 26789 24599 26847 24605
rect 26789 24565 26801 24599
rect 26835 24565 26847 24599
rect 26789 24559 26847 24565
rect 27430 24556 27436 24608
rect 27488 24596 27494 24608
rect 27816 24596 27844 24704
rect 28169 24701 28181 24704
rect 28215 24701 28227 24735
rect 28169 24695 28227 24701
rect 29089 24735 29147 24741
rect 29089 24701 29101 24735
rect 29135 24732 29147 24735
rect 29270 24732 29276 24744
rect 29135 24704 29276 24732
rect 29135 24701 29147 24704
rect 29089 24695 29147 24701
rect 29270 24692 29276 24704
rect 29328 24692 29334 24744
rect 29457 24735 29515 24741
rect 29457 24701 29469 24735
rect 29503 24732 29515 24735
rect 30006 24732 30012 24744
rect 29503 24704 30012 24732
rect 29503 24701 29515 24704
rect 29457 24695 29515 24701
rect 30006 24692 30012 24704
rect 30064 24692 30070 24744
rect 30834 24692 30840 24744
rect 30892 24732 30898 24744
rect 30929 24735 30987 24741
rect 30929 24732 30941 24735
rect 30892 24704 30941 24732
rect 30892 24692 30898 24704
rect 30929 24701 30941 24704
rect 30975 24701 30987 24735
rect 31110 24732 31116 24744
rect 31071 24704 31116 24732
rect 30929 24695 30987 24701
rect 31110 24692 31116 24704
rect 31168 24692 31174 24744
rect 31846 24692 31852 24744
rect 31904 24732 31910 24744
rect 31941 24735 31999 24741
rect 31941 24732 31953 24735
rect 31904 24704 31953 24732
rect 31904 24692 31910 24704
rect 31941 24701 31953 24704
rect 31987 24701 31999 24735
rect 31941 24695 31999 24701
rect 32401 24735 32459 24741
rect 32401 24701 32413 24735
rect 32447 24701 32459 24735
rect 32401 24695 32459 24701
rect 32769 24735 32827 24741
rect 32769 24701 32781 24735
rect 32815 24732 32827 24735
rect 33318 24732 33324 24744
rect 32815 24704 33324 24732
rect 32815 24701 32827 24704
rect 32769 24695 32827 24701
rect 28445 24667 28503 24673
rect 28445 24633 28457 24667
rect 28491 24664 28503 24667
rect 28534 24664 28540 24676
rect 28491 24636 28540 24664
rect 28491 24633 28503 24636
rect 28445 24627 28503 24633
rect 28534 24624 28540 24636
rect 28592 24624 28598 24676
rect 30098 24664 30104 24676
rect 28920 24636 29960 24664
rect 30059 24636 30104 24664
rect 28920 24605 28948 24636
rect 27488 24568 27844 24596
rect 28905 24599 28963 24605
rect 27488 24556 27494 24568
rect 28905 24565 28917 24599
rect 28951 24565 28963 24599
rect 29932 24596 29960 24636
rect 30098 24624 30104 24636
rect 30156 24624 30162 24676
rect 31570 24624 31576 24676
rect 31628 24664 31634 24676
rect 32416 24664 32444 24695
rect 33318 24692 33324 24704
rect 33376 24692 33382 24744
rect 34054 24732 34060 24744
rect 34015 24704 34060 24732
rect 34054 24692 34060 24704
rect 34112 24692 34118 24744
rect 35161 24735 35219 24741
rect 35161 24701 35173 24735
rect 35207 24701 35219 24735
rect 35161 24695 35219 24701
rect 31628 24636 32444 24664
rect 35176 24664 35204 24695
rect 35342 24692 35348 24744
rect 35400 24732 35406 24744
rect 35437 24735 35495 24741
rect 35437 24732 35449 24735
rect 35400 24704 35449 24732
rect 35400 24692 35406 24704
rect 35437 24701 35449 24704
rect 35483 24701 35495 24735
rect 35437 24695 35495 24701
rect 35618 24692 35624 24744
rect 35676 24732 35682 24744
rect 35802 24732 35808 24744
rect 35676 24704 35808 24732
rect 35676 24692 35682 24704
rect 35802 24692 35808 24704
rect 35860 24732 35866 24744
rect 36173 24735 36231 24741
rect 36173 24732 36185 24735
rect 35860 24704 36185 24732
rect 35860 24692 35866 24704
rect 36173 24701 36185 24704
rect 36219 24701 36231 24735
rect 36173 24695 36231 24701
rect 36265 24735 36323 24741
rect 36265 24701 36277 24735
rect 36311 24732 36323 24735
rect 36906 24732 36912 24744
rect 36311 24704 36912 24732
rect 36311 24701 36323 24704
rect 36265 24695 36323 24701
rect 36906 24692 36912 24704
rect 36964 24692 36970 24744
rect 37185 24735 37243 24741
rect 37185 24701 37197 24735
rect 37231 24732 37243 24735
rect 37274 24732 37280 24744
rect 37231 24704 37280 24732
rect 37231 24701 37243 24704
rect 37185 24695 37243 24701
rect 37274 24692 37280 24704
rect 37332 24692 37338 24744
rect 37458 24732 37464 24744
rect 37419 24704 37464 24732
rect 37458 24692 37464 24704
rect 37516 24692 37522 24744
rect 35250 24664 35256 24676
rect 35176 24636 35256 24664
rect 31628 24624 31634 24636
rect 35250 24624 35256 24636
rect 35308 24624 35314 24676
rect 32766 24596 32772 24608
rect 29932 24568 32772 24596
rect 28905 24559 28963 24565
rect 32766 24556 32772 24568
rect 32824 24596 32830 24608
rect 33042 24596 33048 24608
rect 32824 24568 33048 24596
rect 32824 24556 32830 24568
rect 33042 24556 33048 24568
rect 33100 24556 33106 24608
rect 34241 24599 34299 24605
rect 34241 24565 34253 24599
rect 34287 24596 34299 24599
rect 35434 24596 35440 24608
rect 34287 24568 35440 24596
rect 34287 24565 34299 24568
rect 34241 24559 34299 24565
rect 35434 24556 35440 24568
rect 35492 24556 35498 24608
rect 38562 24596 38568 24608
rect 38523 24568 38568 24596
rect 38562 24556 38568 24568
rect 38620 24556 38626 24608
rect 1104 24506 39836 24528
rect 1104 24454 19606 24506
rect 19658 24454 19670 24506
rect 19722 24454 19734 24506
rect 19786 24454 19798 24506
rect 19850 24454 39836 24506
rect 1104 24432 39836 24454
rect 1854 24392 1860 24404
rect 1815 24364 1860 24392
rect 1854 24352 1860 24364
rect 1912 24352 1918 24404
rect 7098 24352 7104 24404
rect 7156 24352 7162 24404
rect 8754 24352 8760 24404
rect 8812 24392 8818 24404
rect 8941 24395 8999 24401
rect 8941 24392 8953 24395
rect 8812 24364 8953 24392
rect 8812 24352 8818 24364
rect 8941 24361 8953 24364
rect 8987 24361 8999 24395
rect 8941 24355 8999 24361
rect 9769 24395 9827 24401
rect 9769 24361 9781 24395
rect 9815 24361 9827 24395
rect 9769 24355 9827 24361
rect 7116 24324 7144 24352
rect 7742 24324 7748 24336
rect 7116 24296 7748 24324
rect 7742 24284 7748 24296
rect 7800 24324 7806 24336
rect 9784 24324 9812 24355
rect 11146 24352 11152 24404
rect 11204 24392 11210 24404
rect 15378 24392 15384 24404
rect 11204 24364 14596 24392
rect 15339 24364 15384 24392
rect 11204 24352 11210 24364
rect 11164 24324 11192 24352
rect 7800 24296 8064 24324
rect 7800 24284 7806 24296
rect 1762 24256 1768 24268
rect 1723 24228 1768 24256
rect 1762 24216 1768 24228
rect 1820 24216 1826 24268
rect 2590 24256 2596 24268
rect 2551 24228 2596 24256
rect 2590 24216 2596 24228
rect 2648 24216 2654 24268
rect 3326 24256 3332 24268
rect 3287 24228 3332 24256
rect 3326 24216 3332 24228
rect 3384 24216 3390 24268
rect 3970 24216 3976 24268
rect 4028 24256 4034 24268
rect 4065 24259 4123 24265
rect 4065 24256 4077 24259
rect 4028 24228 4077 24256
rect 4028 24216 4034 24228
rect 4065 24225 4077 24228
rect 4111 24225 4123 24259
rect 7098 24256 7104 24268
rect 7059 24228 7104 24256
rect 4065 24219 4123 24225
rect 7098 24216 7104 24228
rect 7156 24216 7162 24268
rect 8036 24265 8064 24296
rect 8864 24296 9812 24324
rect 9968 24296 11192 24324
rect 8864 24265 8892 24296
rect 8021 24259 8079 24265
rect 8021 24225 8033 24259
rect 8067 24225 8079 24259
rect 8021 24219 8079 24225
rect 8849 24259 8907 24265
rect 8849 24225 8861 24259
rect 8895 24225 8907 24259
rect 9030 24256 9036 24268
rect 8991 24228 9036 24256
rect 8849 24219 8907 24225
rect 9030 24216 9036 24228
rect 9088 24216 9094 24268
rect 9968 24265 9996 24296
rect 11974 24284 11980 24336
rect 12032 24324 12038 24336
rect 12345 24327 12403 24333
rect 12345 24324 12357 24327
rect 12032 24296 12357 24324
rect 12032 24284 12038 24296
rect 12345 24293 12357 24296
rect 12391 24293 12403 24327
rect 12345 24287 12403 24293
rect 9953 24259 10011 24265
rect 9953 24225 9965 24259
rect 9999 24225 10011 24259
rect 9953 24219 10011 24225
rect 10229 24259 10287 24265
rect 10229 24225 10241 24259
rect 10275 24256 10287 24259
rect 11054 24256 11060 24268
rect 10275 24228 11060 24256
rect 10275 24225 10287 24228
rect 10229 24219 10287 24225
rect 11054 24216 11060 24228
rect 11112 24216 11118 24268
rect 11149 24259 11207 24265
rect 11149 24225 11161 24259
rect 11195 24225 11207 24259
rect 11149 24219 11207 24225
rect 2685 24191 2743 24197
rect 2685 24157 2697 24191
rect 2731 24188 2743 24191
rect 4798 24188 4804 24200
rect 2731 24160 4804 24188
rect 2731 24157 2743 24160
rect 2685 24151 2743 24157
rect 4798 24148 4804 24160
rect 4856 24148 4862 24200
rect 4982 24188 4988 24200
rect 4943 24160 4988 24188
rect 4982 24148 4988 24160
rect 5040 24148 5046 24200
rect 5261 24191 5319 24197
rect 5261 24157 5273 24191
rect 5307 24188 5319 24191
rect 7193 24191 7251 24197
rect 7193 24188 7205 24191
rect 5307 24160 7205 24188
rect 5307 24157 5319 24160
rect 5261 24151 5319 24157
rect 7193 24157 7205 24160
rect 7239 24157 7251 24191
rect 7193 24151 7251 24157
rect 11164 24120 11192 24219
rect 11238 24216 11244 24268
rect 11296 24256 11302 24268
rect 11333 24259 11391 24265
rect 11333 24256 11345 24259
rect 11296 24228 11345 24256
rect 11296 24216 11302 24228
rect 11333 24225 11345 24228
rect 11379 24225 11391 24259
rect 11882 24256 11888 24268
rect 11843 24228 11888 24256
rect 11333 24219 11391 24225
rect 11882 24216 11888 24228
rect 11940 24216 11946 24268
rect 12250 24256 12256 24268
rect 12211 24228 12256 24256
rect 12250 24216 12256 24228
rect 12308 24216 12314 24268
rect 13446 24256 13452 24268
rect 13407 24228 13452 24256
rect 13446 24216 13452 24228
rect 13504 24216 13510 24268
rect 13906 24256 13912 24268
rect 13867 24228 13912 24256
rect 13906 24216 13912 24228
rect 13964 24216 13970 24268
rect 14568 24265 14596 24364
rect 15378 24352 15384 24364
rect 15436 24352 15442 24404
rect 20346 24392 20352 24404
rect 16592 24364 20352 24392
rect 15838 24284 15844 24336
rect 15896 24324 15902 24336
rect 15933 24327 15991 24333
rect 15933 24324 15945 24327
rect 15896 24296 15945 24324
rect 15896 24284 15902 24296
rect 15933 24293 15945 24296
rect 15979 24293 15991 24327
rect 15933 24287 15991 24293
rect 16592 24265 16620 24364
rect 20346 24352 20352 24364
rect 20404 24352 20410 24404
rect 20898 24352 20904 24404
rect 20956 24392 20962 24404
rect 21085 24395 21143 24401
rect 21085 24392 21097 24395
rect 20956 24364 21097 24392
rect 20956 24352 20962 24364
rect 21085 24361 21097 24364
rect 21131 24361 21143 24395
rect 21085 24355 21143 24361
rect 22094 24352 22100 24404
rect 22152 24392 22158 24404
rect 22152 24364 22416 24392
rect 22152 24352 22158 24364
rect 18966 24324 18972 24336
rect 16960 24296 18972 24324
rect 16960 24265 16988 24296
rect 18966 24284 18972 24296
rect 19024 24284 19030 24336
rect 19150 24284 19156 24336
rect 19208 24324 19214 24336
rect 22186 24324 22192 24336
rect 19208 24296 22192 24324
rect 19208 24284 19214 24296
rect 22186 24284 22192 24296
rect 22244 24284 22250 24336
rect 22388 24324 22416 24364
rect 23842 24352 23848 24404
rect 23900 24352 23906 24404
rect 24302 24392 24308 24404
rect 24263 24364 24308 24392
rect 24302 24352 24308 24364
rect 24360 24352 24366 24404
rect 27614 24352 27620 24404
rect 27672 24392 27678 24404
rect 27801 24395 27859 24401
rect 27801 24392 27813 24395
rect 27672 24364 27813 24392
rect 27672 24352 27678 24364
rect 27801 24361 27813 24364
rect 27847 24361 27859 24395
rect 27801 24355 27859 24361
rect 31018 24352 31024 24404
rect 31076 24392 31082 24404
rect 31076 24364 38240 24392
rect 31076 24352 31082 24364
rect 23860 24324 23888 24352
rect 25590 24324 25596 24336
rect 22388 24296 23888 24324
rect 25424 24296 25596 24324
rect 14553 24259 14611 24265
rect 14553 24225 14565 24259
rect 14599 24225 14611 24259
rect 14553 24219 14611 24225
rect 15289 24259 15347 24265
rect 15289 24225 15301 24259
rect 15335 24225 15347 24259
rect 15289 24219 15347 24225
rect 16209 24259 16267 24265
rect 16209 24225 16221 24259
rect 16255 24225 16267 24259
rect 16209 24219 16267 24225
rect 16577 24259 16635 24265
rect 16577 24225 16589 24259
rect 16623 24225 16635 24259
rect 16577 24219 16635 24225
rect 16945 24259 17003 24265
rect 16945 24225 16957 24259
rect 16991 24225 17003 24259
rect 16945 24219 17003 24225
rect 17129 24259 17187 24265
rect 17129 24225 17141 24259
rect 17175 24225 17187 24259
rect 17770 24256 17776 24268
rect 17731 24228 17776 24256
rect 17129 24219 17187 24225
rect 13725 24191 13783 24197
rect 13725 24157 13737 24191
rect 13771 24188 13783 24191
rect 15304 24188 15332 24219
rect 13771 24160 15332 24188
rect 16224 24188 16252 24219
rect 16666 24188 16672 24200
rect 16224 24160 16672 24188
rect 13771 24157 13783 24160
rect 13725 24151 13783 24157
rect 16666 24148 16672 24160
rect 16724 24148 16730 24200
rect 14645 24123 14703 24129
rect 14645 24120 14657 24123
rect 11164 24092 14657 24120
rect 14645 24089 14657 24092
rect 14691 24120 14703 24123
rect 17144 24120 17172 24219
rect 17770 24216 17776 24228
rect 17828 24216 17834 24268
rect 18322 24256 18328 24268
rect 18283 24228 18328 24256
rect 18322 24216 18328 24228
rect 18380 24216 18386 24268
rect 18601 24259 18659 24265
rect 18601 24225 18613 24259
rect 18647 24225 18659 24259
rect 18601 24219 18659 24225
rect 18616 24188 18644 24219
rect 18782 24216 18788 24268
rect 18840 24256 18846 24268
rect 18877 24259 18935 24265
rect 18877 24256 18889 24259
rect 18840 24228 18889 24256
rect 18840 24216 18846 24228
rect 18877 24225 18889 24228
rect 18923 24225 18935 24259
rect 19058 24256 19064 24268
rect 19019 24228 19064 24256
rect 18877 24219 18935 24225
rect 19058 24216 19064 24228
rect 19116 24216 19122 24268
rect 19337 24259 19395 24265
rect 19337 24225 19349 24259
rect 19383 24256 19395 24259
rect 19518 24256 19524 24268
rect 19383 24228 19524 24256
rect 19383 24225 19395 24228
rect 19337 24219 19395 24225
rect 19518 24216 19524 24228
rect 19576 24216 19582 24268
rect 19797 24259 19855 24265
rect 19797 24225 19809 24259
rect 19843 24256 19855 24259
rect 20254 24256 20260 24268
rect 19843 24228 20260 24256
rect 19843 24225 19855 24228
rect 19797 24219 19855 24225
rect 20254 24216 20260 24228
rect 20312 24216 20318 24268
rect 20898 24256 20904 24268
rect 20859 24228 20904 24256
rect 20898 24216 20904 24228
rect 20956 24216 20962 24268
rect 21726 24256 21732 24268
rect 21687 24228 21732 24256
rect 21726 24216 21732 24228
rect 21784 24216 21790 24268
rect 22388 24265 22416 24296
rect 22373 24259 22431 24265
rect 22373 24225 22385 24259
rect 22419 24225 22431 24259
rect 22373 24219 22431 24225
rect 22646 24216 22652 24268
rect 22704 24256 22710 24268
rect 23676 24265 23704 24296
rect 22741 24259 22799 24265
rect 22741 24256 22753 24259
rect 22704 24228 22753 24256
rect 22704 24216 22710 24228
rect 22741 24225 22753 24228
rect 22787 24225 22799 24259
rect 22741 24219 22799 24225
rect 23661 24259 23719 24265
rect 23661 24225 23673 24259
rect 23707 24225 23719 24259
rect 23842 24256 23848 24268
rect 23803 24228 23848 24256
rect 23661 24219 23719 24225
rect 18690 24188 18696 24200
rect 18603 24160 18696 24188
rect 18690 24148 18696 24160
rect 18748 24188 18754 24200
rect 20162 24188 20168 24200
rect 18748 24160 20168 24188
rect 18748 24148 18754 24160
rect 20162 24148 20168 24160
rect 20220 24148 20226 24200
rect 22756 24188 22784 24219
rect 23842 24216 23848 24228
rect 23900 24216 23906 24268
rect 25424 24265 25452 24296
rect 25590 24284 25596 24296
rect 25648 24324 25654 24336
rect 25958 24324 25964 24336
rect 25648 24296 25964 24324
rect 25648 24284 25654 24296
rect 25958 24284 25964 24296
rect 26016 24284 26022 24336
rect 27816 24296 29960 24324
rect 24213 24259 24271 24265
rect 24213 24225 24225 24259
rect 24259 24225 24271 24259
rect 24213 24219 24271 24225
rect 25409 24259 25467 24265
rect 25409 24225 25421 24259
rect 25455 24225 25467 24259
rect 25409 24219 25467 24225
rect 25777 24259 25835 24265
rect 25777 24225 25789 24259
rect 25823 24256 25835 24259
rect 26510 24256 26516 24268
rect 25823 24228 26516 24256
rect 25823 24225 25835 24228
rect 25777 24219 25835 24225
rect 24228 24188 24256 24219
rect 26510 24216 26516 24228
rect 26568 24216 26574 24268
rect 27816 24265 27844 24296
rect 27065 24259 27123 24265
rect 27065 24225 27077 24259
rect 27111 24256 27123 24259
rect 27801 24259 27859 24265
rect 27111 24228 27292 24256
rect 27111 24225 27123 24228
rect 27065 24219 27123 24225
rect 22756 24160 24256 24188
rect 25869 24191 25927 24197
rect 25869 24157 25881 24191
rect 25915 24188 25927 24191
rect 27154 24188 27160 24200
rect 25915 24160 27160 24188
rect 25915 24157 25927 24160
rect 25869 24151 25927 24157
rect 27154 24148 27160 24160
rect 27212 24148 27218 24200
rect 27264 24188 27292 24228
rect 27801 24225 27813 24259
rect 27847 24225 27859 24259
rect 28350 24256 28356 24268
rect 28311 24228 28356 24256
rect 27801 24219 27859 24225
rect 28350 24216 28356 24228
rect 28408 24216 28414 24268
rect 28534 24256 28540 24268
rect 28495 24228 28540 24256
rect 28534 24216 28540 24228
rect 28592 24216 28598 24268
rect 27890 24188 27896 24200
rect 27264 24160 27896 24188
rect 27890 24148 27896 24160
rect 27948 24148 27954 24200
rect 29454 24148 29460 24200
rect 29512 24188 29518 24200
rect 29825 24191 29883 24197
rect 29825 24188 29837 24191
rect 29512 24160 29837 24188
rect 29512 24148 29518 24160
rect 29825 24157 29837 24160
rect 29871 24157 29883 24191
rect 29932 24188 29960 24296
rect 36262 24284 36268 24336
rect 36320 24324 36326 24336
rect 36446 24324 36452 24336
rect 36320 24296 36452 24324
rect 36320 24284 36326 24296
rect 36446 24284 36452 24296
rect 36504 24324 36510 24336
rect 36504 24296 36676 24324
rect 36504 24284 36510 24296
rect 30098 24256 30104 24268
rect 30059 24228 30104 24256
rect 30098 24216 30104 24228
rect 30156 24216 30162 24268
rect 31846 24216 31852 24268
rect 31904 24256 31910 24268
rect 32122 24256 32128 24268
rect 31904 24228 32128 24256
rect 31904 24216 31910 24228
rect 32122 24216 32128 24228
rect 32180 24256 32186 24268
rect 32309 24259 32367 24265
rect 32309 24256 32321 24259
rect 32180 24228 32321 24256
rect 32180 24216 32186 24228
rect 32309 24225 32321 24228
rect 32355 24225 32367 24259
rect 32309 24219 32367 24225
rect 32582 24216 32588 24268
rect 32640 24256 32646 24268
rect 33137 24259 33195 24265
rect 33137 24256 33149 24259
rect 32640 24228 33149 24256
rect 32640 24216 32646 24228
rect 33137 24225 33149 24228
rect 33183 24225 33195 24259
rect 33318 24256 33324 24268
rect 33231 24228 33324 24256
rect 33137 24219 33195 24225
rect 33318 24216 33324 24228
rect 33376 24256 33382 24268
rect 36354 24256 36360 24268
rect 33376 24228 35388 24256
rect 36315 24228 36360 24256
rect 33376 24216 33382 24228
rect 30282 24188 30288 24200
rect 29932 24160 30288 24188
rect 29825 24151 29883 24157
rect 30282 24148 30288 24160
rect 30340 24148 30346 24200
rect 32490 24148 32496 24200
rect 32548 24188 32554 24200
rect 33336 24188 33364 24216
rect 33962 24188 33968 24200
rect 32548 24160 33364 24188
rect 33923 24160 33968 24188
rect 32548 24148 32554 24160
rect 33962 24148 33968 24160
rect 34020 24148 34026 24200
rect 34238 24188 34244 24200
rect 34199 24160 34244 24188
rect 34238 24148 34244 24160
rect 34296 24148 34302 24200
rect 35360 24197 35388 24228
rect 36354 24216 36360 24228
rect 36412 24216 36418 24268
rect 36648 24265 36676 24296
rect 36633 24259 36691 24265
rect 36633 24225 36645 24259
rect 36679 24225 36691 24259
rect 36633 24219 36691 24225
rect 38013 24259 38071 24265
rect 38013 24225 38025 24259
rect 38059 24225 38071 24259
rect 38212 24256 38240 24364
rect 38286 24256 38292 24268
rect 38199 24228 38292 24256
rect 38013 24219 38071 24225
rect 35345 24191 35403 24197
rect 35345 24157 35357 24191
rect 35391 24157 35403 24191
rect 36446 24188 36452 24200
rect 36407 24160 36452 24188
rect 35345 24151 35403 24157
rect 36446 24148 36452 24160
rect 36504 24148 36510 24200
rect 38028 24188 38056 24219
rect 38286 24216 38292 24228
rect 38344 24216 38350 24268
rect 38930 24256 38936 24268
rect 38891 24228 38936 24256
rect 38930 24216 38936 24228
rect 38988 24216 38994 24268
rect 38102 24188 38108 24200
rect 38015 24160 38108 24188
rect 38102 24148 38108 24160
rect 38160 24188 38166 24200
rect 39025 24191 39083 24197
rect 39025 24188 39037 24191
rect 38160 24160 39037 24188
rect 38160 24148 38166 24160
rect 39025 24157 39037 24160
rect 39071 24157 39083 24191
rect 39025 24151 39083 24157
rect 14691 24092 17172 24120
rect 14691 24089 14703 24092
rect 14645 24083 14703 24089
rect 18322 24080 18328 24132
rect 18380 24120 18386 24132
rect 22278 24120 22284 24132
rect 18380 24092 22284 24120
rect 18380 24080 18386 24092
rect 22278 24080 22284 24092
rect 22336 24080 22342 24132
rect 25225 24123 25283 24129
rect 25225 24089 25237 24123
rect 25271 24120 25283 24123
rect 27522 24120 27528 24132
rect 25271 24092 27528 24120
rect 25271 24089 25283 24092
rect 25225 24083 25283 24089
rect 27522 24080 27528 24092
rect 27580 24080 27586 24132
rect 33134 24120 33140 24132
rect 33095 24092 33140 24120
rect 33134 24080 33140 24092
rect 33192 24080 33198 24132
rect 37458 24080 37464 24132
rect 37516 24120 37522 24132
rect 37829 24123 37887 24129
rect 37829 24120 37841 24123
rect 37516 24092 37841 24120
rect 37516 24080 37522 24092
rect 37829 24089 37841 24092
rect 37875 24089 37887 24123
rect 37829 24083 37887 24089
rect 3418 24052 3424 24064
rect 3379 24024 3424 24052
rect 3418 24012 3424 24024
rect 3476 24012 3482 24064
rect 4157 24055 4215 24061
rect 4157 24021 4169 24055
rect 4203 24052 4215 24055
rect 4614 24052 4620 24064
rect 4203 24024 4620 24052
rect 4203 24021 4215 24024
rect 4157 24015 4215 24021
rect 4614 24012 4620 24024
rect 4672 24012 4678 24064
rect 5626 24012 5632 24064
rect 5684 24052 5690 24064
rect 6549 24055 6607 24061
rect 6549 24052 6561 24055
rect 5684 24024 6561 24052
rect 5684 24012 5690 24024
rect 6549 24021 6561 24024
rect 6595 24052 6607 24055
rect 6822 24052 6828 24064
rect 6595 24024 6828 24052
rect 6595 24021 6607 24024
rect 6549 24015 6607 24021
rect 6822 24012 6828 24024
rect 6880 24012 6886 24064
rect 9950 24012 9956 24064
rect 10008 24052 10014 24064
rect 13998 24052 14004 24064
rect 10008 24024 14004 24052
rect 10008 24012 10014 24024
rect 13998 24012 14004 24024
rect 14056 24012 14062 24064
rect 21821 24055 21879 24061
rect 21821 24021 21833 24055
rect 21867 24052 21879 24055
rect 22462 24052 22468 24064
rect 21867 24024 22468 24052
rect 21867 24021 21879 24024
rect 21821 24015 21879 24021
rect 22462 24012 22468 24024
rect 22520 24052 22526 24064
rect 23106 24052 23112 24064
rect 22520 24024 23112 24052
rect 22520 24012 22526 24024
rect 23106 24012 23112 24024
rect 23164 24012 23170 24064
rect 31389 24055 31447 24061
rect 31389 24021 31401 24055
rect 31435 24052 31447 24055
rect 31478 24052 31484 24064
rect 31435 24024 31484 24052
rect 31435 24021 31447 24024
rect 31389 24015 31447 24021
rect 31478 24012 31484 24024
rect 31536 24012 31542 24064
rect 1104 23962 39836 23984
rect 1104 23910 4246 23962
rect 4298 23910 4310 23962
rect 4362 23910 4374 23962
rect 4426 23910 4438 23962
rect 4490 23910 34966 23962
rect 35018 23910 35030 23962
rect 35082 23910 35094 23962
rect 35146 23910 35158 23962
rect 35210 23910 39836 23962
rect 1104 23888 39836 23910
rect 7742 23848 7748 23860
rect 7703 23820 7748 23848
rect 7742 23808 7748 23820
rect 7800 23848 7806 23860
rect 8018 23848 8024 23860
rect 7800 23820 8024 23848
rect 7800 23808 7806 23820
rect 8018 23808 8024 23820
rect 8076 23808 8082 23860
rect 15470 23808 15476 23860
rect 15528 23848 15534 23860
rect 17405 23851 17463 23857
rect 15528 23820 17356 23848
rect 15528 23808 15534 23820
rect 2590 23780 2596 23792
rect 2551 23752 2596 23780
rect 2590 23740 2596 23752
rect 2648 23740 2654 23792
rect 3694 23780 3700 23792
rect 2884 23752 3700 23780
rect 2685 23647 2743 23653
rect 2685 23613 2697 23647
rect 2731 23644 2743 23647
rect 2884 23644 2912 23752
rect 3694 23740 3700 23752
rect 3752 23780 3758 23792
rect 4249 23783 4307 23789
rect 4249 23780 4261 23783
rect 3752 23752 4261 23780
rect 3752 23740 3758 23752
rect 4249 23749 4261 23752
rect 4295 23749 4307 23783
rect 4249 23743 4307 23749
rect 5537 23783 5595 23789
rect 5537 23749 5549 23783
rect 5583 23780 5595 23783
rect 7098 23780 7104 23792
rect 5583 23752 7104 23780
rect 5583 23749 5595 23752
rect 5537 23743 5595 23749
rect 7098 23740 7104 23752
rect 7156 23740 7162 23792
rect 11882 23740 11888 23792
rect 11940 23780 11946 23792
rect 12529 23783 12587 23789
rect 12529 23780 12541 23783
rect 11940 23752 12541 23780
rect 11940 23740 11946 23752
rect 12529 23749 12541 23752
rect 12575 23749 12587 23783
rect 12529 23743 12587 23749
rect 15286 23740 15292 23792
rect 15344 23780 15350 23792
rect 15565 23783 15623 23789
rect 15565 23780 15577 23783
rect 15344 23752 15577 23780
rect 15344 23740 15350 23752
rect 15565 23749 15577 23752
rect 15611 23780 15623 23783
rect 15611 23752 16988 23780
rect 15611 23749 15623 23752
rect 15565 23743 15623 23749
rect 2958 23672 2964 23724
rect 3016 23712 3022 23724
rect 3329 23715 3387 23721
rect 3329 23712 3341 23715
rect 3016 23684 3341 23712
rect 3016 23672 3022 23684
rect 3329 23681 3341 23684
rect 3375 23681 3387 23715
rect 9674 23712 9680 23724
rect 9635 23684 9680 23712
rect 3329 23675 3387 23681
rect 9674 23672 9680 23684
rect 9732 23672 9738 23724
rect 3234 23644 3240 23656
rect 2731 23616 2912 23644
rect 3195 23616 3240 23644
rect 2731 23613 2743 23616
rect 2685 23607 2743 23613
rect 3234 23604 3240 23616
rect 3292 23604 3298 23656
rect 3970 23604 3976 23656
rect 4028 23644 4034 23656
rect 4065 23647 4123 23653
rect 4065 23644 4077 23647
rect 4028 23616 4077 23644
rect 4028 23604 4034 23616
rect 4065 23613 4077 23616
rect 4111 23613 4123 23647
rect 5718 23644 5724 23656
rect 5679 23616 5724 23644
rect 4065 23607 4123 23613
rect 5718 23604 5724 23616
rect 5776 23604 5782 23656
rect 6089 23647 6147 23653
rect 6089 23613 6101 23647
rect 6135 23613 6147 23647
rect 6089 23607 6147 23613
rect 6104 23576 6132 23607
rect 6178 23604 6184 23656
rect 6236 23644 6242 23656
rect 7561 23647 7619 23653
rect 6236 23616 6281 23644
rect 6236 23604 6242 23616
rect 7561 23613 7573 23647
rect 7607 23644 7619 23647
rect 7834 23644 7840 23656
rect 7607 23616 7840 23644
rect 7607 23613 7619 23616
rect 7561 23607 7619 23613
rect 7834 23604 7840 23616
rect 7892 23604 7898 23656
rect 8941 23647 8999 23653
rect 8941 23613 8953 23647
rect 8987 23613 8999 23647
rect 8941 23607 8999 23613
rect 6822 23576 6828 23588
rect 6104 23548 6828 23576
rect 6822 23536 6828 23548
rect 6880 23536 6886 23588
rect 8956 23576 8984 23607
rect 9030 23604 9036 23656
rect 9088 23644 9094 23656
rect 9125 23647 9183 23653
rect 9125 23644 9137 23647
rect 9088 23616 9137 23644
rect 9088 23604 9094 23616
rect 9125 23613 9137 23616
rect 9171 23613 9183 23647
rect 9125 23607 9183 23613
rect 9585 23647 9643 23653
rect 9585 23613 9597 23647
rect 9631 23644 9643 23647
rect 9766 23644 9772 23656
rect 9631 23616 9772 23644
rect 9631 23613 9643 23616
rect 9585 23607 9643 23613
rect 9766 23604 9772 23616
rect 9824 23604 9830 23656
rect 11057 23647 11115 23653
rect 11057 23613 11069 23647
rect 11103 23644 11115 23647
rect 11146 23644 11152 23656
rect 11103 23616 11152 23644
rect 11103 23613 11115 23616
rect 11057 23607 11115 23613
rect 11146 23604 11152 23616
rect 11204 23604 11210 23656
rect 11609 23647 11667 23653
rect 11609 23613 11621 23647
rect 11655 23613 11667 23647
rect 11609 23607 11667 23613
rect 11793 23647 11851 23653
rect 11793 23613 11805 23647
rect 11839 23644 11851 23647
rect 11900 23644 11928 23740
rect 13998 23712 14004 23724
rect 12452 23684 13216 23712
rect 13959 23684 14004 23712
rect 11839 23616 11928 23644
rect 11839 23613 11851 23616
rect 11793 23607 11851 23613
rect 10502 23576 10508 23588
rect 8956 23548 10508 23576
rect 10502 23536 10508 23548
rect 10560 23536 10566 23588
rect 11624 23576 11652 23607
rect 12066 23604 12072 23656
rect 12124 23644 12130 23656
rect 12452 23644 12480 23684
rect 12618 23644 12624 23656
rect 12124 23616 12480 23644
rect 12579 23616 12624 23644
rect 12124 23604 12130 23616
rect 12618 23604 12624 23616
rect 12676 23604 12682 23656
rect 13188 23653 13216 23684
rect 13998 23672 14004 23684
rect 14056 23672 14062 23724
rect 14277 23715 14335 23721
rect 14277 23681 14289 23715
rect 14323 23712 14335 23715
rect 16853 23715 16911 23721
rect 16853 23712 16865 23715
rect 14323 23684 16865 23712
rect 14323 23681 14335 23684
rect 14277 23675 14335 23681
rect 16853 23681 16865 23684
rect 16899 23681 16911 23715
rect 16853 23675 16911 23681
rect 13173 23647 13231 23653
rect 13173 23613 13185 23647
rect 13219 23644 13231 23647
rect 13722 23644 13728 23656
rect 13219 23616 13728 23644
rect 13219 23613 13231 23616
rect 13173 23607 13231 23613
rect 13722 23604 13728 23616
rect 13780 23604 13786 23656
rect 14550 23604 14556 23656
rect 14608 23644 14614 23656
rect 16117 23647 16175 23653
rect 16117 23644 16129 23647
rect 14608 23616 16129 23644
rect 14608 23604 14614 23616
rect 16117 23613 16129 23616
rect 16163 23613 16175 23647
rect 16117 23607 16175 23613
rect 16393 23647 16451 23653
rect 16393 23613 16405 23647
rect 16439 23613 16451 23647
rect 16393 23607 16451 23613
rect 12250 23576 12256 23588
rect 11624 23548 12256 23576
rect 12250 23536 12256 23548
rect 12308 23576 12314 23588
rect 12308 23548 13032 23576
rect 12308 23536 12314 23548
rect 13004 23520 13032 23548
rect 15194 23536 15200 23588
rect 15252 23576 15258 23588
rect 16301 23579 16359 23585
rect 16301 23576 16313 23579
rect 15252 23548 16313 23576
rect 15252 23536 15258 23548
rect 16301 23545 16313 23548
rect 16347 23545 16359 23579
rect 16301 23539 16359 23545
rect 1486 23468 1492 23520
rect 1544 23508 1550 23520
rect 4982 23508 4988 23520
rect 1544 23480 4988 23508
rect 1544 23468 1550 23480
rect 4982 23468 4988 23480
rect 5040 23468 5046 23520
rect 11054 23508 11060 23520
rect 11015 23480 11060 23508
rect 11054 23468 11060 23480
rect 11112 23468 11118 23520
rect 12986 23468 12992 23520
rect 13044 23508 13050 23520
rect 16408 23508 16436 23607
rect 16960 23576 16988 23752
rect 17328 23653 17356 23820
rect 17405 23817 17417 23851
rect 17451 23848 17463 23851
rect 17586 23848 17592 23860
rect 17451 23820 17592 23848
rect 17451 23817 17463 23820
rect 17405 23811 17463 23817
rect 17586 23808 17592 23820
rect 17644 23808 17650 23860
rect 18874 23808 18880 23860
rect 18932 23848 18938 23860
rect 19518 23848 19524 23860
rect 18932 23820 19524 23848
rect 18932 23808 18938 23820
rect 18322 23712 18328 23724
rect 18283 23684 18328 23712
rect 18322 23672 18328 23684
rect 18380 23672 18386 23724
rect 19168 23656 19196 23820
rect 19518 23808 19524 23820
rect 19576 23808 19582 23860
rect 19705 23851 19763 23857
rect 19705 23817 19717 23851
rect 19751 23848 19763 23851
rect 21174 23848 21180 23860
rect 19751 23820 21180 23848
rect 19751 23817 19763 23820
rect 19705 23811 19763 23817
rect 21174 23808 21180 23820
rect 21232 23808 21238 23860
rect 28629 23851 28687 23857
rect 28629 23817 28641 23851
rect 28675 23848 28687 23851
rect 29546 23848 29552 23860
rect 28675 23820 29552 23848
rect 28675 23817 28687 23820
rect 28629 23811 28687 23817
rect 29546 23808 29552 23820
rect 29604 23808 29610 23860
rect 32401 23851 32459 23857
rect 32401 23817 32413 23851
rect 32447 23848 32459 23851
rect 32674 23848 32680 23860
rect 32447 23820 32680 23848
rect 32447 23817 32459 23820
rect 32401 23811 32459 23817
rect 32674 23808 32680 23820
rect 32732 23808 32738 23860
rect 34514 23808 34520 23860
rect 34572 23848 34578 23860
rect 34698 23848 34704 23860
rect 34572 23820 34704 23848
rect 34572 23808 34578 23820
rect 34698 23808 34704 23820
rect 34756 23808 34762 23860
rect 38930 23808 38936 23860
rect 38988 23848 38994 23860
rect 39025 23851 39083 23857
rect 39025 23848 39037 23851
rect 38988 23820 39037 23848
rect 38988 23808 38994 23820
rect 39025 23817 39037 23820
rect 39071 23817 39083 23851
rect 39025 23811 39083 23817
rect 20162 23740 20168 23792
rect 20220 23780 20226 23792
rect 20349 23783 20407 23789
rect 20349 23780 20361 23783
rect 20220 23752 20361 23780
rect 20220 23740 20226 23752
rect 20349 23749 20361 23752
rect 20395 23749 20407 23783
rect 22833 23783 22891 23789
rect 22833 23780 22845 23783
rect 20349 23743 20407 23749
rect 21928 23752 22845 23780
rect 17313 23647 17371 23653
rect 17313 23613 17325 23647
rect 17359 23613 17371 23647
rect 18690 23644 18696 23656
rect 18651 23616 18696 23644
rect 17313 23607 17371 23613
rect 18690 23604 18696 23616
rect 18748 23604 18754 23656
rect 18782 23604 18788 23656
rect 18840 23644 18846 23656
rect 18877 23647 18935 23653
rect 18877 23644 18889 23647
rect 18840 23616 18889 23644
rect 18840 23604 18846 23616
rect 18877 23613 18889 23616
rect 18923 23613 18935 23647
rect 18877 23607 18935 23613
rect 19061 23647 19119 23653
rect 19061 23613 19073 23647
rect 19107 23613 19119 23647
rect 19061 23607 19119 23613
rect 19076 23576 19104 23607
rect 19150 23604 19156 23656
rect 19208 23644 19214 23656
rect 19337 23647 19395 23653
rect 19337 23644 19349 23647
rect 19208 23616 19349 23644
rect 19208 23604 19214 23616
rect 19337 23613 19349 23616
rect 19383 23613 19395 23647
rect 20530 23644 20536 23656
rect 20491 23616 20536 23644
rect 19337 23607 19395 23613
rect 20530 23604 20536 23616
rect 20588 23604 20594 23656
rect 20806 23644 20812 23656
rect 20767 23616 20812 23644
rect 20806 23604 20812 23616
rect 20864 23604 20870 23656
rect 20898 23604 20904 23656
rect 20956 23644 20962 23656
rect 21453 23647 21511 23653
rect 21453 23644 21465 23647
rect 20956 23616 21465 23644
rect 20956 23604 20962 23616
rect 21453 23613 21465 23616
rect 21499 23613 21511 23647
rect 21453 23607 21511 23613
rect 16960 23548 19104 23576
rect 21468 23576 21496 23607
rect 21726 23604 21732 23656
rect 21784 23644 21790 23656
rect 21928 23653 21956 23752
rect 22833 23749 22845 23752
rect 22879 23749 22891 23783
rect 27890 23780 27896 23792
rect 22833 23743 22891 23749
rect 25884 23752 27896 23780
rect 22094 23672 22100 23724
rect 22152 23712 22158 23724
rect 22189 23715 22247 23721
rect 22189 23712 22201 23715
rect 22152 23684 22201 23712
rect 22152 23672 22158 23684
rect 22189 23681 22201 23684
rect 22235 23712 22247 23715
rect 22738 23712 22744 23724
rect 22235 23684 22744 23712
rect 22235 23681 22247 23684
rect 22189 23675 22247 23681
rect 22738 23672 22744 23684
rect 22796 23672 22802 23724
rect 21913 23647 21971 23653
rect 21913 23644 21925 23647
rect 21784 23616 21925 23644
rect 21784 23604 21790 23616
rect 21913 23613 21925 23616
rect 21959 23613 21971 23647
rect 22646 23644 22652 23656
rect 22607 23616 22652 23644
rect 21913 23607 21971 23613
rect 22646 23604 22652 23616
rect 22704 23604 22710 23656
rect 22848 23644 22876 23743
rect 23658 23672 23664 23724
rect 23716 23712 23722 23724
rect 25884 23721 25912 23752
rect 27890 23740 27896 23752
rect 27948 23740 27954 23792
rect 32490 23780 32496 23792
rect 29564 23752 32496 23780
rect 23753 23715 23811 23721
rect 23753 23712 23765 23715
rect 23716 23684 23765 23712
rect 23716 23672 23722 23684
rect 23753 23681 23765 23684
rect 23799 23681 23811 23715
rect 23753 23675 23811 23681
rect 25869 23715 25927 23721
rect 25869 23681 25881 23715
rect 25915 23681 25927 23715
rect 27338 23712 27344 23724
rect 25869 23675 25927 23681
rect 26252 23684 27344 23712
rect 26252 23656 26280 23684
rect 27338 23672 27344 23684
rect 27396 23712 27402 23724
rect 27396 23684 28028 23712
rect 27396 23672 27402 23684
rect 23842 23644 23848 23656
rect 22848 23616 23848 23644
rect 23842 23604 23848 23616
rect 23900 23604 23906 23656
rect 24029 23647 24087 23653
rect 24029 23613 24041 23647
rect 24075 23613 24087 23647
rect 24394 23644 24400 23656
rect 24355 23616 24400 23644
rect 24029 23607 24087 23613
rect 22278 23576 22284 23588
rect 21468 23548 22284 23576
rect 22278 23536 22284 23548
rect 22336 23576 22342 23588
rect 24044 23576 24072 23607
rect 24394 23604 24400 23616
rect 24452 23604 24458 23656
rect 25133 23647 25191 23653
rect 25133 23613 25145 23647
rect 25179 23644 25191 23647
rect 25774 23644 25780 23656
rect 25179 23616 25780 23644
rect 25179 23613 25191 23616
rect 25133 23607 25191 23613
rect 25774 23604 25780 23616
rect 25832 23604 25838 23656
rect 26234 23644 26240 23656
rect 26195 23616 26240 23644
rect 26234 23604 26240 23616
rect 26292 23604 26298 23656
rect 26605 23647 26663 23653
rect 26605 23613 26617 23647
rect 26651 23644 26663 23647
rect 26694 23644 26700 23656
rect 26651 23616 26700 23644
rect 26651 23613 26663 23616
rect 26605 23607 26663 23613
rect 26694 23604 26700 23616
rect 26752 23604 26758 23656
rect 26878 23604 26884 23656
rect 26936 23644 26942 23656
rect 27249 23647 27307 23653
rect 27249 23644 27261 23647
rect 26936 23616 27261 23644
rect 26936 23604 26942 23616
rect 27249 23613 27261 23616
rect 27295 23613 27307 23647
rect 27890 23644 27896 23656
rect 27851 23616 27896 23644
rect 27249 23607 27307 23613
rect 27890 23604 27896 23616
rect 27948 23604 27954 23656
rect 28000 23653 28028 23684
rect 27985 23647 28043 23653
rect 27985 23613 27997 23647
rect 28031 23613 28043 23647
rect 27985 23607 28043 23613
rect 28442 23604 28448 23656
rect 28500 23644 28506 23656
rect 29564 23653 29592 23752
rect 30837 23715 30895 23721
rect 30837 23681 30849 23715
rect 30883 23712 30895 23715
rect 31110 23712 31116 23724
rect 30883 23684 31116 23712
rect 30883 23681 30895 23684
rect 30837 23675 30895 23681
rect 31110 23672 31116 23684
rect 31168 23672 31174 23724
rect 31404 23721 31432 23752
rect 32490 23740 32496 23752
rect 32548 23740 32554 23792
rect 32582 23740 32588 23792
rect 32640 23780 32646 23792
rect 32640 23752 33364 23780
rect 32640 23740 32646 23752
rect 31389 23715 31447 23721
rect 31389 23681 31401 23715
rect 31435 23681 31447 23715
rect 31389 23675 31447 23681
rect 31570 23672 31576 23724
rect 31628 23712 31634 23724
rect 31849 23715 31907 23721
rect 31849 23712 31861 23715
rect 31628 23684 31861 23712
rect 31628 23672 31634 23684
rect 31849 23681 31861 23684
rect 31895 23681 31907 23715
rect 31849 23675 31907 23681
rect 33045 23715 33103 23721
rect 33045 23681 33057 23715
rect 33091 23712 33103 23715
rect 33134 23712 33140 23724
rect 33091 23684 33140 23712
rect 33091 23681 33103 23684
rect 33045 23675 33103 23681
rect 33134 23672 33140 23684
rect 33192 23672 33198 23724
rect 28537 23647 28595 23653
rect 28537 23644 28549 23647
rect 28500 23616 28549 23644
rect 28500 23604 28506 23616
rect 28537 23613 28549 23616
rect 28583 23613 28595 23647
rect 28537 23607 28595 23613
rect 29549 23647 29607 23653
rect 29549 23613 29561 23647
rect 29595 23613 29607 23647
rect 29549 23607 29607 23613
rect 30193 23647 30251 23653
rect 30193 23613 30205 23647
rect 30239 23644 30251 23647
rect 31662 23644 31668 23656
rect 30239 23616 30788 23644
rect 31623 23616 31668 23644
rect 30239 23613 30251 23616
rect 30193 23607 30251 23613
rect 22336 23548 24072 23576
rect 26789 23579 26847 23585
rect 22336 23536 22342 23548
rect 26789 23545 26801 23579
rect 26835 23576 26847 23579
rect 28350 23576 28356 23588
rect 26835 23548 28356 23576
rect 26835 23545 26847 23548
rect 26789 23539 26847 23545
rect 28350 23536 28356 23548
rect 28408 23536 28414 23588
rect 29641 23579 29699 23585
rect 29641 23545 29653 23579
rect 29687 23576 29699 23579
rect 30760 23576 30788 23616
rect 31662 23604 31668 23616
rect 31720 23604 31726 23656
rect 32953 23647 33011 23653
rect 32953 23613 32965 23647
rect 32999 23644 33011 23647
rect 33226 23644 33232 23656
rect 32999 23616 33232 23644
rect 32999 23613 33011 23616
rect 32953 23607 33011 23613
rect 33226 23604 33232 23616
rect 33284 23604 33290 23656
rect 33336 23653 33364 23752
rect 33962 23740 33968 23792
rect 34020 23780 34026 23792
rect 34020 23752 35112 23780
rect 34020 23740 34026 23752
rect 35084 23721 35112 23752
rect 35069 23715 35127 23721
rect 35069 23681 35081 23715
rect 35115 23712 35127 23715
rect 37274 23712 37280 23724
rect 35115 23684 37280 23712
rect 35115 23681 35127 23684
rect 35069 23675 35127 23681
rect 37274 23672 37280 23684
rect 37332 23712 37338 23724
rect 37461 23715 37519 23721
rect 37461 23712 37473 23715
rect 37332 23684 37473 23712
rect 37332 23672 37338 23684
rect 37461 23681 37473 23684
rect 37507 23681 37519 23715
rect 37461 23675 37519 23681
rect 33321 23647 33379 23653
rect 33321 23613 33333 23647
rect 33367 23613 33379 23647
rect 33321 23607 33379 23613
rect 33413 23647 33471 23653
rect 33413 23613 33425 23647
rect 33459 23613 33471 23647
rect 33413 23607 33471 23613
rect 33965 23647 34023 23653
rect 33965 23613 33977 23647
rect 34011 23644 34023 23647
rect 34146 23644 34152 23656
rect 34011 23616 34152 23644
rect 34011 23613 34023 23616
rect 33965 23607 34023 23613
rect 31478 23576 31484 23588
rect 29687 23548 30696 23576
rect 30760 23548 31484 23576
rect 29687 23545 29699 23548
rect 29641 23539 29699 23545
rect 13044 23480 16436 23508
rect 13044 23468 13050 23480
rect 27706 23468 27712 23520
rect 27764 23508 27770 23520
rect 28442 23508 28448 23520
rect 27764 23480 28448 23508
rect 27764 23468 27770 23480
rect 28442 23468 28448 23480
rect 28500 23468 28506 23520
rect 30282 23508 30288 23520
rect 30243 23480 30288 23508
rect 30282 23468 30288 23480
rect 30340 23468 30346 23520
rect 30668 23508 30696 23548
rect 31478 23536 31484 23548
rect 31536 23576 31542 23588
rect 32582 23576 32588 23588
rect 31536 23548 32588 23576
rect 31536 23536 31542 23548
rect 32582 23536 32588 23548
rect 32640 23536 32646 23588
rect 32766 23536 32772 23588
rect 32824 23576 32830 23588
rect 33428 23576 33456 23607
rect 34146 23604 34152 23616
rect 34204 23604 34210 23656
rect 35345 23647 35403 23653
rect 35345 23613 35357 23647
rect 35391 23644 35403 23647
rect 35986 23644 35992 23656
rect 35391 23616 35992 23644
rect 35391 23613 35403 23616
rect 35345 23607 35403 23613
rect 35986 23604 35992 23616
rect 36044 23604 36050 23656
rect 37734 23644 37740 23656
rect 37695 23616 37740 23644
rect 37734 23604 37740 23616
rect 37792 23604 37798 23656
rect 32824 23548 33456 23576
rect 32824 23536 32830 23548
rect 32030 23508 32036 23520
rect 30668 23480 32036 23508
rect 32030 23468 32036 23480
rect 32088 23468 32094 23520
rect 34054 23468 34060 23520
rect 34112 23508 34118 23520
rect 34149 23511 34207 23517
rect 34149 23508 34161 23511
rect 34112 23480 34161 23508
rect 34112 23468 34118 23480
rect 34149 23477 34161 23480
rect 34195 23477 34207 23511
rect 34149 23471 34207 23477
rect 36354 23468 36360 23520
rect 36412 23508 36418 23520
rect 36449 23511 36507 23517
rect 36449 23508 36461 23511
rect 36412 23480 36461 23508
rect 36412 23468 36418 23480
rect 36449 23477 36461 23480
rect 36495 23477 36507 23511
rect 36449 23471 36507 23477
rect 1104 23418 39836 23440
rect 1104 23366 19606 23418
rect 19658 23366 19670 23418
rect 19722 23366 19734 23418
rect 19786 23366 19798 23418
rect 19850 23366 39836 23418
rect 1104 23344 39836 23366
rect 5169 23307 5227 23313
rect 5169 23273 5181 23307
rect 5215 23304 5227 23307
rect 5442 23304 5448 23316
rect 5215 23276 5448 23304
rect 5215 23273 5227 23276
rect 5169 23267 5227 23273
rect 5442 23264 5448 23276
rect 5500 23264 5506 23316
rect 7834 23264 7840 23316
rect 7892 23304 7898 23316
rect 8757 23307 8815 23313
rect 8757 23304 8769 23307
rect 7892 23276 8769 23304
rect 7892 23264 7898 23276
rect 8757 23273 8769 23276
rect 8803 23273 8815 23307
rect 9766 23304 9772 23316
rect 9727 23276 9772 23304
rect 8757 23267 8815 23273
rect 3145 23239 3203 23245
rect 3145 23205 3157 23239
rect 3191 23236 3203 23239
rect 3970 23236 3976 23248
rect 3191 23208 3976 23236
rect 3191 23205 3203 23208
rect 3145 23199 3203 23205
rect 3970 23196 3976 23208
rect 4028 23196 4034 23248
rect 1486 23168 1492 23180
rect 1447 23140 1492 23168
rect 1486 23128 1492 23140
rect 1544 23128 1550 23180
rect 1765 23171 1823 23177
rect 1765 23137 1777 23171
rect 1811 23168 1823 23171
rect 1854 23168 1860 23180
rect 1811 23140 1860 23168
rect 1811 23137 1823 23140
rect 1765 23131 1823 23137
rect 1854 23128 1860 23140
rect 1912 23128 1918 23180
rect 3418 23128 3424 23180
rect 3476 23168 3482 23180
rect 4065 23171 4123 23177
rect 4065 23168 4077 23171
rect 3476 23140 4077 23168
rect 3476 23128 3482 23140
rect 4065 23137 4077 23140
rect 4111 23137 4123 23171
rect 4890 23168 4896 23180
rect 4851 23140 4896 23168
rect 4065 23131 4123 23137
rect 4890 23128 4896 23140
rect 4948 23128 4954 23180
rect 5074 23168 5080 23180
rect 5035 23140 5080 23168
rect 5074 23128 5080 23140
rect 5132 23128 5138 23180
rect 5994 23168 6000 23180
rect 5955 23140 6000 23168
rect 5994 23128 6000 23140
rect 6052 23128 6058 23180
rect 6549 23171 6607 23177
rect 6549 23137 6561 23171
rect 6595 23168 6607 23171
rect 6638 23168 6644 23180
rect 6595 23140 6644 23168
rect 6595 23137 6607 23140
rect 6549 23131 6607 23137
rect 6638 23128 6644 23140
rect 6696 23128 6702 23180
rect 7193 23171 7251 23177
rect 7193 23137 7205 23171
rect 7239 23168 7251 23171
rect 7374 23168 7380 23180
rect 7239 23140 7380 23168
rect 7239 23137 7251 23140
rect 7193 23131 7251 23137
rect 7374 23128 7380 23140
rect 7432 23128 7438 23180
rect 7834 23168 7840 23180
rect 7795 23140 7840 23168
rect 7834 23128 7840 23140
rect 7892 23128 7898 23180
rect 8573 23171 8631 23177
rect 8573 23137 8585 23171
rect 8619 23168 8631 23171
rect 8662 23168 8668 23180
rect 8619 23140 8668 23168
rect 8619 23137 8631 23140
rect 8573 23131 8631 23137
rect 8662 23128 8668 23140
rect 8720 23128 8726 23180
rect 8772 23168 8800 23267
rect 9766 23264 9772 23276
rect 9824 23264 9830 23316
rect 10594 23264 10600 23316
rect 10652 23304 10658 23316
rect 17497 23307 17555 23313
rect 10652 23276 14320 23304
rect 10652 23264 10658 23276
rect 9030 23196 9036 23248
rect 9088 23236 9094 23248
rect 14292 23236 14320 23276
rect 17497 23273 17509 23307
rect 17543 23304 17555 23307
rect 19426 23304 19432 23316
rect 17543 23276 19432 23304
rect 17543 23273 17555 23276
rect 17497 23267 17555 23273
rect 19426 23264 19432 23276
rect 19484 23264 19490 23316
rect 21450 23264 21456 23316
rect 21508 23304 21514 23316
rect 21726 23304 21732 23316
rect 21508 23276 21732 23304
rect 21508 23264 21514 23276
rect 21726 23264 21732 23276
rect 21784 23264 21790 23316
rect 22373 23307 22431 23313
rect 22373 23273 22385 23307
rect 22419 23304 22431 23307
rect 22554 23304 22560 23316
rect 22419 23276 22560 23304
rect 22419 23273 22431 23276
rect 22373 23267 22431 23273
rect 22554 23264 22560 23276
rect 22612 23264 22618 23316
rect 24305 23307 24363 23313
rect 24305 23273 24317 23307
rect 24351 23304 24363 23307
rect 24394 23304 24400 23316
rect 24351 23276 24400 23304
rect 24351 23273 24363 23276
rect 24305 23267 24363 23273
rect 24394 23264 24400 23276
rect 24452 23264 24458 23316
rect 26234 23264 26240 23316
rect 26292 23304 26298 23316
rect 26605 23307 26663 23313
rect 26605 23304 26617 23307
rect 26292 23276 26617 23304
rect 26292 23264 26298 23276
rect 26605 23273 26617 23276
rect 26651 23273 26663 23307
rect 28166 23304 28172 23316
rect 28127 23276 28172 23304
rect 26605 23267 26663 23273
rect 28166 23264 28172 23276
rect 28224 23264 28230 23316
rect 30834 23304 30840 23316
rect 30795 23276 30840 23304
rect 30834 23264 30840 23276
rect 30892 23264 30898 23316
rect 32214 23304 32220 23316
rect 32175 23276 32220 23304
rect 32214 23264 32220 23276
rect 32272 23264 32278 23316
rect 33686 23304 33692 23316
rect 33599 23276 33692 23304
rect 33686 23264 33692 23276
rect 33744 23304 33750 23316
rect 33962 23304 33968 23316
rect 33744 23276 33968 23304
rect 33744 23264 33750 23276
rect 33962 23264 33968 23276
rect 34020 23264 34026 23316
rect 35897 23307 35955 23313
rect 35897 23273 35909 23307
rect 35943 23304 35955 23307
rect 35986 23304 35992 23316
rect 35943 23276 35992 23304
rect 35943 23273 35955 23276
rect 35897 23267 35955 23273
rect 35986 23264 35992 23276
rect 36044 23264 36050 23316
rect 19705 23239 19763 23245
rect 9088 23208 12296 23236
rect 9088 23196 9094 23208
rect 9398 23168 9404 23180
rect 8772 23140 9404 23168
rect 9398 23128 9404 23140
rect 9456 23168 9462 23180
rect 10336 23177 10364 23208
rect 9677 23171 9735 23177
rect 9677 23168 9689 23171
rect 9456 23140 9689 23168
rect 9456 23128 9462 23140
rect 9677 23137 9689 23140
rect 9723 23137 9735 23171
rect 9677 23131 9735 23137
rect 10321 23171 10379 23177
rect 10321 23137 10333 23171
rect 10367 23137 10379 23171
rect 10502 23168 10508 23180
rect 10463 23140 10508 23168
rect 10321 23131 10379 23137
rect 10502 23128 10508 23140
rect 10560 23168 10566 23180
rect 11422 23168 11428 23180
rect 10560 23140 11428 23168
rect 10560 23128 10566 23140
rect 11422 23128 11428 23140
rect 11480 23168 11486 23180
rect 11517 23171 11575 23177
rect 11517 23168 11529 23171
rect 11480 23140 11529 23168
rect 11480 23128 11486 23140
rect 11517 23137 11529 23140
rect 11563 23137 11575 23171
rect 12066 23168 12072 23180
rect 12027 23140 12072 23168
rect 11517 23131 11575 23137
rect 12066 23128 12072 23140
rect 12124 23128 12130 23180
rect 12268 23168 12296 23208
rect 14292 23208 19012 23236
rect 12342 23168 12348 23180
rect 12268 23140 12348 23168
rect 12342 23128 12348 23140
rect 12400 23128 12406 23180
rect 13722 23168 13728 23180
rect 13683 23140 13728 23168
rect 13722 23128 13728 23140
rect 13780 23128 13786 23180
rect 13909 23171 13967 23177
rect 13909 23137 13921 23171
rect 13955 23137 13967 23171
rect 13909 23131 13967 23137
rect 14093 23171 14151 23177
rect 14093 23137 14105 23171
rect 14139 23168 14151 23171
rect 14182 23168 14188 23180
rect 14139 23140 14188 23168
rect 14139 23137 14151 23140
rect 14093 23131 14151 23137
rect 5813 23103 5871 23109
rect 5813 23069 5825 23103
rect 5859 23100 5871 23103
rect 6730 23100 6736 23112
rect 5859 23072 5948 23100
rect 6691 23072 6736 23100
rect 5859 23069 5871 23072
rect 5813 23063 5871 23069
rect 5920 22976 5948 23072
rect 6730 23060 6736 23072
rect 6788 23060 6794 23112
rect 12434 23100 12440 23112
rect 12395 23072 12440 23100
rect 12434 23060 12440 23072
rect 12492 23060 12498 23112
rect 13170 23100 13176 23112
rect 13131 23072 13176 23100
rect 13170 23060 13176 23072
rect 13228 23060 13234 23112
rect 13924 23100 13952 23131
rect 14182 23128 14188 23140
rect 14240 23128 14246 23180
rect 14292 23177 14320 23208
rect 14277 23171 14335 23177
rect 14277 23137 14289 23171
rect 14323 23137 14335 23171
rect 14277 23131 14335 23137
rect 14553 23171 14611 23177
rect 14553 23137 14565 23171
rect 14599 23168 14611 23171
rect 15286 23168 15292 23180
rect 14599 23140 15292 23168
rect 14599 23137 14611 23140
rect 14553 23131 14611 23137
rect 15286 23128 15292 23140
rect 15344 23128 15350 23180
rect 15381 23171 15439 23177
rect 15381 23137 15393 23171
rect 15427 23168 15439 23171
rect 16482 23168 16488 23180
rect 15427 23140 16344 23168
rect 16443 23140 16488 23168
rect 15427 23137 15439 23140
rect 15381 23131 15439 23137
rect 15194 23100 15200 23112
rect 13924 23072 15200 23100
rect 15194 23060 15200 23072
rect 15252 23060 15258 23112
rect 16114 23100 16120 23112
rect 16075 23072 16120 23100
rect 16114 23060 16120 23072
rect 16172 23060 16178 23112
rect 16316 23100 16344 23140
rect 16482 23128 16488 23140
rect 16540 23128 16546 23180
rect 16574 23128 16580 23180
rect 16632 23128 16638 23180
rect 16666 23128 16672 23180
rect 16724 23168 16730 23180
rect 16945 23171 17003 23177
rect 16724 23140 16769 23168
rect 16724 23128 16730 23140
rect 16945 23137 16957 23171
rect 16991 23137 17003 23171
rect 16945 23131 17003 23137
rect 17129 23171 17187 23177
rect 17129 23137 17141 23171
rect 17175 23168 17187 23171
rect 17218 23168 17224 23180
rect 17175 23140 17224 23168
rect 17175 23137 17187 23140
rect 17129 23131 17187 23137
rect 16592 23100 16620 23128
rect 16316 23072 16620 23100
rect 16960 23100 16988 23131
rect 17218 23128 17224 23140
rect 17276 23128 17282 23180
rect 17862 23128 17868 23180
rect 17920 23168 17926 23180
rect 18233 23171 18291 23177
rect 18233 23168 18245 23171
rect 17920 23140 18245 23168
rect 17920 23128 17926 23140
rect 18233 23137 18245 23140
rect 18279 23137 18291 23171
rect 18598 23168 18604 23180
rect 18559 23140 18604 23168
rect 18233 23131 18291 23137
rect 18598 23128 18604 23140
rect 18656 23128 18662 23180
rect 18782 23168 18788 23180
rect 18743 23140 18788 23168
rect 18782 23128 18788 23140
rect 18840 23128 18846 23180
rect 18984 23177 19012 23208
rect 19705 23205 19717 23239
rect 19751 23236 19763 23239
rect 19978 23236 19984 23248
rect 19751 23208 19984 23236
rect 19751 23205 19763 23208
rect 19705 23199 19763 23205
rect 19978 23196 19984 23208
rect 20036 23196 20042 23248
rect 22646 23236 22652 23248
rect 20180 23208 22652 23236
rect 18969 23171 19027 23177
rect 18969 23137 18981 23171
rect 19015 23137 19027 23171
rect 19150 23168 19156 23180
rect 19111 23140 19156 23168
rect 18969 23131 19027 23137
rect 19150 23128 19156 23140
rect 19208 23128 19214 23180
rect 20180 23177 20208 23208
rect 22646 23196 22652 23208
rect 22704 23196 22710 23248
rect 27614 23236 27620 23248
rect 25332 23208 27620 23236
rect 20165 23171 20223 23177
rect 20165 23137 20177 23171
rect 20211 23137 20223 23171
rect 20165 23131 20223 23137
rect 20898 23128 20904 23180
rect 20956 23168 20962 23180
rect 21085 23171 21143 23177
rect 21085 23168 21097 23171
rect 20956 23140 21097 23168
rect 20956 23128 20962 23140
rect 21085 23137 21097 23140
rect 21131 23137 21143 23171
rect 21085 23131 21143 23137
rect 21545 23171 21603 23177
rect 21545 23137 21557 23171
rect 21591 23168 21603 23171
rect 21818 23168 21824 23180
rect 21591 23140 21824 23168
rect 21591 23137 21603 23140
rect 21545 23131 21603 23137
rect 18138 23100 18144 23112
rect 16960 23072 18144 23100
rect 18138 23060 18144 23072
rect 18196 23060 18202 23112
rect 20714 23060 20720 23112
rect 20772 23100 20778 23112
rect 21634 23100 21640 23112
rect 20772 23072 21640 23100
rect 20772 23060 20778 23072
rect 21634 23060 21640 23072
rect 21692 23060 21698 23112
rect 7190 22992 7196 23044
rect 7248 23032 7254 23044
rect 8021 23035 8079 23041
rect 8021 23032 8033 23035
rect 7248 23004 8033 23032
rect 7248 22992 7254 23004
rect 8021 23001 8033 23004
rect 8067 23001 8079 23035
rect 8021 22995 8079 23001
rect 20257 23035 20315 23041
rect 20257 23001 20269 23035
rect 20303 23032 20315 23035
rect 21744 23032 21772 23140
rect 21818 23128 21824 23140
rect 21876 23128 21882 23180
rect 22278 23168 22284 23180
rect 22239 23140 22284 23168
rect 22278 23128 22284 23140
rect 22336 23128 22342 23180
rect 22925 23171 22983 23177
rect 22925 23137 22937 23171
rect 22971 23168 22983 23171
rect 23474 23168 23480 23180
rect 22971 23140 23480 23168
rect 22971 23137 22983 23140
rect 22925 23131 22983 23137
rect 20303 23004 21772 23032
rect 20303 23001 20315 23004
rect 20257 22995 20315 23001
rect 5902 22964 5908 22976
rect 5815 22936 5908 22964
rect 5902 22924 5908 22936
rect 5960 22964 5966 22976
rect 7285 22967 7343 22973
rect 7285 22964 7297 22967
rect 5960 22936 7297 22964
rect 5960 22924 5966 22936
rect 7285 22933 7297 22936
rect 7331 22964 7343 22967
rect 7466 22964 7472 22976
rect 7331 22936 7472 22964
rect 7331 22933 7343 22936
rect 7285 22927 7343 22933
rect 7466 22924 7472 22936
rect 7524 22924 7530 22976
rect 11422 22924 11428 22976
rect 11480 22964 11486 22976
rect 14182 22964 14188 22976
rect 11480 22936 14188 22964
rect 11480 22924 11486 22936
rect 14182 22924 14188 22936
rect 14240 22924 14246 22976
rect 15565 22967 15623 22973
rect 15565 22933 15577 22967
rect 15611 22964 15623 22967
rect 16666 22964 16672 22976
rect 15611 22936 16672 22964
rect 15611 22933 15623 22936
rect 15565 22927 15623 22933
rect 16666 22924 16672 22936
rect 16724 22924 16730 22976
rect 21358 22924 21364 22976
rect 21416 22964 21422 22976
rect 22940 22964 22968 23131
rect 23474 23128 23480 23140
rect 23532 23128 23538 23180
rect 24210 23128 24216 23180
rect 24268 23168 24274 23180
rect 25332 23177 25360 23208
rect 27614 23196 27620 23208
rect 27672 23196 27678 23248
rect 31754 23196 31760 23248
rect 31812 23236 31818 23248
rect 34149 23239 34207 23245
rect 31812 23208 33916 23236
rect 31812 23196 31818 23208
rect 25317 23171 25375 23177
rect 25317 23168 25329 23171
rect 24268 23140 25329 23168
rect 24268 23128 24274 23140
rect 25317 23137 25329 23140
rect 25363 23137 25375 23171
rect 25317 23131 25375 23137
rect 25406 23128 25412 23180
rect 25464 23168 25470 23180
rect 25593 23171 25651 23177
rect 25593 23168 25605 23171
rect 25464 23140 25605 23168
rect 25464 23128 25470 23140
rect 25593 23137 25605 23140
rect 25639 23137 25651 23171
rect 25593 23131 25651 23137
rect 25961 23171 26019 23177
rect 25961 23137 25973 23171
rect 26007 23168 26019 23171
rect 26418 23168 26424 23180
rect 26007 23140 26424 23168
rect 26007 23137 26019 23140
rect 25961 23131 26019 23137
rect 26418 23128 26424 23140
rect 26476 23128 26482 23180
rect 26789 23171 26847 23177
rect 26789 23137 26801 23171
rect 26835 23168 26847 23171
rect 27062 23168 27068 23180
rect 26835 23140 27068 23168
rect 26835 23137 26847 23140
rect 26789 23131 26847 23137
rect 27062 23128 27068 23140
rect 27120 23128 27126 23180
rect 27341 23171 27399 23177
rect 27341 23168 27353 23171
rect 27172 23140 27353 23168
rect 23201 23103 23259 23109
rect 23201 23069 23213 23103
rect 23247 23100 23259 23103
rect 23566 23100 23572 23112
rect 23247 23072 23572 23100
rect 23247 23069 23259 23072
rect 23201 23063 23259 23069
rect 23566 23060 23572 23072
rect 23624 23060 23630 23112
rect 23658 23060 23664 23112
rect 23716 23100 23722 23112
rect 27172 23100 27200 23140
rect 27341 23137 27353 23140
rect 27387 23137 27399 23171
rect 27341 23131 27399 23137
rect 27522 23128 27528 23180
rect 27580 23168 27586 23180
rect 28077 23171 28135 23177
rect 28077 23168 28089 23171
rect 27580 23140 28089 23168
rect 27580 23128 27586 23140
rect 28077 23137 28089 23140
rect 28123 23137 28135 23171
rect 28077 23131 28135 23137
rect 28350 23128 28356 23180
rect 28408 23168 28414 23180
rect 28629 23171 28687 23177
rect 28629 23168 28641 23171
rect 28408 23140 28641 23168
rect 28408 23128 28414 23140
rect 28629 23137 28641 23140
rect 28675 23137 28687 23171
rect 28629 23131 28687 23137
rect 30193 23171 30251 23177
rect 30193 23137 30205 23171
rect 30239 23137 30251 23171
rect 30193 23131 30251 23137
rect 23716 23072 27200 23100
rect 23716 23060 23722 23072
rect 27246 23060 27252 23112
rect 27304 23100 27310 23112
rect 28905 23103 28963 23109
rect 28905 23100 28917 23103
rect 27304 23072 27349 23100
rect 28368 23072 28917 23100
rect 27304 23060 27310 23072
rect 28368 23044 28396 23072
rect 28905 23069 28917 23072
rect 28951 23069 28963 23103
rect 30208 23100 30236 23131
rect 30282 23128 30288 23180
rect 30340 23168 30346 23180
rect 30745 23171 30803 23177
rect 30745 23168 30757 23171
rect 30340 23140 30757 23168
rect 30340 23128 30346 23140
rect 30745 23137 30757 23140
rect 30791 23137 30803 23171
rect 30745 23131 30803 23137
rect 30929 23171 30987 23177
rect 30929 23137 30941 23171
rect 30975 23168 30987 23171
rect 31662 23168 31668 23180
rect 30975 23140 31668 23168
rect 30975 23137 30987 23140
rect 30929 23131 30987 23137
rect 31662 23128 31668 23140
rect 31720 23128 31726 23180
rect 31846 23128 31852 23180
rect 31904 23168 31910 23180
rect 31941 23171 31999 23177
rect 31941 23168 31953 23171
rect 31904 23140 31953 23168
rect 31904 23128 31910 23140
rect 31941 23137 31953 23140
rect 31987 23137 31999 23171
rect 32122 23168 32128 23180
rect 32083 23140 32128 23168
rect 31941 23131 31999 23137
rect 32122 23128 32128 23140
rect 32180 23128 32186 23180
rect 32582 23168 32588 23180
rect 32543 23140 32588 23168
rect 32582 23128 32588 23140
rect 32640 23128 32646 23180
rect 32953 23171 33011 23177
rect 32953 23137 32965 23171
rect 32999 23168 33011 23171
rect 33502 23168 33508 23180
rect 32999 23140 33508 23168
rect 32999 23137 33011 23140
rect 32953 23131 33011 23137
rect 30466 23100 30472 23112
rect 30208 23072 30472 23100
rect 28905 23063 28963 23069
rect 30466 23060 30472 23072
rect 30524 23060 30530 23112
rect 32030 23060 32036 23112
rect 32088 23100 32094 23112
rect 32968 23100 32996 23131
rect 33502 23128 33508 23140
rect 33560 23128 33566 23180
rect 33888 23177 33916 23208
rect 34149 23205 34161 23239
rect 34195 23236 34207 23239
rect 34238 23236 34244 23248
rect 34195 23208 34244 23236
rect 34195 23205 34207 23208
rect 34149 23199 34207 23205
rect 34238 23196 34244 23208
rect 34296 23196 34302 23248
rect 36354 23236 36360 23248
rect 35360 23208 36360 23236
rect 33873 23171 33931 23177
rect 33873 23137 33885 23171
rect 33919 23137 33931 23171
rect 33873 23131 33931 23137
rect 34793 23171 34851 23177
rect 34793 23137 34805 23171
rect 34839 23137 34851 23171
rect 34793 23131 34851 23137
rect 35161 23171 35219 23177
rect 35161 23137 35173 23171
rect 35207 23168 35219 23171
rect 35250 23168 35256 23180
rect 35207 23140 35256 23168
rect 35207 23137 35219 23140
rect 35161 23131 35219 23137
rect 32088 23072 32996 23100
rect 32088 23060 32094 23072
rect 33226 23060 33232 23112
rect 33284 23100 33290 23112
rect 34808 23100 34836 23131
rect 35250 23128 35256 23140
rect 35308 23128 35314 23180
rect 35360 23177 35388 23208
rect 36354 23196 36360 23208
rect 36412 23196 36418 23248
rect 35345 23171 35403 23177
rect 35345 23137 35357 23171
rect 35391 23137 35403 23171
rect 35345 23131 35403 23137
rect 35805 23171 35863 23177
rect 35805 23137 35817 23171
rect 35851 23137 35863 23171
rect 36446 23168 36452 23180
rect 36407 23140 36452 23168
rect 35805 23131 35863 23137
rect 33284 23072 34836 23100
rect 34885 23103 34943 23109
rect 33284 23060 33290 23072
rect 34885 23069 34897 23103
rect 34931 23100 34943 23103
rect 35434 23100 35440 23112
rect 34931 23072 35440 23100
rect 34931 23069 34943 23072
rect 34885 23063 34943 23069
rect 35434 23060 35440 23072
rect 35492 23060 35498 23112
rect 28350 22992 28356 23044
rect 28408 22992 28414 23044
rect 33318 22992 33324 23044
rect 33376 23032 33382 23044
rect 35820 23032 35848 23131
rect 36446 23128 36452 23140
rect 36504 23128 36510 23180
rect 38010 23168 38016 23180
rect 37971 23140 38016 23168
rect 38010 23128 38016 23140
rect 38068 23128 38074 23180
rect 38286 23168 38292 23180
rect 38247 23140 38292 23168
rect 38286 23128 38292 23140
rect 38344 23128 38350 23180
rect 38933 23171 38991 23177
rect 38933 23137 38945 23171
rect 38979 23137 38991 23171
rect 38933 23131 38991 23137
rect 36630 23100 36636 23112
rect 36591 23072 36636 23100
rect 36630 23060 36636 23072
rect 36688 23060 36694 23112
rect 36814 23060 36820 23112
rect 36872 23100 36878 23112
rect 38948 23100 38976 23131
rect 36872 23072 38976 23100
rect 36872 23060 36878 23072
rect 33376 23004 35848 23032
rect 33376 22992 33382 23004
rect 37734 22992 37740 23044
rect 37792 23032 37798 23044
rect 37829 23035 37887 23041
rect 37829 23032 37841 23035
rect 37792 23004 37841 23032
rect 37792 22992 37798 23004
rect 37829 23001 37841 23004
rect 37875 23001 37887 23035
rect 37829 22995 37887 23001
rect 31754 22964 31760 22976
rect 21416 22936 22968 22964
rect 31715 22936 31760 22964
rect 21416 22924 21422 22936
rect 31754 22924 31760 22936
rect 31812 22924 31818 22976
rect 35434 22924 35440 22976
rect 35492 22964 35498 22976
rect 36538 22964 36544 22976
rect 35492 22936 36544 22964
rect 35492 22924 35498 22936
rect 36538 22924 36544 22936
rect 36596 22924 36602 22976
rect 39022 22964 39028 22976
rect 38983 22936 39028 22964
rect 39022 22924 39028 22936
rect 39080 22924 39086 22976
rect 1104 22874 39836 22896
rect 1104 22822 4246 22874
rect 4298 22822 4310 22874
rect 4362 22822 4374 22874
rect 4426 22822 4438 22874
rect 4490 22822 34966 22874
rect 35018 22822 35030 22874
rect 35082 22822 35094 22874
rect 35146 22822 35158 22874
rect 35210 22822 39836 22874
rect 1104 22800 39836 22822
rect 5074 22720 5080 22772
rect 5132 22760 5138 22772
rect 6917 22763 6975 22769
rect 6917 22760 6929 22763
rect 5132 22732 6929 22760
rect 5132 22720 5138 22732
rect 6917 22729 6929 22732
rect 6963 22729 6975 22763
rect 6917 22723 6975 22729
rect 11701 22763 11759 22769
rect 11701 22729 11713 22763
rect 11747 22760 11759 22763
rect 12618 22760 12624 22772
rect 11747 22732 12624 22760
rect 11747 22729 11759 22732
rect 11701 22723 11759 22729
rect 12618 22720 12624 22732
rect 12676 22720 12682 22772
rect 17218 22720 17224 22772
rect 17276 22760 17282 22772
rect 18233 22763 18291 22769
rect 18233 22760 18245 22763
rect 17276 22732 18245 22760
rect 17276 22720 17282 22732
rect 18233 22729 18245 22732
rect 18279 22729 18291 22763
rect 18966 22760 18972 22772
rect 18927 22732 18972 22760
rect 18233 22723 18291 22729
rect 18966 22720 18972 22732
rect 19024 22720 19030 22772
rect 22278 22720 22284 22772
rect 22336 22760 22342 22772
rect 22741 22763 22799 22769
rect 22741 22760 22753 22763
rect 22336 22732 22753 22760
rect 22336 22720 22342 22732
rect 22741 22729 22753 22732
rect 22787 22729 22799 22763
rect 22741 22723 22799 22729
rect 25961 22763 26019 22769
rect 25961 22729 25973 22763
rect 26007 22760 26019 22763
rect 26694 22760 26700 22772
rect 26007 22732 26700 22760
rect 26007 22729 26019 22732
rect 25961 22723 26019 22729
rect 26694 22720 26700 22732
rect 26752 22720 26758 22772
rect 28905 22763 28963 22769
rect 28905 22729 28917 22763
rect 28951 22760 28963 22763
rect 28994 22760 29000 22772
rect 28951 22732 29000 22760
rect 28951 22729 28963 22732
rect 28905 22723 28963 22729
rect 28994 22720 29000 22732
rect 29052 22760 29058 22772
rect 29454 22760 29460 22772
rect 29052 22732 29460 22760
rect 29052 22720 29058 22732
rect 29454 22720 29460 22732
rect 29512 22720 29518 22772
rect 30466 22720 30472 22772
rect 30524 22720 30530 22772
rect 31113 22763 31171 22769
rect 31113 22729 31125 22763
rect 31159 22760 31171 22763
rect 32122 22760 32128 22772
rect 31159 22732 32128 22760
rect 31159 22729 31171 22732
rect 31113 22723 31171 22729
rect 32122 22720 32128 22732
rect 32180 22720 32186 22772
rect 32398 22720 32404 22772
rect 32456 22760 32462 22772
rect 36630 22760 36636 22772
rect 32456 22732 36636 22760
rect 32456 22720 32462 22732
rect 36630 22720 36636 22732
rect 36688 22720 36694 22772
rect 36998 22720 37004 22772
rect 37056 22760 37062 22772
rect 38381 22763 38439 22769
rect 38381 22760 38393 22763
rect 37056 22732 38393 22760
rect 37056 22720 37062 22732
rect 38381 22729 38393 22732
rect 38427 22729 38439 22763
rect 38381 22723 38439 22729
rect 4798 22652 4804 22704
rect 4856 22692 4862 22704
rect 4893 22695 4951 22701
rect 4893 22692 4905 22695
rect 4856 22664 4905 22692
rect 4856 22652 4862 22664
rect 4893 22661 4905 22664
rect 4939 22661 4951 22695
rect 4893 22655 4951 22661
rect 2314 22584 2320 22636
rect 2372 22624 2378 22636
rect 2958 22624 2964 22636
rect 2372 22596 2964 22624
rect 2372 22584 2378 22596
rect 2958 22584 2964 22596
rect 3016 22584 3022 22636
rect 4614 22624 4620 22636
rect 4080 22596 4620 22624
rect 2133 22559 2191 22565
rect 2133 22525 2145 22559
rect 2179 22525 2191 22559
rect 2682 22556 2688 22568
rect 2595 22528 2688 22556
rect 2133 22519 2191 22525
rect 2148 22488 2176 22519
rect 2682 22516 2688 22528
rect 2740 22556 2746 22568
rect 3234 22556 3240 22568
rect 2740 22528 3240 22556
rect 2740 22516 2746 22528
rect 3234 22516 3240 22528
rect 3292 22516 3298 22568
rect 3418 22516 3424 22568
rect 3476 22556 3482 22568
rect 4080 22565 4108 22596
rect 4614 22584 4620 22596
rect 4672 22584 4678 22636
rect 5092 22624 5120 22720
rect 19886 22692 19892 22704
rect 19847 22664 19892 22692
rect 19886 22652 19892 22664
rect 19944 22652 19950 22704
rect 30484 22692 30512 22720
rect 31570 22692 31576 22704
rect 24872 22664 26832 22692
rect 30484 22664 31576 22692
rect 5902 22624 5908 22636
rect 4724 22596 5120 22624
rect 5552 22596 5908 22624
rect 3513 22559 3571 22565
rect 3513 22556 3525 22559
rect 3476 22528 3525 22556
rect 3476 22516 3482 22528
rect 3513 22525 3525 22528
rect 3559 22525 3571 22559
rect 3513 22519 3571 22525
rect 4065 22559 4123 22565
rect 4065 22525 4077 22559
rect 4111 22525 4123 22559
rect 4522 22556 4528 22568
rect 4435 22528 4528 22556
rect 4065 22519 4123 22525
rect 4522 22516 4528 22528
rect 4580 22556 4586 22568
rect 4724 22556 4752 22596
rect 4890 22556 4896 22568
rect 4580 22528 4752 22556
rect 4851 22528 4896 22556
rect 4580 22516 4586 22528
rect 4890 22516 4896 22528
rect 4948 22516 4954 22568
rect 5552 22565 5580 22596
rect 5902 22584 5908 22596
rect 5960 22584 5966 22636
rect 6178 22624 6184 22636
rect 6139 22596 6184 22624
rect 6178 22584 6184 22596
rect 6236 22584 6242 22636
rect 8021 22627 8079 22633
rect 8021 22593 8033 22627
rect 8067 22624 8079 22627
rect 9585 22627 9643 22633
rect 8067 22596 9536 22624
rect 8067 22593 8079 22596
rect 8021 22587 8079 22593
rect 5537 22559 5595 22565
rect 5537 22525 5549 22559
rect 5583 22525 5595 22559
rect 5537 22519 5595 22525
rect 5626 22516 5632 22568
rect 5684 22556 5690 22568
rect 5994 22556 6000 22568
rect 5684 22528 6000 22556
rect 5684 22516 5690 22528
rect 5994 22516 6000 22528
rect 6052 22516 6058 22568
rect 6822 22556 6828 22568
rect 6783 22528 6828 22556
rect 6822 22516 6828 22528
rect 6880 22516 6886 22568
rect 7374 22556 7380 22568
rect 7335 22528 7380 22556
rect 7374 22516 7380 22528
rect 7432 22516 7438 22568
rect 8294 22556 8300 22568
rect 8255 22528 8300 22556
rect 8294 22516 8300 22528
rect 8352 22516 8358 22568
rect 9508 22556 9536 22596
rect 9585 22593 9597 22627
rect 9631 22624 9643 22627
rect 10594 22624 10600 22636
rect 9631 22596 10600 22624
rect 9631 22593 9643 22596
rect 9585 22587 9643 22593
rect 10594 22584 10600 22596
rect 10652 22584 10658 22636
rect 13814 22624 13820 22636
rect 13727 22596 13820 22624
rect 13814 22584 13820 22596
rect 13872 22624 13878 22636
rect 13998 22624 14004 22636
rect 13872 22596 14004 22624
rect 13872 22584 13878 22596
rect 13998 22584 14004 22596
rect 14056 22584 14062 22636
rect 14182 22584 14188 22636
rect 14240 22624 14246 22636
rect 17494 22624 17500 22636
rect 14240 22596 16804 22624
rect 17455 22596 17500 22624
rect 14240 22584 14246 22596
rect 9950 22556 9956 22568
rect 9508 22528 9956 22556
rect 9950 22516 9956 22528
rect 10008 22556 10014 22568
rect 10137 22559 10195 22565
rect 10137 22556 10149 22559
rect 10008 22528 10149 22556
rect 10008 22516 10014 22528
rect 10137 22525 10149 22528
rect 10183 22525 10195 22559
rect 10410 22556 10416 22568
rect 10371 22528 10416 22556
rect 10137 22519 10195 22525
rect 10410 22516 10416 22528
rect 10468 22516 10474 22568
rect 11054 22516 11060 22568
rect 11112 22556 11118 22568
rect 12437 22559 12495 22565
rect 12437 22556 12449 22559
rect 11112 22528 12449 22556
rect 11112 22516 11118 22528
rect 12437 22525 12449 22528
rect 12483 22525 12495 22559
rect 12986 22556 12992 22568
rect 12947 22528 12992 22556
rect 12437 22519 12495 22525
rect 12986 22516 12992 22528
rect 13044 22516 13050 22568
rect 14093 22559 14151 22565
rect 14093 22525 14105 22559
rect 14139 22556 14151 22559
rect 15378 22556 15384 22568
rect 14139 22528 15384 22556
rect 14139 22525 14151 22528
rect 14093 22519 14151 22525
rect 15378 22516 15384 22528
rect 15436 22516 15442 22568
rect 16025 22559 16083 22565
rect 16025 22525 16037 22559
rect 16071 22556 16083 22559
rect 16114 22556 16120 22568
rect 16071 22528 16120 22556
rect 16071 22525 16083 22528
rect 16025 22519 16083 22525
rect 16114 22516 16120 22528
rect 16172 22516 16178 22568
rect 16393 22559 16451 22565
rect 16393 22525 16405 22559
rect 16439 22556 16451 22559
rect 16482 22556 16488 22568
rect 16439 22528 16488 22556
rect 16439 22525 16451 22528
rect 16393 22519 16451 22525
rect 16482 22516 16488 22528
rect 16540 22516 16546 22568
rect 16577 22559 16635 22565
rect 16577 22525 16589 22559
rect 16623 22556 16635 22559
rect 16666 22556 16672 22568
rect 16623 22528 16672 22556
rect 16623 22525 16635 22528
rect 16577 22519 16635 22525
rect 16666 22516 16672 22528
rect 16724 22516 16730 22568
rect 16776 22565 16804 22596
rect 17494 22584 17500 22596
rect 17552 22584 17558 22636
rect 23934 22624 23940 22636
rect 19996 22596 23940 22624
rect 16761 22559 16819 22565
rect 16761 22525 16773 22559
rect 16807 22525 16819 22559
rect 16761 22519 16819 22525
rect 17037 22559 17095 22565
rect 17037 22525 17049 22559
rect 17083 22556 17095 22559
rect 17218 22556 17224 22568
rect 17083 22528 17224 22556
rect 17083 22525 17095 22528
rect 17037 22519 17095 22525
rect 17218 22516 17224 22528
rect 17276 22516 17282 22568
rect 18046 22556 18052 22568
rect 18007 22528 18052 22556
rect 18046 22516 18052 22528
rect 18104 22516 18110 22568
rect 18782 22556 18788 22568
rect 18695 22528 18788 22556
rect 18782 22516 18788 22528
rect 18840 22516 18846 22568
rect 19996 22565 20024 22596
rect 23934 22584 23940 22596
rect 23992 22584 23998 22636
rect 24872 22568 24900 22664
rect 25317 22627 25375 22633
rect 25317 22593 25329 22627
rect 25363 22624 25375 22627
rect 25406 22624 25412 22636
rect 25363 22596 25412 22624
rect 25363 22593 25375 22596
rect 25317 22587 25375 22593
rect 25406 22584 25412 22596
rect 25464 22584 25470 22636
rect 26804 22624 26832 22664
rect 31570 22652 31576 22664
rect 31628 22692 31634 22704
rect 33781 22695 33839 22701
rect 33781 22692 33793 22695
rect 31628 22664 33793 22692
rect 31628 22652 31634 22664
rect 33781 22661 33793 22664
rect 33827 22661 33839 22695
rect 33781 22655 33839 22661
rect 35526 22652 35532 22704
rect 35584 22692 35590 22704
rect 36354 22692 36360 22704
rect 35584 22664 36360 22692
rect 35584 22652 35590 22664
rect 36354 22652 36360 22664
rect 36412 22652 36418 22704
rect 27246 22624 27252 22636
rect 26804 22596 27252 22624
rect 26804 22568 26832 22596
rect 27246 22584 27252 22596
rect 27304 22584 27310 22636
rect 31754 22624 31760 22636
rect 29104 22596 31760 22624
rect 19981 22559 20039 22565
rect 19981 22525 19993 22559
rect 20027 22525 20039 22559
rect 19981 22519 20039 22525
rect 20254 22516 20260 22568
rect 20312 22556 20318 22568
rect 20349 22559 20407 22565
rect 20349 22556 20361 22559
rect 20312 22528 20361 22556
rect 20312 22516 20318 22528
rect 20349 22525 20361 22528
rect 20395 22525 20407 22559
rect 20622 22556 20628 22568
rect 20583 22528 20628 22556
rect 20349 22519 20407 22525
rect 20622 22516 20628 22528
rect 20680 22516 20686 22568
rect 21358 22556 21364 22568
rect 21319 22528 21364 22556
rect 21358 22516 21364 22528
rect 21416 22516 21422 22568
rect 21634 22556 21640 22568
rect 21595 22528 21640 22556
rect 21634 22516 21640 22528
rect 21692 22516 21698 22568
rect 23658 22556 23664 22568
rect 23619 22528 23664 22556
rect 23658 22516 23664 22528
rect 23716 22516 23722 22568
rect 24854 22556 24860 22568
rect 24767 22528 24860 22556
rect 24854 22516 24860 22528
rect 24912 22516 24918 22568
rect 25225 22559 25283 22565
rect 25225 22525 25237 22559
rect 25271 22525 25283 22559
rect 26418 22556 26424 22568
rect 26379 22528 26424 22556
rect 25225 22519 25283 22525
rect 7834 22488 7840 22500
rect 2148 22460 7840 22488
rect 7834 22448 7840 22460
rect 7892 22448 7898 22500
rect 15473 22491 15531 22497
rect 15473 22457 15485 22491
rect 15519 22488 15531 22491
rect 17126 22488 17132 22500
rect 15519 22460 17132 22488
rect 15519 22457 15531 22460
rect 15473 22451 15531 22457
rect 2041 22423 2099 22429
rect 2041 22389 2053 22423
rect 2087 22420 2099 22423
rect 2958 22420 2964 22432
rect 2087 22392 2964 22420
rect 2087 22389 2099 22392
rect 2041 22383 2099 22389
rect 2958 22380 2964 22392
rect 3016 22380 3022 22432
rect 12342 22380 12348 22432
rect 12400 22420 12406 22432
rect 12529 22423 12587 22429
rect 12529 22420 12541 22423
rect 12400 22392 12541 22420
rect 12400 22380 12406 22392
rect 12529 22389 12541 22392
rect 12575 22389 12587 22423
rect 12529 22383 12587 22389
rect 13722 22380 13728 22432
rect 13780 22420 13786 22432
rect 15488 22420 15516 22451
rect 17126 22448 17132 22460
rect 17184 22448 17190 22500
rect 18800 22488 18828 22516
rect 20070 22488 20076 22500
rect 18800 22460 20076 22488
rect 20070 22448 20076 22460
rect 20128 22448 20134 22500
rect 24302 22448 24308 22500
rect 24360 22488 24366 22500
rect 24397 22491 24455 22497
rect 24397 22488 24409 22491
rect 24360 22460 24409 22488
rect 24360 22448 24366 22460
rect 24397 22457 24409 22460
rect 24443 22457 24455 22491
rect 24397 22451 24455 22457
rect 24578 22448 24584 22500
rect 24636 22488 24642 22500
rect 25240 22488 25268 22519
rect 26418 22516 26424 22528
rect 26476 22516 26482 22568
rect 26605 22559 26663 22565
rect 26605 22525 26617 22559
rect 26651 22556 26663 22559
rect 26651 22528 26740 22556
rect 26651 22525 26663 22528
rect 26605 22519 26663 22525
rect 24636 22460 25268 22488
rect 24636 22448 24642 22460
rect 13780 22392 15516 22420
rect 23845 22423 23903 22429
rect 13780 22380 13786 22392
rect 23845 22389 23857 22423
rect 23891 22420 23903 22423
rect 24210 22420 24216 22432
rect 23891 22392 24216 22420
rect 23891 22389 23903 22392
rect 23845 22383 23903 22389
rect 24210 22380 24216 22392
rect 24268 22380 24274 22432
rect 26712 22420 26740 22528
rect 26786 22516 26792 22568
rect 26844 22556 26850 22568
rect 27062 22556 27068 22568
rect 26844 22528 26937 22556
rect 27023 22528 27068 22556
rect 26844 22516 26850 22528
rect 27062 22516 27068 22528
rect 27120 22516 27126 22568
rect 27154 22516 27160 22568
rect 27212 22556 27218 22568
rect 27985 22559 28043 22565
rect 27212 22528 27257 22556
rect 27212 22516 27218 22528
rect 27985 22525 27997 22559
rect 28031 22556 28043 22559
rect 28258 22556 28264 22568
rect 28031 22528 28264 22556
rect 28031 22525 28043 22528
rect 27985 22519 28043 22525
rect 28258 22516 28264 22528
rect 28316 22516 28322 22568
rect 29104 22565 29132 22596
rect 31754 22584 31760 22596
rect 31812 22584 31818 22636
rect 32306 22624 32312 22636
rect 32267 22596 32312 22624
rect 32306 22584 32312 22596
rect 32364 22584 32370 22636
rect 34054 22584 34060 22636
rect 34112 22624 34118 22636
rect 34422 22624 34428 22636
rect 34112 22596 34428 22624
rect 34112 22584 34118 22596
rect 34422 22584 34428 22596
rect 34480 22624 34486 22636
rect 35897 22627 35955 22633
rect 34480 22596 35756 22624
rect 34480 22584 34486 22596
rect 29089 22559 29147 22565
rect 29089 22525 29101 22559
rect 29135 22525 29147 22559
rect 29089 22519 29147 22525
rect 29454 22516 29460 22568
rect 29512 22556 29518 22568
rect 29549 22559 29607 22565
rect 29549 22556 29561 22559
rect 29512 22528 29561 22556
rect 29512 22516 29518 22528
rect 29549 22525 29561 22528
rect 29595 22525 29607 22559
rect 29822 22556 29828 22568
rect 29783 22528 29828 22556
rect 29549 22519 29607 22525
rect 29822 22516 29828 22528
rect 29880 22516 29886 22568
rect 30282 22516 30288 22568
rect 30340 22556 30346 22568
rect 31665 22559 31723 22565
rect 31665 22556 31677 22559
rect 30340 22528 31677 22556
rect 30340 22516 30346 22528
rect 31665 22525 31677 22528
rect 31711 22525 31723 22559
rect 32030 22556 32036 22568
rect 31991 22528 32036 22556
rect 31665 22519 31723 22525
rect 32030 22516 32036 22528
rect 32088 22516 32094 22568
rect 32398 22556 32404 22568
rect 32359 22528 32404 22556
rect 32398 22516 32404 22528
rect 32456 22516 32462 22568
rect 32490 22516 32496 22568
rect 32548 22556 32554 22568
rect 32953 22559 33011 22565
rect 32953 22556 32965 22559
rect 32548 22528 32965 22556
rect 32548 22516 32554 22528
rect 32953 22525 32965 22528
rect 32999 22525 33011 22559
rect 33594 22556 33600 22568
rect 33555 22528 33600 22556
rect 32953 22519 33011 22525
rect 33594 22516 33600 22528
rect 33652 22516 33658 22568
rect 34885 22559 34943 22565
rect 34885 22525 34897 22559
rect 34931 22556 34943 22559
rect 35250 22556 35256 22568
rect 34931 22528 35256 22556
rect 34931 22525 34943 22528
rect 34885 22519 34943 22525
rect 35250 22516 35256 22528
rect 35308 22516 35314 22568
rect 26970 22448 26976 22500
rect 27028 22488 27034 22500
rect 27172 22488 27200 22516
rect 27028 22460 27200 22488
rect 27028 22448 27034 22460
rect 33962 22448 33968 22500
rect 34020 22488 34026 22500
rect 35728 22488 35756 22596
rect 35897 22593 35909 22627
rect 35943 22624 35955 22627
rect 37274 22624 37280 22636
rect 35943 22596 37280 22624
rect 35943 22593 35955 22596
rect 35897 22587 35955 22593
rect 37274 22584 37280 22596
rect 37332 22584 37338 22636
rect 37918 22624 37924 22636
rect 37831 22596 37924 22624
rect 37918 22584 37924 22596
rect 37976 22624 37982 22636
rect 38286 22624 38292 22636
rect 37976 22596 38292 22624
rect 37976 22584 37982 22596
rect 38286 22584 38292 22596
rect 38344 22584 38350 22636
rect 36170 22556 36176 22568
rect 36131 22528 36176 22556
rect 36170 22516 36176 22528
rect 36228 22516 36234 22568
rect 37093 22559 37151 22565
rect 37093 22556 37105 22559
rect 36280 22528 37105 22556
rect 36081 22491 36139 22497
rect 36081 22488 36093 22491
rect 34020 22460 35664 22488
rect 35728 22460 36093 22488
rect 34020 22448 34026 22460
rect 27614 22420 27620 22432
rect 26712 22392 27620 22420
rect 27614 22380 27620 22392
rect 27672 22380 27678 22432
rect 27890 22380 27896 22432
rect 27948 22420 27954 22432
rect 28169 22423 28227 22429
rect 28169 22420 28181 22423
rect 27948 22392 28181 22420
rect 27948 22380 27954 22392
rect 28169 22389 28181 22392
rect 28215 22389 28227 22423
rect 28169 22383 28227 22389
rect 28534 22380 28540 22432
rect 28592 22420 28598 22432
rect 31018 22420 31024 22432
rect 28592 22392 31024 22420
rect 28592 22380 28598 22392
rect 31018 22380 31024 22392
rect 31076 22380 31082 22432
rect 31662 22380 31668 22432
rect 31720 22420 31726 22432
rect 33778 22420 33784 22432
rect 31720 22392 33784 22420
rect 31720 22380 31726 22392
rect 33778 22380 33784 22392
rect 33836 22420 33842 22432
rect 35069 22423 35127 22429
rect 35069 22420 35081 22423
rect 33836 22392 35081 22420
rect 33836 22380 33842 22392
rect 35069 22389 35081 22392
rect 35115 22420 35127 22423
rect 35526 22420 35532 22432
rect 35115 22392 35532 22420
rect 35115 22389 35127 22392
rect 35069 22383 35127 22389
rect 35526 22380 35532 22392
rect 35584 22380 35590 22432
rect 35636 22420 35664 22460
rect 36081 22457 36093 22460
rect 36127 22457 36139 22491
rect 36081 22451 36139 22457
rect 36280 22420 36308 22528
rect 37093 22525 37105 22528
rect 37139 22525 37151 22559
rect 38102 22556 38108 22568
rect 38063 22528 38108 22556
rect 37093 22519 37151 22525
rect 38102 22516 38108 22528
rect 38160 22516 38166 22568
rect 38197 22559 38255 22565
rect 38197 22525 38209 22559
rect 38243 22556 38255 22559
rect 38562 22556 38568 22568
rect 38243 22528 38568 22556
rect 38243 22525 38255 22528
rect 38197 22519 38255 22525
rect 38562 22516 38568 22528
rect 38620 22516 38626 22568
rect 36633 22491 36691 22497
rect 36633 22457 36645 22491
rect 36679 22488 36691 22491
rect 37182 22488 37188 22500
rect 36679 22460 37188 22488
rect 36679 22457 36691 22460
rect 36633 22451 36691 22457
rect 37182 22448 37188 22460
rect 37240 22448 37246 22500
rect 35636 22392 36308 22420
rect 37277 22423 37335 22429
rect 37277 22389 37289 22423
rect 37323 22420 37335 22423
rect 37366 22420 37372 22432
rect 37323 22392 37372 22420
rect 37323 22389 37335 22392
rect 37277 22383 37335 22389
rect 37366 22380 37372 22392
rect 37424 22380 37430 22432
rect 1104 22330 39836 22352
rect 1104 22278 19606 22330
rect 19658 22278 19670 22330
rect 19722 22278 19734 22330
rect 19786 22278 19798 22330
rect 19850 22278 39836 22330
rect 1104 22256 39836 22278
rect 1581 22219 1639 22225
rect 1581 22185 1593 22219
rect 1627 22216 1639 22219
rect 2314 22216 2320 22228
rect 1627 22188 2320 22216
rect 1627 22185 1639 22188
rect 1581 22179 1639 22185
rect 2314 22176 2320 22188
rect 2372 22176 2378 22228
rect 3234 22176 3240 22228
rect 3292 22216 3298 22228
rect 4341 22219 4399 22225
rect 4341 22216 4353 22219
rect 3292 22188 4353 22216
rect 3292 22176 3298 22188
rect 4341 22185 4353 22188
rect 4387 22185 4399 22219
rect 7374 22216 7380 22228
rect 7335 22188 7380 22216
rect 4341 22179 4399 22185
rect 7374 22176 7380 22188
rect 7432 22176 7438 22228
rect 8294 22216 8300 22228
rect 8255 22188 8300 22216
rect 8294 22176 8300 22188
rect 8352 22176 8358 22228
rect 9769 22219 9827 22225
rect 9769 22185 9781 22219
rect 9815 22216 9827 22219
rect 10410 22216 10416 22228
rect 9815 22188 10416 22216
rect 9815 22185 9827 22188
rect 9769 22179 9827 22185
rect 10410 22176 10416 22188
rect 10468 22176 10474 22228
rect 11422 22216 11428 22228
rect 11383 22188 11428 22216
rect 11422 22176 11428 22188
rect 11480 22176 11486 22228
rect 14182 22176 14188 22228
rect 14240 22216 14246 22228
rect 15286 22216 15292 22228
rect 14240 22188 15292 22216
rect 14240 22176 14246 22188
rect 15286 22176 15292 22188
rect 15344 22176 15350 22228
rect 18966 22176 18972 22228
rect 19024 22216 19030 22228
rect 19150 22216 19156 22228
rect 19024 22188 19156 22216
rect 19024 22176 19030 22188
rect 19150 22176 19156 22188
rect 19208 22176 19214 22228
rect 25314 22216 25320 22228
rect 25275 22188 25320 22216
rect 25314 22176 25320 22188
rect 25372 22176 25378 22228
rect 26973 22219 27031 22225
rect 26973 22185 26985 22219
rect 27019 22216 27031 22219
rect 27522 22216 27528 22228
rect 27019 22188 27528 22216
rect 27019 22185 27031 22188
rect 26973 22179 27031 22185
rect 27522 22176 27528 22188
rect 27580 22176 27586 22228
rect 29822 22216 29828 22228
rect 29783 22188 29828 22216
rect 29822 22176 29828 22188
rect 29880 22176 29886 22228
rect 33226 22176 33232 22228
rect 33284 22216 33290 22228
rect 33321 22219 33379 22225
rect 33321 22216 33333 22219
rect 33284 22188 33333 22216
rect 33284 22176 33290 22188
rect 33321 22185 33333 22188
rect 33367 22185 33379 22219
rect 37826 22216 37832 22228
rect 37787 22188 37832 22216
rect 33321 22179 33379 22185
rect 37826 22176 37832 22188
rect 37884 22176 37890 22228
rect 12618 22148 12624 22160
rect 11256 22120 12624 22148
rect 1397 22083 1455 22089
rect 1397 22049 1409 22083
rect 1443 22049 1455 22083
rect 2314 22080 2320 22092
rect 2275 22052 2320 22080
rect 1397 22043 1455 22049
rect 1412 21876 1440 22043
rect 2314 22040 2320 22052
rect 2372 22040 2378 22092
rect 2682 22080 2688 22092
rect 2643 22052 2688 22080
rect 2682 22040 2688 22052
rect 2740 22040 2746 22092
rect 2958 22080 2964 22092
rect 2919 22052 2964 22080
rect 2958 22040 2964 22052
rect 3016 22040 3022 22092
rect 4522 22080 4528 22092
rect 4483 22052 4528 22080
rect 4522 22040 4528 22052
rect 4580 22040 4586 22092
rect 4801 22083 4859 22089
rect 4801 22049 4813 22083
rect 4847 22049 4859 22083
rect 4801 22043 4859 22049
rect 4816 22012 4844 22043
rect 4982 22040 4988 22092
rect 5040 22080 5046 22092
rect 5813 22083 5871 22089
rect 5813 22080 5825 22083
rect 5040 22052 5825 22080
rect 5040 22040 5046 22052
rect 5813 22049 5825 22052
rect 5859 22049 5871 22083
rect 8018 22080 8024 22092
rect 7979 22052 8024 22080
rect 5813 22043 5871 22049
rect 8018 22040 8024 22052
rect 8076 22040 8082 22092
rect 8846 22080 8852 22092
rect 8807 22052 8852 22080
rect 8846 22040 8852 22052
rect 8904 22040 8910 22092
rect 9030 22080 9036 22092
rect 8991 22052 9036 22080
rect 9030 22040 9036 22052
rect 9088 22040 9094 22092
rect 9674 22080 9680 22092
rect 9635 22052 9680 22080
rect 9674 22040 9680 22052
rect 9732 22040 9738 22092
rect 9950 22040 9956 22092
rect 10008 22080 10014 22092
rect 10594 22080 10600 22092
rect 10008 22052 10600 22080
rect 10008 22040 10014 22052
rect 10594 22040 10600 22052
rect 10652 22040 10658 22092
rect 10689 22083 10747 22089
rect 10689 22049 10701 22083
rect 10735 22080 10747 22083
rect 11054 22080 11060 22092
rect 10735 22052 11060 22080
rect 10735 22049 10747 22052
rect 10689 22043 10747 22049
rect 11054 22040 11060 22052
rect 11112 22040 11118 22092
rect 11256 22089 11284 22120
rect 12618 22108 12624 22120
rect 12676 22108 12682 22160
rect 14001 22151 14059 22157
rect 14001 22117 14013 22151
rect 14047 22148 14059 22151
rect 15194 22148 15200 22160
rect 14047 22120 15200 22148
rect 14047 22117 14059 22120
rect 14001 22111 14059 22117
rect 15194 22108 15200 22120
rect 15252 22148 15258 22160
rect 15381 22151 15439 22157
rect 15381 22148 15393 22151
rect 15252 22120 15393 22148
rect 15252 22108 15258 22120
rect 15381 22117 15393 22120
rect 15427 22117 15439 22151
rect 17862 22148 17868 22160
rect 15381 22111 15439 22117
rect 16408 22120 17868 22148
rect 11241 22083 11299 22089
rect 11241 22049 11253 22083
rect 11287 22049 11299 22083
rect 12434 22080 12440 22092
rect 12395 22052 12440 22080
rect 11241 22043 11299 22049
rect 12434 22040 12440 22052
rect 12492 22040 12498 22092
rect 12526 22040 12532 22092
rect 12584 22080 12590 22092
rect 12713 22083 12771 22089
rect 12713 22080 12725 22083
rect 12584 22052 12725 22080
rect 12584 22040 12590 22052
rect 12713 22049 12725 22052
rect 12759 22049 12771 22083
rect 13170 22080 13176 22092
rect 13131 22052 13176 22080
rect 12713 22043 12771 22049
rect 13170 22040 13176 22052
rect 13228 22040 13234 22092
rect 14182 22080 14188 22092
rect 14143 22052 14188 22080
rect 14182 22040 14188 22052
rect 14240 22040 14246 22092
rect 14550 22080 14556 22092
rect 14511 22052 14556 22080
rect 14550 22040 14556 22052
rect 14608 22040 14614 22092
rect 15289 22083 15347 22089
rect 15289 22049 15301 22083
rect 15335 22049 15347 22083
rect 15289 22043 15347 22049
rect 5534 22012 5540 22024
rect 4816 21984 5540 22012
rect 5534 21972 5540 21984
rect 5592 21972 5598 22024
rect 6089 22015 6147 22021
rect 6089 21981 6101 22015
rect 6135 22012 6147 22015
rect 6914 22012 6920 22024
rect 6135 21984 6920 22012
rect 6135 21981 6147 21984
rect 6089 21975 6147 21981
rect 6914 21972 6920 21984
rect 6972 21972 6978 22024
rect 7190 21972 7196 22024
rect 7248 22012 7254 22024
rect 13541 22015 13599 22021
rect 7248 21984 9996 22012
rect 7248 21972 7254 21984
rect 1854 21904 1860 21956
rect 1912 21944 1918 21956
rect 2961 21947 3019 21953
rect 2961 21944 2973 21947
rect 1912 21916 2973 21944
rect 1912 21904 1918 21916
rect 2961 21913 2973 21916
rect 3007 21913 3019 21947
rect 9968 21944 9996 21984
rect 13541 21981 13553 22015
rect 13587 21981 13599 22015
rect 13541 21975 13599 21981
rect 12158 21944 12164 21956
rect 9968 21916 12164 21944
rect 2961 21907 3019 21913
rect 12158 21904 12164 21916
rect 12216 21904 12222 21956
rect 13556 21944 13584 21975
rect 13722 21972 13728 22024
rect 13780 22012 13786 22024
rect 15304 22012 15332 22043
rect 13780 21984 15332 22012
rect 16117 22015 16175 22021
rect 13780 21972 13786 21984
rect 16117 21981 16129 22015
rect 16163 22012 16175 22015
rect 16408 22012 16436 22120
rect 17862 22108 17868 22120
rect 17920 22108 17926 22160
rect 18690 22108 18696 22160
rect 18748 22148 18754 22160
rect 18748 22120 20116 22148
rect 18748 22108 18754 22120
rect 16485 22083 16543 22089
rect 16485 22049 16497 22083
rect 16531 22049 16543 22083
rect 16485 22043 16543 22049
rect 16669 22083 16727 22089
rect 16669 22049 16681 22083
rect 16715 22080 16727 22083
rect 16758 22080 16764 22092
rect 16715 22052 16764 22080
rect 16715 22049 16727 22052
rect 16669 22043 16727 22049
rect 16163 21984 16436 22012
rect 16163 21981 16175 21984
rect 16117 21975 16175 21981
rect 16500 21956 16528 22043
rect 16758 22040 16764 22052
rect 16816 22040 16822 22092
rect 16942 22080 16948 22092
rect 16903 22052 16948 22080
rect 16942 22040 16948 22052
rect 17000 22040 17006 22092
rect 17037 22083 17095 22089
rect 17037 22049 17049 22083
rect 17083 22080 17095 22083
rect 17218 22080 17224 22092
rect 17083 22052 17224 22080
rect 17083 22049 17095 22052
rect 17037 22043 17095 22049
rect 16574 21972 16580 22024
rect 16632 22012 16638 22024
rect 17052 22012 17080 22043
rect 17218 22040 17224 22052
rect 17276 22040 17282 22092
rect 17586 22040 17592 22092
rect 17644 22080 17650 22092
rect 18141 22083 18199 22089
rect 18141 22080 18153 22083
rect 17644 22052 18153 22080
rect 17644 22040 17650 22052
rect 18141 22049 18153 22052
rect 18187 22049 18199 22083
rect 18141 22043 18199 22049
rect 18785 22083 18843 22089
rect 18785 22049 18797 22083
rect 18831 22049 18843 22083
rect 18785 22043 18843 22049
rect 19153 22083 19211 22089
rect 19153 22049 19165 22083
rect 19199 22049 19211 22083
rect 19153 22043 19211 22049
rect 17402 22012 17408 22024
rect 16632 21984 17080 22012
rect 17363 21984 17408 22012
rect 16632 21972 16638 21984
rect 17402 21972 17408 21984
rect 17460 21972 17466 22024
rect 18800 22012 18828 22043
rect 18966 22012 18972 22024
rect 18800 21984 18972 22012
rect 18966 21972 18972 21984
rect 19024 21972 19030 22024
rect 19168 22012 19196 22043
rect 19334 22040 19340 22092
rect 19392 22080 19398 22092
rect 19613 22083 19671 22089
rect 19613 22080 19625 22083
rect 19392 22052 19625 22080
rect 19392 22040 19398 22052
rect 19613 22049 19625 22052
rect 19659 22080 19671 22083
rect 19886 22080 19892 22092
rect 19659 22052 19892 22080
rect 19659 22049 19671 22052
rect 19613 22043 19671 22049
rect 19886 22040 19892 22052
rect 19944 22040 19950 22092
rect 20088 22089 20116 22120
rect 26786 22108 26792 22160
rect 26844 22148 26850 22160
rect 26844 22120 27292 22148
rect 26844 22108 26850 22120
rect 20073 22083 20131 22089
rect 20073 22049 20085 22083
rect 20119 22049 20131 22083
rect 20073 22043 20131 22049
rect 20901 22083 20959 22089
rect 20901 22049 20913 22083
rect 20947 22080 20959 22083
rect 22557 22083 22615 22089
rect 20947 22052 21404 22080
rect 20947 22049 20959 22052
rect 20901 22043 20959 22049
rect 21376 22024 21404 22052
rect 22557 22049 22569 22083
rect 22603 22080 22615 22083
rect 22646 22080 22652 22092
rect 22603 22052 22652 22080
rect 22603 22049 22615 22052
rect 22557 22043 22615 22049
rect 22646 22040 22652 22052
rect 22704 22040 22710 22092
rect 23658 22080 23664 22092
rect 23619 22052 23664 22080
rect 23658 22040 23664 22052
rect 23716 22040 23722 22092
rect 24302 22080 24308 22092
rect 24263 22052 24308 22080
rect 24302 22040 24308 22052
rect 24360 22040 24366 22092
rect 25498 22080 25504 22092
rect 25459 22052 25504 22080
rect 25498 22040 25504 22052
rect 25556 22040 25562 22092
rect 25682 22080 25688 22092
rect 25643 22052 25688 22080
rect 25682 22040 25688 22052
rect 25740 22040 25746 22092
rect 26970 22080 26976 22092
rect 26931 22052 26976 22080
rect 26970 22040 26976 22052
rect 27028 22040 27034 22092
rect 27062 22040 27068 22092
rect 27120 22080 27126 22092
rect 27157 22083 27215 22089
rect 27157 22080 27169 22083
rect 27120 22052 27169 22080
rect 27120 22040 27126 22052
rect 27157 22049 27169 22052
rect 27203 22049 27215 22083
rect 27264 22080 27292 22120
rect 27614 22108 27620 22160
rect 27672 22148 27678 22160
rect 32214 22148 32220 22160
rect 27672 22120 28120 22148
rect 27672 22108 27678 22120
rect 27706 22080 27712 22092
rect 27264 22052 27712 22080
rect 27157 22043 27215 22049
rect 27706 22040 27712 22052
rect 27764 22040 27770 22092
rect 28092 22089 28120 22120
rect 31036 22120 32220 22148
rect 28077 22083 28135 22089
rect 28077 22049 28089 22083
rect 28123 22080 28135 22083
rect 28166 22080 28172 22092
rect 28123 22052 28172 22080
rect 28123 22049 28135 22052
rect 28077 22043 28135 22049
rect 28166 22040 28172 22052
rect 28224 22040 28230 22092
rect 29086 22080 29092 22092
rect 29047 22052 29092 22080
rect 29086 22040 29092 22052
rect 29144 22040 29150 22092
rect 29546 22040 29552 22092
rect 29604 22080 29610 22092
rect 29733 22083 29791 22089
rect 29733 22080 29745 22083
rect 29604 22052 29745 22080
rect 29604 22040 29610 22052
rect 29733 22049 29745 22052
rect 29779 22049 29791 22083
rect 29733 22043 29791 22049
rect 29917 22083 29975 22089
rect 29917 22049 29929 22083
rect 29963 22080 29975 22083
rect 30282 22080 30288 22092
rect 29963 22052 30288 22080
rect 29963 22049 29975 22052
rect 29917 22043 29975 22049
rect 21174 22012 21180 22024
rect 19168 21984 20300 22012
rect 21135 21984 21180 22012
rect 15286 21944 15292 21956
rect 13556 21916 15292 21944
rect 15286 21904 15292 21916
rect 15344 21904 15350 21956
rect 16482 21944 16488 21956
rect 16395 21916 16488 21944
rect 16482 21904 16488 21916
rect 16540 21944 16546 21956
rect 19168 21944 19196 21984
rect 20272 21953 20300 21984
rect 21174 21972 21180 21984
rect 21232 21972 21238 22024
rect 21358 21972 21364 22024
rect 21416 21972 21422 22024
rect 24118 21972 24124 22024
rect 24176 22012 24182 22024
rect 24397 22015 24455 22021
rect 24397 22012 24409 22015
rect 24176 21984 24409 22012
rect 24176 21972 24182 21984
rect 24397 21981 24409 21984
rect 24443 21981 24455 22015
rect 29748 22012 29776 22043
rect 30282 22040 30288 22052
rect 30340 22040 30346 22092
rect 30653 22083 30711 22089
rect 30653 22049 30665 22083
rect 30699 22080 30711 22083
rect 30834 22080 30840 22092
rect 30699 22052 30840 22080
rect 30699 22049 30711 22052
rect 30653 22043 30711 22049
rect 30834 22040 30840 22052
rect 30892 22040 30898 22092
rect 31036 22089 31064 22120
rect 32214 22108 32220 22120
rect 32272 22108 32278 22160
rect 33686 22108 33692 22160
rect 33744 22148 33750 22160
rect 34422 22148 34428 22160
rect 33744 22120 34428 22148
rect 33744 22108 33750 22120
rect 34422 22108 34428 22120
rect 34480 22108 34486 22160
rect 31021 22083 31079 22089
rect 31021 22049 31033 22083
rect 31067 22049 31079 22083
rect 31386 22080 31392 22092
rect 31347 22052 31392 22080
rect 31021 22043 31079 22049
rect 31386 22040 31392 22052
rect 31444 22040 31450 22092
rect 32122 22040 32128 22092
rect 32180 22080 32186 22092
rect 32309 22083 32367 22089
rect 32309 22080 32321 22083
rect 32180 22052 32321 22080
rect 32180 22040 32186 22052
rect 32309 22049 32321 22052
rect 32355 22080 32367 22083
rect 32766 22080 32772 22092
rect 32355 22052 32772 22080
rect 32355 22049 32367 22052
rect 32309 22043 32367 22049
rect 32766 22040 32772 22052
rect 32824 22040 32830 22092
rect 33045 22083 33103 22089
rect 33045 22049 33057 22083
rect 33091 22049 33103 22083
rect 33045 22043 33103 22049
rect 33060 22012 33088 22043
rect 33502 22040 33508 22092
rect 33560 22080 33566 22092
rect 33873 22083 33931 22089
rect 33873 22080 33885 22083
rect 33560 22052 33885 22080
rect 33560 22040 33566 22052
rect 33873 22049 33885 22052
rect 33919 22049 33931 22083
rect 36814 22080 36820 22092
rect 33873 22043 33931 22049
rect 33980 22052 36820 22080
rect 33778 22012 33784 22024
rect 29748 21984 30052 22012
rect 33060 21984 33640 22012
rect 33739 21984 33784 22012
rect 24397 21975 24455 21981
rect 16540 21916 19196 21944
rect 20257 21947 20315 21953
rect 16540 21904 16546 21916
rect 20257 21913 20269 21947
rect 20303 21913 20315 21947
rect 23842 21944 23848 21956
rect 23803 21916 23848 21944
rect 20257 21907 20315 21913
rect 23842 21904 23848 21916
rect 23900 21904 23906 21956
rect 3326 21876 3332 21888
rect 1412 21848 3332 21876
rect 3326 21836 3332 21848
rect 3384 21836 3390 21888
rect 19334 21876 19340 21888
rect 19295 21848 19340 21876
rect 19334 21836 19340 21848
rect 19392 21836 19398 21888
rect 20162 21836 20168 21888
rect 20220 21876 20226 21888
rect 20530 21876 20536 21888
rect 20220 21848 20536 21876
rect 20220 21836 20226 21848
rect 20530 21836 20536 21848
rect 20588 21836 20594 21888
rect 23658 21836 23664 21888
rect 23716 21876 23722 21888
rect 29178 21876 29184 21888
rect 23716 21848 29184 21876
rect 23716 21836 23722 21848
rect 29178 21836 29184 21848
rect 29236 21836 29242 21888
rect 30024 21876 30052 21984
rect 33612 21956 33640 21984
rect 33778 21972 33784 21984
rect 33836 21972 33842 22024
rect 31389 21947 31447 21953
rect 31389 21913 31401 21947
rect 31435 21944 31447 21947
rect 31478 21944 31484 21956
rect 31435 21916 31484 21944
rect 31435 21913 31447 21916
rect 31389 21907 31447 21913
rect 31478 21904 31484 21916
rect 31536 21904 31542 21956
rect 33594 21904 33600 21956
rect 33652 21944 33658 21956
rect 33980 21944 34008 22052
rect 36814 22040 36820 22052
rect 36872 22040 36878 22092
rect 37366 22040 37372 22092
rect 37424 22080 37430 22092
rect 37737 22083 37795 22089
rect 37737 22080 37749 22083
rect 37424 22052 37749 22080
rect 37424 22040 37430 22052
rect 37737 22049 37749 22052
rect 37783 22049 37795 22083
rect 37737 22043 37795 22049
rect 38102 22040 38108 22092
rect 38160 22080 38166 22092
rect 38565 22083 38623 22089
rect 38565 22080 38577 22083
rect 38160 22052 38577 22080
rect 38160 22040 38166 22052
rect 38565 22049 38577 22052
rect 38611 22049 38623 22083
rect 38565 22043 38623 22049
rect 34422 21972 34428 22024
rect 34480 22012 34486 22024
rect 35161 22015 35219 22021
rect 35161 22012 35173 22015
rect 34480 21984 35173 22012
rect 34480 21972 34486 21984
rect 35161 21981 35173 21984
rect 35207 21981 35219 22015
rect 35434 22012 35440 22024
rect 35395 21984 35440 22012
rect 35161 21975 35219 21981
rect 35434 21972 35440 21984
rect 35492 21972 35498 22024
rect 38470 22012 38476 22024
rect 38431 21984 38476 22012
rect 38470 21972 38476 21984
rect 38528 21972 38534 22024
rect 33652 21916 34008 21944
rect 33652 21904 33658 21916
rect 31754 21876 31760 21888
rect 30024 21848 31760 21876
rect 31754 21836 31760 21848
rect 31812 21876 31818 21888
rect 32493 21879 32551 21885
rect 32493 21876 32505 21879
rect 31812 21848 32505 21876
rect 31812 21836 31818 21848
rect 32493 21845 32505 21848
rect 32539 21845 32551 21879
rect 32493 21839 32551 21845
rect 1104 21786 39836 21808
rect 1104 21734 4246 21786
rect 4298 21734 4310 21786
rect 4362 21734 4374 21786
rect 4426 21734 4438 21786
rect 4490 21734 34966 21786
rect 35018 21734 35030 21786
rect 35082 21734 35094 21786
rect 35146 21734 35158 21786
rect 35210 21734 39836 21786
rect 1104 21712 39836 21734
rect 2961 21675 3019 21681
rect 2961 21641 2973 21675
rect 3007 21672 3019 21675
rect 3326 21672 3332 21684
rect 3007 21644 3332 21672
rect 3007 21641 3019 21644
rect 2961 21635 3019 21641
rect 3326 21632 3332 21644
rect 3384 21632 3390 21684
rect 16942 21672 16948 21684
rect 12912 21644 16948 21672
rect 5534 21564 5540 21616
rect 5592 21604 5598 21616
rect 6089 21607 6147 21613
rect 6089 21604 6101 21607
rect 5592 21576 6101 21604
rect 5592 21564 5598 21576
rect 6089 21573 6101 21576
rect 6135 21573 6147 21607
rect 6914 21604 6920 21616
rect 6875 21576 6920 21604
rect 6089 21567 6147 21573
rect 1762 21496 1768 21548
rect 1820 21536 1826 21548
rect 3970 21536 3976 21548
rect 1820 21508 3976 21536
rect 1820 21496 1826 21508
rect 3970 21496 3976 21508
rect 4028 21496 4034 21548
rect 4890 21496 4896 21548
rect 4948 21536 4954 21548
rect 5353 21539 5411 21545
rect 5353 21536 5365 21539
rect 4948 21508 5365 21536
rect 4948 21496 4954 21508
rect 5353 21505 5365 21508
rect 5399 21505 5411 21539
rect 6104 21536 6132 21567
rect 6914 21564 6920 21576
rect 6972 21564 6978 21616
rect 7653 21539 7711 21545
rect 7653 21536 7665 21539
rect 6104 21508 7665 21536
rect 5353 21499 5411 21505
rect 7653 21505 7665 21508
rect 7699 21505 7711 21539
rect 7653 21499 7711 21505
rect 1397 21471 1455 21477
rect 1397 21437 1409 21471
rect 1443 21468 1455 21471
rect 1486 21468 1492 21480
rect 1443 21440 1492 21468
rect 1443 21437 1455 21440
rect 1397 21431 1455 21437
rect 1486 21428 1492 21440
rect 1544 21428 1550 21480
rect 1673 21471 1731 21477
rect 1673 21437 1685 21471
rect 1719 21468 1731 21471
rect 1946 21468 1952 21480
rect 1719 21440 1952 21468
rect 1719 21437 1731 21440
rect 1673 21431 1731 21437
rect 1946 21428 1952 21440
rect 2004 21428 2010 21480
rect 4062 21468 4068 21480
rect 4023 21440 4068 21468
rect 4062 21428 4068 21440
rect 4120 21428 4126 21480
rect 4341 21471 4399 21477
rect 4341 21437 4353 21471
rect 4387 21437 4399 21471
rect 4982 21468 4988 21480
rect 4943 21440 4988 21468
rect 4341 21431 4399 21437
rect 2958 21360 2964 21412
rect 3016 21400 3022 21412
rect 4356 21400 4384 21431
rect 4982 21428 4988 21440
rect 5040 21428 5046 21480
rect 5261 21471 5319 21477
rect 5261 21437 5273 21471
rect 5307 21437 5319 21471
rect 5368 21468 5396 21499
rect 10778 21496 10784 21548
rect 10836 21536 10842 21548
rect 12526 21536 12532 21548
rect 10836 21508 12532 21536
rect 10836 21496 10842 21508
rect 5905 21471 5963 21477
rect 5905 21468 5917 21471
rect 5368 21440 5917 21468
rect 5261 21431 5319 21437
rect 5905 21437 5917 21440
rect 5951 21437 5963 21471
rect 5905 21431 5963 21437
rect 3016 21372 4384 21400
rect 5276 21400 5304 21431
rect 6730 21428 6736 21480
rect 6788 21468 6794 21480
rect 6825 21471 6883 21477
rect 6825 21468 6837 21471
rect 6788 21440 6837 21468
rect 6788 21428 6794 21440
rect 6825 21437 6837 21440
rect 6871 21437 6883 21471
rect 7466 21468 7472 21480
rect 7427 21440 7472 21468
rect 6825 21431 6883 21437
rect 7466 21428 7472 21440
rect 7524 21428 7530 21480
rect 10686 21468 10692 21480
rect 10647 21440 10692 21468
rect 10686 21428 10692 21440
rect 10744 21428 10750 21480
rect 11072 21477 11100 21508
rect 12526 21496 12532 21508
rect 12584 21496 12590 21548
rect 11057 21471 11115 21477
rect 11057 21437 11069 21471
rect 11103 21437 11115 21471
rect 11057 21431 11115 21437
rect 11425 21471 11483 21477
rect 11425 21437 11437 21471
rect 11471 21468 11483 21471
rect 12434 21468 12440 21480
rect 11471 21440 12440 21468
rect 11471 21437 11483 21440
rect 11425 21431 11483 21437
rect 12434 21428 12440 21440
rect 12492 21428 12498 21480
rect 12710 21428 12716 21480
rect 12768 21468 12774 21480
rect 12805 21471 12863 21477
rect 12805 21468 12817 21471
rect 12768 21440 12817 21468
rect 12768 21428 12774 21440
rect 12805 21437 12817 21440
rect 12851 21468 12863 21471
rect 12912 21468 12940 21644
rect 16942 21632 16948 21644
rect 17000 21632 17006 21684
rect 18138 21672 18144 21684
rect 18099 21644 18144 21672
rect 18138 21632 18144 21644
rect 18196 21632 18202 21684
rect 25225 21675 25283 21681
rect 23308 21644 24624 21672
rect 20346 21564 20352 21616
rect 20404 21604 20410 21616
rect 20404 21576 21220 21604
rect 20404 21564 20410 21576
rect 13722 21536 13728 21548
rect 13683 21508 13728 21536
rect 13722 21496 13728 21508
rect 13780 21496 13786 21548
rect 13814 21496 13820 21548
rect 13872 21536 13878 21548
rect 14185 21539 14243 21545
rect 14185 21536 14197 21539
rect 13872 21508 14197 21536
rect 13872 21496 13878 21508
rect 14185 21505 14197 21508
rect 14231 21505 14243 21539
rect 14185 21499 14243 21505
rect 17037 21539 17095 21545
rect 17037 21505 17049 21539
rect 17083 21536 17095 21539
rect 21192 21536 21220 21576
rect 21450 21564 21456 21616
rect 21508 21604 21514 21616
rect 22554 21604 22560 21616
rect 21508 21576 22560 21604
rect 21508 21564 21514 21576
rect 22554 21564 22560 21576
rect 22612 21564 22618 21616
rect 17083 21508 21128 21536
rect 21192 21508 21680 21536
rect 17083 21505 17095 21508
rect 17037 21499 17095 21505
rect 13170 21468 13176 21480
rect 12851 21440 12940 21468
rect 13131 21440 13176 21468
rect 12851 21437 12863 21440
rect 12805 21431 12863 21437
rect 13170 21428 13176 21440
rect 13228 21428 13234 21480
rect 13541 21471 13599 21477
rect 13541 21437 13553 21471
rect 13587 21437 13599 21471
rect 14458 21468 14464 21480
rect 14419 21440 14464 21468
rect 13541 21431 13599 21437
rect 5534 21400 5540 21412
rect 5276 21372 5540 21400
rect 3016 21360 3022 21372
rect 5534 21360 5540 21372
rect 5592 21360 5598 21412
rect 11609 21403 11667 21409
rect 11609 21369 11621 21403
rect 11655 21400 11667 21403
rect 11698 21400 11704 21412
rect 11655 21372 11704 21400
rect 11655 21369 11667 21372
rect 11609 21363 11667 21369
rect 11698 21360 11704 21372
rect 11756 21360 11762 21412
rect 13556 21400 13584 21431
rect 14458 21428 14464 21440
rect 14516 21428 14522 21480
rect 16574 21468 16580 21480
rect 16535 21440 16580 21468
rect 16574 21428 16580 21440
rect 16632 21428 16638 21480
rect 16761 21471 16819 21477
rect 16761 21437 16773 21471
rect 16807 21437 16819 21471
rect 16761 21431 16819 21437
rect 13722 21400 13728 21412
rect 13556 21372 13728 21400
rect 13722 21360 13728 21372
rect 13780 21360 13786 21412
rect 15841 21403 15899 21409
rect 15841 21369 15853 21403
rect 15887 21400 15899 21403
rect 16114 21400 16120 21412
rect 15887 21372 16120 21400
rect 15887 21369 15899 21372
rect 15841 21363 15899 21369
rect 16114 21360 16120 21372
rect 16172 21360 16178 21412
rect 16482 21360 16488 21412
rect 16540 21400 16546 21412
rect 16776 21400 16804 21431
rect 17126 21428 17132 21480
rect 17184 21468 17190 21480
rect 18049 21471 18107 21477
rect 18049 21468 18061 21471
rect 17184 21440 18061 21468
rect 17184 21428 17190 21440
rect 18049 21437 18061 21440
rect 18095 21437 18107 21471
rect 18049 21431 18107 21437
rect 18877 21471 18935 21477
rect 18877 21437 18889 21471
rect 18923 21437 18935 21471
rect 19150 21468 19156 21480
rect 19111 21440 19156 21468
rect 18877 21431 18935 21437
rect 16540 21372 16804 21400
rect 16540 21360 16546 21372
rect 13078 21292 13084 21344
rect 13136 21332 13142 21344
rect 18892 21332 18920 21431
rect 19150 21428 19156 21440
rect 19208 21428 19214 21480
rect 20898 21360 20904 21412
rect 20956 21400 20962 21412
rect 20993 21403 21051 21409
rect 20993 21400 21005 21403
rect 20956 21372 21005 21400
rect 20956 21360 20962 21372
rect 20993 21369 21005 21372
rect 21039 21369 21051 21403
rect 21100 21400 21128 21508
rect 21450 21468 21456 21480
rect 21411 21440 21456 21468
rect 21450 21428 21456 21440
rect 21508 21428 21514 21480
rect 21652 21477 21680 21508
rect 21744 21508 23244 21536
rect 21637 21471 21695 21477
rect 21637 21437 21649 21471
rect 21683 21437 21695 21471
rect 21637 21431 21695 21437
rect 21744 21400 21772 21508
rect 21821 21471 21879 21477
rect 21821 21437 21833 21471
rect 21867 21468 21879 21471
rect 21867 21440 22508 21468
rect 21867 21437 21879 21440
rect 21821 21431 21879 21437
rect 21100 21372 21772 21400
rect 20993 21363 21051 21369
rect 21910 21360 21916 21412
rect 21968 21400 21974 21412
rect 22097 21403 22155 21409
rect 22097 21400 22109 21403
rect 21968 21372 22109 21400
rect 21968 21360 21974 21372
rect 22097 21369 22109 21372
rect 22143 21369 22155 21403
rect 22480 21400 22508 21440
rect 22554 21428 22560 21480
rect 22612 21468 22618 21480
rect 22741 21471 22799 21477
rect 22612 21440 22657 21468
rect 22612 21428 22618 21440
rect 22741 21437 22753 21471
rect 22787 21468 22799 21471
rect 22830 21468 22836 21480
rect 22787 21440 22836 21468
rect 22787 21437 22799 21440
rect 22741 21431 22799 21437
rect 22830 21428 22836 21440
rect 22888 21428 22894 21480
rect 23216 21477 23244 21508
rect 22925 21471 22983 21477
rect 22925 21437 22937 21471
rect 22971 21437 22983 21471
rect 22925 21431 22983 21437
rect 23201 21471 23259 21477
rect 23201 21437 23213 21471
rect 23247 21437 23259 21471
rect 23201 21431 23259 21437
rect 22940 21400 22968 21431
rect 23308 21400 23336 21644
rect 24596 21604 24624 21644
rect 25225 21641 25237 21675
rect 25271 21672 25283 21675
rect 25682 21672 25688 21684
rect 25271 21644 25688 21672
rect 25271 21641 25283 21644
rect 25225 21635 25283 21641
rect 25682 21632 25688 21644
rect 25740 21632 25746 21684
rect 25774 21632 25780 21684
rect 25832 21672 25838 21684
rect 34146 21672 34152 21684
rect 25832 21644 34152 21672
rect 25832 21632 25838 21644
rect 34146 21632 34152 21644
rect 34204 21632 34210 21684
rect 36170 21672 36176 21684
rect 34992 21644 36176 21672
rect 26786 21604 26792 21616
rect 24596 21576 26792 21604
rect 26786 21564 26792 21576
rect 26844 21564 26850 21616
rect 31481 21607 31539 21613
rect 31481 21573 31493 21607
rect 31527 21573 31539 21607
rect 31481 21567 31539 21573
rect 33597 21607 33655 21613
rect 33597 21573 33609 21607
rect 33643 21604 33655 21607
rect 34330 21604 34336 21616
rect 33643 21576 34336 21604
rect 33643 21573 33655 21576
rect 33597 21567 33655 21573
rect 23474 21496 23480 21548
rect 23532 21536 23538 21548
rect 23661 21539 23719 21545
rect 23661 21536 23673 21539
rect 23532 21508 23673 21536
rect 23532 21496 23538 21508
rect 23661 21505 23673 21508
rect 23707 21505 23719 21539
rect 23661 21499 23719 21505
rect 23676 21468 23704 21499
rect 23842 21496 23848 21548
rect 23900 21536 23906 21548
rect 23937 21539 23995 21545
rect 23937 21536 23949 21539
rect 23900 21508 23949 21536
rect 23900 21496 23906 21508
rect 23937 21505 23949 21508
rect 23983 21505 23995 21539
rect 28994 21536 29000 21548
rect 23937 21499 23995 21505
rect 26436 21508 29000 21536
rect 26142 21468 26148 21480
rect 23676 21440 26004 21468
rect 26103 21440 26148 21468
rect 22480 21372 23336 21400
rect 25976 21400 26004 21440
rect 26142 21428 26148 21440
rect 26200 21428 26206 21480
rect 26436 21412 26464 21508
rect 28994 21496 29000 21508
rect 29052 21536 29058 21548
rect 29273 21539 29331 21545
rect 29273 21536 29285 21539
rect 29052 21508 29285 21536
rect 29052 21496 29058 21508
rect 29273 21505 29285 21508
rect 29319 21505 29331 21539
rect 29273 21499 29331 21505
rect 29549 21539 29607 21545
rect 29549 21505 29561 21539
rect 29595 21536 29607 21539
rect 31496 21536 31524 21567
rect 34330 21564 34336 21576
rect 34388 21604 34394 21616
rect 34388 21576 34928 21604
rect 34388 21564 34394 21576
rect 32306 21536 32312 21548
rect 29595 21508 31524 21536
rect 32267 21508 32312 21536
rect 29595 21505 29607 21508
rect 29549 21499 29607 21505
rect 32306 21496 32312 21508
rect 32364 21496 32370 21548
rect 32950 21496 32956 21548
rect 33008 21536 33014 21548
rect 33962 21536 33968 21548
rect 33008 21508 33968 21536
rect 33008 21496 33014 21508
rect 26789 21471 26847 21477
rect 26789 21437 26801 21471
rect 26835 21437 26847 21471
rect 26970 21468 26976 21480
rect 26931 21440 26976 21468
rect 26789 21431 26847 21437
rect 26418 21400 26424 21412
rect 25976 21372 26424 21400
rect 22097 21363 22155 21369
rect 26418 21360 26424 21372
rect 26476 21360 26482 21412
rect 26804 21400 26832 21431
rect 26970 21428 26976 21440
rect 27028 21428 27034 21480
rect 27706 21468 27712 21480
rect 27667 21440 27712 21468
rect 27706 21428 27712 21440
rect 27764 21428 27770 21480
rect 28166 21468 28172 21480
rect 28127 21440 28172 21468
rect 28166 21428 28172 21440
rect 28224 21428 28230 21480
rect 29178 21428 29184 21480
rect 29236 21468 29242 21480
rect 31389 21471 31447 21477
rect 31389 21468 31401 21471
rect 29236 21440 31401 21468
rect 29236 21428 29242 21440
rect 31389 21437 31401 21440
rect 31435 21437 31447 21471
rect 31389 21431 31447 21437
rect 27982 21400 27988 21412
rect 26804 21372 27988 21400
rect 27982 21360 27988 21372
rect 28040 21360 28046 21412
rect 31404 21400 31432 21431
rect 31478 21428 31484 21480
rect 31536 21468 31542 21480
rect 31941 21471 31999 21477
rect 31941 21468 31953 21471
rect 31536 21440 31953 21468
rect 31536 21428 31542 21440
rect 31941 21437 31953 21440
rect 31987 21437 31999 21471
rect 33226 21468 33232 21480
rect 33187 21440 33232 21468
rect 31941 21431 31999 21437
rect 33226 21428 33232 21440
rect 33284 21428 33290 21480
rect 33796 21477 33824 21508
rect 33962 21496 33968 21508
rect 34020 21496 34026 21548
rect 33781 21471 33839 21477
rect 33781 21437 33793 21471
rect 33827 21437 33839 21471
rect 34146 21468 34152 21480
rect 34107 21440 34152 21468
rect 33781 21431 33839 21437
rect 34146 21428 34152 21440
rect 34204 21428 34210 21480
rect 34900 21477 34928 21576
rect 34241 21471 34299 21477
rect 34241 21437 34253 21471
rect 34287 21437 34299 21471
rect 34241 21431 34299 21437
rect 34885 21471 34943 21477
rect 34885 21437 34897 21471
rect 34931 21437 34943 21471
rect 34885 21431 34943 21437
rect 34256 21400 34284 21431
rect 34992 21400 35020 21644
rect 36170 21632 36176 21644
rect 36228 21672 36234 21684
rect 38841 21675 38899 21681
rect 38841 21672 38853 21675
rect 36228 21644 38853 21672
rect 36228 21632 36234 21644
rect 38841 21641 38853 21644
rect 38887 21641 38899 21675
rect 38841 21635 38899 21641
rect 35618 21564 35624 21616
rect 35676 21604 35682 21616
rect 35802 21604 35808 21616
rect 35676 21576 35808 21604
rect 35676 21564 35682 21576
rect 35802 21564 35808 21576
rect 35860 21564 35866 21616
rect 35434 21536 35440 21548
rect 35395 21508 35440 21536
rect 35434 21496 35440 21508
rect 35492 21496 35498 21548
rect 36446 21496 36452 21548
rect 36504 21536 36510 21548
rect 37461 21539 37519 21545
rect 37461 21536 37473 21539
rect 36504 21508 37473 21536
rect 36504 21496 36510 21508
rect 37461 21505 37473 21508
rect 37507 21505 37519 21539
rect 37461 21499 37519 21505
rect 37737 21539 37795 21545
rect 37737 21505 37749 21539
rect 37783 21536 37795 21539
rect 37826 21536 37832 21548
rect 37783 21508 37832 21536
rect 37783 21505 37795 21508
rect 37737 21499 37795 21505
rect 37826 21496 37832 21508
rect 37884 21496 37890 21548
rect 35529 21471 35587 21477
rect 35529 21437 35541 21471
rect 35575 21437 35587 21471
rect 35802 21468 35808 21480
rect 35763 21440 35808 21468
rect 35529 21431 35587 21437
rect 31404 21372 34100 21400
rect 34256 21372 35020 21400
rect 34072 21344 34100 21372
rect 13136 21304 18920 21332
rect 20441 21335 20499 21341
rect 13136 21292 13142 21304
rect 20441 21301 20453 21335
rect 20487 21332 20499 21335
rect 22554 21332 22560 21344
rect 20487 21304 22560 21332
rect 20487 21301 20499 21304
rect 20441 21295 20499 21301
rect 22554 21292 22560 21304
rect 22612 21292 22618 21344
rect 23290 21332 23296 21344
rect 23251 21304 23296 21332
rect 23290 21292 23296 21304
rect 23348 21292 23354 21344
rect 23382 21292 23388 21344
rect 23440 21332 23446 21344
rect 25774 21332 25780 21344
rect 23440 21304 25780 21332
rect 23440 21292 23446 21304
rect 25774 21292 25780 21304
rect 25832 21292 25838 21344
rect 26234 21332 26240 21344
rect 26195 21304 26240 21332
rect 26234 21292 26240 21304
rect 26292 21292 26298 21344
rect 27614 21292 27620 21344
rect 27672 21332 27678 21344
rect 27801 21335 27859 21341
rect 27801 21332 27813 21335
rect 27672 21304 27813 21332
rect 27672 21292 27678 21304
rect 27801 21301 27813 21304
rect 27847 21301 27859 21335
rect 27801 21295 27859 21301
rect 29362 21292 29368 21344
rect 29420 21332 29426 21344
rect 30006 21332 30012 21344
rect 29420 21304 30012 21332
rect 29420 21292 29426 21304
rect 30006 21292 30012 21304
rect 30064 21332 30070 21344
rect 30653 21335 30711 21341
rect 30653 21332 30665 21335
rect 30064 21304 30665 21332
rect 30064 21292 30070 21304
rect 30653 21301 30665 21304
rect 30699 21301 30711 21335
rect 30653 21295 30711 21301
rect 31846 21292 31852 21344
rect 31904 21332 31910 21344
rect 33042 21332 33048 21344
rect 31904 21304 33048 21332
rect 31904 21292 31910 21304
rect 33042 21292 33048 21304
rect 33100 21292 33106 21344
rect 34054 21292 34060 21344
rect 34112 21292 34118 21344
rect 35544 21332 35572 21431
rect 35802 21428 35808 21440
rect 35860 21428 35866 21480
rect 35986 21428 35992 21480
rect 36044 21468 36050 21480
rect 36081 21471 36139 21477
rect 36081 21468 36093 21471
rect 36044 21440 36093 21468
rect 36044 21428 36050 21440
rect 36081 21437 36093 21440
rect 36127 21468 36139 21471
rect 36262 21468 36268 21480
rect 36127 21440 36268 21468
rect 36127 21437 36139 21440
rect 36081 21431 36139 21437
rect 36262 21428 36268 21440
rect 36320 21428 36326 21480
rect 36538 21428 36544 21480
rect 36596 21468 36602 21480
rect 36817 21471 36875 21477
rect 36817 21468 36829 21471
rect 36596 21440 36829 21468
rect 36596 21428 36602 21440
rect 36817 21437 36829 21440
rect 36863 21468 36875 21471
rect 36906 21468 36912 21480
rect 36863 21440 36912 21468
rect 36863 21437 36875 21440
rect 36817 21431 36875 21437
rect 36906 21428 36912 21440
rect 36964 21428 36970 21480
rect 39022 21400 39028 21412
rect 38672 21372 39028 21400
rect 38672 21344 38700 21372
rect 39022 21360 39028 21372
rect 39080 21360 39086 21412
rect 38654 21332 38660 21344
rect 35544 21304 38660 21332
rect 38654 21292 38660 21304
rect 38712 21292 38718 21344
rect 1104 21242 39836 21264
rect 1104 21190 19606 21242
rect 19658 21190 19670 21242
rect 19722 21190 19734 21242
rect 19786 21190 19798 21242
rect 19850 21190 39836 21242
rect 1104 21168 39836 21190
rect 1946 21128 1952 21140
rect 1907 21100 1952 21128
rect 1946 21088 1952 21100
rect 2004 21088 2010 21140
rect 5534 21088 5540 21140
rect 5592 21128 5598 21140
rect 5902 21128 5908 21140
rect 5592 21100 5908 21128
rect 5592 21088 5598 21100
rect 5902 21088 5908 21100
rect 5960 21128 5966 21140
rect 7193 21131 7251 21137
rect 7193 21128 7205 21131
rect 5960 21100 7205 21128
rect 5960 21088 5966 21100
rect 7193 21097 7205 21100
rect 7239 21097 7251 21131
rect 9858 21128 9864 21140
rect 7193 21091 7251 21097
rect 8036 21100 9864 21128
rect 1762 21020 1768 21072
rect 1820 21060 1826 21072
rect 2498 21060 2504 21072
rect 1820 21032 2504 21060
rect 1820 21020 1826 21032
rect 2498 21020 2504 21032
rect 2556 21060 2562 21072
rect 4801 21063 4859 21069
rect 4801 21060 4813 21063
rect 2556 21032 4813 21060
rect 2556 21020 2562 21032
rect 4801 21029 4813 21032
rect 4847 21029 4859 21063
rect 4801 21023 4859 21029
rect 1854 20992 1860 21004
rect 1815 20964 1860 20992
rect 1854 20952 1860 20964
rect 1912 20952 1918 21004
rect 2958 20992 2964 21004
rect 2919 20964 2964 20992
rect 2958 20952 2964 20964
rect 3016 20952 3022 21004
rect 3326 20992 3332 21004
rect 3287 20964 3332 20992
rect 3326 20952 3332 20964
rect 3384 20952 3390 21004
rect 4893 20995 4951 21001
rect 4893 20961 4905 20995
rect 4939 20992 4951 20995
rect 5626 20992 5632 21004
rect 4939 20964 5632 20992
rect 4939 20961 4951 20964
rect 4893 20955 4951 20961
rect 5626 20952 5632 20964
rect 5684 20952 5690 21004
rect 8036 21001 8064 21100
rect 9858 21088 9864 21100
rect 9916 21088 9922 21140
rect 15378 21128 15384 21140
rect 10888 21100 13492 21128
rect 15339 21100 15384 21128
rect 8846 21020 8852 21072
rect 8904 21060 8910 21072
rect 10045 21063 10103 21069
rect 10045 21060 10057 21063
rect 8904 21032 10057 21060
rect 8904 21020 8910 21032
rect 10045 21029 10057 21032
rect 10091 21029 10103 21063
rect 10045 21023 10103 21029
rect 8021 20995 8079 21001
rect 8021 20992 8033 20995
rect 5736 20964 8033 20992
rect 1670 20884 1676 20936
rect 1728 20924 1734 20936
rect 2501 20927 2559 20933
rect 2501 20924 2513 20927
rect 1728 20896 2513 20924
rect 1728 20884 1734 20896
rect 2501 20893 2513 20896
rect 2547 20893 2559 20927
rect 2501 20887 2559 20893
rect 3421 20927 3479 20933
rect 3421 20893 3433 20927
rect 3467 20924 3479 20927
rect 4982 20924 4988 20936
rect 3467 20896 4988 20924
rect 3467 20893 3479 20896
rect 3421 20887 3479 20893
rect 4982 20884 4988 20896
rect 5040 20884 5046 20936
rect 3970 20816 3976 20868
rect 4028 20856 4034 20868
rect 5736 20856 5764 20964
rect 8021 20961 8033 20964
rect 8067 20961 8079 20995
rect 8021 20955 8079 20961
rect 8757 20995 8815 21001
rect 8757 20961 8769 20995
rect 8803 20992 8815 20995
rect 9950 20992 9956 21004
rect 8803 20964 9628 20992
rect 9911 20964 9956 20992
rect 8803 20961 8815 20964
rect 8757 20955 8815 20961
rect 5810 20884 5816 20936
rect 5868 20924 5874 20936
rect 6089 20927 6147 20933
rect 5868 20896 5913 20924
rect 5868 20884 5874 20896
rect 6089 20893 6101 20927
rect 6135 20924 6147 20927
rect 6914 20924 6920 20936
rect 6135 20896 6920 20924
rect 6135 20893 6147 20896
rect 6089 20887 6147 20893
rect 6914 20884 6920 20896
rect 6972 20884 6978 20936
rect 9033 20927 9091 20933
rect 9033 20893 9045 20927
rect 9079 20924 9091 20927
rect 9122 20924 9128 20936
rect 9079 20896 9128 20924
rect 9079 20893 9091 20896
rect 9033 20887 9091 20893
rect 9122 20884 9128 20896
rect 9180 20884 9186 20936
rect 4028 20828 5764 20856
rect 8297 20859 8355 20865
rect 4028 20816 4034 20828
rect 8297 20825 8309 20859
rect 8343 20856 8355 20859
rect 8662 20856 8668 20868
rect 8343 20828 8668 20856
rect 8343 20825 8355 20828
rect 8297 20819 8355 20825
rect 8662 20816 8668 20828
rect 8720 20816 8726 20868
rect 9600 20856 9628 20964
rect 9950 20952 9956 20964
rect 10008 20952 10014 21004
rect 10410 20992 10416 21004
rect 10371 20964 10416 20992
rect 10410 20952 10416 20964
rect 10468 20952 10474 21004
rect 10888 21001 10916 21100
rect 13170 21060 13176 21072
rect 11164 21032 13176 21060
rect 11164 21004 11192 21032
rect 13170 21020 13176 21032
rect 13228 21020 13234 21072
rect 13464 21060 13492 21100
rect 15378 21088 15384 21100
rect 15436 21088 15442 21140
rect 17586 21088 17592 21140
rect 17644 21128 17650 21140
rect 21177 21131 21235 21137
rect 17644 21100 20024 21128
rect 17644 21088 17650 21100
rect 19996 21072 20024 21100
rect 21177 21097 21189 21131
rect 21223 21128 21235 21131
rect 21634 21128 21640 21140
rect 21223 21100 21640 21128
rect 21223 21097 21235 21100
rect 21177 21091 21235 21097
rect 21634 21088 21640 21100
rect 21692 21088 21698 21140
rect 23569 21131 23627 21137
rect 23569 21097 23581 21131
rect 23615 21128 23627 21131
rect 24854 21128 24860 21140
rect 23615 21100 24860 21128
rect 23615 21097 23627 21100
rect 23569 21091 23627 21097
rect 24854 21088 24860 21100
rect 24912 21088 24918 21140
rect 26510 21088 26516 21140
rect 26568 21128 26574 21140
rect 26973 21131 27031 21137
rect 26973 21128 26985 21131
rect 26568 21100 26985 21128
rect 26568 21088 26574 21100
rect 26973 21097 26985 21100
rect 27019 21097 27031 21131
rect 26973 21091 27031 21097
rect 28258 21088 28264 21140
rect 28316 21128 28322 21140
rect 29365 21131 29423 21137
rect 29365 21128 29377 21131
rect 28316 21100 29377 21128
rect 28316 21088 28322 21100
rect 29365 21097 29377 21100
rect 29411 21097 29423 21131
rect 29365 21091 29423 21097
rect 31481 21131 31539 21137
rect 31481 21097 31493 21131
rect 31527 21128 31539 21131
rect 32214 21128 32220 21140
rect 31527 21100 32220 21128
rect 31527 21097 31539 21100
rect 31481 21091 31539 21097
rect 32214 21088 32220 21100
rect 32272 21088 32278 21140
rect 32585 21131 32643 21137
rect 32585 21097 32597 21131
rect 32631 21128 32643 21131
rect 34146 21128 34152 21140
rect 32631 21100 34152 21128
rect 32631 21097 32643 21100
rect 32585 21091 32643 21097
rect 34146 21088 34152 21100
rect 34204 21088 34210 21140
rect 35434 21088 35440 21140
rect 35492 21128 35498 21140
rect 35802 21128 35808 21140
rect 35492 21100 35808 21128
rect 35492 21088 35498 21100
rect 35802 21088 35808 21100
rect 35860 21128 35866 21140
rect 35860 21100 37780 21128
rect 35860 21088 35866 21100
rect 14182 21060 14188 21072
rect 13464 21032 14188 21060
rect 10873 20995 10931 21001
rect 10873 20961 10885 20995
rect 10919 20961 10931 20995
rect 11146 20992 11152 21004
rect 11059 20964 11152 20992
rect 10873 20955 10931 20961
rect 11146 20952 11152 20964
rect 11204 20952 11210 21004
rect 11606 20992 11612 21004
rect 11567 20964 11612 20992
rect 11606 20952 11612 20964
rect 11664 20952 11670 21004
rect 12710 20992 12716 21004
rect 12671 20964 12716 20992
rect 12710 20952 12716 20964
rect 12768 20952 12774 21004
rect 13464 21001 13492 21032
rect 14182 21020 14188 21032
rect 14240 21020 14246 21072
rect 14274 21020 14280 21072
rect 14332 21060 14338 21072
rect 16209 21063 16267 21069
rect 16209 21060 16221 21063
rect 14332 21032 16221 21060
rect 14332 21020 14338 21032
rect 16209 21029 16221 21032
rect 16255 21029 16267 21063
rect 18877 21063 18935 21069
rect 16209 21023 16267 21029
rect 17144 21032 18736 21060
rect 17144 21004 17172 21032
rect 12805 20995 12863 21001
rect 12805 20961 12817 20995
rect 12851 20961 12863 20995
rect 12805 20955 12863 20961
rect 13449 20995 13507 21001
rect 13449 20961 13461 20995
rect 13495 20961 13507 20995
rect 13722 20992 13728 21004
rect 13683 20964 13728 20992
rect 13449 20955 13507 20961
rect 12820 20924 12848 20955
rect 13722 20952 13728 20964
rect 13780 20952 13786 21004
rect 14369 20995 14427 21001
rect 14369 20961 14381 20995
rect 14415 20961 14427 20995
rect 15286 20992 15292 21004
rect 15247 20964 15292 20992
rect 14369 20955 14427 20961
rect 13078 20924 13084 20936
rect 12820 20896 13084 20924
rect 13078 20884 13084 20896
rect 13136 20924 13142 20936
rect 14384 20924 14412 20955
rect 15286 20952 15292 20964
rect 15344 20952 15350 21004
rect 16666 20992 16672 21004
rect 16627 20964 16672 20992
rect 16666 20952 16672 20964
rect 16724 20952 16730 21004
rect 16850 20992 16856 21004
rect 16811 20964 16856 20992
rect 16850 20952 16856 20964
rect 16908 20952 16914 21004
rect 17126 20992 17132 21004
rect 17039 20964 17132 20992
rect 17126 20952 17132 20964
rect 17184 20952 17190 21004
rect 17310 20992 17316 21004
rect 17271 20964 17316 20992
rect 17310 20952 17316 20964
rect 17368 20952 17374 21004
rect 17586 20992 17592 21004
rect 17547 20964 17592 20992
rect 17586 20952 17592 20964
rect 17644 20952 17650 21004
rect 18141 20995 18199 21001
rect 18141 20961 18153 20995
rect 18187 20961 18199 20995
rect 18141 20955 18199 20961
rect 18601 20995 18659 21001
rect 18601 20961 18613 20995
rect 18647 20961 18659 20995
rect 18708 20992 18736 21032
rect 18877 21029 18889 21063
rect 18923 21060 18935 21063
rect 19150 21060 19156 21072
rect 18923 21032 19156 21060
rect 18923 21029 18935 21032
rect 18877 21023 18935 21029
rect 19150 21020 19156 21032
rect 19208 21020 19214 21072
rect 19426 21020 19432 21072
rect 19484 21060 19490 21072
rect 19797 21063 19855 21069
rect 19797 21060 19809 21063
rect 19484 21032 19809 21060
rect 19484 21020 19490 21032
rect 19797 21029 19809 21032
rect 19843 21029 19855 21063
rect 19978 21060 19984 21072
rect 19939 21032 19984 21060
rect 19797 21023 19855 21029
rect 19978 21020 19984 21032
rect 20036 21020 20042 21072
rect 22830 21060 22836 21072
rect 20824 21032 22836 21060
rect 19886 20992 19892 21004
rect 18708 20964 19748 20992
rect 19847 20964 19892 20992
rect 18601 20955 18659 20961
rect 13136 20896 14412 20924
rect 13136 20884 13142 20896
rect 10410 20856 10416 20868
rect 9600 20828 10416 20856
rect 10410 20816 10416 20828
rect 10468 20816 10474 20868
rect 12158 20816 12164 20868
rect 12216 20856 12222 20868
rect 18156 20856 18184 20955
rect 18616 20924 18644 20955
rect 18874 20924 18880 20936
rect 18616 20896 18880 20924
rect 18874 20884 18880 20896
rect 18932 20884 18938 20936
rect 19613 20927 19671 20933
rect 19613 20893 19625 20927
rect 19659 20893 19671 20927
rect 19720 20924 19748 20964
rect 19886 20952 19892 20964
rect 19944 20952 19950 21004
rect 20162 20992 20168 21004
rect 19996 20964 20168 20992
rect 19996 20924 20024 20964
rect 20162 20952 20168 20964
rect 20220 20992 20226 21004
rect 20824 20992 20852 21032
rect 22830 21020 22836 21032
rect 22888 21020 22894 21072
rect 25682 21060 25688 21072
rect 23492 21032 25688 21060
rect 20220 20964 20852 20992
rect 20220 20952 20226 20964
rect 20898 20952 20904 21004
rect 20956 20992 20962 21004
rect 21085 20995 21143 21001
rect 21085 20992 21097 20995
rect 20956 20964 21097 20992
rect 20956 20952 20962 20964
rect 21085 20961 21097 20964
rect 21131 20961 21143 20995
rect 21085 20955 21143 20961
rect 21266 20952 21272 21004
rect 21324 20992 21330 21004
rect 21637 20995 21695 21001
rect 21637 20992 21649 20995
rect 21324 20964 21649 20992
rect 21324 20952 21330 20964
rect 21637 20961 21649 20964
rect 21683 20961 21695 20995
rect 22554 20992 22560 21004
rect 22515 20964 22560 20992
rect 21637 20955 21695 20961
rect 22554 20952 22560 20964
rect 22612 20952 22618 21004
rect 23109 20995 23167 21001
rect 23109 20961 23121 20995
rect 23155 20992 23167 20995
rect 23382 20992 23388 21004
rect 23155 20964 23388 20992
rect 23155 20961 23167 20964
rect 23109 20955 23167 20961
rect 23382 20952 23388 20964
rect 23440 20952 23446 21004
rect 23492 21001 23520 21032
rect 25682 21020 25688 21032
rect 25740 21020 25746 21072
rect 23477 20995 23535 21001
rect 23477 20961 23489 20995
rect 23523 20961 23535 20995
rect 23750 20992 23756 21004
rect 23711 20964 23756 20992
rect 23477 20955 23535 20961
rect 23750 20952 23756 20964
rect 23808 20952 23814 21004
rect 24118 20992 24124 21004
rect 24079 20964 24124 20992
rect 24118 20952 24124 20964
rect 24176 20952 24182 21004
rect 24489 20995 24547 21001
rect 24489 20961 24501 20995
rect 24535 20992 24547 20995
rect 24578 20992 24584 21004
rect 24535 20964 24584 20992
rect 24535 20961 24547 20964
rect 24489 20955 24547 20961
rect 24578 20952 24584 20964
rect 24636 20952 24642 21004
rect 25409 20995 25467 21001
rect 25409 20961 25421 20995
rect 25455 20992 25467 20995
rect 25590 20992 25596 21004
rect 25455 20964 25596 20992
rect 25455 20961 25467 20964
rect 25409 20955 25467 20961
rect 19720 20896 20024 20924
rect 20349 20927 20407 20933
rect 19613 20887 19671 20893
rect 20349 20893 20361 20927
rect 20395 20924 20407 20927
rect 20395 20896 21312 20924
rect 20395 20893 20407 20896
rect 20349 20887 20407 20893
rect 12216 20828 18184 20856
rect 12216 20816 12222 20828
rect 4614 20788 4620 20800
rect 4575 20760 4620 20788
rect 4614 20748 4620 20760
rect 4672 20748 4678 20800
rect 5074 20788 5080 20800
rect 5035 20760 5080 20788
rect 5074 20748 5080 20760
rect 5132 20748 5138 20800
rect 12529 20791 12587 20797
rect 12529 20757 12541 20791
rect 12575 20788 12587 20791
rect 12986 20788 12992 20800
rect 12575 20760 12992 20788
rect 12575 20757 12587 20760
rect 12529 20751 12587 20757
rect 12986 20748 12992 20760
rect 13044 20748 13050 20800
rect 13170 20748 13176 20800
rect 13228 20788 13234 20800
rect 14553 20791 14611 20797
rect 14553 20788 14565 20791
rect 13228 20760 14565 20788
rect 13228 20748 13234 20760
rect 14553 20757 14565 20760
rect 14599 20788 14611 20791
rect 19058 20788 19064 20800
rect 14599 20760 19064 20788
rect 14599 20757 14611 20760
rect 14553 20751 14611 20757
rect 19058 20748 19064 20760
rect 19116 20748 19122 20800
rect 19628 20788 19656 20887
rect 21284 20856 21312 20896
rect 21818 20884 21824 20936
rect 21876 20924 21882 20936
rect 21913 20927 21971 20933
rect 21913 20924 21925 20927
rect 21876 20896 21925 20924
rect 21876 20884 21882 20896
rect 21913 20893 21925 20896
rect 21959 20893 21971 20927
rect 21913 20887 21971 20893
rect 22370 20884 22376 20936
rect 22428 20924 22434 20936
rect 22465 20927 22523 20933
rect 22465 20924 22477 20927
rect 22428 20896 22477 20924
rect 22428 20884 22434 20896
rect 22465 20893 22477 20896
rect 22511 20893 22523 20927
rect 22465 20887 22523 20893
rect 22646 20884 22652 20936
rect 22704 20924 22710 20936
rect 25424 20924 25452 20955
rect 25590 20952 25596 20964
rect 25648 20952 25654 21004
rect 25777 20995 25835 21001
rect 25777 20961 25789 20995
rect 25823 20992 25835 20995
rect 26528 20992 26556 21088
rect 28442 21020 28448 21072
rect 28500 21060 28506 21072
rect 28902 21060 28908 21072
rect 28500 21032 28908 21060
rect 28500 21020 28506 21032
rect 28902 21020 28908 21032
rect 28960 21060 28966 21072
rect 29273 21063 29331 21069
rect 29273 21060 29285 21063
rect 28960 21032 29285 21060
rect 28960 21020 28966 21032
rect 29273 21029 29285 21032
rect 29319 21029 29331 21063
rect 29273 21023 29331 21029
rect 29457 21063 29515 21069
rect 29457 21029 29469 21063
rect 29503 21029 29515 21063
rect 29457 21023 29515 21029
rect 26786 20992 26792 21004
rect 25823 20964 26556 20992
rect 26747 20964 26792 20992
rect 25823 20961 25835 20964
rect 25777 20955 25835 20961
rect 26786 20952 26792 20964
rect 26844 20952 26850 21004
rect 27525 20995 27583 21001
rect 27525 20992 27537 20995
rect 27448 20964 27537 20992
rect 22704 20896 25452 20924
rect 25869 20927 25927 20933
rect 22704 20884 22710 20896
rect 23106 20856 23112 20868
rect 21284 20828 23112 20856
rect 23106 20816 23112 20828
rect 23164 20816 23170 20868
rect 23308 20865 23336 20896
rect 25869 20893 25881 20927
rect 25915 20924 25927 20927
rect 25958 20924 25964 20936
rect 25915 20896 25964 20924
rect 25915 20893 25927 20896
rect 25869 20887 25927 20893
rect 25958 20884 25964 20896
rect 26016 20924 26022 20936
rect 27062 20924 27068 20936
rect 26016 20896 27068 20924
rect 26016 20884 26022 20896
rect 27062 20884 27068 20896
rect 27120 20884 27126 20936
rect 23293 20859 23351 20865
rect 23293 20825 23305 20859
rect 23339 20825 23351 20859
rect 23293 20819 23351 20825
rect 25225 20859 25283 20865
rect 25225 20825 25237 20859
rect 25271 20856 25283 20859
rect 26142 20856 26148 20868
rect 25271 20828 26148 20856
rect 25271 20825 25283 20828
rect 25225 20819 25283 20825
rect 26142 20816 26148 20828
rect 26200 20816 26206 20868
rect 22094 20788 22100 20800
rect 19628 20760 22100 20788
rect 22094 20748 22100 20760
rect 22152 20748 22158 20800
rect 22738 20788 22744 20800
rect 22699 20760 22744 20788
rect 22738 20748 22744 20760
rect 22796 20748 22802 20800
rect 24762 20748 24768 20800
rect 24820 20788 24826 20800
rect 27448 20788 27476 20964
rect 27525 20961 27537 20964
rect 27571 20961 27583 20995
rect 27525 20955 27583 20961
rect 27614 20952 27620 21004
rect 27672 20992 27678 21004
rect 28077 20995 28135 21001
rect 28077 20992 28089 20995
rect 27672 20964 28089 20992
rect 27672 20952 27678 20964
rect 28077 20961 28089 20964
rect 28123 20992 28135 20995
rect 29089 20995 29147 21001
rect 29089 20992 29101 20995
rect 28123 20964 29101 20992
rect 28123 20961 28135 20964
rect 28077 20955 28135 20961
rect 29089 20961 29101 20964
rect 29135 20961 29147 20995
rect 29089 20955 29147 20961
rect 27706 20884 27712 20936
rect 27764 20924 27770 20936
rect 28353 20927 28411 20933
rect 28353 20924 28365 20927
rect 27764 20896 28365 20924
rect 27764 20884 27770 20896
rect 28353 20893 28365 20896
rect 28399 20924 28411 20927
rect 29472 20924 29500 21023
rect 30282 21020 30288 21072
rect 30340 21060 30346 21072
rect 32950 21060 32956 21072
rect 30340 21032 32956 21060
rect 30340 21020 30346 21032
rect 32950 21020 32956 21032
rect 33008 21020 33014 21072
rect 34790 21060 34796 21072
rect 34703 21032 34796 21060
rect 34790 21020 34796 21032
rect 34848 21060 34854 21072
rect 35250 21060 35256 21072
rect 34848 21032 35256 21060
rect 34848 21020 34854 21032
rect 35250 21020 35256 21032
rect 35308 21020 35314 21072
rect 30561 20995 30619 21001
rect 30561 20961 30573 20995
rect 30607 20961 30619 20995
rect 30561 20955 30619 20961
rect 31297 20995 31355 21001
rect 31297 20961 31309 20995
rect 31343 20992 31355 20995
rect 32306 20992 32312 21004
rect 31343 20964 32312 20992
rect 31343 20961 31355 20964
rect 31297 20955 31355 20961
rect 29822 20924 29828 20936
rect 28399 20896 29500 20924
rect 29783 20896 29828 20924
rect 28399 20893 28411 20896
rect 28353 20887 28411 20893
rect 29822 20884 29828 20896
rect 29880 20884 29886 20936
rect 30576 20924 30604 20955
rect 32306 20952 32312 20964
rect 32364 20952 32370 21004
rect 32401 20995 32459 21001
rect 32401 20961 32413 20995
rect 32447 20961 32459 20995
rect 32401 20955 32459 20961
rect 33137 20995 33195 21001
rect 33137 20961 33149 20995
rect 33183 20992 33195 20995
rect 33686 20992 33692 21004
rect 33183 20964 33692 20992
rect 33183 20961 33195 20964
rect 33137 20955 33195 20961
rect 32122 20924 32128 20936
rect 30576 20896 32128 20924
rect 32122 20884 32128 20896
rect 32180 20884 32186 20936
rect 32416 20924 32444 20955
rect 33686 20952 33692 20964
rect 33744 20952 33750 21004
rect 35805 20995 35863 21001
rect 35805 20961 35817 20995
rect 35851 20992 35863 20995
rect 36998 20992 37004 21004
rect 35851 20964 37004 20992
rect 35851 20961 35863 20964
rect 35805 20955 35863 20961
rect 36998 20952 37004 20964
rect 37056 20952 37062 21004
rect 37752 21001 37780 21100
rect 37737 20995 37795 21001
rect 37737 20961 37749 20995
rect 37783 20961 37795 20995
rect 37737 20955 37795 20961
rect 38105 20995 38163 21001
rect 38105 20961 38117 20995
rect 38151 20961 38163 20995
rect 38654 20992 38660 21004
rect 38615 20964 38660 20992
rect 38105 20955 38163 20961
rect 33410 20924 33416 20936
rect 32416 20896 33180 20924
rect 33371 20896 33416 20924
rect 33152 20868 33180 20896
rect 33410 20884 33416 20896
rect 33468 20884 33474 20936
rect 35529 20927 35587 20933
rect 35529 20893 35541 20927
rect 35575 20924 35587 20927
rect 36446 20924 36452 20936
rect 35575 20896 36452 20924
rect 35575 20893 35587 20896
rect 35529 20887 35587 20893
rect 36446 20884 36452 20896
rect 36504 20884 36510 20936
rect 37274 20884 37280 20936
rect 37332 20924 37338 20936
rect 37829 20927 37887 20933
rect 37829 20924 37841 20927
rect 37332 20896 37841 20924
rect 37332 20884 37338 20896
rect 37829 20893 37841 20896
rect 37875 20893 37887 20927
rect 37829 20887 37887 20893
rect 27801 20859 27859 20865
rect 27801 20825 27813 20859
rect 27847 20856 27859 20859
rect 27890 20856 27896 20868
rect 27847 20828 27896 20856
rect 27847 20825 27859 20828
rect 27801 20819 27859 20825
rect 27890 20816 27896 20828
rect 27948 20816 27954 20868
rect 29546 20856 29552 20868
rect 29012 20828 29552 20856
rect 29012 20788 29040 20828
rect 29546 20816 29552 20828
rect 29604 20816 29610 20868
rect 33134 20816 33140 20868
rect 33192 20816 33198 20868
rect 36538 20816 36544 20868
rect 36596 20856 36602 20868
rect 38120 20856 38148 20955
rect 38654 20952 38660 20964
rect 38712 20952 38718 21004
rect 36596 20828 38148 20856
rect 36596 20816 36602 20828
rect 24820 20760 29040 20788
rect 30745 20791 30803 20797
rect 24820 20748 24826 20760
rect 30745 20757 30757 20791
rect 30791 20788 30803 20791
rect 31202 20788 31208 20800
rect 30791 20760 31208 20788
rect 30791 20757 30803 20760
rect 30745 20751 30803 20757
rect 31202 20748 31208 20760
rect 31260 20748 31266 20800
rect 34238 20748 34244 20800
rect 34296 20788 34302 20800
rect 36630 20788 36636 20800
rect 34296 20760 36636 20788
rect 34296 20748 34302 20760
rect 36630 20748 36636 20760
rect 36688 20748 36694 20800
rect 36814 20748 36820 20800
rect 36872 20788 36878 20800
rect 36909 20791 36967 20797
rect 36909 20788 36921 20791
rect 36872 20760 36921 20788
rect 36872 20748 36878 20760
rect 36909 20757 36921 20760
rect 36955 20757 36967 20791
rect 36909 20751 36967 20757
rect 1104 20698 39836 20720
rect 1104 20646 4246 20698
rect 4298 20646 4310 20698
rect 4362 20646 4374 20698
rect 4426 20646 4438 20698
rect 4490 20646 34966 20698
rect 35018 20646 35030 20698
rect 35082 20646 35094 20698
rect 35146 20646 35158 20698
rect 35210 20646 39836 20698
rect 1104 20624 39836 20646
rect 2958 20584 2964 20596
rect 2919 20556 2964 20584
rect 2958 20544 2964 20556
rect 3016 20544 3022 20596
rect 3881 20587 3939 20593
rect 3881 20553 3893 20587
rect 3927 20584 3939 20587
rect 4614 20584 4620 20596
rect 3927 20556 4620 20584
rect 3927 20553 3939 20556
rect 3881 20547 3939 20553
rect 4614 20544 4620 20556
rect 4672 20544 4678 20596
rect 9493 20587 9551 20593
rect 9493 20553 9505 20587
rect 9539 20584 9551 20587
rect 9950 20584 9956 20596
rect 9539 20556 9956 20584
rect 9539 20553 9551 20556
rect 9493 20547 9551 20553
rect 9950 20544 9956 20556
rect 10008 20584 10014 20596
rect 12710 20584 12716 20596
rect 10008 20556 12716 20584
rect 10008 20544 10014 20556
rect 12710 20544 12716 20556
rect 12768 20544 12774 20596
rect 16298 20584 16304 20596
rect 16259 20556 16304 20584
rect 16298 20544 16304 20556
rect 16356 20544 16362 20596
rect 18598 20544 18604 20596
rect 18656 20584 18662 20596
rect 30282 20584 30288 20596
rect 18656 20556 30288 20584
rect 18656 20544 18662 20556
rect 30282 20544 30288 20556
rect 30340 20544 30346 20596
rect 38102 20584 38108 20596
rect 30392 20556 38108 20584
rect 10410 20476 10416 20528
rect 10468 20516 10474 20528
rect 10468 20488 10916 20516
rect 10468 20476 10474 20488
rect 4893 20451 4951 20457
rect 4893 20417 4905 20451
rect 4939 20448 4951 20451
rect 5074 20448 5080 20460
rect 4939 20420 5080 20448
rect 4939 20417 4951 20420
rect 4893 20411 4951 20417
rect 5074 20408 5080 20420
rect 5132 20408 5138 20460
rect 6822 20408 6828 20460
rect 6880 20448 6886 20460
rect 7929 20451 7987 20457
rect 7929 20448 7941 20451
rect 6880 20420 7941 20448
rect 6880 20408 6886 20420
rect 7929 20417 7941 20420
rect 7975 20448 7987 20451
rect 10226 20448 10232 20460
rect 7975 20420 10232 20448
rect 7975 20417 7987 20420
rect 7929 20411 7987 20417
rect 10226 20408 10232 20420
rect 10284 20408 10290 20460
rect 10686 20448 10692 20460
rect 10647 20420 10692 20448
rect 10686 20408 10692 20420
rect 10744 20408 10750 20460
rect 10888 20392 10916 20488
rect 15102 20476 15108 20528
rect 15160 20516 15166 20528
rect 20717 20519 20775 20525
rect 20717 20516 20729 20519
rect 15160 20488 20729 20516
rect 15160 20476 15166 20488
rect 20717 20485 20729 20488
rect 20763 20485 20775 20519
rect 23750 20516 23756 20528
rect 23711 20488 23756 20516
rect 20717 20479 20775 20485
rect 23750 20476 23756 20488
rect 23808 20476 23814 20528
rect 12434 20408 12440 20460
rect 12492 20448 12498 20460
rect 13170 20448 13176 20460
rect 12492 20420 12537 20448
rect 12912 20420 13176 20448
rect 12492 20408 12498 20420
rect 1394 20380 1400 20392
rect 1355 20352 1400 20380
rect 1394 20340 1400 20352
rect 1452 20340 1458 20392
rect 1673 20383 1731 20389
rect 1673 20349 1685 20383
rect 1719 20380 1731 20383
rect 2038 20380 2044 20392
rect 1719 20352 2044 20380
rect 1719 20349 1731 20352
rect 1673 20343 1731 20349
rect 2038 20340 2044 20352
rect 2096 20340 2102 20392
rect 3789 20383 3847 20389
rect 3789 20349 3801 20383
rect 3835 20380 3847 20383
rect 4062 20380 4068 20392
rect 3835 20352 4068 20380
rect 3835 20349 3847 20352
rect 3789 20343 3847 20349
rect 4062 20340 4068 20352
rect 4120 20380 4126 20392
rect 4617 20383 4675 20389
rect 4120 20352 4568 20380
rect 4120 20340 4126 20352
rect 3605 20315 3663 20321
rect 3605 20281 3617 20315
rect 3651 20312 3663 20315
rect 4154 20312 4160 20324
rect 3651 20284 4160 20312
rect 3651 20281 3663 20284
rect 3605 20275 3663 20281
rect 4154 20272 4160 20284
rect 4212 20272 4218 20324
rect 4540 20244 4568 20352
rect 4617 20349 4629 20383
rect 4663 20380 4675 20383
rect 5810 20380 5816 20392
rect 4663 20352 5816 20380
rect 4663 20349 4675 20352
rect 4617 20343 4675 20349
rect 5810 20340 5816 20352
rect 5868 20340 5874 20392
rect 8202 20380 8208 20392
rect 8163 20352 8208 20380
rect 8202 20340 8208 20352
rect 8260 20340 8266 20392
rect 10321 20383 10379 20389
rect 10321 20349 10333 20383
rect 10367 20349 10379 20383
rect 10321 20343 10379 20349
rect 10597 20383 10655 20389
rect 10597 20349 10609 20383
rect 10643 20349 10655 20383
rect 10870 20380 10876 20392
rect 10831 20352 10876 20380
rect 10597 20343 10655 20349
rect 5997 20247 6055 20253
rect 5997 20244 6009 20247
rect 4540 20216 6009 20244
rect 5997 20213 6009 20216
rect 6043 20213 6055 20247
rect 5997 20207 6055 20213
rect 9122 20204 9128 20256
rect 9180 20244 9186 20256
rect 10134 20244 10140 20256
rect 9180 20216 10140 20244
rect 9180 20204 9186 20216
rect 10134 20204 10140 20216
rect 10192 20244 10198 20256
rect 10336 20244 10364 20343
rect 10612 20312 10640 20343
rect 10870 20340 10876 20352
rect 10928 20340 10934 20392
rect 11698 20380 11704 20392
rect 11659 20352 11704 20380
rect 11698 20340 11704 20352
rect 11756 20340 11762 20392
rect 12912 20389 12940 20420
rect 13170 20408 13176 20420
rect 13228 20408 13234 20460
rect 13446 20408 13452 20460
rect 13504 20448 13510 20460
rect 14185 20451 14243 20457
rect 14185 20448 14197 20451
rect 13504 20420 14197 20448
rect 13504 20408 13510 20420
rect 14185 20417 14197 20420
rect 14231 20417 14243 20451
rect 14185 20411 14243 20417
rect 19058 20408 19064 20460
rect 19116 20448 19122 20460
rect 19426 20448 19432 20460
rect 19116 20420 19432 20448
rect 19116 20408 19122 20420
rect 19426 20408 19432 20420
rect 19484 20408 19490 20460
rect 26234 20408 26240 20460
rect 26292 20448 26298 20460
rect 26697 20451 26755 20457
rect 26697 20448 26709 20451
rect 26292 20420 26709 20448
rect 26292 20408 26298 20420
rect 26697 20417 26709 20420
rect 26743 20417 26755 20451
rect 26697 20411 26755 20417
rect 26786 20408 26792 20460
rect 26844 20448 26850 20460
rect 30098 20448 30104 20460
rect 26844 20420 30104 20448
rect 26844 20408 26850 20420
rect 12897 20383 12955 20389
rect 12897 20349 12909 20383
rect 12943 20349 12955 20383
rect 12897 20343 12955 20349
rect 13081 20383 13139 20389
rect 13081 20349 13093 20383
rect 13127 20349 13139 20383
rect 13262 20380 13268 20392
rect 13223 20352 13268 20380
rect 13081 20343 13139 20349
rect 11146 20312 11152 20324
rect 10612 20284 11152 20312
rect 11146 20272 11152 20284
rect 11204 20272 11210 20324
rect 11606 20272 11612 20324
rect 11664 20312 11670 20324
rect 13096 20312 13124 20343
rect 13262 20340 13268 20352
rect 13320 20380 13326 20392
rect 13722 20380 13728 20392
rect 13320 20352 13728 20380
rect 13320 20340 13326 20352
rect 13722 20340 13728 20352
rect 13780 20340 13786 20392
rect 13814 20340 13820 20392
rect 13872 20380 13878 20392
rect 13909 20383 13967 20389
rect 13909 20380 13921 20383
rect 13872 20352 13921 20380
rect 13872 20340 13878 20352
rect 13909 20349 13921 20352
rect 13955 20349 13967 20383
rect 13909 20343 13967 20349
rect 15010 20340 15016 20392
rect 15068 20380 15074 20392
rect 16025 20383 16083 20389
rect 16025 20380 16037 20383
rect 15068 20352 16037 20380
rect 15068 20340 15074 20352
rect 16025 20349 16037 20352
rect 16071 20349 16083 20383
rect 16025 20343 16083 20349
rect 16114 20340 16120 20392
rect 16172 20380 16178 20392
rect 17221 20383 17279 20389
rect 16172 20352 16217 20380
rect 16172 20340 16178 20352
rect 17221 20349 17233 20383
rect 17267 20380 17279 20383
rect 17494 20380 17500 20392
rect 17267 20352 17500 20380
rect 17267 20349 17279 20352
rect 17221 20343 17279 20349
rect 17494 20340 17500 20352
rect 17552 20340 17558 20392
rect 22922 20340 22928 20392
rect 22980 20380 22986 20392
rect 23661 20383 23719 20389
rect 23661 20380 23673 20383
rect 22980 20352 23673 20380
rect 22980 20340 22986 20352
rect 23661 20349 23673 20352
rect 23707 20349 23719 20383
rect 23661 20343 23719 20349
rect 24121 20383 24179 20389
rect 24121 20349 24133 20383
rect 24167 20349 24179 20383
rect 24121 20343 24179 20349
rect 11664 20284 13124 20312
rect 11664 20272 11670 20284
rect 18506 20272 18512 20324
rect 18564 20312 18570 20324
rect 18782 20312 18788 20324
rect 18564 20284 18788 20312
rect 18564 20272 18570 20284
rect 18782 20272 18788 20284
rect 18840 20272 18846 20324
rect 19426 20312 19432 20324
rect 19387 20284 19432 20312
rect 19426 20272 19432 20284
rect 19484 20272 19490 20324
rect 21634 20312 21640 20324
rect 21595 20284 21640 20312
rect 21634 20272 21640 20284
rect 21692 20272 21698 20324
rect 23385 20315 23443 20321
rect 23385 20281 23397 20315
rect 23431 20281 23443 20315
rect 24136 20312 24164 20343
rect 24210 20340 24216 20392
rect 24268 20380 24274 20392
rect 24397 20383 24455 20389
rect 24397 20380 24409 20383
rect 24268 20352 24409 20380
rect 24268 20340 24274 20352
rect 24397 20349 24409 20352
rect 24443 20349 24455 20383
rect 24854 20380 24860 20392
rect 24815 20352 24860 20380
rect 24397 20343 24455 20349
rect 24854 20340 24860 20352
rect 24912 20340 24918 20392
rect 25593 20383 25651 20389
rect 25593 20349 25605 20383
rect 25639 20380 25651 20383
rect 25682 20380 25688 20392
rect 25639 20352 25688 20380
rect 25639 20349 25651 20352
rect 25593 20343 25651 20349
rect 25682 20340 25688 20352
rect 25740 20340 25746 20392
rect 26418 20380 26424 20392
rect 26379 20352 26424 20380
rect 26418 20340 26424 20352
rect 26476 20340 26482 20392
rect 28552 20389 28580 20420
rect 30098 20408 30104 20420
rect 30156 20408 30162 20460
rect 30392 20457 30420 20556
rect 38102 20544 38108 20556
rect 38160 20544 38166 20596
rect 31386 20516 31392 20528
rect 31347 20488 31392 20516
rect 31386 20476 31392 20488
rect 31444 20476 31450 20528
rect 30377 20451 30435 20457
rect 30377 20417 30389 20451
rect 30423 20417 30435 20451
rect 32122 20448 32128 20460
rect 32083 20420 32128 20448
rect 30377 20411 30435 20417
rect 32122 20408 32128 20420
rect 32180 20408 32186 20460
rect 33134 20448 33140 20460
rect 32600 20420 33140 20448
rect 28537 20383 28595 20389
rect 28537 20349 28549 20383
rect 28583 20349 28595 20383
rect 28537 20343 28595 20349
rect 29178 20340 29184 20392
rect 29236 20340 29242 20392
rect 29546 20380 29552 20392
rect 29507 20352 29552 20380
rect 29546 20340 29552 20352
rect 29604 20340 29610 20392
rect 30466 20380 30472 20392
rect 30427 20352 30472 20380
rect 30466 20340 30472 20352
rect 30524 20340 30530 20392
rect 30558 20340 30564 20392
rect 30616 20380 30622 20392
rect 30929 20383 30987 20389
rect 30929 20380 30941 20383
rect 30616 20352 30941 20380
rect 30616 20340 30622 20352
rect 30929 20349 30941 20352
rect 30975 20349 30987 20383
rect 30929 20343 30987 20349
rect 31018 20340 31024 20392
rect 31076 20380 31082 20392
rect 31478 20380 31484 20392
rect 31076 20352 31484 20380
rect 31076 20340 31082 20352
rect 31478 20340 31484 20352
rect 31536 20340 31542 20392
rect 32600 20389 32628 20420
rect 33134 20408 33140 20420
rect 33192 20448 33198 20460
rect 34238 20448 34244 20460
rect 33192 20420 34244 20448
rect 33192 20408 33198 20420
rect 34238 20408 34244 20420
rect 34296 20408 34302 20460
rect 36446 20448 36452 20460
rect 36407 20420 36452 20448
rect 36446 20408 36452 20420
rect 36504 20408 36510 20460
rect 32585 20383 32643 20389
rect 32585 20349 32597 20383
rect 32631 20349 32643 20383
rect 32585 20343 32643 20349
rect 32769 20383 32827 20389
rect 32769 20349 32781 20383
rect 32815 20380 32827 20383
rect 32858 20380 32864 20392
rect 32815 20352 32864 20380
rect 32815 20349 32827 20352
rect 32769 20343 32827 20349
rect 32858 20340 32864 20352
rect 32916 20340 32922 20392
rect 32953 20383 33011 20389
rect 32953 20349 32965 20383
rect 32999 20349 33011 20383
rect 32953 20343 33011 20349
rect 24486 20312 24492 20324
rect 24136 20284 24492 20312
rect 23385 20275 23443 20281
rect 11624 20244 11652 20272
rect 11790 20244 11796 20256
rect 10192 20216 11652 20244
rect 11751 20216 11796 20244
rect 10192 20204 10198 20216
rect 11790 20204 11796 20216
rect 11848 20204 11854 20256
rect 15286 20244 15292 20256
rect 15247 20216 15292 20244
rect 15286 20204 15292 20216
rect 15344 20204 15350 20256
rect 17405 20247 17463 20253
rect 17405 20213 17417 20247
rect 17451 20244 17463 20247
rect 18690 20244 18696 20256
rect 17451 20216 18696 20244
rect 17451 20213 17463 20216
rect 17405 20207 17463 20213
rect 18690 20204 18696 20216
rect 18748 20204 18754 20256
rect 18800 20244 18828 20272
rect 22830 20244 22836 20256
rect 18800 20216 22836 20244
rect 22830 20204 22836 20216
rect 22888 20204 22894 20256
rect 23400 20244 23428 20275
rect 24486 20272 24492 20284
rect 24544 20272 24550 20324
rect 29196 20312 29224 20340
rect 27356 20284 29224 20312
rect 24394 20244 24400 20256
rect 23400 20216 24400 20244
rect 24394 20204 24400 20216
rect 24452 20244 24458 20256
rect 27356 20244 27384 20284
rect 29270 20272 29276 20324
rect 29328 20312 29334 20324
rect 30576 20312 30604 20340
rect 29328 20284 30604 20312
rect 29328 20272 29334 20284
rect 32306 20272 32312 20324
rect 32364 20312 32370 20324
rect 32968 20312 32996 20343
rect 33502 20340 33508 20392
rect 33560 20380 33566 20392
rect 33597 20383 33655 20389
rect 33597 20380 33609 20383
rect 33560 20352 33609 20380
rect 33560 20340 33566 20352
rect 33597 20349 33609 20352
rect 33643 20349 33655 20383
rect 33597 20343 33655 20349
rect 34149 20383 34207 20389
rect 34149 20349 34161 20383
rect 34195 20380 34207 20383
rect 34790 20380 34796 20392
rect 34195 20352 34796 20380
rect 34195 20349 34207 20352
rect 34149 20343 34207 20349
rect 34790 20340 34796 20352
rect 34848 20340 34854 20392
rect 35161 20383 35219 20389
rect 35161 20349 35173 20383
rect 35207 20380 35219 20383
rect 35250 20380 35256 20392
rect 35207 20352 35256 20380
rect 35207 20349 35219 20352
rect 35161 20343 35219 20349
rect 35250 20340 35256 20352
rect 35308 20340 35314 20392
rect 35437 20383 35495 20389
rect 35437 20349 35449 20383
rect 35483 20380 35495 20383
rect 36170 20380 36176 20392
rect 35483 20352 36176 20380
rect 35483 20349 35495 20352
rect 35437 20343 35495 20349
rect 36170 20340 36176 20352
rect 36228 20340 36234 20392
rect 36725 20383 36783 20389
rect 36725 20349 36737 20383
rect 36771 20380 36783 20383
rect 37734 20380 37740 20392
rect 36771 20352 37740 20380
rect 36771 20349 36783 20352
rect 36725 20343 36783 20349
rect 37734 20340 37740 20352
rect 37792 20340 37798 20392
rect 38286 20340 38292 20392
rect 38344 20380 38350 20392
rect 38565 20383 38623 20389
rect 38565 20380 38577 20383
rect 38344 20352 38577 20380
rect 38344 20340 38350 20352
rect 38565 20349 38577 20352
rect 38611 20349 38623 20383
rect 38565 20343 38623 20349
rect 32364 20284 33732 20312
rect 32364 20272 32370 20284
rect 24452 20216 27384 20244
rect 24452 20204 24458 20216
rect 27706 20204 27712 20256
rect 27764 20244 27770 20256
rect 27801 20247 27859 20253
rect 27801 20244 27813 20247
rect 27764 20216 27813 20244
rect 27764 20204 27770 20216
rect 27801 20213 27813 20216
rect 27847 20213 27859 20247
rect 27801 20207 27859 20213
rect 28629 20247 28687 20253
rect 28629 20213 28641 20247
rect 28675 20244 28687 20247
rect 29178 20244 29184 20256
rect 28675 20216 29184 20244
rect 28675 20213 28687 20216
rect 28629 20207 28687 20213
rect 29178 20204 29184 20216
rect 29236 20204 29242 20256
rect 29733 20247 29791 20253
rect 29733 20213 29745 20247
rect 29779 20244 29791 20247
rect 30006 20244 30012 20256
rect 29779 20216 30012 20244
rect 29779 20213 29791 20216
rect 29733 20207 29791 20213
rect 30006 20204 30012 20216
rect 30064 20204 30070 20256
rect 33704 20253 33732 20284
rect 33689 20247 33747 20253
rect 33689 20213 33701 20247
rect 33735 20213 33747 20247
rect 33689 20207 33747 20213
rect 34698 20204 34704 20256
rect 34756 20244 34762 20256
rect 34977 20247 35035 20253
rect 34977 20244 34989 20247
rect 34756 20216 34989 20244
rect 34756 20204 34762 20216
rect 34977 20213 34989 20216
rect 35023 20213 35035 20247
rect 34977 20207 35035 20213
rect 36998 20204 37004 20256
rect 37056 20244 37062 20256
rect 37829 20247 37887 20253
rect 37829 20244 37841 20247
rect 37056 20216 37841 20244
rect 37056 20204 37062 20216
rect 37829 20213 37841 20216
rect 37875 20213 37887 20247
rect 37829 20207 37887 20213
rect 38657 20247 38715 20253
rect 38657 20213 38669 20247
rect 38703 20244 38715 20247
rect 38746 20244 38752 20256
rect 38703 20216 38752 20244
rect 38703 20213 38715 20216
rect 38657 20207 38715 20213
rect 38746 20204 38752 20216
rect 38804 20204 38810 20256
rect 1104 20154 39836 20176
rect 1104 20102 19606 20154
rect 19658 20102 19670 20154
rect 19722 20102 19734 20154
rect 19786 20102 19798 20154
rect 19850 20102 39836 20154
rect 1104 20080 39836 20102
rect 10134 20040 10140 20052
rect 10095 20012 10140 20040
rect 10134 20000 10140 20012
rect 10192 20000 10198 20052
rect 11422 20000 11428 20052
rect 11480 20040 11486 20052
rect 11480 20012 16160 20040
rect 11480 20000 11486 20012
rect 2958 19972 2964 19984
rect 2608 19944 2964 19972
rect 2608 19913 2636 19944
rect 2958 19932 2964 19944
rect 3016 19932 3022 19984
rect 8113 19975 8171 19981
rect 3160 19944 5028 19972
rect 2593 19907 2651 19913
rect 2593 19873 2605 19907
rect 2639 19873 2651 19907
rect 2593 19867 2651 19873
rect 2869 19907 2927 19913
rect 2869 19873 2881 19907
rect 2915 19873 2927 19907
rect 2869 19867 2927 19873
rect 2884 19836 2912 19867
rect 3160 19836 3188 19944
rect 5000 19916 5028 19944
rect 8113 19941 8125 19975
rect 8159 19972 8171 19975
rect 8202 19972 8208 19984
rect 8159 19944 8208 19972
rect 8159 19941 8171 19944
rect 8113 19935 8171 19941
rect 8202 19932 8208 19944
rect 8260 19932 8266 19984
rect 9122 19932 9128 19984
rect 9180 19932 9186 19984
rect 13078 19932 13084 19984
rect 13136 19972 13142 19984
rect 16132 19981 16160 20012
rect 17218 20000 17224 20052
rect 17276 20040 17282 20052
rect 17770 20040 17776 20052
rect 17276 20012 17776 20040
rect 17276 20000 17282 20012
rect 17770 20000 17776 20012
rect 17828 20040 17834 20052
rect 17828 20012 19196 20040
rect 17828 20000 17834 20012
rect 13173 19975 13231 19981
rect 13173 19972 13185 19975
rect 13136 19944 13185 19972
rect 13136 19932 13142 19944
rect 13173 19941 13185 19944
rect 13219 19941 13231 19975
rect 13173 19935 13231 19941
rect 16117 19975 16175 19981
rect 16117 19941 16129 19975
rect 16163 19941 16175 19975
rect 16117 19935 16175 19941
rect 17310 19932 17316 19984
rect 17368 19972 17374 19984
rect 19168 19972 19196 20012
rect 19978 20000 19984 20052
rect 20036 20040 20042 20052
rect 20349 20043 20407 20049
rect 20349 20040 20361 20043
rect 20036 20012 20361 20040
rect 20036 20000 20042 20012
rect 20349 20009 20361 20012
rect 20395 20009 20407 20043
rect 24762 20040 24768 20052
rect 20349 20003 20407 20009
rect 22756 20012 24768 20040
rect 19702 19972 19708 19984
rect 17368 19944 18920 19972
rect 17368 19932 17374 19944
rect 3326 19904 3332 19916
rect 3239 19876 3332 19904
rect 3326 19864 3332 19876
rect 3384 19904 3390 19916
rect 4062 19904 4068 19916
rect 3384 19876 3924 19904
rect 4023 19876 4068 19904
rect 3384 19864 3390 19876
rect 3510 19836 3516 19848
rect 2884 19808 3188 19836
rect 3471 19808 3516 19836
rect 3510 19796 3516 19808
rect 3568 19796 3574 19848
rect 3896 19836 3924 19876
rect 4062 19864 4068 19876
rect 4120 19864 4126 19916
rect 4798 19904 4804 19916
rect 4759 19876 4804 19904
rect 4798 19864 4804 19876
rect 4856 19864 4862 19916
rect 4982 19904 4988 19916
rect 4943 19876 4988 19904
rect 4982 19864 4988 19876
rect 5040 19864 5046 19916
rect 5721 19907 5779 19913
rect 5721 19873 5733 19907
rect 5767 19904 5779 19907
rect 5810 19904 5816 19916
rect 5767 19876 5816 19904
rect 5767 19873 5779 19876
rect 5721 19867 5779 19873
rect 5810 19864 5816 19876
rect 5868 19904 5874 19916
rect 6822 19904 6828 19916
rect 5868 19876 6828 19904
rect 5868 19864 5874 19876
rect 6822 19864 6828 19876
rect 6880 19864 6886 19916
rect 8662 19904 8668 19916
rect 8623 19876 8668 19904
rect 8662 19864 8668 19876
rect 8720 19864 8726 19916
rect 8941 19907 8999 19913
rect 8941 19873 8953 19907
rect 8987 19904 8999 19907
rect 9140 19904 9168 19932
rect 9950 19904 9956 19916
rect 8987 19876 9168 19904
rect 9911 19876 9956 19904
rect 8987 19873 8999 19876
rect 8941 19867 8999 19873
rect 9950 19864 9956 19876
rect 10008 19864 10014 19916
rect 10686 19904 10692 19916
rect 10647 19876 10692 19904
rect 10686 19864 10692 19876
rect 10744 19864 10750 19916
rect 11790 19904 11796 19916
rect 11751 19876 11796 19904
rect 11790 19864 11796 19876
rect 11848 19864 11854 19916
rect 14182 19904 14188 19916
rect 14143 19876 14188 19904
rect 14182 19864 14188 19876
rect 14240 19864 14246 19916
rect 15194 19864 15200 19916
rect 15252 19904 15258 19916
rect 15289 19907 15347 19913
rect 15289 19904 15301 19907
rect 15252 19876 15301 19904
rect 15252 19864 15258 19876
rect 15289 19873 15301 19876
rect 15335 19873 15347 19907
rect 15289 19867 15347 19873
rect 16206 19864 16212 19916
rect 16264 19904 16270 19916
rect 16577 19907 16635 19913
rect 16577 19904 16589 19907
rect 16264 19876 16589 19904
rect 16264 19864 16270 19876
rect 16577 19873 16589 19876
rect 16623 19873 16635 19907
rect 16850 19904 16856 19916
rect 16811 19876 16856 19904
rect 16577 19867 16635 19873
rect 3970 19836 3976 19848
rect 3883 19808 3976 19836
rect 3970 19796 3976 19808
rect 4028 19836 4034 19848
rect 4816 19836 4844 19864
rect 5994 19836 6000 19848
rect 4028 19808 4844 19836
rect 5955 19808 6000 19836
rect 4028 19796 4034 19808
rect 5994 19796 6000 19808
rect 6052 19796 6058 19848
rect 9125 19839 9183 19845
rect 9125 19805 9137 19839
rect 9171 19836 9183 19839
rect 10870 19836 10876 19848
rect 9171 19808 10876 19836
rect 9171 19805 9183 19808
rect 9125 19799 9183 19805
rect 10870 19796 10876 19808
rect 10928 19796 10934 19848
rect 11517 19839 11575 19845
rect 11517 19805 11529 19839
rect 11563 19805 11575 19839
rect 11517 19799 11575 19805
rect 4341 19771 4399 19777
rect 4341 19737 4353 19771
rect 4387 19768 4399 19771
rect 4706 19768 4712 19780
rect 4387 19740 4712 19768
rect 4387 19737 4399 19740
rect 4341 19731 4399 19737
rect 4706 19728 4712 19740
rect 4764 19728 4770 19780
rect 10226 19728 10232 19780
rect 10284 19768 10290 19780
rect 11532 19768 11560 19799
rect 12434 19796 12440 19848
rect 12492 19836 12498 19848
rect 14093 19839 14151 19845
rect 14093 19836 14105 19839
rect 12492 19808 14105 19836
rect 12492 19796 12498 19808
rect 14093 19805 14105 19808
rect 14139 19836 14151 19839
rect 14734 19836 14740 19848
rect 14139 19808 14740 19836
rect 14139 19805 14151 19808
rect 14093 19799 14151 19805
rect 14734 19796 14740 19808
rect 14792 19836 14798 19848
rect 16592 19836 16620 19867
rect 16850 19864 16856 19876
rect 16908 19864 16914 19916
rect 16942 19864 16948 19916
rect 17000 19904 17006 19916
rect 17126 19904 17132 19916
rect 17000 19876 17045 19904
rect 17087 19876 17132 19904
rect 17000 19864 17006 19876
rect 17126 19864 17132 19876
rect 17184 19864 17190 19916
rect 17494 19904 17500 19916
rect 17455 19876 17500 19904
rect 17494 19864 17500 19876
rect 17552 19864 17558 19916
rect 17678 19904 17684 19916
rect 17591 19876 17684 19904
rect 16666 19836 16672 19848
rect 14792 19808 15516 19836
rect 16579 19808 16672 19836
rect 14792 19796 14798 19808
rect 14826 19768 14832 19780
rect 10284 19740 11560 19768
rect 14016 19740 14832 19768
rect 10284 19728 10290 19740
rect 7098 19700 7104 19712
rect 7059 19672 7104 19700
rect 7098 19660 7104 19672
rect 7156 19660 7162 19712
rect 10873 19703 10931 19709
rect 10873 19669 10885 19703
rect 10919 19700 10931 19703
rect 14016 19700 14044 19740
rect 14826 19728 14832 19740
rect 14884 19728 14890 19780
rect 15488 19777 15516 19808
rect 16666 19796 16672 19808
rect 16724 19836 16730 19848
rect 17604 19836 17632 19876
rect 17678 19864 17684 19876
rect 17736 19864 17742 19916
rect 18598 19904 18604 19916
rect 18559 19876 18604 19904
rect 18598 19864 18604 19876
rect 18656 19864 18662 19916
rect 18892 19913 18920 19944
rect 19168 19944 19708 19972
rect 19168 19913 19196 19944
rect 19702 19932 19708 19944
rect 19760 19932 19766 19984
rect 20180 19944 22048 19972
rect 20180 19913 20208 19944
rect 18693 19907 18751 19913
rect 18693 19873 18705 19907
rect 18739 19873 18751 19907
rect 18693 19867 18751 19873
rect 18877 19907 18935 19913
rect 18877 19873 18889 19907
rect 18923 19873 18935 19907
rect 18877 19867 18935 19873
rect 19153 19907 19211 19913
rect 19153 19873 19165 19907
rect 19199 19873 19211 19907
rect 19153 19867 19211 19873
rect 19337 19907 19395 19913
rect 19337 19873 19349 19907
rect 19383 19873 19395 19907
rect 19337 19867 19395 19873
rect 20165 19907 20223 19913
rect 20165 19873 20177 19907
rect 20211 19873 20223 19907
rect 20165 19867 20223 19873
rect 16724 19808 17632 19836
rect 18049 19839 18107 19845
rect 16724 19796 16730 19808
rect 18049 19805 18061 19839
rect 18095 19836 18107 19839
rect 18138 19836 18144 19848
rect 18095 19808 18144 19836
rect 18095 19805 18107 19808
rect 18049 19799 18107 19805
rect 18138 19796 18144 19808
rect 18196 19796 18202 19848
rect 18506 19796 18512 19848
rect 18564 19836 18570 19848
rect 18708 19836 18736 19867
rect 18564 19808 18736 19836
rect 18564 19796 18570 19808
rect 18782 19796 18788 19848
rect 18840 19836 18846 19848
rect 19352 19836 19380 19867
rect 20346 19864 20352 19916
rect 20404 19904 20410 19916
rect 20901 19907 20959 19913
rect 20901 19904 20913 19907
rect 20404 19876 20913 19904
rect 20404 19864 20410 19876
rect 20901 19873 20913 19876
rect 20947 19873 20959 19907
rect 22020 19904 22048 19944
rect 22557 19907 22615 19913
rect 22020 19876 22508 19904
rect 20901 19867 20959 19873
rect 18840 19808 19380 19836
rect 18840 19796 18846 19808
rect 19794 19796 19800 19848
rect 19852 19836 19858 19848
rect 20806 19836 20812 19848
rect 19852 19808 20812 19836
rect 19852 19796 19858 19808
rect 20806 19796 20812 19808
rect 20864 19796 20870 19848
rect 21910 19836 21916 19848
rect 21871 19808 21916 19836
rect 21910 19796 21916 19808
rect 21968 19796 21974 19848
rect 22278 19796 22284 19848
rect 22336 19836 22342 19848
rect 22373 19839 22431 19845
rect 22373 19836 22385 19839
rect 22336 19808 22385 19836
rect 22336 19796 22342 19808
rect 22373 19805 22385 19808
rect 22419 19805 22431 19839
rect 22373 19799 22431 19805
rect 15473 19771 15531 19777
rect 15473 19737 15485 19771
rect 15519 19737 15531 19771
rect 15473 19731 15531 19737
rect 17494 19728 17500 19780
rect 17552 19768 17558 19780
rect 20346 19768 20352 19780
rect 17552 19740 20352 19768
rect 17552 19728 17558 19740
rect 20346 19728 20352 19740
rect 20404 19728 20410 19780
rect 22480 19768 22508 19876
rect 22557 19873 22569 19907
rect 22603 19873 22615 19907
rect 22756 19904 22784 20012
rect 24762 20000 24768 20012
rect 24820 20000 24826 20052
rect 25869 20043 25927 20049
rect 25869 20009 25881 20043
rect 25915 20040 25927 20043
rect 25958 20040 25964 20052
rect 25915 20012 25964 20040
rect 25915 20009 25927 20012
rect 25869 20003 25927 20009
rect 25958 20000 25964 20012
rect 26016 20000 26022 20052
rect 29362 20040 29368 20052
rect 26068 20012 29368 20040
rect 22830 19932 22836 19984
rect 22888 19972 22894 19984
rect 26068 19972 26096 20012
rect 29362 20000 29368 20012
rect 29420 20000 29426 20052
rect 31662 20040 31668 20052
rect 29656 20012 31668 20040
rect 27706 19972 27712 19984
rect 22888 19944 24256 19972
rect 22888 19932 22894 19944
rect 22925 19907 22983 19913
rect 22925 19904 22937 19907
rect 22756 19876 22937 19904
rect 22557 19867 22615 19873
rect 22925 19873 22937 19876
rect 22971 19873 22983 19907
rect 22925 19867 22983 19873
rect 22572 19836 22600 19867
rect 23014 19864 23020 19916
rect 23072 19904 23078 19916
rect 24228 19913 24256 19944
rect 24504 19944 26096 19972
rect 27080 19944 27712 19972
rect 24213 19907 24271 19913
rect 23072 19876 23117 19904
rect 23072 19864 23078 19876
rect 24213 19873 24225 19907
rect 24259 19873 24271 19907
rect 24213 19867 24271 19873
rect 22830 19836 22836 19848
rect 22572 19808 22836 19836
rect 22830 19796 22836 19808
rect 22888 19796 22894 19848
rect 24504 19836 24532 19944
rect 24578 19864 24584 19916
rect 24636 19904 24642 19916
rect 24636 19876 24681 19904
rect 24636 19864 24642 19876
rect 25498 19864 25504 19916
rect 25556 19904 25562 19916
rect 27080 19913 27108 19944
rect 27706 19932 27712 19944
rect 27764 19932 27770 19984
rect 25777 19907 25835 19913
rect 25777 19904 25789 19907
rect 25556 19876 25789 19904
rect 25556 19864 25562 19876
rect 25777 19873 25789 19876
rect 25823 19904 25835 19907
rect 27065 19907 27123 19913
rect 27065 19904 27077 19907
rect 25823 19876 27077 19904
rect 25823 19873 25835 19876
rect 25777 19867 25835 19873
rect 27065 19873 27077 19876
rect 27111 19873 27123 19907
rect 27614 19904 27620 19916
rect 27575 19876 27620 19904
rect 27065 19867 27123 19873
rect 27614 19864 27620 19876
rect 27672 19864 27678 19916
rect 27890 19904 27896 19916
rect 27851 19876 27896 19904
rect 27890 19864 27896 19876
rect 27948 19864 27954 19916
rect 29656 19913 29684 20012
rect 31662 20000 31668 20012
rect 31720 20000 31726 20052
rect 34330 20040 34336 20052
rect 33336 20012 34336 20040
rect 30098 19932 30104 19984
rect 30156 19972 30162 19984
rect 32677 19975 32735 19981
rect 32677 19972 32689 19975
rect 30156 19944 32689 19972
rect 30156 19932 30162 19944
rect 32677 19941 32689 19944
rect 32723 19941 32735 19975
rect 32677 19935 32735 19941
rect 29641 19907 29699 19913
rect 29641 19873 29653 19907
rect 29687 19873 29699 19907
rect 29641 19867 29699 19873
rect 29730 19864 29736 19916
rect 29788 19904 29794 19916
rect 29917 19907 29975 19913
rect 29917 19904 29929 19907
rect 29788 19876 29929 19904
rect 29788 19864 29794 19876
rect 29917 19873 29929 19876
rect 29963 19873 29975 19907
rect 30650 19904 30656 19916
rect 30611 19876 30656 19904
rect 29917 19867 29975 19873
rect 30650 19864 30656 19876
rect 30708 19864 30714 19916
rect 30742 19864 30748 19916
rect 30800 19904 30806 19916
rect 31205 19907 31263 19913
rect 31205 19904 31217 19907
rect 30800 19876 31217 19904
rect 30800 19864 30806 19876
rect 31205 19873 31217 19876
rect 31251 19873 31263 19907
rect 32214 19904 32220 19916
rect 32175 19876 32220 19904
rect 31205 19867 31263 19873
rect 32214 19864 32220 19876
rect 32272 19864 32278 19916
rect 33336 19913 33364 20012
rect 34330 20000 34336 20012
rect 34388 20000 34394 20052
rect 35621 20043 35679 20049
rect 35621 20009 35633 20043
rect 35667 20040 35679 20043
rect 36906 20040 36912 20052
rect 35667 20012 36912 20040
rect 35667 20009 35679 20012
rect 35621 20003 35679 20009
rect 36906 20000 36912 20012
rect 36964 20040 36970 20052
rect 36964 20012 38424 20040
rect 36964 20000 36970 20012
rect 36538 19972 36544 19984
rect 33888 19944 36544 19972
rect 33888 19913 33916 19944
rect 36538 19932 36544 19944
rect 36596 19932 36602 19984
rect 36814 19972 36820 19984
rect 36648 19944 36820 19972
rect 33321 19907 33379 19913
rect 33321 19873 33333 19907
rect 33367 19873 33379 19907
rect 33321 19867 33379 19873
rect 33873 19907 33931 19913
rect 33873 19873 33885 19907
rect 33919 19873 33931 19907
rect 33873 19867 33931 19873
rect 33965 19907 34023 19913
rect 33965 19873 33977 19907
rect 34011 19873 34023 19907
rect 34422 19904 34428 19916
rect 34383 19876 34428 19904
rect 33965 19867 34023 19873
rect 23860 19808 24532 19836
rect 24673 19839 24731 19845
rect 23860 19768 23888 19808
rect 24673 19805 24685 19839
rect 24719 19805 24731 19839
rect 27982 19836 27988 19848
rect 27943 19808 27988 19836
rect 24673 19799 24731 19805
rect 24026 19768 24032 19780
rect 22480 19740 23888 19768
rect 23987 19740 24032 19768
rect 24026 19728 24032 19740
rect 24084 19728 24090 19780
rect 24118 19728 24124 19780
rect 24176 19768 24182 19780
rect 24688 19768 24716 19799
rect 27982 19796 27988 19808
rect 28040 19796 28046 19848
rect 29273 19839 29331 19845
rect 29273 19805 29285 19839
rect 29319 19836 29331 19839
rect 30466 19836 30472 19848
rect 29319 19808 30472 19836
rect 29319 19805 29331 19808
rect 29273 19799 29331 19805
rect 30466 19796 30472 19808
rect 30524 19796 30530 19848
rect 31021 19839 31079 19845
rect 31021 19805 31033 19839
rect 31067 19805 31079 19839
rect 32122 19836 32128 19848
rect 32083 19808 32128 19836
rect 31021 19799 31079 19805
rect 29917 19771 29975 19777
rect 29917 19768 29929 19771
rect 24176 19740 29929 19768
rect 24176 19728 24182 19740
rect 29917 19737 29929 19740
rect 29963 19737 29975 19771
rect 31036 19768 31064 19799
rect 32122 19796 32128 19808
rect 32180 19796 32186 19848
rect 33410 19836 33416 19848
rect 33371 19808 33416 19836
rect 33410 19796 33416 19808
rect 33468 19796 33474 19848
rect 32030 19768 32036 19780
rect 31036 19740 32036 19768
rect 29917 19731 29975 19737
rect 32030 19728 32036 19740
rect 32088 19768 32094 19780
rect 33980 19768 34008 19867
rect 34422 19864 34428 19876
rect 34480 19864 34486 19916
rect 35161 19907 35219 19913
rect 35161 19873 35173 19907
rect 35207 19904 35219 19907
rect 35621 19907 35679 19913
rect 35621 19904 35633 19907
rect 35207 19876 35633 19904
rect 35207 19873 35219 19876
rect 35161 19867 35219 19873
rect 35621 19873 35633 19876
rect 35667 19873 35679 19907
rect 35621 19867 35679 19873
rect 35713 19907 35771 19913
rect 35713 19873 35725 19907
rect 35759 19873 35771 19907
rect 35713 19867 35771 19873
rect 35728 19836 35756 19867
rect 35802 19864 35808 19916
rect 35860 19904 35866 19916
rect 36648 19913 36676 19944
rect 36814 19932 36820 19944
rect 36872 19972 36878 19984
rect 37734 19972 37740 19984
rect 36872 19944 37136 19972
rect 37695 19944 37740 19972
rect 36872 19932 36878 19944
rect 36265 19907 36323 19913
rect 36265 19904 36277 19907
rect 35860 19876 36277 19904
rect 35860 19864 35866 19876
rect 36265 19873 36277 19876
rect 36311 19873 36323 19907
rect 36265 19867 36323 19873
rect 36633 19907 36691 19913
rect 36633 19873 36645 19907
rect 36679 19873 36691 19907
rect 36633 19867 36691 19873
rect 36909 19907 36967 19913
rect 36909 19873 36921 19907
rect 36955 19904 36967 19907
rect 36998 19904 37004 19916
rect 36955 19876 37004 19904
rect 36955 19873 36967 19876
rect 36909 19867 36967 19873
rect 35894 19836 35900 19848
rect 35728 19808 35900 19836
rect 35894 19796 35900 19808
rect 35952 19796 35958 19848
rect 36173 19839 36231 19845
rect 36173 19805 36185 19839
rect 36219 19836 36231 19839
rect 36722 19836 36728 19848
rect 36219 19808 36728 19836
rect 36219 19805 36231 19808
rect 36173 19799 36231 19805
rect 36722 19796 36728 19808
rect 36780 19796 36786 19848
rect 32088 19740 34008 19768
rect 32088 19728 32094 19740
rect 36262 19728 36268 19780
rect 36320 19768 36326 19780
rect 36924 19768 36952 19867
rect 36998 19864 37004 19876
rect 37056 19864 37062 19916
rect 37108 19836 37136 19944
rect 37734 19932 37740 19944
rect 37792 19932 37798 19984
rect 38396 19972 38424 20012
rect 38396 19944 38516 19972
rect 37182 19864 37188 19916
rect 37240 19904 37246 19916
rect 38488 19913 38516 19944
rect 38381 19907 38439 19913
rect 38381 19904 38393 19907
rect 37240 19876 38393 19904
rect 37240 19864 37246 19876
rect 38381 19873 38393 19876
rect 38427 19873 38439 19907
rect 38381 19867 38439 19873
rect 38473 19907 38531 19913
rect 38473 19873 38485 19907
rect 38519 19873 38531 19907
rect 38746 19904 38752 19916
rect 38707 19876 38752 19904
rect 38473 19867 38531 19873
rect 38746 19864 38752 19876
rect 38804 19864 38810 19916
rect 38286 19836 38292 19848
rect 37108 19808 38292 19836
rect 38286 19796 38292 19808
rect 38344 19796 38350 19848
rect 38841 19839 38899 19845
rect 38841 19805 38853 19839
rect 38887 19805 38899 19839
rect 38841 19799 38899 19805
rect 38856 19768 38884 19799
rect 38930 19768 38936 19780
rect 36320 19740 38936 19768
rect 36320 19728 36326 19740
rect 38930 19728 38936 19740
rect 38988 19728 38994 19780
rect 10919 19672 14044 19700
rect 10919 19669 10931 19672
rect 10873 19663 10931 19669
rect 14090 19660 14096 19712
rect 14148 19700 14154 19712
rect 14369 19703 14427 19709
rect 14369 19700 14381 19703
rect 14148 19672 14381 19700
rect 14148 19660 14154 19672
rect 14369 19669 14381 19672
rect 14415 19669 14427 19703
rect 14369 19663 14427 19669
rect 17865 19703 17923 19709
rect 17865 19669 17877 19703
rect 17911 19700 17923 19703
rect 19334 19700 19340 19712
rect 17911 19672 19340 19700
rect 17911 19669 17923 19672
rect 17865 19663 17923 19669
rect 19334 19660 19340 19672
rect 19392 19660 19398 19712
rect 19702 19660 19708 19712
rect 19760 19700 19766 19712
rect 20162 19700 20168 19712
rect 19760 19672 20168 19700
rect 19760 19660 19766 19672
rect 20162 19660 20168 19672
rect 20220 19660 20226 19712
rect 20806 19660 20812 19712
rect 20864 19700 20870 19712
rect 21085 19703 21143 19709
rect 21085 19700 21097 19703
rect 20864 19672 21097 19700
rect 20864 19660 20870 19672
rect 21085 19669 21097 19672
rect 21131 19700 21143 19703
rect 22186 19700 22192 19712
rect 21131 19672 22192 19700
rect 21131 19669 21143 19672
rect 21085 19663 21143 19669
rect 22186 19660 22192 19672
rect 22244 19660 22250 19712
rect 28994 19660 29000 19712
rect 29052 19700 29058 19712
rect 29730 19700 29736 19712
rect 29052 19672 29736 19700
rect 29052 19660 29058 19672
rect 29730 19660 29736 19672
rect 29788 19660 29794 19712
rect 1104 19610 39836 19632
rect 1104 19558 4246 19610
rect 4298 19558 4310 19610
rect 4362 19558 4374 19610
rect 4426 19558 4438 19610
rect 4490 19558 34966 19610
rect 35018 19558 35030 19610
rect 35082 19558 35094 19610
rect 35146 19558 35158 19610
rect 35210 19558 39836 19610
rect 1104 19536 39836 19558
rect 2038 19496 2044 19508
rect 1999 19468 2044 19496
rect 2038 19456 2044 19468
rect 2096 19456 2102 19508
rect 4341 19499 4399 19505
rect 4341 19465 4353 19499
rect 4387 19496 4399 19499
rect 4614 19496 4620 19508
rect 4387 19468 4620 19496
rect 4387 19465 4399 19468
rect 4341 19459 4399 19465
rect 4614 19456 4620 19468
rect 4672 19496 4678 19508
rect 4982 19496 4988 19508
rect 4672 19468 4988 19496
rect 4672 19456 4678 19468
rect 4982 19456 4988 19468
rect 5040 19456 5046 19508
rect 9861 19499 9919 19505
rect 9861 19465 9873 19499
rect 9907 19496 9919 19499
rect 10686 19496 10692 19508
rect 9907 19468 10692 19496
rect 9907 19465 9919 19468
rect 9861 19459 9919 19465
rect 10686 19456 10692 19468
rect 10744 19456 10750 19508
rect 14001 19499 14059 19505
rect 11532 19468 13952 19496
rect 3510 19360 3516 19372
rect 2700 19332 3516 19360
rect 1670 19292 1676 19304
rect 1631 19264 1676 19292
rect 1670 19252 1676 19264
rect 1728 19252 1734 19304
rect 1762 19252 1768 19304
rect 1820 19292 1826 19304
rect 1898 19295 1956 19301
rect 1820 19264 1865 19292
rect 1820 19252 1826 19264
rect 1898 19261 1910 19295
rect 1944 19292 1956 19295
rect 2700 19292 2728 19332
rect 3510 19320 3516 19332
rect 3568 19320 3574 19372
rect 10704 19360 10732 19456
rect 11532 19360 11560 19468
rect 12434 19428 12440 19440
rect 5736 19332 6040 19360
rect 1944 19264 2728 19292
rect 2777 19295 2835 19301
rect 1944 19261 1956 19264
rect 1898 19255 1956 19261
rect 2777 19261 2789 19295
rect 2823 19261 2835 19295
rect 3050 19292 3056 19304
rect 3011 19264 3056 19292
rect 2777 19255 2835 19261
rect 1394 19116 1400 19168
rect 1452 19156 1458 19168
rect 2792 19156 2820 19255
rect 3050 19252 3056 19264
rect 3108 19252 3114 19304
rect 3878 19252 3884 19304
rect 3936 19292 3942 19304
rect 5736 19292 5764 19332
rect 5902 19292 5908 19304
rect 3936 19264 5764 19292
rect 5863 19264 5908 19292
rect 3936 19252 3942 19264
rect 5902 19252 5908 19264
rect 5960 19252 5966 19304
rect 6012 19292 6040 19332
rect 7024 19332 7420 19360
rect 10704 19332 11560 19360
rect 7024 19292 7052 19332
rect 6012 19264 7052 19292
rect 7101 19295 7159 19301
rect 7101 19261 7113 19295
rect 7147 19292 7159 19295
rect 7190 19292 7196 19304
rect 7147 19264 7196 19292
rect 7147 19261 7159 19264
rect 7101 19255 7159 19261
rect 7190 19252 7196 19264
rect 7248 19252 7254 19304
rect 7285 19295 7343 19301
rect 7285 19261 7297 19295
rect 7331 19261 7343 19295
rect 7285 19255 7343 19261
rect 4798 19184 4804 19236
rect 4856 19224 4862 19236
rect 7300 19224 7328 19255
rect 4856 19196 7328 19224
rect 7392 19224 7420 19332
rect 8389 19295 8447 19301
rect 8389 19261 8401 19295
rect 8435 19292 8447 19295
rect 8570 19292 8576 19304
rect 8435 19264 8576 19292
rect 8435 19261 8447 19264
rect 8389 19255 8447 19261
rect 8570 19252 8576 19264
rect 8628 19252 8634 19304
rect 9030 19252 9036 19304
rect 9088 19292 9094 19304
rect 9677 19295 9735 19301
rect 9677 19292 9689 19295
rect 9088 19264 9689 19292
rect 9088 19252 9094 19264
rect 9677 19261 9689 19264
rect 9723 19261 9735 19295
rect 9677 19255 9735 19261
rect 10413 19295 10471 19301
rect 10413 19261 10425 19295
rect 10459 19292 10471 19295
rect 10505 19295 10563 19301
rect 10505 19292 10517 19295
rect 10459 19264 10517 19292
rect 10459 19261 10471 19264
rect 10413 19255 10471 19261
rect 10505 19261 10517 19264
rect 10551 19261 10563 19295
rect 10505 19255 10563 19261
rect 10597 19295 10655 19301
rect 10597 19261 10609 19295
rect 10643 19292 10655 19295
rect 11238 19292 11244 19304
rect 10643 19264 11244 19292
rect 10643 19261 10655 19264
rect 10597 19255 10655 19261
rect 11238 19252 11244 19264
rect 11296 19252 11302 19304
rect 11532 19301 11560 19332
rect 12360 19400 12440 19428
rect 11517 19295 11575 19301
rect 11517 19261 11529 19295
rect 11563 19261 11575 19295
rect 11517 19255 11575 19261
rect 11057 19227 11115 19233
rect 11057 19224 11069 19227
rect 7392 19196 11069 19224
rect 4856 19184 4862 19196
rect 6104 19165 6132 19196
rect 11057 19193 11069 19196
rect 11103 19193 11115 19227
rect 12360 19224 12388 19400
rect 12434 19388 12440 19400
rect 12492 19388 12498 19440
rect 13924 19428 13952 19468
rect 14001 19465 14013 19499
rect 14047 19496 14059 19499
rect 14182 19496 14188 19508
rect 14047 19468 14188 19496
rect 14047 19465 14059 19468
rect 14001 19459 14059 19465
rect 14182 19456 14188 19468
rect 14240 19456 14246 19508
rect 17034 19496 17040 19508
rect 16776 19468 17040 19496
rect 15194 19428 15200 19440
rect 13924 19400 15200 19428
rect 15194 19388 15200 19400
rect 15252 19388 15258 19440
rect 12636 19332 13124 19360
rect 12437 19295 12495 19301
rect 12437 19261 12449 19295
rect 12483 19292 12495 19295
rect 12636 19292 12664 19332
rect 12483 19264 12664 19292
rect 12713 19295 12771 19301
rect 12483 19261 12495 19264
rect 12437 19255 12495 19261
rect 12713 19261 12725 19295
rect 12759 19292 12771 19295
rect 12986 19292 12992 19304
rect 12759 19264 12992 19292
rect 12759 19261 12771 19264
rect 12713 19255 12771 19261
rect 12986 19252 12992 19264
rect 13044 19252 13050 19304
rect 13096 19292 13124 19332
rect 14734 19320 14740 19372
rect 14792 19360 14798 19372
rect 14918 19360 14924 19372
rect 14792 19332 14924 19360
rect 14792 19320 14798 19332
rect 14918 19320 14924 19332
rect 14976 19320 14982 19372
rect 15488 19332 16160 19360
rect 13814 19292 13820 19304
rect 13096 19264 13820 19292
rect 13814 19252 13820 19264
rect 13872 19252 13878 19304
rect 15010 19292 15016 19304
rect 14971 19264 15016 19292
rect 15010 19252 15016 19264
rect 15068 19252 15074 19304
rect 15105 19295 15163 19301
rect 15105 19261 15117 19295
rect 15151 19292 15163 19295
rect 15286 19292 15292 19304
rect 15151 19264 15292 19292
rect 15151 19261 15163 19264
rect 15105 19255 15163 19261
rect 15286 19252 15292 19264
rect 15344 19252 15350 19304
rect 11057 19187 11115 19193
rect 11164 19196 12388 19224
rect 1452 19128 2820 19156
rect 6089 19159 6147 19165
rect 1452 19116 1458 19128
rect 6089 19125 6101 19159
rect 6135 19125 6147 19159
rect 6914 19156 6920 19168
rect 6875 19128 6920 19156
rect 6089 19119 6147 19125
rect 6914 19116 6920 19128
rect 6972 19116 6978 19168
rect 8573 19159 8631 19165
rect 8573 19125 8585 19159
rect 8619 19156 8631 19159
rect 9858 19156 9864 19168
rect 8619 19128 9864 19156
rect 8619 19125 8631 19128
rect 8573 19119 8631 19125
rect 9858 19116 9864 19128
rect 9916 19116 9922 19168
rect 10413 19159 10471 19165
rect 10413 19125 10425 19159
rect 10459 19156 10471 19159
rect 11164 19156 11192 19196
rect 13538 19184 13544 19236
rect 13596 19224 13602 19236
rect 15488 19224 15516 19332
rect 15565 19295 15623 19301
rect 15565 19261 15577 19295
rect 15611 19292 15623 19295
rect 15930 19292 15936 19304
rect 15611 19264 15936 19292
rect 15611 19261 15623 19264
rect 15565 19255 15623 19261
rect 15930 19252 15936 19264
rect 15988 19252 15994 19304
rect 13596 19196 15516 19224
rect 16025 19227 16083 19233
rect 13596 19184 13602 19196
rect 16025 19193 16037 19227
rect 16071 19193 16083 19227
rect 16132 19224 16160 19332
rect 16206 19252 16212 19304
rect 16264 19292 16270 19304
rect 16776 19301 16804 19468
rect 17034 19456 17040 19468
rect 17092 19496 17098 19508
rect 18506 19496 18512 19508
rect 17092 19468 18512 19496
rect 17092 19456 17098 19468
rect 18506 19456 18512 19468
rect 18564 19456 18570 19508
rect 19150 19456 19156 19508
rect 19208 19496 19214 19508
rect 20714 19496 20720 19508
rect 19208 19468 20720 19496
rect 19208 19456 19214 19468
rect 20714 19456 20720 19468
rect 20772 19456 20778 19508
rect 29546 19456 29552 19508
rect 29604 19496 29610 19508
rect 31297 19499 31355 19505
rect 31297 19496 31309 19499
rect 29604 19468 31309 19496
rect 29604 19456 29610 19468
rect 31297 19465 31309 19468
rect 31343 19496 31355 19499
rect 32214 19496 32220 19508
rect 31343 19468 32220 19496
rect 31343 19465 31355 19468
rect 31297 19459 31355 19465
rect 32214 19456 32220 19468
rect 32272 19456 32278 19508
rect 34238 19496 34244 19508
rect 34199 19468 34244 19496
rect 34238 19456 34244 19468
rect 34296 19456 34302 19508
rect 35069 19499 35127 19505
rect 35069 19465 35081 19499
rect 35115 19496 35127 19499
rect 35250 19496 35256 19508
rect 35115 19468 35256 19496
rect 35115 19465 35127 19468
rect 35069 19459 35127 19465
rect 16942 19428 16948 19440
rect 16855 19400 16948 19428
rect 16942 19388 16948 19400
rect 17000 19428 17006 19440
rect 19610 19428 19616 19440
rect 17000 19400 19616 19428
rect 17000 19388 17006 19400
rect 19610 19388 19616 19400
rect 19668 19428 19674 19440
rect 20438 19428 20444 19440
rect 19668 19400 20444 19428
rect 19668 19388 19674 19400
rect 20438 19388 20444 19400
rect 20496 19388 20502 19440
rect 21082 19388 21088 19440
rect 21140 19428 21146 19440
rect 21726 19428 21732 19440
rect 21140 19400 21732 19428
rect 21140 19388 21146 19400
rect 21726 19388 21732 19400
rect 21784 19388 21790 19440
rect 22186 19388 22192 19440
rect 22244 19428 22250 19440
rect 32490 19428 32496 19440
rect 22244 19400 32496 19428
rect 22244 19388 22250 19400
rect 32490 19388 32496 19400
rect 32548 19388 32554 19440
rect 35084 19428 35112 19459
rect 35250 19456 35256 19468
rect 35308 19456 35314 19508
rect 34532 19400 35112 19428
rect 16960 19301 16988 19388
rect 19334 19320 19340 19372
rect 19392 19360 19398 19372
rect 23382 19360 23388 19372
rect 19392 19332 23388 19360
rect 19392 19320 19398 19332
rect 16485 19295 16543 19301
rect 16485 19292 16497 19295
rect 16264 19264 16497 19292
rect 16264 19252 16270 19264
rect 16485 19261 16497 19264
rect 16531 19261 16543 19295
rect 16485 19255 16543 19261
rect 16761 19295 16819 19301
rect 16761 19261 16773 19295
rect 16807 19261 16819 19295
rect 16761 19255 16819 19261
rect 16945 19295 17003 19301
rect 16945 19261 16957 19295
rect 16991 19261 17003 19295
rect 16945 19255 17003 19261
rect 17129 19295 17187 19301
rect 17129 19261 17141 19295
rect 17175 19292 17187 19295
rect 17218 19292 17224 19304
rect 17175 19264 17224 19292
rect 17175 19261 17187 19264
rect 17129 19255 17187 19261
rect 17218 19252 17224 19264
rect 17276 19252 17282 19304
rect 17405 19295 17463 19301
rect 17405 19261 17417 19295
rect 17451 19292 17463 19295
rect 17494 19292 17500 19304
rect 17451 19264 17500 19292
rect 17451 19261 17463 19264
rect 17405 19255 17463 19261
rect 17494 19252 17500 19264
rect 17552 19252 17558 19304
rect 17678 19252 17684 19304
rect 17736 19292 17742 19304
rect 18049 19295 18107 19301
rect 18049 19292 18061 19295
rect 17736 19264 18061 19292
rect 17736 19252 17742 19264
rect 18049 19261 18061 19264
rect 18095 19261 18107 19295
rect 18049 19255 18107 19261
rect 18601 19295 18659 19301
rect 18601 19261 18613 19295
rect 18647 19292 18659 19295
rect 18782 19292 18788 19304
rect 18647 19264 18788 19292
rect 18647 19261 18659 19264
rect 18601 19255 18659 19261
rect 18782 19252 18788 19264
rect 18840 19252 18846 19304
rect 19444 19301 19472 19332
rect 23382 19320 23388 19332
rect 23440 19320 23446 19372
rect 25866 19360 25872 19372
rect 25827 19332 25872 19360
rect 25866 19320 25872 19332
rect 25924 19320 25930 19372
rect 28184 19332 28580 19360
rect 19429 19295 19487 19301
rect 19429 19261 19441 19295
rect 19475 19261 19487 19295
rect 19610 19292 19616 19304
rect 19571 19264 19616 19292
rect 19429 19255 19487 19261
rect 19610 19252 19616 19264
rect 19668 19252 19674 19304
rect 19702 19252 19708 19304
rect 19760 19292 19766 19304
rect 19760 19264 19805 19292
rect 19760 19252 19766 19264
rect 19978 19252 19984 19304
rect 20036 19292 20042 19304
rect 20257 19295 20315 19301
rect 20036 19264 20081 19292
rect 20036 19252 20042 19264
rect 20257 19261 20269 19295
rect 20303 19292 20315 19295
rect 20346 19292 20352 19304
rect 20303 19264 20352 19292
rect 20303 19261 20315 19264
rect 20257 19255 20315 19261
rect 20346 19252 20352 19264
rect 20404 19252 20410 19304
rect 20625 19295 20683 19301
rect 20625 19261 20637 19295
rect 20671 19292 20683 19295
rect 20898 19292 20904 19304
rect 20671 19264 20904 19292
rect 20671 19261 20683 19264
rect 20625 19255 20683 19261
rect 20898 19252 20904 19264
rect 20956 19252 20962 19304
rect 21177 19295 21235 19301
rect 21177 19261 21189 19295
rect 21223 19292 21235 19295
rect 21266 19292 21272 19304
rect 21223 19264 21272 19292
rect 21223 19261 21235 19264
rect 21177 19255 21235 19261
rect 21266 19252 21272 19264
rect 21324 19252 21330 19304
rect 21453 19295 21511 19301
rect 21453 19261 21465 19295
rect 21499 19292 21511 19295
rect 21818 19292 21824 19304
rect 21499 19264 21824 19292
rect 21499 19261 21511 19264
rect 21453 19255 21511 19261
rect 21818 19252 21824 19264
rect 21876 19252 21882 19304
rect 22094 19252 22100 19304
rect 22152 19292 22158 19304
rect 22281 19295 22339 19301
rect 22281 19292 22293 19295
rect 22152 19264 22293 19292
rect 22152 19252 22158 19264
rect 22281 19261 22293 19264
rect 22327 19261 22339 19295
rect 22281 19255 22339 19261
rect 22465 19295 22523 19301
rect 22465 19261 22477 19295
rect 22511 19261 22523 19295
rect 22830 19292 22836 19304
rect 22791 19264 22836 19292
rect 22465 19255 22523 19261
rect 18877 19227 18935 19233
rect 16132 19196 18276 19224
rect 16025 19187 16083 19193
rect 11698 19156 11704 19168
rect 10459 19128 11192 19156
rect 11659 19128 11704 19156
rect 10459 19125 10471 19128
rect 10413 19119 10471 19125
rect 11698 19116 11704 19128
rect 11756 19116 11762 19168
rect 14550 19116 14556 19168
rect 14608 19156 14614 19168
rect 15838 19156 15844 19168
rect 14608 19128 15844 19156
rect 14608 19116 14614 19128
rect 15838 19116 15844 19128
rect 15896 19116 15902 19168
rect 16040 19156 16068 19187
rect 16850 19156 16856 19168
rect 16040 19128 16856 19156
rect 16850 19116 16856 19128
rect 16908 19116 16914 19168
rect 16942 19116 16948 19168
rect 17000 19156 17006 19168
rect 18141 19159 18199 19165
rect 18141 19156 18153 19159
rect 17000 19128 18153 19156
rect 17000 19116 17006 19128
rect 18141 19125 18153 19128
rect 18187 19125 18199 19159
rect 18248 19156 18276 19196
rect 18877 19193 18889 19227
rect 18923 19224 18935 19227
rect 22480 19224 22508 19255
rect 22830 19252 22836 19264
rect 22888 19252 22894 19304
rect 22922 19252 22928 19304
rect 22980 19292 22986 19304
rect 23658 19292 23664 19304
rect 22980 19264 23025 19292
rect 23619 19264 23664 19292
rect 22980 19252 22986 19264
rect 23658 19252 23664 19264
rect 23716 19252 23722 19304
rect 24026 19252 24032 19304
rect 24084 19292 24090 19304
rect 24213 19295 24271 19301
rect 24213 19292 24225 19295
rect 24084 19264 24225 19292
rect 24084 19252 24090 19264
rect 24213 19261 24225 19264
rect 24259 19261 24271 19295
rect 24670 19292 24676 19304
rect 24631 19264 24676 19292
rect 24213 19255 24271 19261
rect 24670 19252 24676 19264
rect 24728 19252 24734 19304
rect 26053 19295 26111 19301
rect 26053 19261 26065 19295
rect 26099 19292 26111 19295
rect 26513 19295 26571 19301
rect 26099 19264 26464 19292
rect 26099 19261 26111 19264
rect 26053 19255 26111 19261
rect 24118 19224 24124 19236
rect 18923 19196 22416 19224
rect 22480 19196 24124 19224
rect 18923 19193 18935 19196
rect 18877 19187 18935 19193
rect 20533 19159 20591 19165
rect 20533 19156 20545 19159
rect 18248 19128 20545 19156
rect 18141 19119 18199 19125
rect 20533 19125 20545 19128
rect 20579 19125 20591 19159
rect 22388 19156 22416 19196
rect 24118 19184 24124 19196
rect 24176 19184 24182 19236
rect 23474 19156 23480 19168
rect 22388 19128 23480 19156
rect 20533 19119 20591 19125
rect 23474 19116 23480 19128
rect 23532 19116 23538 19168
rect 23566 19116 23572 19168
rect 23624 19156 23630 19168
rect 23753 19159 23811 19165
rect 23753 19156 23765 19159
rect 23624 19128 23765 19156
rect 23624 19116 23630 19128
rect 23753 19125 23765 19128
rect 23799 19125 23811 19159
rect 26436 19156 26464 19264
rect 26513 19261 26525 19295
rect 26559 19261 26571 19295
rect 26513 19255 26571 19261
rect 26528 19224 26556 19255
rect 26602 19252 26608 19304
rect 26660 19292 26666 19304
rect 27249 19295 27307 19301
rect 26660 19264 26705 19292
rect 26660 19252 26666 19264
rect 27249 19261 27261 19295
rect 27295 19292 27307 19295
rect 27706 19292 27712 19304
rect 27295 19264 27712 19292
rect 27295 19261 27307 19264
rect 27249 19255 27307 19261
rect 27706 19252 27712 19264
rect 27764 19252 27770 19304
rect 27154 19224 27160 19236
rect 26528 19196 27160 19224
rect 27154 19184 27160 19196
rect 27212 19184 27218 19236
rect 26786 19156 26792 19168
rect 26436 19128 26792 19156
rect 23753 19119 23811 19125
rect 26786 19116 26792 19128
rect 26844 19116 26850 19168
rect 27062 19116 27068 19168
rect 27120 19156 27126 19168
rect 28184 19156 28212 19332
rect 28261 19295 28319 19301
rect 28261 19261 28273 19295
rect 28307 19261 28319 19295
rect 28442 19292 28448 19304
rect 28403 19264 28448 19292
rect 28261 19255 28319 19261
rect 27120 19128 28212 19156
rect 28276 19156 28304 19255
rect 28442 19252 28448 19264
rect 28500 19252 28506 19304
rect 28552 19292 28580 19332
rect 29730 19320 29736 19372
rect 29788 19360 29794 19372
rect 30193 19363 30251 19369
rect 30193 19360 30205 19363
rect 29788 19332 30205 19360
rect 29788 19320 29794 19332
rect 30193 19329 30205 19332
rect 30239 19329 30251 19363
rect 30193 19323 30251 19329
rect 30742 19320 30748 19372
rect 30800 19360 30806 19372
rect 32858 19360 32864 19372
rect 30800 19332 31708 19360
rect 30800 19320 30806 19332
rect 31680 19304 31708 19332
rect 31864 19332 32864 19360
rect 29086 19292 29092 19304
rect 28552 19264 29092 19292
rect 29086 19252 29092 19264
rect 29144 19252 29150 19304
rect 29457 19295 29515 19301
rect 29457 19261 29469 19295
rect 29503 19261 29515 19295
rect 29638 19292 29644 19304
rect 29599 19264 29644 19292
rect 29457 19255 29515 19261
rect 28721 19227 28779 19233
rect 28721 19193 28733 19227
rect 28767 19224 28779 19227
rect 29362 19224 29368 19236
rect 28767 19196 29368 19224
rect 28767 19193 28779 19196
rect 28721 19187 28779 19193
rect 29362 19184 29368 19196
rect 29420 19184 29426 19236
rect 29472 19224 29500 19255
rect 29638 19252 29644 19264
rect 29696 19252 29702 19304
rect 30098 19292 30104 19304
rect 30059 19264 30104 19292
rect 30098 19252 30104 19264
rect 30156 19252 30162 19304
rect 31386 19292 31392 19304
rect 31347 19264 31392 19292
rect 31386 19252 31392 19264
rect 31444 19252 31450 19304
rect 31573 19295 31631 19301
rect 31573 19261 31585 19295
rect 31619 19261 31631 19295
rect 31573 19255 31631 19261
rect 30650 19224 30656 19236
rect 29472 19196 30656 19224
rect 30650 19184 30656 19196
rect 30708 19184 30714 19236
rect 31294 19184 31300 19236
rect 31352 19224 31358 19236
rect 31588 19224 31616 19255
rect 31662 19252 31668 19304
rect 31720 19252 31726 19304
rect 31864 19224 31892 19332
rect 32858 19320 32864 19332
rect 32916 19320 32922 19372
rect 34532 19360 34560 19400
rect 34072 19332 34560 19360
rect 32214 19292 32220 19304
rect 32175 19264 32220 19292
rect 32214 19252 32220 19264
rect 32272 19252 32278 19304
rect 33134 19292 33140 19304
rect 33095 19264 33140 19292
rect 33134 19252 33140 19264
rect 33192 19252 33198 19304
rect 33318 19292 33324 19304
rect 33279 19264 33324 19292
rect 33318 19252 33324 19264
rect 33376 19252 33382 19304
rect 33689 19295 33747 19301
rect 33689 19261 33701 19295
rect 33735 19292 33747 19295
rect 33962 19292 33968 19304
rect 33735 19264 33968 19292
rect 33735 19261 33747 19264
rect 33689 19255 33747 19261
rect 33962 19252 33968 19264
rect 34020 19292 34026 19304
rect 34072 19292 34100 19332
rect 34790 19320 34796 19372
rect 34848 19360 34854 19372
rect 34848 19332 35664 19360
rect 34848 19320 34854 19332
rect 34020 19264 34100 19292
rect 34020 19252 34026 19264
rect 34146 19252 34152 19304
rect 34204 19292 34210 19304
rect 35636 19301 35664 19332
rect 36446 19320 36452 19372
rect 36504 19360 36510 19372
rect 36504 19332 36860 19360
rect 36504 19320 36510 19332
rect 34885 19295 34943 19301
rect 34885 19292 34897 19295
rect 34204 19264 34897 19292
rect 34204 19252 34210 19264
rect 34885 19261 34897 19264
rect 34931 19261 34943 19295
rect 34885 19255 34943 19261
rect 35621 19295 35679 19301
rect 35621 19261 35633 19295
rect 35667 19261 35679 19295
rect 36354 19292 36360 19304
rect 36315 19264 36360 19292
rect 35621 19255 35679 19261
rect 36354 19252 36360 19264
rect 36412 19252 36418 19304
rect 36722 19292 36728 19304
rect 36683 19264 36728 19292
rect 36722 19252 36728 19264
rect 36780 19252 36786 19304
rect 36832 19292 36860 19332
rect 36906 19292 36912 19304
rect 36832 19264 36912 19292
rect 36906 19252 36912 19264
rect 36964 19292 36970 19304
rect 37461 19295 37519 19301
rect 37461 19292 37473 19295
rect 36964 19264 37473 19292
rect 36964 19252 36970 19264
rect 37461 19261 37473 19264
rect 37507 19261 37519 19295
rect 37737 19295 37795 19301
rect 37737 19292 37749 19295
rect 37461 19255 37519 19261
rect 37568 19264 37749 19292
rect 31352 19196 31892 19224
rect 37001 19227 37059 19233
rect 31352 19184 31358 19196
rect 37001 19193 37013 19227
rect 37047 19224 37059 19227
rect 37568 19224 37596 19264
rect 37737 19261 37749 19264
rect 37783 19261 37795 19295
rect 37737 19255 37795 19261
rect 37047 19196 37596 19224
rect 37047 19193 37059 19196
rect 37001 19187 37059 19193
rect 30374 19156 30380 19168
rect 28276 19128 30380 19156
rect 27120 19116 27126 19128
rect 30374 19116 30380 19128
rect 30432 19116 30438 19168
rect 32122 19116 32128 19168
rect 32180 19156 32186 19168
rect 34514 19156 34520 19168
rect 32180 19128 34520 19156
rect 32180 19116 32186 19128
rect 34514 19116 34520 19128
rect 34572 19116 34578 19168
rect 35713 19159 35771 19165
rect 35713 19125 35725 19159
rect 35759 19156 35771 19159
rect 36538 19156 36544 19168
rect 35759 19128 36544 19156
rect 35759 19125 35771 19128
rect 35713 19119 35771 19125
rect 36538 19116 36544 19128
rect 36596 19116 36602 19168
rect 36722 19116 36728 19168
rect 36780 19156 36786 19168
rect 38841 19159 38899 19165
rect 38841 19156 38853 19159
rect 36780 19128 38853 19156
rect 36780 19116 36786 19128
rect 38841 19125 38853 19128
rect 38887 19125 38899 19159
rect 38841 19119 38899 19125
rect 1104 19066 39836 19088
rect 1104 19014 19606 19066
rect 19658 19014 19670 19066
rect 19722 19014 19734 19066
rect 19786 19014 19798 19066
rect 19850 19014 39836 19066
rect 1104 18992 39836 19014
rect 2774 18912 2780 18964
rect 2832 18952 2838 18964
rect 4154 18952 4160 18964
rect 2832 18924 2877 18952
rect 4115 18924 4160 18952
rect 2832 18912 2838 18924
rect 4154 18912 4160 18924
rect 4212 18912 4218 18964
rect 5994 18912 6000 18964
rect 6052 18952 6058 18964
rect 9030 18952 9036 18964
rect 6052 18924 8892 18952
rect 8991 18924 9036 18952
rect 6052 18912 6058 18924
rect 8864 18884 8892 18924
rect 9030 18912 9036 18924
rect 9088 18912 9094 18964
rect 14366 18952 14372 18964
rect 9232 18924 14372 18952
rect 9232 18884 9260 18924
rect 14366 18912 14372 18924
rect 14424 18912 14430 18964
rect 14476 18924 17080 18952
rect 8864 18856 9260 18884
rect 1394 18816 1400 18828
rect 1355 18788 1400 18816
rect 1394 18776 1400 18788
rect 1452 18776 1458 18828
rect 3510 18776 3516 18828
rect 3568 18816 3574 18828
rect 4065 18819 4123 18825
rect 4065 18816 4077 18819
rect 3568 18788 4077 18816
rect 3568 18776 3574 18788
rect 4065 18785 4077 18788
rect 4111 18785 4123 18819
rect 5166 18816 5172 18828
rect 5127 18788 5172 18816
rect 4065 18779 4123 18785
rect 5166 18776 5172 18788
rect 5224 18776 5230 18828
rect 6270 18816 6276 18828
rect 6231 18788 6276 18816
rect 6270 18776 6276 18788
rect 6328 18776 6334 18828
rect 6822 18816 6828 18828
rect 6783 18788 6828 18816
rect 6822 18776 6828 18788
rect 6880 18776 6886 18828
rect 7098 18816 7104 18828
rect 7059 18788 7104 18816
rect 7098 18776 7104 18788
rect 7156 18776 7162 18828
rect 8941 18819 8999 18825
rect 8941 18816 8953 18819
rect 8220 18788 8953 18816
rect 1673 18751 1731 18757
rect 1673 18717 1685 18751
rect 1719 18748 1731 18751
rect 5074 18748 5080 18760
rect 1719 18720 2728 18748
rect 5035 18720 5080 18748
rect 1719 18717 1731 18720
rect 1673 18711 1731 18717
rect 2700 18680 2728 18720
rect 5074 18708 5080 18720
rect 5132 18708 5138 18760
rect 6089 18683 6147 18689
rect 2700 18652 5396 18680
rect 5368 18621 5396 18652
rect 6089 18649 6101 18683
rect 6135 18680 6147 18683
rect 6840 18680 6868 18776
rect 6135 18652 6868 18680
rect 6135 18649 6147 18652
rect 6089 18643 6147 18649
rect 5353 18615 5411 18621
rect 5353 18581 5365 18615
rect 5399 18581 5411 18615
rect 5353 18575 5411 18581
rect 7926 18572 7932 18624
rect 7984 18612 7990 18624
rect 8220 18621 8248 18788
rect 8941 18785 8953 18788
rect 8987 18785 8999 18819
rect 8941 18779 8999 18785
rect 9677 18819 9735 18825
rect 9677 18785 9689 18819
rect 9723 18816 9735 18819
rect 14476 18816 14504 18924
rect 15378 18844 15384 18896
rect 15436 18844 15442 18896
rect 9723 18788 14504 18816
rect 9723 18785 9735 18788
rect 9677 18779 9735 18785
rect 14550 18776 14556 18828
rect 14608 18816 14614 18828
rect 15396 18816 15424 18844
rect 15565 18819 15623 18825
rect 15565 18816 15577 18819
rect 14608 18788 14653 18816
rect 15396 18788 15577 18816
rect 14608 18776 14614 18788
rect 15565 18785 15577 18788
rect 15611 18785 15623 18819
rect 15565 18779 15623 18785
rect 15838 18776 15844 18828
rect 15896 18816 15902 18828
rect 16942 18816 16948 18828
rect 15896 18788 16948 18816
rect 15896 18776 15902 18788
rect 16942 18776 16948 18788
rect 17000 18776 17006 18828
rect 10226 18708 10232 18760
rect 10284 18748 10290 18760
rect 10321 18751 10379 18757
rect 10321 18748 10333 18751
rect 10284 18720 10333 18748
rect 10284 18708 10290 18720
rect 10321 18717 10333 18720
rect 10367 18717 10379 18751
rect 10594 18748 10600 18760
rect 10555 18720 10600 18748
rect 10321 18711 10379 18717
rect 10594 18708 10600 18720
rect 10652 18708 10658 18760
rect 12434 18748 12440 18760
rect 12395 18720 12440 18748
rect 12434 18708 12440 18720
rect 12492 18708 12498 18760
rect 12713 18751 12771 18757
rect 12713 18717 12725 18751
rect 12759 18748 12771 18751
rect 13538 18748 13544 18760
rect 12759 18720 13544 18748
rect 12759 18717 12771 18720
rect 12713 18711 12771 18717
rect 13538 18708 13544 18720
rect 13596 18708 13602 18760
rect 15289 18751 15347 18757
rect 15289 18717 15301 18751
rect 15335 18748 15347 18751
rect 16758 18748 16764 18760
rect 15335 18720 16764 18748
rect 15335 18717 15347 18720
rect 15289 18711 15347 18717
rect 16758 18708 16764 18720
rect 16816 18708 16822 18760
rect 17052 18748 17080 18924
rect 19058 18912 19064 18964
rect 19116 18952 19122 18964
rect 19797 18955 19855 18961
rect 19797 18952 19809 18955
rect 19116 18924 19809 18952
rect 19116 18912 19122 18924
rect 19797 18921 19809 18924
rect 19843 18921 19855 18955
rect 19797 18915 19855 18921
rect 19889 18955 19947 18961
rect 19889 18921 19901 18955
rect 19935 18952 19947 18955
rect 20070 18952 20076 18964
rect 19935 18924 20076 18952
rect 19935 18921 19947 18924
rect 19889 18915 19947 18921
rect 20070 18912 20076 18924
rect 20128 18912 20134 18964
rect 20993 18955 21051 18961
rect 20993 18921 21005 18955
rect 21039 18952 21051 18955
rect 21174 18952 21180 18964
rect 21039 18924 21180 18952
rect 21039 18921 21051 18924
rect 20993 18915 21051 18921
rect 21174 18912 21180 18924
rect 21232 18912 21238 18964
rect 21450 18912 21456 18964
rect 21508 18952 21514 18964
rect 21508 18924 30328 18952
rect 21508 18912 21514 18924
rect 19518 18884 19524 18896
rect 19076 18856 19524 18884
rect 17310 18776 17316 18828
rect 17368 18816 17374 18828
rect 17681 18819 17739 18825
rect 17681 18816 17693 18819
rect 17368 18788 17693 18816
rect 17368 18776 17374 18788
rect 17681 18785 17693 18788
rect 17727 18785 17739 18819
rect 18414 18816 18420 18828
rect 18375 18788 18420 18816
rect 17681 18779 17739 18785
rect 18414 18776 18420 18788
rect 18472 18776 18478 18828
rect 18693 18819 18751 18825
rect 18693 18785 18705 18819
rect 18739 18816 18751 18819
rect 18782 18816 18788 18828
rect 18739 18788 18788 18816
rect 18739 18785 18751 18788
rect 18693 18779 18751 18785
rect 18782 18776 18788 18788
rect 18840 18776 18846 18828
rect 19076 18825 19104 18856
rect 19518 18844 19524 18856
rect 19576 18844 19582 18896
rect 19610 18844 19616 18896
rect 19668 18884 19674 18896
rect 19981 18887 20039 18893
rect 19981 18884 19993 18887
rect 19668 18856 19713 18884
rect 19904 18856 19993 18884
rect 19668 18844 19674 18856
rect 19061 18819 19119 18825
rect 19061 18785 19073 18819
rect 19107 18785 19119 18819
rect 19061 18779 19119 18785
rect 19245 18819 19303 18825
rect 19245 18785 19257 18819
rect 19291 18816 19303 18819
rect 19904 18816 19932 18856
rect 19981 18853 19993 18856
rect 20027 18884 20039 18887
rect 20162 18884 20168 18896
rect 20027 18856 20168 18884
rect 20027 18853 20039 18856
rect 19981 18847 20039 18853
rect 20162 18844 20168 18856
rect 20220 18844 20226 18896
rect 21358 18884 21364 18896
rect 21100 18856 21364 18884
rect 21100 18825 21128 18856
rect 21358 18844 21364 18856
rect 21416 18884 21422 18896
rect 22002 18884 22008 18896
rect 21416 18856 22008 18884
rect 21416 18844 21422 18856
rect 22002 18844 22008 18856
rect 22060 18844 22066 18896
rect 22830 18844 22836 18896
rect 22888 18884 22894 18896
rect 25130 18884 25136 18896
rect 22888 18856 25136 18884
rect 22888 18844 22894 18856
rect 25130 18844 25136 18856
rect 25188 18884 25194 18896
rect 25188 18856 28948 18884
rect 25188 18844 25194 18856
rect 19291 18788 19932 18816
rect 21085 18819 21143 18825
rect 19291 18785 19303 18788
rect 19245 18779 19303 18785
rect 21085 18785 21097 18819
rect 21131 18785 21143 18819
rect 21085 18779 21143 18785
rect 21266 18776 21272 18828
rect 21324 18816 21330 18828
rect 21453 18819 21511 18825
rect 21453 18816 21465 18819
rect 21324 18788 21465 18816
rect 21324 18776 21330 18788
rect 21453 18785 21465 18788
rect 21499 18785 21511 18819
rect 21910 18816 21916 18828
rect 21871 18788 21916 18816
rect 21453 18779 21511 18785
rect 20349 18751 20407 18757
rect 20349 18748 20361 18751
rect 17052 18720 20361 18748
rect 20349 18717 20361 18720
rect 20395 18717 20407 18751
rect 21468 18748 21496 18779
rect 21910 18776 21916 18788
rect 21968 18776 21974 18828
rect 22462 18816 22468 18828
rect 22423 18788 22468 18816
rect 22462 18776 22468 18788
rect 22520 18776 22526 18828
rect 23661 18819 23719 18825
rect 23661 18785 23673 18819
rect 23707 18785 23719 18819
rect 24026 18816 24032 18828
rect 23987 18788 24032 18816
rect 23661 18779 23719 18785
rect 21818 18748 21824 18760
rect 21468 18720 21824 18748
rect 20349 18711 20407 18717
rect 21818 18708 21824 18720
rect 21876 18708 21882 18760
rect 23676 18748 23704 18779
rect 24026 18776 24032 18788
rect 24084 18776 24090 18828
rect 25041 18819 25099 18825
rect 25041 18785 25053 18819
rect 25087 18816 25099 18819
rect 25498 18816 25504 18828
rect 25087 18788 25504 18816
rect 25087 18785 25099 18788
rect 25041 18779 25099 18785
rect 25498 18776 25504 18788
rect 25556 18776 25562 18828
rect 25682 18816 25688 18828
rect 25643 18788 25688 18816
rect 25682 18776 25688 18788
rect 25740 18776 25746 18828
rect 26786 18816 26792 18828
rect 26747 18788 26792 18816
rect 26786 18776 26792 18788
rect 26844 18776 26850 18828
rect 26970 18816 26976 18828
rect 26896 18788 26976 18816
rect 24489 18751 24547 18757
rect 23676 18720 23980 18748
rect 11974 18680 11980 18692
rect 11256 18652 11980 18680
rect 8205 18615 8263 18621
rect 8205 18612 8217 18615
rect 7984 18584 8217 18612
rect 7984 18572 7990 18584
rect 8205 18581 8217 18584
rect 8251 18581 8263 18615
rect 8205 18575 8263 18581
rect 9769 18615 9827 18621
rect 9769 18581 9781 18615
rect 9815 18612 9827 18615
rect 11256 18612 11284 18652
rect 11974 18640 11980 18652
rect 12032 18640 12038 18692
rect 14645 18683 14703 18689
rect 14645 18680 14657 18683
rect 13372 18652 14657 18680
rect 11882 18612 11888 18624
rect 9815 18584 11284 18612
rect 11843 18584 11888 18612
rect 9815 18581 9827 18584
rect 9769 18575 9827 18581
rect 11882 18572 11888 18584
rect 11940 18572 11946 18624
rect 12618 18572 12624 18624
rect 12676 18612 12682 18624
rect 13372 18612 13400 18652
rect 14645 18649 14657 18652
rect 14691 18649 14703 18683
rect 14645 18643 14703 18649
rect 16853 18683 16911 18689
rect 16853 18649 16865 18683
rect 16899 18680 16911 18683
rect 17494 18680 17500 18692
rect 16899 18652 17500 18680
rect 16899 18649 16911 18652
rect 16853 18643 16911 18649
rect 17494 18640 17500 18652
rect 17552 18640 17558 18692
rect 18966 18640 18972 18692
rect 19024 18680 19030 18692
rect 19061 18683 19119 18689
rect 19061 18680 19073 18683
rect 19024 18652 19073 18680
rect 19024 18640 19030 18652
rect 19061 18649 19073 18652
rect 19107 18649 19119 18683
rect 23753 18683 23811 18689
rect 19061 18643 19119 18649
rect 19168 18652 23612 18680
rect 12676 18584 13400 18612
rect 12676 18572 12682 18584
rect 13722 18572 13728 18624
rect 13780 18612 13786 18624
rect 13817 18615 13875 18621
rect 13817 18612 13829 18615
rect 13780 18584 13829 18612
rect 13780 18572 13786 18584
rect 13817 18581 13829 18584
rect 13863 18581 13875 18615
rect 13817 18575 13875 18581
rect 14366 18572 14372 18624
rect 14424 18612 14430 18624
rect 19168 18612 19196 18652
rect 14424 18584 19196 18612
rect 19429 18615 19487 18621
rect 14424 18572 14430 18584
rect 19429 18581 19441 18615
rect 19475 18612 19487 18615
rect 20346 18612 20352 18624
rect 19475 18584 20352 18612
rect 19475 18581 19487 18584
rect 19429 18575 19487 18581
rect 20346 18572 20352 18584
rect 20404 18572 20410 18624
rect 20530 18572 20536 18624
rect 20588 18612 20594 18624
rect 21174 18612 21180 18624
rect 20588 18584 21180 18612
rect 20588 18572 20594 18584
rect 21174 18572 21180 18584
rect 21232 18572 21238 18624
rect 22370 18572 22376 18624
rect 22428 18612 22434 18624
rect 22649 18615 22707 18621
rect 22649 18612 22661 18615
rect 22428 18584 22661 18612
rect 22428 18572 22434 18584
rect 22649 18581 22661 18584
rect 22695 18581 22707 18615
rect 23584 18612 23612 18652
rect 23753 18649 23765 18683
rect 23799 18680 23811 18683
rect 23842 18680 23848 18692
rect 23799 18652 23848 18680
rect 23799 18649 23811 18652
rect 23753 18643 23811 18649
rect 23842 18640 23848 18652
rect 23900 18640 23906 18692
rect 23952 18680 23980 18720
rect 24489 18717 24501 18751
rect 24535 18748 24547 18751
rect 24670 18748 24676 18760
rect 24535 18720 24676 18748
rect 24535 18717 24547 18720
rect 24489 18711 24547 18717
rect 24670 18708 24676 18720
rect 24728 18748 24734 18760
rect 26234 18748 26240 18760
rect 24728 18720 26240 18748
rect 24728 18708 24734 18720
rect 26234 18708 26240 18720
rect 26292 18708 26298 18760
rect 26896 18757 26924 18788
rect 26970 18776 26976 18788
rect 27028 18776 27034 18828
rect 27154 18816 27160 18828
rect 27115 18788 27160 18816
rect 27154 18776 27160 18788
rect 27212 18776 27218 18828
rect 27430 18816 27436 18828
rect 27391 18788 27436 18816
rect 27430 18776 27436 18788
rect 27488 18776 27494 18828
rect 27706 18816 27712 18828
rect 27667 18788 27712 18816
rect 27706 18776 27712 18788
rect 27764 18776 27770 18828
rect 28460 18825 28488 18856
rect 28445 18819 28503 18825
rect 28445 18785 28457 18819
rect 28491 18785 28503 18819
rect 28920 18816 28948 18856
rect 29362 18816 29368 18828
rect 28920 18788 29224 18816
rect 29323 18788 29368 18816
rect 28445 18779 28503 18785
rect 26881 18751 26939 18757
rect 26881 18717 26893 18751
rect 26927 18717 26939 18751
rect 29086 18748 29092 18760
rect 29047 18720 29092 18748
rect 26881 18711 26939 18717
rect 29086 18708 29092 18720
rect 29144 18708 29150 18760
rect 29196 18748 29224 18788
rect 29362 18776 29368 18788
rect 29420 18776 29426 18828
rect 30300 18816 30328 18924
rect 30650 18912 30656 18964
rect 30708 18952 30714 18964
rect 30708 18924 31892 18952
rect 30708 18912 30714 18924
rect 30742 18884 30748 18896
rect 30703 18856 30748 18884
rect 30742 18844 30748 18856
rect 30800 18844 30806 18896
rect 31570 18884 31576 18896
rect 30852 18856 31576 18884
rect 30852 18816 30880 18856
rect 31570 18844 31576 18856
rect 31628 18844 31634 18896
rect 30300 18788 30880 18816
rect 31205 18819 31263 18825
rect 31205 18785 31217 18819
rect 31251 18816 31263 18819
rect 31294 18816 31300 18828
rect 31251 18788 31300 18816
rect 31251 18785 31263 18788
rect 31205 18779 31263 18785
rect 31294 18776 31300 18788
rect 31352 18776 31358 18828
rect 31864 18816 31892 18924
rect 35710 18912 35716 18964
rect 35768 18952 35774 18964
rect 37366 18952 37372 18964
rect 35768 18924 37372 18952
rect 35768 18912 35774 18924
rect 37366 18912 37372 18924
rect 37424 18912 37430 18964
rect 37734 18912 37740 18964
rect 37792 18952 37798 18964
rect 37829 18955 37887 18961
rect 37829 18952 37841 18955
rect 37792 18924 37841 18952
rect 37792 18912 37798 18924
rect 37829 18921 37841 18924
rect 37875 18921 37887 18955
rect 37829 18915 37887 18921
rect 32858 18884 32864 18896
rect 32819 18856 32864 18884
rect 32858 18844 32864 18856
rect 32916 18844 32922 18896
rect 32950 18844 32956 18896
rect 33008 18884 33014 18896
rect 33008 18856 33732 18884
rect 33008 18844 33014 18856
rect 32125 18819 32183 18825
rect 32125 18816 32137 18819
rect 31864 18788 32137 18816
rect 32125 18785 32137 18788
rect 32171 18785 32183 18819
rect 32582 18816 32588 18828
rect 32543 18788 32588 18816
rect 32125 18779 32183 18785
rect 32140 18748 32168 18779
rect 32582 18776 32588 18788
rect 32640 18776 32646 18828
rect 33042 18776 33048 18828
rect 33100 18816 33106 18828
rect 33597 18819 33655 18825
rect 33597 18816 33609 18819
rect 33100 18788 33609 18816
rect 33100 18776 33106 18788
rect 33597 18785 33609 18788
rect 33643 18785 33655 18819
rect 33597 18779 33655 18785
rect 33502 18748 33508 18760
rect 29196 18720 31432 18748
rect 32140 18720 33508 18748
rect 27062 18680 27068 18692
rect 23952 18652 27068 18680
rect 27062 18640 27068 18652
rect 27120 18640 27126 18692
rect 28258 18680 28264 18692
rect 27632 18652 28264 18680
rect 25133 18615 25191 18621
rect 25133 18612 25145 18615
rect 23584 18584 25145 18612
rect 22649 18575 22707 18581
rect 25133 18581 25145 18584
rect 25179 18581 25191 18615
rect 25133 18575 25191 18581
rect 25869 18615 25927 18621
rect 25869 18581 25881 18615
rect 25915 18612 25927 18615
rect 27632 18612 27660 18652
rect 28258 18640 28264 18652
rect 28316 18640 28322 18692
rect 31404 18689 31432 18720
rect 33502 18708 33508 18720
rect 33560 18708 33566 18760
rect 33704 18748 33732 18856
rect 33778 18844 33784 18896
rect 33836 18884 33842 18896
rect 34425 18887 34483 18893
rect 34425 18884 34437 18887
rect 33836 18856 34437 18884
rect 33836 18844 33842 18856
rect 34425 18853 34437 18856
rect 34471 18853 34483 18887
rect 39025 18887 39083 18893
rect 39025 18884 39037 18887
rect 34425 18847 34483 18853
rect 35268 18856 39037 18884
rect 35268 18828 35296 18856
rect 39025 18853 39037 18856
rect 39071 18853 39083 18887
rect 39025 18847 39083 18853
rect 33962 18816 33968 18828
rect 33923 18788 33968 18816
rect 33962 18776 33968 18788
rect 34020 18776 34026 18828
rect 34241 18819 34299 18825
rect 34241 18785 34253 18819
rect 34287 18816 34299 18819
rect 34514 18816 34520 18828
rect 34287 18788 34520 18816
rect 34287 18785 34299 18788
rect 34241 18779 34299 18785
rect 34514 18776 34520 18788
rect 34572 18776 34578 18828
rect 35250 18816 35256 18828
rect 35163 18788 35256 18816
rect 35250 18776 35256 18788
rect 35308 18776 35314 18828
rect 35434 18816 35440 18828
rect 35395 18788 35440 18816
rect 35434 18776 35440 18788
rect 35492 18776 35498 18828
rect 35713 18819 35771 18825
rect 35713 18785 35725 18819
rect 35759 18785 35771 18819
rect 35713 18779 35771 18785
rect 36449 18819 36507 18825
rect 36449 18785 36461 18819
rect 36495 18816 36507 18819
rect 36538 18816 36544 18828
rect 36495 18788 36544 18816
rect 36495 18785 36507 18788
rect 36449 18779 36507 18785
rect 35728 18748 35756 18779
rect 36538 18776 36544 18788
rect 36596 18776 36602 18828
rect 36630 18776 36636 18828
rect 36688 18816 36694 18828
rect 36909 18819 36967 18825
rect 36909 18816 36921 18819
rect 36688 18788 36921 18816
rect 36688 18776 36694 18788
rect 36909 18785 36921 18788
rect 36955 18816 36967 18819
rect 37737 18819 37795 18825
rect 37737 18816 37749 18819
rect 36955 18788 37749 18816
rect 36955 18785 36967 18788
rect 36909 18779 36967 18785
rect 37737 18785 37749 18788
rect 37783 18785 37795 18819
rect 38286 18816 38292 18828
rect 38247 18788 38292 18816
rect 37737 18779 37795 18785
rect 38286 18776 38292 18788
rect 38344 18776 38350 18828
rect 38930 18816 38936 18828
rect 38891 18788 38936 18816
rect 38930 18776 38936 18788
rect 38988 18776 38994 18828
rect 33704 18720 35756 18748
rect 31389 18683 31447 18689
rect 31389 18649 31401 18683
rect 31435 18649 31447 18683
rect 31389 18643 31447 18649
rect 32490 18640 32496 18692
rect 32548 18680 32554 18692
rect 33413 18683 33471 18689
rect 33413 18680 33425 18683
rect 32548 18652 33425 18680
rect 32548 18640 32554 18652
rect 33413 18649 33425 18652
rect 33459 18680 33471 18683
rect 37182 18680 37188 18692
rect 33459 18652 37188 18680
rect 33459 18649 33471 18652
rect 33413 18643 33471 18649
rect 37182 18640 37188 18652
rect 37240 18640 37246 18692
rect 25915 18584 27660 18612
rect 25915 18581 25927 18584
rect 25869 18575 25927 18581
rect 27706 18572 27712 18624
rect 27764 18612 27770 18624
rect 28537 18615 28595 18621
rect 28537 18612 28549 18615
rect 27764 18584 28549 18612
rect 27764 18572 27770 18584
rect 28537 18581 28549 18584
rect 28583 18581 28595 18615
rect 28537 18575 28595 18581
rect 28902 18572 28908 18624
rect 28960 18612 28966 18624
rect 31202 18612 31208 18624
rect 28960 18584 31208 18612
rect 28960 18572 28966 18584
rect 31202 18572 31208 18584
rect 31260 18572 31266 18624
rect 36357 18615 36415 18621
rect 36357 18581 36369 18615
rect 36403 18612 36415 18615
rect 36538 18612 36544 18624
rect 36403 18584 36544 18612
rect 36403 18581 36415 18584
rect 36357 18575 36415 18581
rect 36538 18572 36544 18584
rect 36596 18572 36602 18624
rect 36630 18572 36636 18624
rect 36688 18612 36694 18624
rect 37093 18615 37151 18621
rect 37093 18612 37105 18615
rect 36688 18584 37105 18612
rect 36688 18572 36694 18584
rect 37093 18581 37105 18584
rect 37139 18581 37151 18615
rect 37093 18575 37151 18581
rect 1104 18522 39836 18544
rect 1104 18470 4246 18522
rect 4298 18470 4310 18522
rect 4362 18470 4374 18522
rect 4426 18470 4438 18522
rect 4490 18470 34966 18522
rect 35018 18470 35030 18522
rect 35082 18470 35094 18522
rect 35146 18470 35158 18522
rect 35210 18470 39836 18522
rect 1104 18448 39836 18470
rect 5166 18368 5172 18420
rect 5224 18408 5230 18420
rect 5905 18411 5963 18417
rect 5905 18408 5917 18411
rect 5224 18380 5917 18408
rect 5224 18368 5230 18380
rect 5905 18377 5917 18380
rect 5951 18377 5963 18411
rect 10226 18408 10232 18420
rect 5905 18371 5963 18377
rect 9876 18380 10232 18408
rect 2961 18275 3019 18281
rect 2961 18241 2973 18275
rect 3007 18272 3019 18275
rect 3050 18272 3056 18284
rect 3007 18244 3056 18272
rect 3007 18241 3019 18244
rect 2961 18235 3019 18241
rect 3050 18232 3056 18244
rect 3108 18232 3114 18284
rect 3513 18275 3571 18281
rect 3513 18241 3525 18275
rect 3559 18272 3571 18275
rect 4706 18272 4712 18284
rect 3559 18244 4712 18272
rect 3559 18241 3571 18244
rect 3513 18235 3571 18241
rect 4706 18232 4712 18244
rect 4764 18232 4770 18284
rect 8386 18272 8392 18284
rect 7116 18244 8392 18272
rect 3789 18207 3847 18213
rect 3789 18173 3801 18207
rect 3835 18173 3847 18207
rect 3970 18204 3976 18216
rect 3931 18176 3976 18204
rect 3789 18167 3847 18173
rect 3804 18136 3832 18167
rect 3970 18164 3976 18176
rect 4028 18164 4034 18216
rect 4433 18207 4491 18213
rect 4433 18173 4445 18207
rect 4479 18204 4491 18207
rect 4525 18207 4583 18213
rect 4525 18204 4537 18207
rect 4479 18176 4537 18204
rect 4479 18173 4491 18176
rect 4433 18167 4491 18173
rect 4525 18173 4537 18176
rect 4571 18173 4583 18207
rect 4525 18167 4583 18173
rect 4801 18207 4859 18213
rect 4801 18173 4813 18207
rect 4847 18204 4859 18207
rect 5442 18204 5448 18216
rect 4847 18176 5448 18204
rect 4847 18173 4859 18176
rect 4801 18167 4859 18173
rect 5442 18164 5448 18176
rect 5500 18164 5506 18216
rect 7116 18213 7144 18244
rect 8386 18232 8392 18244
rect 8444 18232 8450 18284
rect 9876 18281 9904 18380
rect 10226 18368 10232 18380
rect 10284 18368 10290 18420
rect 11238 18408 11244 18420
rect 11199 18380 11244 18408
rect 11238 18368 11244 18380
rect 11296 18368 11302 18420
rect 15378 18368 15384 18420
rect 15436 18408 15442 18420
rect 15436 18380 21588 18408
rect 15436 18368 15442 18380
rect 16206 18340 16212 18352
rect 16167 18312 16212 18340
rect 16206 18300 16212 18312
rect 16264 18300 16270 18352
rect 16761 18343 16819 18349
rect 16761 18309 16773 18343
rect 16807 18340 16819 18343
rect 19150 18340 19156 18352
rect 16807 18312 19156 18340
rect 16807 18309 16819 18312
rect 16761 18303 16819 18309
rect 19150 18300 19156 18312
rect 19208 18300 19214 18352
rect 21450 18300 21456 18352
rect 21508 18300 21514 18352
rect 21560 18349 21588 18380
rect 26786 18368 26792 18420
rect 26844 18408 26850 18420
rect 27430 18408 27436 18420
rect 26844 18380 27436 18408
rect 26844 18368 26850 18380
rect 27430 18368 27436 18380
rect 27488 18408 27494 18420
rect 28534 18408 28540 18420
rect 27488 18380 28540 18408
rect 27488 18368 27494 18380
rect 28534 18368 28540 18380
rect 28592 18368 28598 18420
rect 28629 18411 28687 18417
rect 28629 18377 28641 18411
rect 28675 18377 28687 18411
rect 28629 18371 28687 18377
rect 21545 18343 21603 18349
rect 21545 18309 21557 18343
rect 21591 18309 21603 18343
rect 21545 18303 21603 18309
rect 22830 18300 22836 18352
rect 22888 18340 22894 18352
rect 25682 18340 25688 18352
rect 22888 18312 25688 18340
rect 22888 18300 22894 18312
rect 25682 18300 25688 18312
rect 25740 18340 25746 18352
rect 28644 18340 28672 18371
rect 30282 18368 30288 18420
rect 30340 18408 30346 18420
rect 30340 18380 32536 18408
rect 30340 18368 30346 18380
rect 32306 18340 32312 18352
rect 25740 18312 28488 18340
rect 25740 18300 25746 18312
rect 9861 18275 9919 18281
rect 9861 18241 9873 18275
rect 9907 18241 9919 18275
rect 9861 18235 9919 18241
rect 11882 18232 11888 18284
rect 11940 18272 11946 18284
rect 14093 18275 14151 18281
rect 11940 18244 12572 18272
rect 11940 18232 11946 18244
rect 7101 18207 7159 18213
rect 7101 18173 7113 18207
rect 7147 18173 7159 18207
rect 7101 18167 7159 18173
rect 7745 18207 7803 18213
rect 7745 18173 7757 18207
rect 7791 18173 7803 18207
rect 8018 18204 8024 18216
rect 7979 18176 8024 18204
rect 7745 18167 7803 18173
rect 4614 18136 4620 18148
rect 3804 18108 4620 18136
rect 4614 18096 4620 18108
rect 4672 18096 4678 18148
rect 6086 18096 6092 18148
rect 6144 18136 6150 18148
rect 7760 18136 7788 18167
rect 8018 18164 8024 18176
rect 8076 18164 8082 18216
rect 10137 18207 10195 18213
rect 10137 18173 10149 18207
rect 10183 18204 10195 18207
rect 10226 18204 10232 18216
rect 10183 18176 10232 18204
rect 10183 18173 10195 18176
rect 10137 18167 10195 18173
rect 10226 18164 10232 18176
rect 10284 18164 10290 18216
rect 11698 18164 11704 18216
rect 11756 18204 11762 18216
rect 12544 18213 12572 18244
rect 12912 18244 14044 18272
rect 12437 18207 12495 18213
rect 12437 18204 12449 18207
rect 11756 18176 12449 18204
rect 11756 18164 11762 18176
rect 12437 18173 12449 18176
rect 12483 18173 12495 18207
rect 12437 18167 12495 18173
rect 12529 18207 12587 18213
rect 12529 18173 12541 18207
rect 12575 18173 12587 18207
rect 12529 18167 12587 18173
rect 9398 18136 9404 18148
rect 6144 18108 7788 18136
rect 6144 18096 6150 18108
rect 4433 18071 4491 18077
rect 4433 18037 4445 18071
rect 4479 18068 4491 18071
rect 6822 18068 6828 18080
rect 4479 18040 6828 18068
rect 4479 18037 4491 18040
rect 4433 18031 4491 18037
rect 6822 18028 6828 18040
rect 6880 18028 6886 18080
rect 7193 18071 7251 18077
rect 7193 18037 7205 18071
rect 7239 18068 7251 18071
rect 7374 18068 7380 18080
rect 7239 18040 7380 18068
rect 7239 18037 7251 18040
rect 7193 18031 7251 18037
rect 7374 18028 7380 18040
rect 7432 18028 7438 18080
rect 7760 18068 7788 18108
rect 8680 18108 9404 18136
rect 8680 18068 8708 18108
rect 9398 18096 9404 18108
rect 9456 18096 9462 18148
rect 12912 18136 12940 18244
rect 13814 18204 13820 18216
rect 13775 18176 13820 18204
rect 13814 18164 13820 18176
rect 13872 18164 13878 18216
rect 14016 18204 14044 18244
rect 14093 18241 14105 18275
rect 14139 18272 14151 18275
rect 16114 18272 16120 18284
rect 14139 18244 16120 18272
rect 14139 18241 14151 18244
rect 14093 18235 14151 18241
rect 16114 18232 16120 18244
rect 16172 18232 16178 18284
rect 17310 18272 17316 18284
rect 16776 18244 17316 18272
rect 16025 18207 16083 18213
rect 16025 18204 16037 18207
rect 14016 18176 16037 18204
rect 16025 18173 16037 18176
rect 16071 18204 16083 18207
rect 16776 18204 16804 18244
rect 17310 18232 17316 18244
rect 17368 18232 17374 18284
rect 19610 18272 19616 18284
rect 17420 18244 19196 18272
rect 19571 18244 19616 18272
rect 16942 18204 16948 18216
rect 16071 18176 16804 18204
rect 16903 18176 16948 18204
rect 16071 18173 16083 18176
rect 16025 18167 16083 18173
rect 16942 18164 16948 18176
rect 17000 18164 17006 18216
rect 17034 18164 17040 18216
rect 17092 18204 17098 18216
rect 17092 18176 17137 18204
rect 17092 18164 17098 18176
rect 10796 18108 12940 18136
rect 12989 18139 13047 18145
rect 7760 18040 8708 18068
rect 9309 18071 9367 18077
rect 9309 18037 9321 18071
rect 9355 18068 9367 18071
rect 10796 18068 10824 18108
rect 12989 18105 13001 18139
rect 13035 18105 13047 18139
rect 17420 18136 17448 18244
rect 19168 18216 19196 18244
rect 19610 18232 19616 18244
rect 19668 18232 19674 18284
rect 19702 18232 19708 18284
rect 19760 18272 19766 18284
rect 21468 18272 21496 18300
rect 19760 18244 21496 18272
rect 19760 18232 19766 18244
rect 21910 18232 21916 18284
rect 21968 18272 21974 18284
rect 22281 18275 22339 18281
rect 22281 18272 22293 18275
rect 21968 18244 22293 18272
rect 21968 18232 21974 18244
rect 22281 18241 22293 18244
rect 22327 18241 22339 18275
rect 25866 18272 25872 18284
rect 22281 18235 22339 18241
rect 24044 18244 25872 18272
rect 18414 18164 18420 18216
rect 18472 18204 18478 18216
rect 18601 18207 18659 18213
rect 18601 18204 18613 18207
rect 18472 18176 18613 18204
rect 18472 18164 18478 18176
rect 18601 18173 18613 18176
rect 18647 18173 18659 18207
rect 18601 18167 18659 18173
rect 19150 18164 19156 18216
rect 19208 18164 19214 18216
rect 19337 18207 19395 18213
rect 19337 18173 19349 18207
rect 19383 18204 19395 18207
rect 20530 18204 20536 18216
rect 19383 18176 20536 18204
rect 19383 18173 19395 18176
rect 19337 18167 19395 18173
rect 12989 18099 13047 18105
rect 15028 18108 17448 18136
rect 17497 18139 17555 18145
rect 9355 18040 10824 18068
rect 13004 18068 13032 18099
rect 15028 18068 15056 18108
rect 17497 18105 17509 18139
rect 17543 18136 17555 18139
rect 17678 18136 17684 18148
rect 17543 18108 17684 18136
rect 17543 18105 17555 18108
rect 17497 18099 17555 18105
rect 17678 18096 17684 18108
rect 17736 18096 17742 18148
rect 17770 18096 17776 18148
rect 17828 18136 17834 18148
rect 19352 18136 19380 18167
rect 20530 18164 20536 18176
rect 20588 18164 20594 18216
rect 21358 18164 21364 18216
rect 21416 18204 21422 18216
rect 21453 18207 21511 18213
rect 21453 18204 21465 18207
rect 21416 18176 21465 18204
rect 21416 18164 21422 18176
rect 21453 18173 21465 18176
rect 21499 18173 21511 18207
rect 21453 18167 21511 18173
rect 21818 18164 21824 18216
rect 21876 18204 21882 18216
rect 22189 18207 22247 18213
rect 22189 18204 22201 18207
rect 21876 18176 22201 18204
rect 21876 18164 21882 18176
rect 22189 18173 22201 18176
rect 22235 18204 22247 18207
rect 24044 18204 24072 18244
rect 25866 18232 25872 18244
rect 25924 18232 25930 18284
rect 26881 18275 26939 18281
rect 26881 18241 26893 18275
rect 26927 18272 26939 18275
rect 28350 18272 28356 18284
rect 26927 18244 28356 18272
rect 26927 18241 26939 18244
rect 26881 18235 26939 18241
rect 28350 18232 28356 18244
rect 28408 18232 28414 18284
rect 22235 18176 24072 18204
rect 24121 18207 24179 18213
rect 22235 18173 22247 18176
rect 22189 18167 22247 18173
rect 24121 18173 24133 18207
rect 24167 18173 24179 18207
rect 24121 18167 24179 18173
rect 24397 18207 24455 18213
rect 24397 18173 24409 18207
rect 24443 18204 24455 18207
rect 24581 18207 24639 18213
rect 24443 18176 24532 18204
rect 24443 18173 24455 18176
rect 24397 18167 24455 18173
rect 24136 18136 24164 18167
rect 17828 18108 19380 18136
rect 20272 18108 24164 18136
rect 17828 18096 17834 18108
rect 15194 18068 15200 18080
rect 13004 18040 15056 18068
rect 15155 18040 15200 18068
rect 9355 18037 9367 18040
rect 9309 18031 9367 18037
rect 15194 18028 15200 18040
rect 15252 18028 15258 18080
rect 15930 18028 15936 18080
rect 15988 18068 15994 18080
rect 18785 18071 18843 18077
rect 18785 18068 18797 18071
rect 15988 18040 18797 18068
rect 15988 18028 15994 18040
rect 18785 18037 18797 18040
rect 18831 18068 18843 18071
rect 20272 18068 20300 18108
rect 18831 18040 20300 18068
rect 18831 18037 18843 18040
rect 18785 18031 18843 18037
rect 20346 18028 20352 18080
rect 20404 18068 20410 18080
rect 20717 18071 20775 18077
rect 20717 18068 20729 18071
rect 20404 18040 20729 18068
rect 20404 18028 20410 18040
rect 20717 18037 20729 18040
rect 20763 18037 20775 18071
rect 20717 18031 20775 18037
rect 21174 18028 21180 18080
rect 21232 18068 21238 18080
rect 24504 18068 24532 18176
rect 24581 18173 24593 18207
rect 24627 18204 24639 18207
rect 24762 18204 24768 18216
rect 24627 18176 24768 18204
rect 24627 18173 24639 18176
rect 24581 18167 24639 18173
rect 24762 18164 24768 18176
rect 24820 18164 24826 18216
rect 24857 18207 24915 18213
rect 24857 18173 24869 18207
rect 24903 18204 24915 18207
rect 24946 18204 24952 18216
rect 24903 18176 24952 18204
rect 24903 18173 24915 18176
rect 24857 18167 24915 18173
rect 24946 18164 24952 18176
rect 25004 18164 25010 18216
rect 25130 18213 25136 18216
rect 25110 18207 25136 18213
rect 25110 18173 25122 18207
rect 25110 18167 25136 18173
rect 25130 18164 25136 18167
rect 25188 18164 25194 18216
rect 26418 18204 26424 18216
rect 25608 18176 26424 18204
rect 24780 18136 24808 18164
rect 25608 18136 25636 18176
rect 26418 18164 26424 18176
rect 26476 18164 26482 18216
rect 26697 18207 26755 18213
rect 26697 18173 26709 18207
rect 26743 18204 26755 18207
rect 26786 18204 26792 18216
rect 26743 18176 26792 18204
rect 26743 18173 26755 18176
rect 26697 18167 26755 18173
rect 26786 18164 26792 18176
rect 26844 18164 26850 18216
rect 27154 18204 27160 18216
rect 27115 18176 27160 18204
rect 27154 18164 27160 18176
rect 27212 18164 27218 18216
rect 27249 18207 27307 18213
rect 27249 18173 27261 18207
rect 27295 18173 27307 18207
rect 27706 18204 27712 18216
rect 27667 18176 27712 18204
rect 27249 18167 27307 18173
rect 24780 18108 25636 18136
rect 25685 18139 25743 18145
rect 25685 18105 25697 18139
rect 25731 18136 25743 18139
rect 26878 18136 26884 18148
rect 25731 18108 26884 18136
rect 25731 18105 25743 18108
rect 25685 18099 25743 18105
rect 26878 18096 26884 18108
rect 26936 18096 26942 18148
rect 27062 18096 27068 18148
rect 27120 18136 27126 18148
rect 27264 18136 27292 18167
rect 27706 18164 27712 18176
rect 27764 18164 27770 18216
rect 28460 18213 28488 18312
rect 28552 18312 28672 18340
rect 28920 18312 29868 18340
rect 32267 18312 32312 18340
rect 28445 18207 28503 18213
rect 28445 18173 28457 18207
rect 28491 18173 28503 18207
rect 28445 18167 28503 18173
rect 27120 18108 27292 18136
rect 28552 18136 28580 18312
rect 28626 18164 28632 18216
rect 28684 18204 28690 18216
rect 28920 18204 28948 18312
rect 29546 18272 29552 18284
rect 29472 18244 29552 18272
rect 29472 18213 29500 18244
rect 29546 18232 29552 18244
rect 29604 18232 29610 18284
rect 28684 18176 28948 18204
rect 29457 18207 29515 18213
rect 28684 18164 28690 18176
rect 29457 18173 29469 18207
rect 29503 18173 29515 18207
rect 29638 18204 29644 18216
rect 29599 18176 29644 18204
rect 29457 18167 29515 18173
rect 29638 18164 29644 18176
rect 29696 18164 29702 18216
rect 29840 18213 29868 18312
rect 32306 18300 32312 18312
rect 32364 18300 32370 18352
rect 30006 18232 30012 18284
rect 30064 18272 30070 18284
rect 31481 18275 31539 18281
rect 31481 18272 31493 18275
rect 30064 18244 31493 18272
rect 30064 18232 30070 18244
rect 31481 18241 31493 18244
rect 31527 18241 31539 18275
rect 32508 18272 32536 18380
rect 36906 18368 36912 18420
rect 36964 18408 36970 18420
rect 37001 18411 37059 18417
rect 37001 18408 37013 18411
rect 36964 18380 37013 18408
rect 36964 18368 36970 18380
rect 37001 18377 37013 18380
rect 37047 18408 37059 18411
rect 37366 18408 37372 18420
rect 37047 18380 37372 18408
rect 37047 18377 37059 18380
rect 37001 18371 37059 18377
rect 37366 18368 37372 18380
rect 37424 18368 37430 18420
rect 32674 18340 32680 18352
rect 32635 18312 32680 18340
rect 32674 18300 32680 18312
rect 32732 18300 32738 18352
rect 32508 18244 32628 18272
rect 31481 18235 31539 18241
rect 29825 18207 29883 18213
rect 29825 18173 29837 18207
rect 29871 18173 29883 18207
rect 29825 18167 29883 18173
rect 30837 18207 30895 18213
rect 30837 18173 30849 18207
rect 30883 18204 30895 18207
rect 30883 18176 31156 18204
rect 30883 18173 30895 18176
rect 30837 18167 30895 18173
rect 31128 18136 31156 18176
rect 31202 18164 31208 18216
rect 31260 18204 31266 18216
rect 32490 18204 32496 18216
rect 31260 18176 31305 18204
rect 32451 18176 32496 18204
rect 31260 18164 31266 18176
rect 32490 18164 32496 18176
rect 32548 18164 32554 18216
rect 32600 18213 32628 18244
rect 33318 18232 33324 18284
rect 33376 18272 33382 18284
rect 33413 18275 33471 18281
rect 33413 18272 33425 18275
rect 33376 18244 33425 18272
rect 33376 18232 33382 18244
rect 33413 18241 33425 18244
rect 33459 18241 33471 18275
rect 36078 18272 36084 18284
rect 36039 18244 36084 18272
rect 33413 18235 33471 18241
rect 36078 18232 36084 18244
rect 36136 18232 36142 18284
rect 36170 18232 36176 18284
rect 36228 18272 36234 18284
rect 37369 18275 37427 18281
rect 37369 18272 37381 18275
rect 36228 18244 37381 18272
rect 36228 18232 36234 18244
rect 37369 18241 37381 18244
rect 37415 18241 37427 18275
rect 37369 18235 37427 18241
rect 32585 18207 32643 18213
rect 32585 18173 32597 18207
rect 32631 18204 32643 18207
rect 33042 18204 33048 18216
rect 32631 18176 33048 18204
rect 32631 18173 32643 18176
rect 32585 18167 32643 18173
rect 33042 18164 33048 18176
rect 33100 18164 33106 18216
rect 33226 18204 33232 18216
rect 33187 18176 33232 18204
rect 33226 18164 33232 18176
rect 33284 18164 33290 18216
rect 33502 18164 33508 18216
rect 33560 18204 33566 18216
rect 34149 18207 34207 18213
rect 34149 18204 34161 18207
rect 33560 18176 34161 18204
rect 33560 18164 33566 18176
rect 34149 18173 34161 18176
rect 34195 18173 34207 18207
rect 35250 18204 35256 18216
rect 35211 18176 35256 18204
rect 34149 18167 34207 18173
rect 35250 18164 35256 18176
rect 35308 18164 35314 18216
rect 35434 18204 35440 18216
rect 35395 18176 35440 18204
rect 35434 18164 35440 18176
rect 35492 18164 35498 18216
rect 35802 18164 35808 18216
rect 35860 18204 35866 18216
rect 35897 18207 35955 18213
rect 35897 18204 35909 18207
rect 35860 18176 35909 18204
rect 35860 18164 35866 18176
rect 35897 18173 35909 18176
rect 35943 18173 35955 18207
rect 36446 18204 36452 18216
rect 36407 18176 36452 18204
rect 35897 18167 35955 18173
rect 36446 18164 36452 18176
rect 36504 18164 36510 18216
rect 37182 18204 37188 18216
rect 37143 18176 37188 18204
rect 37182 18164 37188 18176
rect 37240 18164 37246 18216
rect 37642 18204 37648 18216
rect 37603 18176 37648 18204
rect 37642 18164 37648 18176
rect 37700 18164 37706 18216
rect 32950 18136 32956 18148
rect 28552 18108 31064 18136
rect 31128 18108 32956 18136
rect 27120 18096 27126 18108
rect 28994 18068 29000 18080
rect 21232 18040 29000 18068
rect 21232 18028 21238 18040
rect 28994 18028 29000 18040
rect 29052 18028 29058 18080
rect 30558 18028 30564 18080
rect 30616 18068 30622 18080
rect 30745 18071 30803 18077
rect 30745 18068 30757 18071
rect 30616 18040 30757 18068
rect 30616 18028 30622 18040
rect 30745 18037 30757 18040
rect 30791 18037 30803 18071
rect 31036 18068 31064 18108
rect 32950 18096 32956 18108
rect 33008 18096 33014 18148
rect 34241 18139 34299 18145
rect 34241 18105 34253 18139
rect 34287 18136 34299 18139
rect 34514 18136 34520 18148
rect 34287 18108 34520 18136
rect 34287 18105 34299 18108
rect 34241 18099 34299 18105
rect 34514 18096 34520 18108
rect 34572 18136 34578 18148
rect 35820 18136 35848 18164
rect 34572 18108 35848 18136
rect 34572 18096 34578 18108
rect 33870 18068 33876 18080
rect 31036 18040 33876 18068
rect 30745 18031 30803 18037
rect 33870 18028 33876 18040
rect 33928 18028 33934 18080
rect 38286 18028 38292 18080
rect 38344 18068 38350 18080
rect 38749 18071 38807 18077
rect 38749 18068 38761 18071
rect 38344 18040 38761 18068
rect 38344 18028 38350 18040
rect 38749 18037 38761 18040
rect 38795 18037 38807 18071
rect 38749 18031 38807 18037
rect 1104 17978 39836 18000
rect 1104 17926 19606 17978
rect 19658 17926 19670 17978
rect 19722 17926 19734 17978
rect 19786 17926 19798 17978
rect 19850 17926 39836 17978
rect 1104 17904 39836 17926
rect 9582 17824 9588 17876
rect 9640 17864 9646 17876
rect 22462 17864 22468 17876
rect 9640 17836 14780 17864
rect 9640 17824 9646 17836
rect 3053 17799 3111 17805
rect 3053 17765 3065 17799
rect 3099 17796 3111 17799
rect 3142 17796 3148 17808
rect 3099 17768 3148 17796
rect 3099 17765 3111 17768
rect 3053 17759 3111 17765
rect 3142 17756 3148 17768
rect 3200 17756 3206 17808
rect 7745 17799 7803 17805
rect 7745 17765 7757 17799
rect 7791 17796 7803 17799
rect 8018 17796 8024 17808
rect 7791 17768 8024 17796
rect 7791 17765 7803 17768
rect 7745 17759 7803 17765
rect 8018 17756 8024 17768
rect 8076 17756 8082 17808
rect 10229 17799 10287 17805
rect 10229 17765 10241 17799
rect 10275 17796 10287 17799
rect 10778 17796 10784 17808
rect 10275 17768 10784 17796
rect 10275 17765 10287 17768
rect 10229 17759 10287 17765
rect 10778 17756 10784 17768
rect 10836 17756 10842 17808
rect 14752 17805 14780 17836
rect 18524 17836 22468 17864
rect 14737 17799 14795 17805
rect 14737 17765 14749 17799
rect 14783 17765 14795 17799
rect 14737 17759 14795 17765
rect 15657 17799 15715 17805
rect 15657 17765 15669 17799
rect 15703 17796 15715 17799
rect 15703 17768 17632 17796
rect 15703 17765 15715 17768
rect 15657 17759 15715 17765
rect 1394 17728 1400 17740
rect 1355 17700 1400 17728
rect 1394 17688 1400 17700
rect 1452 17688 1458 17740
rect 5169 17731 5227 17737
rect 5169 17697 5181 17731
rect 5215 17728 5227 17731
rect 5258 17728 5264 17740
rect 5215 17700 5264 17728
rect 5215 17697 5227 17700
rect 5169 17691 5227 17697
rect 5258 17688 5264 17700
rect 5316 17688 5322 17740
rect 5353 17731 5411 17737
rect 5353 17697 5365 17731
rect 5399 17728 5411 17731
rect 7374 17728 7380 17740
rect 5399 17700 7380 17728
rect 5399 17697 5411 17700
rect 5353 17691 5411 17697
rect 7374 17688 7380 17700
rect 7432 17688 7438 17740
rect 7926 17688 7932 17740
rect 7984 17728 7990 17740
rect 8389 17731 8447 17737
rect 8389 17728 8401 17731
rect 7984 17700 8401 17728
rect 7984 17688 7990 17700
rect 8389 17697 8401 17700
rect 8435 17697 8447 17731
rect 8389 17691 8447 17697
rect 8846 17688 8852 17740
rect 8904 17728 8910 17740
rect 9769 17731 9827 17737
rect 9769 17728 9781 17731
rect 8904 17700 9781 17728
rect 8904 17688 8910 17700
rect 9769 17697 9781 17700
rect 9815 17697 9827 17731
rect 11422 17728 11428 17740
rect 11383 17700 11428 17728
rect 9769 17691 9827 17697
rect 11422 17688 11428 17700
rect 11480 17688 11486 17740
rect 11790 17728 11796 17740
rect 11751 17700 11796 17728
rect 11790 17688 11796 17700
rect 11848 17688 11854 17740
rect 11974 17728 11980 17740
rect 11935 17700 11980 17728
rect 11974 17688 11980 17700
rect 12032 17688 12038 17740
rect 12618 17728 12624 17740
rect 12579 17700 12624 17728
rect 12618 17688 12624 17700
rect 12676 17688 12682 17740
rect 13170 17728 13176 17740
rect 13131 17700 13176 17728
rect 13170 17688 13176 17700
rect 13228 17688 13234 17740
rect 14277 17731 14335 17737
rect 14277 17697 14289 17731
rect 14323 17728 14335 17731
rect 15194 17728 15200 17740
rect 14323 17700 15200 17728
rect 14323 17697 14335 17700
rect 14277 17691 14335 17697
rect 15194 17688 15200 17700
rect 15252 17688 15258 17740
rect 15838 17728 15844 17740
rect 15799 17700 15844 17728
rect 15838 17688 15844 17700
rect 15896 17688 15902 17740
rect 17604 17737 17632 17768
rect 17313 17731 17371 17737
rect 17313 17697 17325 17731
rect 17359 17697 17371 17731
rect 17313 17691 17371 17697
rect 17589 17731 17647 17737
rect 17589 17697 17601 17731
rect 17635 17728 17647 17731
rect 18046 17728 18052 17740
rect 17635 17700 18052 17728
rect 17635 17697 17647 17700
rect 17589 17691 17647 17697
rect 1673 17663 1731 17669
rect 1673 17629 1685 17663
rect 1719 17660 1731 17663
rect 4062 17660 4068 17672
rect 1719 17632 4068 17660
rect 1719 17629 1731 17632
rect 1673 17623 1731 17629
rect 4062 17620 4068 17632
rect 4120 17620 4126 17672
rect 5442 17660 5448 17672
rect 5403 17632 5448 17660
rect 5442 17620 5448 17632
rect 5500 17620 5506 17672
rect 6086 17660 6092 17672
rect 6047 17632 6092 17660
rect 6086 17620 6092 17632
rect 6144 17620 6150 17672
rect 6365 17663 6423 17669
rect 6365 17629 6377 17663
rect 6411 17660 6423 17663
rect 7190 17660 7196 17672
rect 6411 17632 7196 17660
rect 6411 17629 6423 17632
rect 6365 17623 6423 17629
rect 7190 17620 7196 17632
rect 7248 17620 7254 17672
rect 9677 17663 9735 17669
rect 9677 17629 9689 17663
rect 9723 17660 9735 17663
rect 11698 17660 11704 17672
rect 9723 17632 11704 17660
rect 9723 17629 9735 17632
rect 9677 17623 9735 17629
rect 8570 17592 8576 17604
rect 8531 17564 8576 17592
rect 8570 17552 8576 17564
rect 8628 17552 8634 17604
rect 5074 17484 5080 17536
rect 5132 17524 5138 17536
rect 9692 17524 9720 17623
rect 11698 17620 11704 17632
rect 11756 17620 11762 17672
rect 12253 17663 12311 17669
rect 12253 17629 12265 17663
rect 12299 17660 12311 17663
rect 12710 17660 12716 17672
rect 12299 17632 12716 17660
rect 12299 17629 12311 17632
rect 12253 17623 12311 17629
rect 12710 17620 12716 17632
rect 12768 17620 12774 17672
rect 14185 17663 14243 17669
rect 14185 17629 14197 17663
rect 14231 17629 14243 17663
rect 14185 17623 14243 17629
rect 11330 17552 11336 17604
rect 11388 17592 11394 17604
rect 13262 17592 13268 17604
rect 11388 17564 13268 17592
rect 11388 17552 11394 17564
rect 13262 17552 13268 17564
rect 13320 17552 13326 17604
rect 14200 17592 14228 17623
rect 15654 17620 15660 17672
rect 15712 17660 15718 17672
rect 15749 17663 15807 17669
rect 15749 17660 15761 17663
rect 15712 17632 15761 17660
rect 15712 17620 15718 17632
rect 15749 17629 15761 17632
rect 15795 17629 15807 17663
rect 15749 17623 15807 17629
rect 16206 17592 16212 17604
rect 14200 17564 16212 17592
rect 16206 17552 16212 17564
rect 16264 17552 16270 17604
rect 17034 17552 17040 17604
rect 17092 17592 17098 17604
rect 17221 17595 17279 17601
rect 17221 17592 17233 17595
rect 17092 17564 17233 17592
rect 17092 17552 17098 17564
rect 17221 17561 17233 17564
rect 17267 17561 17279 17595
rect 17328 17592 17356 17691
rect 18046 17688 18052 17700
rect 18104 17688 18110 17740
rect 18524 17737 18552 17836
rect 22462 17824 22468 17836
rect 22520 17824 22526 17876
rect 25866 17864 25872 17876
rect 25779 17836 25872 17864
rect 25866 17824 25872 17836
rect 25924 17864 25930 17876
rect 25924 17836 28764 17864
rect 25924 17824 25930 17836
rect 19334 17756 19340 17808
rect 19392 17796 19398 17808
rect 20162 17796 20168 17808
rect 19392 17768 20168 17796
rect 19392 17756 19398 17768
rect 18141 17731 18199 17737
rect 18141 17697 18153 17731
rect 18187 17697 18199 17731
rect 18141 17691 18199 17697
rect 18509 17731 18567 17737
rect 18509 17697 18521 17731
rect 18555 17697 18567 17731
rect 18509 17691 18567 17697
rect 18156 17660 18184 17691
rect 18782 17688 18788 17740
rect 18840 17728 18846 17740
rect 19061 17731 19119 17737
rect 19061 17728 19073 17731
rect 18840 17700 19073 17728
rect 18840 17688 18846 17700
rect 19061 17697 19073 17700
rect 19107 17728 19119 17731
rect 19702 17728 19708 17740
rect 19107 17700 19708 17728
rect 19107 17697 19119 17700
rect 19061 17691 19119 17697
rect 19702 17688 19708 17700
rect 19760 17688 19766 17740
rect 20088 17737 20116 17768
rect 20162 17756 20168 17768
rect 20220 17756 20226 17808
rect 26234 17756 26240 17808
rect 26292 17796 26298 17808
rect 26513 17799 26571 17805
rect 26513 17796 26525 17799
rect 26292 17768 26525 17796
rect 26292 17756 26298 17768
rect 26513 17765 26525 17768
rect 26559 17765 26571 17799
rect 26513 17759 26571 17765
rect 27062 17756 27068 17808
rect 27120 17796 27126 17808
rect 28626 17796 28632 17808
rect 27120 17768 28632 17796
rect 27120 17756 27126 17768
rect 28626 17756 28632 17768
rect 28684 17756 28690 17808
rect 19797 17731 19855 17737
rect 19797 17697 19809 17731
rect 19843 17697 19855 17731
rect 19797 17691 19855 17697
rect 20073 17731 20131 17737
rect 20073 17697 20085 17731
rect 20119 17697 20131 17731
rect 22554 17728 22560 17740
rect 20073 17691 20131 17697
rect 20180 17700 22560 17728
rect 18690 17660 18696 17672
rect 18156 17632 18696 17660
rect 18690 17620 18696 17632
rect 18748 17620 18754 17672
rect 19812 17660 19840 17691
rect 20180 17660 20208 17700
rect 22554 17688 22560 17700
rect 22612 17688 22618 17740
rect 23842 17728 23848 17740
rect 23803 17700 23848 17728
rect 23842 17688 23848 17700
rect 23900 17688 23906 17740
rect 24578 17688 24584 17740
rect 24636 17728 24642 17740
rect 25685 17731 25743 17737
rect 25685 17728 25697 17731
rect 24636 17700 25697 17728
rect 24636 17688 24642 17700
rect 25685 17697 25697 17700
rect 25731 17697 25743 17731
rect 25685 17691 25743 17697
rect 19812 17632 20208 17660
rect 20530 17620 20536 17672
rect 20588 17660 20594 17672
rect 21453 17663 21511 17669
rect 21453 17660 21465 17663
rect 20588 17632 21465 17660
rect 20588 17620 20594 17632
rect 21453 17629 21465 17632
rect 21499 17629 21511 17663
rect 21453 17623 21511 17629
rect 21729 17663 21787 17669
rect 21729 17629 21741 17663
rect 21775 17660 21787 17663
rect 21818 17660 21824 17672
rect 21775 17632 21824 17660
rect 21775 17629 21787 17632
rect 21729 17623 21787 17629
rect 21818 17620 21824 17632
rect 21876 17620 21882 17672
rect 23569 17663 23627 17669
rect 23569 17629 23581 17663
rect 23615 17660 23627 17663
rect 24762 17660 24768 17672
rect 23615 17632 24768 17660
rect 23615 17629 23627 17632
rect 23569 17623 23627 17629
rect 24762 17620 24768 17632
rect 24820 17620 24826 17672
rect 19150 17592 19156 17604
rect 17328 17564 19156 17592
rect 17221 17555 17279 17561
rect 19150 17552 19156 17564
rect 19208 17592 19214 17604
rect 19613 17595 19671 17601
rect 19613 17592 19625 17595
rect 19208 17564 19625 17592
rect 19208 17552 19214 17564
rect 19613 17561 19625 17564
rect 19659 17561 19671 17595
rect 25700 17592 25728 17691
rect 26878 17688 26884 17740
rect 26936 17728 26942 17740
rect 26973 17731 27031 17737
rect 26973 17728 26985 17731
rect 26936 17700 26985 17728
rect 26936 17688 26942 17700
rect 26973 17697 26985 17700
rect 27019 17697 27031 17731
rect 26973 17691 27031 17697
rect 27154 17688 27160 17740
rect 27212 17728 27218 17740
rect 27341 17731 27399 17737
rect 27341 17728 27353 17731
rect 27212 17700 27353 17728
rect 27212 17688 27218 17700
rect 27341 17697 27353 17700
rect 27387 17697 27399 17731
rect 27341 17691 27399 17697
rect 27430 17688 27436 17740
rect 27488 17728 27494 17740
rect 28534 17728 28540 17740
rect 27488 17700 27533 17728
rect 28495 17700 28540 17728
rect 27488 17688 27494 17700
rect 28534 17688 28540 17700
rect 28592 17688 28598 17740
rect 28736 17737 28764 17836
rect 28994 17824 29000 17876
rect 29052 17864 29058 17876
rect 29362 17864 29368 17876
rect 29052 17836 29368 17864
rect 29052 17824 29058 17836
rect 29362 17824 29368 17836
rect 29420 17824 29426 17876
rect 32582 17824 32588 17876
rect 32640 17864 32646 17876
rect 32640 17836 33272 17864
rect 32640 17824 32646 17836
rect 29178 17756 29184 17808
rect 29236 17796 29242 17808
rect 30650 17796 30656 17808
rect 29236 17768 30656 17796
rect 29236 17756 29242 17768
rect 30650 17756 30656 17768
rect 30708 17756 30714 17808
rect 33244 17796 33272 17836
rect 33502 17824 33508 17876
rect 33560 17864 33566 17876
rect 33689 17867 33747 17873
rect 33689 17864 33701 17867
rect 33560 17836 33701 17864
rect 33560 17824 33566 17836
rect 33689 17833 33701 17836
rect 33735 17833 33747 17867
rect 33689 17827 33747 17833
rect 35894 17824 35900 17876
rect 35952 17864 35958 17876
rect 36909 17867 36967 17873
rect 36909 17864 36921 17867
rect 35952 17836 36921 17864
rect 35952 17824 35958 17836
rect 36909 17833 36921 17836
rect 36955 17833 36967 17867
rect 36909 17827 36967 17833
rect 37642 17824 37648 17876
rect 37700 17864 37706 17876
rect 37829 17867 37887 17873
rect 37829 17864 37841 17867
rect 37700 17836 37841 17864
rect 37700 17824 37706 17836
rect 37829 17833 37841 17836
rect 37875 17833 37887 17867
rect 37829 17827 37887 17833
rect 38010 17824 38016 17876
rect 38068 17864 38074 17876
rect 39025 17867 39083 17873
rect 39025 17864 39037 17867
rect 38068 17836 39037 17864
rect 38068 17824 38074 17836
rect 39025 17833 39037 17836
rect 39071 17833 39083 17867
rect 39025 17827 39083 17833
rect 33244 17768 36768 17796
rect 28721 17731 28779 17737
rect 28721 17697 28733 17731
rect 28767 17697 28779 17731
rect 28721 17691 28779 17697
rect 28626 17660 28632 17672
rect 28587 17632 28632 17660
rect 28626 17620 28632 17632
rect 28684 17620 28690 17672
rect 29196 17660 29224 17756
rect 36740 17740 36768 17768
rect 29362 17728 29368 17740
rect 29323 17700 29368 17728
rect 29362 17688 29368 17700
rect 29420 17688 29426 17740
rect 29546 17728 29552 17740
rect 29507 17700 29552 17728
rect 29546 17688 29552 17700
rect 29604 17688 29610 17740
rect 29638 17688 29644 17740
rect 29696 17728 29702 17740
rect 29917 17731 29975 17737
rect 29917 17728 29929 17731
rect 29696 17700 29929 17728
rect 29696 17688 29702 17700
rect 29917 17697 29929 17700
rect 29963 17697 29975 17731
rect 30834 17728 30840 17740
rect 30795 17700 30840 17728
rect 29917 17691 29975 17697
rect 30834 17688 30840 17700
rect 30892 17688 30898 17740
rect 31389 17731 31447 17737
rect 31389 17728 31401 17731
rect 30944 17700 31401 17728
rect 28736 17632 29224 17660
rect 28736 17592 28764 17632
rect 25700 17564 28764 17592
rect 19613 17555 19671 17561
rect 29270 17552 29276 17604
rect 29328 17592 29334 17604
rect 30098 17592 30104 17604
rect 29328 17564 30104 17592
rect 29328 17552 29334 17564
rect 30098 17552 30104 17564
rect 30156 17552 30162 17604
rect 5132 17496 9720 17524
rect 5132 17484 5138 17496
rect 10318 17484 10324 17536
rect 10376 17524 10382 17536
rect 15657 17527 15715 17533
rect 15657 17524 15669 17527
rect 10376 17496 15669 17524
rect 10376 17484 10382 17496
rect 15657 17493 15669 17496
rect 15703 17493 15715 17527
rect 15657 17487 15715 17493
rect 15746 17484 15752 17536
rect 15804 17524 15810 17536
rect 16025 17527 16083 17533
rect 16025 17524 16037 17527
rect 15804 17496 16037 17524
rect 15804 17484 15810 17496
rect 16025 17493 16037 17496
rect 16071 17493 16083 17527
rect 16025 17487 16083 17493
rect 19058 17484 19064 17536
rect 19116 17524 19122 17536
rect 22830 17524 22836 17536
rect 19116 17496 22836 17524
rect 19116 17484 19122 17496
rect 22830 17484 22836 17496
rect 22888 17484 22894 17536
rect 23017 17527 23075 17533
rect 23017 17493 23029 17527
rect 23063 17524 23075 17527
rect 23382 17524 23388 17536
rect 23063 17496 23388 17524
rect 23063 17493 23075 17496
rect 23017 17487 23075 17493
rect 23382 17484 23388 17496
rect 23440 17484 23446 17536
rect 23842 17484 23848 17536
rect 23900 17524 23906 17536
rect 24949 17527 25007 17533
rect 24949 17524 24961 17527
rect 23900 17496 24961 17524
rect 23900 17484 23906 17496
rect 24949 17493 24961 17496
rect 24995 17493 25007 17527
rect 24949 17487 25007 17493
rect 25406 17484 25412 17536
rect 25464 17524 25470 17536
rect 26602 17524 26608 17536
rect 25464 17496 26608 17524
rect 25464 17484 25470 17496
rect 26602 17484 26608 17496
rect 26660 17524 26666 17536
rect 30944 17524 30972 17700
rect 31389 17697 31401 17700
rect 31435 17697 31447 17731
rect 32306 17728 32312 17740
rect 32267 17700 32312 17728
rect 31389 17691 31447 17697
rect 32306 17688 32312 17700
rect 32364 17688 32370 17740
rect 32585 17731 32643 17737
rect 32585 17697 32597 17731
rect 32631 17728 32643 17731
rect 32674 17728 32680 17740
rect 32631 17700 32680 17728
rect 32631 17697 32643 17700
rect 32585 17691 32643 17697
rect 32674 17688 32680 17700
rect 32732 17688 32738 17740
rect 34790 17688 34796 17740
rect 34848 17728 34854 17740
rect 35253 17731 35311 17737
rect 35253 17728 35265 17731
rect 34848 17700 35265 17728
rect 34848 17688 34854 17700
rect 35253 17697 35265 17700
rect 35299 17697 35311 17731
rect 35253 17691 35311 17697
rect 35437 17731 35495 17737
rect 35437 17697 35449 17731
rect 35483 17728 35495 17731
rect 35526 17728 35532 17740
rect 35483 17700 35532 17728
rect 35483 17697 35495 17700
rect 35437 17691 35495 17697
rect 35526 17688 35532 17700
rect 35584 17688 35590 17740
rect 35894 17688 35900 17740
rect 35952 17728 35958 17740
rect 35989 17731 36047 17737
rect 35989 17728 36001 17731
rect 35952 17700 36001 17728
rect 35952 17688 35958 17700
rect 35989 17697 36001 17700
rect 36035 17728 36047 17731
rect 36630 17728 36636 17740
rect 36035 17700 36636 17728
rect 36035 17697 36047 17700
rect 35989 17691 36047 17697
rect 36630 17688 36636 17700
rect 36688 17688 36694 17740
rect 36722 17688 36728 17740
rect 36780 17728 36786 17740
rect 37737 17731 37795 17737
rect 36780 17700 36825 17728
rect 36780 17688 36786 17700
rect 37737 17697 37749 17731
rect 37783 17697 37795 17731
rect 37737 17691 37795 17697
rect 38289 17731 38347 17737
rect 38289 17697 38301 17731
rect 38335 17728 38347 17731
rect 38654 17728 38660 17740
rect 38335 17700 38660 17728
rect 38335 17697 38347 17700
rect 38289 17691 38347 17697
rect 31205 17663 31263 17669
rect 31205 17629 31217 17663
rect 31251 17660 31263 17663
rect 31754 17660 31760 17672
rect 31251 17632 31760 17660
rect 31251 17629 31263 17632
rect 31205 17623 31263 17629
rect 31754 17620 31760 17632
rect 31812 17620 31818 17672
rect 34146 17620 34152 17672
rect 34204 17660 34210 17672
rect 34425 17663 34483 17669
rect 34425 17660 34437 17663
rect 34204 17632 34437 17660
rect 34204 17620 34210 17632
rect 34425 17629 34437 17632
rect 34471 17629 34483 17663
rect 34425 17623 34483 17629
rect 34698 17620 34704 17672
rect 34756 17660 34762 17672
rect 34977 17663 35035 17669
rect 34977 17660 34989 17663
rect 34756 17632 34989 17660
rect 34756 17620 34762 17632
rect 34977 17629 34989 17632
rect 35023 17629 35035 17663
rect 37752 17660 37780 17691
rect 38654 17688 38660 17700
rect 38712 17688 38718 17740
rect 38930 17728 38936 17740
rect 38891 17700 38936 17728
rect 38930 17688 38936 17700
rect 38988 17688 38994 17740
rect 34977 17623 35035 17629
rect 36372 17632 37780 17660
rect 36372 17604 36400 17632
rect 36173 17595 36231 17601
rect 36173 17561 36185 17595
rect 36219 17592 36231 17595
rect 36354 17592 36360 17604
rect 36219 17564 36360 17592
rect 36219 17561 36231 17564
rect 36173 17555 36231 17561
rect 36354 17552 36360 17564
rect 36412 17552 36418 17604
rect 26660 17496 30972 17524
rect 26660 17484 26666 17496
rect 32766 17484 32772 17536
rect 32824 17524 32830 17536
rect 37458 17524 37464 17536
rect 32824 17496 37464 17524
rect 32824 17484 32830 17496
rect 37458 17484 37464 17496
rect 37516 17484 37522 17536
rect 1104 17434 39836 17456
rect 1104 17382 4246 17434
rect 4298 17382 4310 17434
rect 4362 17382 4374 17434
rect 4426 17382 4438 17434
rect 4490 17382 34966 17434
rect 35018 17382 35030 17434
rect 35082 17382 35094 17434
rect 35146 17382 35158 17434
rect 35210 17382 39836 17434
rect 1104 17360 39836 17382
rect 2777 17323 2835 17329
rect 2777 17289 2789 17323
rect 2823 17320 2835 17323
rect 2866 17320 2872 17332
rect 2823 17292 2872 17320
rect 2823 17289 2835 17292
rect 2777 17283 2835 17289
rect 2866 17280 2872 17292
rect 2924 17280 2930 17332
rect 5905 17323 5963 17329
rect 5905 17320 5917 17323
rect 4448 17292 5917 17320
rect 1394 17184 1400 17196
rect 1355 17156 1400 17184
rect 1394 17144 1400 17156
rect 1452 17144 1458 17196
rect 1673 17187 1731 17193
rect 1673 17153 1685 17187
rect 1719 17184 1731 17187
rect 4448 17184 4476 17292
rect 5905 17289 5917 17292
rect 5951 17289 5963 17323
rect 8846 17320 8852 17332
rect 8807 17292 8852 17320
rect 5905 17283 5963 17289
rect 8846 17280 8852 17292
rect 8904 17280 8910 17332
rect 9030 17280 9036 17332
rect 9088 17320 9094 17332
rect 9088 17292 15792 17320
rect 9088 17280 9094 17292
rect 9769 17255 9827 17261
rect 9769 17221 9781 17255
rect 9815 17252 9827 17255
rect 15764 17252 15792 17292
rect 15838 17280 15844 17332
rect 15896 17320 15902 17332
rect 16117 17323 16175 17329
rect 16117 17320 16129 17323
rect 15896 17292 16129 17320
rect 15896 17280 15902 17292
rect 16117 17289 16129 17292
rect 16163 17289 16175 17323
rect 16117 17283 16175 17289
rect 16206 17280 16212 17332
rect 16264 17320 16270 17332
rect 26142 17320 26148 17332
rect 16264 17292 26148 17320
rect 16264 17280 16270 17292
rect 26142 17280 26148 17292
rect 26200 17280 26206 17332
rect 26421 17323 26479 17329
rect 26421 17289 26433 17323
rect 26467 17320 26479 17323
rect 32766 17320 32772 17332
rect 26467 17292 32772 17320
rect 26467 17289 26479 17292
rect 26421 17283 26479 17289
rect 32766 17280 32772 17292
rect 32824 17280 32830 17332
rect 32950 17280 32956 17332
rect 33008 17320 33014 17332
rect 33045 17323 33103 17329
rect 33045 17320 33057 17323
rect 33008 17292 33057 17320
rect 33008 17280 33014 17292
rect 33045 17289 33057 17292
rect 33091 17289 33103 17323
rect 33045 17283 33103 17289
rect 34977 17323 35035 17329
rect 34977 17289 34989 17323
rect 35023 17320 35035 17323
rect 35434 17320 35440 17332
rect 35023 17292 35440 17320
rect 35023 17289 35035 17292
rect 34977 17283 35035 17289
rect 35434 17280 35440 17292
rect 35492 17280 35498 17332
rect 38930 17320 38936 17332
rect 36464 17292 38936 17320
rect 17405 17255 17463 17261
rect 9815 17224 11560 17252
rect 15764 17224 15976 17252
rect 9815 17221 9827 17224
rect 9769 17215 9827 17221
rect 1719 17156 4476 17184
rect 1719 17153 1731 17156
rect 1673 17147 1731 17153
rect 4706 17144 4712 17196
rect 4764 17184 4770 17196
rect 5074 17184 5080 17196
rect 4764 17156 5080 17184
rect 4764 17144 4770 17156
rect 5074 17144 5080 17156
rect 5132 17184 5138 17196
rect 5629 17187 5687 17193
rect 5629 17184 5641 17187
rect 5132 17156 5641 17184
rect 5132 17144 5138 17156
rect 5629 17153 5641 17156
rect 5675 17153 5687 17187
rect 5629 17147 5687 17153
rect 6822 17144 6828 17196
rect 6880 17184 6886 17196
rect 7285 17187 7343 17193
rect 7285 17184 7297 17187
rect 6880 17156 7297 17184
rect 6880 17144 6886 17156
rect 7285 17153 7297 17156
rect 7331 17153 7343 17187
rect 7285 17147 7343 17153
rect 1412 17116 1440 17144
rect 11532 17128 11560 17224
rect 12434 17184 12440 17196
rect 12395 17156 12440 17184
rect 12434 17144 12440 17156
rect 12492 17144 12498 17196
rect 12710 17184 12716 17196
rect 12671 17156 12716 17184
rect 12710 17144 12716 17156
rect 12768 17144 12774 17196
rect 13814 17144 13820 17196
rect 13872 17184 13878 17196
rect 14737 17187 14795 17193
rect 14737 17184 14749 17187
rect 13872 17156 14749 17184
rect 13872 17144 13878 17156
rect 14737 17153 14749 17156
rect 14783 17184 14795 17187
rect 15470 17184 15476 17196
rect 14783 17156 15476 17184
rect 14783 17153 14795 17156
rect 14737 17147 14795 17153
rect 15470 17144 15476 17156
rect 15528 17144 15534 17196
rect 2498 17116 2504 17128
rect 1412 17088 2504 17116
rect 2498 17076 2504 17088
rect 2556 17116 2562 17128
rect 3513 17119 3571 17125
rect 3513 17116 3525 17119
rect 2556 17088 3525 17116
rect 2556 17076 2562 17088
rect 3513 17085 3525 17088
rect 3559 17085 3571 17119
rect 3513 17079 3571 17085
rect 3789 17119 3847 17125
rect 3789 17085 3801 17119
rect 3835 17116 3847 17119
rect 5534 17116 5540 17128
rect 3835 17088 5540 17116
rect 3835 17085 3847 17088
rect 3789 17079 3847 17085
rect 5534 17076 5540 17088
rect 5592 17076 5598 17128
rect 5721 17119 5779 17125
rect 5721 17085 5733 17119
rect 5767 17085 5779 17119
rect 7558 17116 7564 17128
rect 7519 17088 7564 17116
rect 5721 17079 5779 17085
rect 5169 17051 5227 17057
rect 5169 17017 5181 17051
rect 5215 17048 5227 17051
rect 5736 17048 5764 17079
rect 7558 17076 7564 17088
rect 7616 17076 7622 17128
rect 8570 17076 8576 17128
rect 8628 17116 8634 17128
rect 9585 17119 9643 17125
rect 9585 17116 9597 17119
rect 8628 17088 9597 17116
rect 8628 17076 8634 17088
rect 9585 17085 9597 17088
rect 9631 17085 9643 17119
rect 9585 17079 9643 17085
rect 10689 17119 10747 17125
rect 10689 17085 10701 17119
rect 10735 17085 10747 17119
rect 10689 17079 10747 17085
rect 10965 17119 11023 17125
rect 10965 17085 10977 17119
rect 11011 17085 11023 17119
rect 10965 17079 11023 17085
rect 5215 17020 5764 17048
rect 5215 17017 5227 17020
rect 5169 17011 5227 17017
rect 10704 16992 10732 17079
rect 10980 17048 11008 17079
rect 11514 17076 11520 17128
rect 11572 17116 11578 17128
rect 11609 17119 11667 17125
rect 11609 17116 11621 17119
rect 11572 17088 11621 17116
rect 11572 17076 11578 17088
rect 11609 17085 11621 17088
rect 11655 17085 11667 17119
rect 11609 17079 11667 17085
rect 11790 17076 11796 17128
rect 11848 17076 11854 17128
rect 15013 17119 15071 17125
rect 15013 17085 15025 17119
rect 15059 17116 15071 17119
rect 15059 17088 15884 17116
rect 15059 17085 15071 17088
rect 15013 17079 15071 17085
rect 11808 17048 11836 17076
rect 10980 17020 11836 17048
rect 10505 16983 10563 16989
rect 10505 16949 10517 16983
rect 10551 16980 10563 16983
rect 10594 16980 10600 16992
rect 10551 16952 10600 16980
rect 10551 16949 10563 16952
rect 10505 16943 10563 16949
rect 10594 16940 10600 16952
rect 10652 16940 10658 16992
rect 10686 16940 10692 16992
rect 10744 16980 10750 16992
rect 11793 16983 11851 16989
rect 11793 16980 11805 16983
rect 10744 16952 11805 16980
rect 10744 16940 10750 16952
rect 11793 16949 11805 16952
rect 11839 16949 11851 16983
rect 13814 16980 13820 16992
rect 13775 16952 13820 16980
rect 11793 16943 11851 16949
rect 13814 16940 13820 16952
rect 13872 16940 13878 16992
rect 15856 16980 15884 17088
rect 15948 17048 15976 17224
rect 17405 17221 17417 17255
rect 17451 17252 17463 17255
rect 19058 17252 19064 17264
rect 17451 17224 19064 17252
rect 17451 17221 17463 17224
rect 17405 17215 17463 17221
rect 19058 17212 19064 17224
rect 19116 17212 19122 17264
rect 19426 17212 19432 17264
rect 19484 17252 19490 17264
rect 19521 17255 19579 17261
rect 19521 17252 19533 17255
rect 19484 17224 19533 17252
rect 19484 17212 19490 17224
rect 19521 17221 19533 17224
rect 19567 17221 19579 17255
rect 19521 17215 19579 17221
rect 19702 17212 19708 17264
rect 19760 17252 19766 17264
rect 28994 17252 29000 17264
rect 19760 17224 22048 17252
rect 19760 17212 19766 17224
rect 16114 17144 16120 17196
rect 16172 17184 16178 17196
rect 18509 17187 18567 17193
rect 18509 17184 18521 17187
rect 16172 17156 18521 17184
rect 16172 17144 16178 17156
rect 18509 17153 18521 17156
rect 18555 17153 18567 17187
rect 22020 17184 22048 17224
rect 24964 17224 29000 17252
rect 24964 17184 24992 17224
rect 28994 17212 29000 17224
rect 29052 17212 29058 17264
rect 32582 17252 32588 17264
rect 29472 17224 32588 17252
rect 26142 17184 26148 17196
rect 18509 17147 18567 17153
rect 18616 17156 19932 17184
rect 17310 17116 17316 17128
rect 17271 17088 17316 17116
rect 17310 17076 17316 17088
rect 17368 17076 17374 17128
rect 18322 17116 18328 17128
rect 18283 17088 18328 17116
rect 18322 17076 18328 17088
rect 18380 17076 18386 17128
rect 18616 17125 18644 17156
rect 18601 17119 18659 17125
rect 18601 17085 18613 17119
rect 18647 17085 18659 17119
rect 18601 17079 18659 17085
rect 19334 17076 19340 17128
rect 19392 17116 19398 17128
rect 19904 17125 19932 17156
rect 22020 17156 24992 17184
rect 26103 17156 26148 17184
rect 19429 17119 19487 17125
rect 19429 17116 19441 17119
rect 19392 17088 19441 17116
rect 19392 17076 19398 17088
rect 19429 17085 19441 17088
rect 19475 17085 19487 17119
rect 19429 17079 19487 17085
rect 19889 17119 19947 17125
rect 19889 17085 19901 17119
rect 19935 17116 19947 17119
rect 19978 17116 19984 17128
rect 19935 17088 19984 17116
rect 19935 17085 19947 17088
rect 19889 17079 19947 17085
rect 19978 17076 19984 17088
rect 20036 17076 20042 17128
rect 20070 17076 20076 17128
rect 20128 17116 20134 17128
rect 20165 17119 20223 17125
rect 20165 17116 20177 17119
rect 20128 17088 20177 17116
rect 20128 17076 20134 17088
rect 20165 17085 20177 17088
rect 20211 17085 20223 17119
rect 20714 17116 20720 17128
rect 20675 17088 20720 17116
rect 20165 17079 20223 17085
rect 20714 17076 20720 17088
rect 20772 17076 20778 17128
rect 21266 17116 21272 17128
rect 21227 17088 21272 17116
rect 21266 17076 21272 17088
rect 21324 17076 21330 17128
rect 22020 17125 22048 17156
rect 26142 17144 26148 17156
rect 26200 17144 26206 17196
rect 27246 17144 27252 17196
rect 27304 17184 27310 17196
rect 27433 17187 27491 17193
rect 27433 17184 27445 17187
rect 27304 17156 27445 17184
rect 27304 17144 27310 17156
rect 27433 17153 27445 17156
rect 27479 17153 27491 17187
rect 27798 17184 27804 17196
rect 27433 17147 27491 17153
rect 27724 17156 27804 17184
rect 22005 17119 22063 17125
rect 22005 17085 22017 17119
rect 22051 17085 22063 17119
rect 22830 17116 22836 17128
rect 22791 17088 22836 17116
rect 22005 17079 22063 17085
rect 22830 17076 22836 17088
rect 22888 17076 22894 17128
rect 24026 17116 24032 17128
rect 23987 17088 24032 17116
rect 24026 17076 24032 17088
rect 24084 17076 24090 17128
rect 24302 17116 24308 17128
rect 24263 17088 24308 17116
rect 24302 17076 24308 17088
rect 24360 17076 24366 17128
rect 26237 17119 26295 17125
rect 26237 17085 26249 17119
rect 26283 17085 26295 17119
rect 27614 17116 27620 17128
rect 27575 17088 27620 17116
rect 26237 17079 26295 17085
rect 25685 17051 25743 17057
rect 15948 17020 23980 17048
rect 17218 16980 17224 16992
rect 15856 16952 17224 16980
rect 17218 16940 17224 16952
rect 17276 16940 17282 16992
rect 21266 16940 21272 16992
rect 21324 16980 21330 16992
rect 22186 16980 22192 16992
rect 21324 16952 22192 16980
rect 21324 16940 21330 16952
rect 22186 16940 22192 16952
rect 22244 16940 22250 16992
rect 22554 16940 22560 16992
rect 22612 16980 22618 16992
rect 23017 16983 23075 16989
rect 23017 16980 23029 16983
rect 22612 16952 23029 16980
rect 22612 16940 22618 16952
rect 23017 16949 23029 16952
rect 23063 16949 23075 16983
rect 23952 16980 23980 17020
rect 25685 17017 25697 17051
rect 25731 17048 25743 17051
rect 26252 17048 26280 17079
rect 27614 17076 27620 17088
rect 27672 17076 27678 17128
rect 27724 17125 27752 17156
rect 27798 17144 27804 17156
rect 27856 17144 27862 17196
rect 29472 17125 29500 17224
rect 32582 17212 32588 17224
rect 32640 17212 32646 17264
rect 29546 17144 29552 17196
rect 29604 17184 29610 17196
rect 32030 17184 32036 17196
rect 29604 17156 32036 17184
rect 29604 17144 29610 17156
rect 27709 17119 27767 17125
rect 27709 17085 27721 17119
rect 27755 17085 27767 17119
rect 27709 17079 27767 17085
rect 29457 17119 29515 17125
rect 29457 17085 29469 17119
rect 29503 17085 29515 17119
rect 29457 17079 29515 17085
rect 30193 17119 30251 17125
rect 30193 17085 30205 17119
rect 30239 17116 30251 17119
rect 30374 17116 30380 17128
rect 30239 17088 30380 17116
rect 30239 17085 30251 17088
rect 30193 17079 30251 17085
rect 30374 17076 30380 17088
rect 30432 17076 30438 17128
rect 30650 17116 30656 17128
rect 30611 17088 30656 17116
rect 30650 17076 30656 17088
rect 30708 17076 30714 17128
rect 31294 17116 31300 17128
rect 31255 17088 31300 17116
rect 31294 17076 31300 17088
rect 31352 17076 31358 17128
rect 31404 17125 31432 17156
rect 32030 17144 32036 17156
rect 32088 17144 32094 17196
rect 33042 17144 33048 17196
rect 33100 17184 33106 17196
rect 35710 17184 35716 17196
rect 33100 17156 35716 17184
rect 33100 17144 33106 17156
rect 31389 17119 31447 17125
rect 31389 17085 31401 17119
rect 31435 17085 31447 17119
rect 31389 17079 31447 17085
rect 31754 17076 31760 17128
rect 31812 17116 31818 17128
rect 32048 17116 32076 17144
rect 32953 17119 33011 17125
rect 32953 17116 32965 17119
rect 31812 17088 31857 17116
rect 32048 17088 32965 17116
rect 31812 17076 31818 17088
rect 32953 17085 32965 17088
rect 32999 17085 33011 17119
rect 33778 17116 33784 17128
rect 33739 17088 33784 17116
rect 32953 17079 33011 17085
rect 33778 17076 33784 17088
rect 33836 17076 33842 17128
rect 34146 17116 34152 17128
rect 34107 17088 34152 17116
rect 34146 17076 34152 17088
rect 34204 17076 34210 17128
rect 34790 17076 34796 17128
rect 34848 17116 34854 17128
rect 35544 17125 35572 17156
rect 35710 17144 35716 17156
rect 35768 17144 35774 17196
rect 36464 17184 36492 17292
rect 38930 17280 38936 17292
rect 38988 17280 38994 17332
rect 38470 17212 38476 17264
rect 38528 17252 38534 17264
rect 38841 17255 38899 17261
rect 38841 17252 38853 17255
rect 38528 17224 38853 17252
rect 38528 17212 38534 17224
rect 38841 17221 38853 17224
rect 38887 17221 38899 17255
rect 38841 17215 38899 17221
rect 38194 17184 38200 17196
rect 36188 17156 36492 17184
rect 36556 17156 38200 17184
rect 36188 17125 36216 17156
rect 36556 17125 36584 17156
rect 38194 17144 38200 17156
rect 38252 17144 38258 17196
rect 34885 17119 34943 17125
rect 34885 17116 34897 17119
rect 34848 17088 34897 17116
rect 34848 17076 34854 17088
rect 34885 17085 34897 17088
rect 34931 17085 34943 17119
rect 34885 17079 34943 17085
rect 35529 17119 35587 17125
rect 35529 17085 35541 17119
rect 35575 17085 35587 17119
rect 35529 17079 35587 17085
rect 36173 17119 36231 17125
rect 36173 17085 36185 17119
rect 36219 17085 36231 17119
rect 36173 17079 36231 17085
rect 36541 17119 36599 17125
rect 36541 17085 36553 17119
rect 36587 17085 36599 17119
rect 36541 17079 36599 17085
rect 36909 17119 36967 17125
rect 36909 17085 36921 17119
rect 36955 17116 36967 17119
rect 36955 17088 37412 17116
rect 36955 17085 36967 17088
rect 36909 17079 36967 17085
rect 25731 17020 26280 17048
rect 27801 17051 27859 17057
rect 25731 17017 25743 17020
rect 25685 17011 25743 17017
rect 27801 17017 27813 17051
rect 27847 17048 27859 17051
rect 27890 17048 27896 17060
rect 27847 17020 27896 17048
rect 27847 17017 27859 17020
rect 27801 17011 27859 17017
rect 27890 17008 27896 17020
rect 27948 17008 27954 17060
rect 28169 17051 28227 17057
rect 28169 17017 28181 17051
rect 28215 17048 28227 17051
rect 30282 17048 30288 17060
rect 28215 17020 30288 17048
rect 28215 17017 28227 17020
rect 28169 17011 28227 17017
rect 30282 17008 30288 17020
rect 30340 17008 30346 17060
rect 30466 17048 30472 17060
rect 30427 17020 30472 17048
rect 30466 17008 30472 17020
rect 30524 17008 30530 17060
rect 34333 17051 34391 17057
rect 34333 17017 34345 17051
rect 34379 17048 34391 17051
rect 36262 17048 36268 17060
rect 34379 17020 36268 17048
rect 34379 17017 34391 17020
rect 34333 17011 34391 17017
rect 36262 17008 36268 17020
rect 36320 17008 36326 17060
rect 24946 16980 24952 16992
rect 23952 16952 24952 16980
rect 23017 16943 23075 16949
rect 24946 16940 24952 16952
rect 25004 16940 25010 16992
rect 26418 16940 26424 16992
rect 26476 16980 26482 16992
rect 26786 16980 26792 16992
rect 26476 16952 26792 16980
rect 26476 16940 26482 16952
rect 26786 16940 26792 16952
rect 26844 16940 26850 16992
rect 28258 16940 28264 16992
rect 28316 16980 28322 16992
rect 28810 16980 28816 16992
rect 28316 16952 28816 16980
rect 28316 16940 28322 16952
rect 28810 16940 28816 16952
rect 28868 16940 28874 16992
rect 29549 16983 29607 16989
rect 29549 16949 29561 16983
rect 29595 16980 29607 16983
rect 32122 16980 32128 16992
rect 29595 16952 32128 16980
rect 29595 16949 29607 16952
rect 29549 16943 29607 16949
rect 32122 16940 32128 16952
rect 32180 16940 32186 16992
rect 34054 16940 34060 16992
rect 34112 16980 34118 16992
rect 36170 16980 36176 16992
rect 34112 16952 36176 16980
rect 34112 16940 34118 16952
rect 36170 16940 36176 16952
rect 36228 16940 36234 16992
rect 36354 16940 36360 16992
rect 36412 16980 36418 16992
rect 36725 16983 36783 16989
rect 36725 16980 36737 16983
rect 36412 16952 36737 16980
rect 36412 16940 36418 16952
rect 36725 16949 36737 16952
rect 36771 16949 36783 16983
rect 37384 16980 37412 17088
rect 37458 17076 37464 17128
rect 37516 17116 37522 17128
rect 37737 17119 37795 17125
rect 37516 17088 37561 17116
rect 37516 17076 37522 17088
rect 37737 17085 37749 17119
rect 37783 17116 37795 17119
rect 38562 17116 38568 17128
rect 37783 17088 38568 17116
rect 37783 17085 37795 17088
rect 37737 17079 37795 17085
rect 38562 17076 38568 17088
rect 38620 17076 38626 17128
rect 38654 16980 38660 16992
rect 37384 16952 38660 16980
rect 36725 16943 36783 16949
rect 38654 16940 38660 16952
rect 38712 16940 38718 16992
rect 1104 16890 39836 16912
rect 1104 16838 19606 16890
rect 19658 16838 19670 16890
rect 19722 16838 19734 16890
rect 19786 16838 19798 16890
rect 19850 16838 39836 16890
rect 1104 16816 39836 16838
rect 1946 16776 1952 16788
rect 1907 16748 1952 16776
rect 1946 16736 1952 16748
rect 2004 16736 2010 16788
rect 2498 16776 2504 16788
rect 2459 16748 2504 16776
rect 2498 16736 2504 16748
rect 2556 16736 2562 16788
rect 5258 16776 5264 16788
rect 2700 16748 4200 16776
rect 5219 16748 5264 16776
rect 1762 16640 1768 16652
rect 1723 16612 1768 16640
rect 1762 16600 1768 16612
rect 1820 16600 1826 16652
rect 2700 16649 2728 16748
rect 4172 16708 4200 16748
rect 5258 16736 5264 16748
rect 5316 16736 5322 16788
rect 6365 16779 6423 16785
rect 6365 16745 6377 16779
rect 6411 16745 6423 16779
rect 10686 16776 10692 16788
rect 6365 16739 6423 16745
rect 6840 16748 10692 16776
rect 6270 16708 6276 16720
rect 4172 16680 6276 16708
rect 6270 16668 6276 16680
rect 6328 16708 6334 16720
rect 6380 16708 6408 16739
rect 6328 16680 6408 16708
rect 6328 16668 6334 16680
rect 2685 16643 2743 16649
rect 2685 16609 2697 16643
rect 2731 16609 2743 16643
rect 2685 16603 2743 16609
rect 4157 16643 4215 16649
rect 4157 16609 4169 16643
rect 4203 16640 4215 16643
rect 4614 16640 4620 16652
rect 4203 16612 4620 16640
rect 4203 16609 4215 16612
rect 4157 16603 4215 16609
rect 4614 16600 4620 16612
rect 4672 16600 4678 16652
rect 4706 16600 4712 16652
rect 4764 16600 4770 16652
rect 5353 16643 5411 16649
rect 5353 16609 5365 16643
rect 5399 16609 5411 16643
rect 5718 16640 5724 16652
rect 5679 16612 5724 16640
rect 5353 16603 5411 16609
rect 4065 16575 4123 16581
rect 4065 16541 4077 16575
rect 4111 16572 4123 16575
rect 4724 16572 4752 16600
rect 4111 16544 4752 16572
rect 4111 16541 4123 16544
rect 4065 16535 4123 16541
rect 5368 16516 5396 16603
rect 5718 16600 5724 16612
rect 5776 16600 5782 16652
rect 6546 16640 6552 16652
rect 6507 16612 6552 16640
rect 6546 16600 6552 16612
rect 6604 16600 6610 16652
rect 6840 16649 6868 16748
rect 10686 16736 10692 16748
rect 10744 16736 10750 16788
rect 11517 16779 11575 16785
rect 11517 16745 11529 16779
rect 11563 16745 11575 16779
rect 11517 16739 11575 16745
rect 7377 16711 7435 16717
rect 7377 16677 7389 16711
rect 7423 16708 7435 16711
rect 7558 16708 7564 16720
rect 7423 16680 7564 16708
rect 7423 16677 7435 16680
rect 7377 16671 7435 16677
rect 7558 16668 7564 16680
rect 7616 16668 7622 16720
rect 9030 16708 9036 16720
rect 8220 16680 9036 16708
rect 6825 16643 6883 16649
rect 6825 16640 6837 16643
rect 6656 16612 6837 16640
rect 5350 16504 5356 16516
rect 5263 16476 5356 16504
rect 5350 16464 5356 16476
rect 5408 16504 5414 16516
rect 6656 16504 6684 16612
rect 6825 16609 6837 16612
rect 6871 16609 6883 16643
rect 6825 16603 6883 16609
rect 7193 16643 7251 16649
rect 7193 16609 7205 16643
rect 7239 16640 7251 16643
rect 7282 16640 7288 16652
rect 7239 16612 7288 16640
rect 7239 16609 7251 16612
rect 7193 16603 7251 16609
rect 7282 16600 7288 16612
rect 7340 16600 7346 16652
rect 8220 16649 8248 16680
rect 9030 16668 9036 16680
rect 9088 16668 9094 16720
rect 10870 16708 10876 16720
rect 9968 16680 10876 16708
rect 9968 16649 9996 16680
rect 10870 16668 10876 16680
rect 10928 16708 10934 16720
rect 11532 16708 11560 16739
rect 11790 16736 11796 16788
rect 11848 16776 11854 16788
rect 14645 16779 14703 16785
rect 14645 16776 14657 16779
rect 11848 16748 14657 16776
rect 11848 16736 11854 16748
rect 14645 16745 14657 16748
rect 14691 16745 14703 16779
rect 14645 16739 14703 16745
rect 15473 16779 15531 16785
rect 15473 16745 15485 16779
rect 15519 16776 15531 16779
rect 15654 16776 15660 16788
rect 15519 16748 15660 16776
rect 15519 16745 15531 16748
rect 15473 16739 15531 16745
rect 15654 16736 15660 16748
rect 15712 16776 15718 16788
rect 15838 16776 15844 16788
rect 15712 16748 15844 16776
rect 15712 16736 15718 16748
rect 15838 16736 15844 16748
rect 15896 16736 15902 16788
rect 16206 16776 16212 16788
rect 16167 16748 16212 16776
rect 16206 16736 16212 16748
rect 16264 16736 16270 16788
rect 19978 16736 19984 16788
rect 20036 16776 20042 16788
rect 20257 16779 20315 16785
rect 20257 16776 20269 16779
rect 20036 16748 20269 16776
rect 20036 16736 20042 16748
rect 20257 16745 20269 16748
rect 20303 16745 20315 16779
rect 23566 16776 23572 16788
rect 20257 16739 20315 16745
rect 21744 16748 23572 16776
rect 10928 16680 11560 16708
rect 10928 16668 10934 16680
rect 13814 16668 13820 16720
rect 13872 16708 13878 16720
rect 21744 16708 21772 16748
rect 23566 16736 23572 16748
rect 23624 16736 23630 16788
rect 26786 16736 26792 16788
rect 26844 16776 26850 16788
rect 30834 16776 30840 16788
rect 26844 16748 30840 16776
rect 26844 16736 26850 16748
rect 30834 16736 30840 16748
rect 30892 16736 30898 16788
rect 31205 16779 31263 16785
rect 31205 16745 31217 16779
rect 31251 16776 31263 16779
rect 31754 16776 31760 16788
rect 31251 16748 31760 16776
rect 31251 16745 31263 16748
rect 31205 16739 31263 16745
rect 31754 16736 31760 16748
rect 31812 16736 31818 16788
rect 32309 16779 32367 16785
rect 32309 16745 32321 16779
rect 32355 16745 32367 16779
rect 32309 16739 32367 16745
rect 33137 16779 33195 16785
rect 33137 16745 33149 16779
rect 33183 16776 33195 16779
rect 33410 16776 33416 16788
rect 33183 16748 33416 16776
rect 33183 16745 33195 16748
rect 33137 16739 33195 16745
rect 13872 16680 14596 16708
rect 13872 16668 13878 16680
rect 8205 16643 8263 16649
rect 8205 16609 8217 16643
rect 8251 16609 8263 16643
rect 8389 16643 8447 16649
rect 8389 16640 8401 16643
rect 8205 16603 8263 16609
rect 8312 16612 8401 16640
rect 8110 16532 8116 16584
rect 8168 16572 8174 16584
rect 8312 16572 8340 16612
rect 8389 16609 8401 16612
rect 8435 16609 8447 16643
rect 8389 16603 8447 16609
rect 8941 16643 8999 16649
rect 8941 16609 8953 16643
rect 8987 16640 8999 16643
rect 9953 16643 10011 16649
rect 8987 16612 9628 16640
rect 8987 16609 8999 16612
rect 8941 16603 8999 16609
rect 9122 16572 9128 16584
rect 8168 16544 8340 16572
rect 9083 16544 9128 16572
rect 8168 16532 8174 16544
rect 9122 16532 9128 16544
rect 9180 16532 9186 16584
rect 9600 16572 9628 16612
rect 9953 16609 9965 16643
rect 9999 16609 10011 16643
rect 9953 16603 10011 16609
rect 10042 16600 10048 16652
rect 10100 16640 10106 16652
rect 10410 16640 10416 16652
rect 10100 16612 10145 16640
rect 10371 16612 10416 16640
rect 10100 16600 10106 16612
rect 10410 16600 10416 16612
rect 10468 16600 10474 16652
rect 11330 16640 11336 16652
rect 11291 16612 11336 16640
rect 11330 16600 11336 16612
rect 11388 16600 11394 16652
rect 12434 16640 12440 16652
rect 12395 16612 12440 16640
rect 12434 16600 12440 16612
rect 12492 16600 12498 16652
rect 12713 16643 12771 16649
rect 12713 16609 12725 16643
rect 12759 16640 12771 16643
rect 13998 16640 14004 16652
rect 12759 16612 14004 16640
rect 12759 16609 12771 16612
rect 12713 16603 12771 16609
rect 13998 16600 14004 16612
rect 14056 16600 14062 16652
rect 14568 16649 14596 16680
rect 21652 16680 21772 16708
rect 14553 16643 14611 16649
rect 14553 16609 14565 16643
rect 14599 16609 14611 16643
rect 15286 16640 15292 16652
rect 15247 16612 15292 16640
rect 14553 16603 14611 16609
rect 15286 16600 15292 16612
rect 15344 16640 15350 16652
rect 16025 16643 16083 16649
rect 16025 16640 16037 16643
rect 15344 16612 16037 16640
rect 15344 16600 15350 16612
rect 16025 16609 16037 16612
rect 16071 16609 16083 16643
rect 17034 16640 17040 16652
rect 16995 16612 17040 16640
rect 16025 16603 16083 16609
rect 17034 16600 17040 16612
rect 17092 16600 17098 16652
rect 19150 16640 19156 16652
rect 19111 16612 19156 16640
rect 19150 16600 19156 16612
rect 19208 16600 19214 16652
rect 20165 16643 20223 16649
rect 20165 16609 20177 16643
rect 20211 16640 20223 16643
rect 20346 16640 20352 16652
rect 20211 16612 20352 16640
rect 20211 16609 20223 16612
rect 20165 16603 20223 16609
rect 20346 16600 20352 16612
rect 20404 16600 20410 16652
rect 20530 16600 20536 16652
rect 20588 16640 20594 16652
rect 21652 16649 21680 16680
rect 22186 16668 22192 16720
rect 22244 16708 22250 16720
rect 27338 16708 27344 16720
rect 22244 16680 22692 16708
rect 22244 16668 22250 16680
rect 22664 16652 22692 16680
rect 27172 16680 27344 16708
rect 20993 16643 21051 16649
rect 20993 16640 21005 16643
rect 20588 16612 21005 16640
rect 20588 16600 20594 16612
rect 20993 16609 21005 16612
rect 21039 16609 21051 16643
rect 20993 16603 21051 16609
rect 21637 16643 21695 16649
rect 21637 16609 21649 16643
rect 21683 16609 21695 16643
rect 21910 16640 21916 16652
rect 21871 16612 21916 16640
rect 21637 16603 21695 16609
rect 21910 16600 21916 16612
rect 21968 16600 21974 16652
rect 22370 16640 22376 16652
rect 22331 16612 22376 16640
rect 22370 16600 22376 16612
rect 22428 16600 22434 16652
rect 22646 16640 22652 16652
rect 22559 16612 22652 16640
rect 22646 16600 22652 16612
rect 22704 16600 22710 16652
rect 23382 16640 23388 16652
rect 23343 16612 23388 16640
rect 23382 16600 23388 16612
rect 23440 16600 23446 16652
rect 23474 16600 23480 16652
rect 23532 16640 23538 16652
rect 24305 16643 24363 16649
rect 24305 16640 24317 16643
rect 23532 16612 24317 16640
rect 23532 16600 23538 16612
rect 24305 16609 24317 16612
rect 24351 16609 24363 16643
rect 24305 16603 24363 16609
rect 25685 16643 25743 16649
rect 25685 16609 25697 16643
rect 25731 16640 25743 16643
rect 26602 16640 26608 16652
rect 25731 16612 26608 16640
rect 25731 16609 25743 16612
rect 25685 16603 25743 16609
rect 26602 16600 26608 16612
rect 26660 16600 26666 16652
rect 26786 16640 26792 16652
rect 26747 16612 26792 16640
rect 26786 16600 26792 16612
rect 26844 16600 26850 16652
rect 27172 16649 27200 16680
rect 27338 16668 27344 16680
rect 27396 16668 27402 16720
rect 30852 16708 30880 16736
rect 32324 16708 32352 16739
rect 33410 16736 33416 16748
rect 33468 16736 33474 16788
rect 35989 16779 36047 16785
rect 33520 16748 35848 16776
rect 30852 16680 32352 16708
rect 27157 16643 27215 16649
rect 27157 16609 27169 16643
rect 27203 16609 27215 16643
rect 27157 16603 27215 16609
rect 27246 16600 27252 16652
rect 27304 16640 27310 16652
rect 27433 16643 27491 16649
rect 27433 16640 27445 16643
rect 27304 16612 27445 16640
rect 27304 16600 27310 16612
rect 27433 16609 27445 16612
rect 27479 16609 27491 16643
rect 27798 16640 27804 16652
rect 27759 16612 27804 16640
rect 27433 16603 27491 16609
rect 27798 16600 27804 16612
rect 27856 16600 27862 16652
rect 28258 16640 28264 16652
rect 28219 16612 28264 16640
rect 28258 16600 28264 16612
rect 28316 16600 28322 16652
rect 28626 16600 28632 16652
rect 28684 16640 28690 16652
rect 29181 16643 29239 16649
rect 29181 16640 29193 16643
rect 28684 16612 29193 16640
rect 28684 16600 28690 16612
rect 29181 16609 29193 16612
rect 29227 16609 29239 16643
rect 29181 16603 29239 16609
rect 30282 16600 30288 16652
rect 30340 16640 30346 16652
rect 31021 16643 31079 16649
rect 31021 16640 31033 16643
rect 30340 16612 31033 16640
rect 30340 16600 30346 16612
rect 31021 16609 31033 16612
rect 31067 16609 31079 16643
rect 31021 16603 31079 16609
rect 32125 16643 32183 16649
rect 32125 16609 32137 16643
rect 32171 16640 32183 16643
rect 32214 16640 32220 16652
rect 32171 16612 32220 16640
rect 32171 16609 32183 16612
rect 32125 16603 32183 16609
rect 32214 16600 32220 16612
rect 32272 16640 32278 16652
rect 32398 16640 32404 16652
rect 32272 16612 32404 16640
rect 32272 16600 32278 16612
rect 32398 16600 32404 16612
rect 32456 16600 32462 16652
rect 32953 16643 33011 16649
rect 32953 16609 32965 16643
rect 32999 16640 33011 16643
rect 33520 16640 33548 16748
rect 33686 16640 33692 16652
rect 32999 16612 33548 16640
rect 33647 16612 33692 16640
rect 32999 16609 33011 16612
rect 32953 16603 33011 16609
rect 33686 16600 33692 16612
rect 33744 16600 33750 16652
rect 33965 16643 34023 16649
rect 33965 16609 33977 16643
rect 34011 16640 34023 16643
rect 34606 16640 34612 16652
rect 34011 16612 34612 16640
rect 34011 16609 34023 16612
rect 33965 16603 34023 16609
rect 34606 16600 34612 16612
rect 34664 16600 34670 16652
rect 35820 16649 35848 16748
rect 35989 16745 36001 16779
rect 36035 16776 36047 16779
rect 36170 16776 36176 16788
rect 36035 16748 36176 16776
rect 36035 16745 36047 16748
rect 35989 16739 36047 16745
rect 36170 16736 36176 16748
rect 36228 16736 36234 16788
rect 38010 16736 38016 16788
rect 38068 16776 38074 16788
rect 38105 16779 38163 16785
rect 38105 16776 38117 16779
rect 38068 16748 38117 16776
rect 38068 16736 38074 16748
rect 38105 16745 38117 16748
rect 38151 16745 38163 16779
rect 38105 16739 38163 16745
rect 38197 16711 38255 16717
rect 38197 16677 38209 16711
rect 38243 16708 38255 16711
rect 38286 16708 38292 16720
rect 38243 16680 38292 16708
rect 38243 16677 38255 16680
rect 38197 16671 38255 16677
rect 38286 16668 38292 16680
rect 38344 16668 38350 16720
rect 38562 16708 38568 16720
rect 38523 16680 38568 16708
rect 38562 16668 38568 16680
rect 38620 16668 38626 16720
rect 35805 16643 35863 16649
rect 35805 16609 35817 16643
rect 35851 16640 35863 16643
rect 35894 16640 35900 16652
rect 35851 16612 35900 16640
rect 35851 16609 35863 16612
rect 35805 16603 35863 16609
rect 35894 16600 35900 16612
rect 35952 16600 35958 16652
rect 36630 16640 36636 16652
rect 36591 16612 36636 16640
rect 36630 16600 36636 16612
rect 36688 16600 36694 16652
rect 36814 16640 36820 16652
rect 36775 16612 36820 16640
rect 36814 16600 36820 16612
rect 36872 16600 36878 16652
rect 38013 16643 38071 16649
rect 38013 16609 38025 16643
rect 38059 16640 38071 16643
rect 38654 16640 38660 16652
rect 38059 16612 38660 16640
rect 38059 16609 38071 16612
rect 38013 16603 38071 16609
rect 38654 16600 38660 16612
rect 38712 16600 38718 16652
rect 9769 16575 9827 16581
rect 9769 16572 9781 16575
rect 9600 16544 9781 16572
rect 9769 16541 9781 16544
rect 9815 16541 9827 16575
rect 16758 16572 16764 16584
rect 16671 16544 16764 16572
rect 9769 16535 9827 16541
rect 16758 16532 16764 16544
rect 16816 16572 16822 16584
rect 17770 16572 17776 16584
rect 16816 16544 17776 16572
rect 16816 16532 16822 16544
rect 17770 16532 17776 16544
rect 17828 16532 17834 16584
rect 21818 16572 21824 16584
rect 21779 16544 21824 16572
rect 21818 16532 21824 16544
rect 21876 16532 21882 16584
rect 22462 16532 22468 16584
rect 22520 16572 22526 16584
rect 23290 16572 23296 16584
rect 22520 16544 23296 16572
rect 22520 16532 22526 16544
rect 23290 16532 23296 16544
rect 23348 16532 23354 16584
rect 24026 16572 24032 16584
rect 23987 16544 24032 16572
rect 24026 16532 24032 16544
rect 24084 16532 24090 16584
rect 26878 16572 26884 16584
rect 26839 16544 26884 16572
rect 26878 16532 26884 16544
rect 26936 16532 26942 16584
rect 28905 16575 28963 16581
rect 28905 16541 28917 16575
rect 28951 16572 28963 16575
rect 29086 16572 29092 16584
rect 28951 16544 29092 16572
rect 28951 16541 28963 16544
rect 28905 16535 28963 16541
rect 29086 16532 29092 16544
rect 29144 16572 29150 16584
rect 30098 16572 30104 16584
rect 29144 16544 30104 16572
rect 29144 16532 29150 16544
rect 30098 16532 30104 16544
rect 30156 16532 30162 16584
rect 37185 16575 37243 16581
rect 37185 16541 37197 16575
rect 37231 16572 37243 16575
rect 37550 16572 37556 16584
rect 37231 16544 37556 16572
rect 37231 16541 37243 16544
rect 37185 16535 37243 16541
rect 37550 16532 37556 16544
rect 37608 16532 37614 16584
rect 37829 16575 37887 16581
rect 37829 16541 37841 16575
rect 37875 16572 37887 16575
rect 38378 16572 38384 16584
rect 37875 16544 38384 16572
rect 37875 16541 37887 16544
rect 37829 16535 37887 16541
rect 38378 16532 38384 16544
rect 38436 16532 38442 16584
rect 23382 16504 23388 16516
rect 5408 16476 6684 16504
rect 13740 16476 16344 16504
rect 5408 16464 5414 16476
rect 4062 16396 4068 16448
rect 4120 16436 4126 16448
rect 4341 16439 4399 16445
rect 4341 16436 4353 16439
rect 4120 16408 4353 16436
rect 4120 16396 4126 16408
rect 4341 16405 4353 16408
rect 4387 16405 4399 16439
rect 4341 16399 4399 16405
rect 10042 16396 10048 16448
rect 10100 16436 10106 16448
rect 13740 16436 13768 16476
rect 10100 16408 13768 16436
rect 10100 16396 10106 16408
rect 13906 16396 13912 16448
rect 13964 16436 13970 16448
rect 14001 16439 14059 16445
rect 14001 16436 14013 16439
rect 13964 16408 14013 16436
rect 13964 16396 13970 16408
rect 14001 16405 14013 16408
rect 14047 16405 14059 16439
rect 16316 16436 16344 16476
rect 17696 16476 23388 16504
rect 17696 16436 17724 16476
rect 23382 16464 23388 16476
rect 23440 16464 23446 16516
rect 16316 16408 17724 16436
rect 14001 16399 14059 16405
rect 17954 16396 17960 16448
rect 18012 16436 18018 16448
rect 18141 16439 18199 16445
rect 18141 16436 18153 16439
rect 18012 16408 18153 16436
rect 18012 16396 18018 16408
rect 18141 16405 18153 16408
rect 18187 16405 18199 16439
rect 19334 16436 19340 16448
rect 19295 16408 19340 16436
rect 18141 16399 18199 16405
rect 19334 16396 19340 16408
rect 19392 16396 19398 16448
rect 19426 16396 19432 16448
rect 19484 16436 19490 16448
rect 21634 16436 21640 16448
rect 19484 16408 21640 16436
rect 19484 16396 19490 16408
rect 21634 16396 21640 16408
rect 21692 16396 21698 16448
rect 23477 16439 23535 16445
rect 23477 16405 23489 16439
rect 23523 16436 23535 16439
rect 23566 16436 23572 16448
rect 23523 16408 23572 16436
rect 23523 16405 23535 16408
rect 23477 16399 23535 16405
rect 23566 16396 23572 16408
rect 23624 16436 23630 16448
rect 24210 16436 24216 16448
rect 23624 16408 24216 16436
rect 23624 16396 23630 16408
rect 24210 16396 24216 16408
rect 24268 16396 24274 16448
rect 30282 16436 30288 16448
rect 30243 16408 30288 16436
rect 30282 16396 30288 16408
rect 30340 16396 30346 16448
rect 34790 16396 34796 16448
rect 34848 16436 34854 16448
rect 35069 16439 35127 16445
rect 35069 16436 35081 16439
rect 34848 16408 35081 16436
rect 34848 16396 34854 16408
rect 35069 16405 35081 16408
rect 35115 16405 35127 16439
rect 35069 16399 35127 16405
rect 1104 16346 39836 16368
rect 1104 16294 4246 16346
rect 4298 16294 4310 16346
rect 4362 16294 4374 16346
rect 4426 16294 4438 16346
rect 4490 16294 34966 16346
rect 35018 16294 35030 16346
rect 35082 16294 35094 16346
rect 35146 16294 35158 16346
rect 35210 16294 39836 16346
rect 1104 16272 39836 16294
rect 4525 16235 4583 16241
rect 4525 16201 4537 16235
rect 4571 16232 4583 16235
rect 4614 16232 4620 16244
rect 4571 16204 4620 16232
rect 4571 16201 4583 16204
rect 4525 16195 4583 16201
rect 4614 16192 4620 16204
rect 4672 16192 4678 16244
rect 10965 16235 11023 16241
rect 10965 16201 10977 16235
rect 11011 16232 11023 16235
rect 11330 16232 11336 16244
rect 11011 16204 11336 16232
rect 11011 16201 11023 16204
rect 10965 16195 11023 16201
rect 11330 16192 11336 16204
rect 11388 16192 11394 16244
rect 16853 16235 16911 16241
rect 16853 16201 16865 16235
rect 16899 16232 16911 16235
rect 18322 16232 18328 16244
rect 16899 16204 18328 16232
rect 16899 16201 16911 16204
rect 16853 16195 16911 16201
rect 18322 16192 18328 16204
rect 18380 16232 18386 16244
rect 18380 16204 22692 16232
rect 18380 16192 18386 16204
rect 7098 16164 7104 16176
rect 7059 16136 7104 16164
rect 7098 16124 7104 16136
rect 7156 16124 7162 16176
rect 11701 16167 11759 16173
rect 11701 16133 11713 16167
rect 11747 16164 11759 16167
rect 13998 16164 14004 16176
rect 11747 16136 12848 16164
rect 13959 16136 14004 16164
rect 11747 16133 11759 16136
rect 11701 16127 11759 16133
rect 2498 16056 2504 16108
rect 2556 16096 2562 16108
rect 2961 16099 3019 16105
rect 2961 16096 2973 16099
rect 2556 16068 2973 16096
rect 2556 16056 2562 16068
rect 2961 16065 2973 16068
rect 3007 16065 3019 16099
rect 2961 16059 3019 16065
rect 3237 16099 3295 16105
rect 3237 16065 3249 16099
rect 3283 16096 3295 16099
rect 5258 16096 5264 16108
rect 3283 16068 5264 16096
rect 3283 16065 3295 16068
rect 3237 16059 3295 16065
rect 5258 16056 5264 16068
rect 5316 16056 5322 16108
rect 5534 16056 5540 16108
rect 5592 16096 5598 16108
rect 5721 16099 5779 16105
rect 5721 16096 5733 16099
rect 5592 16068 5733 16096
rect 5592 16056 5598 16068
rect 5721 16065 5733 16068
rect 5767 16065 5779 16099
rect 5721 16059 5779 16065
rect 9122 16056 9128 16108
rect 9180 16096 9186 16108
rect 9677 16099 9735 16105
rect 9677 16096 9689 16099
rect 9180 16068 9689 16096
rect 9180 16056 9186 16068
rect 9677 16065 9689 16068
rect 9723 16065 9735 16099
rect 9677 16059 9735 16065
rect 12820 16040 12848 16136
rect 13998 16124 14004 16136
rect 14056 16124 14062 16176
rect 16114 16164 16120 16176
rect 14936 16136 16120 16164
rect 13280 16068 14596 16096
rect 5350 16028 5356 16040
rect 5311 16000 5356 16028
rect 5350 15988 5356 16000
rect 5408 15988 5414 16040
rect 5629 16031 5687 16037
rect 5629 15997 5641 16031
rect 5675 16028 5687 16031
rect 6178 16028 6184 16040
rect 5675 16000 6184 16028
rect 5675 15997 5687 16000
rect 5629 15991 5687 15997
rect 6178 15988 6184 16000
rect 6236 15988 6242 16040
rect 6825 16031 6883 16037
rect 6825 15997 6837 16031
rect 6871 15997 6883 16031
rect 7374 16028 7380 16040
rect 7335 16000 7380 16028
rect 6825 15991 6883 15997
rect 5994 15920 6000 15972
rect 6052 15960 6058 15972
rect 6840 15960 6868 15991
rect 7374 15988 7380 16000
rect 7432 15988 7438 16040
rect 7558 16028 7564 16040
rect 7519 16000 7564 16028
rect 7558 15988 7564 16000
rect 7616 15988 7622 16040
rect 8202 16028 8208 16040
rect 8163 16000 8208 16028
rect 8202 15988 8208 16000
rect 8260 15988 8266 16040
rect 8757 16031 8815 16037
rect 8757 15997 8769 16031
rect 8803 16028 8815 16031
rect 9030 16028 9036 16040
rect 8803 16000 9036 16028
rect 8803 15997 8815 16000
rect 8757 15991 8815 15997
rect 9030 15988 9036 16000
rect 9088 15988 9094 16040
rect 9398 16028 9404 16040
rect 9359 16000 9404 16028
rect 9398 15988 9404 16000
rect 9456 15988 9462 16040
rect 11514 16028 11520 16040
rect 11475 16000 11520 16028
rect 11514 15988 11520 16000
rect 11572 15988 11578 16040
rect 12802 16028 12808 16040
rect 12763 16000 12808 16028
rect 12802 15988 12808 16000
rect 12860 15988 12866 16040
rect 13280 16037 13308 16068
rect 14568 16040 14596 16068
rect 13265 16031 13323 16037
rect 13265 15997 13277 16031
rect 13311 15997 13323 16031
rect 13446 16028 13452 16040
rect 13407 16000 13452 16028
rect 13265 15991 13323 15997
rect 13446 15988 13452 16000
rect 13504 15988 13510 16040
rect 14093 16031 14151 16037
rect 14093 15997 14105 16031
rect 14139 16028 14151 16031
rect 14274 16028 14280 16040
rect 14139 16000 14280 16028
rect 14139 15997 14151 16000
rect 14093 15991 14151 15997
rect 14274 15988 14280 16000
rect 14332 15988 14338 16040
rect 14550 16028 14556 16040
rect 14511 16000 14556 16028
rect 14550 15988 14556 16000
rect 14608 15988 14614 16040
rect 14936 16037 14964 16136
rect 16114 16124 16120 16136
rect 16172 16124 16178 16176
rect 18046 16124 18052 16176
rect 18104 16164 18110 16176
rect 18141 16167 18199 16173
rect 18141 16164 18153 16167
rect 18104 16136 18153 16164
rect 18104 16124 18110 16136
rect 18141 16133 18153 16136
rect 18187 16133 18199 16167
rect 21358 16164 21364 16176
rect 18141 16127 18199 16133
rect 19812 16136 21364 16164
rect 19812 16096 19840 16136
rect 21358 16124 21364 16136
rect 21416 16164 21422 16176
rect 21910 16164 21916 16176
rect 21416 16136 21916 16164
rect 21416 16124 21422 16136
rect 21910 16124 21916 16136
rect 21968 16124 21974 16176
rect 19978 16096 19984 16108
rect 15304 16068 19840 16096
rect 19939 16068 19984 16096
rect 15304 16037 15332 16068
rect 19978 16056 19984 16068
rect 20036 16056 20042 16108
rect 22370 16096 22376 16108
rect 20732 16068 22376 16096
rect 20732 16040 20760 16068
rect 22370 16056 22376 16068
rect 22428 16056 22434 16108
rect 22664 16096 22692 16204
rect 34606 16192 34612 16244
rect 34664 16232 34670 16244
rect 34977 16235 35035 16241
rect 34977 16232 34989 16235
rect 34664 16204 34989 16232
rect 34664 16192 34670 16204
rect 34977 16201 34989 16204
rect 35023 16201 35035 16235
rect 34977 16195 35035 16201
rect 38841 16235 38899 16241
rect 38841 16201 38853 16235
rect 38887 16232 38899 16235
rect 38930 16232 38936 16244
rect 38887 16204 38936 16232
rect 38887 16201 38899 16204
rect 38841 16195 38899 16201
rect 38930 16192 38936 16204
rect 38988 16192 38994 16244
rect 28902 16164 28908 16176
rect 26344 16136 28908 16164
rect 23109 16099 23167 16105
rect 22664 16068 23060 16096
rect 14921 16031 14979 16037
rect 14921 15997 14933 16031
rect 14967 15997 14979 16031
rect 14921 15991 14979 15997
rect 15289 16031 15347 16037
rect 15289 15997 15301 16031
rect 15335 15997 15347 16031
rect 15289 15991 15347 15997
rect 15841 16031 15899 16037
rect 15841 15997 15853 16031
rect 15887 16028 15899 16031
rect 15930 16028 15936 16040
rect 15887 16000 15936 16028
rect 15887 15997 15899 16000
rect 15841 15991 15899 15997
rect 15930 15988 15936 16000
rect 15988 15988 15994 16040
rect 16669 16031 16727 16037
rect 16669 15997 16681 16031
rect 16715 15997 16727 16031
rect 16669 15991 16727 15997
rect 6052 15932 6868 15960
rect 11532 15960 11560 15988
rect 16684 15960 16712 15991
rect 17954 15988 17960 16040
rect 18012 16028 18018 16040
rect 18049 16031 18107 16037
rect 18049 16028 18061 16031
rect 18012 16000 18061 16028
rect 18012 15988 18018 16000
rect 18049 15997 18061 16000
rect 18095 15997 18107 16031
rect 18049 15991 18107 15997
rect 18414 15988 18420 16040
rect 18472 16028 18478 16040
rect 18693 16031 18751 16037
rect 18693 16028 18705 16031
rect 18472 16000 18705 16028
rect 18472 15988 18478 16000
rect 18693 15997 18705 16000
rect 18739 15997 18751 16031
rect 18693 15991 18751 15997
rect 19334 15988 19340 16040
rect 19392 16028 19398 16040
rect 19613 16031 19671 16037
rect 19613 16028 19625 16031
rect 19392 16000 19625 16028
rect 19392 15988 19398 16000
rect 19613 15997 19625 16000
rect 19659 15997 19671 16031
rect 19613 15991 19671 15997
rect 20073 16031 20131 16037
rect 20073 15997 20085 16031
rect 20119 15997 20131 16031
rect 20254 16028 20260 16040
rect 20215 16000 20260 16028
rect 20073 15991 20131 15997
rect 19426 15960 19432 15972
rect 11532 15932 16712 15960
rect 16776 15932 19432 15960
rect 6052 15920 6058 15932
rect 6840 15892 6868 15932
rect 11422 15892 11428 15904
rect 6840 15864 11428 15892
rect 11422 15852 11428 15864
rect 11480 15852 11486 15904
rect 13170 15852 13176 15904
rect 13228 15892 13234 15904
rect 16776 15892 16804 15932
rect 19426 15920 19432 15932
rect 19484 15920 19490 15972
rect 18782 15892 18788 15904
rect 13228 15864 16804 15892
rect 18743 15864 18788 15892
rect 13228 15852 13234 15864
rect 18782 15852 18788 15864
rect 18840 15852 18846 15904
rect 19628 15892 19656 15991
rect 20088 15960 20116 15991
rect 20254 15988 20260 16000
rect 20312 15988 20318 16040
rect 20714 16028 20720 16040
rect 20675 16000 20720 16028
rect 20714 15988 20720 16000
rect 20772 15988 20778 16040
rect 20990 15988 20996 16040
rect 21048 16028 21054 16040
rect 21085 16031 21143 16037
rect 21085 16028 21097 16031
rect 21048 16000 21097 16028
rect 21048 15988 21054 16000
rect 21085 15997 21097 16000
rect 21131 15997 21143 16031
rect 21085 15991 21143 15997
rect 21174 15988 21180 16040
rect 21232 16028 21238 16040
rect 22462 16028 22468 16040
rect 21232 16000 22468 16028
rect 21232 15988 21238 16000
rect 22462 15988 22468 16000
rect 22520 15988 22526 16040
rect 22664 16037 22692 16068
rect 22649 16031 22707 16037
rect 22649 15997 22661 16031
rect 22695 15997 22707 16031
rect 22649 15991 22707 15997
rect 22833 16031 22891 16037
rect 22833 15997 22845 16031
rect 22879 15997 22891 16031
rect 23032 16028 23060 16068
rect 23109 16065 23121 16099
rect 23155 16096 23167 16099
rect 23474 16096 23480 16108
rect 23155 16068 23480 16096
rect 23155 16065 23167 16068
rect 23109 16059 23167 16065
rect 23474 16056 23480 16068
rect 23532 16056 23538 16108
rect 24302 16096 24308 16108
rect 24263 16068 24308 16096
rect 24302 16056 24308 16068
rect 24360 16056 24366 16108
rect 26344 16105 26372 16136
rect 28902 16124 28908 16136
rect 28960 16124 28966 16176
rect 26329 16099 26387 16105
rect 26329 16065 26341 16099
rect 26375 16065 26387 16099
rect 26329 16059 26387 16065
rect 26878 16056 26884 16108
rect 26936 16096 26942 16108
rect 27801 16099 27859 16105
rect 27801 16096 27813 16099
rect 26936 16068 27813 16096
rect 26936 16056 26942 16068
rect 27801 16065 27813 16068
rect 27847 16065 27859 16099
rect 27801 16059 27859 16065
rect 30466 16056 30472 16108
rect 30524 16096 30530 16108
rect 30561 16099 30619 16105
rect 30561 16096 30573 16099
rect 30524 16068 30573 16096
rect 30524 16056 30530 16068
rect 30561 16065 30573 16068
rect 30607 16065 30619 16099
rect 32306 16096 32312 16108
rect 30561 16059 30619 16065
rect 32048 16068 32312 16096
rect 23658 16028 23664 16040
rect 23032 16000 23664 16028
rect 22833 15991 22891 15997
rect 21818 15960 21824 15972
rect 20088 15932 21824 15960
rect 21818 15920 21824 15932
rect 21876 15960 21882 15972
rect 22848 15960 22876 15991
rect 23658 15988 23664 16000
rect 23716 15988 23722 16040
rect 24210 16028 24216 16040
rect 24171 16000 24216 16028
rect 24210 15988 24216 16000
rect 24268 15988 24274 16040
rect 26605 16031 26663 16037
rect 26605 15997 26617 16031
rect 26651 15997 26663 16031
rect 26605 15991 26663 15997
rect 26789 16031 26847 16037
rect 26789 15997 26801 16031
rect 26835 16028 26847 16031
rect 27614 16028 27620 16040
rect 26835 16000 27620 16028
rect 26835 15997 26847 16000
rect 26789 15991 26847 15997
rect 21876 15932 22876 15960
rect 25777 15963 25835 15969
rect 21876 15920 21882 15932
rect 25777 15929 25789 15963
rect 25823 15960 25835 15963
rect 26510 15960 26516 15972
rect 25823 15932 26516 15960
rect 25823 15929 25835 15932
rect 25777 15923 25835 15929
rect 26510 15920 26516 15932
rect 26568 15920 26574 15972
rect 26620 15960 26648 15991
rect 27614 15988 27620 16000
rect 27672 15988 27678 16040
rect 28074 16028 28080 16040
rect 28035 16000 28080 16028
rect 28074 15988 28080 16000
rect 28132 15988 28138 16040
rect 28258 16028 28264 16040
rect 28219 16000 28264 16028
rect 28258 15988 28264 16000
rect 28316 15988 28322 16040
rect 30098 15988 30104 16040
rect 30156 16028 30162 16040
rect 30285 16031 30343 16037
rect 30285 16028 30297 16031
rect 30156 16000 30297 16028
rect 30156 15988 30162 16000
rect 30285 15997 30297 16000
rect 30331 16028 30343 16031
rect 32048 16028 32076 16068
rect 32306 16056 32312 16068
rect 32364 16056 32370 16108
rect 34790 16096 34796 16108
rect 33336 16068 34796 16096
rect 32398 16028 32404 16040
rect 30331 16000 32076 16028
rect 32359 16000 32404 16028
rect 30331 15997 30343 16000
rect 30285 15991 30343 15997
rect 32398 15988 32404 16000
rect 32456 15988 32462 16040
rect 33336 16037 33364 16068
rect 34790 16056 34796 16068
rect 34848 16056 34854 16108
rect 35894 16056 35900 16108
rect 35952 16096 35958 16108
rect 37550 16096 37556 16108
rect 35952 16068 36584 16096
rect 37511 16068 37556 16096
rect 35952 16056 35958 16068
rect 33321 16031 33379 16037
rect 33321 15997 33333 16031
rect 33367 15997 33379 16031
rect 33502 16028 33508 16040
rect 33463 16000 33508 16028
rect 33321 15991 33379 15997
rect 33502 15988 33508 16000
rect 33560 15988 33566 16040
rect 34149 16031 34207 16037
rect 34149 15997 34161 16031
rect 34195 15997 34207 16031
rect 34149 15991 34207 15997
rect 34333 16031 34391 16037
rect 34333 15997 34345 16031
rect 34379 16028 34391 16031
rect 34885 16031 34943 16037
rect 34885 16028 34897 16031
rect 34379 16000 34897 16028
rect 34379 15997 34391 16000
rect 34333 15991 34391 15997
rect 34885 15997 34897 16000
rect 34931 15997 34943 16031
rect 34885 15991 34943 15997
rect 35621 16031 35679 16037
rect 35621 15997 35633 16031
rect 35667 16028 35679 16031
rect 35802 16028 35808 16040
rect 35667 16000 35808 16028
rect 35667 15997 35679 16000
rect 35621 15991 35679 15997
rect 27249 15963 27307 15969
rect 27249 15960 27261 15963
rect 26620 15932 27261 15960
rect 27249 15929 27261 15932
rect 27295 15929 27307 15963
rect 34164 15960 34192 15991
rect 35802 15988 35808 16000
rect 35860 15988 35866 16040
rect 35986 16028 35992 16040
rect 35947 16000 35992 16028
rect 35986 15988 35992 16000
rect 36044 15988 36050 16040
rect 36556 16037 36584 16068
rect 37550 16056 37556 16068
rect 37608 16056 37614 16108
rect 36173 16031 36231 16037
rect 36173 15997 36185 16031
rect 36219 15997 36231 16031
rect 36173 15991 36231 15997
rect 36541 16031 36599 16037
rect 36541 15997 36553 16031
rect 36587 15997 36599 16031
rect 36541 15991 36599 15997
rect 37277 16031 37335 16037
rect 37277 15997 37289 16031
rect 37323 16028 37335 16031
rect 37366 16028 37372 16040
rect 37323 16000 37372 16028
rect 37323 15997 37335 16000
rect 37277 15991 37335 15997
rect 34698 15960 34704 15972
rect 34164 15932 34704 15960
rect 27249 15923 27307 15929
rect 34698 15920 34704 15932
rect 34756 15920 34762 15972
rect 20530 15892 20536 15904
rect 19628 15864 20536 15892
rect 20530 15852 20536 15864
rect 20588 15852 20594 15904
rect 20990 15852 20996 15904
rect 21048 15892 21054 15904
rect 21266 15892 21272 15904
rect 21048 15864 21272 15892
rect 21048 15852 21054 15864
rect 21266 15852 21272 15864
rect 21324 15852 21330 15904
rect 21634 15852 21640 15904
rect 21692 15892 21698 15904
rect 22922 15892 22928 15904
rect 21692 15864 22928 15892
rect 21692 15852 21698 15864
rect 22922 15852 22928 15864
rect 22980 15852 22986 15904
rect 23382 15852 23388 15904
rect 23440 15892 23446 15904
rect 30098 15892 30104 15904
rect 23440 15864 30104 15892
rect 23440 15852 23446 15864
rect 30098 15852 30104 15864
rect 30156 15852 30162 15904
rect 31662 15892 31668 15904
rect 31623 15864 31668 15892
rect 31662 15852 31668 15864
rect 31720 15852 31726 15904
rect 32214 15852 32220 15904
rect 32272 15892 32278 15904
rect 32493 15895 32551 15901
rect 32493 15892 32505 15895
rect 32272 15864 32505 15892
rect 32272 15852 32278 15864
rect 32493 15861 32505 15864
rect 32539 15861 32551 15895
rect 32493 15855 32551 15861
rect 34330 15852 34336 15904
rect 34388 15892 34394 15904
rect 36188 15892 36216 15991
rect 37366 15988 37372 16000
rect 37424 15988 37430 16040
rect 34388 15864 36216 15892
rect 34388 15852 34394 15864
rect 1104 15802 39836 15824
rect 1104 15750 19606 15802
rect 19658 15750 19670 15802
rect 19722 15750 19734 15802
rect 19786 15750 19798 15802
rect 19850 15750 39836 15802
rect 1104 15728 39836 15750
rect 2424 15660 7144 15688
rect 1394 15552 1400 15564
rect 1355 15524 1400 15552
rect 1394 15512 1400 15524
rect 1452 15512 1458 15564
rect 1673 15555 1731 15561
rect 1673 15521 1685 15555
rect 1719 15552 1731 15555
rect 2424 15552 2452 15660
rect 7116 15620 7144 15660
rect 7190 15648 7196 15700
rect 7248 15688 7254 15700
rect 7561 15691 7619 15697
rect 7561 15688 7573 15691
rect 7248 15660 7573 15688
rect 7248 15648 7254 15660
rect 7561 15657 7573 15660
rect 7607 15657 7619 15691
rect 7561 15651 7619 15657
rect 13906 15648 13912 15700
rect 13964 15688 13970 15700
rect 14277 15691 14335 15697
rect 13964 15660 14228 15688
rect 13964 15648 13970 15660
rect 7926 15620 7932 15632
rect 7116 15592 7932 15620
rect 7926 15580 7932 15592
rect 7984 15580 7990 15632
rect 8202 15580 8208 15632
rect 8260 15620 8266 15632
rect 12618 15620 12624 15632
rect 8260 15592 12624 15620
rect 8260 15580 8266 15592
rect 1719 15524 2452 15552
rect 1719 15521 1731 15524
rect 1673 15515 1731 15521
rect 2498 15512 2504 15564
rect 2556 15552 2562 15564
rect 2682 15552 2688 15564
rect 2556 15524 2688 15552
rect 2556 15512 2562 15524
rect 2682 15512 2688 15524
rect 2740 15552 2746 15564
rect 8312 15561 8340 15592
rect 12618 15580 12624 15592
rect 12676 15580 12682 15632
rect 12802 15580 12808 15632
rect 12860 15620 12866 15632
rect 14200 15620 14228 15660
rect 14277 15657 14289 15691
rect 14323 15688 14335 15691
rect 14458 15688 14464 15700
rect 14323 15660 14464 15688
rect 14323 15657 14335 15660
rect 14277 15651 14335 15657
rect 14458 15648 14464 15660
rect 14516 15648 14522 15700
rect 14550 15648 14556 15700
rect 14608 15688 14614 15700
rect 16025 15691 16083 15697
rect 16025 15688 16037 15691
rect 14608 15660 16037 15688
rect 14608 15648 14614 15660
rect 16025 15657 16037 15660
rect 16071 15657 16083 15691
rect 16025 15651 16083 15657
rect 16114 15648 16120 15700
rect 16172 15688 16178 15700
rect 21174 15688 21180 15700
rect 16172 15660 21180 15688
rect 16172 15648 16178 15660
rect 21174 15648 21180 15660
rect 21232 15648 21238 15700
rect 28718 15648 28724 15700
rect 28776 15688 28782 15700
rect 28776 15660 30052 15688
rect 28776 15648 28782 15660
rect 18414 15620 18420 15632
rect 12860 15592 14044 15620
rect 14200 15592 15976 15620
rect 18375 15592 18420 15620
rect 12860 15580 12866 15592
rect 4065 15555 4123 15561
rect 4065 15552 4077 15555
rect 2740 15524 4077 15552
rect 2740 15512 2746 15524
rect 4065 15521 4077 15524
rect 4111 15521 4123 15555
rect 4065 15515 4123 15521
rect 5721 15555 5779 15561
rect 5721 15521 5733 15555
rect 5767 15552 5779 15555
rect 6457 15555 6515 15561
rect 6457 15552 6469 15555
rect 5767 15524 6469 15552
rect 5767 15521 5779 15524
rect 5721 15515 5779 15521
rect 6457 15521 6469 15524
rect 6503 15521 6515 15555
rect 6457 15515 6515 15521
rect 8297 15555 8355 15561
rect 8297 15521 8309 15555
rect 8343 15521 8355 15555
rect 8297 15515 8355 15521
rect 8386 15512 8392 15564
rect 8444 15552 8450 15564
rect 10137 15555 10195 15561
rect 10137 15552 10149 15555
rect 8444 15524 10149 15552
rect 8444 15512 8450 15524
rect 10137 15521 10149 15524
rect 10183 15521 10195 15555
rect 10870 15552 10876 15564
rect 10831 15524 10876 15552
rect 10137 15515 10195 15521
rect 10870 15512 10876 15524
rect 10928 15512 10934 15564
rect 11422 15552 11428 15564
rect 11383 15524 11428 15552
rect 11422 15512 11428 15524
rect 11480 15512 11486 15564
rect 11790 15552 11796 15564
rect 11751 15524 11796 15552
rect 11790 15512 11796 15524
rect 11848 15512 11854 15564
rect 11974 15552 11980 15564
rect 11887 15524 11980 15552
rect 11974 15512 11980 15524
rect 12032 15552 12038 15564
rect 12069 15555 12127 15561
rect 12069 15552 12081 15555
rect 12032 15524 12081 15552
rect 12032 15512 12038 15524
rect 12069 15521 12081 15524
rect 12115 15521 12127 15555
rect 12636 15552 12664 15580
rect 14016 15561 14044 15592
rect 12713 15555 12771 15561
rect 12713 15552 12725 15555
rect 12636 15524 12725 15552
rect 12069 15515 12127 15521
rect 12713 15521 12725 15524
rect 12759 15521 12771 15555
rect 12713 15515 12771 15521
rect 13265 15555 13323 15561
rect 13265 15521 13277 15555
rect 13311 15552 13323 15555
rect 13909 15555 13967 15561
rect 13311 15524 13860 15552
rect 13311 15521 13323 15524
rect 13265 15515 13323 15521
rect 4341 15487 4399 15493
rect 4341 15453 4353 15487
rect 4387 15484 4399 15487
rect 5166 15484 5172 15496
rect 4387 15456 5172 15484
rect 4387 15453 4399 15456
rect 4341 15447 4399 15453
rect 5166 15444 5172 15456
rect 5224 15444 5230 15496
rect 6181 15487 6239 15493
rect 6181 15453 6193 15487
rect 6227 15484 6239 15487
rect 6822 15484 6828 15496
rect 6227 15456 6828 15484
rect 6227 15453 6239 15456
rect 6181 15447 6239 15453
rect 6822 15444 6828 15456
rect 6880 15444 6886 15496
rect 7558 15444 7564 15496
rect 7616 15484 7622 15496
rect 10505 15487 10563 15493
rect 7616 15456 10456 15484
rect 7616 15444 7622 15456
rect 2777 15351 2835 15357
rect 2777 15317 2789 15351
rect 2823 15348 2835 15351
rect 2866 15348 2872 15360
rect 2823 15320 2872 15348
rect 2823 15317 2835 15320
rect 2777 15311 2835 15317
rect 2866 15308 2872 15320
rect 2924 15308 2930 15360
rect 8202 15308 8208 15360
rect 8260 15348 8266 15360
rect 8481 15351 8539 15357
rect 8481 15348 8493 15351
rect 8260 15320 8493 15348
rect 8260 15308 8266 15320
rect 8481 15317 8493 15320
rect 8527 15317 8539 15351
rect 10428 15348 10456 15456
rect 10505 15453 10517 15487
rect 10551 15484 10563 15487
rect 11882 15484 11888 15496
rect 10551 15456 11888 15484
rect 10551 15453 10563 15456
rect 10505 15447 10563 15453
rect 11882 15444 11888 15456
rect 11940 15444 11946 15496
rect 11606 15416 11612 15428
rect 11567 15388 11612 15416
rect 11606 15376 11612 15388
rect 11664 15376 11670 15428
rect 11992 15348 12020 15512
rect 10428 15320 12020 15348
rect 8481 15311 8539 15317
rect 13630 15308 13636 15360
rect 13688 15348 13694 15360
rect 13725 15351 13783 15357
rect 13725 15348 13737 15351
rect 13688 15320 13737 15348
rect 13688 15308 13694 15320
rect 13725 15317 13737 15320
rect 13771 15317 13783 15351
rect 13832 15348 13860 15524
rect 13909 15521 13921 15555
rect 13955 15521 13967 15555
rect 13909 15515 13967 15521
rect 14001 15555 14059 15561
rect 14001 15521 14013 15555
rect 14047 15521 14059 15555
rect 14001 15515 14059 15521
rect 14553 15555 14611 15561
rect 14553 15521 14565 15555
rect 14599 15552 14611 15555
rect 14642 15552 14648 15564
rect 14599 15524 14648 15552
rect 14599 15521 14611 15524
rect 14553 15515 14611 15521
rect 13924 15416 13952 15515
rect 14642 15512 14648 15524
rect 14700 15512 14706 15564
rect 15948 15561 15976 15592
rect 18414 15580 18420 15592
rect 18472 15580 18478 15632
rect 18782 15580 18788 15632
rect 18840 15620 18846 15632
rect 27065 15623 27123 15629
rect 18840 15592 19840 15620
rect 18840 15580 18846 15592
rect 15289 15555 15347 15561
rect 15289 15521 15301 15555
rect 15335 15552 15347 15555
rect 15933 15555 15991 15561
rect 15335 15524 15884 15552
rect 15335 15521 15347 15524
rect 15289 15515 15347 15521
rect 14660 15484 14688 15512
rect 15381 15487 15439 15493
rect 15381 15484 15393 15487
rect 14660 15456 15393 15484
rect 15381 15453 15393 15456
rect 15427 15453 15439 15487
rect 15856 15484 15884 15524
rect 15933 15521 15945 15555
rect 15979 15521 15991 15555
rect 16758 15552 16764 15564
rect 16719 15524 16764 15552
rect 15933 15515 15991 15521
rect 16758 15512 16764 15524
rect 16816 15512 16822 15564
rect 18966 15552 18972 15564
rect 16868 15524 18972 15552
rect 16298 15484 16304 15496
rect 15856 15456 16304 15484
rect 15381 15447 15439 15453
rect 16298 15444 16304 15456
rect 16356 15444 16362 15496
rect 16868 15484 16896 15524
rect 18966 15512 18972 15524
rect 19024 15552 19030 15564
rect 19061 15555 19119 15561
rect 19061 15552 19073 15555
rect 19024 15524 19073 15552
rect 19024 15512 19030 15524
rect 19061 15521 19073 15524
rect 19107 15521 19119 15555
rect 19061 15515 19119 15521
rect 19150 15512 19156 15564
rect 19208 15552 19214 15564
rect 19812 15561 19840 15592
rect 27065 15589 27077 15623
rect 27111 15620 27123 15623
rect 27111 15592 29868 15620
rect 27111 15589 27123 15592
rect 27065 15583 27123 15589
rect 19613 15555 19671 15561
rect 19613 15552 19625 15555
rect 19208 15524 19625 15552
rect 19208 15512 19214 15524
rect 19613 15521 19625 15524
rect 19659 15521 19671 15555
rect 19613 15515 19671 15521
rect 19797 15555 19855 15561
rect 19797 15521 19809 15555
rect 19843 15521 19855 15555
rect 19797 15515 19855 15521
rect 20530 15512 20536 15564
rect 20588 15552 20594 15564
rect 21269 15555 21327 15561
rect 21269 15552 21281 15555
rect 20588 15524 21281 15552
rect 20588 15512 20594 15524
rect 21269 15521 21281 15524
rect 21315 15521 21327 15555
rect 21269 15515 21327 15521
rect 21913 15555 21971 15561
rect 21913 15521 21925 15555
rect 21959 15552 21971 15555
rect 22094 15552 22100 15564
rect 21959 15524 22100 15552
rect 21959 15521 21971 15524
rect 21913 15515 21971 15521
rect 22094 15512 22100 15524
rect 22152 15512 22158 15564
rect 22281 15555 22339 15561
rect 22281 15521 22293 15555
rect 22327 15552 22339 15555
rect 22370 15552 22376 15564
rect 22327 15524 22376 15552
rect 22327 15521 22339 15524
rect 22281 15515 22339 15521
rect 22370 15512 22376 15524
rect 22428 15512 22434 15564
rect 22462 15512 22468 15564
rect 22520 15552 22526 15564
rect 22520 15524 22565 15552
rect 22520 15512 22526 15524
rect 22646 15512 22652 15564
rect 22704 15552 22710 15564
rect 22925 15555 22983 15561
rect 22925 15552 22937 15555
rect 22704 15524 22937 15552
rect 22704 15512 22710 15524
rect 22925 15521 22937 15524
rect 22971 15521 22983 15555
rect 23658 15552 23664 15564
rect 23619 15524 23664 15552
rect 22925 15515 22983 15521
rect 23658 15512 23664 15524
rect 23716 15512 23722 15564
rect 24121 15555 24179 15561
rect 24121 15521 24133 15555
rect 24167 15521 24179 15555
rect 26602 15552 26608 15564
rect 26563 15524 26608 15552
rect 24121 15515 24179 15521
rect 16776 15456 16896 15484
rect 17037 15487 17095 15493
rect 15102 15416 15108 15428
rect 13924 15388 15108 15416
rect 15102 15376 15108 15388
rect 15160 15376 15166 15428
rect 15470 15376 15476 15428
rect 15528 15416 15534 15428
rect 16776 15416 16804 15456
rect 17037 15453 17049 15487
rect 17083 15484 17095 15487
rect 18874 15484 18880 15496
rect 17083 15456 18552 15484
rect 18835 15456 18880 15484
rect 17083 15453 17095 15456
rect 17037 15447 17095 15453
rect 15528 15388 16804 15416
rect 18524 15416 18552 15456
rect 18874 15444 18880 15456
rect 18932 15444 18938 15496
rect 22186 15484 22192 15496
rect 22147 15456 22192 15484
rect 22186 15444 22192 15456
rect 22244 15444 22250 15496
rect 23014 15444 23020 15496
rect 23072 15484 23078 15496
rect 24136 15484 24164 15515
rect 26602 15512 26608 15524
rect 26660 15512 26666 15564
rect 28445 15555 28503 15561
rect 28445 15521 28457 15555
rect 28491 15552 28503 15555
rect 28718 15552 28724 15564
rect 28491 15524 28724 15552
rect 28491 15521 28503 15524
rect 28445 15515 28503 15521
rect 28718 15512 28724 15524
rect 28776 15512 28782 15564
rect 28813 15555 28871 15561
rect 28813 15521 28825 15555
rect 28859 15552 28871 15555
rect 29178 15552 29184 15564
rect 28859 15524 29184 15552
rect 28859 15521 28871 15524
rect 28813 15515 28871 15521
rect 29178 15512 29184 15524
rect 29236 15512 29242 15564
rect 24394 15484 24400 15496
rect 23072 15456 24164 15484
rect 24355 15456 24400 15484
rect 23072 15444 23078 15456
rect 24394 15444 24400 15456
rect 24452 15444 24458 15496
rect 26142 15444 26148 15496
rect 26200 15484 26206 15496
rect 26513 15487 26571 15493
rect 26513 15484 26525 15487
rect 26200 15456 26525 15484
rect 26200 15444 26206 15456
rect 26513 15453 26525 15456
rect 26559 15453 26571 15487
rect 26513 15447 26571 15453
rect 28077 15487 28135 15493
rect 28077 15453 28089 15487
rect 28123 15484 28135 15487
rect 28994 15484 29000 15496
rect 28123 15456 29000 15484
rect 28123 15453 28135 15456
rect 28077 15447 28135 15453
rect 28994 15444 29000 15456
rect 29052 15444 29058 15496
rect 29733 15487 29791 15493
rect 29733 15453 29745 15487
rect 29779 15453 29791 15487
rect 29840 15484 29868 15592
rect 30024 15561 30052 15660
rect 30098 15648 30104 15700
rect 30156 15688 30162 15700
rect 33502 15688 33508 15700
rect 30156 15660 33508 15688
rect 30156 15648 30162 15660
rect 33502 15648 33508 15660
rect 33560 15648 33566 15700
rect 33594 15648 33600 15700
rect 33652 15688 33658 15700
rect 33965 15691 34023 15697
rect 33965 15688 33977 15691
rect 33652 15660 33977 15688
rect 33652 15648 33658 15660
rect 33965 15657 33977 15660
rect 34011 15688 34023 15691
rect 34422 15688 34428 15700
rect 34011 15660 34428 15688
rect 34011 15657 34023 15660
rect 33965 15651 34023 15657
rect 34422 15648 34428 15660
rect 34480 15648 34486 15700
rect 35894 15688 35900 15700
rect 34716 15660 35900 15688
rect 30009 15555 30067 15561
rect 30009 15521 30021 15555
rect 30055 15521 30067 15555
rect 30009 15515 30067 15521
rect 30098 15512 30104 15564
rect 30156 15552 30162 15564
rect 30469 15555 30527 15561
rect 30469 15552 30481 15555
rect 30156 15524 30481 15552
rect 30156 15512 30162 15524
rect 30469 15521 30481 15524
rect 30515 15521 30527 15555
rect 30469 15515 30527 15521
rect 31205 15555 31263 15561
rect 31205 15521 31217 15555
rect 31251 15552 31263 15555
rect 31303 15555 31361 15561
rect 31303 15552 31315 15555
rect 31251 15524 31315 15552
rect 31251 15521 31263 15524
rect 31205 15515 31263 15521
rect 31303 15521 31315 15524
rect 31349 15521 31361 15555
rect 31303 15515 31361 15521
rect 31846 15512 31852 15564
rect 31904 15552 31910 15564
rect 32030 15552 32036 15564
rect 31904 15524 32036 15552
rect 31904 15512 31910 15524
rect 32030 15512 32036 15524
rect 32088 15552 32094 15564
rect 32125 15555 32183 15561
rect 32125 15552 32137 15555
rect 32088 15524 32137 15552
rect 32088 15512 32094 15524
rect 32125 15521 32137 15524
rect 32171 15521 32183 15555
rect 32766 15552 32772 15564
rect 32727 15524 32772 15552
rect 32125 15515 32183 15521
rect 32766 15512 32772 15524
rect 32824 15512 32830 15564
rect 33873 15555 33931 15561
rect 33873 15521 33885 15555
rect 33919 15552 33931 15555
rect 34330 15552 34336 15564
rect 33919 15524 34336 15552
rect 33919 15521 33931 15524
rect 33873 15515 33931 15521
rect 34330 15512 34336 15524
rect 34388 15512 34394 15564
rect 34514 15552 34520 15564
rect 34475 15524 34520 15552
rect 34514 15512 34520 15524
rect 34572 15512 34578 15564
rect 34716 15561 34744 15660
rect 35894 15648 35900 15660
rect 35952 15648 35958 15700
rect 36630 15648 36636 15700
rect 36688 15688 36694 15700
rect 36909 15691 36967 15697
rect 36909 15688 36921 15691
rect 36688 15660 36921 15688
rect 36688 15648 36694 15660
rect 36909 15657 36921 15660
rect 36955 15657 36967 15691
rect 36909 15651 36967 15657
rect 34701 15555 34759 15561
rect 34701 15521 34713 15555
rect 34747 15521 34759 15555
rect 34701 15515 34759 15521
rect 35069 15555 35127 15561
rect 35069 15521 35081 15555
rect 35115 15552 35127 15555
rect 35805 15555 35863 15561
rect 35805 15552 35817 15555
rect 35115 15524 35817 15552
rect 35115 15521 35127 15524
rect 35069 15515 35127 15521
rect 35805 15521 35817 15524
rect 35851 15521 35863 15555
rect 37918 15552 37924 15564
rect 37879 15524 37924 15552
rect 35805 15515 35863 15521
rect 37918 15512 37924 15524
rect 37976 15512 37982 15564
rect 38470 15552 38476 15564
rect 38431 15524 38476 15552
rect 38470 15512 38476 15524
rect 38528 15512 38534 15564
rect 31938 15484 31944 15496
rect 29840 15456 31944 15484
rect 29733 15447 29791 15453
rect 19981 15419 20039 15425
rect 19981 15416 19993 15419
rect 18524 15388 19993 15416
rect 15528 15376 15534 15388
rect 19981 15385 19993 15388
rect 20027 15385 20039 15419
rect 19981 15379 20039 15385
rect 28534 15376 28540 15428
rect 28592 15416 28598 15428
rect 28721 15419 28779 15425
rect 28721 15416 28733 15419
rect 28592 15388 28733 15416
rect 28592 15376 28598 15388
rect 28721 15385 28733 15388
rect 28767 15385 28779 15419
rect 28721 15379 28779 15385
rect 22278 15348 22284 15360
rect 13832 15320 22284 15348
rect 13725 15311 13783 15317
rect 22278 15308 22284 15320
rect 22336 15348 22342 15360
rect 27154 15348 27160 15360
rect 22336 15320 27160 15348
rect 22336 15308 22342 15320
rect 27154 15308 27160 15320
rect 27212 15308 27218 15360
rect 29748 15348 29776 15447
rect 31938 15444 31944 15456
rect 31996 15444 32002 15496
rect 32306 15444 32312 15496
rect 32364 15484 32370 15496
rect 32953 15487 33011 15493
rect 32953 15484 32965 15487
rect 32364 15456 32965 15484
rect 32364 15444 32370 15456
rect 32953 15453 32965 15456
rect 32999 15453 33011 15487
rect 32953 15447 33011 15453
rect 35529 15487 35587 15493
rect 35529 15453 35541 15487
rect 35575 15484 35587 15487
rect 37366 15484 37372 15496
rect 35575 15456 37372 15484
rect 35575 15453 35587 15456
rect 35529 15447 35587 15453
rect 37366 15444 37372 15456
rect 37424 15444 37430 15496
rect 38378 15484 38384 15496
rect 38339 15456 38384 15484
rect 38378 15444 38384 15456
rect 38436 15444 38442 15496
rect 30374 15376 30380 15428
rect 30432 15416 30438 15428
rect 30469 15419 30527 15425
rect 30469 15416 30481 15419
rect 30432 15388 30481 15416
rect 30432 15376 30438 15388
rect 30469 15385 30481 15388
rect 30515 15385 30527 15419
rect 30469 15379 30527 15385
rect 31205 15419 31263 15425
rect 31205 15385 31217 15419
rect 31251 15416 31263 15419
rect 32214 15416 32220 15428
rect 31251 15388 32220 15416
rect 31251 15385 31263 15388
rect 31205 15379 31263 15385
rect 32214 15376 32220 15388
rect 32272 15376 32278 15428
rect 32401 15419 32459 15425
rect 32401 15385 32413 15419
rect 32447 15416 32459 15419
rect 33318 15416 33324 15428
rect 32447 15388 33324 15416
rect 32447 15385 32459 15388
rect 32401 15379 32459 15385
rect 33318 15376 33324 15388
rect 33376 15376 33382 15428
rect 31386 15348 31392 15360
rect 29748 15320 31392 15348
rect 31386 15308 31392 15320
rect 31444 15308 31450 15360
rect 31478 15308 31484 15360
rect 31536 15348 31542 15360
rect 31536 15320 31581 15348
rect 31536 15308 31542 15320
rect 37918 15308 37924 15360
rect 37976 15348 37982 15360
rect 38657 15351 38715 15357
rect 38657 15348 38669 15351
rect 37976 15320 38669 15348
rect 37976 15308 37982 15320
rect 38657 15317 38669 15320
rect 38703 15317 38715 15351
rect 38657 15311 38715 15317
rect 1104 15258 39836 15280
rect 1104 15206 4246 15258
rect 4298 15206 4310 15258
rect 4362 15206 4374 15258
rect 4426 15206 4438 15258
rect 4490 15206 34966 15258
rect 35018 15206 35030 15258
rect 35082 15206 35094 15258
rect 35146 15206 35158 15258
rect 35210 15206 39836 15258
rect 1104 15184 39836 15206
rect 4062 15104 4068 15156
rect 4120 15144 4126 15156
rect 5166 15144 5172 15156
rect 4120 15116 4752 15144
rect 5127 15116 5172 15144
rect 4120 15104 4126 15116
rect 4724 15076 4752 15116
rect 5166 15104 5172 15116
rect 5224 15104 5230 15156
rect 8386 15144 8392 15156
rect 5276 15116 7788 15144
rect 8347 15116 8392 15144
rect 5276 15076 5304 15116
rect 4724 15048 5304 15076
rect 7760 15076 7788 15116
rect 8386 15104 8392 15116
rect 8444 15104 8450 15156
rect 9214 15104 9220 15156
rect 9272 15144 9278 15156
rect 9398 15144 9404 15156
rect 9272 15116 9404 15144
rect 9272 15104 9278 15116
rect 9398 15104 9404 15116
rect 9456 15144 9462 15156
rect 11422 15144 11428 15156
rect 9456 15116 11428 15144
rect 9456 15104 9462 15116
rect 11422 15104 11428 15116
rect 11480 15144 11486 15156
rect 11885 15147 11943 15153
rect 11885 15144 11897 15147
rect 11480 15116 11897 15144
rect 11480 15104 11486 15116
rect 11885 15113 11897 15116
rect 11931 15144 11943 15147
rect 12434 15144 12440 15156
rect 11931 15116 12440 15144
rect 11931 15113 11943 15116
rect 11885 15107 11943 15113
rect 12434 15104 12440 15116
rect 12492 15104 12498 15156
rect 12894 15104 12900 15156
rect 12952 15144 12958 15156
rect 17494 15144 17500 15156
rect 12952 15116 17500 15144
rect 12952 15104 12958 15116
rect 17494 15104 17500 15116
rect 17552 15104 17558 15156
rect 19426 15104 19432 15156
rect 19484 15144 19490 15156
rect 19886 15144 19892 15156
rect 19484 15116 19892 15144
rect 19484 15104 19490 15116
rect 19886 15104 19892 15116
rect 19944 15104 19950 15156
rect 20162 15104 20168 15156
rect 20220 15144 20226 15156
rect 20530 15144 20536 15156
rect 20220 15116 20536 15144
rect 20220 15104 20226 15116
rect 20530 15104 20536 15116
rect 20588 15104 20594 15156
rect 21818 15144 21824 15156
rect 21779 15116 21824 15144
rect 21818 15104 21824 15116
rect 21876 15104 21882 15156
rect 28994 15104 29000 15156
rect 29052 15144 29058 15156
rect 30282 15144 30288 15156
rect 29052 15116 30288 15144
rect 29052 15104 29058 15116
rect 30282 15104 30288 15116
rect 30340 15104 30346 15156
rect 31386 15104 31392 15156
rect 31444 15144 31450 15156
rect 31481 15147 31539 15153
rect 31481 15144 31493 15147
rect 31444 15116 31493 15144
rect 31444 15104 31450 15116
rect 31481 15113 31493 15116
rect 31527 15113 31539 15147
rect 31481 15107 31539 15113
rect 33226 15104 33232 15156
rect 33284 15144 33290 15156
rect 34057 15147 34115 15153
rect 34057 15144 34069 15147
rect 33284 15116 34069 15144
rect 33284 15104 33290 15116
rect 34057 15113 34069 15116
rect 34103 15113 34115 15147
rect 34057 15107 34115 15113
rect 38102 15104 38108 15156
rect 38160 15144 38166 15156
rect 38841 15147 38899 15153
rect 38841 15144 38853 15147
rect 38160 15116 38853 15144
rect 38160 15104 38166 15116
rect 38841 15113 38853 15116
rect 38887 15113 38899 15147
rect 38841 15107 38899 15113
rect 12158 15076 12164 15088
rect 7760 15048 12164 15076
rect 12158 15036 12164 15048
rect 12216 15036 12222 15088
rect 13814 15076 13820 15088
rect 13372 15048 13820 15076
rect 3329 15011 3387 15017
rect 3329 14977 3341 15011
rect 3375 15008 3387 15011
rect 4065 15011 4123 15017
rect 4065 15008 4077 15011
rect 3375 14980 4077 15008
rect 3375 14977 3387 14980
rect 3329 14971 3387 14977
rect 4065 14977 4077 14980
rect 4111 14977 4123 15011
rect 7098 15008 7104 15020
rect 7059 14980 7104 15008
rect 4065 14971 4123 14977
rect 7098 14968 7104 14980
rect 7156 14968 7162 15020
rect 9125 15011 9183 15017
rect 9125 14977 9137 15011
rect 9171 15008 9183 15011
rect 13170 15008 13176 15020
rect 9171 14980 13176 15008
rect 9171 14977 9183 14980
rect 9125 14971 9183 14977
rect 13170 14968 13176 14980
rect 13228 14968 13234 15020
rect 1394 14900 1400 14952
rect 1452 14940 1458 14952
rect 1673 14943 1731 14949
rect 1673 14940 1685 14943
rect 1452 14912 1685 14940
rect 1452 14900 1458 14912
rect 1673 14909 1685 14912
rect 1719 14909 1731 14943
rect 1946 14940 1952 14952
rect 1907 14912 1952 14940
rect 1673 14903 1731 14909
rect 1946 14900 1952 14912
rect 2004 14900 2010 14952
rect 2682 14900 2688 14952
rect 2740 14940 2746 14952
rect 3789 14943 3847 14949
rect 3789 14940 3801 14943
rect 2740 14912 3801 14940
rect 2740 14900 2746 14912
rect 3789 14909 3801 14912
rect 3835 14909 3847 14943
rect 3789 14903 3847 14909
rect 5997 14943 6055 14949
rect 5997 14909 6009 14943
rect 6043 14909 6055 14943
rect 6822 14940 6828 14952
rect 6783 14912 6828 14940
rect 5997 14903 6055 14909
rect 6012 14872 6040 14903
rect 6822 14900 6828 14912
rect 6880 14900 6886 14952
rect 7558 14940 7564 14952
rect 6932 14912 7564 14940
rect 6932 14872 6960 14912
rect 7558 14900 7564 14912
rect 7616 14900 7622 14952
rect 8846 14900 8852 14952
rect 8904 14940 8910 14952
rect 9309 14943 9367 14949
rect 9309 14940 9321 14943
rect 8904 14912 9321 14940
rect 8904 14900 8910 14912
rect 9309 14909 9321 14912
rect 9355 14909 9367 14943
rect 9766 14940 9772 14952
rect 9727 14912 9772 14940
rect 9309 14903 9367 14909
rect 6012 14844 6960 14872
rect 6181 14807 6239 14813
rect 6181 14773 6193 14807
rect 6227 14804 6239 14807
rect 6730 14804 6736 14816
rect 6227 14776 6736 14804
rect 6227 14773 6239 14776
rect 6181 14767 6239 14773
rect 6730 14764 6736 14776
rect 6788 14764 6794 14816
rect 6914 14764 6920 14816
rect 6972 14804 6978 14816
rect 9214 14804 9220 14816
rect 6972 14776 9220 14804
rect 6972 14764 6978 14776
rect 9214 14764 9220 14776
rect 9272 14764 9278 14816
rect 9324 14804 9352 14903
rect 9766 14900 9772 14912
rect 9824 14900 9830 14952
rect 10686 14940 10692 14952
rect 10647 14912 10692 14940
rect 10686 14900 10692 14912
rect 10744 14900 10750 14952
rect 11054 14940 11060 14952
rect 11015 14912 11060 14940
rect 11054 14900 11060 14912
rect 11112 14900 11118 14952
rect 11330 14940 11336 14952
rect 11291 14912 11336 14940
rect 11330 14900 11336 14912
rect 11388 14900 11394 14952
rect 12066 14940 12072 14952
rect 12027 14912 12072 14940
rect 12066 14900 12072 14912
rect 12124 14900 12130 14952
rect 12434 14900 12440 14952
rect 12492 14940 12498 14952
rect 13372 14949 13400 15048
rect 13814 15036 13820 15048
rect 13872 15036 13878 15088
rect 30006 15036 30012 15088
rect 30064 15036 30070 15088
rect 13449 15011 13507 15017
rect 13449 14977 13461 15011
rect 13495 15008 13507 15011
rect 14090 15008 14096 15020
rect 13495 14980 14096 15008
rect 13495 14977 13507 14980
rect 13449 14971 13507 14977
rect 14090 14968 14096 14980
rect 14148 14968 14154 15020
rect 14277 15011 14335 15017
rect 14277 14977 14289 15011
rect 14323 15008 14335 15011
rect 16577 15011 16635 15017
rect 14323 14980 14688 15008
rect 14323 14977 14335 14980
rect 14277 14971 14335 14977
rect 13357 14943 13415 14949
rect 12492 14912 12537 14940
rect 12492 14900 12498 14912
rect 13357 14909 13369 14943
rect 13403 14909 13415 14943
rect 13357 14903 13415 14909
rect 13725 14943 13783 14949
rect 13725 14909 13737 14943
rect 13771 14940 13783 14943
rect 13998 14940 14004 14952
rect 13771 14912 14004 14940
rect 13771 14909 13783 14912
rect 13725 14903 13783 14909
rect 13998 14900 14004 14912
rect 14056 14900 14062 14952
rect 14550 14940 14556 14952
rect 14511 14912 14556 14940
rect 14550 14900 14556 14912
rect 14608 14900 14614 14952
rect 14660 14940 14688 14980
rect 16577 14977 16589 15011
rect 16623 15008 16635 15011
rect 17034 15008 17040 15020
rect 16623 14980 17040 15008
rect 16623 14977 16635 14980
rect 16577 14971 16635 14977
rect 17034 14968 17040 14980
rect 17092 14968 17098 15020
rect 18322 14968 18328 15020
rect 18380 15008 18386 15020
rect 19429 15011 19487 15017
rect 19429 15008 19441 15011
rect 18380 14980 19441 15008
rect 18380 14968 18386 14980
rect 19429 14977 19441 14980
rect 19475 14977 19487 15011
rect 20162 15008 20168 15020
rect 19429 14971 19487 14977
rect 19812 14980 20168 15008
rect 15286 14940 15292 14952
rect 14660 14912 15292 14940
rect 15286 14900 15292 14912
rect 15344 14940 15350 14952
rect 16758 14940 16764 14952
rect 15344 14912 16764 14940
rect 15344 14900 15350 14912
rect 16758 14900 16764 14912
rect 16816 14900 16822 14952
rect 16942 14940 16948 14952
rect 16903 14912 16948 14940
rect 16942 14900 16948 14912
rect 17000 14900 17006 14952
rect 17221 14943 17279 14949
rect 17221 14909 17233 14943
rect 17267 14909 17279 14943
rect 18230 14940 18236 14952
rect 18191 14912 18236 14940
rect 17221 14903 17279 14909
rect 9398 14832 9404 14884
rect 9456 14872 9462 14884
rect 10045 14875 10103 14881
rect 10045 14872 10057 14875
rect 9456 14844 10057 14872
rect 9456 14832 9462 14844
rect 10045 14841 10057 14844
rect 10091 14841 10103 14875
rect 17236 14872 17264 14903
rect 18230 14900 18236 14912
rect 18288 14900 18294 14952
rect 18693 14943 18751 14949
rect 18693 14909 18705 14943
rect 18739 14909 18751 14943
rect 19334 14940 19340 14952
rect 19295 14912 19340 14940
rect 18693 14903 18751 14909
rect 10045 14835 10103 14841
rect 15212 14844 17264 14872
rect 17497 14875 17555 14881
rect 11238 14804 11244 14816
rect 9324 14776 11244 14804
rect 11238 14764 11244 14776
rect 11296 14764 11302 14816
rect 11330 14764 11336 14816
rect 11388 14804 11394 14816
rect 11790 14804 11796 14816
rect 11388 14776 11796 14804
rect 11388 14764 11394 14776
rect 11790 14764 11796 14776
rect 11848 14804 11854 14816
rect 12529 14807 12587 14813
rect 12529 14804 12541 14807
rect 11848 14776 12541 14804
rect 11848 14764 11854 14776
rect 12529 14773 12541 14776
rect 12575 14773 12587 14807
rect 12529 14767 12587 14773
rect 13538 14764 13544 14816
rect 13596 14804 13602 14816
rect 15212 14804 15240 14844
rect 17497 14841 17509 14875
rect 17543 14872 17555 14875
rect 18046 14872 18052 14884
rect 17543 14844 18052 14872
rect 17543 14841 17555 14844
rect 17497 14835 17555 14841
rect 18046 14832 18052 14844
rect 18104 14832 18110 14884
rect 18708 14872 18736 14903
rect 19334 14900 19340 14912
rect 19392 14900 19398 14952
rect 19812 14949 19840 14980
rect 20162 14968 20168 14980
rect 20220 14968 20226 15020
rect 21266 15008 21272 15020
rect 20548 14980 21272 15008
rect 19797 14943 19855 14949
rect 19797 14909 19809 14943
rect 19843 14909 19855 14943
rect 19797 14903 19855 14909
rect 20349 14943 20407 14949
rect 20349 14909 20361 14943
rect 20395 14940 20407 14943
rect 20548 14940 20576 14980
rect 21266 14968 21272 14980
rect 21324 14968 21330 15020
rect 24302 14968 24308 15020
rect 24360 15008 24366 15020
rect 24397 15011 24455 15017
rect 24397 15008 24409 15011
rect 24360 14980 24409 15008
rect 24360 14968 24366 14980
rect 24397 14977 24409 14980
rect 24443 14977 24455 15011
rect 24397 14971 24455 14977
rect 24486 14968 24492 15020
rect 24544 15008 24550 15020
rect 24762 15008 24768 15020
rect 24544 14980 24768 15008
rect 24544 14968 24550 14980
rect 24762 14968 24768 14980
rect 24820 15008 24826 15020
rect 26237 15011 26295 15017
rect 26237 15008 26249 15011
rect 24820 14980 26249 15008
rect 24820 14968 24826 14980
rect 26237 14977 26249 14980
rect 26283 14977 26295 15011
rect 26510 15008 26516 15020
rect 26471 14980 26516 15008
rect 26237 14971 26295 14977
rect 26510 14968 26516 14980
rect 26568 14968 26574 15020
rect 28902 14968 28908 15020
rect 28960 15008 28966 15020
rect 29457 15011 29515 15017
rect 29457 15008 29469 15011
rect 28960 14980 29469 15008
rect 28960 14968 28966 14980
rect 29457 14977 29469 14980
rect 29503 14977 29515 15011
rect 30024 15008 30052 15036
rect 30469 15011 30527 15017
rect 30469 15008 30481 15011
rect 30024 14980 30481 15008
rect 29457 14971 29515 14977
rect 30469 14977 30481 14980
rect 30515 14977 30527 15011
rect 31570 15008 31576 15020
rect 30469 14971 30527 14977
rect 30576 14980 31576 15008
rect 30576 14952 30604 14980
rect 31570 14968 31576 14980
rect 31628 14968 31634 15020
rect 33042 15008 33048 15020
rect 33003 14980 33048 15008
rect 33042 14968 33048 14980
rect 33100 14968 33106 15020
rect 37366 14968 37372 15020
rect 37424 15008 37430 15020
rect 37461 15011 37519 15017
rect 37461 15008 37473 15011
rect 37424 14980 37473 15008
rect 37424 14968 37430 14980
rect 37461 14977 37473 14980
rect 37507 14977 37519 15011
rect 37461 14971 37519 14977
rect 20714 14940 20720 14952
rect 20395 14912 20576 14940
rect 20675 14912 20720 14940
rect 20395 14909 20407 14912
rect 20349 14903 20407 14909
rect 20714 14900 20720 14912
rect 20772 14900 20778 14952
rect 20990 14940 20996 14952
rect 20951 14912 20996 14940
rect 20990 14900 20996 14912
rect 21048 14900 21054 14952
rect 21082 14900 21088 14952
rect 21140 14940 21146 14952
rect 21729 14943 21787 14949
rect 21729 14940 21741 14943
rect 21140 14912 21741 14940
rect 21140 14900 21146 14912
rect 21729 14909 21741 14912
rect 21775 14909 21787 14943
rect 22922 14940 22928 14952
rect 22883 14912 22928 14940
rect 21729 14903 21787 14909
rect 22922 14900 22928 14912
rect 22980 14900 22986 14952
rect 24118 14940 24124 14952
rect 24079 14912 24124 14940
rect 24118 14900 24124 14912
rect 24176 14900 24182 14952
rect 24854 14900 24860 14952
rect 24912 14940 24918 14952
rect 24912 14912 29040 14940
rect 24912 14900 24918 14912
rect 22830 14872 22836 14884
rect 18708 14844 22836 14872
rect 22830 14832 22836 14844
rect 22888 14832 22894 14884
rect 27890 14872 27896 14884
rect 27803 14844 27896 14872
rect 27890 14832 27896 14844
rect 27948 14872 27954 14884
rect 28350 14872 28356 14884
rect 27948 14844 28356 14872
rect 27948 14832 27954 14844
rect 28350 14832 28356 14844
rect 28408 14832 28414 14884
rect 13596 14776 15240 14804
rect 15841 14807 15899 14813
rect 13596 14764 13602 14776
rect 15841 14773 15853 14807
rect 15887 14804 15899 14807
rect 17126 14804 17132 14816
rect 15887 14776 17132 14804
rect 15887 14773 15899 14776
rect 15841 14767 15899 14773
rect 17126 14764 17132 14776
rect 17184 14764 17190 14816
rect 17402 14764 17408 14816
rect 17460 14804 17466 14816
rect 18233 14807 18291 14813
rect 18233 14804 18245 14807
rect 17460 14776 18245 14804
rect 17460 14764 17466 14776
rect 18233 14773 18245 14776
rect 18279 14773 18291 14807
rect 18233 14767 18291 14773
rect 22094 14764 22100 14816
rect 22152 14804 22158 14816
rect 23014 14804 23020 14816
rect 22152 14776 23020 14804
rect 22152 14764 22158 14776
rect 23014 14764 23020 14776
rect 23072 14764 23078 14816
rect 25685 14807 25743 14813
rect 25685 14773 25697 14807
rect 25731 14804 25743 14807
rect 26602 14804 26608 14816
rect 25731 14776 26608 14804
rect 25731 14773 25743 14776
rect 25685 14767 25743 14773
rect 26602 14764 26608 14776
rect 26660 14764 26666 14816
rect 28902 14764 28908 14816
rect 28960 14804 28966 14816
rect 29012 14804 29040 14912
rect 29178 14900 29184 14952
rect 29236 14940 29242 14952
rect 30009 14943 30067 14949
rect 30009 14940 30021 14943
rect 29236 14912 30021 14940
rect 29236 14900 29242 14912
rect 30009 14909 30021 14912
rect 30055 14940 30067 14943
rect 30098 14940 30104 14952
rect 30055 14912 30104 14940
rect 30055 14909 30067 14912
rect 30009 14903 30067 14909
rect 30098 14900 30104 14912
rect 30156 14900 30162 14952
rect 30285 14943 30343 14949
rect 30285 14909 30297 14943
rect 30331 14940 30343 14943
rect 30558 14940 30564 14952
rect 30331 14912 30564 14940
rect 30331 14909 30343 14912
rect 30285 14903 30343 14909
rect 30558 14900 30564 14912
rect 30616 14900 30622 14952
rect 30742 14900 30748 14952
rect 30800 14940 30806 14952
rect 31297 14943 31355 14949
rect 31297 14940 31309 14943
rect 30800 14912 31309 14940
rect 30800 14900 30806 14912
rect 31297 14909 31309 14912
rect 31343 14940 31355 14943
rect 31662 14940 31668 14952
rect 31343 14912 31668 14940
rect 31343 14909 31355 14912
rect 31297 14903 31355 14909
rect 31662 14900 31668 14912
rect 31720 14900 31726 14952
rect 32306 14940 32312 14952
rect 32267 14912 32312 14940
rect 32306 14900 32312 14912
rect 32364 14900 32370 14952
rect 32401 14943 32459 14949
rect 32401 14909 32413 14943
rect 32447 14909 32459 14943
rect 32766 14940 32772 14952
rect 32727 14912 32772 14940
rect 32401 14903 32459 14909
rect 32214 14832 32220 14884
rect 32272 14872 32278 14884
rect 32416 14872 32444 14903
rect 32766 14900 32772 14912
rect 32824 14900 32830 14952
rect 33505 14943 33563 14949
rect 33505 14909 33517 14943
rect 33551 14940 33563 14943
rect 33594 14940 33600 14952
rect 33551 14912 33600 14940
rect 33551 14909 33563 14912
rect 33505 14903 33563 14909
rect 33594 14900 33600 14912
rect 33652 14900 33658 14952
rect 33778 14900 33784 14952
rect 33836 14940 33842 14952
rect 33965 14943 34023 14949
rect 33965 14940 33977 14943
rect 33836 14912 33977 14940
rect 33836 14900 33842 14912
rect 33965 14909 33977 14912
rect 34011 14909 34023 14943
rect 33965 14903 34023 14909
rect 35897 14943 35955 14949
rect 35897 14909 35909 14943
rect 35943 14909 35955 14943
rect 36078 14940 36084 14952
rect 36039 14912 36084 14940
rect 35897 14903 35955 14909
rect 32272 14844 32444 14872
rect 35437 14875 35495 14881
rect 32272 14832 32278 14844
rect 35437 14841 35449 14875
rect 35483 14872 35495 14875
rect 35802 14872 35808 14884
rect 35483 14844 35808 14872
rect 35483 14841 35495 14844
rect 35437 14835 35495 14841
rect 35802 14832 35808 14844
rect 35860 14832 35866 14884
rect 34514 14804 34520 14816
rect 28960 14776 34520 14804
rect 28960 14764 28966 14776
rect 34514 14764 34520 14776
rect 34572 14764 34578 14816
rect 35912 14804 35940 14903
rect 36078 14900 36084 14912
rect 36136 14900 36142 14952
rect 36262 14940 36268 14952
rect 36223 14912 36268 14940
rect 36262 14900 36268 14912
rect 36320 14900 36326 14952
rect 37734 14940 37740 14952
rect 37695 14912 37740 14940
rect 37734 14900 37740 14912
rect 37792 14900 37798 14952
rect 38470 14804 38476 14816
rect 35912 14776 38476 14804
rect 38470 14764 38476 14776
rect 38528 14764 38534 14816
rect 1104 14714 39836 14736
rect 1104 14662 19606 14714
rect 19658 14662 19670 14714
rect 19722 14662 19734 14714
rect 19786 14662 19798 14714
rect 19850 14662 39836 14714
rect 1104 14640 39836 14662
rect 1946 14560 1952 14612
rect 2004 14600 2010 14612
rect 2777 14603 2835 14609
rect 2777 14600 2789 14603
rect 2004 14572 2789 14600
rect 2004 14560 2010 14572
rect 2777 14569 2789 14572
rect 2823 14569 2835 14603
rect 2777 14563 2835 14569
rect 9490 14560 9496 14612
rect 9548 14600 9554 14612
rect 13538 14600 13544 14612
rect 9548 14572 13400 14600
rect 13499 14572 13544 14600
rect 9548 14560 9554 14572
rect 10686 14532 10692 14544
rect 9048 14504 10692 14532
rect 1670 14464 1676 14476
rect 1631 14436 1676 14464
rect 1670 14424 1676 14436
rect 1728 14424 1734 14476
rect 3878 14464 3884 14476
rect 3839 14436 3884 14464
rect 3878 14424 3884 14436
rect 3936 14424 3942 14476
rect 6181 14467 6239 14473
rect 6181 14433 6193 14467
rect 6227 14464 6239 14467
rect 6914 14464 6920 14476
rect 6227 14436 6920 14464
rect 6227 14433 6239 14436
rect 6181 14427 6239 14433
rect 6914 14424 6920 14436
rect 6972 14424 6978 14476
rect 8665 14467 8723 14473
rect 8665 14433 8677 14467
rect 8711 14464 8723 14467
rect 9048 14464 9076 14504
rect 10686 14492 10692 14504
rect 10744 14492 10750 14544
rect 8711 14436 9076 14464
rect 8711 14433 8723 14436
rect 8665 14427 8723 14433
rect 9048 14408 9076 14436
rect 9125 14467 9183 14473
rect 9125 14433 9137 14467
rect 9171 14464 9183 14467
rect 9950 14464 9956 14476
rect 9171 14436 9956 14464
rect 9171 14433 9183 14436
rect 9125 14427 9183 14433
rect 9950 14424 9956 14436
rect 10008 14424 10014 14476
rect 10042 14424 10048 14476
rect 10100 14464 10106 14476
rect 10410 14464 10416 14476
rect 10100 14436 10145 14464
rect 10371 14436 10416 14464
rect 10100 14424 10106 14436
rect 10410 14424 10416 14436
rect 10468 14424 10474 14476
rect 11333 14467 11391 14473
rect 11333 14433 11345 14467
rect 11379 14464 11391 14467
rect 11422 14464 11428 14476
rect 11379 14436 11428 14464
rect 11379 14433 11391 14436
rect 11333 14427 11391 14433
rect 11422 14424 11428 14436
rect 11480 14424 11486 14476
rect 11606 14464 11612 14476
rect 11567 14436 11612 14464
rect 11606 14424 11612 14436
rect 11664 14424 11670 14476
rect 13372 14464 13400 14572
rect 13538 14560 13544 14572
rect 13596 14560 13602 14612
rect 14550 14560 14556 14612
rect 14608 14600 14614 14612
rect 16485 14603 16543 14609
rect 16485 14600 16497 14603
rect 14608 14572 16497 14600
rect 14608 14560 14614 14572
rect 16485 14569 16497 14572
rect 16531 14569 16543 14603
rect 16485 14563 16543 14569
rect 17957 14603 18015 14609
rect 17957 14569 17969 14603
rect 18003 14600 18015 14603
rect 18003 14572 22876 14600
rect 18003 14569 18015 14572
rect 17957 14563 18015 14569
rect 17221 14535 17279 14541
rect 17221 14532 17233 14535
rect 15948 14504 17233 14532
rect 15948 14476 15976 14504
rect 17221 14501 17233 14504
rect 17267 14501 17279 14535
rect 22848 14532 22876 14572
rect 22922 14560 22928 14612
rect 22980 14600 22986 14612
rect 23293 14603 23351 14609
rect 23293 14600 23305 14603
rect 22980 14572 23305 14600
rect 22980 14560 22986 14572
rect 23293 14569 23305 14572
rect 23339 14569 23351 14603
rect 24670 14600 24676 14612
rect 23293 14563 23351 14569
rect 23400 14572 24676 14600
rect 23400 14532 23428 14572
rect 24670 14560 24676 14572
rect 24728 14600 24734 14612
rect 27798 14600 27804 14612
rect 24728 14572 27804 14600
rect 24728 14560 24734 14572
rect 27798 14560 27804 14572
rect 27856 14560 27862 14612
rect 29822 14560 29828 14612
rect 29880 14600 29886 14612
rect 29880 14572 31340 14600
rect 29880 14560 29886 14572
rect 22848 14504 23428 14532
rect 17221 14495 17279 14501
rect 28074 14492 28080 14544
rect 28132 14532 28138 14544
rect 31202 14532 31208 14544
rect 28132 14504 31208 14532
rect 28132 14492 28138 14504
rect 28552 14476 28580 14504
rect 31202 14492 31208 14504
rect 31260 14492 31266 14544
rect 13538 14464 13544 14476
rect 13372 14436 13544 14464
rect 13538 14424 13544 14436
rect 13596 14424 13602 14476
rect 13633 14467 13691 14473
rect 13633 14433 13645 14467
rect 13679 14464 13691 14467
rect 13722 14464 13728 14476
rect 13679 14436 13728 14464
rect 13679 14433 13691 14436
rect 13633 14427 13691 14433
rect 13722 14424 13728 14436
rect 13780 14424 13786 14476
rect 13906 14424 13912 14476
rect 13964 14464 13970 14476
rect 14001 14467 14059 14473
rect 14001 14464 14013 14467
rect 13964 14436 14013 14464
rect 13964 14424 13970 14436
rect 14001 14433 14013 14436
rect 14047 14433 14059 14467
rect 14001 14427 14059 14433
rect 15378 14424 15384 14476
rect 15436 14464 15442 14476
rect 15473 14467 15531 14473
rect 15473 14464 15485 14467
rect 15436 14436 15485 14464
rect 15436 14424 15442 14436
rect 15473 14433 15485 14436
rect 15519 14433 15531 14467
rect 15473 14427 15531 14433
rect 15565 14467 15623 14473
rect 15565 14433 15577 14467
rect 15611 14464 15623 14467
rect 15654 14464 15660 14476
rect 15611 14436 15660 14464
rect 15611 14433 15623 14436
rect 15565 14427 15623 14433
rect 15654 14424 15660 14436
rect 15712 14424 15718 14476
rect 15930 14464 15936 14476
rect 15891 14436 15936 14464
rect 15930 14424 15936 14436
rect 15988 14424 15994 14476
rect 16025 14467 16083 14473
rect 16025 14433 16037 14467
rect 16071 14464 16083 14467
rect 17126 14464 17132 14476
rect 16071 14436 16988 14464
rect 17087 14436 17132 14464
rect 16071 14433 16083 14436
rect 16025 14427 16083 14433
rect 1394 14396 1400 14408
rect 1355 14368 1400 14396
rect 1394 14356 1400 14368
rect 1452 14356 1458 14408
rect 4062 14396 4068 14408
rect 4023 14368 4068 14396
rect 4062 14356 4068 14368
rect 4120 14356 4126 14408
rect 4341 14399 4399 14405
rect 4341 14365 4353 14399
rect 4387 14396 4399 14399
rect 5626 14396 5632 14408
rect 4387 14368 5632 14396
rect 4387 14365 4399 14368
rect 4341 14359 4399 14365
rect 5626 14356 5632 14368
rect 5684 14356 5690 14408
rect 6454 14396 6460 14408
rect 6415 14368 6460 14396
rect 6454 14356 6460 14368
rect 6512 14356 6518 14408
rect 8757 14399 8815 14405
rect 8757 14365 8769 14399
rect 8803 14365 8815 14399
rect 8757 14359 8815 14365
rect 5074 14288 5080 14340
rect 5132 14328 5138 14340
rect 5445 14331 5503 14337
rect 5445 14328 5457 14331
rect 5132 14300 5457 14328
rect 5132 14288 5138 14300
rect 5445 14297 5457 14300
rect 5491 14297 5503 14331
rect 8772 14328 8800 14359
rect 9030 14356 9036 14408
rect 9088 14356 9094 14408
rect 9766 14396 9772 14408
rect 9727 14368 9772 14396
rect 9766 14356 9772 14368
rect 9824 14356 9830 14408
rect 12434 14356 12440 14408
rect 12492 14396 12498 14408
rect 12989 14399 13047 14405
rect 12989 14396 13001 14399
rect 12492 14368 13001 14396
rect 12492 14356 12498 14368
rect 12989 14365 13001 14368
rect 13035 14396 13047 14399
rect 14277 14399 14335 14405
rect 14277 14396 14289 14399
rect 13035 14368 14289 14396
rect 13035 14365 13047 14368
rect 12989 14359 13047 14365
rect 14277 14365 14289 14368
rect 14323 14365 14335 14399
rect 16960 14396 16988 14436
rect 17126 14424 17132 14436
rect 17184 14424 17190 14476
rect 18138 14464 18144 14476
rect 17972 14436 18144 14464
rect 17972 14396 18000 14436
rect 18138 14424 18144 14436
rect 18196 14424 18202 14476
rect 18322 14464 18328 14476
rect 18283 14436 18328 14464
rect 18322 14424 18328 14436
rect 18380 14424 18386 14476
rect 19426 14424 19432 14476
rect 19484 14464 19490 14476
rect 20165 14467 20223 14473
rect 20165 14464 20177 14467
rect 19484 14436 20177 14464
rect 19484 14424 19490 14436
rect 20165 14433 20177 14436
rect 20211 14433 20223 14467
rect 22186 14464 22192 14476
rect 22147 14436 22192 14464
rect 20165 14427 20223 14433
rect 22186 14424 22192 14436
rect 22244 14424 22250 14476
rect 24394 14464 24400 14476
rect 24355 14436 24400 14464
rect 24394 14424 24400 14436
rect 24452 14424 24458 14476
rect 26602 14464 26608 14476
rect 26563 14436 26608 14464
rect 26602 14424 26608 14436
rect 26660 14424 26666 14476
rect 27706 14424 27712 14476
rect 27764 14464 27770 14476
rect 27801 14467 27859 14473
rect 27801 14464 27813 14467
rect 27764 14436 27813 14464
rect 27764 14424 27770 14436
rect 27801 14433 27813 14436
rect 27847 14433 27859 14467
rect 27801 14427 27859 14433
rect 28258 14424 28264 14476
rect 28316 14464 28322 14476
rect 28353 14467 28411 14473
rect 28353 14464 28365 14467
rect 28316 14436 28365 14464
rect 28316 14424 28322 14436
rect 28353 14433 28365 14436
rect 28399 14433 28411 14467
rect 28534 14464 28540 14476
rect 28447 14436 28540 14464
rect 28353 14427 28411 14433
rect 16960 14368 18000 14396
rect 18049 14399 18107 14405
rect 14277 14359 14335 14365
rect 18049 14365 18061 14399
rect 18095 14365 18107 14399
rect 18156 14396 18184 14424
rect 19150 14396 19156 14408
rect 18156 14368 19156 14396
rect 18049 14359 18107 14365
rect 11146 14328 11152 14340
rect 8772 14300 11152 14328
rect 5445 14291 5503 14297
rect 11146 14288 11152 14300
rect 11204 14288 11210 14340
rect 16206 14288 16212 14340
rect 16264 14328 16270 14340
rect 16758 14328 16764 14340
rect 16264 14300 16764 14328
rect 16264 14288 16270 14300
rect 16758 14288 16764 14300
rect 16816 14328 16822 14340
rect 18064 14328 18092 14359
rect 19150 14356 19156 14368
rect 19208 14356 19214 14408
rect 21913 14399 21971 14405
rect 21913 14365 21925 14399
rect 21959 14365 21971 14399
rect 21913 14359 21971 14365
rect 21928 14328 21956 14359
rect 23474 14356 23480 14408
rect 23532 14396 23538 14408
rect 24118 14396 24124 14408
rect 23532 14368 24124 14396
rect 23532 14356 23538 14368
rect 24118 14356 24124 14368
rect 24176 14356 24182 14408
rect 26142 14356 26148 14408
rect 26200 14396 26206 14408
rect 26513 14399 26571 14405
rect 26513 14396 26525 14399
rect 26200 14368 26525 14396
rect 26200 14356 26206 14368
rect 26513 14365 26525 14368
rect 26559 14365 26571 14399
rect 26513 14359 26571 14365
rect 27614 14356 27620 14408
rect 27672 14396 27678 14408
rect 28074 14396 28080 14408
rect 27672 14368 28080 14396
rect 27672 14356 27678 14368
rect 28074 14356 28080 14368
rect 28132 14356 28138 14408
rect 16816 14300 18092 14328
rect 16816 14288 16822 14300
rect 3697 14263 3755 14269
rect 3697 14229 3709 14263
rect 3743 14260 3755 14263
rect 4706 14260 4712 14272
rect 3743 14232 4712 14260
rect 3743 14229 3755 14232
rect 3697 14223 3755 14229
rect 4706 14220 4712 14232
rect 4764 14260 4770 14272
rect 6546 14260 6552 14272
rect 4764 14232 6552 14260
rect 4764 14220 4770 14232
rect 6546 14220 6552 14232
rect 6604 14220 6610 14272
rect 7742 14260 7748 14272
rect 7703 14232 7748 14260
rect 7742 14220 7748 14232
rect 7800 14220 7806 14272
rect 8754 14220 8760 14272
rect 8812 14260 8818 14272
rect 17957 14263 18015 14269
rect 17957 14260 17969 14263
rect 8812 14232 17969 14260
rect 8812 14220 8818 14232
rect 17957 14229 17969 14232
rect 18003 14229 18015 14263
rect 18064 14260 18092 14300
rect 19168 14300 21956 14328
rect 19168 14272 19196 14300
rect 19150 14260 19156 14272
rect 18064 14232 19156 14260
rect 17957 14223 18015 14229
rect 19150 14220 19156 14232
rect 19208 14220 19214 14272
rect 19426 14260 19432 14272
rect 19387 14232 19432 14260
rect 19426 14220 19432 14232
rect 19484 14220 19490 14272
rect 20162 14220 20168 14272
rect 20220 14260 20226 14272
rect 20257 14263 20315 14269
rect 20257 14260 20269 14263
rect 20220 14232 20269 14260
rect 20220 14220 20226 14232
rect 20257 14229 20269 14232
rect 20303 14260 20315 14263
rect 24118 14260 24124 14272
rect 20303 14232 24124 14260
rect 20303 14229 20315 14232
rect 20257 14223 20315 14229
rect 24118 14220 24124 14232
rect 24176 14220 24182 14272
rect 25038 14220 25044 14272
rect 25096 14260 25102 14272
rect 25501 14263 25559 14269
rect 25501 14260 25513 14263
rect 25096 14232 25513 14260
rect 25096 14220 25102 14232
rect 25501 14229 25513 14232
rect 25547 14229 25559 14263
rect 26786 14260 26792 14272
rect 26747 14232 26792 14260
rect 25501 14223 25559 14229
rect 26786 14220 26792 14232
rect 26844 14220 26850 14272
rect 26878 14220 26884 14272
rect 26936 14260 26942 14272
rect 27893 14263 27951 14269
rect 27893 14260 27905 14263
rect 26936 14232 27905 14260
rect 26936 14220 26942 14232
rect 27893 14229 27905 14232
rect 27939 14229 27951 14263
rect 28368 14260 28396 14427
rect 28534 14424 28540 14436
rect 28592 14424 28598 14476
rect 29086 14464 29092 14476
rect 29047 14436 29092 14464
rect 29086 14424 29092 14436
rect 29144 14424 29150 14476
rect 30006 14424 30012 14476
rect 30064 14464 30070 14476
rect 31312 14473 31340 14572
rect 34330 14560 34336 14612
rect 34388 14600 34394 14612
rect 34977 14603 35035 14609
rect 34977 14600 34989 14603
rect 34388 14572 34989 14600
rect 34388 14560 34394 14572
rect 34977 14569 34989 14572
rect 35023 14569 35035 14603
rect 34977 14563 35035 14569
rect 37734 14560 37740 14612
rect 37792 14600 37798 14612
rect 37829 14603 37887 14609
rect 37829 14600 37841 14603
rect 37792 14572 37841 14600
rect 37792 14560 37798 14572
rect 37829 14569 37841 14572
rect 37875 14569 37887 14603
rect 37829 14563 37887 14569
rect 31570 14492 31576 14544
rect 31628 14532 31634 14544
rect 31628 14504 32996 14532
rect 31628 14492 31634 14504
rect 30101 14467 30159 14473
rect 30101 14464 30113 14467
rect 30064 14436 30113 14464
rect 30064 14424 30070 14436
rect 30101 14433 30113 14436
rect 30147 14433 30159 14467
rect 30101 14427 30159 14433
rect 30653 14467 30711 14473
rect 30653 14433 30665 14467
rect 30699 14433 30711 14467
rect 30653 14427 30711 14433
rect 31297 14467 31355 14473
rect 31297 14433 31309 14467
rect 31343 14433 31355 14467
rect 32122 14464 32128 14476
rect 31297 14427 31355 14433
rect 31404 14436 31984 14464
rect 32083 14436 32128 14464
rect 29917 14399 29975 14405
rect 29917 14365 29929 14399
rect 29963 14396 29975 14399
rect 30282 14396 30288 14408
rect 29963 14368 30288 14396
rect 29963 14365 29975 14368
rect 29917 14359 29975 14365
rect 30282 14356 30288 14368
rect 30340 14356 30346 14408
rect 30668 14396 30696 14427
rect 31404 14396 31432 14436
rect 30668 14368 31432 14396
rect 31956 14396 31984 14436
rect 32122 14424 32128 14436
rect 32180 14424 32186 14476
rect 32968 14473 32996 14504
rect 32953 14467 33011 14473
rect 32953 14433 32965 14467
rect 32999 14433 33011 14467
rect 32953 14427 33011 14433
rect 33597 14467 33655 14473
rect 33597 14433 33609 14467
rect 33643 14464 33655 14467
rect 34606 14464 34612 14476
rect 33643 14436 34612 14464
rect 33643 14433 33655 14436
rect 33597 14427 33655 14433
rect 34606 14424 34612 14436
rect 34664 14464 34670 14476
rect 35526 14464 35532 14476
rect 34664 14436 35532 14464
rect 34664 14424 34670 14436
rect 35526 14424 35532 14436
rect 35584 14424 35590 14476
rect 35713 14467 35771 14473
rect 35713 14433 35725 14467
rect 35759 14433 35771 14467
rect 35713 14427 35771 14433
rect 33318 14396 33324 14408
rect 31956 14368 33324 14396
rect 33318 14356 33324 14368
rect 33376 14356 33382 14408
rect 33870 14396 33876 14408
rect 33831 14368 33876 14396
rect 33870 14356 33876 14368
rect 33928 14356 33934 14408
rect 34054 14356 34060 14408
rect 34112 14396 34118 14408
rect 35728 14396 35756 14427
rect 35802 14424 35808 14476
rect 35860 14464 35866 14476
rect 36265 14467 36323 14473
rect 36265 14464 36277 14467
rect 35860 14436 36277 14464
rect 35860 14424 35866 14436
rect 36265 14433 36277 14436
rect 36311 14433 36323 14467
rect 36538 14464 36544 14476
rect 36499 14436 36544 14464
rect 36265 14427 36323 14433
rect 36538 14424 36544 14436
rect 36596 14424 36602 14476
rect 37734 14464 37740 14476
rect 37695 14436 37740 14464
rect 37734 14424 37740 14436
rect 37792 14424 37798 14476
rect 37826 14424 37832 14476
rect 37884 14464 37890 14476
rect 38289 14467 38347 14473
rect 38289 14464 38301 14467
rect 37884 14436 38301 14464
rect 37884 14424 37890 14436
rect 38289 14433 38301 14436
rect 38335 14433 38347 14467
rect 38289 14427 38347 14433
rect 38562 14396 38568 14408
rect 34112 14368 35756 14396
rect 38523 14368 38568 14396
rect 34112 14356 34118 14368
rect 38562 14356 38568 14368
rect 38620 14356 38626 14408
rect 29362 14288 29368 14340
rect 29420 14328 29426 14340
rect 30561 14331 30619 14337
rect 30561 14328 30573 14331
rect 29420 14300 30573 14328
rect 29420 14288 29426 14300
rect 30561 14297 30573 14300
rect 30607 14297 30619 14331
rect 30561 14291 30619 14297
rect 31202 14288 31208 14340
rect 31260 14328 31266 14340
rect 31481 14331 31539 14337
rect 31481 14328 31493 14331
rect 31260 14300 31493 14328
rect 31260 14288 31266 14300
rect 31481 14297 31493 14300
rect 31527 14328 31539 14331
rect 32766 14328 32772 14340
rect 31527 14300 32772 14328
rect 31527 14297 31539 14300
rect 31481 14291 31539 14297
rect 32766 14288 32772 14300
rect 32824 14288 32830 14340
rect 35802 14328 35808 14340
rect 35763 14300 35808 14328
rect 35802 14288 35808 14300
rect 35860 14288 35866 14340
rect 30098 14260 30104 14272
rect 28368 14232 30104 14260
rect 27893 14223 27951 14229
rect 30098 14220 30104 14232
rect 30156 14220 30162 14272
rect 32309 14263 32367 14269
rect 32309 14229 32321 14263
rect 32355 14260 32367 14263
rect 32582 14260 32588 14272
rect 32355 14232 32588 14260
rect 32355 14229 32367 14232
rect 32309 14223 32367 14229
rect 32582 14220 32588 14232
rect 32640 14220 32646 14272
rect 33045 14263 33103 14269
rect 33045 14229 33057 14263
rect 33091 14260 33103 14263
rect 33226 14260 33232 14272
rect 33091 14232 33232 14260
rect 33091 14229 33103 14232
rect 33045 14223 33103 14229
rect 33226 14220 33232 14232
rect 33284 14220 33290 14272
rect 1104 14170 39836 14192
rect 1104 14118 4246 14170
rect 4298 14118 4310 14170
rect 4362 14118 4374 14170
rect 4426 14118 4438 14170
rect 4490 14118 34966 14170
rect 35018 14118 35030 14170
rect 35082 14118 35094 14170
rect 35146 14118 35158 14170
rect 35210 14118 39836 14170
rect 1104 14096 39836 14118
rect 9950 14016 9956 14068
rect 10008 14056 10014 14068
rect 10597 14059 10655 14065
rect 10597 14056 10609 14059
rect 10008 14028 10609 14056
rect 10008 14016 10014 14028
rect 10597 14025 10609 14028
rect 10643 14025 10655 14059
rect 10597 14019 10655 14025
rect 11238 14016 11244 14068
rect 11296 14056 11302 14068
rect 11517 14059 11575 14065
rect 11517 14056 11529 14059
rect 11296 14028 11529 14056
rect 11296 14016 11302 14028
rect 11517 14025 11529 14028
rect 11563 14025 11575 14059
rect 12066 14056 12072 14068
rect 12027 14028 12072 14056
rect 11517 14019 11575 14025
rect 12066 14016 12072 14028
rect 12124 14016 12130 14068
rect 12158 14016 12164 14068
rect 12216 14056 12222 14068
rect 24854 14056 24860 14068
rect 12216 14028 24860 14056
rect 12216 14016 12222 14028
rect 24854 14016 24860 14028
rect 24912 14016 24918 14068
rect 26142 14056 26148 14068
rect 24964 14028 26148 14056
rect 5534 13948 5540 14000
rect 5592 13988 5598 14000
rect 6181 13991 6239 13997
rect 6181 13988 6193 13991
rect 5592 13960 6193 13988
rect 5592 13948 5598 13960
rect 6181 13957 6193 13960
rect 6227 13957 6239 13991
rect 6181 13951 6239 13957
rect 2682 13861 2688 13864
rect 2677 13852 2688 13861
rect 2643 13824 2688 13852
rect 2677 13815 2688 13824
rect 2682 13812 2688 13815
rect 2740 13812 2746 13864
rect 3145 13855 3203 13861
rect 3145 13821 3157 13855
rect 3191 13852 3203 13855
rect 3421 13855 3479 13861
rect 3191 13824 3280 13852
rect 3191 13821 3203 13824
rect 3145 13815 3203 13821
rect 2501 13719 2559 13725
rect 2501 13685 2513 13719
rect 2547 13716 2559 13719
rect 3252 13716 3280 13824
rect 3421 13821 3433 13855
rect 3467 13852 3479 13855
rect 4890 13852 4896 13864
rect 3467 13824 4896 13852
rect 3467 13821 3479 13824
rect 3421 13815 3479 13821
rect 4890 13812 4896 13824
rect 4948 13812 4954 13864
rect 5994 13852 6000 13864
rect 5955 13824 6000 13852
rect 5994 13812 6000 13824
rect 6052 13812 6058 13864
rect 6196 13852 6224 13951
rect 6454 13948 6460 14000
rect 6512 13988 6518 14000
rect 6917 13991 6975 13997
rect 6917 13988 6929 13991
rect 6512 13960 6929 13988
rect 6512 13948 6518 13960
rect 6917 13957 6929 13960
rect 6963 13957 6975 13991
rect 12084 13988 12112 14016
rect 12084 13960 14964 13988
rect 6917 13951 6975 13957
rect 6730 13880 6736 13932
rect 6788 13920 6794 13932
rect 6788 13892 7604 13920
rect 6788 13880 6794 13892
rect 6825 13855 6883 13861
rect 6825 13852 6837 13855
rect 6196 13824 6837 13852
rect 6825 13821 6837 13824
rect 6871 13821 6883 13855
rect 7282 13852 7288 13864
rect 7243 13824 7288 13852
rect 6825 13815 6883 13821
rect 7282 13812 7288 13824
rect 7340 13812 7346 13864
rect 7576 13861 7604 13892
rect 7742 13880 7748 13932
rect 7800 13920 7806 13932
rect 7800 13892 9352 13920
rect 7800 13880 7806 13892
rect 7561 13855 7619 13861
rect 7561 13821 7573 13855
rect 7607 13821 7619 13855
rect 8202 13852 8208 13864
rect 8163 13824 8208 13852
rect 7561 13815 7619 13821
rect 8202 13812 8208 13824
rect 8260 13812 8266 13864
rect 8754 13852 8760 13864
rect 8715 13824 8760 13852
rect 8754 13812 8760 13824
rect 8812 13812 8818 13864
rect 9214 13852 9220 13864
rect 9175 13824 9220 13852
rect 9214 13812 9220 13824
rect 9272 13812 9278 13864
rect 9324 13852 9352 13892
rect 9398 13880 9404 13932
rect 9456 13920 9462 13932
rect 9493 13923 9551 13929
rect 9493 13920 9505 13923
rect 9456 13892 9505 13920
rect 9456 13880 9462 13892
rect 9493 13889 9505 13892
rect 9539 13889 9551 13923
rect 14001 13923 14059 13929
rect 14001 13920 14013 13923
rect 9493 13883 9551 13889
rect 9600 13892 14013 13920
rect 9600 13852 9628 13892
rect 14001 13889 14013 13892
rect 14047 13889 14059 13923
rect 14001 13883 14059 13889
rect 9324 13824 9628 13852
rect 10410 13812 10416 13864
rect 10468 13852 10474 13864
rect 11333 13855 11391 13861
rect 11333 13852 11345 13855
rect 10468 13824 11345 13852
rect 10468 13812 10474 13824
rect 11333 13821 11345 13824
rect 11379 13821 11391 13855
rect 11333 13815 11391 13821
rect 12253 13855 12311 13861
rect 12253 13821 12265 13855
rect 12299 13852 12311 13855
rect 12434 13852 12440 13864
rect 12299 13824 12440 13852
rect 12299 13821 12311 13824
rect 12253 13815 12311 13821
rect 12434 13812 12440 13824
rect 12492 13812 12498 13864
rect 12529 13855 12587 13861
rect 12529 13821 12541 13855
rect 12575 13821 12587 13855
rect 12529 13815 12587 13821
rect 12621 13855 12679 13861
rect 12621 13821 12633 13855
rect 12667 13852 12679 13855
rect 13262 13852 13268 13864
rect 12667 13824 13268 13852
rect 12667 13821 12679 13824
rect 12621 13815 12679 13821
rect 12544 13784 12572 13815
rect 13262 13812 13268 13824
rect 13320 13812 13326 13864
rect 13354 13812 13360 13864
rect 13412 13852 13418 13864
rect 13722 13852 13728 13864
rect 13412 13824 13728 13852
rect 13412 13812 13418 13824
rect 13722 13812 13728 13824
rect 13780 13812 13786 13864
rect 13906 13852 13912 13864
rect 13867 13824 13912 13852
rect 13906 13812 13912 13824
rect 13964 13812 13970 13864
rect 14936 13861 14964 13960
rect 15562 13948 15568 14000
rect 15620 13988 15626 14000
rect 16114 13988 16120 14000
rect 15620 13960 16120 13988
rect 15620 13948 15626 13960
rect 16114 13948 16120 13960
rect 16172 13948 16178 14000
rect 16574 13948 16580 14000
rect 16632 13988 16638 14000
rect 22097 13991 22155 13997
rect 16632 13960 18644 13988
rect 16632 13948 16638 13960
rect 17037 13923 17095 13929
rect 15028 13892 15976 13920
rect 14921 13855 14979 13861
rect 14921 13821 14933 13855
rect 14967 13821 14979 13855
rect 14921 13815 14979 13821
rect 12894 13784 12900 13796
rect 12544 13756 12900 13784
rect 12894 13744 12900 13756
rect 12952 13744 12958 13796
rect 15028 13784 15056 13892
rect 15194 13852 15200 13864
rect 15155 13824 15200 13852
rect 15194 13812 15200 13824
rect 15252 13812 15258 13864
rect 15948 13861 15976 13892
rect 17037 13889 17049 13923
rect 17083 13920 17095 13923
rect 18506 13920 18512 13932
rect 17083 13892 18512 13920
rect 17083 13889 17095 13892
rect 17037 13883 17095 13889
rect 18506 13880 18512 13892
rect 18564 13880 18570 13932
rect 15657 13855 15715 13861
rect 15657 13821 15669 13855
rect 15703 13821 15715 13855
rect 15657 13815 15715 13821
rect 15933 13855 15991 13861
rect 15933 13821 15945 13855
rect 15979 13821 15991 13855
rect 15933 13815 15991 13821
rect 16209 13855 16267 13861
rect 16209 13821 16221 13855
rect 16255 13852 16267 13855
rect 16669 13855 16727 13861
rect 16669 13852 16681 13855
rect 16255 13824 16681 13852
rect 16255 13821 16267 13824
rect 16209 13815 16267 13821
rect 16669 13821 16681 13824
rect 16715 13821 16727 13855
rect 16669 13815 16727 13821
rect 13280 13756 15056 13784
rect 15672 13784 15700 13815
rect 16758 13812 16764 13864
rect 16816 13852 16822 13864
rect 17221 13855 17279 13861
rect 17221 13852 17233 13855
rect 16816 13824 17233 13852
rect 16816 13812 16822 13824
rect 17221 13821 17233 13824
rect 17267 13821 17279 13855
rect 18046 13852 18052 13864
rect 18007 13824 18052 13852
rect 17221 13815 17279 13821
rect 18046 13812 18052 13824
rect 18104 13812 18110 13864
rect 18414 13852 18420 13864
rect 18375 13824 18420 13852
rect 18414 13812 18420 13824
rect 18472 13812 18478 13864
rect 18616 13861 18644 13960
rect 22097 13957 22109 13991
rect 22143 13988 22155 13991
rect 23198 13988 23204 14000
rect 22143 13960 23204 13988
rect 22143 13957 22155 13960
rect 22097 13951 22155 13957
rect 23198 13948 23204 13960
rect 23256 13948 23262 14000
rect 19150 13880 19156 13932
rect 19208 13920 19214 13932
rect 19429 13923 19487 13929
rect 19429 13920 19441 13923
rect 19208 13892 19441 13920
rect 19208 13880 19214 13892
rect 19429 13889 19441 13892
rect 19475 13889 19487 13923
rect 21082 13920 21088 13932
rect 21043 13892 21088 13920
rect 19429 13883 19487 13889
rect 21082 13880 21088 13892
rect 21140 13880 21146 13932
rect 21821 13923 21879 13929
rect 21821 13889 21833 13923
rect 21867 13920 21879 13923
rect 22186 13920 22192 13932
rect 21867 13892 22192 13920
rect 21867 13889 21879 13892
rect 21821 13883 21879 13889
rect 22186 13880 22192 13892
rect 22244 13880 22250 13932
rect 22278 13880 22284 13932
rect 22336 13920 22342 13932
rect 22833 13923 22891 13929
rect 22833 13920 22845 13923
rect 22336 13892 22845 13920
rect 22336 13880 22342 13892
rect 22833 13889 22845 13892
rect 22879 13889 22891 13923
rect 24302 13920 24308 13932
rect 24263 13892 24308 13920
rect 22833 13883 22891 13889
rect 24302 13880 24308 13892
rect 24360 13880 24366 13932
rect 24964 13929 24992 14028
rect 26142 14016 26148 14028
rect 26200 14016 26206 14068
rect 31478 14056 31484 14068
rect 26252 14028 31484 14056
rect 24949 13923 25007 13929
rect 24949 13889 24961 13923
rect 24995 13889 25007 13923
rect 24949 13883 25007 13889
rect 18601 13855 18659 13861
rect 18601 13821 18613 13855
rect 18647 13821 18659 13855
rect 18601 13815 18659 13821
rect 19705 13855 19763 13861
rect 19705 13821 19717 13855
rect 19751 13852 19763 13855
rect 19978 13852 19984 13864
rect 19751 13824 19984 13852
rect 19751 13821 19763 13824
rect 19705 13815 19763 13821
rect 19978 13812 19984 13824
rect 20036 13812 20042 13864
rect 22554 13852 22560 13864
rect 22515 13824 22560 13852
rect 22554 13812 22560 13824
rect 22612 13812 22618 13864
rect 23658 13852 23664 13864
rect 23619 13824 23664 13852
rect 23658 13812 23664 13824
rect 23716 13812 23722 13864
rect 24118 13852 24124 13864
rect 24079 13824 24124 13852
rect 24118 13812 24124 13824
rect 24176 13812 24182 13864
rect 25038 13812 25044 13864
rect 25096 13852 25102 13864
rect 26252 13861 26280 14028
rect 31478 14016 31484 14028
rect 31536 14016 31542 14068
rect 33410 14016 33416 14068
rect 33468 14056 33474 14068
rect 37734 14056 37740 14068
rect 33468 14028 37740 14056
rect 33468 14016 33474 14028
rect 37734 14016 37740 14028
rect 37792 14016 37798 14068
rect 27246 13948 27252 14000
rect 27304 13988 27310 14000
rect 34698 13988 34704 14000
rect 27304 13960 34704 13988
rect 27304 13948 27310 13960
rect 34698 13948 34704 13960
rect 34756 13948 34762 14000
rect 27614 13920 27620 13932
rect 26620 13892 27620 13920
rect 26237 13855 26295 13861
rect 25096 13824 25141 13852
rect 25096 13812 25102 13824
rect 26237 13821 26249 13855
rect 26283 13821 26295 13855
rect 26237 13815 26295 13821
rect 26329 13855 26387 13861
rect 26329 13821 26341 13855
rect 26375 13852 26387 13855
rect 26620 13852 26648 13892
rect 27614 13880 27620 13892
rect 27672 13880 27678 13932
rect 28074 13920 28080 13932
rect 28035 13892 28080 13920
rect 28074 13880 28080 13892
rect 28132 13880 28138 13932
rect 28534 13880 28540 13932
rect 28592 13920 28598 13932
rect 29273 13923 29331 13929
rect 29273 13920 29285 13923
rect 28592 13892 29285 13920
rect 28592 13880 28598 13892
rect 29273 13889 29285 13892
rect 29319 13889 29331 13923
rect 30006 13920 30012 13932
rect 29967 13892 30012 13920
rect 29273 13883 29331 13889
rect 30006 13880 30012 13892
rect 30064 13880 30070 13932
rect 30834 13920 30840 13932
rect 30795 13892 30840 13920
rect 30834 13880 30840 13892
rect 30892 13880 30898 13932
rect 34146 13920 34152 13932
rect 34107 13892 34152 13920
rect 34146 13880 34152 13892
rect 34204 13880 34210 13932
rect 35526 13920 35532 13932
rect 35487 13892 35532 13920
rect 35526 13880 35532 13892
rect 35584 13880 35590 13932
rect 35802 13920 35808 13932
rect 35763 13892 35808 13920
rect 35802 13880 35808 13892
rect 35860 13880 35866 13932
rect 38289 13923 38347 13929
rect 38289 13889 38301 13923
rect 38335 13920 38347 13923
rect 38562 13920 38568 13932
rect 38335 13892 38568 13920
rect 38335 13889 38347 13892
rect 38289 13883 38347 13889
rect 38562 13880 38568 13892
rect 38620 13880 38626 13932
rect 26375 13824 26648 13852
rect 26697 13855 26755 13861
rect 26375 13821 26387 13824
rect 26329 13815 26387 13821
rect 26697 13821 26709 13855
rect 26743 13852 26755 13855
rect 26878 13852 26884 13864
rect 26743 13824 26884 13852
rect 26743 13821 26755 13824
rect 26697 13815 26755 13821
rect 26878 13812 26884 13824
rect 26936 13812 26942 13864
rect 27154 13852 27160 13864
rect 27115 13824 27160 13852
rect 27154 13812 27160 13824
rect 27212 13852 27218 13864
rect 27430 13852 27436 13864
rect 27212 13824 27436 13852
rect 27212 13812 27218 13824
rect 27430 13812 27436 13824
rect 27488 13812 27494 13864
rect 27709 13855 27767 13861
rect 27709 13821 27721 13855
rect 27755 13852 27767 13855
rect 27890 13852 27896 13864
rect 27755 13824 27896 13852
rect 27755 13821 27767 13824
rect 27709 13815 27767 13821
rect 27890 13812 27896 13824
rect 27948 13812 27954 13864
rect 27985 13855 28043 13861
rect 27985 13821 27997 13855
rect 28031 13852 28043 13855
rect 28718 13852 28724 13864
rect 28031 13824 28724 13852
rect 28031 13821 28043 13824
rect 27985 13815 28043 13821
rect 28552 13796 28580 13824
rect 28718 13812 28724 13824
rect 28776 13812 28782 13864
rect 28902 13812 28908 13864
rect 28960 13812 28966 13864
rect 29086 13812 29092 13864
rect 29144 13852 29150 13864
rect 29362 13852 29368 13864
rect 29144 13824 29368 13852
rect 29144 13812 29150 13824
rect 29362 13812 29368 13824
rect 29420 13852 29426 13864
rect 29457 13855 29515 13861
rect 29457 13852 29469 13855
rect 29420 13824 29469 13852
rect 29420 13812 29426 13824
rect 29457 13821 29469 13824
rect 29503 13821 29515 13855
rect 31386 13852 31392 13864
rect 31347 13824 31392 13852
rect 29457 13815 29515 13821
rect 31386 13812 31392 13824
rect 31444 13812 31450 13864
rect 31754 13812 31760 13864
rect 31812 13852 31818 13864
rect 32125 13855 32183 13861
rect 31812 13824 31857 13852
rect 31812 13812 31818 13824
rect 32125 13821 32137 13855
rect 32171 13821 32183 13855
rect 32490 13852 32496 13864
rect 32451 13824 32496 13852
rect 32125 13815 32183 13821
rect 16942 13784 16948 13796
rect 15672 13756 16948 13784
rect 4062 13716 4068 13728
rect 2547 13688 4068 13716
rect 2547 13685 2559 13688
rect 2501 13679 2559 13685
rect 4062 13676 4068 13688
rect 4120 13676 4126 13728
rect 4338 13676 4344 13728
rect 4396 13716 4402 13728
rect 13280 13725 13308 13756
rect 16684 13728 16712 13756
rect 16942 13744 16948 13756
rect 17000 13744 17006 13796
rect 25501 13787 25559 13793
rect 25501 13753 25513 13787
rect 25547 13784 25559 13787
rect 27246 13784 27252 13796
rect 25547 13756 27252 13784
rect 25547 13753 25559 13756
rect 25501 13747 25559 13753
rect 27246 13744 27252 13756
rect 27304 13744 27310 13796
rect 28534 13744 28540 13796
rect 28592 13744 28598 13796
rect 28920 13784 28948 13812
rect 29641 13787 29699 13793
rect 29641 13784 29653 13787
rect 28736 13756 28948 13784
rect 29380 13756 29653 13784
rect 28736 13728 28764 13756
rect 4525 13719 4583 13725
rect 4525 13716 4537 13719
rect 4396 13688 4537 13716
rect 4396 13676 4402 13688
rect 4525 13685 4537 13688
rect 4571 13685 4583 13719
rect 4525 13679 4583 13685
rect 13265 13719 13323 13725
rect 13265 13685 13277 13719
rect 13311 13685 13323 13719
rect 13265 13679 13323 13685
rect 14737 13719 14795 13725
rect 14737 13685 14749 13719
rect 14783 13716 14795 13719
rect 15286 13716 15292 13728
rect 14783 13688 15292 13716
rect 14783 13685 14795 13688
rect 14737 13679 14795 13685
rect 15286 13676 15292 13688
rect 15344 13676 15350 13728
rect 16666 13676 16672 13728
rect 16724 13676 16730 13728
rect 28718 13676 28724 13728
rect 28776 13676 28782 13728
rect 28902 13676 28908 13728
rect 28960 13716 28966 13728
rect 29380 13716 29408 13756
rect 29641 13753 29653 13756
rect 29687 13753 29699 13787
rect 31202 13784 31208 13796
rect 31163 13756 31208 13784
rect 29641 13747 29699 13753
rect 31202 13744 31208 13756
rect 31260 13744 31266 13796
rect 31662 13744 31668 13796
rect 31720 13784 31726 13796
rect 32140 13784 32168 13815
rect 32490 13812 32496 13824
rect 32548 13812 32554 13864
rect 33226 13852 33232 13864
rect 33187 13824 33232 13852
rect 33226 13812 33232 13824
rect 33284 13812 33290 13864
rect 33318 13812 33324 13864
rect 33376 13852 33382 13864
rect 33597 13855 33655 13861
rect 33597 13852 33609 13855
rect 33376 13824 33609 13852
rect 33376 13812 33382 13824
rect 33597 13821 33609 13824
rect 33643 13821 33655 13855
rect 33597 13815 33655 13821
rect 34057 13855 34115 13861
rect 34057 13821 34069 13855
rect 34103 13852 34115 13855
rect 34330 13852 34336 13864
rect 34103 13824 34336 13852
rect 34103 13821 34115 13824
rect 34057 13815 34115 13821
rect 34330 13812 34336 13824
rect 34388 13812 34394 13864
rect 38102 13852 38108 13864
rect 38063 13824 38108 13852
rect 38102 13812 38108 13824
rect 38160 13812 38166 13864
rect 38470 13852 38476 13864
rect 38431 13824 38476 13852
rect 38470 13812 38476 13824
rect 38528 13812 38534 13864
rect 31720 13756 32168 13784
rect 31720 13744 31726 13756
rect 28960 13688 29408 13716
rect 28960 13676 28966 13688
rect 29546 13676 29552 13728
rect 29604 13716 29610 13728
rect 29604 13688 29649 13716
rect 29604 13676 29610 13688
rect 36538 13676 36544 13728
rect 36596 13716 36602 13728
rect 36909 13719 36967 13725
rect 36909 13716 36921 13719
rect 36596 13688 36921 13716
rect 36596 13676 36602 13688
rect 36909 13685 36921 13688
rect 36955 13685 36967 13719
rect 36909 13679 36967 13685
rect 1104 13626 39836 13648
rect 1104 13574 19606 13626
rect 19658 13574 19670 13626
rect 19722 13574 19734 13626
rect 19786 13574 19798 13626
rect 19850 13574 39836 13626
rect 1104 13552 39836 13574
rect 5626 13512 5632 13524
rect 5587 13484 5632 13512
rect 5626 13472 5632 13484
rect 5684 13472 5690 13524
rect 6365 13515 6423 13521
rect 6365 13481 6377 13515
rect 6411 13512 6423 13515
rect 7282 13512 7288 13524
rect 6411 13484 7288 13512
rect 6411 13481 6423 13484
rect 6365 13475 6423 13481
rect 7282 13472 7288 13484
rect 7340 13472 7346 13524
rect 8110 13472 8116 13524
rect 8168 13512 8174 13524
rect 9033 13515 9091 13521
rect 9033 13512 9045 13515
rect 8168 13484 9045 13512
rect 8168 13472 8174 13484
rect 9033 13481 9045 13484
rect 9079 13481 9091 13515
rect 9674 13512 9680 13524
rect 9033 13475 9091 13481
rect 9140 13484 9680 13512
rect 7742 13444 7748 13456
rect 6288 13416 7748 13444
rect 4062 13376 4068 13388
rect 4023 13348 4068 13376
rect 4062 13336 4068 13348
rect 4120 13336 4126 13388
rect 4338 13376 4344 13388
rect 4299 13348 4344 13376
rect 4338 13336 4344 13348
rect 4396 13336 4402 13388
rect 6288 13385 6316 13416
rect 7742 13404 7748 13416
rect 7800 13404 7806 13456
rect 6273 13379 6331 13385
rect 6273 13345 6285 13379
rect 6319 13345 6331 13379
rect 6273 13339 6331 13345
rect 7469 13379 7527 13385
rect 7469 13345 7481 13379
rect 7515 13345 7527 13379
rect 7469 13339 7527 13345
rect 7837 13379 7895 13385
rect 7837 13345 7849 13379
rect 7883 13376 7895 13379
rect 8294 13376 8300 13388
rect 7883 13348 8300 13376
rect 7883 13345 7895 13348
rect 7837 13339 7895 13345
rect 1394 13308 1400 13320
rect 1355 13280 1400 13308
rect 1394 13268 1400 13280
rect 1452 13268 1458 13320
rect 1670 13308 1676 13320
rect 1631 13280 1676 13308
rect 1670 13268 1676 13280
rect 1728 13268 1734 13320
rect 7098 13308 7104 13320
rect 7059 13280 7104 13308
rect 7098 13268 7104 13280
rect 7156 13268 7162 13320
rect 7374 13268 7380 13320
rect 7432 13308 7438 13320
rect 7484 13308 7512 13339
rect 8294 13336 8300 13348
rect 8352 13336 8358 13388
rect 8849 13379 8907 13385
rect 8849 13345 8861 13379
rect 8895 13376 8907 13379
rect 9140 13376 9168 13484
rect 9674 13472 9680 13484
rect 9732 13512 9738 13524
rect 10410 13512 10416 13524
rect 9732 13484 10416 13512
rect 9732 13472 9738 13484
rect 10410 13472 10416 13484
rect 10468 13472 10474 13524
rect 16942 13472 16948 13524
rect 17000 13512 17006 13524
rect 17218 13512 17224 13524
rect 17000 13484 17224 13512
rect 17000 13472 17006 13484
rect 17218 13472 17224 13484
rect 17276 13472 17282 13524
rect 20622 13472 20628 13524
rect 20680 13512 20686 13524
rect 20993 13515 21051 13521
rect 20993 13512 21005 13515
rect 20680 13484 21005 13512
rect 20680 13472 20686 13484
rect 20993 13481 21005 13484
rect 21039 13481 21051 13515
rect 20993 13475 21051 13481
rect 22186 13472 22192 13524
rect 22244 13512 22250 13524
rect 22244 13484 25360 13512
rect 22244 13472 22250 13484
rect 23934 13444 23940 13456
rect 10428 13416 23244 13444
rect 10134 13376 10140 13388
rect 8895 13348 9168 13376
rect 10095 13348 10140 13376
rect 8895 13345 8907 13348
rect 8849 13339 8907 13345
rect 10134 13336 10140 13348
rect 10192 13336 10198 13388
rect 10428 13385 10456 13416
rect 10413 13379 10471 13385
rect 10413 13345 10425 13379
rect 10459 13345 10471 13379
rect 10778 13376 10784 13388
rect 10739 13348 10784 13376
rect 10413 13339 10471 13345
rect 10778 13336 10784 13348
rect 10836 13336 10842 13388
rect 11054 13336 11060 13388
rect 11112 13376 11118 13388
rect 11425 13379 11483 13385
rect 11425 13376 11437 13379
rect 11112 13348 11437 13376
rect 11112 13336 11118 13348
rect 11425 13345 11437 13348
rect 11471 13345 11483 13379
rect 11974 13376 11980 13388
rect 11935 13348 11980 13376
rect 11425 13339 11483 13345
rect 11974 13336 11980 13348
rect 12032 13336 12038 13388
rect 12437 13379 12495 13385
rect 12437 13345 12449 13379
rect 12483 13376 12495 13379
rect 13357 13379 13415 13385
rect 12483 13348 12848 13376
rect 12483 13345 12495 13348
rect 12437 13339 12495 13345
rect 8110 13308 8116 13320
rect 7432 13280 8116 13308
rect 7432 13268 7438 13280
rect 8110 13268 8116 13280
rect 8168 13268 8174 13320
rect 12621 13311 12679 13317
rect 12621 13277 12633 13311
rect 12667 13277 12679 13311
rect 12820 13308 12848 13348
rect 13357 13345 13369 13379
rect 13403 13345 13415 13379
rect 13722 13376 13728 13388
rect 13683 13348 13728 13376
rect 13357 13339 13415 13345
rect 13372 13308 13400 13339
rect 13722 13336 13728 13348
rect 13780 13336 13786 13388
rect 14461 13379 14519 13385
rect 14461 13345 14473 13379
rect 14507 13345 14519 13379
rect 15746 13376 15752 13388
rect 15707 13348 15752 13376
rect 14461 13339 14519 13345
rect 13814 13308 13820 13320
rect 12820 13280 13216 13308
rect 13372 13280 13820 13308
rect 12621 13271 12679 13277
rect 7282 13200 7288 13252
rect 7340 13240 7346 13252
rect 7745 13243 7803 13249
rect 7745 13240 7757 13243
rect 7340 13212 7757 13240
rect 7340 13200 7346 13212
rect 7745 13209 7757 13212
rect 7791 13209 7803 13243
rect 7745 13203 7803 13209
rect 2961 13175 3019 13181
rect 2961 13141 2973 13175
rect 3007 13172 3019 13175
rect 3786 13172 3792 13184
rect 3007 13144 3792 13172
rect 3007 13141 3019 13144
rect 2961 13135 3019 13141
rect 3786 13132 3792 13144
rect 3844 13132 3850 13184
rect 12636 13172 12664 13271
rect 13188 13249 13216 13280
rect 13814 13268 13820 13280
rect 13872 13268 13878 13320
rect 13173 13243 13231 13249
rect 13173 13209 13185 13243
rect 13219 13209 13231 13243
rect 13173 13203 13231 13209
rect 13262 13200 13268 13252
rect 13320 13240 13326 13252
rect 13998 13240 14004 13252
rect 13320 13212 14004 13240
rect 13320 13200 13326 13212
rect 13998 13200 14004 13212
rect 14056 13240 14062 13252
rect 14476 13240 14504 13339
rect 15746 13336 15752 13348
rect 15804 13336 15810 13388
rect 16114 13376 16120 13388
rect 16075 13348 16120 13376
rect 16114 13336 16120 13348
rect 16172 13336 16178 13388
rect 16393 13379 16451 13385
rect 16393 13345 16405 13379
rect 16439 13376 16451 13379
rect 16758 13376 16764 13388
rect 16439 13348 16764 13376
rect 16439 13345 16451 13348
rect 16393 13339 16451 13345
rect 16758 13336 16764 13348
rect 16816 13336 16822 13388
rect 16853 13379 16911 13385
rect 16853 13345 16865 13379
rect 16899 13345 16911 13379
rect 16853 13339 16911 13345
rect 15473 13311 15531 13317
rect 15473 13277 15485 13311
rect 15519 13308 15531 13311
rect 15930 13308 15936 13320
rect 15519 13280 15936 13308
rect 15519 13277 15531 13280
rect 15473 13271 15531 13277
rect 15930 13268 15936 13280
rect 15988 13268 15994 13320
rect 16868 13240 16896 13339
rect 18506 13336 18512 13388
rect 18564 13376 18570 13388
rect 18601 13379 18659 13385
rect 18601 13376 18613 13379
rect 18564 13348 18613 13376
rect 18564 13336 18570 13348
rect 18601 13345 18613 13348
rect 18647 13345 18659 13379
rect 19334 13376 19340 13388
rect 18601 13339 18659 13345
rect 18984 13348 19340 13376
rect 17865 13311 17923 13317
rect 17865 13277 17877 13311
rect 17911 13308 17923 13311
rect 18230 13308 18236 13320
rect 17911 13280 18236 13308
rect 17911 13277 17923 13280
rect 17865 13271 17923 13277
rect 18230 13268 18236 13280
rect 18288 13268 18294 13320
rect 18325 13243 18383 13249
rect 14056 13212 16896 13240
rect 16960 13212 17264 13240
rect 14056 13200 14062 13212
rect 13538 13172 13544 13184
rect 12636 13144 13544 13172
rect 13538 13132 13544 13144
rect 13596 13132 13602 13184
rect 14645 13175 14703 13181
rect 14645 13141 14657 13175
rect 14691 13172 14703 13175
rect 15102 13172 15108 13184
rect 14691 13144 15108 13172
rect 14691 13141 14703 13144
rect 14645 13135 14703 13141
rect 15102 13132 15108 13144
rect 15160 13172 15166 13184
rect 15746 13172 15752 13184
rect 15160 13144 15752 13172
rect 15160 13132 15166 13144
rect 15746 13132 15752 13144
rect 15804 13172 15810 13184
rect 16960 13172 16988 13212
rect 15804 13144 16988 13172
rect 17037 13175 17095 13181
rect 15804 13132 15810 13144
rect 17037 13141 17049 13175
rect 17083 13172 17095 13175
rect 17126 13172 17132 13184
rect 17083 13144 17132 13172
rect 17083 13141 17095 13144
rect 17037 13135 17095 13141
rect 17126 13132 17132 13144
rect 17184 13132 17190 13184
rect 17236 13172 17264 13212
rect 18325 13209 18337 13243
rect 18371 13240 18383 13243
rect 18984 13240 19012 13348
rect 19334 13336 19340 13348
rect 19392 13336 19398 13388
rect 19886 13376 19892 13388
rect 19847 13348 19892 13376
rect 19886 13336 19892 13348
rect 19944 13336 19950 13388
rect 20346 13376 20352 13388
rect 20307 13348 20352 13376
rect 20346 13336 20352 13348
rect 20404 13336 20410 13388
rect 20438 13336 20444 13388
rect 20496 13376 20502 13388
rect 20622 13376 20628 13388
rect 20496 13348 20628 13376
rect 20496 13336 20502 13348
rect 20622 13336 20628 13348
rect 20680 13336 20686 13388
rect 21085 13379 21143 13385
rect 21085 13345 21097 13379
rect 21131 13376 21143 13379
rect 21174 13376 21180 13388
rect 21131 13348 21180 13376
rect 21131 13345 21143 13348
rect 21085 13339 21143 13345
rect 21174 13336 21180 13348
rect 21232 13336 21238 13388
rect 21450 13376 21456 13388
rect 21411 13348 21456 13376
rect 21450 13336 21456 13348
rect 21508 13336 21514 13388
rect 23216 13385 23244 13416
rect 23308 13416 23940 13444
rect 23201 13379 23259 13385
rect 23201 13345 23213 13379
rect 23247 13345 23259 13379
rect 23201 13339 23259 13345
rect 19061 13311 19119 13317
rect 19061 13277 19073 13311
rect 19107 13277 19119 13311
rect 19061 13271 19119 13277
rect 19981 13311 20039 13317
rect 19981 13277 19993 13311
rect 20027 13308 20039 13311
rect 21729 13311 21787 13317
rect 21729 13308 21741 13311
rect 20027 13280 21741 13308
rect 20027 13277 20039 13280
rect 19981 13271 20039 13277
rect 21729 13277 21741 13280
rect 21775 13277 21787 13311
rect 21729 13271 21787 13277
rect 22465 13311 22523 13317
rect 22465 13277 22477 13311
rect 22511 13308 22523 13311
rect 22646 13308 22652 13320
rect 22511 13280 22652 13308
rect 22511 13277 22523 13280
rect 22465 13271 22523 13277
rect 19076 13240 19104 13271
rect 22646 13268 22652 13280
rect 22704 13268 22710 13320
rect 23308 13308 23336 13416
rect 23934 13404 23940 13416
rect 23992 13404 23998 13456
rect 25332 13453 25360 13484
rect 26418 13472 26424 13524
rect 26476 13512 26482 13524
rect 29362 13512 29368 13524
rect 26476 13484 29368 13512
rect 26476 13472 26482 13484
rect 29362 13472 29368 13484
rect 29420 13472 29426 13524
rect 32306 13512 32312 13524
rect 29840 13484 32168 13512
rect 32267 13484 32312 13512
rect 25317 13447 25375 13453
rect 25317 13413 25329 13447
rect 25363 13413 25375 13447
rect 25317 13407 25375 13413
rect 26970 13404 26976 13456
rect 27028 13404 27034 13456
rect 27338 13404 27344 13456
rect 27396 13444 27402 13456
rect 29457 13447 29515 13453
rect 29457 13444 29469 13447
rect 27396 13416 27844 13444
rect 27396 13404 27402 13416
rect 23477 13379 23535 13385
rect 23477 13345 23489 13379
rect 23523 13345 23535 13379
rect 23477 13339 23535 13345
rect 22940 13280 23336 13308
rect 19150 13240 19156 13252
rect 18371 13212 19012 13240
rect 19063 13212 19156 13240
rect 18371 13209 18383 13212
rect 18325 13203 18383 13209
rect 19150 13200 19156 13212
rect 19208 13240 19214 13252
rect 22278 13240 22284 13252
rect 19208 13212 22284 13240
rect 19208 13200 19214 13212
rect 22278 13200 22284 13212
rect 22336 13200 22342 13252
rect 22940 13249 22968 13280
rect 22925 13243 22983 13249
rect 22925 13209 22937 13243
rect 22971 13209 22983 13243
rect 22925 13203 22983 13209
rect 21910 13172 21916 13184
rect 17236 13144 21916 13172
rect 21910 13132 21916 13144
rect 21968 13132 21974 13184
rect 22296 13172 22324 13200
rect 23492 13172 23520 13339
rect 23566 13336 23572 13388
rect 23624 13376 23630 13388
rect 24581 13379 24639 13385
rect 24581 13376 24593 13379
rect 23624 13348 24593 13376
rect 23624 13336 23630 13348
rect 24581 13345 24593 13348
rect 24627 13345 24639 13379
rect 24581 13339 24639 13345
rect 25041 13379 25099 13385
rect 25041 13345 25053 13379
rect 25087 13345 25099 13379
rect 26988 13376 27016 13404
rect 27433 13379 27491 13385
rect 27433 13376 27445 13379
rect 26988 13348 27445 13376
rect 25041 13339 25099 13345
rect 27433 13345 27445 13348
rect 27479 13345 27491 13379
rect 27433 13339 27491 13345
rect 24210 13268 24216 13320
rect 24268 13308 24274 13320
rect 24305 13311 24363 13317
rect 24305 13308 24317 13311
rect 24268 13280 24317 13308
rect 24268 13268 24274 13280
rect 24305 13277 24317 13280
rect 24351 13277 24363 13311
rect 24305 13271 24363 13277
rect 23658 13200 23664 13252
rect 23716 13240 23722 13252
rect 25056 13240 25084 13339
rect 27522 13336 27528 13388
rect 27580 13376 27586 13388
rect 27816 13385 27844 13416
rect 28368 13416 29469 13444
rect 27617 13379 27675 13385
rect 27617 13376 27629 13379
rect 27580 13348 27629 13376
rect 27580 13336 27586 13348
rect 27617 13345 27629 13348
rect 27663 13345 27675 13379
rect 27617 13339 27675 13345
rect 27801 13379 27859 13385
rect 27801 13345 27813 13379
rect 27847 13345 27859 13379
rect 28074 13376 28080 13388
rect 28035 13348 28080 13376
rect 27801 13339 27859 13345
rect 28074 13336 28080 13348
rect 28132 13336 28138 13388
rect 28368 13385 28396 13416
rect 29457 13413 29469 13416
rect 29503 13444 29515 13447
rect 29546 13444 29552 13456
rect 29503 13416 29552 13444
rect 29503 13413 29515 13416
rect 29457 13407 29515 13413
rect 29546 13404 29552 13416
rect 29604 13404 29610 13456
rect 29840 13453 29868 13484
rect 29825 13447 29883 13453
rect 29825 13413 29837 13447
rect 29871 13413 29883 13447
rect 29825 13407 29883 13413
rect 28353 13379 28411 13385
rect 28353 13345 28365 13379
rect 28399 13345 28411 13379
rect 28353 13339 28411 13345
rect 28994 13336 29000 13388
rect 29052 13376 29058 13388
rect 29273 13379 29331 13385
rect 29273 13376 29285 13379
rect 29052 13348 29285 13376
rect 29052 13336 29058 13348
rect 29273 13345 29285 13348
rect 29319 13376 29331 13379
rect 30282 13376 30288 13388
rect 29319 13348 30288 13376
rect 29319 13345 29331 13348
rect 29273 13339 29331 13345
rect 30282 13336 30288 13348
rect 30340 13336 30346 13388
rect 30834 13376 30840 13388
rect 30795 13348 30840 13376
rect 30834 13336 30840 13348
rect 30892 13336 30898 13388
rect 31202 13336 31208 13388
rect 31260 13376 31266 13388
rect 32140 13385 32168 13484
rect 32306 13472 32312 13484
rect 32364 13472 32370 13524
rect 33229 13515 33287 13521
rect 33229 13481 33241 13515
rect 33275 13512 33287 13515
rect 33870 13512 33876 13524
rect 33275 13484 33876 13512
rect 33275 13481 33287 13484
rect 33229 13475 33287 13481
rect 33870 13472 33876 13484
rect 33928 13472 33934 13524
rect 33962 13472 33968 13524
rect 34020 13512 34026 13524
rect 34020 13484 34836 13512
rect 34020 13472 34026 13484
rect 34054 13444 34060 13456
rect 33336 13416 34060 13444
rect 33336 13385 33364 13416
rect 34054 13404 34060 13416
rect 34112 13404 34118 13456
rect 31297 13379 31355 13385
rect 31297 13376 31309 13379
rect 31260 13348 31309 13376
rect 31260 13336 31266 13348
rect 31297 13345 31309 13348
rect 31343 13345 31355 13379
rect 31297 13339 31355 13345
rect 32125 13379 32183 13385
rect 32125 13345 32137 13379
rect 32171 13345 32183 13379
rect 32125 13339 32183 13345
rect 33321 13379 33379 13385
rect 33321 13345 33333 13379
rect 33367 13345 33379 13379
rect 33686 13376 33692 13388
rect 33647 13348 33692 13376
rect 33321 13339 33379 13345
rect 33686 13336 33692 13348
rect 33744 13336 33750 13388
rect 34146 13376 34152 13388
rect 34107 13348 34152 13376
rect 34146 13336 34152 13348
rect 34204 13336 34210 13388
rect 34808 13385 34836 13484
rect 37185 13447 37243 13453
rect 37185 13413 37197 13447
rect 37231 13444 37243 13447
rect 37826 13444 37832 13456
rect 37231 13416 37832 13444
rect 37231 13413 37243 13416
rect 37185 13407 37243 13413
rect 37826 13404 37832 13416
rect 37884 13404 37890 13456
rect 34793 13379 34851 13385
rect 34793 13345 34805 13379
rect 34839 13345 34851 13379
rect 36078 13376 36084 13388
rect 36039 13348 36084 13376
rect 34793 13339 34851 13345
rect 36078 13336 36084 13348
rect 36136 13336 36142 13388
rect 36538 13376 36544 13388
rect 36499 13348 36544 13376
rect 36538 13336 36544 13348
rect 36596 13336 36602 13388
rect 36722 13376 36728 13388
rect 36683 13348 36728 13376
rect 36722 13336 36728 13348
rect 36780 13336 36786 13388
rect 37734 13376 37740 13388
rect 37695 13348 37740 13376
rect 37734 13336 37740 13348
rect 37792 13336 37798 13388
rect 38194 13336 38200 13388
rect 38252 13376 38258 13388
rect 38289 13379 38347 13385
rect 38289 13376 38301 13379
rect 38252 13348 38301 13376
rect 38252 13336 38258 13348
rect 38289 13345 38301 13348
rect 38335 13345 38347 13379
rect 38289 13339 38347 13345
rect 26973 13311 27031 13317
rect 26973 13277 26985 13311
rect 27019 13277 27031 13311
rect 26973 13271 27031 13277
rect 23716 13212 25084 13240
rect 26988 13240 27016 13271
rect 27706 13268 27712 13320
rect 27764 13308 27770 13320
rect 28902 13308 28908 13320
rect 27764 13280 28908 13308
rect 27764 13268 27770 13280
rect 28902 13268 28908 13280
rect 28960 13308 28966 13320
rect 29089 13311 29147 13317
rect 29089 13308 29101 13311
rect 28960 13280 29101 13308
rect 28960 13268 28966 13280
rect 29089 13277 29101 13280
rect 29135 13277 29147 13311
rect 30650 13308 30656 13320
rect 30563 13280 30656 13308
rect 29089 13271 29147 13277
rect 30650 13268 30656 13280
rect 30708 13308 30714 13320
rect 31386 13308 31392 13320
rect 30708 13280 31392 13308
rect 30708 13268 30714 13280
rect 31386 13268 31392 13280
rect 31444 13268 31450 13320
rect 32030 13268 32036 13320
rect 32088 13308 32094 13320
rect 32306 13308 32312 13320
rect 32088 13280 32312 13308
rect 32088 13268 32094 13280
rect 32306 13268 32312 13280
rect 32364 13268 32370 13320
rect 38562 13308 38568 13320
rect 38523 13280 38568 13308
rect 38562 13268 38568 13280
rect 38620 13268 38626 13320
rect 29730 13240 29736 13252
rect 26988 13212 29736 13240
rect 23716 13200 23722 13212
rect 29730 13200 29736 13212
rect 29788 13200 29794 13252
rect 31294 13240 31300 13252
rect 31255 13212 31300 13240
rect 31294 13200 31300 13212
rect 31352 13200 31358 13252
rect 37734 13200 37740 13252
rect 37792 13240 37798 13252
rect 37829 13243 37887 13249
rect 37829 13240 37841 13243
rect 37792 13212 37841 13240
rect 37792 13200 37798 13212
rect 37829 13209 37841 13212
rect 37875 13209 37887 13243
rect 37829 13203 37887 13209
rect 22296 13144 23520 13172
rect 34977 13175 35035 13181
rect 34977 13141 34989 13175
rect 35023 13172 35035 13175
rect 35802 13172 35808 13184
rect 35023 13144 35808 13172
rect 35023 13141 35035 13144
rect 34977 13135 35035 13141
rect 35802 13132 35808 13144
rect 35860 13132 35866 13184
rect 1104 13082 39836 13104
rect 1104 13030 4246 13082
rect 4298 13030 4310 13082
rect 4362 13030 4374 13082
rect 4426 13030 4438 13082
rect 4490 13030 34966 13082
rect 35018 13030 35030 13082
rect 35082 13030 35094 13082
rect 35146 13030 35158 13082
rect 35210 13030 39836 13082
rect 1104 13008 39836 13030
rect 1670 12928 1676 12980
rect 1728 12968 1734 12980
rect 2777 12971 2835 12977
rect 2777 12968 2789 12971
rect 1728 12940 2789 12968
rect 1728 12928 1734 12940
rect 2777 12937 2789 12940
rect 2823 12937 2835 12971
rect 4890 12968 4896 12980
rect 4851 12940 4896 12968
rect 2777 12931 2835 12937
rect 4890 12928 4896 12940
rect 4948 12928 4954 12980
rect 6178 12968 6184 12980
rect 6139 12940 6184 12968
rect 6178 12928 6184 12940
rect 6236 12928 6242 12980
rect 14093 12971 14151 12977
rect 14093 12937 14105 12971
rect 14139 12968 14151 12971
rect 16758 12968 16764 12980
rect 14139 12940 16764 12968
rect 14139 12937 14151 12940
rect 14093 12931 14151 12937
rect 16758 12928 16764 12940
rect 16816 12928 16822 12980
rect 20990 12968 20996 12980
rect 20364 12940 20996 12968
rect 11054 12860 11060 12912
rect 11112 12900 11118 12912
rect 12529 12903 12587 12909
rect 12529 12900 12541 12903
rect 11112 12872 12541 12900
rect 11112 12860 11118 12872
rect 12529 12869 12541 12872
rect 12575 12869 12587 12903
rect 12529 12863 12587 12869
rect 13722 12860 13728 12912
rect 13780 12900 13786 12912
rect 18509 12903 18567 12909
rect 13780 12872 16988 12900
rect 13780 12860 13786 12872
rect 1394 12832 1400 12844
rect 1307 12804 1400 12832
rect 1394 12792 1400 12804
rect 1452 12832 1458 12844
rect 1854 12832 1860 12844
rect 1452 12804 1860 12832
rect 1452 12792 1458 12804
rect 1854 12792 1860 12804
rect 1912 12832 1918 12844
rect 3786 12832 3792 12844
rect 1912 12804 3556 12832
rect 3747 12804 3792 12832
rect 1912 12792 1918 12804
rect 1673 12767 1731 12773
rect 1673 12733 1685 12767
rect 1719 12764 1731 12767
rect 3234 12764 3240 12776
rect 1719 12736 3240 12764
rect 1719 12733 1731 12736
rect 1673 12727 1731 12733
rect 3234 12724 3240 12736
rect 3292 12724 3298 12776
rect 3528 12773 3556 12804
rect 3786 12792 3792 12804
rect 3844 12792 3850 12844
rect 6914 12792 6920 12844
rect 6972 12832 6978 12844
rect 7009 12835 7067 12841
rect 7009 12832 7021 12835
rect 6972 12804 7021 12832
rect 6972 12792 6978 12804
rect 7009 12801 7021 12804
rect 7055 12801 7067 12835
rect 7282 12832 7288 12844
rect 7243 12804 7288 12832
rect 7009 12795 7067 12801
rect 7282 12792 7288 12804
rect 7340 12792 7346 12844
rect 9493 12835 9551 12841
rect 9493 12801 9505 12835
rect 9539 12832 9551 12835
rect 9858 12832 9864 12844
rect 9539 12804 9864 12832
rect 9539 12801 9551 12804
rect 9493 12795 9551 12801
rect 9858 12792 9864 12804
rect 9916 12792 9922 12844
rect 13814 12832 13820 12844
rect 10888 12804 13820 12832
rect 10888 12776 10916 12804
rect 13814 12792 13820 12804
rect 13872 12792 13878 12844
rect 14829 12835 14887 12841
rect 14829 12801 14841 12835
rect 14875 12832 14887 12835
rect 15749 12835 15807 12841
rect 14875 12804 15700 12832
rect 14875 12801 14887 12804
rect 14829 12795 14887 12801
rect 3513 12767 3571 12773
rect 3513 12733 3525 12767
rect 3559 12764 3571 12767
rect 4062 12764 4068 12776
rect 3559 12736 4068 12764
rect 3559 12733 3571 12736
rect 3513 12727 3571 12733
rect 4062 12724 4068 12736
rect 4120 12724 4126 12776
rect 6089 12767 6147 12773
rect 6089 12733 6101 12767
rect 6135 12733 6147 12767
rect 9122 12764 9128 12776
rect 9083 12736 9128 12764
rect 6089 12727 6147 12733
rect 6104 12628 6132 12727
rect 9122 12724 9128 12736
rect 9180 12724 9186 12776
rect 9677 12767 9735 12773
rect 9677 12733 9689 12767
rect 9723 12733 9735 12767
rect 9677 12727 9735 12733
rect 10321 12767 10379 12773
rect 10321 12733 10333 12767
rect 10367 12733 10379 12767
rect 10686 12764 10692 12776
rect 10647 12736 10692 12764
rect 10321 12727 10379 12733
rect 8018 12656 8024 12708
rect 8076 12696 8082 12708
rect 8665 12699 8723 12705
rect 8665 12696 8677 12699
rect 8076 12668 8677 12696
rect 8076 12656 8082 12668
rect 8665 12665 8677 12668
rect 8711 12696 8723 12699
rect 9692 12696 9720 12727
rect 8711 12668 9720 12696
rect 8711 12665 8723 12668
rect 8665 12659 8723 12665
rect 8478 12628 8484 12640
rect 6104 12600 8484 12628
rect 8478 12588 8484 12600
rect 8536 12628 8542 12640
rect 10336 12628 10364 12727
rect 10686 12724 10692 12736
rect 10744 12724 10750 12776
rect 10870 12764 10876 12776
rect 10831 12736 10876 12764
rect 10870 12724 10876 12736
rect 10928 12724 10934 12776
rect 11701 12767 11759 12773
rect 11701 12733 11713 12767
rect 11747 12764 11759 12767
rect 11790 12764 11796 12776
rect 11747 12736 11796 12764
rect 11747 12733 11759 12736
rect 11701 12727 11759 12733
rect 11790 12724 11796 12736
rect 11848 12764 11854 12776
rect 12713 12767 12771 12773
rect 11848 12736 12664 12764
rect 11848 12724 11854 12736
rect 8536 12600 10364 12628
rect 11793 12631 11851 12637
rect 8536 12588 8542 12600
rect 11793 12597 11805 12631
rect 11839 12628 11851 12631
rect 12434 12628 12440 12640
rect 11839 12600 12440 12628
rect 11839 12597 11851 12600
rect 11793 12591 11851 12597
rect 12434 12588 12440 12600
rect 12492 12588 12498 12640
rect 12636 12628 12664 12736
rect 12713 12733 12725 12767
rect 12759 12733 12771 12767
rect 12713 12727 12771 12733
rect 13173 12767 13231 12773
rect 13173 12733 13185 12767
rect 13219 12764 13231 12767
rect 13722 12764 13728 12776
rect 13219 12736 13728 12764
rect 13219 12733 13231 12736
rect 13173 12727 13231 12733
rect 12728 12696 12756 12727
rect 13722 12724 13728 12736
rect 13780 12724 13786 12776
rect 13909 12767 13967 12773
rect 13909 12733 13921 12767
rect 13955 12764 13967 12767
rect 13998 12764 14004 12776
rect 13955 12736 14004 12764
rect 13955 12733 13967 12736
rect 13909 12727 13967 12733
rect 13998 12724 14004 12736
rect 14056 12764 14062 12776
rect 14182 12764 14188 12776
rect 14056 12736 14188 12764
rect 14056 12724 14062 12736
rect 14182 12724 14188 12736
rect 14240 12724 14246 12776
rect 15102 12764 15108 12776
rect 15063 12736 15108 12764
rect 15102 12724 15108 12736
rect 15160 12724 15166 12776
rect 15565 12767 15623 12773
rect 15565 12733 15577 12767
rect 15611 12733 15623 12767
rect 15565 12727 15623 12733
rect 13262 12696 13268 12708
rect 12728 12668 13268 12696
rect 13262 12656 13268 12668
rect 13320 12656 13326 12708
rect 13354 12628 13360 12640
rect 12636 12600 13360 12628
rect 13354 12588 13360 12600
rect 13412 12588 13418 12640
rect 13998 12588 14004 12640
rect 14056 12628 14062 12640
rect 14274 12628 14280 12640
rect 14056 12600 14280 12628
rect 14056 12588 14062 12600
rect 14274 12588 14280 12600
rect 14332 12588 14338 12640
rect 15580 12628 15608 12727
rect 15672 12696 15700 12804
rect 15749 12801 15761 12835
rect 15795 12832 15807 12835
rect 16574 12832 16580 12844
rect 15795 12804 16580 12832
rect 15795 12801 15807 12804
rect 15749 12795 15807 12801
rect 16574 12792 16580 12804
rect 16632 12792 16638 12844
rect 15838 12724 15844 12776
rect 15896 12764 15902 12776
rect 16960 12773 16988 12872
rect 18509 12869 18521 12903
rect 18555 12900 18567 12903
rect 19242 12900 19248 12912
rect 18555 12872 19248 12900
rect 18555 12869 18567 12872
rect 18509 12863 18567 12869
rect 19242 12860 19248 12872
rect 19300 12860 19306 12912
rect 17221 12835 17279 12841
rect 17221 12801 17233 12835
rect 17267 12832 17279 12835
rect 18138 12832 18144 12844
rect 17267 12804 18144 12832
rect 17267 12801 17279 12804
rect 17221 12795 17279 12801
rect 18138 12792 18144 12804
rect 18196 12792 18202 12844
rect 19150 12832 19156 12844
rect 19111 12804 19156 12832
rect 19150 12792 19156 12804
rect 19208 12792 19214 12844
rect 20364 12832 20392 12940
rect 20990 12928 20996 12940
rect 21048 12928 21054 12980
rect 22278 12928 22284 12980
rect 22336 12968 22342 12980
rect 22462 12968 22468 12980
rect 22336 12940 22468 12968
rect 22336 12928 22342 12940
rect 22462 12928 22468 12940
rect 22520 12928 22526 12980
rect 22830 12928 22836 12980
rect 22888 12968 22894 12980
rect 24581 12971 24639 12977
rect 24581 12968 24593 12971
rect 22888 12940 24593 12968
rect 22888 12928 22894 12940
rect 24581 12937 24593 12940
rect 24627 12937 24639 12971
rect 32030 12968 32036 12980
rect 24581 12931 24639 12937
rect 31128 12940 32036 12968
rect 20898 12900 20904 12912
rect 20456 12872 20904 12900
rect 20456 12841 20484 12872
rect 20898 12860 20904 12872
rect 20956 12860 20962 12912
rect 22646 12900 22652 12912
rect 22607 12872 22652 12900
rect 22646 12860 22652 12872
rect 22704 12860 22710 12912
rect 28350 12900 28356 12912
rect 27264 12872 28356 12900
rect 19260 12804 20392 12832
rect 20441 12835 20499 12841
rect 16209 12767 16267 12773
rect 16209 12764 16221 12767
rect 15896 12736 16221 12764
rect 15896 12724 15902 12736
rect 16209 12733 16221 12736
rect 16255 12733 16267 12767
rect 16209 12727 16267 12733
rect 16945 12767 17003 12773
rect 16945 12733 16957 12767
rect 16991 12733 17003 12767
rect 18046 12764 18052 12776
rect 18007 12736 18052 12764
rect 16945 12727 17003 12733
rect 16960 12696 16988 12727
rect 18046 12724 18052 12736
rect 18104 12724 18110 12776
rect 18414 12724 18420 12776
rect 18472 12764 18478 12776
rect 18785 12767 18843 12773
rect 18785 12764 18797 12767
rect 18472 12736 18797 12764
rect 18472 12724 18478 12736
rect 18785 12733 18797 12736
rect 18831 12733 18843 12767
rect 18785 12727 18843 12733
rect 17126 12696 17132 12708
rect 15672 12668 16896 12696
rect 16960 12668 17132 12696
rect 16301 12631 16359 12637
rect 16301 12628 16313 12631
rect 15580 12600 16313 12628
rect 16301 12597 16313 12600
rect 16347 12597 16359 12631
rect 16868 12628 16896 12668
rect 17126 12656 17132 12668
rect 17184 12696 17190 12708
rect 19260 12696 19288 12804
rect 20441 12801 20453 12835
rect 20487 12801 20499 12835
rect 20441 12795 20499 12801
rect 22005 12835 22063 12841
rect 22005 12801 22017 12835
rect 22051 12832 22063 12835
rect 22094 12832 22100 12844
rect 22051 12804 22100 12832
rect 22051 12801 22063 12804
rect 22005 12795 22063 12801
rect 22094 12792 22100 12804
rect 22152 12792 22158 12844
rect 19978 12764 19984 12776
rect 19939 12736 19984 12764
rect 19978 12724 19984 12736
rect 20036 12724 20042 12776
rect 20070 12724 20076 12776
rect 20128 12764 20134 12776
rect 20346 12764 20352 12776
rect 20128 12736 20352 12764
rect 20128 12724 20134 12736
rect 20346 12724 20352 12736
rect 20404 12724 20410 12776
rect 20530 12764 20536 12776
rect 20491 12736 20536 12764
rect 20530 12724 20536 12736
rect 20588 12724 20594 12776
rect 20898 12764 20904 12776
rect 20859 12736 20904 12764
rect 20898 12724 20904 12736
rect 20956 12724 20962 12776
rect 21085 12767 21143 12773
rect 21085 12733 21097 12767
rect 21131 12733 21143 12767
rect 21085 12727 21143 12733
rect 21100 12696 21128 12727
rect 21910 12724 21916 12776
rect 21968 12764 21974 12776
rect 22189 12767 22247 12773
rect 22189 12764 22201 12767
rect 21968 12736 22201 12764
rect 21968 12724 21974 12736
rect 22189 12733 22201 12736
rect 22235 12733 22247 12767
rect 22646 12764 22652 12776
rect 22607 12736 22652 12764
rect 22189 12727 22247 12733
rect 22646 12724 22652 12736
rect 22704 12724 22710 12776
rect 24489 12767 24547 12773
rect 24489 12733 24501 12767
rect 24535 12764 24547 12767
rect 25774 12764 25780 12776
rect 24535 12736 25780 12764
rect 24535 12733 24547 12736
rect 24489 12727 24547 12733
rect 25774 12724 25780 12736
rect 25832 12724 25838 12776
rect 26513 12767 26571 12773
rect 26513 12733 26525 12767
rect 26559 12764 26571 12767
rect 27264 12764 27292 12872
rect 28350 12860 28356 12872
rect 28408 12900 28414 12912
rect 28408 12872 29316 12900
rect 28408 12860 28414 12872
rect 27338 12792 27344 12844
rect 27396 12792 27402 12844
rect 27522 12792 27528 12844
rect 27580 12832 27586 12844
rect 27617 12835 27675 12841
rect 27617 12832 27629 12835
rect 27580 12804 27629 12832
rect 27580 12792 27586 12804
rect 27617 12801 27629 12804
rect 27663 12801 27675 12835
rect 27617 12795 27675 12801
rect 26559 12736 27292 12764
rect 27356 12764 27384 12792
rect 29288 12773 29316 12872
rect 29822 12792 29828 12844
rect 29880 12832 29886 12844
rect 30101 12835 30159 12841
rect 30101 12832 30113 12835
rect 29880 12804 30113 12832
rect 29880 12792 29886 12804
rect 30101 12801 30113 12804
rect 30147 12801 30159 12835
rect 30834 12832 30840 12844
rect 30795 12804 30840 12832
rect 30101 12795 30159 12801
rect 30834 12792 30840 12804
rect 30892 12792 30898 12844
rect 27801 12767 27859 12773
rect 27801 12764 27813 12767
rect 27356 12736 27813 12764
rect 26559 12733 26571 12736
rect 26513 12727 26571 12733
rect 27801 12733 27813 12736
rect 27847 12733 27859 12767
rect 27801 12727 27859 12733
rect 29273 12767 29331 12773
rect 29273 12733 29285 12767
rect 29319 12733 29331 12767
rect 29273 12727 29331 12733
rect 30377 12767 30435 12773
rect 30377 12733 30389 12767
rect 30423 12764 30435 12767
rect 31128 12764 31156 12940
rect 32030 12928 32036 12940
rect 32088 12968 32094 12980
rect 32490 12968 32496 12980
rect 32088 12940 32496 12968
rect 32088 12928 32094 12940
rect 32490 12928 32496 12940
rect 32548 12928 32554 12980
rect 36909 12971 36967 12977
rect 36909 12937 36921 12971
rect 36955 12968 36967 12971
rect 38194 12968 38200 12980
rect 36955 12940 38200 12968
rect 36955 12937 36967 12940
rect 36909 12931 36967 12937
rect 38194 12928 38200 12940
rect 38252 12928 38258 12980
rect 31202 12860 31208 12912
rect 31260 12900 31266 12912
rect 31260 12872 33640 12900
rect 31260 12860 31266 12872
rect 31386 12792 31392 12844
rect 31444 12832 31450 12844
rect 31444 12804 32628 12832
rect 31444 12792 31450 12804
rect 31297 12767 31355 12773
rect 31297 12764 31309 12767
rect 30423 12736 31309 12764
rect 30423 12733 30435 12736
rect 30377 12727 30435 12733
rect 31297 12733 31309 12736
rect 31343 12733 31355 12767
rect 31297 12727 31355 12733
rect 31665 12767 31723 12773
rect 31665 12733 31677 12767
rect 31711 12733 31723 12767
rect 31665 12727 31723 12733
rect 17184 12668 19288 12696
rect 20088 12668 21128 12696
rect 27065 12699 27123 12705
rect 17184 12656 17190 12668
rect 18782 12628 18788 12640
rect 16868 12600 18788 12628
rect 16301 12591 16359 12597
rect 18782 12588 18788 12600
rect 18840 12588 18846 12640
rect 19334 12588 19340 12640
rect 19392 12628 19398 12640
rect 20088 12628 20116 12668
rect 27065 12665 27077 12699
rect 27111 12696 27123 12699
rect 27338 12696 27344 12708
rect 27111 12668 27344 12696
rect 27111 12665 27123 12668
rect 27065 12659 27123 12665
rect 27338 12656 27344 12668
rect 27396 12656 27402 12708
rect 27706 12656 27712 12708
rect 27764 12696 27770 12708
rect 27985 12699 28043 12705
rect 27985 12696 27997 12699
rect 27764 12668 27997 12696
rect 27764 12656 27770 12668
rect 27985 12665 27997 12668
rect 28031 12665 28043 12699
rect 28350 12696 28356 12708
rect 28311 12668 28356 12696
rect 27985 12659 28043 12665
rect 28350 12656 28356 12668
rect 28408 12656 28414 12708
rect 29086 12656 29092 12708
rect 29144 12696 29150 12708
rect 30098 12696 30104 12708
rect 29144 12668 30104 12696
rect 29144 12656 29150 12668
rect 30098 12656 30104 12668
rect 30156 12696 30162 12708
rect 30469 12699 30527 12705
rect 30469 12696 30481 12699
rect 30156 12668 30481 12696
rect 30156 12656 30162 12668
rect 30469 12665 30481 12668
rect 30515 12665 30527 12699
rect 30469 12659 30527 12665
rect 31680 12640 31708 12727
rect 31754 12724 31760 12776
rect 31812 12764 31818 12776
rect 32033 12767 32091 12773
rect 32033 12764 32045 12767
rect 31812 12736 32045 12764
rect 31812 12724 31818 12736
rect 32033 12733 32045 12736
rect 32079 12764 32091 12767
rect 32490 12764 32496 12776
rect 32079 12736 32496 12764
rect 32079 12733 32091 12736
rect 32033 12727 32091 12733
rect 32490 12724 32496 12736
rect 32548 12724 32554 12776
rect 32600 12773 32628 12804
rect 32674 12792 32680 12844
rect 32732 12832 32738 12844
rect 32732 12804 32777 12832
rect 32732 12792 32738 12804
rect 32585 12767 32643 12773
rect 32585 12733 32597 12767
rect 32631 12733 32643 12767
rect 33226 12764 33232 12776
rect 33187 12736 33232 12764
rect 32585 12727 32643 12733
rect 33226 12724 33232 12736
rect 33284 12724 33290 12776
rect 33612 12773 33640 12872
rect 37734 12832 37740 12844
rect 37695 12804 37740 12832
rect 37734 12792 37740 12804
rect 37792 12792 37798 12844
rect 39114 12832 39120 12844
rect 39075 12804 39120 12832
rect 39114 12792 39120 12804
rect 39172 12792 39178 12844
rect 33597 12767 33655 12773
rect 33597 12733 33609 12767
rect 33643 12733 33655 12767
rect 34054 12764 34060 12776
rect 34015 12736 34060 12764
rect 33597 12727 33655 12733
rect 34054 12724 34060 12736
rect 34112 12724 34118 12776
rect 34885 12767 34943 12773
rect 34885 12764 34897 12767
rect 34164 12736 34897 12764
rect 31846 12656 31852 12708
rect 31904 12696 31910 12708
rect 34164 12696 34192 12736
rect 34885 12733 34897 12736
rect 34931 12733 34943 12767
rect 34885 12727 34943 12733
rect 35250 12724 35256 12776
rect 35308 12764 35314 12776
rect 35529 12767 35587 12773
rect 35529 12764 35541 12767
rect 35308 12736 35541 12764
rect 35308 12724 35314 12736
rect 35529 12733 35541 12736
rect 35575 12733 35587 12767
rect 36078 12764 36084 12776
rect 36039 12736 36084 12764
rect 35529 12727 35587 12733
rect 36078 12724 36084 12736
rect 36136 12724 36142 12776
rect 36265 12767 36323 12773
rect 36265 12733 36277 12767
rect 36311 12733 36323 12767
rect 36265 12727 36323 12733
rect 31904 12668 34192 12696
rect 31904 12656 31910 12668
rect 34238 12656 34244 12708
rect 34296 12696 34302 12708
rect 34333 12699 34391 12705
rect 34333 12696 34345 12699
rect 34296 12668 34345 12696
rect 34296 12656 34302 12668
rect 34333 12665 34345 12668
rect 34379 12665 34391 12699
rect 34333 12659 34391 12665
rect 34977 12699 35035 12705
rect 34977 12665 34989 12699
rect 35023 12696 35035 12699
rect 36170 12696 36176 12708
rect 35023 12668 36176 12696
rect 35023 12665 35035 12668
rect 34977 12659 35035 12665
rect 36170 12656 36176 12668
rect 36228 12696 36234 12708
rect 36280 12696 36308 12727
rect 36538 12724 36544 12776
rect 36596 12764 36602 12776
rect 36817 12767 36875 12773
rect 36817 12764 36829 12767
rect 36596 12736 36829 12764
rect 36596 12724 36602 12736
rect 36817 12733 36829 12736
rect 36863 12733 36875 12767
rect 36817 12727 36875 12733
rect 37182 12724 37188 12776
rect 37240 12764 37246 12776
rect 37461 12767 37519 12773
rect 37461 12764 37473 12767
rect 37240 12736 37473 12764
rect 37240 12724 37246 12736
rect 37461 12733 37473 12736
rect 37507 12733 37519 12767
rect 37461 12727 37519 12733
rect 36228 12668 36308 12696
rect 36228 12656 36234 12668
rect 19392 12600 20116 12628
rect 19392 12588 19398 12600
rect 20622 12588 20628 12640
rect 20680 12628 20686 12640
rect 23566 12628 23572 12640
rect 20680 12600 23572 12628
rect 20680 12588 20686 12600
rect 23566 12588 23572 12600
rect 23624 12588 23630 12640
rect 27893 12631 27951 12637
rect 27893 12597 27905 12631
rect 27939 12628 27951 12631
rect 29457 12631 29515 12637
rect 29457 12628 29469 12631
rect 27939 12600 29469 12628
rect 27939 12597 27951 12600
rect 27893 12591 27951 12597
rect 29457 12597 29469 12600
rect 29503 12628 29515 12631
rect 29546 12628 29552 12640
rect 29503 12600 29552 12628
rect 29503 12597 29515 12600
rect 29457 12591 29515 12597
rect 29546 12588 29552 12600
rect 29604 12588 29610 12640
rect 30285 12631 30343 12637
rect 30285 12597 30297 12631
rect 30331 12628 30343 12631
rect 31662 12628 31668 12640
rect 30331 12600 31668 12628
rect 30331 12597 30343 12600
rect 30285 12591 30343 12597
rect 31662 12588 31668 12600
rect 31720 12588 31726 12640
rect 1104 12538 39836 12560
rect 1104 12486 19606 12538
rect 19658 12486 19670 12538
rect 19722 12486 19734 12538
rect 19786 12486 19798 12538
rect 19850 12486 39836 12538
rect 1104 12464 39836 12486
rect 3234 12424 3240 12436
rect 3195 12396 3240 12424
rect 3234 12384 3240 12396
rect 3292 12384 3298 12436
rect 10042 12384 10048 12436
rect 10100 12384 10106 12436
rect 11974 12384 11980 12436
rect 12032 12424 12038 12436
rect 12032 12396 13400 12424
rect 12032 12384 12038 12396
rect 6178 12356 6184 12368
rect 6012 12328 6184 12356
rect 1854 12288 1860 12300
rect 1815 12260 1860 12288
rect 1854 12248 1860 12260
rect 1912 12248 1918 12300
rect 4617 12291 4675 12297
rect 4617 12257 4629 12291
rect 4663 12288 4675 12291
rect 4706 12288 4712 12300
rect 4663 12260 4712 12288
rect 4663 12257 4675 12260
rect 4617 12251 4675 12257
rect 4706 12248 4712 12260
rect 4764 12248 4770 12300
rect 5534 12288 5540 12300
rect 5495 12260 5540 12288
rect 5534 12248 5540 12260
rect 5592 12248 5598 12300
rect 6012 12297 6040 12328
rect 6178 12316 6184 12328
rect 6236 12316 6242 12368
rect 6730 12356 6736 12368
rect 6288 12328 6736 12356
rect 6288 12300 6316 12328
rect 6730 12316 6736 12328
rect 6788 12316 6794 12368
rect 7006 12356 7012 12368
rect 6840 12328 7012 12356
rect 5997 12291 6055 12297
rect 5997 12257 6009 12291
rect 6043 12257 6055 12291
rect 6270 12288 6276 12300
rect 6231 12260 6276 12288
rect 5997 12251 6055 12257
rect 6270 12248 6276 12260
rect 6328 12248 6334 12300
rect 6641 12291 6699 12297
rect 6641 12257 6653 12291
rect 6687 12288 6699 12291
rect 6840 12288 6868 12328
rect 7006 12316 7012 12328
rect 7064 12356 7070 12368
rect 8202 12356 8208 12368
rect 7064 12328 8208 12356
rect 7064 12316 7070 12328
rect 8202 12316 8208 12328
rect 8260 12316 8266 12368
rect 10060 12356 10088 12384
rect 8404 12328 10088 12356
rect 6687 12260 6868 12288
rect 6687 12257 6699 12260
rect 6641 12251 6699 12257
rect 7190 12248 7196 12300
rect 7248 12288 7254 12300
rect 7285 12291 7343 12297
rect 7285 12288 7297 12291
rect 7248 12260 7297 12288
rect 7248 12248 7254 12260
rect 7285 12257 7297 12260
rect 7331 12288 7343 12291
rect 7834 12288 7840 12300
rect 7331 12260 7840 12288
rect 7331 12257 7343 12260
rect 7285 12251 7343 12257
rect 7834 12248 7840 12260
rect 7892 12248 7898 12300
rect 8018 12288 8024 12300
rect 7979 12260 8024 12288
rect 8018 12248 8024 12260
rect 8076 12248 8082 12300
rect 8404 12297 8432 12328
rect 11146 12316 11152 12368
rect 11204 12356 11210 12368
rect 11204 12328 13032 12356
rect 11204 12316 11210 12328
rect 8389 12291 8447 12297
rect 8389 12257 8401 12291
rect 8435 12257 8447 12291
rect 8754 12288 8760 12300
rect 8715 12260 8760 12288
rect 8389 12251 8447 12257
rect 8754 12248 8760 12260
rect 8812 12248 8818 12300
rect 9953 12291 10011 12297
rect 9953 12257 9965 12291
rect 9999 12257 10011 12291
rect 9953 12251 10011 12257
rect 10321 12291 10379 12297
rect 10321 12257 10333 12291
rect 10367 12288 10379 12291
rect 10410 12288 10416 12300
rect 10367 12260 10416 12288
rect 10367 12257 10379 12260
rect 10321 12251 10379 12257
rect 2130 12220 2136 12232
rect 2091 12192 2136 12220
rect 2130 12180 2136 12192
rect 2188 12180 2194 12232
rect 6365 12223 6423 12229
rect 6365 12189 6377 12223
rect 6411 12220 6423 12223
rect 7098 12220 7104 12232
rect 6411 12192 7104 12220
rect 6411 12189 6423 12192
rect 6365 12183 6423 12189
rect 7098 12180 7104 12192
rect 7156 12180 7162 12232
rect 8294 12220 8300 12232
rect 8255 12192 8300 12220
rect 8294 12180 8300 12192
rect 8352 12180 8358 12232
rect 9968 12152 9996 12251
rect 10410 12248 10416 12260
rect 10468 12248 10474 12300
rect 10686 12288 10692 12300
rect 10647 12260 10692 12288
rect 10686 12248 10692 12260
rect 10744 12248 10750 12300
rect 11514 12288 11520 12300
rect 11475 12260 11520 12288
rect 11514 12248 11520 12260
rect 11572 12248 11578 12300
rect 11793 12291 11851 12297
rect 11793 12257 11805 12291
rect 11839 12257 11851 12291
rect 11793 12251 11851 12257
rect 10134 12220 10140 12232
rect 10095 12192 10140 12220
rect 10134 12180 10140 12192
rect 10192 12180 10198 12232
rect 10428 12220 10456 12248
rect 11808 12220 11836 12251
rect 11882 12248 11888 12300
rect 11940 12288 11946 12300
rect 13004 12297 13032 12328
rect 13372 12297 13400 12396
rect 13630 12384 13636 12436
rect 13688 12424 13694 12436
rect 17126 12424 17132 12436
rect 13688 12396 17132 12424
rect 13688 12384 13694 12396
rect 17126 12384 17132 12396
rect 17184 12384 17190 12436
rect 18874 12384 18880 12436
rect 18932 12424 18938 12436
rect 23014 12424 23020 12436
rect 18932 12396 21588 12424
rect 18932 12384 18938 12396
rect 13906 12316 13912 12368
rect 13964 12356 13970 12368
rect 14366 12356 14372 12368
rect 13964 12328 14372 12356
rect 13964 12316 13970 12328
rect 14366 12316 14372 12328
rect 14424 12356 14430 12368
rect 16761 12359 16819 12365
rect 14424 12328 15884 12356
rect 14424 12316 14430 12328
rect 12069 12291 12127 12297
rect 12069 12288 12081 12291
rect 11940 12260 12081 12288
rect 11940 12248 11946 12260
rect 12069 12257 12081 12260
rect 12115 12257 12127 12291
rect 12069 12251 12127 12257
rect 12989 12291 13047 12297
rect 12989 12257 13001 12291
rect 13035 12257 13047 12291
rect 12989 12251 13047 12257
rect 13357 12291 13415 12297
rect 13357 12257 13369 12291
rect 13403 12257 13415 12291
rect 13357 12251 13415 12257
rect 14001 12291 14059 12297
rect 14001 12257 14013 12291
rect 14047 12257 14059 12291
rect 14001 12251 14059 12257
rect 14185 12291 14243 12297
rect 14185 12257 14197 12291
rect 14231 12288 14243 12291
rect 14274 12288 14280 12300
rect 14231 12260 14280 12288
rect 14231 12257 14243 12260
rect 14185 12251 14243 12257
rect 12342 12220 12348 12232
rect 10428 12192 12348 12220
rect 12342 12180 12348 12192
rect 12400 12180 12406 12232
rect 12526 12220 12532 12232
rect 12487 12192 12532 12220
rect 12526 12180 12532 12192
rect 12584 12180 12590 12232
rect 14016 12220 14044 12251
rect 14274 12248 14280 12260
rect 14332 12248 14338 12300
rect 14550 12248 14556 12300
rect 14608 12288 14614 12300
rect 15856 12297 15884 12328
rect 16761 12325 16773 12359
rect 16807 12356 16819 12359
rect 18046 12356 18052 12368
rect 16807 12328 18052 12356
rect 16807 12325 16819 12328
rect 16761 12319 16819 12325
rect 18046 12316 18052 12328
rect 18104 12316 18110 12368
rect 18230 12316 18236 12368
rect 18288 12356 18294 12368
rect 18417 12359 18475 12365
rect 18417 12356 18429 12359
rect 18288 12328 18429 12356
rect 18288 12316 18294 12328
rect 18417 12325 18429 12328
rect 18463 12325 18475 12359
rect 18417 12319 18475 12325
rect 19518 12316 19524 12368
rect 19576 12356 19582 12368
rect 20254 12356 20260 12368
rect 19576 12328 20260 12356
rect 19576 12316 19582 12328
rect 20254 12316 20260 12328
rect 20312 12316 20318 12368
rect 15289 12291 15347 12297
rect 15289 12288 15301 12291
rect 14608 12260 15301 12288
rect 14608 12248 14614 12260
rect 15289 12257 15301 12260
rect 15335 12257 15347 12291
rect 15289 12251 15347 12257
rect 15841 12291 15899 12297
rect 15841 12257 15853 12291
rect 15887 12257 15899 12291
rect 17402 12288 17408 12300
rect 17363 12260 17408 12288
rect 15841 12251 15899 12257
rect 17402 12248 17408 12260
rect 17460 12248 17466 12300
rect 17773 12291 17831 12297
rect 17773 12257 17785 12291
rect 17819 12288 17831 12291
rect 17954 12288 17960 12300
rect 17819 12260 17960 12288
rect 17819 12257 17831 12260
rect 17773 12251 17831 12257
rect 17954 12248 17960 12260
rect 18012 12248 18018 12300
rect 19058 12288 19064 12300
rect 19019 12260 19064 12288
rect 19058 12248 19064 12260
rect 19116 12248 19122 12300
rect 19426 12288 19432 12300
rect 19387 12260 19432 12288
rect 19426 12248 19432 12260
rect 19484 12248 19490 12300
rect 20070 12288 20076 12300
rect 20031 12260 20076 12288
rect 20070 12248 20076 12260
rect 20128 12248 20134 12300
rect 20901 12291 20959 12297
rect 20901 12257 20913 12291
rect 20947 12257 20959 12291
rect 20901 12251 20959 12257
rect 14016 12192 15424 12220
rect 11514 12152 11520 12164
rect 9968 12124 11520 12152
rect 11514 12112 11520 12124
rect 11572 12112 11578 12164
rect 15396 12161 15424 12192
rect 17218 12180 17224 12232
rect 17276 12220 17282 12232
rect 17313 12223 17371 12229
rect 17313 12220 17325 12223
rect 17276 12192 17325 12220
rect 17276 12180 17282 12192
rect 17313 12189 17325 12192
rect 17359 12189 17371 12223
rect 17313 12183 17371 12189
rect 17865 12223 17923 12229
rect 17865 12189 17877 12223
rect 17911 12220 17923 12223
rect 18230 12220 18236 12232
rect 17911 12192 18236 12220
rect 17911 12189 17923 12192
rect 17865 12183 17923 12189
rect 15381 12155 15439 12161
rect 15381 12121 15393 12155
rect 15427 12121 15439 12155
rect 17328 12152 17356 12183
rect 18230 12180 18236 12192
rect 18288 12180 18294 12232
rect 18969 12223 19027 12229
rect 18969 12189 18981 12223
rect 19015 12220 19027 12223
rect 19242 12220 19248 12232
rect 19015 12192 19248 12220
rect 19015 12189 19027 12192
rect 18969 12183 19027 12189
rect 18984 12152 19012 12183
rect 19242 12180 19248 12192
rect 19300 12180 19306 12232
rect 19521 12223 19579 12229
rect 19521 12189 19533 12223
rect 19567 12220 19579 12223
rect 19886 12220 19892 12232
rect 19567 12192 19892 12220
rect 19567 12189 19579 12192
rect 19521 12183 19579 12189
rect 19886 12180 19892 12192
rect 19944 12220 19950 12232
rect 20162 12220 20168 12232
rect 19944 12192 20168 12220
rect 19944 12180 19950 12192
rect 20162 12180 20168 12192
rect 20220 12220 20226 12232
rect 20916 12220 20944 12251
rect 21082 12248 21088 12300
rect 21140 12288 21146 12300
rect 21453 12291 21511 12297
rect 21453 12288 21465 12291
rect 21140 12260 21465 12288
rect 21140 12248 21146 12260
rect 21453 12257 21465 12260
rect 21499 12257 21511 12291
rect 21453 12251 21511 12257
rect 20220 12192 20944 12220
rect 21560 12220 21588 12396
rect 22756 12396 23020 12424
rect 22465 12291 22523 12297
rect 22465 12257 22477 12291
rect 22511 12288 22523 12291
rect 22756 12288 22784 12396
rect 23014 12384 23020 12396
rect 23072 12384 23078 12436
rect 26786 12384 26792 12436
rect 26844 12424 26850 12436
rect 27522 12424 27528 12436
rect 26844 12396 27528 12424
rect 26844 12384 26850 12396
rect 27522 12384 27528 12396
rect 27580 12384 27586 12436
rect 27706 12384 27712 12436
rect 27764 12424 27770 12436
rect 28074 12424 28080 12436
rect 27764 12396 28080 12424
rect 27764 12384 27770 12396
rect 28074 12384 28080 12396
rect 28132 12424 28138 12436
rect 28132 12396 28488 12424
rect 28132 12384 28138 12396
rect 23750 12356 23756 12368
rect 23032 12328 23756 12356
rect 22511 12260 22784 12288
rect 22511 12257 22523 12260
rect 22465 12251 22523 12257
rect 22830 12248 22836 12300
rect 22888 12288 22894 12300
rect 23032 12297 23060 12328
rect 23750 12316 23756 12328
rect 23808 12316 23814 12368
rect 25774 12356 25780 12368
rect 25735 12328 25780 12356
rect 25774 12316 25780 12328
rect 25832 12316 25838 12368
rect 28350 12356 28356 12368
rect 26988 12328 28356 12356
rect 26988 12297 27016 12328
rect 28350 12316 28356 12328
rect 28408 12316 28414 12368
rect 28460 12356 28488 12396
rect 29086 12384 29092 12436
rect 29144 12424 29150 12436
rect 29365 12427 29423 12433
rect 29365 12424 29377 12427
rect 29144 12396 29377 12424
rect 29144 12384 29150 12396
rect 29365 12393 29377 12396
rect 29411 12393 29423 12427
rect 29365 12387 29423 12393
rect 29822 12384 29828 12436
rect 29880 12424 29886 12436
rect 30193 12427 30251 12433
rect 30193 12424 30205 12427
rect 29880 12396 30205 12424
rect 29880 12384 29886 12396
rect 30193 12393 30205 12396
rect 30239 12424 30251 12427
rect 30742 12424 30748 12436
rect 30239 12396 30748 12424
rect 30239 12393 30251 12396
rect 30193 12387 30251 12393
rect 30742 12384 30748 12396
rect 30800 12384 30806 12436
rect 32306 12384 32312 12436
rect 32364 12424 32370 12436
rect 32364 12396 33364 12424
rect 32364 12384 32370 12396
rect 30377 12359 30435 12365
rect 30377 12356 30389 12359
rect 28460 12328 30389 12356
rect 30377 12325 30389 12328
rect 30423 12356 30435 12359
rect 30423 12328 31248 12356
rect 30423 12325 30435 12328
rect 30377 12319 30435 12325
rect 22925 12291 22983 12297
rect 22925 12288 22937 12291
rect 22888 12260 22937 12288
rect 22888 12248 22894 12260
rect 22925 12257 22937 12260
rect 22971 12257 22983 12291
rect 22925 12251 22983 12257
rect 23017 12291 23075 12297
rect 23017 12257 23029 12291
rect 23063 12257 23075 12291
rect 24397 12291 24455 12297
rect 24397 12288 24409 12291
rect 23017 12251 23075 12257
rect 23584 12260 24409 12288
rect 23584 12229 23612 12260
rect 24397 12257 24409 12260
rect 24443 12257 24455 12291
rect 24397 12251 24455 12257
rect 26973 12291 27031 12297
rect 26973 12257 26985 12291
rect 27019 12257 27031 12291
rect 27614 12288 27620 12300
rect 27575 12260 27620 12288
rect 26973 12251 27031 12257
rect 27614 12248 27620 12260
rect 27672 12248 27678 12300
rect 28258 12288 28264 12300
rect 28219 12260 28264 12288
rect 28258 12248 28264 12260
rect 28316 12248 28322 12300
rect 29181 12291 29239 12297
rect 29181 12257 29193 12291
rect 29227 12288 29239 12291
rect 29546 12288 29552 12300
rect 29227 12260 29552 12288
rect 29227 12257 29239 12260
rect 29181 12251 29239 12257
rect 29546 12248 29552 12260
rect 29604 12248 29610 12300
rect 30282 12288 30288 12300
rect 30243 12260 30288 12288
rect 30282 12248 30288 12260
rect 30340 12248 30346 12300
rect 31220 12297 31248 12328
rect 31205 12291 31263 12297
rect 31205 12257 31217 12291
rect 31251 12288 31263 12291
rect 31386 12288 31392 12300
rect 31251 12260 31392 12288
rect 31251 12257 31263 12260
rect 31205 12251 31263 12257
rect 31386 12248 31392 12260
rect 31444 12248 31450 12300
rect 32122 12288 32128 12300
rect 32083 12260 32128 12288
rect 32122 12248 32128 12260
rect 32180 12248 32186 12300
rect 32585 12291 32643 12297
rect 32585 12257 32597 12291
rect 32631 12257 32643 12291
rect 32585 12251 32643 12257
rect 22373 12223 22431 12229
rect 22373 12220 22385 12223
rect 21560 12192 22385 12220
rect 20220 12180 20226 12192
rect 22373 12189 22385 12192
rect 22419 12189 22431 12223
rect 22373 12183 22431 12189
rect 23569 12223 23627 12229
rect 23569 12189 23581 12223
rect 23615 12189 23627 12223
rect 24118 12220 24124 12232
rect 24079 12192 24124 12220
rect 23569 12183 23627 12189
rect 17328 12124 19012 12152
rect 19076 12124 20852 12152
rect 15381 12115 15439 12121
rect 2774 12044 2780 12096
rect 2832 12084 2838 12096
rect 3694 12084 3700 12096
rect 2832 12056 3700 12084
rect 2832 12044 2838 12056
rect 3694 12044 3700 12056
rect 3752 12084 3758 12096
rect 4433 12087 4491 12093
rect 4433 12084 4445 12087
rect 3752 12056 4445 12084
rect 3752 12044 3758 12056
rect 4433 12053 4445 12056
rect 4479 12053 4491 12087
rect 4433 12047 4491 12053
rect 13630 12044 13636 12096
rect 13688 12084 13694 12096
rect 19076 12084 19104 12124
rect 13688 12056 19104 12084
rect 13688 12044 13694 12056
rect 19242 12044 19248 12096
rect 19300 12084 19306 12096
rect 20254 12084 20260 12096
rect 19300 12056 20260 12084
rect 19300 12044 19306 12056
rect 20254 12044 20260 12056
rect 20312 12044 20318 12096
rect 20824 12084 20852 12124
rect 20898 12112 20904 12164
rect 20956 12152 20962 12164
rect 20993 12155 21051 12161
rect 20993 12152 21005 12155
rect 20956 12124 21005 12152
rect 20956 12112 20962 12124
rect 20993 12121 21005 12124
rect 21039 12121 21051 12155
rect 22388 12152 22416 12183
rect 24118 12180 24124 12192
rect 24176 12220 24182 12232
rect 24486 12220 24492 12232
rect 24176 12192 24492 12220
rect 24176 12180 24182 12192
rect 24486 12180 24492 12192
rect 24544 12180 24550 12232
rect 27065 12223 27123 12229
rect 27065 12189 27077 12223
rect 27111 12220 27123 12223
rect 28445 12223 28503 12229
rect 28445 12220 28457 12223
rect 27111 12192 28457 12220
rect 27111 12189 27123 12192
rect 27065 12183 27123 12189
rect 28445 12189 28457 12192
rect 28491 12189 28503 12223
rect 28445 12183 28503 12189
rect 30009 12223 30067 12229
rect 30009 12189 30021 12223
rect 30055 12220 30067 12223
rect 30558 12220 30564 12232
rect 30055 12192 30564 12220
rect 30055 12189 30067 12192
rect 30009 12183 30067 12189
rect 30558 12180 30564 12192
rect 30616 12180 30622 12232
rect 30745 12223 30803 12229
rect 30745 12189 30757 12223
rect 30791 12189 30803 12223
rect 32600 12220 32628 12251
rect 32674 12248 32680 12300
rect 32732 12288 32738 12300
rect 33336 12297 33364 12396
rect 39114 12356 39120 12368
rect 38396 12328 39120 12356
rect 32861 12291 32919 12297
rect 32861 12288 32873 12291
rect 32732 12260 32873 12288
rect 32732 12248 32738 12260
rect 32861 12257 32873 12260
rect 32907 12257 32919 12291
rect 32861 12251 32919 12257
rect 33321 12291 33379 12297
rect 33321 12257 33333 12291
rect 33367 12257 33379 12291
rect 34054 12288 34060 12300
rect 33967 12260 34060 12288
rect 33321 12251 33379 12257
rect 34054 12248 34060 12260
rect 34112 12288 34118 12300
rect 34112 12260 35940 12288
rect 34112 12248 34118 12260
rect 30745 12183 30803 12189
rect 30852 12192 32628 12220
rect 33045 12223 33103 12229
rect 22830 12152 22836 12164
rect 22388 12124 22836 12152
rect 20993 12115 21051 12121
rect 22830 12112 22836 12124
rect 22888 12112 22894 12164
rect 27893 12155 27951 12161
rect 27893 12121 27905 12155
rect 27939 12152 27951 12155
rect 28074 12152 28080 12164
rect 27939 12124 28080 12152
rect 27939 12121 27951 12124
rect 27893 12115 27951 12121
rect 28074 12112 28080 12124
rect 28132 12112 28138 12164
rect 28902 12112 28908 12164
rect 28960 12152 28966 12164
rect 30760 12152 30788 12183
rect 28960 12124 30788 12152
rect 28960 12112 28966 12124
rect 22554 12084 22560 12096
rect 20824 12056 22560 12084
rect 22554 12044 22560 12056
rect 22612 12044 22618 12096
rect 27798 12044 27804 12096
rect 27856 12084 27862 12096
rect 30852 12084 30880 12192
rect 33045 12189 33057 12223
rect 33091 12220 33103 12223
rect 33226 12220 33232 12232
rect 33091 12192 33232 12220
rect 33091 12189 33103 12192
rect 33045 12183 33103 12189
rect 33226 12180 33232 12192
rect 33284 12180 33290 12232
rect 34514 12220 34520 12232
rect 34475 12192 34520 12220
rect 34514 12180 34520 12192
rect 34572 12180 34578 12232
rect 34790 12220 34796 12232
rect 34751 12192 34796 12220
rect 34790 12180 34796 12192
rect 34848 12180 34854 12232
rect 35912 12229 35940 12260
rect 36538 12248 36544 12300
rect 36596 12288 36602 12300
rect 38396 12297 38424 12328
rect 39114 12316 39120 12328
rect 39172 12316 39178 12368
rect 37001 12291 37059 12297
rect 37001 12288 37013 12291
rect 36596 12260 37013 12288
rect 36596 12248 36602 12260
rect 37001 12257 37013 12260
rect 37047 12257 37059 12291
rect 37001 12251 37059 12257
rect 38381 12291 38439 12297
rect 38381 12257 38393 12291
rect 38427 12257 38439 12291
rect 38562 12288 38568 12300
rect 38523 12260 38568 12288
rect 38381 12251 38439 12257
rect 38562 12248 38568 12260
rect 38620 12248 38626 12300
rect 38749 12291 38807 12297
rect 38749 12257 38761 12291
rect 38795 12257 38807 12291
rect 38749 12251 38807 12257
rect 35897 12223 35955 12229
rect 35897 12189 35909 12223
rect 35943 12189 35955 12223
rect 35897 12183 35955 12189
rect 37093 12223 37151 12229
rect 37093 12189 37105 12223
rect 37139 12220 37151 12223
rect 38470 12220 38476 12232
rect 37139 12192 38476 12220
rect 37139 12189 37151 12192
rect 37093 12183 37151 12189
rect 38470 12180 38476 12192
rect 38528 12220 38534 12232
rect 38764 12220 38792 12251
rect 38528 12192 38792 12220
rect 38528 12180 38534 12192
rect 31294 12084 31300 12096
rect 27856 12056 30880 12084
rect 31255 12056 31300 12084
rect 27856 12044 27862 12056
rect 31294 12044 31300 12056
rect 31352 12044 31358 12096
rect 1104 11994 39836 12016
rect 1104 11942 4246 11994
rect 4298 11942 4310 11994
rect 4362 11942 4374 11994
rect 4426 11942 4438 11994
rect 4490 11942 34966 11994
rect 35018 11942 35030 11994
rect 35082 11942 35094 11994
rect 35146 11942 35158 11994
rect 35210 11942 39836 11994
rect 1104 11920 39836 11942
rect 2130 11840 2136 11892
rect 2188 11880 2194 11892
rect 4709 11883 4767 11889
rect 4709 11880 4721 11883
rect 2188 11852 4721 11880
rect 2188 11840 2194 11852
rect 4709 11849 4721 11852
rect 4755 11849 4767 11883
rect 4709 11843 4767 11849
rect 8389 11883 8447 11889
rect 8389 11849 8401 11883
rect 8435 11880 8447 11883
rect 8478 11880 8484 11892
rect 8435 11852 8484 11880
rect 8435 11849 8447 11852
rect 8389 11843 8447 11849
rect 8478 11840 8484 11852
rect 8536 11840 8542 11892
rect 9309 11883 9367 11889
rect 9309 11849 9321 11883
rect 9355 11880 9367 11883
rect 9674 11880 9680 11892
rect 9355 11852 9680 11880
rect 9355 11849 9367 11852
rect 9309 11843 9367 11849
rect 9674 11840 9680 11852
rect 9732 11840 9738 11892
rect 12342 11840 12348 11892
rect 12400 11880 12406 11892
rect 12621 11883 12679 11889
rect 12621 11880 12633 11883
rect 12400 11852 12633 11880
rect 12400 11840 12406 11852
rect 12621 11849 12633 11852
rect 12667 11849 12679 11883
rect 15378 11880 15384 11892
rect 12621 11843 12679 11849
rect 14016 11852 15384 11880
rect 14016 11812 14044 11852
rect 15378 11840 15384 11852
rect 15436 11840 15442 11892
rect 18230 11880 18236 11892
rect 18191 11852 18236 11880
rect 18230 11840 18236 11852
rect 18288 11840 18294 11892
rect 19610 11880 19616 11892
rect 18432 11852 19616 11880
rect 9232 11784 14044 11812
rect 15749 11815 15807 11821
rect 3329 11747 3387 11753
rect 3329 11713 3341 11747
rect 3375 11744 3387 11747
rect 3510 11744 3516 11756
rect 3375 11716 3516 11744
rect 3375 11713 3387 11716
rect 3329 11707 3387 11713
rect 3510 11704 3516 11716
rect 3568 11704 3574 11756
rect 7098 11744 7104 11756
rect 7059 11716 7104 11744
rect 7098 11704 7104 11716
rect 7156 11704 7162 11756
rect 2682 11676 2688 11688
rect 2643 11648 2688 11676
rect 2682 11636 2688 11648
rect 2740 11636 2746 11688
rect 3605 11679 3663 11685
rect 3605 11645 3617 11679
rect 3651 11676 3663 11679
rect 4890 11676 4896 11688
rect 3651 11648 4896 11676
rect 3651 11645 3663 11648
rect 3605 11639 3663 11645
rect 4890 11636 4896 11648
rect 4948 11636 4954 11688
rect 6825 11679 6883 11685
rect 6825 11645 6837 11679
rect 6871 11676 6883 11679
rect 6914 11676 6920 11688
rect 6871 11648 6920 11676
rect 6871 11645 6883 11648
rect 6825 11639 6883 11645
rect 6914 11636 6920 11648
rect 6972 11636 6978 11688
rect 9232 11685 9260 11784
rect 15749 11781 15761 11815
rect 15795 11812 15807 11815
rect 16114 11812 16120 11824
rect 15795 11784 16120 11812
rect 15795 11781 15807 11784
rect 15749 11775 15807 11781
rect 16114 11772 16120 11784
rect 16172 11772 16178 11824
rect 16574 11772 16580 11824
rect 16632 11812 16638 11824
rect 18432 11812 18460 11852
rect 19610 11840 19616 11852
rect 19668 11880 19674 11892
rect 20622 11880 20628 11892
rect 19668 11852 20628 11880
rect 19668 11840 19674 11852
rect 20622 11840 20628 11852
rect 20680 11840 20686 11892
rect 23658 11880 23664 11892
rect 20732 11852 23664 11880
rect 16632 11784 18460 11812
rect 19153 11815 19211 11821
rect 16632 11772 16638 11784
rect 19153 11781 19165 11815
rect 19199 11812 19211 11815
rect 19334 11812 19340 11824
rect 19199 11784 19340 11812
rect 19199 11781 19211 11784
rect 19153 11775 19211 11781
rect 19334 11772 19340 11784
rect 19392 11772 19398 11824
rect 20732 11821 20760 11852
rect 23658 11840 23664 11852
rect 23716 11840 23722 11892
rect 26878 11880 26884 11892
rect 24228 11852 26884 11880
rect 20717 11815 20775 11821
rect 20717 11781 20729 11815
rect 20763 11781 20775 11815
rect 20717 11775 20775 11781
rect 22281 11815 22339 11821
rect 22281 11781 22293 11815
rect 22327 11812 22339 11815
rect 22646 11812 22652 11824
rect 22327 11784 22652 11812
rect 22327 11781 22339 11784
rect 22281 11775 22339 11781
rect 22646 11772 22652 11784
rect 22704 11772 22710 11824
rect 10778 11744 10784 11756
rect 10739 11716 10784 11744
rect 10778 11704 10784 11716
rect 10836 11704 10842 11756
rect 13814 11744 13820 11756
rect 13775 11716 13820 11744
rect 13814 11704 13820 11716
rect 13872 11704 13878 11756
rect 14090 11704 14096 11756
rect 14148 11744 14154 11756
rect 16592 11744 16620 11772
rect 19978 11744 19984 11756
rect 14148 11716 14228 11744
rect 14148 11704 14154 11716
rect 9217 11679 9275 11685
rect 9217 11645 9229 11679
rect 9263 11645 9275 11679
rect 9858 11676 9864 11688
rect 9819 11648 9864 11676
rect 9217 11639 9275 11645
rect 9858 11636 9864 11648
rect 9916 11636 9922 11688
rect 10134 11636 10140 11688
rect 10192 11676 10198 11688
rect 10229 11679 10287 11685
rect 10229 11676 10241 11679
rect 10192 11648 10241 11676
rect 10192 11636 10198 11648
rect 10229 11645 10241 11648
rect 10275 11645 10287 11679
rect 10229 11639 10287 11645
rect 10873 11679 10931 11685
rect 10873 11645 10885 11679
rect 10919 11676 10931 11679
rect 11054 11676 11060 11688
rect 10919 11648 11060 11676
rect 10919 11645 10931 11648
rect 10873 11639 10931 11645
rect 11054 11636 11060 11648
rect 11112 11636 11118 11688
rect 11517 11679 11575 11685
rect 11517 11645 11529 11679
rect 11563 11645 11575 11679
rect 12434 11676 12440 11688
rect 12347 11648 12440 11676
rect 11517 11639 11575 11645
rect 11532 11608 11560 11639
rect 12434 11636 12440 11648
rect 12492 11676 12498 11688
rect 13449 11679 13507 11685
rect 12492 11648 13400 11676
rect 12492 11636 12498 11648
rect 12894 11608 12900 11620
rect 11532 11580 12900 11608
rect 12894 11568 12900 11580
rect 12952 11568 12958 11620
rect 2774 11500 2780 11552
rect 2832 11540 2838 11552
rect 2832 11512 2877 11540
rect 2832 11500 2838 11512
rect 8386 11500 8392 11552
rect 8444 11540 8450 11552
rect 9122 11540 9128 11552
rect 8444 11512 9128 11540
rect 8444 11500 8450 11512
rect 9122 11500 9128 11512
rect 9180 11540 9186 11552
rect 11701 11543 11759 11549
rect 11701 11540 11713 11543
rect 9180 11512 11713 11540
rect 9180 11500 9186 11512
rect 11701 11509 11713 11512
rect 11747 11540 11759 11543
rect 11882 11540 11888 11552
rect 11747 11512 11888 11540
rect 11747 11509 11759 11512
rect 11701 11503 11759 11509
rect 11882 11500 11888 11512
rect 11940 11500 11946 11552
rect 13372 11540 13400 11648
rect 13449 11645 13461 11679
rect 13495 11645 13507 11679
rect 13906 11676 13912 11688
rect 13867 11648 13912 11676
rect 13449 11639 13507 11645
rect 13464 11608 13492 11639
rect 13906 11636 13912 11648
rect 13964 11636 13970 11688
rect 14200 11685 14228 11716
rect 16224 11716 16620 11744
rect 19076 11716 19984 11744
rect 14185 11679 14243 11685
rect 14185 11645 14197 11679
rect 14231 11645 14243 11679
rect 14185 11639 14243 11645
rect 15381 11679 15439 11685
rect 15381 11645 15393 11679
rect 15427 11676 15439 11679
rect 15657 11679 15715 11685
rect 15657 11676 15669 11679
rect 15427 11648 15669 11676
rect 15427 11645 15439 11648
rect 15381 11639 15439 11645
rect 15657 11645 15669 11648
rect 15703 11676 15715 11679
rect 15838 11676 15844 11688
rect 15703 11648 15844 11676
rect 15703 11645 15715 11648
rect 15657 11639 15715 11645
rect 15838 11636 15844 11648
rect 15896 11636 15902 11688
rect 16224 11685 16252 11716
rect 16209 11679 16267 11685
rect 16209 11645 16221 11679
rect 16255 11645 16267 11679
rect 16209 11639 16267 11645
rect 16298 11636 16304 11688
rect 16356 11676 16362 11688
rect 17218 11676 17224 11688
rect 16356 11648 16401 11676
rect 17179 11648 17224 11676
rect 16356 11636 16362 11648
rect 17218 11636 17224 11648
rect 17276 11636 17282 11688
rect 17954 11636 17960 11688
rect 18012 11676 18018 11688
rect 19076 11685 19104 11716
rect 19978 11704 19984 11716
rect 20036 11704 20042 11756
rect 20254 11704 20260 11756
rect 20312 11704 20318 11756
rect 24228 11744 24256 11852
rect 26878 11840 26884 11852
rect 26936 11840 26942 11892
rect 27614 11840 27620 11892
rect 27672 11880 27678 11892
rect 27798 11880 27804 11892
rect 27672 11852 27804 11880
rect 27672 11840 27678 11852
rect 27798 11840 27804 11852
rect 27856 11840 27862 11892
rect 28537 11883 28595 11889
rect 28537 11849 28549 11883
rect 28583 11880 28595 11883
rect 31846 11880 31852 11892
rect 28583 11852 31852 11880
rect 28583 11849 28595 11852
rect 28537 11843 28595 11849
rect 31846 11840 31852 11852
rect 31904 11840 31910 11892
rect 32125 11883 32183 11889
rect 32125 11849 32137 11883
rect 32171 11880 32183 11883
rect 33686 11880 33692 11892
rect 32171 11852 33692 11880
rect 32171 11849 32183 11852
rect 32125 11843 32183 11849
rect 33686 11840 33692 11852
rect 33744 11840 33750 11892
rect 24302 11772 24308 11824
rect 24360 11812 24366 11824
rect 24360 11784 29316 11812
rect 24360 11772 24366 11784
rect 28994 11744 29000 11756
rect 21008 11716 22600 11744
rect 18049 11679 18107 11685
rect 18049 11676 18061 11679
rect 18012 11648 18061 11676
rect 18012 11636 18018 11648
rect 18049 11645 18061 11648
rect 18095 11645 18107 11679
rect 18049 11639 18107 11645
rect 19061 11679 19119 11685
rect 19061 11645 19073 11679
rect 19107 11645 19119 11679
rect 19610 11676 19616 11688
rect 19571 11648 19616 11676
rect 19061 11639 19119 11645
rect 19610 11636 19616 11648
rect 19668 11636 19674 11688
rect 19889 11679 19947 11685
rect 19889 11645 19901 11679
rect 19935 11645 19947 11679
rect 20272 11676 20300 11704
rect 21008 11688 21036 11716
rect 20622 11676 20628 11688
rect 20272 11648 20628 11676
rect 19889 11639 19947 11645
rect 17770 11608 17776 11620
rect 13464 11580 17776 11608
rect 17770 11568 17776 11580
rect 17828 11568 17834 11620
rect 19904 11608 19932 11639
rect 20622 11636 20628 11648
rect 20680 11636 20686 11688
rect 20990 11676 20996 11688
rect 20951 11648 20996 11676
rect 20990 11636 20996 11648
rect 21048 11636 21054 11688
rect 21453 11679 21511 11685
rect 21453 11645 21465 11679
rect 21499 11676 21511 11679
rect 22002 11676 22008 11688
rect 21499 11648 22008 11676
rect 21499 11645 21511 11648
rect 21453 11639 21511 11645
rect 22002 11636 22008 11648
rect 22060 11636 22066 11688
rect 22572 11685 22600 11716
rect 22664 11716 24256 11744
rect 26620 11716 29000 11744
rect 22664 11688 22692 11716
rect 22097 11679 22155 11685
rect 22097 11645 22109 11679
rect 22143 11645 22155 11679
rect 22097 11639 22155 11645
rect 22557 11679 22615 11685
rect 22557 11645 22569 11679
rect 22603 11645 22615 11679
rect 22557 11639 22615 11645
rect 21542 11608 21548 11620
rect 19904 11580 21548 11608
rect 21542 11568 21548 11580
rect 21600 11568 21606 11620
rect 22112 11608 22140 11639
rect 22646 11636 22652 11688
rect 22704 11636 22710 11688
rect 22922 11676 22928 11688
rect 22883 11648 22928 11676
rect 22922 11636 22928 11648
rect 22980 11636 22986 11688
rect 23198 11636 23204 11688
rect 23256 11676 23262 11688
rect 23842 11676 23848 11688
rect 23256 11648 23848 11676
rect 23256 11636 23262 11648
rect 23842 11636 23848 11648
rect 23900 11636 23906 11688
rect 25409 11679 25467 11685
rect 25409 11645 25421 11679
rect 25455 11645 25467 11679
rect 25409 11639 25467 11645
rect 26145 11679 26203 11685
rect 26145 11645 26157 11679
rect 26191 11676 26203 11679
rect 26620 11676 26648 11716
rect 28994 11704 29000 11716
rect 29052 11704 29058 11756
rect 29288 11688 29316 11784
rect 30466 11772 30472 11824
rect 30524 11812 30530 11824
rect 31481 11815 31539 11821
rect 31481 11812 31493 11815
rect 30524 11784 31493 11812
rect 30524 11772 30530 11784
rect 31481 11781 31493 11784
rect 31527 11812 31539 11815
rect 31662 11812 31668 11824
rect 31527 11784 31668 11812
rect 31527 11781 31539 11784
rect 31481 11775 31539 11781
rect 31662 11772 31668 11784
rect 31720 11772 31726 11824
rect 33505 11815 33563 11821
rect 33505 11781 33517 11815
rect 33551 11812 33563 11815
rect 34790 11812 34796 11824
rect 33551 11784 34796 11812
rect 33551 11781 33563 11784
rect 33505 11775 33563 11781
rect 34790 11772 34796 11784
rect 34848 11772 34854 11824
rect 35621 11815 35679 11821
rect 35621 11781 35633 11815
rect 35667 11812 35679 11815
rect 36722 11812 36728 11824
rect 35667 11784 36728 11812
rect 35667 11781 35679 11784
rect 35621 11775 35679 11781
rect 36722 11772 36728 11784
rect 36780 11772 36786 11824
rect 29454 11744 29460 11756
rect 29415 11716 29460 11744
rect 29454 11704 29460 11716
rect 29512 11704 29518 11756
rect 30650 11744 30656 11756
rect 30116 11716 30656 11744
rect 26191 11648 26648 11676
rect 26697 11679 26755 11685
rect 26191 11645 26203 11648
rect 26145 11639 26203 11645
rect 26697 11645 26709 11679
rect 26743 11676 26755 11679
rect 27157 11679 27215 11685
rect 27157 11676 27169 11679
rect 26743 11648 27169 11676
rect 26743 11645 26755 11648
rect 26697 11639 26755 11645
rect 27157 11645 27169 11648
rect 27203 11645 27215 11679
rect 27338 11676 27344 11688
rect 27299 11648 27344 11676
rect 27157 11639 27215 11645
rect 21652 11580 22140 11608
rect 13906 11540 13912 11552
rect 13372 11512 13912 11540
rect 13906 11500 13912 11512
rect 13964 11540 13970 11552
rect 15381 11543 15439 11549
rect 15381 11540 15393 11543
rect 13964 11512 15393 11540
rect 13964 11500 13970 11512
rect 15381 11509 15393 11512
rect 15427 11509 15439 11543
rect 15381 11503 15439 11509
rect 17405 11543 17463 11549
rect 17405 11509 17417 11543
rect 17451 11540 17463 11543
rect 19150 11540 19156 11552
rect 17451 11512 19156 11540
rect 17451 11509 17463 11512
rect 17405 11503 17463 11509
rect 19150 11500 19156 11512
rect 19208 11500 19214 11552
rect 20622 11500 20628 11552
rect 20680 11540 20686 11552
rect 21652 11540 21680 11580
rect 22186 11568 22192 11620
rect 22244 11608 22250 11620
rect 23934 11608 23940 11620
rect 22244 11580 23940 11608
rect 22244 11568 22250 11580
rect 23934 11568 23940 11580
rect 23992 11568 23998 11620
rect 20680 11512 21680 11540
rect 20680 11500 20686 11512
rect 22002 11500 22008 11552
rect 22060 11540 22066 11552
rect 25424 11540 25452 11639
rect 27338 11636 27344 11648
rect 27396 11636 27402 11688
rect 27706 11676 27712 11688
rect 27667 11648 27712 11676
rect 27706 11636 27712 11648
rect 27764 11636 27770 11688
rect 27798 11636 27804 11688
rect 27856 11676 27862 11688
rect 27893 11679 27951 11685
rect 27893 11676 27905 11679
rect 27856 11648 27905 11676
rect 27856 11636 27862 11648
rect 27893 11645 27905 11648
rect 27939 11645 27951 11679
rect 27893 11639 27951 11645
rect 27982 11636 27988 11688
rect 28040 11676 28046 11688
rect 28077 11679 28135 11685
rect 28077 11676 28089 11679
rect 28040 11648 28089 11676
rect 28040 11636 28046 11648
rect 28077 11645 28089 11648
rect 28123 11645 28135 11679
rect 28077 11639 28135 11645
rect 29270 11636 29276 11688
rect 29328 11676 29334 11688
rect 30116 11685 30144 11716
rect 30650 11704 30656 11716
rect 30708 11704 30714 11756
rect 34054 11744 34060 11756
rect 30760 11716 34060 11744
rect 29365 11679 29423 11685
rect 29365 11676 29377 11679
rect 29328 11648 29377 11676
rect 29328 11636 29334 11648
rect 29365 11645 29377 11648
rect 29411 11645 29423 11679
rect 29365 11639 29423 11645
rect 30101 11679 30159 11685
rect 30101 11645 30113 11679
rect 30147 11645 30159 11679
rect 30101 11639 30159 11645
rect 30193 11679 30251 11685
rect 30193 11645 30205 11679
rect 30239 11645 30251 11679
rect 30558 11676 30564 11688
rect 30519 11648 30564 11676
rect 30193 11639 30251 11645
rect 30208 11608 30236 11639
rect 30558 11636 30564 11648
rect 30616 11676 30622 11688
rect 30760 11676 30788 11716
rect 34054 11704 34060 11716
rect 34112 11704 34118 11756
rect 34238 11744 34244 11756
rect 34199 11716 34244 11744
rect 34238 11704 34244 11716
rect 34296 11704 34302 11756
rect 35250 11704 35256 11756
rect 35308 11744 35314 11756
rect 35710 11744 35716 11756
rect 35308 11716 35716 11744
rect 35308 11704 35314 11716
rect 35710 11704 35716 11716
rect 35768 11744 35774 11756
rect 35768 11716 36032 11744
rect 35768 11704 35774 11716
rect 30616 11648 30788 11676
rect 31297 11679 31355 11685
rect 30616 11636 30622 11648
rect 31297 11645 31309 11679
rect 31343 11676 31355 11679
rect 31478 11676 31484 11688
rect 31343 11648 31484 11676
rect 31343 11645 31355 11648
rect 31297 11639 31355 11645
rect 31478 11636 31484 11648
rect 31536 11636 31542 11688
rect 32306 11676 32312 11688
rect 32267 11648 32312 11676
rect 32306 11636 32312 11648
rect 32364 11636 32370 11688
rect 32766 11676 32772 11688
rect 32727 11648 32772 11676
rect 32766 11636 32772 11648
rect 32824 11636 32830 11688
rect 33410 11676 33416 11688
rect 33323 11648 33416 11676
rect 33410 11636 33416 11648
rect 33468 11676 33474 11688
rect 33686 11676 33692 11688
rect 33468 11648 33692 11676
rect 33468 11636 33474 11648
rect 33686 11636 33692 11648
rect 33744 11636 33750 11688
rect 33965 11679 34023 11685
rect 33965 11645 33977 11679
rect 34011 11676 34023 11679
rect 34790 11676 34796 11688
rect 34011 11648 34796 11676
rect 34011 11645 34023 11648
rect 33965 11639 34023 11645
rect 34790 11636 34796 11648
rect 34848 11636 34854 11688
rect 36004 11685 36032 11716
rect 37182 11704 37188 11756
rect 37240 11744 37246 11756
rect 37461 11747 37519 11753
rect 37461 11744 37473 11747
rect 37240 11716 37473 11744
rect 37240 11704 37246 11716
rect 37461 11713 37473 11716
rect 37507 11713 37519 11747
rect 37461 11707 37519 11713
rect 37737 11747 37795 11753
rect 37737 11713 37749 11747
rect 37783 11744 37795 11747
rect 37918 11744 37924 11756
rect 37783 11716 37924 11744
rect 37783 11713 37795 11716
rect 37737 11707 37795 11713
rect 37918 11704 37924 11716
rect 37976 11704 37982 11756
rect 35805 11679 35863 11685
rect 35805 11645 35817 11679
rect 35851 11645 35863 11679
rect 35805 11639 35863 11645
rect 35989 11679 36047 11685
rect 35989 11645 36001 11679
rect 36035 11645 36047 11679
rect 36170 11676 36176 11688
rect 36131 11648 36176 11676
rect 35989 11639 36047 11645
rect 30116 11580 30236 11608
rect 22060 11512 25452 11540
rect 22060 11500 22066 11512
rect 25498 11500 25504 11552
rect 25556 11540 25562 11552
rect 30116 11540 30144 11580
rect 32398 11568 32404 11620
rect 32456 11608 32462 11620
rect 35820 11608 35848 11639
rect 36170 11636 36176 11648
rect 36228 11636 36234 11688
rect 32456 11580 35848 11608
rect 32456 11568 32462 11580
rect 30834 11540 30840 11552
rect 25556 11512 30840 11540
rect 25556 11500 25562 11512
rect 30834 11500 30840 11512
rect 30892 11500 30898 11552
rect 37826 11500 37832 11552
rect 37884 11540 37890 11552
rect 38841 11543 38899 11549
rect 38841 11540 38853 11543
rect 37884 11512 38853 11540
rect 37884 11500 37890 11512
rect 38841 11509 38853 11512
rect 38887 11509 38899 11543
rect 38841 11503 38899 11509
rect 1104 11450 39836 11472
rect 1104 11398 19606 11450
rect 19658 11398 19670 11450
rect 19722 11398 19734 11450
rect 19786 11398 19798 11450
rect 19850 11398 39836 11450
rect 1104 11376 39836 11398
rect 7834 11336 7840 11348
rect 7795 11308 7840 11336
rect 7834 11296 7840 11308
rect 7892 11296 7898 11348
rect 11057 11339 11115 11345
rect 11057 11305 11069 11339
rect 11103 11336 11115 11339
rect 12710 11336 12716 11348
rect 11103 11308 12716 11336
rect 11103 11305 11115 11308
rect 11057 11299 11115 11305
rect 12710 11296 12716 11308
rect 12768 11336 12774 11348
rect 13354 11336 13360 11348
rect 12768 11308 13360 11336
rect 12768 11296 12774 11308
rect 13354 11296 13360 11308
rect 13412 11296 13418 11348
rect 14366 11336 14372 11348
rect 14327 11308 14372 11336
rect 14366 11296 14372 11308
rect 14424 11296 14430 11348
rect 14476 11308 16252 11336
rect 7006 11268 7012 11280
rect 6656 11240 7012 11268
rect 1670 11160 1676 11212
rect 1728 11200 1734 11212
rect 1949 11203 2007 11209
rect 1949 11200 1961 11203
rect 1728 11172 1961 11200
rect 1728 11160 1734 11172
rect 1949 11169 1961 11172
rect 1995 11169 2007 11203
rect 1949 11163 2007 11169
rect 2774 11160 2780 11212
rect 2832 11200 2838 11212
rect 2958 11200 2964 11212
rect 2832 11172 2877 11200
rect 2919 11172 2964 11200
rect 2832 11160 2838 11172
rect 2958 11160 2964 11172
rect 3016 11160 3022 11212
rect 5445 11203 5503 11209
rect 5445 11169 5457 11203
rect 5491 11200 5503 11203
rect 5534 11200 5540 11212
rect 5491 11172 5540 11200
rect 5491 11169 5503 11172
rect 5445 11163 5503 11169
rect 5534 11160 5540 11172
rect 5592 11160 5598 11212
rect 5718 11160 5724 11212
rect 5776 11200 5782 11212
rect 5905 11203 5963 11209
rect 5905 11200 5917 11203
rect 5776 11172 5917 11200
rect 5776 11160 5782 11172
rect 5905 11169 5917 11172
rect 5951 11169 5963 11203
rect 5905 11163 5963 11169
rect 6273 11203 6331 11209
rect 6273 11169 6285 11203
rect 6319 11200 6331 11203
rect 6362 11200 6368 11212
rect 6319 11172 6368 11200
rect 6319 11169 6331 11172
rect 6273 11163 6331 11169
rect 5920 11132 5948 11163
rect 6362 11160 6368 11172
rect 6420 11160 6426 11212
rect 6656 11209 6684 11240
rect 7006 11228 7012 11240
rect 7064 11228 7070 11280
rect 10413 11271 10471 11277
rect 7300 11240 10180 11268
rect 6641 11203 6699 11209
rect 6641 11169 6653 11203
rect 6687 11169 6699 11203
rect 7190 11200 7196 11212
rect 7151 11172 7196 11200
rect 6641 11163 6699 11169
rect 7190 11160 7196 11172
rect 7248 11160 7254 11212
rect 5994 11132 6000 11144
rect 5907 11104 6000 11132
rect 5994 11092 6000 11104
rect 6052 11132 6058 11144
rect 7300 11132 7328 11240
rect 7745 11203 7803 11209
rect 7745 11169 7757 11203
rect 7791 11169 7803 11203
rect 8386 11200 8392 11212
rect 8347 11172 8392 11200
rect 7745 11163 7803 11169
rect 6052 11104 7328 11132
rect 6052 11092 6058 11104
rect 2590 11024 2596 11076
rect 2648 11064 2654 11076
rect 2685 11067 2743 11073
rect 2685 11064 2697 11067
rect 2648 11036 2697 11064
rect 2648 11024 2654 11036
rect 2685 11033 2697 11036
rect 2731 11033 2743 11067
rect 5534 11064 5540 11076
rect 5495 11036 5540 11064
rect 2685 11027 2743 11033
rect 5534 11024 5540 11036
rect 5592 11024 5598 11076
rect 7760 11064 7788 11163
rect 8386 11160 8392 11172
rect 8444 11160 8450 11212
rect 8478 11160 8484 11212
rect 8536 11200 8542 11212
rect 8849 11203 8907 11209
rect 8849 11200 8861 11203
rect 8536 11172 8861 11200
rect 8536 11160 8542 11172
rect 8849 11169 8861 11172
rect 8895 11169 8907 11203
rect 9674 11200 9680 11212
rect 9635 11172 9680 11200
rect 8849 11163 8907 11169
rect 9674 11160 9680 11172
rect 9732 11160 9738 11212
rect 10152 11209 10180 11240
rect 10413 11237 10425 11271
rect 10459 11268 10471 11271
rect 10459 11240 12020 11268
rect 10459 11237 10471 11240
rect 10413 11231 10471 11237
rect 10137 11203 10195 11209
rect 10137 11169 10149 11203
rect 10183 11169 10195 11203
rect 11238 11200 11244 11212
rect 11199 11172 11244 11200
rect 10137 11163 10195 11169
rect 11238 11160 11244 11172
rect 11296 11160 11302 11212
rect 11992 11209 12020 11240
rect 12066 11228 12072 11280
rect 12124 11268 12130 11280
rect 14476 11268 14504 11308
rect 12124 11240 14504 11268
rect 16224 11268 16252 11308
rect 16298 11296 16304 11348
rect 16356 11336 16362 11348
rect 16669 11339 16727 11345
rect 16669 11336 16681 11339
rect 16356 11308 16681 11336
rect 16356 11296 16362 11308
rect 16669 11305 16681 11308
rect 16715 11305 16727 11339
rect 16669 11299 16727 11305
rect 18230 11296 18236 11348
rect 18288 11296 18294 11348
rect 19058 11296 19064 11348
rect 19116 11336 19122 11348
rect 19153 11339 19211 11345
rect 19153 11336 19165 11339
rect 19116 11308 19165 11336
rect 19116 11296 19122 11308
rect 19153 11305 19165 11308
rect 19199 11305 19211 11339
rect 19153 11299 19211 11305
rect 20070 11296 20076 11348
rect 20128 11336 20134 11348
rect 21085 11339 21143 11345
rect 20128 11308 20208 11336
rect 20128 11296 20134 11308
rect 18248 11268 18276 11296
rect 16224 11240 18276 11268
rect 12124 11228 12130 11240
rect 11977 11203 12035 11209
rect 11977 11169 11989 11203
rect 12023 11169 12035 11203
rect 12342 11200 12348 11212
rect 12303 11172 12348 11200
rect 11977 11163 12035 11169
rect 12342 11160 12348 11172
rect 12400 11160 12406 11212
rect 12452 11209 12480 11240
rect 18322 11228 18328 11280
rect 18380 11268 18386 11280
rect 20180 11268 20208 11308
rect 21085 11305 21097 11339
rect 21131 11336 21143 11339
rect 21450 11336 21456 11348
rect 21131 11308 21456 11336
rect 21131 11305 21143 11308
rect 21085 11299 21143 11305
rect 21450 11296 21456 11308
rect 21508 11296 21514 11348
rect 21542 11296 21548 11348
rect 21600 11336 21606 11348
rect 25130 11336 25136 11348
rect 21600 11308 25136 11336
rect 21600 11296 21606 11308
rect 25130 11296 25136 11308
rect 25188 11296 25194 11348
rect 25225 11339 25283 11345
rect 25225 11305 25237 11339
rect 25271 11336 25283 11339
rect 27982 11336 27988 11348
rect 25271 11308 27988 11336
rect 25271 11305 25283 11308
rect 25225 11299 25283 11305
rect 23198 11268 23204 11280
rect 18380 11240 19104 11268
rect 20180 11240 22140 11268
rect 18380 11228 18386 11240
rect 19076 11212 19104 11240
rect 12437 11203 12495 11209
rect 12437 11169 12449 11203
rect 12483 11169 12495 11203
rect 12437 11163 12495 11169
rect 12526 11160 12532 11212
rect 12584 11200 12590 11212
rect 12989 11203 13047 11209
rect 12989 11200 13001 11203
rect 12584 11172 13001 11200
rect 12584 11160 12590 11172
rect 12989 11169 13001 11172
rect 13035 11169 13047 11203
rect 13538 11200 13544 11212
rect 13499 11172 13544 11200
rect 12989 11163 13047 11169
rect 13538 11160 13544 11172
rect 13596 11160 13602 11212
rect 14182 11200 14188 11212
rect 14143 11172 14188 11200
rect 14182 11160 14188 11172
rect 14240 11160 14246 11212
rect 15102 11160 15108 11212
rect 15160 11200 15166 11212
rect 15565 11203 15623 11209
rect 15565 11200 15577 11203
rect 15160 11172 15577 11200
rect 15160 11160 15166 11172
rect 15565 11169 15577 11172
rect 15611 11169 15623 11203
rect 17954 11200 17960 11212
rect 17915 11172 17960 11200
rect 15565 11163 15623 11169
rect 17954 11160 17960 11172
rect 18012 11160 18018 11212
rect 18417 11203 18475 11209
rect 18417 11169 18429 11203
rect 18463 11200 18475 11203
rect 18782 11200 18788 11212
rect 18463 11172 18788 11200
rect 18463 11169 18475 11172
rect 18417 11163 18475 11169
rect 18782 11160 18788 11172
rect 18840 11160 18846 11212
rect 19058 11200 19064 11212
rect 19019 11172 19064 11200
rect 19058 11160 19064 11172
rect 19116 11160 19122 11212
rect 19429 11203 19487 11209
rect 19429 11169 19441 11203
rect 19475 11200 19487 11203
rect 19794 11200 19800 11212
rect 19475 11172 19800 11200
rect 19475 11169 19487 11172
rect 19429 11163 19487 11169
rect 19794 11160 19800 11172
rect 19852 11160 19858 11212
rect 20070 11200 20076 11212
rect 20031 11172 20076 11200
rect 20070 11160 20076 11172
rect 20128 11160 20134 11212
rect 20990 11200 20996 11212
rect 20272 11172 20996 11200
rect 9125 11135 9183 11141
rect 9125 11101 9137 11135
rect 9171 11132 9183 11135
rect 10870 11132 10876 11144
rect 9171 11104 10876 11132
rect 9171 11101 9183 11104
rect 9125 11095 9183 11101
rect 10870 11092 10876 11104
rect 10928 11092 10934 11144
rect 11885 11135 11943 11141
rect 11885 11132 11897 11135
rect 11256 11104 11897 11132
rect 7760 11036 10088 11064
rect 10060 10996 10088 11036
rect 10134 11024 10140 11076
rect 10192 11064 10198 11076
rect 11256 11064 11284 11104
rect 11885 11101 11897 11104
rect 11931 11101 11943 11135
rect 11885 11095 11943 11101
rect 13357 11135 13415 11141
rect 13357 11101 13369 11135
rect 13403 11132 13415 11135
rect 13630 11132 13636 11144
rect 13403 11104 13636 11132
rect 13403 11101 13415 11104
rect 13357 11095 13415 11101
rect 11422 11064 11428 11076
rect 10192 11036 11284 11064
rect 11383 11036 11428 11064
rect 10192 11024 10198 11036
rect 11422 11024 11428 11036
rect 11480 11024 11486 11076
rect 11900 11064 11928 11095
rect 13630 11092 13636 11104
rect 13688 11092 13694 11144
rect 15289 11135 15347 11141
rect 15289 11101 15301 11135
rect 15335 11132 15347 11135
rect 16206 11132 16212 11144
rect 15335 11104 16212 11132
rect 15335 11101 15347 11104
rect 15289 11095 15347 11101
rect 16206 11092 16212 11104
rect 16264 11092 16270 11144
rect 11974 11064 11980 11076
rect 11900 11036 11980 11064
rect 11974 11024 11980 11036
rect 12032 11024 12038 11076
rect 17770 11064 17776 11076
rect 17731 11036 17776 11064
rect 17770 11024 17776 11036
rect 17828 11024 17834 11076
rect 19978 11024 19984 11076
rect 20036 11064 20042 11076
rect 20272 11073 20300 11172
rect 20990 11160 20996 11172
rect 21048 11160 21054 11212
rect 21545 11203 21603 11209
rect 21545 11169 21557 11203
rect 21591 11169 21603 11203
rect 21545 11163 21603 11169
rect 21560 11132 21588 11163
rect 21910 11132 21916 11144
rect 21560 11104 21916 11132
rect 21910 11092 21916 11104
rect 21968 11092 21974 11144
rect 22005 11135 22063 11141
rect 22005 11101 22017 11135
rect 22051 11101 22063 11135
rect 22112 11132 22140 11240
rect 22572 11240 23204 11268
rect 22186 11160 22192 11212
rect 22244 11200 22250 11212
rect 22572 11209 22600 11240
rect 23198 11228 23204 11240
rect 23256 11228 23262 11280
rect 25240 11268 25268 11299
rect 27982 11296 27988 11308
rect 28040 11296 28046 11348
rect 30558 11296 30564 11348
rect 30616 11296 30622 11348
rect 32306 11296 32312 11348
rect 32364 11336 32370 11348
rect 33594 11336 33600 11348
rect 32364 11308 33600 11336
rect 32364 11296 32370 11308
rect 33594 11296 33600 11308
rect 33652 11296 33658 11348
rect 35802 11336 35808 11348
rect 34532 11308 35808 11336
rect 24228 11240 25268 11268
rect 25869 11271 25927 11277
rect 22557 11203 22615 11209
rect 22557 11200 22569 11203
rect 22244 11172 22569 11200
rect 22244 11160 22250 11172
rect 22557 11169 22569 11172
rect 22603 11169 22615 11203
rect 22557 11163 22615 11169
rect 23014 11160 23020 11212
rect 23072 11200 23078 11212
rect 23477 11203 23535 11209
rect 23477 11200 23489 11203
rect 23072 11172 23489 11200
rect 23072 11160 23078 11172
rect 23477 11169 23489 11172
rect 23523 11169 23535 11203
rect 23477 11163 23535 11169
rect 23842 11160 23848 11212
rect 23900 11200 23906 11212
rect 24228 11209 24256 11240
rect 25869 11237 25881 11271
rect 25915 11268 25927 11271
rect 27249 11271 27307 11277
rect 25915 11240 27200 11268
rect 25915 11237 25927 11240
rect 25869 11231 25927 11237
rect 24029 11203 24087 11209
rect 24029 11200 24041 11203
rect 23900 11172 24041 11200
rect 23900 11160 23906 11172
rect 24029 11169 24041 11172
rect 24075 11169 24087 11203
rect 24029 11163 24087 11169
rect 24213 11203 24271 11209
rect 24213 11169 24225 11203
rect 24259 11169 24271 11203
rect 25130 11200 25136 11212
rect 25091 11172 25136 11200
rect 24213 11163 24271 11169
rect 25130 11160 25136 11172
rect 25188 11200 25194 11212
rect 25682 11200 25688 11212
rect 25188 11172 25688 11200
rect 25188 11160 25194 11172
rect 25682 11160 25688 11172
rect 25740 11160 25746 11212
rect 25777 11203 25835 11209
rect 25777 11169 25789 11203
rect 25823 11169 25835 11203
rect 25777 11163 25835 11169
rect 22649 11135 22707 11141
rect 22649 11132 22661 11135
rect 22112 11104 22661 11132
rect 22005 11095 22063 11101
rect 22649 11101 22661 11104
rect 22695 11101 22707 11135
rect 23290 11132 23296 11144
rect 23251 11104 23296 11132
rect 22649 11095 22707 11101
rect 20257 11067 20315 11073
rect 20257 11064 20269 11067
rect 20036 11036 20269 11064
rect 20036 11024 20042 11036
rect 20257 11033 20269 11036
rect 20303 11033 20315 11067
rect 22020 11064 22048 11095
rect 23290 11092 23296 11104
rect 23348 11092 23354 11144
rect 25792 11132 25820 11163
rect 26418 11160 26424 11212
rect 26476 11200 26482 11212
rect 26513 11203 26571 11209
rect 26513 11200 26525 11203
rect 26476 11172 26525 11200
rect 26476 11160 26482 11172
rect 26513 11169 26525 11172
rect 26559 11169 26571 11203
rect 26513 11163 26571 11169
rect 26602 11160 26608 11212
rect 26660 11200 26666 11212
rect 26973 11203 27031 11209
rect 26973 11200 26985 11203
rect 26660 11172 26985 11200
rect 26660 11160 26666 11172
rect 26973 11169 26985 11172
rect 27019 11169 27031 11203
rect 26973 11163 27031 11169
rect 27172 11132 27200 11240
rect 27249 11237 27261 11271
rect 27295 11268 27307 11271
rect 27706 11268 27712 11280
rect 27295 11240 27712 11268
rect 27295 11237 27307 11240
rect 27249 11231 27307 11237
rect 27706 11228 27712 11240
rect 27764 11228 27770 11280
rect 30576 11268 30604 11296
rect 28092 11240 28948 11268
rect 30576 11240 31064 11268
rect 27338 11160 27344 11212
rect 27396 11200 27402 11212
rect 28092 11200 28120 11240
rect 28920 11209 28948 11240
rect 27396 11172 28120 11200
rect 28169 11203 28227 11209
rect 27396 11160 27402 11172
rect 28169 11169 28181 11203
rect 28215 11200 28227 11203
rect 28905 11203 28963 11209
rect 28215 11172 28856 11200
rect 28215 11169 28227 11172
rect 28169 11163 28227 11169
rect 28258 11132 28264 11144
rect 25792 11104 27016 11132
rect 27172 11104 28264 11132
rect 26988 11076 27016 11104
rect 28258 11092 28264 11104
rect 28316 11132 28322 11144
rect 28721 11135 28779 11141
rect 28721 11132 28733 11135
rect 28316 11104 28733 11132
rect 28316 11092 28322 11104
rect 28721 11101 28733 11104
rect 28767 11101 28779 11135
rect 28828 11132 28856 11172
rect 28905 11169 28917 11203
rect 28951 11169 28963 11203
rect 29270 11200 29276 11212
rect 29231 11172 29276 11200
rect 28905 11163 28963 11169
rect 29270 11160 29276 11172
rect 29328 11160 29334 11212
rect 29457 11203 29515 11209
rect 29457 11169 29469 11203
rect 29503 11200 29515 11203
rect 29822 11200 29828 11212
rect 29503 11172 29828 11200
rect 29503 11169 29515 11172
rect 29457 11163 29515 11169
rect 29822 11160 29828 11172
rect 29880 11160 29886 11212
rect 30558 11200 30564 11212
rect 30519 11172 30564 11200
rect 30558 11160 30564 11172
rect 30616 11160 30622 11212
rect 30834 11160 30840 11212
rect 30892 11200 30898 11212
rect 31036 11209 31064 11240
rect 32950 11228 32956 11280
rect 33008 11268 33014 11280
rect 34532 11268 34560 11308
rect 35802 11296 35808 11308
rect 35860 11296 35866 11348
rect 36078 11296 36084 11348
rect 36136 11336 36142 11348
rect 36909 11339 36967 11345
rect 36909 11336 36921 11339
rect 36136 11308 36921 11336
rect 36136 11296 36142 11308
rect 36909 11305 36921 11308
rect 36955 11305 36967 11339
rect 36909 11299 36967 11305
rect 38654 11296 38660 11348
rect 38712 11336 38718 11348
rect 38841 11339 38899 11345
rect 38841 11336 38853 11339
rect 38712 11308 38853 11336
rect 38712 11296 38718 11308
rect 38841 11305 38853 11308
rect 38887 11305 38899 11339
rect 38841 11299 38899 11305
rect 38289 11271 38347 11277
rect 38289 11268 38301 11271
rect 33008 11240 34560 11268
rect 36832 11240 38301 11268
rect 33008 11228 33014 11240
rect 30929 11203 30987 11209
rect 30929 11200 30941 11203
rect 30892 11172 30941 11200
rect 30892 11160 30898 11172
rect 30929 11169 30941 11172
rect 30975 11169 30987 11203
rect 30929 11163 30987 11169
rect 31021 11203 31079 11209
rect 31021 11169 31033 11203
rect 31067 11169 31079 11203
rect 32122 11200 32128 11212
rect 32083 11172 32128 11200
rect 31021 11163 31079 11169
rect 32122 11160 32128 11172
rect 32180 11160 32186 11212
rect 32306 11160 32312 11212
rect 32364 11200 32370 11212
rect 32493 11203 32551 11209
rect 32493 11200 32505 11203
rect 32364 11172 32505 11200
rect 32364 11160 32370 11172
rect 32493 11169 32505 11172
rect 32539 11200 32551 11203
rect 32582 11200 32588 11212
rect 32539 11172 32588 11200
rect 32539 11169 32551 11172
rect 32493 11163 32551 11169
rect 32582 11160 32588 11172
rect 32640 11160 32646 11212
rect 33042 11200 33048 11212
rect 33003 11172 33048 11200
rect 33042 11160 33048 11172
rect 33100 11160 33106 11212
rect 33686 11200 33692 11212
rect 33647 11172 33692 11200
rect 33686 11160 33692 11172
rect 33744 11160 33750 11212
rect 33778 11160 33784 11212
rect 33836 11200 33842 11212
rect 34241 11203 34299 11209
rect 34241 11200 34253 11203
rect 33836 11172 34253 11200
rect 33836 11160 33842 11172
rect 34241 11169 34253 11172
rect 34287 11169 34299 11203
rect 34241 11163 34299 11169
rect 35805 11203 35863 11209
rect 35805 11169 35817 11203
rect 35851 11200 35863 11203
rect 36832 11200 36860 11240
rect 38289 11237 38301 11240
rect 38335 11237 38347 11271
rect 38289 11231 38347 11237
rect 37826 11200 37832 11212
rect 35851 11172 36860 11200
rect 37787 11172 37832 11200
rect 35851 11169 35863 11172
rect 35805 11163 35863 11169
rect 37826 11160 37832 11172
rect 37884 11160 37890 11212
rect 37918 11160 37924 11212
rect 37976 11200 37982 11212
rect 38749 11203 38807 11209
rect 38749 11200 38761 11203
rect 37976 11172 38761 11200
rect 37976 11160 37982 11172
rect 38749 11169 38761 11172
rect 38795 11169 38807 11203
rect 38749 11163 38807 11169
rect 28828 11104 29776 11132
rect 28721 11095 28779 11101
rect 22554 11064 22560 11076
rect 22020 11036 22560 11064
rect 20257 11027 20315 11033
rect 22554 11024 22560 11036
rect 22612 11024 22618 11076
rect 26970 11024 26976 11076
rect 27028 11024 27034 11076
rect 27985 11067 28043 11073
rect 27985 11033 27997 11067
rect 28031 11033 28043 11067
rect 27985 11027 28043 11033
rect 28537 11067 28595 11073
rect 28537 11033 28549 11067
rect 28583 11064 28595 11067
rect 28994 11064 29000 11076
rect 28583 11036 29000 11064
rect 28583 11033 28595 11036
rect 28537 11027 28595 11033
rect 10502 10996 10508 11008
rect 10060 10968 10508 10996
rect 10502 10956 10508 10968
rect 10560 10956 10566 11008
rect 18046 10956 18052 11008
rect 18104 10996 18110 11008
rect 20714 10996 20720 11008
rect 18104 10968 20720 10996
rect 18104 10956 18110 10968
rect 20714 10956 20720 10968
rect 20772 10996 20778 11008
rect 21266 10996 21272 11008
rect 20772 10968 21272 10996
rect 20772 10956 20778 10968
rect 21266 10956 21272 10968
rect 21324 10956 21330 11008
rect 24486 10996 24492 11008
rect 24447 10968 24492 10996
rect 24486 10956 24492 10968
rect 24544 10956 24550 11008
rect 28000 10996 28028 11027
rect 28994 11024 29000 11036
rect 29052 11024 29058 11076
rect 29748 11064 29776 11104
rect 30282 11092 30288 11144
rect 30340 11132 30346 11144
rect 30653 11135 30711 11141
rect 30653 11132 30665 11135
rect 30340 11104 30665 11132
rect 30340 11092 30346 11104
rect 30653 11101 30665 11104
rect 30699 11132 30711 11135
rect 31478 11132 31484 11144
rect 30699 11104 31484 11132
rect 30699 11101 30711 11104
rect 30653 11095 30711 11101
rect 31478 11092 31484 11104
rect 31536 11092 31542 11144
rect 32766 11092 32772 11144
rect 32824 11132 32830 11144
rect 32953 11135 33011 11141
rect 32953 11132 32965 11135
rect 32824 11104 32965 11132
rect 32824 11092 32830 11104
rect 32953 11101 32965 11104
rect 32999 11101 33011 11135
rect 34517 11135 34575 11141
rect 34517 11132 34529 11135
rect 32953 11095 33011 11101
rect 33060 11104 34529 11132
rect 30834 11064 30840 11076
rect 29748 11036 30840 11064
rect 30834 11024 30840 11036
rect 30892 11024 30898 11076
rect 32582 11024 32588 11076
rect 32640 11064 32646 11076
rect 33060 11064 33088 11104
rect 34517 11101 34529 11104
rect 34563 11101 34575 11135
rect 34517 11095 34575 11101
rect 34606 11092 34612 11144
rect 34664 11132 34670 11144
rect 35529 11135 35587 11141
rect 35529 11132 35541 11135
rect 34664 11104 35541 11132
rect 34664 11092 34670 11104
rect 35529 11101 35541 11104
rect 35575 11132 35587 11135
rect 36170 11132 36176 11144
rect 35575 11104 36176 11132
rect 35575 11101 35587 11104
rect 35529 11095 35587 11101
rect 36170 11092 36176 11104
rect 36228 11092 36234 11144
rect 37737 11135 37795 11141
rect 37737 11101 37749 11135
rect 37783 11101 37795 11135
rect 37737 11095 37795 11101
rect 33962 11064 33968 11076
rect 32640 11036 33088 11064
rect 33923 11036 33968 11064
rect 32640 11024 32646 11036
rect 33962 11024 33968 11036
rect 34020 11024 34026 11076
rect 28902 10996 28908 11008
rect 28000 10968 28908 10996
rect 28902 10956 28908 10968
rect 28960 10956 28966 11008
rect 29086 10956 29092 11008
rect 29144 10996 29150 11008
rect 30193 10999 30251 11005
rect 30193 10996 30205 10999
rect 29144 10968 30205 10996
rect 29144 10956 29150 10968
rect 30193 10965 30205 10968
rect 30239 10965 30251 10999
rect 30193 10959 30251 10965
rect 33134 10956 33140 11008
rect 33192 10996 33198 11008
rect 34330 10996 34336 11008
rect 33192 10968 34336 10996
rect 33192 10956 33198 10968
rect 34330 10956 34336 10968
rect 34388 10996 34394 11008
rect 34624 10996 34652 11092
rect 37752 11064 37780 11095
rect 36464 11036 37780 11064
rect 34388 10968 34652 10996
rect 34388 10956 34394 10968
rect 35802 10956 35808 11008
rect 35860 10996 35866 11008
rect 36464 10996 36492 11036
rect 35860 10968 36492 10996
rect 35860 10956 35866 10968
rect 1104 10906 39836 10928
rect 1104 10854 4246 10906
rect 4298 10854 4310 10906
rect 4362 10854 4374 10906
rect 4426 10854 4438 10906
rect 4490 10854 34966 10906
rect 35018 10854 35030 10906
rect 35082 10854 35094 10906
rect 35146 10854 35158 10906
rect 35210 10854 39836 10906
rect 1104 10832 39836 10854
rect 2682 10752 2688 10804
rect 2740 10792 2746 10804
rect 2777 10795 2835 10801
rect 2777 10792 2789 10795
rect 2740 10764 2789 10792
rect 2740 10752 2746 10764
rect 2777 10761 2789 10764
rect 2823 10761 2835 10795
rect 4890 10792 4896 10804
rect 4851 10764 4896 10792
rect 2777 10755 2835 10761
rect 4890 10752 4896 10764
rect 4948 10752 4954 10804
rect 5994 10792 6000 10804
rect 5955 10764 6000 10792
rect 5994 10752 6000 10764
rect 6052 10752 6058 10804
rect 16758 10792 16764 10804
rect 11072 10764 16436 10792
rect 16719 10764 16764 10792
rect 4614 10616 4620 10668
rect 4672 10656 4678 10668
rect 6825 10659 6883 10665
rect 6825 10656 6837 10659
rect 4672 10628 6837 10656
rect 4672 10616 4678 10628
rect 6825 10625 6837 10628
rect 6871 10625 6883 10659
rect 6825 10619 6883 10625
rect 9677 10659 9735 10665
rect 9677 10625 9689 10659
rect 9723 10656 9735 10659
rect 11072 10656 11100 10764
rect 11149 10727 11207 10733
rect 11149 10693 11161 10727
rect 11195 10693 11207 10727
rect 11149 10687 11207 10693
rect 9723 10628 11100 10656
rect 11164 10656 11192 10687
rect 11514 10684 11520 10736
rect 11572 10724 11578 10736
rect 12529 10727 12587 10733
rect 12529 10724 12541 10727
rect 11572 10696 12541 10724
rect 11572 10684 11578 10696
rect 12529 10693 12541 10696
rect 12575 10693 12587 10727
rect 16408 10724 16436 10764
rect 16758 10752 16764 10764
rect 16816 10752 16822 10804
rect 17126 10752 17132 10804
rect 17184 10792 17190 10804
rect 20806 10792 20812 10804
rect 17184 10764 20812 10792
rect 17184 10752 17190 10764
rect 20806 10752 20812 10764
rect 20864 10752 20870 10804
rect 26234 10792 26240 10804
rect 20916 10764 26240 10792
rect 17218 10724 17224 10736
rect 12529 10687 12587 10693
rect 13096 10696 16160 10724
rect 16408 10696 17224 10724
rect 13096 10656 13124 10696
rect 11164 10628 13124 10656
rect 9723 10625 9735 10628
rect 9677 10619 9735 10625
rect 13170 10616 13176 10668
rect 13228 10656 13234 10668
rect 13909 10659 13967 10665
rect 13909 10656 13921 10659
rect 13228 10628 13921 10656
rect 13228 10616 13234 10628
rect 13909 10625 13921 10628
rect 13955 10625 13967 10659
rect 15562 10656 15568 10668
rect 13909 10619 13967 10625
rect 14844 10628 15568 10656
rect 1394 10588 1400 10600
rect 1355 10560 1400 10588
rect 1394 10548 1400 10560
rect 1452 10548 1458 10600
rect 1670 10588 1676 10600
rect 1631 10560 1676 10588
rect 1670 10548 1676 10560
rect 1728 10548 1734 10600
rect 3510 10588 3516 10600
rect 3471 10560 3516 10588
rect 3510 10548 3516 10560
rect 3568 10548 3574 10600
rect 3786 10588 3792 10600
rect 3747 10560 3792 10588
rect 3786 10548 3792 10560
rect 3844 10548 3850 10600
rect 5902 10588 5908 10600
rect 5863 10560 5908 10588
rect 5902 10548 5908 10560
rect 5960 10548 5966 10600
rect 7098 10588 7104 10600
rect 7059 10560 7104 10588
rect 7098 10548 7104 10560
rect 7156 10548 7162 10600
rect 9306 10588 9312 10600
rect 9267 10560 9312 10588
rect 9306 10548 9312 10560
rect 9364 10548 9370 10600
rect 9858 10588 9864 10600
rect 9819 10560 9864 10588
rect 9858 10548 9864 10560
rect 9916 10548 9922 10600
rect 11238 10548 11244 10600
rect 11296 10588 11302 10600
rect 11333 10591 11391 10597
rect 11333 10588 11345 10591
rect 11296 10560 11345 10588
rect 11296 10548 11302 10560
rect 11333 10557 11345 10560
rect 11379 10557 11391 10591
rect 11514 10588 11520 10600
rect 11475 10560 11520 10588
rect 11333 10551 11391 10557
rect 11514 10548 11520 10560
rect 11572 10548 11578 10600
rect 11698 10588 11704 10600
rect 11659 10560 11704 10588
rect 11698 10548 11704 10560
rect 11756 10548 11762 10600
rect 11882 10548 11888 10600
rect 11940 10588 11946 10600
rect 12437 10591 12495 10597
rect 12437 10588 12449 10591
rect 11940 10560 12449 10588
rect 11940 10548 11946 10560
rect 12437 10557 12449 10560
rect 12483 10557 12495 10591
rect 12437 10551 12495 10557
rect 12989 10591 13047 10597
rect 12989 10557 13001 10591
rect 13035 10557 13047 10591
rect 13998 10588 14004 10600
rect 13959 10560 14004 10588
rect 12989 10551 13047 10557
rect 8481 10523 8539 10529
rect 8481 10489 8493 10523
rect 8527 10520 8539 10523
rect 8938 10520 8944 10532
rect 8527 10492 8944 10520
rect 8527 10489 8539 10492
rect 8481 10483 8539 10489
rect 8938 10480 8944 10492
rect 8996 10480 9002 10532
rect 10594 10480 10600 10532
rect 10652 10520 10658 10532
rect 13004 10520 13032 10551
rect 13998 10548 14004 10560
rect 14056 10548 14062 10600
rect 14844 10597 14872 10628
rect 15562 10616 15568 10628
rect 15620 10616 15626 10668
rect 16022 10656 16028 10668
rect 15764 10628 16028 10656
rect 14277 10591 14335 10597
rect 14277 10557 14289 10591
rect 14323 10557 14335 10591
rect 14277 10551 14335 10557
rect 14829 10591 14887 10597
rect 14829 10557 14841 10591
rect 14875 10557 14887 10591
rect 14829 10551 14887 10557
rect 15105 10591 15163 10597
rect 15105 10557 15117 10591
rect 15151 10588 15163 10591
rect 15286 10588 15292 10600
rect 15151 10560 15292 10588
rect 15151 10557 15163 10560
rect 15105 10551 15163 10557
rect 10652 10492 13032 10520
rect 10652 10480 10658 10492
rect 8846 10412 8852 10464
rect 8904 10452 8910 10464
rect 14292 10452 14320 10551
rect 15286 10548 15292 10560
rect 15344 10548 15350 10600
rect 15764 10597 15792 10628
rect 16022 10616 16028 10628
rect 16080 10616 16086 10668
rect 15749 10591 15807 10597
rect 15749 10557 15761 10591
rect 15795 10557 15807 10591
rect 15749 10551 15807 10557
rect 16132 10520 16160 10696
rect 17218 10684 17224 10696
rect 17276 10684 17282 10736
rect 19245 10727 19303 10733
rect 19245 10693 19257 10727
rect 19291 10724 19303 10727
rect 20916 10724 20944 10764
rect 26234 10752 26240 10764
rect 26292 10752 26298 10804
rect 26418 10752 26424 10804
rect 26476 10792 26482 10804
rect 27154 10792 27160 10804
rect 26476 10764 27160 10792
rect 26476 10752 26482 10764
rect 27154 10752 27160 10764
rect 27212 10752 27218 10804
rect 31478 10752 31484 10804
rect 31536 10792 31542 10804
rect 33318 10792 33324 10804
rect 31536 10764 33324 10792
rect 31536 10752 31542 10764
rect 33318 10752 33324 10764
rect 33376 10752 33382 10804
rect 34790 10752 34796 10804
rect 34848 10792 34854 10804
rect 34977 10795 35035 10801
rect 34977 10792 34989 10795
rect 34848 10764 34989 10792
rect 34848 10752 34854 10764
rect 34977 10761 34989 10764
rect 35023 10761 35035 10795
rect 34977 10755 35035 10761
rect 37737 10795 37795 10801
rect 37737 10761 37749 10795
rect 37783 10792 37795 10795
rect 37918 10792 37924 10804
rect 37783 10764 37924 10792
rect 37783 10761 37795 10764
rect 37737 10755 37795 10761
rect 37918 10752 37924 10764
rect 37976 10752 37982 10804
rect 19291 10696 20944 10724
rect 23937 10727 23995 10733
rect 19291 10693 19303 10696
rect 19245 10687 19303 10693
rect 23937 10693 23949 10727
rect 23983 10724 23995 10727
rect 24854 10724 24860 10736
rect 23983 10696 24860 10724
rect 23983 10693 23995 10696
rect 23937 10687 23995 10693
rect 24854 10684 24860 10696
rect 24912 10684 24918 10736
rect 25038 10684 25044 10736
rect 25096 10724 25102 10736
rect 25314 10724 25320 10736
rect 25096 10696 25320 10724
rect 25096 10684 25102 10696
rect 25314 10684 25320 10696
rect 25372 10684 25378 10736
rect 26142 10684 26148 10736
rect 26200 10724 26206 10736
rect 26200 10696 28856 10724
rect 26200 10684 26206 10696
rect 17402 10616 17408 10668
rect 17460 10656 17466 10668
rect 22002 10656 22008 10668
rect 17460 10628 19656 10656
rect 21963 10628 22008 10656
rect 17460 10616 17466 10628
rect 16206 10548 16212 10600
rect 16264 10588 16270 10600
rect 16393 10591 16451 10597
rect 16393 10588 16405 10591
rect 16264 10560 16405 10588
rect 16264 10548 16270 10560
rect 16393 10557 16405 10560
rect 16439 10557 16451 10591
rect 16393 10551 16451 10557
rect 16945 10591 17003 10597
rect 16945 10557 16957 10591
rect 16991 10557 17003 10591
rect 17310 10588 17316 10600
rect 17271 10560 17316 10588
rect 16945 10551 17003 10557
rect 16960 10520 16988 10551
rect 17310 10548 17316 10560
rect 17368 10548 17374 10600
rect 17494 10548 17500 10600
rect 17552 10588 17558 10600
rect 18049 10591 18107 10597
rect 18049 10588 18061 10591
rect 17552 10560 18061 10588
rect 17552 10548 17558 10560
rect 18049 10557 18061 10560
rect 18095 10557 18107 10591
rect 18049 10551 18107 10557
rect 18877 10591 18935 10597
rect 18877 10557 18889 10591
rect 18923 10588 18935 10591
rect 18966 10588 18972 10600
rect 18923 10560 18972 10588
rect 18923 10557 18935 10560
rect 18877 10551 18935 10557
rect 18966 10548 18972 10560
rect 19024 10548 19030 10600
rect 19628 10597 19656 10628
rect 22002 10616 22008 10628
rect 22060 10616 22066 10668
rect 23017 10659 23075 10665
rect 23017 10625 23029 10659
rect 23063 10656 23075 10659
rect 24302 10656 24308 10668
rect 23063 10628 24308 10656
rect 23063 10625 23075 10628
rect 23017 10619 23075 10625
rect 24302 10616 24308 10628
rect 24360 10616 24366 10668
rect 24872 10656 24900 10684
rect 24872 10628 25176 10656
rect 19613 10591 19671 10597
rect 19613 10557 19625 10591
rect 19659 10557 19671 10591
rect 19613 10551 19671 10557
rect 19889 10591 19947 10597
rect 19889 10557 19901 10591
rect 19935 10557 19947 10591
rect 20806 10588 20812 10600
rect 20767 10560 20812 10588
rect 19889 10551 19947 10557
rect 17126 10520 17132 10532
rect 16132 10492 16896 10520
rect 16960 10492 17132 10520
rect 8904 10424 14320 10452
rect 8904 10412 8910 10424
rect 15470 10412 15476 10464
rect 15528 10452 15534 10464
rect 16209 10455 16267 10461
rect 16209 10452 16221 10455
rect 15528 10424 16221 10452
rect 15528 10412 15534 10424
rect 16209 10421 16221 10424
rect 16255 10421 16267 10455
rect 16868 10452 16896 10492
rect 17126 10480 17132 10492
rect 17184 10520 17190 10532
rect 17954 10520 17960 10532
rect 17184 10492 17960 10520
rect 17184 10480 17190 10492
rect 17954 10480 17960 10492
rect 18012 10520 18018 10532
rect 18012 10492 18276 10520
rect 18012 10480 18018 10492
rect 18248 10464 18276 10492
rect 19150 10480 19156 10532
rect 19208 10520 19214 10532
rect 19904 10520 19932 10551
rect 20806 10548 20812 10560
rect 20864 10548 20870 10600
rect 20990 10588 20996 10600
rect 20951 10560 20996 10588
rect 20990 10548 20996 10560
rect 21048 10548 21054 10600
rect 21729 10591 21787 10597
rect 21729 10557 21741 10591
rect 21775 10588 21787 10591
rect 21910 10588 21916 10600
rect 21775 10560 21916 10588
rect 21775 10557 21787 10560
rect 21729 10551 21787 10557
rect 21910 10548 21916 10560
rect 21968 10548 21974 10600
rect 22833 10591 22891 10597
rect 22833 10557 22845 10591
rect 22879 10557 22891 10591
rect 22833 10551 22891 10557
rect 19208 10492 19932 10520
rect 22848 10520 22876 10551
rect 22922 10548 22928 10600
rect 22980 10588 22986 10600
rect 23750 10588 23756 10600
rect 22980 10560 23025 10588
rect 23711 10560 23756 10588
rect 22980 10548 22986 10560
rect 23750 10548 23756 10560
rect 23808 10548 23814 10600
rect 24578 10548 24584 10600
rect 24636 10588 24642 10600
rect 24673 10591 24731 10597
rect 24673 10588 24685 10591
rect 24636 10560 24685 10588
rect 24636 10548 24642 10560
rect 24673 10557 24685 10560
rect 24719 10557 24731 10591
rect 24903 10591 24961 10597
rect 24903 10588 24915 10591
rect 24673 10551 24731 10557
rect 24780 10560 24915 10588
rect 23198 10520 23204 10532
rect 22848 10492 23204 10520
rect 19208 10480 19214 10492
rect 23198 10480 23204 10492
rect 23256 10480 23262 10532
rect 23842 10480 23848 10532
rect 23900 10520 23906 10532
rect 24780 10520 24808 10560
rect 24903 10557 24915 10560
rect 24949 10557 24961 10591
rect 25038 10588 25044 10600
rect 24999 10560 25044 10588
rect 24903 10551 24961 10557
rect 25038 10548 25044 10560
rect 25096 10548 25102 10600
rect 25148 10588 25176 10628
rect 27154 10616 27160 10668
rect 27212 10656 27218 10668
rect 28721 10659 28779 10665
rect 28721 10656 28733 10659
rect 27212 10628 28733 10656
rect 27212 10616 27218 10628
rect 28721 10625 28733 10628
rect 28767 10625 28779 10659
rect 28721 10619 28779 10625
rect 25501 10591 25559 10597
rect 25501 10588 25513 10591
rect 25148 10560 25513 10588
rect 25501 10557 25513 10560
rect 25547 10557 25559 10591
rect 25501 10551 25559 10557
rect 25685 10591 25743 10597
rect 25685 10557 25697 10591
rect 25731 10588 25743 10591
rect 26602 10588 26608 10600
rect 25731 10560 26608 10588
rect 25731 10557 25743 10560
rect 25685 10551 25743 10557
rect 26602 10548 26608 10560
rect 26660 10548 26666 10600
rect 26970 10588 26976 10600
rect 26931 10560 26976 10588
rect 26970 10548 26976 10560
rect 27028 10548 27034 10600
rect 28261 10591 28319 10597
rect 28261 10557 28273 10591
rect 28307 10557 28319 10591
rect 28534 10588 28540 10600
rect 28495 10560 28540 10588
rect 28261 10551 28319 10557
rect 23900 10492 24808 10520
rect 23900 10480 23906 10492
rect 25774 10480 25780 10532
rect 25832 10520 25838 10532
rect 27709 10523 27767 10529
rect 25832 10492 26096 10520
rect 25832 10480 25838 10492
rect 17218 10452 17224 10464
rect 16868 10424 17224 10452
rect 16209 10415 16267 10421
rect 17218 10412 17224 10424
rect 17276 10412 17282 10464
rect 18230 10452 18236 10464
rect 18143 10424 18236 10452
rect 18230 10412 18236 10424
rect 18288 10412 18294 10464
rect 19334 10412 19340 10464
rect 19392 10452 19398 10464
rect 20622 10452 20628 10464
rect 19392 10424 20628 10452
rect 19392 10412 19398 10424
rect 20622 10412 20628 10424
rect 20680 10412 20686 10464
rect 21082 10452 21088 10464
rect 21043 10424 21088 10452
rect 21082 10412 21088 10424
rect 21140 10412 21146 10464
rect 22649 10455 22707 10461
rect 22649 10421 22661 10455
rect 22695 10452 22707 10455
rect 23474 10452 23480 10464
rect 22695 10424 23480 10452
rect 22695 10421 22707 10424
rect 22649 10415 22707 10421
rect 23474 10412 23480 10424
rect 23532 10412 23538 10464
rect 24394 10412 24400 10464
rect 24452 10452 24458 10464
rect 24489 10455 24547 10461
rect 24489 10452 24501 10455
rect 24452 10424 24501 10452
rect 24452 10412 24458 10424
rect 24489 10421 24501 10424
rect 24535 10452 24547 10455
rect 24578 10452 24584 10464
rect 24535 10424 24584 10452
rect 24535 10421 24547 10424
rect 24489 10415 24547 10421
rect 24578 10412 24584 10424
rect 24636 10412 24642 10464
rect 25958 10452 25964 10464
rect 25919 10424 25964 10452
rect 25958 10412 25964 10424
rect 26016 10412 26022 10464
rect 26068 10452 26096 10492
rect 27709 10489 27721 10523
rect 27755 10520 27767 10523
rect 27798 10520 27804 10532
rect 27755 10492 27804 10520
rect 27755 10489 27767 10492
rect 27709 10483 27767 10489
rect 27798 10480 27804 10492
rect 27856 10480 27862 10532
rect 28276 10520 28304 10551
rect 28534 10548 28540 10560
rect 28592 10548 28598 10600
rect 28828 10588 28856 10696
rect 29822 10684 29828 10736
rect 29880 10724 29886 10736
rect 35710 10724 35716 10736
rect 29880 10696 35716 10724
rect 29880 10684 29886 10696
rect 35710 10684 35716 10696
rect 35768 10684 35774 10736
rect 29362 10616 29368 10668
rect 29420 10656 29426 10668
rect 29733 10659 29791 10665
rect 29733 10656 29745 10659
rect 29420 10628 29745 10656
rect 29420 10616 29426 10628
rect 29733 10625 29745 10628
rect 29779 10625 29791 10659
rect 30558 10656 30564 10668
rect 29733 10619 29791 10625
rect 30208 10628 30564 10656
rect 29641 10591 29699 10597
rect 29641 10588 29653 10591
rect 28828 10560 29653 10588
rect 29641 10557 29653 10560
rect 29687 10588 29699 10591
rect 30208 10588 30236 10628
rect 30558 10616 30564 10628
rect 30616 10616 30622 10668
rect 31294 10656 31300 10668
rect 30668 10628 31300 10656
rect 29687 10560 30236 10588
rect 30285 10591 30343 10597
rect 29687 10557 29699 10560
rect 29641 10551 29699 10557
rect 30285 10557 30297 10591
rect 30331 10588 30343 10591
rect 30466 10588 30472 10600
rect 30331 10560 30472 10588
rect 30331 10557 30343 10560
rect 30285 10551 30343 10557
rect 30466 10548 30472 10560
rect 30524 10548 30530 10600
rect 30668 10597 30696 10628
rect 31294 10616 31300 10628
rect 31352 10616 31358 10668
rect 32766 10656 32772 10668
rect 32324 10628 32628 10656
rect 32727 10628 32772 10656
rect 30653 10591 30711 10597
rect 30653 10557 30665 10591
rect 30699 10557 30711 10591
rect 30653 10551 30711 10557
rect 30837 10591 30895 10597
rect 30837 10557 30849 10591
rect 30883 10557 30895 10591
rect 30837 10551 30895 10557
rect 32033 10591 32091 10597
rect 32033 10557 32045 10591
rect 32079 10588 32091 10591
rect 32214 10588 32220 10600
rect 32079 10560 32220 10588
rect 32079 10557 32091 10560
rect 32033 10551 32091 10557
rect 29178 10520 29184 10532
rect 28276 10492 29184 10520
rect 29178 10480 29184 10492
rect 29236 10480 29242 10532
rect 30852 10452 30880 10551
rect 32214 10548 32220 10560
rect 32272 10548 32278 10600
rect 32324 10597 32352 10628
rect 32309 10591 32367 10597
rect 32309 10557 32321 10591
rect 32355 10557 32367 10591
rect 32490 10588 32496 10600
rect 32451 10560 32496 10588
rect 32309 10551 32367 10557
rect 32490 10548 32496 10560
rect 32548 10548 32554 10600
rect 32600 10588 32628 10628
rect 32766 10616 32772 10628
rect 32824 10616 32830 10668
rect 33226 10616 33232 10668
rect 33284 10656 33290 10668
rect 36170 10656 36176 10668
rect 33284 10628 35480 10656
rect 36083 10628 36176 10656
rect 33284 10616 33290 10628
rect 32674 10588 32680 10600
rect 32600 10560 32680 10588
rect 32674 10548 32680 10560
rect 32732 10548 32738 10600
rect 32858 10548 32864 10600
rect 32916 10588 32922 10600
rect 35452 10597 35480 10628
rect 36170 10616 36176 10628
rect 36228 10656 36234 10668
rect 36538 10656 36544 10668
rect 36228 10628 36544 10656
rect 36228 10616 36234 10628
rect 36538 10616 36544 10628
rect 36596 10656 36602 10668
rect 37182 10656 37188 10668
rect 36596 10628 37188 10656
rect 36596 10616 36602 10628
rect 37182 10616 37188 10628
rect 37240 10616 37246 10668
rect 33045 10591 33103 10597
rect 33045 10588 33057 10591
rect 32916 10560 33057 10588
rect 32916 10548 32922 10560
rect 33045 10557 33057 10560
rect 33091 10557 33103 10591
rect 33045 10551 33103 10557
rect 33689 10591 33747 10597
rect 33689 10557 33701 10591
rect 33735 10557 33747 10591
rect 34885 10591 34943 10597
rect 34885 10588 34897 10591
rect 33689 10551 33747 10557
rect 33888 10560 34897 10588
rect 31570 10480 31576 10532
rect 31628 10520 31634 10532
rect 33704 10520 33732 10551
rect 31628 10492 33732 10520
rect 31628 10480 31634 10492
rect 26068 10424 30880 10452
rect 33594 10412 33600 10464
rect 33652 10452 33658 10464
rect 33888 10461 33916 10560
rect 34885 10557 34897 10560
rect 34931 10557 34943 10591
rect 34885 10551 34943 10557
rect 35437 10591 35495 10597
rect 35437 10557 35449 10591
rect 35483 10557 35495 10591
rect 36446 10588 36452 10600
rect 36407 10560 36452 10588
rect 35437 10551 35495 10557
rect 36446 10548 36452 10560
rect 36504 10548 36510 10600
rect 33873 10455 33931 10461
rect 33873 10452 33885 10455
rect 33652 10424 33885 10452
rect 33652 10412 33658 10424
rect 33873 10421 33885 10424
rect 33919 10421 33931 10455
rect 33873 10415 33931 10421
rect 1104 10362 39836 10384
rect 1104 10310 19606 10362
rect 19658 10310 19670 10362
rect 19722 10310 19734 10362
rect 19786 10310 19798 10362
rect 19850 10310 39836 10362
rect 1104 10288 39836 10310
rect 1670 10208 1676 10260
rect 1728 10248 1734 10260
rect 2777 10251 2835 10257
rect 2777 10248 2789 10251
rect 1728 10220 2789 10248
rect 1728 10208 1734 10220
rect 2777 10217 2789 10220
rect 2823 10217 2835 10251
rect 2777 10211 2835 10217
rect 5902 10208 5908 10260
rect 5960 10248 5966 10260
rect 5997 10251 6055 10257
rect 5997 10248 6009 10251
rect 5960 10220 6009 10248
rect 5960 10208 5966 10220
rect 5997 10217 6009 10220
rect 6043 10217 6055 10251
rect 5997 10211 6055 10217
rect 7006 10208 7012 10260
rect 7064 10248 7070 10260
rect 9766 10248 9772 10260
rect 7064 10220 7696 10248
rect 9727 10220 9772 10248
rect 7064 10208 7070 10220
rect 6362 10140 6368 10192
rect 6420 10180 6426 10192
rect 6420 10152 7328 10180
rect 6420 10140 6426 10152
rect 1673 10115 1731 10121
rect 1673 10081 1685 10115
rect 1719 10112 1731 10115
rect 2866 10112 2872 10124
rect 1719 10084 2872 10112
rect 1719 10081 1731 10084
rect 1673 10075 1731 10081
rect 2866 10072 2872 10084
rect 2924 10072 2930 10124
rect 3694 10072 3700 10124
rect 3752 10112 3758 10124
rect 3789 10115 3847 10121
rect 3789 10112 3801 10115
rect 3752 10084 3801 10112
rect 3752 10072 3758 10084
rect 3789 10081 3801 10084
rect 3835 10081 3847 10115
rect 3789 10075 3847 10081
rect 4709 10115 4767 10121
rect 4709 10081 4721 10115
rect 4755 10112 4767 10115
rect 5534 10112 5540 10124
rect 4755 10084 5540 10112
rect 4755 10081 4767 10084
rect 4709 10075 4767 10081
rect 5534 10072 5540 10084
rect 5592 10072 5598 10124
rect 5626 10072 5632 10124
rect 5684 10112 5690 10124
rect 7300 10121 7328 10152
rect 6549 10115 6607 10121
rect 6549 10112 6561 10115
rect 5684 10084 6561 10112
rect 5684 10072 5690 10084
rect 6549 10081 6561 10084
rect 6595 10081 6607 10115
rect 6549 10075 6607 10081
rect 7193 10115 7251 10121
rect 7193 10081 7205 10115
rect 7239 10081 7251 10115
rect 7193 10075 7251 10081
rect 7285 10115 7343 10121
rect 7285 10081 7297 10115
rect 7331 10081 7343 10115
rect 7668 10112 7696 10220
rect 9766 10208 9772 10220
rect 9824 10208 9830 10260
rect 17218 10208 17224 10260
rect 17276 10248 17282 10260
rect 22554 10248 22560 10260
rect 17276 10220 22560 10248
rect 17276 10208 17282 10220
rect 22554 10208 22560 10220
rect 22612 10208 22618 10260
rect 22922 10208 22928 10260
rect 22980 10248 22986 10260
rect 23569 10251 23627 10257
rect 23569 10248 23581 10251
rect 22980 10220 23581 10248
rect 22980 10208 22986 10220
rect 23569 10217 23581 10220
rect 23615 10217 23627 10251
rect 25682 10248 25688 10260
rect 25643 10220 25688 10248
rect 23569 10211 23627 10217
rect 25682 10208 25688 10220
rect 25740 10208 25746 10260
rect 26970 10208 26976 10260
rect 27028 10248 27034 10260
rect 28261 10251 28319 10257
rect 28261 10248 28273 10251
rect 27028 10220 28273 10248
rect 27028 10208 27034 10220
rect 28261 10217 28273 10220
rect 28307 10217 28319 10251
rect 28261 10211 28319 10217
rect 29086 10208 29092 10260
rect 29144 10248 29150 10260
rect 29181 10251 29239 10257
rect 29181 10248 29193 10251
rect 29144 10220 29193 10248
rect 29144 10208 29150 10220
rect 29181 10217 29193 10220
rect 29227 10217 29239 10251
rect 29181 10211 29239 10217
rect 29273 10251 29331 10257
rect 29273 10217 29285 10251
rect 29319 10248 29331 10251
rect 29454 10248 29460 10260
rect 29319 10220 29460 10248
rect 29319 10217 29331 10220
rect 29273 10211 29331 10217
rect 29454 10208 29460 10220
rect 29512 10208 29518 10260
rect 33134 10248 33140 10260
rect 33095 10220 33140 10248
rect 33134 10208 33140 10220
rect 33192 10208 33198 10260
rect 33318 10208 33324 10260
rect 33376 10248 33382 10260
rect 34793 10251 34851 10257
rect 34793 10248 34805 10251
rect 33376 10220 34805 10248
rect 33376 10208 33382 10220
rect 34793 10217 34805 10220
rect 34839 10217 34851 10251
rect 34793 10211 34851 10217
rect 9950 10180 9956 10192
rect 8496 10152 9956 10180
rect 8496 10121 8524 10152
rect 9950 10140 9956 10152
rect 10008 10140 10014 10192
rect 11241 10183 11299 10189
rect 11241 10149 11253 10183
rect 11287 10180 11299 10183
rect 11514 10180 11520 10192
rect 11287 10152 11520 10180
rect 11287 10149 11299 10152
rect 11241 10143 11299 10149
rect 11514 10140 11520 10152
rect 11572 10140 11578 10192
rect 14550 10180 14556 10192
rect 14511 10152 14556 10180
rect 14550 10140 14556 10152
rect 14608 10140 14614 10192
rect 15562 10140 15568 10192
rect 15620 10180 15626 10192
rect 18690 10180 18696 10192
rect 15620 10152 16620 10180
rect 15620 10140 15626 10152
rect 7745 10115 7803 10121
rect 7745 10112 7757 10115
rect 7668 10084 7757 10112
rect 7285 10075 7343 10081
rect 7745 10081 7757 10084
rect 7791 10081 7803 10115
rect 7745 10075 7803 10081
rect 8481 10115 8539 10121
rect 8481 10081 8493 10115
rect 8527 10081 8539 10115
rect 8938 10112 8944 10124
rect 8899 10084 8944 10112
rect 8481 10075 8539 10081
rect 1394 10044 1400 10056
rect 1307 10016 1400 10044
rect 1394 10004 1400 10016
rect 1452 10004 1458 10056
rect 4433 10047 4491 10053
rect 4433 10013 4445 10047
rect 4479 10044 4491 10047
rect 4614 10044 4620 10056
rect 4479 10016 4620 10044
rect 4479 10013 4491 10016
rect 4433 10007 4491 10013
rect 4614 10004 4620 10016
rect 4672 10004 4678 10056
rect 5350 10004 5356 10056
rect 5408 10044 5414 10056
rect 5644 10044 5672 10072
rect 7098 10044 7104 10056
rect 5408 10016 5672 10044
rect 7059 10016 7104 10044
rect 5408 10004 5414 10016
rect 7098 10004 7104 10016
rect 7156 10004 7162 10056
rect 7208 10044 7236 10075
rect 8938 10072 8944 10084
rect 8996 10072 9002 10124
rect 9674 10112 9680 10124
rect 9635 10084 9680 10112
rect 9674 10072 9680 10084
rect 9732 10112 9738 10124
rect 10042 10112 10048 10124
rect 9732 10084 10048 10112
rect 9732 10072 9738 10084
rect 10042 10072 10048 10084
rect 10100 10072 10106 10124
rect 10137 10115 10195 10121
rect 10137 10081 10149 10115
rect 10183 10081 10195 10115
rect 10137 10075 10195 10081
rect 9033 10047 9091 10053
rect 9033 10044 9045 10047
rect 7208 10016 9045 10044
rect 9033 10013 9045 10016
rect 9079 10044 9091 10047
rect 10152 10044 10180 10075
rect 10870 10072 10876 10124
rect 10928 10112 10934 10124
rect 11885 10115 11943 10121
rect 11885 10112 11897 10115
rect 10928 10084 11897 10112
rect 10928 10072 10934 10084
rect 11885 10081 11897 10084
rect 11931 10081 11943 10115
rect 11885 10075 11943 10081
rect 12253 10115 12311 10121
rect 12253 10081 12265 10115
rect 12299 10112 12311 10115
rect 12802 10112 12808 10124
rect 12299 10084 12808 10112
rect 12299 10081 12311 10084
rect 12253 10075 12311 10081
rect 12802 10072 12808 10084
rect 12860 10072 12866 10124
rect 13170 10112 13176 10124
rect 13131 10084 13176 10112
rect 13170 10072 13176 10084
rect 13228 10072 13234 10124
rect 13998 10072 14004 10124
rect 14056 10112 14062 10124
rect 15841 10115 15899 10121
rect 15841 10112 15853 10115
rect 14056 10084 15853 10112
rect 14056 10072 14062 10084
rect 15841 10081 15853 10084
rect 15887 10081 15899 10115
rect 16482 10112 16488 10124
rect 16443 10084 16488 10112
rect 15841 10075 15899 10081
rect 11790 10044 11796 10056
rect 9079 10016 10180 10044
rect 11751 10016 11796 10044
rect 9079 10013 9091 10016
rect 9033 10007 9091 10013
rect 11790 10004 11796 10016
rect 11848 10004 11854 10056
rect 12345 10047 12403 10053
rect 12345 10013 12357 10047
rect 12391 10044 12403 10047
rect 12618 10044 12624 10056
rect 12391 10016 12624 10044
rect 12391 10013 12403 10016
rect 12345 10007 12403 10013
rect 12618 10004 12624 10016
rect 12676 10004 12682 10056
rect 12897 10047 12955 10053
rect 12897 10013 12909 10047
rect 12943 10013 12955 10047
rect 12897 10007 12955 10013
rect 1412 9908 1440 10004
rect 12434 9936 12440 9988
rect 12492 9976 12498 9988
rect 12912 9976 12940 10007
rect 12492 9948 12940 9976
rect 12492 9936 12498 9948
rect 2958 9908 2964 9920
rect 1412 9880 2964 9908
rect 2958 9868 2964 9880
rect 3016 9908 3022 9920
rect 3510 9908 3516 9920
rect 3016 9880 3516 9908
rect 3016 9868 3022 9880
rect 3510 9868 3516 9880
rect 3568 9908 3574 9920
rect 3605 9911 3663 9917
rect 3605 9908 3617 9911
rect 3568 9880 3617 9908
rect 3568 9868 3574 9880
rect 3605 9877 3617 9880
rect 3651 9877 3663 9911
rect 15856 9908 15884 10075
rect 16482 10072 16488 10084
rect 16540 10072 16546 10124
rect 16592 10121 16620 10152
rect 17144 10152 18696 10180
rect 17144 10121 17172 10152
rect 18690 10140 18696 10152
rect 18748 10140 18754 10192
rect 18966 10180 18972 10192
rect 18927 10152 18972 10180
rect 18966 10140 18972 10152
rect 19024 10140 19030 10192
rect 24118 10180 24124 10192
rect 23400 10152 24124 10180
rect 16577 10115 16635 10121
rect 16577 10081 16589 10115
rect 16623 10081 16635 10115
rect 16577 10075 16635 10081
rect 17129 10115 17187 10121
rect 17129 10081 17141 10115
rect 17175 10081 17187 10115
rect 17129 10075 17187 10081
rect 17497 10115 17555 10121
rect 17497 10081 17509 10115
rect 17543 10081 17555 10115
rect 18230 10112 18236 10124
rect 18191 10084 18236 10112
rect 17497 10075 17555 10081
rect 16022 10004 16028 10056
rect 16080 10044 16086 10056
rect 17512 10044 17540 10075
rect 18230 10072 18236 10084
rect 18288 10072 18294 10124
rect 19426 10072 19432 10124
rect 19484 10112 19490 10124
rect 19613 10115 19671 10121
rect 19613 10112 19625 10115
rect 19484 10084 19625 10112
rect 19484 10072 19490 10084
rect 19613 10081 19625 10084
rect 19659 10081 19671 10115
rect 19978 10112 19984 10124
rect 19939 10084 19984 10112
rect 19613 10075 19671 10081
rect 19978 10072 19984 10084
rect 20036 10072 20042 10124
rect 20901 10115 20959 10121
rect 20901 10112 20913 10115
rect 20088 10084 20913 10112
rect 20088 10056 20116 10084
rect 20901 10081 20913 10084
rect 20947 10081 20959 10115
rect 21450 10112 21456 10124
rect 21411 10084 21456 10112
rect 20901 10075 20959 10081
rect 21450 10072 21456 10084
rect 21508 10072 21514 10124
rect 22189 10115 22247 10121
rect 22189 10081 22201 10115
rect 22235 10112 22247 10115
rect 23400 10112 23428 10152
rect 24118 10140 24124 10152
rect 24176 10140 24182 10192
rect 28994 10180 29000 10192
rect 28955 10152 29000 10180
rect 28994 10140 29000 10152
rect 29052 10140 29058 10192
rect 29362 10180 29368 10192
rect 29323 10152 29368 10180
rect 29362 10140 29368 10152
rect 29420 10140 29426 10192
rect 29733 10183 29791 10189
rect 29733 10149 29745 10183
rect 29779 10180 29791 10183
rect 29822 10180 29828 10192
rect 29779 10152 29828 10180
rect 29779 10149 29791 10152
rect 29733 10143 29791 10149
rect 29822 10140 29828 10152
rect 29880 10140 29886 10192
rect 29932 10152 33548 10180
rect 22235 10084 23428 10112
rect 22235 10081 22247 10084
rect 22189 10075 22247 10081
rect 23474 10072 23480 10124
rect 23532 10112 23538 10124
rect 29932 10112 29960 10152
rect 23532 10084 29960 10112
rect 30193 10115 30251 10121
rect 23532 10072 23538 10084
rect 30193 10081 30205 10115
rect 30239 10081 30251 10115
rect 30193 10075 30251 10081
rect 30929 10115 30987 10121
rect 30929 10081 30941 10115
rect 30975 10112 30987 10115
rect 31018 10112 31024 10124
rect 30975 10084 31024 10112
rect 30975 10081 30987 10084
rect 30929 10075 30987 10081
rect 16080 10016 17540 10044
rect 19705 10047 19763 10053
rect 16080 10004 16086 10016
rect 19705 10013 19717 10047
rect 19751 10044 19763 10047
rect 19886 10044 19892 10056
rect 19751 10016 19892 10044
rect 19751 10013 19763 10016
rect 19705 10007 19763 10013
rect 19886 10004 19892 10016
rect 19944 10004 19950 10056
rect 20070 10044 20076 10056
rect 20031 10016 20076 10044
rect 20070 10004 20076 10016
rect 20128 10004 20134 10056
rect 21266 10044 21272 10056
rect 21227 10016 21272 10044
rect 21266 10004 21272 10016
rect 21324 10004 21330 10056
rect 22465 10047 22523 10053
rect 22465 10013 22477 10047
rect 22511 10044 22523 10047
rect 24210 10044 24216 10056
rect 22511 10016 24216 10044
rect 22511 10013 22523 10016
rect 22465 10007 22523 10013
rect 24210 10004 24216 10016
rect 24268 10004 24274 10056
rect 24305 10047 24363 10053
rect 24305 10013 24317 10047
rect 24351 10013 24363 10047
rect 24305 10007 24363 10013
rect 16114 9976 16120 9988
rect 16075 9948 16120 9976
rect 16114 9936 16120 9948
rect 16172 9936 16178 9988
rect 17402 9936 17408 9988
rect 17460 9976 17466 9988
rect 22186 9976 22192 9988
rect 17460 9948 22192 9976
rect 17460 9936 17466 9948
rect 22186 9936 22192 9948
rect 22244 9936 22250 9988
rect 24118 9936 24124 9988
rect 24176 9976 24182 9988
rect 24320 9976 24348 10007
rect 24486 10004 24492 10056
rect 24544 10044 24550 10056
rect 24581 10047 24639 10053
rect 24581 10044 24593 10047
rect 24544 10016 24593 10044
rect 24544 10004 24550 10016
rect 24581 10013 24593 10016
rect 24627 10013 24639 10047
rect 24581 10007 24639 10013
rect 26881 10047 26939 10053
rect 26881 10013 26893 10047
rect 26927 10013 26939 10047
rect 27154 10044 27160 10056
rect 27115 10016 27160 10044
rect 26881 10007 26939 10013
rect 24176 9948 24348 9976
rect 24176 9936 24182 9948
rect 16758 9908 16764 9920
rect 15856 9880 16764 9908
rect 3605 9871 3663 9877
rect 16758 9868 16764 9880
rect 16816 9868 16822 9920
rect 17310 9868 17316 9920
rect 17368 9908 17374 9920
rect 18322 9908 18328 9920
rect 17368 9880 18328 9908
rect 17368 9868 17374 9880
rect 18322 9868 18328 9880
rect 18380 9868 18386 9920
rect 18417 9911 18475 9917
rect 18417 9877 18429 9911
rect 18463 9908 18475 9911
rect 20070 9908 20076 9920
rect 18463 9880 20076 9908
rect 18463 9877 18475 9880
rect 18417 9871 18475 9877
rect 20070 9868 20076 9880
rect 20128 9868 20134 9920
rect 24320 9908 24348 9948
rect 25682 9908 25688 9920
rect 24320 9880 25688 9908
rect 25682 9868 25688 9880
rect 25740 9908 25746 9920
rect 26896 9908 26924 10007
rect 27154 10004 27160 10016
rect 27212 10004 27218 10056
rect 29730 10004 29736 10056
rect 29788 10044 29794 10056
rect 30208 10044 30236 10075
rect 31018 10072 31024 10084
rect 31076 10072 31082 10124
rect 31205 10115 31263 10121
rect 31205 10081 31217 10115
rect 31251 10112 31263 10115
rect 31294 10112 31300 10124
rect 31251 10084 31300 10112
rect 31251 10081 31263 10084
rect 31205 10075 31263 10081
rect 31294 10072 31300 10084
rect 31352 10072 31358 10124
rect 32214 10072 32220 10124
rect 32272 10121 32278 10124
rect 32272 10115 32295 10121
rect 32283 10081 32295 10115
rect 32272 10075 32295 10081
rect 33321 10115 33379 10121
rect 33321 10081 33333 10115
rect 33367 10081 33379 10115
rect 33520 10112 33548 10152
rect 33689 10115 33747 10121
rect 33520 10084 33640 10112
rect 33321 10075 33379 10081
rect 32272 10072 32278 10075
rect 29788 10016 30236 10044
rect 32125 10047 32183 10053
rect 29788 10004 29794 10016
rect 32125 10013 32137 10047
rect 32171 10044 32183 10047
rect 32950 10044 32956 10056
rect 32171 10016 32956 10044
rect 32171 10013 32183 10016
rect 32125 10007 32183 10013
rect 32950 10004 32956 10016
rect 33008 10004 33014 10056
rect 28902 9976 28908 9988
rect 27816 9948 28908 9976
rect 27816 9908 27844 9948
rect 28902 9936 28908 9948
rect 28960 9936 28966 9988
rect 30374 9976 30380 9988
rect 30335 9948 30380 9976
rect 30374 9936 30380 9948
rect 30432 9936 30438 9988
rect 30834 9936 30840 9988
rect 30892 9976 30898 9988
rect 33336 9976 33364 10075
rect 33410 10004 33416 10056
rect 33468 10044 33474 10056
rect 33612 10044 33640 10084
rect 33689 10081 33701 10115
rect 33735 10112 33747 10115
rect 33962 10112 33968 10124
rect 33735 10084 33968 10112
rect 33735 10081 33747 10084
rect 33689 10075 33747 10081
rect 33962 10072 33968 10084
rect 34020 10072 34026 10124
rect 34698 10072 34704 10124
rect 34756 10112 34762 10124
rect 35805 10115 35863 10121
rect 35805 10112 35817 10115
rect 34756 10084 35817 10112
rect 34756 10072 34762 10084
rect 35805 10081 35817 10084
rect 35851 10081 35863 10115
rect 37182 10112 37188 10124
rect 37143 10084 37188 10112
rect 35805 10075 35863 10081
rect 37182 10072 37188 10084
rect 37240 10072 37246 10124
rect 37918 10112 37924 10124
rect 37879 10084 37924 10112
rect 37918 10072 37924 10084
rect 37976 10072 37982 10124
rect 38102 10112 38108 10124
rect 38063 10084 38108 10112
rect 38102 10072 38108 10084
rect 38160 10072 38166 10124
rect 38378 10112 38384 10124
rect 38339 10084 38384 10112
rect 38378 10072 38384 10084
rect 38436 10072 38442 10124
rect 38933 10115 38991 10121
rect 38933 10081 38945 10115
rect 38979 10081 38991 10115
rect 38933 10075 38991 10081
rect 35529 10047 35587 10053
rect 35529 10044 35541 10047
rect 33468 10016 33513 10044
rect 33612 10016 35541 10044
rect 33468 10004 33474 10016
rect 35529 10013 35541 10016
rect 35575 10044 35587 10047
rect 35575 10016 36952 10044
rect 35575 10013 35587 10016
rect 35529 10007 35587 10013
rect 30892 9948 33364 9976
rect 36924 9976 36952 10016
rect 36998 10004 37004 10056
rect 37056 10044 37062 10056
rect 38948 10044 38976 10075
rect 37056 10016 38976 10044
rect 37056 10004 37062 10016
rect 37458 9976 37464 9988
rect 36924 9948 37464 9976
rect 30892 9936 30898 9948
rect 37458 9936 37464 9948
rect 37516 9936 37522 9988
rect 25740 9880 27844 9908
rect 25740 9868 25746 9880
rect 28166 9868 28172 9920
rect 28224 9908 28230 9920
rect 32214 9908 32220 9920
rect 28224 9880 32220 9908
rect 28224 9868 28230 9880
rect 32214 9868 32220 9880
rect 32272 9868 32278 9920
rect 32398 9908 32404 9920
rect 32359 9880 32404 9908
rect 32398 9868 32404 9880
rect 32456 9868 32462 9920
rect 38286 9868 38292 9920
rect 38344 9908 38350 9920
rect 39025 9911 39083 9917
rect 39025 9908 39037 9911
rect 38344 9880 39037 9908
rect 38344 9868 38350 9880
rect 39025 9877 39037 9880
rect 39071 9877 39083 9911
rect 39025 9871 39083 9877
rect 1104 9818 39836 9840
rect 1104 9766 4246 9818
rect 4298 9766 4310 9818
rect 4362 9766 4374 9818
rect 4426 9766 4438 9818
rect 4490 9766 34966 9818
rect 35018 9766 35030 9818
rect 35082 9766 35094 9818
rect 35146 9766 35158 9818
rect 35210 9766 39836 9818
rect 1104 9744 39836 9766
rect 3786 9664 3792 9716
rect 3844 9704 3850 9716
rect 3881 9707 3939 9713
rect 3881 9704 3893 9707
rect 3844 9676 3893 9704
rect 3844 9664 3850 9676
rect 3881 9673 3893 9676
rect 3927 9673 3939 9707
rect 9306 9704 9312 9716
rect 9267 9676 9312 9704
rect 3881 9667 3939 9673
rect 9306 9664 9312 9676
rect 9364 9664 9370 9716
rect 11072 9676 11284 9704
rect 8018 9636 8024 9648
rect 5552 9608 8024 9636
rect 2593 9571 2651 9577
rect 2593 9537 2605 9571
rect 2639 9568 2651 9571
rect 2682 9568 2688 9580
rect 2639 9540 2688 9568
rect 2639 9537 2651 9540
rect 2593 9531 2651 9537
rect 2682 9528 2688 9540
rect 2740 9528 2746 9580
rect 4062 9528 4068 9580
rect 4120 9568 4126 9580
rect 5552 9568 5580 9608
rect 8018 9596 8024 9608
rect 8076 9596 8082 9648
rect 4120 9540 5580 9568
rect 4120 9528 4126 9540
rect 5626 9528 5632 9580
rect 5684 9568 5690 9580
rect 7653 9571 7711 9577
rect 7653 9568 7665 9571
rect 5684 9540 7665 9568
rect 5684 9528 5690 9540
rect 7653 9537 7665 9540
rect 7699 9537 7711 9571
rect 11072 9568 11100 9676
rect 11256 9636 11284 9676
rect 12268 9676 12756 9704
rect 12268 9636 12296 9676
rect 11256 9608 12296 9636
rect 12526 9596 12532 9648
rect 12584 9636 12590 9648
rect 12621 9639 12679 9645
rect 12621 9636 12633 9639
rect 12584 9608 12633 9636
rect 12584 9596 12590 9608
rect 12621 9605 12633 9608
rect 12667 9605 12679 9639
rect 12728 9636 12756 9676
rect 15286 9664 15292 9716
rect 15344 9704 15350 9716
rect 18325 9707 18383 9713
rect 18325 9704 18337 9707
rect 15344 9676 18337 9704
rect 15344 9664 15350 9676
rect 18325 9673 18337 9676
rect 18371 9704 18383 9707
rect 19518 9704 19524 9716
rect 18371 9676 19524 9704
rect 18371 9673 18383 9676
rect 18325 9667 18383 9673
rect 19518 9664 19524 9676
rect 19576 9664 19582 9716
rect 20732 9676 21588 9704
rect 20162 9636 20168 9648
rect 12728 9608 20168 9636
rect 12621 9599 12679 9605
rect 20162 9596 20168 9608
rect 20220 9596 20226 9648
rect 20732 9636 20760 9676
rect 20548 9608 20760 9636
rect 20809 9639 20867 9645
rect 7653 9531 7711 9537
rect 7944 9540 11100 9568
rect 2317 9503 2375 9509
rect 2317 9469 2329 9503
rect 2363 9500 2375 9503
rect 2958 9500 2964 9512
rect 2363 9472 2964 9500
rect 2363 9469 2375 9472
rect 2317 9463 2375 9469
rect 2958 9460 2964 9472
rect 3016 9460 3022 9512
rect 4614 9500 4620 9512
rect 4575 9472 4620 9500
rect 4614 9460 4620 9472
rect 4672 9460 4678 9512
rect 4890 9500 4896 9512
rect 4851 9472 4896 9500
rect 4890 9460 4896 9472
rect 4948 9460 4954 9512
rect 7009 9503 7067 9509
rect 7009 9469 7021 9503
rect 7055 9469 7067 9503
rect 7374 9500 7380 9512
rect 7335 9472 7380 9500
rect 7009 9463 7067 9469
rect 7024 9432 7052 9463
rect 7374 9460 7380 9472
rect 7432 9460 7438 9512
rect 7745 9503 7803 9509
rect 7745 9469 7757 9503
rect 7791 9500 7803 9503
rect 7834 9500 7840 9512
rect 7791 9472 7840 9500
rect 7791 9469 7803 9472
rect 7745 9463 7803 9469
rect 7834 9460 7840 9472
rect 7892 9460 7898 9512
rect 7190 9432 7196 9444
rect 7024 9404 7196 9432
rect 7190 9392 7196 9404
rect 7248 9432 7254 9444
rect 7944 9432 7972 9540
rect 11146 9528 11152 9580
rect 11204 9568 11210 9580
rect 11204 9540 11744 9568
rect 11204 9528 11210 9540
rect 8570 9500 8576 9512
rect 8531 9472 8576 9500
rect 8570 9460 8576 9472
rect 8628 9460 8634 9512
rect 9766 9460 9772 9512
rect 9824 9500 9830 9512
rect 9861 9503 9919 9509
rect 9861 9500 9873 9503
rect 9824 9472 9873 9500
rect 9824 9460 9830 9472
rect 9861 9469 9873 9472
rect 9907 9469 9919 9503
rect 9861 9463 9919 9469
rect 9953 9503 10011 9509
rect 9953 9469 9965 9503
rect 9999 9500 10011 9503
rect 10134 9500 10140 9512
rect 9999 9472 10140 9500
rect 9999 9469 10011 9472
rect 9953 9463 10011 9469
rect 10134 9460 10140 9472
rect 10192 9460 10198 9512
rect 10229 9503 10287 9509
rect 10229 9469 10241 9503
rect 10275 9469 10287 9503
rect 10229 9463 10287 9469
rect 10413 9503 10471 9509
rect 10413 9469 10425 9503
rect 10459 9500 10471 9503
rect 11054 9500 11060 9512
rect 10459 9472 11060 9500
rect 10459 9469 10471 9472
rect 10413 9463 10471 9469
rect 7248 9404 7972 9432
rect 7248 9392 7254 9404
rect 9490 9392 9496 9444
rect 9548 9432 9554 9444
rect 10244 9432 10272 9463
rect 11054 9460 11060 9472
rect 11112 9460 11118 9512
rect 11238 9460 11244 9512
rect 11296 9500 11302 9512
rect 11333 9503 11391 9509
rect 11333 9500 11345 9503
rect 11296 9472 11345 9500
rect 11296 9460 11302 9472
rect 11333 9469 11345 9472
rect 11379 9469 11391 9503
rect 11333 9463 11391 9469
rect 11422 9460 11428 9512
rect 11480 9500 11486 9512
rect 11716 9509 11744 9540
rect 11790 9528 11796 9580
rect 11848 9568 11854 9580
rect 15102 9568 15108 9580
rect 11848 9540 13216 9568
rect 15063 9540 15108 9568
rect 11848 9528 11854 9540
rect 11517 9503 11575 9509
rect 11517 9500 11529 9503
rect 11480 9472 11529 9500
rect 11480 9460 11486 9472
rect 11517 9469 11529 9472
rect 11563 9469 11575 9503
rect 11517 9463 11575 9469
rect 11701 9503 11759 9509
rect 11701 9469 11713 9503
rect 11747 9469 11759 9503
rect 11701 9463 11759 9469
rect 12437 9503 12495 9509
rect 12437 9469 12449 9503
rect 12483 9500 12495 9503
rect 12526 9500 12532 9512
rect 12483 9472 12532 9500
rect 12483 9469 12495 9472
rect 12437 9463 12495 9469
rect 12526 9460 12532 9472
rect 12584 9460 12590 9512
rect 13188 9509 13216 9540
rect 15102 9528 15108 9540
rect 15160 9528 15166 9580
rect 18046 9568 18052 9580
rect 15488 9540 18052 9568
rect 13173 9503 13231 9509
rect 13173 9469 13185 9503
rect 13219 9469 13231 9503
rect 14366 9500 14372 9512
rect 14327 9472 14372 9500
rect 13173 9463 13231 9469
rect 14366 9460 14372 9472
rect 14424 9460 14430 9512
rect 14642 9500 14648 9512
rect 14603 9472 14648 9500
rect 14642 9460 14648 9472
rect 14700 9460 14706 9512
rect 14734 9460 14740 9512
rect 14792 9500 14798 9512
rect 15488 9509 15516 9540
rect 18046 9528 18052 9540
rect 18104 9528 18110 9580
rect 20548 9568 20576 9608
rect 20809 9605 20821 9639
rect 20855 9636 20867 9639
rect 20855 9608 21496 9636
rect 20855 9605 20867 9608
rect 20809 9599 20867 9605
rect 21174 9568 21180 9580
rect 18248 9540 20576 9568
rect 20640 9540 21180 9568
rect 14921 9503 14979 9509
rect 14921 9500 14933 9503
rect 14792 9472 14933 9500
rect 14792 9460 14798 9472
rect 14921 9469 14933 9472
rect 14967 9469 14979 9503
rect 14921 9463 14979 9469
rect 15473 9503 15531 9509
rect 15473 9469 15485 9503
rect 15519 9469 15531 9503
rect 15473 9463 15531 9469
rect 15562 9460 15568 9512
rect 15620 9500 15626 9512
rect 15841 9503 15899 9509
rect 15841 9500 15853 9503
rect 15620 9472 15853 9500
rect 15620 9460 15626 9472
rect 15841 9469 15853 9472
rect 15887 9469 15899 9503
rect 16574 9500 16580 9512
rect 16535 9472 16580 9500
rect 15841 9463 15899 9469
rect 16574 9460 16580 9472
rect 16632 9460 16638 9512
rect 16666 9460 16672 9512
rect 16724 9500 16730 9512
rect 16724 9472 16769 9500
rect 16724 9460 16730 9472
rect 17126 9460 17132 9512
rect 17184 9500 17190 9512
rect 17221 9503 17279 9509
rect 17221 9500 17233 9503
rect 17184 9472 17233 9500
rect 17184 9460 17190 9472
rect 17221 9469 17233 9472
rect 17267 9469 17279 9503
rect 17221 9463 17279 9469
rect 17862 9460 17868 9512
rect 17920 9500 17926 9512
rect 18248 9509 18276 9540
rect 18233 9503 18291 9509
rect 18233 9500 18245 9503
rect 17920 9472 18245 9500
rect 17920 9460 17926 9472
rect 18233 9469 18245 9472
rect 18279 9469 18291 9503
rect 18598 9500 18604 9512
rect 18559 9472 18604 9500
rect 18233 9463 18291 9469
rect 18598 9460 18604 9472
rect 18656 9460 18662 9512
rect 18966 9500 18972 9512
rect 18927 9472 18972 9500
rect 18966 9460 18972 9472
rect 19024 9460 19030 9512
rect 19904 9509 19932 9540
rect 20640 9509 20668 9540
rect 21174 9528 21180 9540
rect 21232 9528 21238 9580
rect 21266 9528 21272 9580
rect 21324 9568 21330 9580
rect 21361 9571 21419 9577
rect 21361 9568 21373 9571
rect 21324 9540 21373 9568
rect 21324 9528 21330 9540
rect 21361 9537 21373 9540
rect 21407 9537 21419 9571
rect 21361 9531 21419 9537
rect 19889 9503 19947 9509
rect 19889 9469 19901 9503
rect 19935 9469 19947 9503
rect 19889 9463 19947 9469
rect 20625 9503 20683 9509
rect 20625 9469 20637 9503
rect 20671 9469 20683 9503
rect 21082 9500 21088 9512
rect 21043 9472 21088 9500
rect 20625 9463 20683 9469
rect 21082 9460 21088 9472
rect 21140 9460 21146 9512
rect 21468 9500 21496 9608
rect 21560 9568 21588 9676
rect 24578 9664 24584 9716
rect 24636 9704 24642 9716
rect 28994 9704 29000 9716
rect 24636 9676 29000 9704
rect 24636 9664 24642 9676
rect 28994 9664 29000 9676
rect 29052 9664 29058 9716
rect 33410 9704 33416 9716
rect 29104 9676 33416 9704
rect 21634 9596 21640 9648
rect 21692 9636 21698 9648
rect 21692 9608 24072 9636
rect 21692 9596 21698 9608
rect 23290 9568 23296 9580
rect 21560 9540 23296 9568
rect 23290 9528 23296 9540
rect 23348 9528 23354 9580
rect 22097 9503 22155 9509
rect 22097 9500 22109 9503
rect 21468 9472 22109 9500
rect 22097 9469 22109 9472
rect 22143 9469 22155 9503
rect 22097 9463 22155 9469
rect 22465 9503 22523 9509
rect 22465 9469 22477 9503
rect 22511 9469 22523 9503
rect 22465 9463 22523 9469
rect 9548 9404 10272 9432
rect 10873 9435 10931 9441
rect 9548 9392 9554 9404
rect 10873 9401 10885 9435
rect 10919 9432 10931 9435
rect 19981 9435 20039 9441
rect 10919 9404 19196 9432
rect 10919 9401 10931 9404
rect 10873 9395 10931 9401
rect 6181 9367 6239 9373
rect 6181 9333 6193 9367
rect 6227 9364 6239 9367
rect 7742 9364 7748 9376
rect 6227 9336 7748 9364
rect 6227 9333 6239 9336
rect 6181 9327 6239 9333
rect 7742 9324 7748 9336
rect 7800 9324 7806 9376
rect 8665 9367 8723 9373
rect 8665 9333 8677 9367
rect 8711 9364 8723 9367
rect 8846 9364 8852 9376
rect 8711 9336 8852 9364
rect 8711 9333 8723 9336
rect 8665 9327 8723 9333
rect 8846 9324 8852 9336
rect 8904 9324 8910 9376
rect 10134 9324 10140 9376
rect 10192 9364 10198 9376
rect 13357 9367 13415 9373
rect 13357 9364 13369 9367
rect 10192 9336 13369 9364
rect 10192 9324 10198 9336
rect 13357 9333 13369 9336
rect 13403 9333 13415 9367
rect 13357 9327 13415 9333
rect 15838 9324 15844 9376
rect 15896 9364 15902 9376
rect 17405 9367 17463 9373
rect 17405 9364 17417 9367
rect 15896 9336 17417 9364
rect 15896 9324 15902 9336
rect 17405 9333 17417 9336
rect 17451 9364 17463 9367
rect 19058 9364 19064 9376
rect 17451 9336 19064 9364
rect 17451 9333 17463 9336
rect 17405 9327 17463 9333
rect 19058 9324 19064 9336
rect 19116 9324 19122 9376
rect 19168 9364 19196 9404
rect 19981 9401 19993 9435
rect 20027 9432 20039 9435
rect 21634 9432 21640 9444
rect 20027 9404 21640 9432
rect 20027 9401 20039 9404
rect 19981 9395 20039 9401
rect 21634 9392 21640 9404
rect 21692 9392 21698 9444
rect 21818 9392 21824 9444
rect 21876 9432 21882 9444
rect 22480 9432 22508 9463
rect 22554 9460 22560 9512
rect 22612 9500 22618 9512
rect 22649 9503 22707 9509
rect 22649 9500 22661 9503
rect 22612 9472 22661 9500
rect 22612 9460 22618 9472
rect 22649 9469 22661 9472
rect 22695 9469 22707 9503
rect 22649 9463 22707 9469
rect 23477 9503 23535 9509
rect 23477 9469 23489 9503
rect 23523 9469 23535 9503
rect 23658 9500 23664 9512
rect 23619 9472 23664 9500
rect 23477 9463 23535 9469
rect 23492 9432 23520 9463
rect 23658 9460 23664 9472
rect 23716 9460 23722 9512
rect 23842 9500 23848 9512
rect 23803 9472 23848 9500
rect 23842 9460 23848 9472
rect 23900 9460 23906 9512
rect 21876 9404 22508 9432
rect 22756 9404 23520 9432
rect 24044 9432 24072 9608
rect 24210 9596 24216 9648
rect 24268 9636 24274 9648
rect 24857 9639 24915 9645
rect 24857 9636 24869 9639
rect 24268 9608 24869 9636
rect 24268 9596 24274 9608
rect 24857 9605 24869 9608
rect 24903 9605 24915 9639
rect 26878 9636 26884 9648
rect 26839 9608 26884 9636
rect 24857 9599 24915 9605
rect 26878 9596 26884 9608
rect 26936 9596 26942 9648
rect 28442 9596 28448 9648
rect 28500 9636 28506 9648
rect 28537 9639 28595 9645
rect 28537 9636 28549 9639
rect 28500 9608 28549 9636
rect 28500 9596 28506 9608
rect 28537 9605 28549 9608
rect 28583 9605 28595 9639
rect 28537 9599 28595 9605
rect 28902 9596 28908 9648
rect 28960 9636 28966 9648
rect 29104 9636 29132 9676
rect 33410 9664 33416 9676
rect 33468 9664 33474 9716
rect 37476 9676 38424 9704
rect 30834 9636 30840 9648
rect 28960 9608 29132 9636
rect 29656 9608 30696 9636
rect 30795 9608 30840 9636
rect 28960 9596 28966 9608
rect 25501 9571 25559 9577
rect 25501 9537 25513 9571
rect 25547 9568 25559 9571
rect 25682 9568 25688 9580
rect 25547 9540 25688 9568
rect 25547 9537 25559 9540
rect 25501 9531 25559 9537
rect 25682 9528 25688 9540
rect 25740 9528 25746 9580
rect 25777 9571 25835 9577
rect 25777 9537 25789 9571
rect 25823 9568 25835 9571
rect 25958 9568 25964 9580
rect 25823 9540 25964 9568
rect 25823 9537 25835 9540
rect 25777 9531 25835 9537
rect 25958 9528 25964 9540
rect 26016 9528 26022 9580
rect 28000 9540 29040 9568
rect 24302 9500 24308 9512
rect 24263 9472 24308 9500
rect 24302 9460 24308 9472
rect 24360 9460 24366 9512
rect 24397 9503 24455 9509
rect 24397 9469 24409 9503
rect 24443 9500 24455 9503
rect 24854 9500 24860 9512
rect 24443 9472 24860 9500
rect 24443 9469 24455 9472
rect 24397 9463 24455 9469
rect 24854 9460 24860 9472
rect 24912 9500 24918 9512
rect 25314 9500 25320 9512
rect 24912 9472 25320 9500
rect 24912 9460 24918 9472
rect 25314 9460 25320 9472
rect 25372 9460 25378 9512
rect 27338 9500 27344 9512
rect 25424 9472 27344 9500
rect 25424 9432 25452 9472
rect 27338 9460 27344 9472
rect 27396 9460 27402 9512
rect 27617 9503 27675 9509
rect 27617 9469 27629 9503
rect 27663 9469 27675 9503
rect 27617 9463 27675 9469
rect 24044 9404 25452 9432
rect 21876 9392 21882 9404
rect 20254 9364 20260 9376
rect 19168 9336 20260 9364
rect 20254 9324 20260 9336
rect 20312 9324 20318 9376
rect 20622 9324 20628 9376
rect 20680 9364 20686 9376
rect 22756 9364 22784 9404
rect 20680 9336 22784 9364
rect 20680 9324 20686 9336
rect 23198 9324 23204 9376
rect 23256 9364 23262 9376
rect 23293 9367 23351 9373
rect 23293 9364 23305 9367
rect 23256 9336 23305 9364
rect 23256 9324 23262 9336
rect 23293 9333 23305 9336
rect 23339 9333 23351 9367
rect 23293 9327 23351 9333
rect 23382 9324 23388 9376
rect 23440 9364 23446 9376
rect 27632 9364 27660 9463
rect 27890 9460 27896 9512
rect 27948 9500 27954 9512
rect 28000 9509 28028 9540
rect 27985 9503 28043 9509
rect 27985 9500 27997 9503
rect 27948 9472 27997 9500
rect 27948 9460 27954 9472
rect 27985 9469 27997 9472
rect 28031 9469 28043 9503
rect 27985 9463 28043 9469
rect 28537 9503 28595 9509
rect 28537 9469 28549 9503
rect 28583 9500 28595 9503
rect 29012 9500 29040 9540
rect 29086 9528 29092 9580
rect 29144 9568 29150 9580
rect 29365 9571 29423 9577
rect 29365 9568 29377 9571
rect 29144 9540 29377 9568
rect 29144 9528 29150 9540
rect 29365 9537 29377 9540
rect 29411 9537 29423 9571
rect 29365 9531 29423 9537
rect 29656 9509 29684 9608
rect 29822 9528 29828 9580
rect 29880 9568 29886 9580
rect 30193 9571 30251 9577
rect 30193 9568 30205 9571
rect 29880 9540 30205 9568
rect 29880 9528 29886 9540
rect 30193 9537 30205 9540
rect 30239 9537 30251 9571
rect 30668 9568 30696 9608
rect 30834 9596 30840 9608
rect 30892 9596 30898 9648
rect 32030 9596 32036 9648
rect 32088 9636 32094 9648
rect 32674 9636 32680 9648
rect 32088 9608 32680 9636
rect 32088 9596 32094 9608
rect 32674 9596 32680 9608
rect 32732 9636 32738 9648
rect 35069 9639 35127 9645
rect 35069 9636 35081 9639
rect 32732 9608 35081 9636
rect 32732 9596 32738 9608
rect 35069 9605 35081 9608
rect 35115 9605 35127 9639
rect 37476 9636 37504 9676
rect 35069 9599 35127 9605
rect 36004 9608 37504 9636
rect 38396 9636 38424 9676
rect 38746 9636 38752 9648
rect 38396 9608 38752 9636
rect 32306 9568 32312 9580
rect 30668 9540 32312 9568
rect 30193 9531 30251 9537
rect 29641 9503 29699 9509
rect 29641 9500 29653 9503
rect 28583 9472 28764 9500
rect 29012 9472 29653 9500
rect 28583 9469 28595 9472
rect 28537 9463 28595 9469
rect 28736 9432 28764 9472
rect 29641 9469 29653 9472
rect 29687 9469 29699 9503
rect 29641 9463 29699 9469
rect 30101 9503 30159 9509
rect 30101 9469 30113 9503
rect 30147 9469 30159 9503
rect 30101 9463 30159 9469
rect 30116 9432 30144 9463
rect 30282 9460 30288 9512
rect 30340 9500 30346 9512
rect 31021 9503 31079 9509
rect 31021 9500 31033 9503
rect 30340 9472 31033 9500
rect 30340 9460 30346 9472
rect 31021 9469 31033 9472
rect 31067 9469 31079 9503
rect 31021 9463 31079 9469
rect 31110 9460 31116 9512
rect 31168 9500 31174 9512
rect 31570 9500 31576 9512
rect 31168 9472 31576 9500
rect 31168 9460 31174 9472
rect 31570 9460 31576 9472
rect 31628 9460 31634 9512
rect 31846 9500 31852 9512
rect 31807 9472 31852 9500
rect 31846 9460 31852 9472
rect 31904 9460 31910 9512
rect 32232 9509 32260 9540
rect 32306 9528 32312 9540
rect 32364 9528 32370 9580
rect 32953 9571 33011 9577
rect 32953 9537 32965 9571
rect 32999 9568 33011 9571
rect 32999 9540 34008 9568
rect 32999 9537 33011 9540
rect 32953 9531 33011 9537
rect 32217 9503 32275 9509
rect 32217 9469 32229 9503
rect 32263 9469 32275 9503
rect 32766 9500 32772 9512
rect 32727 9472 32772 9500
rect 32217 9463 32275 9469
rect 32766 9460 32772 9472
rect 32824 9460 32830 9512
rect 33413 9503 33471 9509
rect 33413 9469 33425 9503
rect 33459 9500 33471 9503
rect 33594 9500 33600 9512
rect 33459 9472 33600 9500
rect 33459 9469 33471 9472
rect 33413 9463 33471 9469
rect 33428 9432 33456 9463
rect 33594 9460 33600 9472
rect 33652 9460 33658 9512
rect 33778 9500 33784 9512
rect 33739 9472 33784 9500
rect 33778 9460 33784 9472
rect 33836 9460 33842 9512
rect 33980 9509 34008 9540
rect 36004 9509 36032 9608
rect 38746 9596 38752 9608
rect 38804 9596 38810 9648
rect 36998 9568 37004 9580
rect 36959 9540 37004 9568
rect 36998 9528 37004 9540
rect 37056 9528 37062 9580
rect 38102 9568 38108 9580
rect 37384 9540 38108 9568
rect 33965 9503 34023 9509
rect 33965 9469 33977 9503
rect 34011 9469 34023 9503
rect 33965 9463 34023 9469
rect 34885 9503 34943 9509
rect 34885 9469 34897 9503
rect 34931 9469 34943 9503
rect 34885 9463 34943 9469
rect 35989 9503 36047 9509
rect 35989 9469 36001 9503
rect 36035 9469 36047 9503
rect 36170 9500 36176 9512
rect 36131 9472 36176 9500
rect 35989 9463 36047 9469
rect 28736 9404 33456 9432
rect 23440 9336 27660 9364
rect 23440 9324 23446 9336
rect 28534 9324 28540 9376
rect 28592 9364 28598 9376
rect 31294 9364 31300 9376
rect 28592 9336 31300 9364
rect 28592 9324 28598 9336
rect 31294 9324 31300 9336
rect 31352 9324 31358 9376
rect 31386 9324 31392 9376
rect 31444 9364 31450 9376
rect 34900 9364 34928 9463
rect 36170 9460 36176 9472
rect 36228 9460 36234 9512
rect 36817 9503 36875 9509
rect 36817 9469 36829 9503
rect 36863 9500 36875 9503
rect 37384 9500 37412 9540
rect 38102 9528 38108 9540
rect 38160 9528 38166 9580
rect 36863 9472 37412 9500
rect 36863 9469 36875 9472
rect 36817 9463 36875 9469
rect 37458 9460 37464 9512
rect 37516 9500 37522 9512
rect 37734 9500 37740 9512
rect 37516 9472 37561 9500
rect 37695 9472 37740 9500
rect 37516 9460 37522 9472
rect 37734 9460 37740 9472
rect 37792 9460 37798 9512
rect 37274 9364 37280 9376
rect 31444 9336 34928 9364
rect 37235 9336 37280 9364
rect 31444 9324 31450 9336
rect 37274 9324 37280 9336
rect 37332 9364 37338 9376
rect 37734 9364 37740 9376
rect 37332 9336 37740 9364
rect 37332 9324 37338 9336
rect 37734 9324 37740 9336
rect 37792 9324 37798 9376
rect 38562 9324 38568 9376
rect 38620 9364 38626 9376
rect 38841 9367 38899 9373
rect 38841 9364 38853 9367
rect 38620 9336 38853 9364
rect 38620 9324 38626 9336
rect 38841 9333 38853 9336
rect 38887 9333 38899 9367
rect 38841 9327 38899 9333
rect 1104 9274 39836 9296
rect 1104 9222 19606 9274
rect 19658 9222 19670 9274
rect 19722 9222 19734 9274
rect 19786 9222 19798 9274
rect 19850 9222 39836 9274
rect 1104 9200 39836 9222
rect 2866 9160 2872 9172
rect 2827 9132 2872 9160
rect 2866 9120 2872 9132
rect 2924 9120 2930 9172
rect 3050 9120 3056 9172
rect 3108 9120 3114 9172
rect 7837 9163 7895 9169
rect 7837 9129 7849 9163
rect 7883 9160 7895 9163
rect 8478 9160 8484 9172
rect 7883 9132 8484 9160
rect 7883 9129 7895 9132
rect 7837 9123 7895 9129
rect 2774 9092 2780 9104
rect 1780 9064 2780 9092
rect 1780 9033 1808 9064
rect 2774 9052 2780 9064
rect 2832 9092 2838 9104
rect 3068 9092 3096 9120
rect 7852 9092 7880 9123
rect 8478 9120 8484 9132
rect 8536 9120 8542 9172
rect 8570 9120 8576 9172
rect 8628 9160 8634 9172
rect 14550 9160 14556 9172
rect 8628 9132 14556 9160
rect 8628 9120 8634 9132
rect 14550 9120 14556 9132
rect 14608 9120 14614 9172
rect 17405 9163 17463 9169
rect 17405 9129 17417 9163
rect 17451 9160 17463 9163
rect 18138 9160 18144 9172
rect 17451 9132 18144 9160
rect 17451 9129 17463 9132
rect 17405 9123 17463 9129
rect 18138 9120 18144 9132
rect 18196 9120 18202 9172
rect 19426 9120 19432 9172
rect 19484 9160 19490 9172
rect 19705 9163 19763 9169
rect 19705 9160 19717 9163
rect 19484 9132 19717 9160
rect 19484 9120 19490 9132
rect 19705 9129 19717 9132
rect 19751 9129 19763 9163
rect 19705 9123 19763 9129
rect 22278 9120 22284 9172
rect 22336 9160 22342 9172
rect 22649 9163 22707 9169
rect 22649 9160 22661 9163
rect 22336 9132 22661 9160
rect 22336 9120 22342 9132
rect 22649 9129 22661 9132
rect 22695 9160 22707 9163
rect 23106 9160 23112 9172
rect 22695 9132 23112 9160
rect 22695 9129 22707 9132
rect 22649 9123 22707 9129
rect 23106 9120 23112 9132
rect 23164 9120 23170 9172
rect 23385 9163 23443 9169
rect 23385 9129 23397 9163
rect 23431 9160 23443 9163
rect 23474 9160 23480 9172
rect 23431 9132 23480 9160
rect 23431 9129 23443 9132
rect 23385 9123 23443 9129
rect 23474 9120 23480 9132
rect 23532 9160 23538 9172
rect 23842 9160 23848 9172
rect 23532 9132 23848 9160
rect 23532 9120 23538 9132
rect 23842 9120 23848 9132
rect 23900 9120 23906 9172
rect 26142 9160 26148 9172
rect 24688 9132 26148 9160
rect 2832 9064 3096 9092
rect 6012 9064 7880 9092
rect 9677 9095 9735 9101
rect 2832 9052 2838 9064
rect 1765 9027 1823 9033
rect 1765 8993 1777 9027
rect 1811 8993 1823 9027
rect 1765 8987 1823 8993
rect 2225 9027 2283 9033
rect 2225 8993 2237 9027
rect 2271 8993 2283 9027
rect 2225 8987 2283 8993
rect 1854 8956 1860 8968
rect 1815 8928 1860 8956
rect 1854 8916 1860 8928
rect 1912 8916 1918 8968
rect 2240 8956 2268 8987
rect 2590 8984 2596 9036
rect 2648 9024 2654 9036
rect 3053 9027 3111 9033
rect 3053 9024 3065 9027
rect 2648 8996 3065 9024
rect 2648 8984 2654 8996
rect 3053 8993 3065 8996
rect 3099 8993 3111 9027
rect 3326 9024 3332 9036
rect 3287 8996 3332 9024
rect 3053 8987 3111 8993
rect 2958 8956 2964 8968
rect 2240 8928 2964 8956
rect 2958 8916 2964 8928
rect 3016 8916 3022 8968
rect 3068 8956 3096 8987
rect 3326 8984 3332 8996
rect 3384 8984 3390 9036
rect 4062 9024 4068 9036
rect 4023 8996 4068 9024
rect 4062 8984 4068 8996
rect 4120 8984 4126 9036
rect 4341 9027 4399 9033
rect 4341 8993 4353 9027
rect 4387 9024 4399 9027
rect 5166 9024 5172 9036
rect 4387 8996 5172 9024
rect 4387 8993 4399 8996
rect 4341 8987 4399 8993
rect 5166 8984 5172 8996
rect 5224 8984 5230 9036
rect 5350 9024 5356 9036
rect 5311 8996 5356 9024
rect 5350 8984 5356 8996
rect 5408 8984 5414 9036
rect 6012 9033 6040 9064
rect 9677 9061 9689 9095
rect 9723 9092 9735 9095
rect 9858 9092 9864 9104
rect 9723 9064 9864 9092
rect 9723 9061 9735 9064
rect 9677 9055 9735 9061
rect 9858 9052 9864 9064
rect 9916 9052 9922 9104
rect 10962 9092 10968 9104
rect 10428 9064 10968 9092
rect 10428 9036 10456 9064
rect 10962 9052 10968 9064
rect 11020 9092 11026 9104
rect 11517 9095 11575 9101
rect 11020 9064 11376 9092
rect 11020 9052 11026 9064
rect 5997 9027 6055 9033
rect 5997 8993 6009 9027
rect 6043 8993 6055 9027
rect 6362 9024 6368 9036
rect 6323 8996 6368 9024
rect 5997 8987 6055 8993
rect 6362 8984 6368 8996
rect 6420 8984 6426 9036
rect 6733 9027 6791 9033
rect 6733 8993 6745 9027
rect 6779 9024 6791 9027
rect 6914 9024 6920 9036
rect 6779 8996 6920 9024
rect 6779 8993 6791 8996
rect 6733 8987 6791 8993
rect 6914 8984 6920 8996
rect 6972 8984 6978 9036
rect 7190 9024 7196 9036
rect 7151 8996 7196 9024
rect 7190 8984 7196 8996
rect 7248 8984 7254 9036
rect 7742 9024 7748 9036
rect 7703 8996 7748 9024
rect 7742 8984 7748 8996
rect 7800 8984 7806 9036
rect 9493 9027 9551 9033
rect 9493 8993 9505 9027
rect 9539 8993 9551 9027
rect 10318 9024 10324 9036
rect 10279 8996 10324 9024
rect 9493 8987 9551 8993
rect 4157 8959 4215 8965
rect 4157 8956 4169 8959
rect 3068 8928 4169 8956
rect 4157 8925 4169 8928
rect 4203 8925 4215 8959
rect 4614 8956 4620 8968
rect 4575 8928 4620 8956
rect 4157 8919 4215 8925
rect 4614 8916 4620 8928
rect 4672 8916 4678 8968
rect 4890 8916 4896 8968
rect 4948 8956 4954 8968
rect 5445 8959 5503 8965
rect 5445 8956 5457 8959
rect 4948 8928 5457 8956
rect 4948 8916 4954 8928
rect 5445 8925 5457 8928
rect 5491 8925 5503 8959
rect 5445 8919 5503 8925
rect 1762 8848 1768 8900
rect 1820 8888 1826 8900
rect 9508 8888 9536 8987
rect 10318 8984 10324 8996
rect 10376 8984 10382 9036
rect 10410 8984 10416 9036
rect 10468 9024 10474 9036
rect 10689 9027 10747 9033
rect 10468 8996 10513 9024
rect 10468 8984 10474 8996
rect 10689 8993 10701 9027
rect 10735 8993 10747 9027
rect 11348 9024 11376 9064
rect 11517 9061 11529 9095
rect 11563 9092 11575 9095
rect 11698 9092 11704 9104
rect 11563 9064 11704 9092
rect 11563 9061 11575 9064
rect 11517 9055 11575 9061
rect 11698 9052 11704 9064
rect 11756 9052 11762 9104
rect 15838 9092 15844 9104
rect 11992 9064 12296 9092
rect 11992 9024 12020 9064
rect 12158 9024 12164 9036
rect 11348 8996 12020 9024
rect 12119 8996 12164 9024
rect 10689 8987 10747 8993
rect 9858 8916 9864 8968
rect 9916 8956 9922 8968
rect 10704 8956 10732 8987
rect 12158 8984 12164 8996
rect 12216 8984 12222 9036
rect 12268 9033 12296 9064
rect 12636 9064 15844 9092
rect 12636 9036 12664 9064
rect 15838 9052 15844 9064
rect 15896 9052 15902 9104
rect 17218 9052 17224 9104
rect 17276 9092 17282 9104
rect 19886 9092 19892 9104
rect 17276 9064 19892 9092
rect 17276 9052 17282 9064
rect 19886 9052 19892 9064
rect 19944 9052 19950 9104
rect 21910 9092 21916 9104
rect 20180 9064 21916 9092
rect 12253 9027 12311 9033
rect 12253 8993 12265 9027
rect 12299 8993 12311 9027
rect 12526 9024 12532 9036
rect 12487 8996 12532 9024
rect 12253 8987 12311 8993
rect 12526 8984 12532 8996
rect 12584 8984 12590 9036
rect 12618 8984 12624 9036
rect 12676 9024 12682 9036
rect 13170 9024 13176 9036
rect 12676 8996 12721 9024
rect 12912 8996 13176 9024
rect 12676 8984 12682 8996
rect 9916 8928 10732 8956
rect 10781 8959 10839 8965
rect 9916 8916 9922 8928
rect 10781 8925 10793 8959
rect 10827 8956 10839 8959
rect 11054 8956 11060 8968
rect 10827 8928 11060 8956
rect 10827 8925 10839 8928
rect 10781 8919 10839 8925
rect 11054 8916 11060 8928
rect 11112 8956 11118 8968
rect 12066 8956 12072 8968
rect 11112 8928 12072 8956
rect 11112 8916 11118 8928
rect 12066 8916 12072 8928
rect 12124 8916 12130 8968
rect 12912 8888 12940 8996
rect 13170 8984 13176 8996
rect 13228 8984 13234 9036
rect 13354 9024 13360 9036
rect 13315 8996 13360 9024
rect 13354 8984 13360 8996
rect 13412 8984 13418 9036
rect 13814 9024 13820 9036
rect 13775 8996 13820 9024
rect 13814 8984 13820 8996
rect 13872 8984 13878 9036
rect 14274 9024 14280 9036
rect 14235 8996 14280 9024
rect 14274 8984 14280 8996
rect 14332 8984 14338 9036
rect 16114 9024 16120 9036
rect 16075 8996 16120 9024
rect 16114 8984 16120 8996
rect 16172 8984 16178 9036
rect 17957 9027 18015 9033
rect 17957 8993 17969 9027
rect 18003 8993 18015 9027
rect 18598 9024 18604 9036
rect 18559 8996 18604 9024
rect 17957 8987 18015 8993
rect 15286 8916 15292 8968
rect 15344 8956 15350 8968
rect 15841 8959 15899 8965
rect 15841 8956 15853 8959
rect 15344 8928 15853 8956
rect 15344 8916 15350 8928
rect 15841 8925 15853 8928
rect 15887 8925 15899 8959
rect 15841 8919 15899 8925
rect 16298 8916 16304 8968
rect 16356 8956 16362 8968
rect 17972 8956 18000 8987
rect 18598 8984 18604 8996
rect 18656 8984 18662 9036
rect 18969 9027 19027 9033
rect 18969 8993 18981 9027
rect 19015 9024 19027 9027
rect 19058 9024 19064 9036
rect 19015 8996 19064 9024
rect 19015 8993 19027 8996
rect 18969 8987 19027 8993
rect 19058 8984 19064 8996
rect 19116 8984 19122 9036
rect 20180 9033 20208 9064
rect 21910 9052 21916 9064
rect 21968 9052 21974 9104
rect 24688 9036 24716 9132
rect 26142 9120 26148 9132
rect 26200 9120 26206 9172
rect 26602 9160 26608 9172
rect 26563 9132 26608 9160
rect 26602 9120 26608 9132
rect 26660 9120 26666 9172
rect 28905 9163 28963 9169
rect 28905 9129 28917 9163
rect 28951 9160 28963 9163
rect 29178 9160 29184 9172
rect 28951 9132 29184 9160
rect 28951 9129 28963 9132
rect 28905 9123 28963 9129
rect 29178 9120 29184 9132
rect 29236 9120 29242 9172
rect 29549 9163 29607 9169
rect 29549 9129 29561 9163
rect 29595 9160 29607 9163
rect 30282 9160 30288 9172
rect 29595 9132 30288 9160
rect 29595 9129 29607 9132
rect 29549 9123 29607 9129
rect 30282 9120 30288 9132
rect 30340 9120 30346 9172
rect 32217 9163 32275 9169
rect 32217 9129 32229 9163
rect 32263 9160 32275 9163
rect 37274 9160 37280 9172
rect 32263 9132 37280 9160
rect 32263 9129 32275 9132
rect 32217 9123 32275 9129
rect 37274 9120 37280 9132
rect 37332 9120 37338 9172
rect 25314 9092 25320 9104
rect 24872 9064 25320 9092
rect 19613 9027 19671 9033
rect 19613 8993 19625 9027
rect 19659 8993 19671 9027
rect 19613 8987 19671 8993
rect 20165 9027 20223 9033
rect 20165 8993 20177 9027
rect 20211 8993 20223 9027
rect 20165 8987 20223 8993
rect 18874 8956 18880 8968
rect 16356 8928 18880 8956
rect 16356 8916 16362 8928
rect 18874 8916 18880 8928
rect 18932 8916 18938 8968
rect 14090 8888 14096 8900
rect 1820 8860 9444 8888
rect 9508 8860 12940 8888
rect 13004 8860 14096 8888
rect 1820 8848 1826 8860
rect 8570 8780 8576 8832
rect 8628 8820 8634 8832
rect 9309 8823 9367 8829
rect 9309 8820 9321 8823
rect 8628 8792 9321 8820
rect 8628 8780 8634 8792
rect 9309 8789 9321 8792
rect 9355 8789 9367 8823
rect 9416 8820 9444 8860
rect 13004 8820 13032 8860
rect 14090 8848 14096 8860
rect 14148 8888 14154 8900
rect 15102 8888 15108 8900
rect 14148 8860 15108 8888
rect 14148 8848 14154 8860
rect 15102 8848 15108 8860
rect 15160 8848 15166 8900
rect 18049 8891 18107 8897
rect 18049 8857 18061 8891
rect 18095 8888 18107 8891
rect 18690 8888 18696 8900
rect 18095 8860 18696 8888
rect 18095 8857 18107 8860
rect 18049 8851 18107 8857
rect 18690 8848 18696 8860
rect 18748 8848 18754 8900
rect 19150 8848 19156 8900
rect 19208 8888 19214 8900
rect 19628 8888 19656 8987
rect 20254 8984 20260 9036
rect 20312 9024 20318 9036
rect 20530 9024 20536 9036
rect 20312 8996 20536 9024
rect 20312 8984 20318 8996
rect 20530 8984 20536 8996
rect 20588 8984 20594 9036
rect 21269 9027 21327 9033
rect 21269 9024 21281 9027
rect 20824 8996 21281 9024
rect 19702 8916 19708 8968
rect 19760 8956 19766 8968
rect 20824 8956 20852 8996
rect 21269 8993 21281 8996
rect 21315 8993 21327 9027
rect 21726 9024 21732 9036
rect 21687 8996 21732 9024
rect 21269 8987 21327 8993
rect 21726 8984 21732 8996
rect 21784 8984 21790 9036
rect 22186 8984 22192 9036
rect 22244 9024 22250 9036
rect 22465 9027 22523 9033
rect 22465 9024 22477 9027
rect 22244 8996 22477 9024
rect 22244 8984 22250 8996
rect 22465 8993 22477 8996
rect 22511 8993 22523 9027
rect 22465 8987 22523 8993
rect 23106 8984 23112 9036
rect 23164 9024 23170 9036
rect 23201 9027 23259 9033
rect 23201 9024 23213 9027
rect 23164 8996 23213 9024
rect 23164 8984 23170 8996
rect 23201 8993 23213 8996
rect 23247 8993 23259 9027
rect 23201 8987 23259 8993
rect 23842 8984 23848 9036
rect 23900 9024 23906 9036
rect 24305 9027 24363 9033
rect 24305 9024 24317 9027
rect 23900 8996 24317 9024
rect 23900 8984 23906 8996
rect 24305 8993 24317 8996
rect 24351 8993 24363 9027
rect 24305 8987 24363 8993
rect 24394 8984 24400 9036
rect 24452 9024 24458 9036
rect 24452 8996 24497 9024
rect 24452 8984 24458 8996
rect 24670 8984 24676 9036
rect 24728 9024 24734 9036
rect 24872 9033 24900 9064
rect 25314 9052 25320 9064
rect 25372 9052 25378 9104
rect 27154 9052 27160 9104
rect 27212 9092 27218 9104
rect 27249 9095 27307 9101
rect 27249 9092 27261 9095
rect 27212 9064 27261 9092
rect 27212 9052 27218 9064
rect 27249 9061 27261 9064
rect 27295 9061 27307 9095
rect 27249 9055 27307 9061
rect 27338 9052 27344 9104
rect 27396 9092 27402 9104
rect 29086 9092 29092 9104
rect 27396 9064 29092 9092
rect 27396 9052 27402 9064
rect 29086 9052 29092 9064
rect 29144 9052 29150 9104
rect 29196 9092 29224 9120
rect 29196 9064 29868 9092
rect 24765 9027 24823 9033
rect 24765 9024 24777 9027
rect 24728 8996 24777 9024
rect 24728 8984 24734 8996
rect 24765 8993 24777 8996
rect 24811 8993 24823 9027
rect 24765 8987 24823 8993
rect 24857 9027 24915 9033
rect 24857 8993 24869 9027
rect 24903 8993 24915 9027
rect 24857 8987 24915 8993
rect 26513 9027 26571 9033
rect 26513 8993 26525 9027
rect 26559 9024 26571 9027
rect 26878 9024 26884 9036
rect 26559 8996 26884 9024
rect 26559 8993 26571 8996
rect 26513 8987 26571 8993
rect 26878 8984 26884 8996
rect 26936 8984 26942 9036
rect 27798 9024 27804 9036
rect 27759 8996 27804 9024
rect 27798 8984 27804 8996
rect 27856 8984 27862 9036
rect 28074 9024 28080 9036
rect 28035 8996 28080 9024
rect 28074 8984 28080 8996
rect 28132 8984 28138 9036
rect 28261 9027 28319 9033
rect 28261 8993 28273 9027
rect 28307 9024 28319 9027
rect 28442 9024 28448 9036
rect 28307 8996 28448 9024
rect 28307 8993 28319 8996
rect 28261 8987 28319 8993
rect 28442 8984 28448 8996
rect 28500 8984 28506 9036
rect 28721 9027 28779 9033
rect 28721 8993 28733 9027
rect 28767 9024 28779 9027
rect 28810 9024 28816 9036
rect 28767 8996 28816 9024
rect 28767 8993 28779 8996
rect 28721 8987 28779 8993
rect 28810 8984 28816 8996
rect 28868 8984 28874 9036
rect 28994 8984 29000 9036
rect 29052 9024 29058 9036
rect 29733 9027 29791 9033
rect 29733 9024 29745 9027
rect 29052 8996 29745 9024
rect 29052 8984 29058 8996
rect 29733 8993 29745 8996
rect 29779 8993 29791 9027
rect 29840 9024 29868 9064
rect 30650 9052 30656 9104
rect 30708 9092 30714 9104
rect 30708 9064 31432 9092
rect 30708 9052 30714 9064
rect 30745 9027 30803 9033
rect 29840 8996 30512 9024
rect 29733 8987 29791 8993
rect 19760 8928 20852 8956
rect 20993 8959 21051 8965
rect 19760 8916 19766 8928
rect 20993 8925 21005 8959
rect 21039 8925 21051 8959
rect 20993 8919 21051 8925
rect 19208 8860 19656 8888
rect 19208 8848 19214 8860
rect 20438 8848 20444 8900
rect 20496 8888 20502 8900
rect 21008 8888 21036 8919
rect 25406 8916 25412 8968
rect 25464 8956 25470 8968
rect 29362 8956 29368 8968
rect 25464 8928 29368 8956
rect 25464 8916 25470 8928
rect 29362 8916 29368 8928
rect 29420 8916 29426 8968
rect 29914 8956 29920 8968
rect 29875 8928 29920 8956
rect 29914 8916 29920 8928
rect 29972 8916 29978 8968
rect 30484 8965 30512 8996
rect 30745 8993 30757 9027
rect 30791 9024 30803 9027
rect 31110 9024 31116 9036
rect 30791 8996 31116 9024
rect 30791 8993 30803 8996
rect 30745 8987 30803 8993
rect 31110 8984 31116 8996
rect 31168 8984 31174 9036
rect 31404 9033 31432 9064
rect 37918 9052 37924 9104
rect 37976 9092 37982 9104
rect 37976 9064 38608 9092
rect 37976 9052 37982 9064
rect 31389 9027 31447 9033
rect 31389 8993 31401 9027
rect 31435 8993 31447 9027
rect 31389 8987 31447 8993
rect 31481 9027 31539 9033
rect 31481 8993 31493 9027
rect 31527 9024 31539 9027
rect 32769 9027 32827 9033
rect 32769 9024 32781 9027
rect 31527 8996 32781 9024
rect 31527 8993 31539 8996
rect 31481 8987 31539 8993
rect 32769 8993 32781 8996
rect 32815 9024 32827 9027
rect 32858 9024 32864 9036
rect 32815 8996 32864 9024
rect 32815 8993 32827 8996
rect 32769 8987 32827 8993
rect 32858 8984 32864 8996
rect 32916 8984 32922 9036
rect 32953 9027 33011 9033
rect 32953 8993 32965 9027
rect 32999 8993 33011 9027
rect 33134 9024 33140 9036
rect 33095 8996 33140 9024
rect 32953 8987 33011 8993
rect 30469 8959 30527 8965
rect 30469 8925 30481 8959
rect 30515 8925 30527 8959
rect 30469 8919 30527 8925
rect 30929 8959 30987 8965
rect 30929 8925 30941 8959
rect 30975 8956 30987 8959
rect 32030 8956 32036 8968
rect 30975 8928 32036 8956
rect 30975 8925 30987 8928
rect 30929 8919 30987 8925
rect 32030 8916 32036 8928
rect 32088 8916 32094 8968
rect 20496 8860 21036 8888
rect 20496 8848 20502 8860
rect 21174 8848 21180 8900
rect 21232 8888 21238 8900
rect 21729 8891 21787 8897
rect 21729 8888 21741 8891
rect 21232 8860 21741 8888
rect 21232 8848 21238 8860
rect 21729 8857 21741 8860
rect 21775 8857 21787 8891
rect 21729 8851 21787 8857
rect 22738 8848 22744 8900
rect 22796 8888 22802 8900
rect 22796 8860 23612 8888
rect 22796 8848 22802 8860
rect 13170 8820 13176 8832
rect 9416 8792 13032 8820
rect 13131 8792 13176 8820
rect 9309 8783 9367 8789
rect 13170 8780 13176 8792
rect 13228 8780 13234 8832
rect 13817 8823 13875 8829
rect 13817 8789 13829 8823
rect 13863 8820 13875 8823
rect 20254 8820 20260 8832
rect 13863 8792 20260 8820
rect 13863 8789 13875 8792
rect 13817 8783 13875 8789
rect 20254 8780 20260 8792
rect 20312 8780 20318 8832
rect 23584 8820 23612 8860
rect 24946 8848 24952 8900
rect 25004 8888 25010 8900
rect 25225 8891 25283 8897
rect 25225 8888 25237 8891
rect 25004 8860 25237 8888
rect 25004 8848 25010 8860
rect 25225 8857 25237 8860
rect 25271 8857 25283 8891
rect 25225 8851 25283 8857
rect 29454 8848 29460 8900
rect 29512 8888 29518 8900
rect 29638 8888 29644 8900
rect 29512 8860 29644 8888
rect 29512 8848 29518 8860
rect 29638 8848 29644 8860
rect 29696 8848 29702 8900
rect 32217 8891 32275 8897
rect 32217 8888 32229 8891
rect 31220 8860 32229 8888
rect 31220 8820 31248 8860
rect 32217 8857 32229 8860
rect 32263 8857 32275 8891
rect 32582 8888 32588 8900
rect 32543 8860 32588 8888
rect 32217 8851 32275 8857
rect 32582 8848 32588 8860
rect 32640 8848 32646 8900
rect 23584 8792 31248 8820
rect 31294 8780 31300 8832
rect 31352 8820 31358 8832
rect 32968 8820 32996 8987
rect 33134 8984 33140 8996
rect 33192 8984 33198 9036
rect 34330 9024 34336 9036
rect 34291 8996 34336 9024
rect 34330 8984 34336 8996
rect 34388 8984 34394 9036
rect 35989 9027 36047 9033
rect 35989 8993 36001 9027
rect 36035 9024 36047 9027
rect 36541 9027 36599 9033
rect 36541 9024 36553 9027
rect 36035 8996 36553 9024
rect 36035 8993 36047 8996
rect 35989 8987 36047 8993
rect 36541 8993 36553 8996
rect 36587 8993 36599 9027
rect 36541 8987 36599 8993
rect 37090 8984 37096 9036
rect 37148 9024 37154 9036
rect 38286 9024 38292 9036
rect 37148 8996 38148 9024
rect 38247 8996 38292 9024
rect 37148 8984 37154 8996
rect 34514 8916 34520 8968
rect 34572 8956 34578 8968
rect 34609 8959 34667 8965
rect 34609 8956 34621 8959
rect 34572 8928 34621 8956
rect 34572 8916 34578 8928
rect 34609 8925 34621 8928
rect 34655 8925 34667 8959
rect 34609 8919 34667 8925
rect 35802 8916 35808 8968
rect 35860 8956 35866 8968
rect 36449 8959 36507 8965
rect 36449 8956 36461 8959
rect 35860 8928 36461 8956
rect 35860 8916 35866 8928
rect 36449 8925 36461 8928
rect 36495 8925 36507 8959
rect 36449 8919 36507 8925
rect 36814 8916 36820 8968
rect 36872 8956 36878 8968
rect 37737 8959 37795 8965
rect 37737 8956 37749 8959
rect 36872 8928 37749 8956
rect 36872 8916 36878 8928
rect 37737 8925 37749 8928
rect 37783 8925 37795 8959
rect 38120 8956 38148 8996
rect 38286 8984 38292 8996
rect 38344 8984 38350 9036
rect 38580 9033 38608 9064
rect 38565 9027 38623 9033
rect 38565 8993 38577 9027
rect 38611 8993 38623 9027
rect 38565 8987 38623 8993
rect 38427 8959 38485 8965
rect 38427 8956 38439 8959
rect 38120 8928 38439 8956
rect 37737 8919 37795 8925
rect 38427 8925 38439 8928
rect 38473 8925 38485 8959
rect 38427 8919 38485 8925
rect 31352 8792 32996 8820
rect 31352 8780 31358 8792
rect 36446 8780 36452 8832
rect 36504 8820 36510 8832
rect 36725 8823 36783 8829
rect 36725 8820 36737 8823
rect 36504 8792 36737 8820
rect 36504 8780 36510 8792
rect 36725 8789 36737 8792
rect 36771 8789 36783 8823
rect 36725 8783 36783 8789
rect 1104 8730 39836 8752
rect 1104 8678 4246 8730
rect 4298 8678 4310 8730
rect 4362 8678 4374 8730
rect 4426 8678 4438 8730
rect 4490 8678 34966 8730
rect 35018 8678 35030 8730
rect 35082 8678 35094 8730
rect 35146 8678 35158 8730
rect 35210 8678 39836 8730
rect 1104 8656 39836 8678
rect 10781 8619 10839 8625
rect 6932 8588 9812 8616
rect 3326 8508 3332 8560
rect 3384 8548 3390 8560
rect 3513 8551 3571 8557
rect 3513 8548 3525 8551
rect 3384 8520 3525 8548
rect 3384 8508 3390 8520
rect 3513 8517 3525 8520
rect 3559 8517 3571 8551
rect 3513 8511 3571 8517
rect 3234 8412 3240 8424
rect 3195 8384 3240 8412
rect 3234 8372 3240 8384
rect 3292 8372 3298 8424
rect 3602 8412 3608 8424
rect 3515 8384 3608 8412
rect 3602 8372 3608 8384
rect 3660 8412 3666 8424
rect 4062 8412 4068 8424
rect 3660 8384 4068 8412
rect 3660 8372 3666 8384
rect 4062 8372 4068 8384
rect 4120 8372 4126 8424
rect 6932 8421 6960 8588
rect 7834 8480 7840 8492
rect 7795 8452 7840 8480
rect 7834 8440 7840 8452
rect 7892 8440 7898 8492
rect 8386 8480 8392 8492
rect 7944 8452 8392 8480
rect 7944 8421 7972 8452
rect 8386 8440 8392 8452
rect 8444 8480 8450 8492
rect 8754 8480 8760 8492
rect 8444 8452 8760 8480
rect 8444 8440 8450 8452
rect 8754 8440 8760 8452
rect 8812 8440 8818 8492
rect 6917 8415 6975 8421
rect 6917 8381 6929 8415
rect 6963 8381 6975 8415
rect 6917 8375 6975 8381
rect 7561 8415 7619 8421
rect 7561 8381 7573 8415
rect 7607 8381 7619 8415
rect 7561 8375 7619 8381
rect 7929 8415 7987 8421
rect 7929 8381 7941 8415
rect 7975 8381 7987 8415
rect 8570 8412 8576 8424
rect 8531 8384 8576 8412
rect 7929 8375 7987 8381
rect 3418 8304 3424 8356
rect 3476 8344 3482 8356
rect 6454 8344 6460 8356
rect 3476 8316 6460 8344
rect 3476 8304 3482 8316
rect 6454 8304 6460 8316
rect 6512 8344 6518 8356
rect 6932 8344 6960 8375
rect 6512 8316 6960 8344
rect 7576 8344 7604 8375
rect 8570 8372 8576 8384
rect 8628 8372 8634 8424
rect 8849 8415 8907 8421
rect 8849 8381 8861 8415
rect 8895 8412 8907 8415
rect 9674 8412 9680 8424
rect 8895 8384 9680 8412
rect 8895 8381 8907 8384
rect 8849 8375 8907 8381
rect 9674 8372 9680 8384
rect 9732 8372 9738 8424
rect 8018 8344 8024 8356
rect 7576 8316 8024 8344
rect 6512 8304 6518 8316
rect 8018 8304 8024 8316
rect 8076 8304 8082 8356
rect 9784 8344 9812 8588
rect 10781 8585 10793 8619
rect 10827 8616 10839 8619
rect 11146 8616 11152 8628
rect 10827 8588 11152 8616
rect 10827 8585 10839 8588
rect 10781 8579 10839 8585
rect 11146 8576 11152 8588
rect 11204 8576 11210 8628
rect 16206 8576 16212 8628
rect 16264 8616 16270 8628
rect 17497 8619 17555 8625
rect 17497 8616 17509 8619
rect 16264 8588 17509 8616
rect 16264 8576 16270 8588
rect 17497 8585 17509 8588
rect 17543 8585 17555 8619
rect 17497 8579 17555 8585
rect 21269 8619 21327 8625
rect 21269 8585 21281 8619
rect 21315 8616 21327 8619
rect 21450 8616 21456 8628
rect 21315 8588 21456 8616
rect 21315 8585 21327 8588
rect 21269 8579 21327 8585
rect 21450 8576 21456 8588
rect 21508 8576 21514 8628
rect 22646 8576 22652 8628
rect 22704 8616 22710 8628
rect 27893 8619 27951 8625
rect 27893 8616 27905 8619
rect 22704 8588 27905 8616
rect 22704 8576 22710 8588
rect 27893 8585 27905 8588
rect 27939 8616 27951 8619
rect 36170 8616 36176 8628
rect 27939 8588 36176 8616
rect 27939 8585 27951 8588
rect 27893 8579 27951 8585
rect 36170 8576 36176 8588
rect 36228 8576 36234 8628
rect 37918 8616 37924 8628
rect 37879 8588 37924 8616
rect 37918 8576 37924 8588
rect 37976 8576 37982 8628
rect 10502 8508 10508 8560
rect 10560 8548 10566 8560
rect 17218 8548 17224 8560
rect 10560 8520 17224 8548
rect 10560 8508 10566 8520
rect 10796 8492 10824 8520
rect 17218 8508 17224 8520
rect 17276 8508 17282 8560
rect 24026 8548 24032 8560
rect 22204 8520 24032 8548
rect 9858 8440 9864 8492
rect 9916 8480 9922 8492
rect 9953 8483 10011 8489
rect 9953 8480 9965 8483
rect 9916 8452 9965 8480
rect 9916 8440 9922 8452
rect 9953 8449 9965 8452
rect 9999 8449 10011 8483
rect 9953 8443 10011 8449
rect 10778 8440 10784 8492
rect 10836 8440 10842 8492
rect 10962 8440 10968 8492
rect 11020 8480 11026 8492
rect 11241 8483 11299 8489
rect 11241 8480 11253 8483
rect 11020 8452 11253 8480
rect 11020 8440 11026 8452
rect 11241 8449 11253 8452
rect 11287 8449 11299 8483
rect 11241 8443 11299 8449
rect 12158 8440 12164 8492
rect 12216 8480 12222 8492
rect 12989 8483 13047 8489
rect 12989 8480 13001 8483
rect 12216 8452 13001 8480
rect 12216 8440 12222 8452
rect 12989 8449 13001 8452
rect 13035 8449 13047 8483
rect 13814 8480 13820 8492
rect 13775 8452 13820 8480
rect 12989 8443 13047 8449
rect 13814 8440 13820 8452
rect 13872 8440 13878 8492
rect 14366 8480 14372 8492
rect 14016 8452 14372 8480
rect 11330 8412 11336 8424
rect 11291 8384 11336 8412
rect 11330 8372 11336 8384
rect 11388 8372 11394 8424
rect 11701 8415 11759 8421
rect 11701 8412 11713 8415
rect 11440 8384 11713 8412
rect 11440 8344 11468 8384
rect 11701 8381 11713 8384
rect 11747 8381 11759 8415
rect 11701 8375 11759 8381
rect 11885 8415 11943 8421
rect 11885 8381 11897 8415
rect 11931 8412 11943 8415
rect 12066 8412 12072 8424
rect 11931 8384 12072 8412
rect 11931 8381 11943 8384
rect 11885 8375 11943 8381
rect 12066 8372 12072 8384
rect 12124 8372 12130 8424
rect 12437 8415 12495 8421
rect 12437 8381 12449 8415
rect 12483 8381 12495 8415
rect 12437 8375 12495 8381
rect 12897 8415 12955 8421
rect 12897 8381 12909 8415
rect 12943 8412 12955 8415
rect 13538 8412 13544 8424
rect 12943 8384 13544 8412
rect 12943 8381 12955 8384
rect 12897 8375 12955 8381
rect 9784 8316 11468 8344
rect 11790 8304 11796 8356
rect 11848 8344 11854 8356
rect 12250 8344 12256 8356
rect 11848 8316 12256 8344
rect 11848 8304 11854 8316
rect 12250 8304 12256 8316
rect 12308 8344 12314 8356
rect 12452 8344 12480 8375
rect 13538 8372 13544 8384
rect 13596 8372 13602 8424
rect 13725 8415 13783 8421
rect 13725 8381 13737 8415
rect 13771 8412 13783 8415
rect 13906 8412 13912 8424
rect 13771 8384 13912 8412
rect 13771 8381 13783 8384
rect 13725 8375 13783 8381
rect 13906 8372 13912 8384
rect 13964 8412 13970 8424
rect 14016 8412 14044 8452
rect 14366 8440 14372 8452
rect 14424 8440 14430 8492
rect 18141 8483 18199 8489
rect 18141 8480 18153 8483
rect 15028 8452 18153 8480
rect 13964 8384 14044 8412
rect 14093 8415 14151 8421
rect 13964 8372 13970 8384
rect 14093 8381 14105 8415
rect 14139 8381 14151 8415
rect 14093 8375 14151 8381
rect 12308 8316 12480 8344
rect 13556 8344 13584 8372
rect 14108 8344 14136 8375
rect 13556 8316 14136 8344
rect 14384 8344 14412 8440
rect 14642 8412 14648 8424
rect 14603 8384 14648 8412
rect 14642 8372 14648 8384
rect 14700 8372 14706 8424
rect 15028 8421 15056 8452
rect 18141 8449 18153 8452
rect 18187 8480 18199 8483
rect 19426 8480 19432 8492
rect 18187 8452 19432 8480
rect 18187 8449 18199 8452
rect 18141 8443 18199 8449
rect 19426 8440 19432 8452
rect 19484 8440 19490 8492
rect 19978 8480 19984 8492
rect 19939 8452 19984 8480
rect 19978 8440 19984 8452
rect 20036 8440 20042 8492
rect 20162 8440 20168 8492
rect 20220 8480 20226 8492
rect 20220 8452 21128 8480
rect 20220 8440 20226 8452
rect 15013 8415 15071 8421
rect 15013 8381 15025 8415
rect 15059 8381 15071 8415
rect 15562 8412 15568 8424
rect 15523 8384 15568 8412
rect 15013 8375 15071 8381
rect 15562 8372 15568 8384
rect 15620 8372 15626 8424
rect 16022 8412 16028 8424
rect 15983 8384 16028 8412
rect 16022 8372 16028 8384
rect 16080 8372 16086 8424
rect 16758 8412 16764 8424
rect 16719 8384 16764 8412
rect 16758 8372 16764 8384
rect 16816 8372 16822 8424
rect 17681 8415 17739 8421
rect 17681 8381 17693 8415
rect 17727 8381 17739 8415
rect 18230 8412 18236 8424
rect 18191 8384 18236 8412
rect 17681 8375 17739 8381
rect 17696 8344 17724 8375
rect 18230 8372 18236 8384
rect 18288 8372 18294 8424
rect 18598 8412 18604 8424
rect 18559 8384 18604 8412
rect 18598 8372 18604 8384
rect 18656 8372 18662 8424
rect 19058 8412 19064 8424
rect 19019 8384 19064 8412
rect 19058 8372 19064 8384
rect 19116 8372 19122 8424
rect 19705 8415 19763 8421
rect 19705 8381 19717 8415
rect 19751 8412 19763 8415
rect 19751 8384 21036 8412
rect 19751 8381 19763 8384
rect 19705 8375 19763 8381
rect 19334 8344 19340 8356
rect 14384 8316 16988 8344
rect 17696 8316 19340 8344
rect 12308 8304 12314 8316
rect 7374 8236 7380 8288
rect 7432 8276 7438 8288
rect 10042 8276 10048 8288
rect 7432 8248 10048 8276
rect 7432 8236 7438 8248
rect 10042 8236 10048 8248
rect 10100 8236 10106 8288
rect 15562 8236 15568 8288
rect 15620 8276 15626 8288
rect 16960 8285 16988 8316
rect 19334 8304 19340 8316
rect 19392 8304 19398 8356
rect 21008 8288 21036 8384
rect 21100 8344 21128 8452
rect 21910 8440 21916 8492
rect 21968 8480 21974 8492
rect 22204 8480 22232 8520
rect 24026 8508 24032 8520
rect 24084 8508 24090 8560
rect 24121 8551 24179 8557
rect 24121 8517 24133 8551
rect 24167 8548 24179 8551
rect 24670 8548 24676 8560
rect 24167 8520 24676 8548
rect 24167 8517 24179 8520
rect 24121 8511 24179 8517
rect 24670 8508 24676 8520
rect 24728 8508 24734 8560
rect 28626 8548 28632 8560
rect 28587 8520 28632 8548
rect 28626 8508 28632 8520
rect 28684 8508 28690 8560
rect 22370 8480 22376 8492
rect 21968 8452 22232 8480
rect 22331 8452 22376 8480
rect 21968 8440 21974 8452
rect 22370 8440 22376 8452
rect 22428 8440 22434 8492
rect 23658 8440 23664 8492
rect 23716 8480 23722 8492
rect 24946 8480 24952 8492
rect 23716 8452 24716 8480
rect 24907 8452 24952 8480
rect 23716 8440 23722 8452
rect 22002 8412 22008 8424
rect 21963 8384 22008 8412
rect 22002 8372 22008 8384
rect 22060 8372 22066 8424
rect 22278 8412 22284 8424
rect 22239 8384 22284 8412
rect 22278 8372 22284 8384
rect 22336 8372 22342 8424
rect 22554 8412 22560 8424
rect 22515 8384 22560 8412
rect 22554 8372 22560 8384
rect 22612 8372 22618 8424
rect 23934 8372 23940 8424
rect 23992 8412 23998 8424
rect 24688 8421 24716 8452
rect 24946 8440 24952 8452
rect 25004 8440 25010 8492
rect 25590 8440 25596 8492
rect 25648 8480 25654 8492
rect 27157 8483 27215 8489
rect 27157 8480 27169 8483
rect 25648 8452 27169 8480
rect 25648 8440 25654 8452
rect 27157 8449 27169 8452
rect 27203 8449 27215 8483
rect 27157 8443 27215 8449
rect 28902 8440 28908 8492
rect 28960 8480 28966 8492
rect 29273 8483 29331 8489
rect 29273 8480 29285 8483
rect 28960 8452 29285 8480
rect 28960 8440 28966 8452
rect 29273 8449 29285 8452
rect 29319 8449 29331 8483
rect 29273 8443 29331 8449
rect 30929 8483 30987 8489
rect 30929 8449 30941 8483
rect 30975 8480 30987 8483
rect 31386 8480 31392 8492
rect 30975 8452 31392 8480
rect 30975 8449 30987 8452
rect 30929 8443 30987 8449
rect 31386 8440 31392 8452
rect 31444 8440 31450 8492
rect 32033 8483 32091 8489
rect 32033 8449 32045 8483
rect 32079 8480 32091 8483
rect 32769 8483 32827 8489
rect 32769 8480 32781 8483
rect 32079 8452 32781 8480
rect 32079 8449 32091 8452
rect 32033 8443 32091 8449
rect 32769 8449 32781 8452
rect 32815 8449 32827 8483
rect 32769 8443 32827 8449
rect 35989 8483 36047 8489
rect 35989 8449 36001 8483
rect 36035 8480 36047 8483
rect 36814 8480 36820 8492
rect 36035 8452 36676 8480
rect 36775 8452 36820 8480
rect 36035 8449 36047 8452
rect 35989 8443 36047 8449
rect 36648 8424 36676 8452
rect 36814 8440 36820 8452
rect 36872 8440 36878 8492
rect 38749 8483 38807 8489
rect 38749 8480 38761 8483
rect 36924 8452 38761 8480
rect 24029 8415 24087 8421
rect 24029 8412 24041 8415
rect 23992 8384 24041 8412
rect 23992 8372 23998 8384
rect 24029 8381 24041 8384
rect 24075 8381 24087 8415
rect 24029 8375 24087 8381
rect 24673 8415 24731 8421
rect 24673 8381 24685 8415
rect 24719 8381 24731 8415
rect 26329 8415 26387 8421
rect 26329 8412 26341 8415
rect 24673 8375 24731 8381
rect 24780 8384 26341 8412
rect 23382 8344 23388 8356
rect 21100 8316 23388 8344
rect 23382 8304 23388 8316
rect 23440 8304 23446 8356
rect 24044 8344 24072 8375
rect 24780 8344 24808 8384
rect 26329 8381 26341 8384
rect 26375 8381 26387 8415
rect 26329 8375 26387 8381
rect 27065 8415 27123 8421
rect 27065 8381 27077 8415
rect 27111 8412 27123 8415
rect 27614 8412 27620 8424
rect 27111 8384 27620 8412
rect 27111 8381 27123 8384
rect 27065 8375 27123 8381
rect 27614 8372 27620 8384
rect 27672 8372 27678 8424
rect 27709 8415 27767 8421
rect 27709 8381 27721 8415
rect 27755 8412 27767 8415
rect 28445 8415 28503 8421
rect 28445 8412 28457 8415
rect 27755 8384 28457 8412
rect 27755 8381 27767 8384
rect 27709 8375 27767 8381
rect 28445 8381 28457 8384
rect 28491 8412 28503 8415
rect 28810 8412 28816 8424
rect 28491 8384 28816 8412
rect 28491 8381 28503 8384
rect 28445 8375 28503 8381
rect 28810 8372 28816 8384
rect 28868 8412 28874 8424
rect 29178 8412 29184 8424
rect 28868 8384 29184 8412
rect 28868 8372 28874 8384
rect 29178 8372 29184 8384
rect 29236 8372 29242 8424
rect 29546 8412 29552 8424
rect 29507 8384 29552 8412
rect 29546 8372 29552 8384
rect 29604 8372 29610 8424
rect 31481 8415 31539 8421
rect 31481 8381 31493 8415
rect 31527 8381 31539 8415
rect 31481 8375 31539 8381
rect 24044 8316 24808 8344
rect 31496 8344 31524 8375
rect 31570 8372 31576 8424
rect 31628 8412 31634 8424
rect 32493 8415 32551 8421
rect 31628 8384 31673 8412
rect 31628 8372 31634 8384
rect 32493 8381 32505 8415
rect 32539 8381 32551 8415
rect 32493 8375 32551 8381
rect 32306 8344 32312 8356
rect 31496 8316 32312 8344
rect 32306 8304 32312 8316
rect 32364 8304 32370 8356
rect 16209 8279 16267 8285
rect 16209 8276 16221 8279
rect 15620 8248 16221 8276
rect 15620 8236 15626 8248
rect 16209 8245 16221 8248
rect 16255 8245 16267 8279
rect 16209 8239 16267 8245
rect 16945 8279 17003 8285
rect 16945 8245 16957 8279
rect 16991 8245 17003 8279
rect 16945 8239 17003 8245
rect 20990 8236 20996 8288
rect 21048 8236 21054 8288
rect 21082 8236 21088 8288
rect 21140 8276 21146 8288
rect 22186 8276 22192 8288
rect 21140 8248 22192 8276
rect 21140 8236 21146 8248
rect 22186 8236 22192 8248
rect 22244 8236 22250 8288
rect 22830 8236 22836 8288
rect 22888 8276 22894 8288
rect 28534 8276 28540 8288
rect 22888 8248 28540 8276
rect 22888 8236 22894 8248
rect 28534 8236 28540 8248
rect 28592 8236 28598 8288
rect 28718 8236 28724 8288
rect 28776 8276 28782 8288
rect 28902 8276 28908 8288
rect 28776 8248 28908 8276
rect 28776 8236 28782 8248
rect 28902 8236 28908 8248
rect 28960 8236 28966 8288
rect 32508 8276 32536 8375
rect 32582 8372 32588 8424
rect 32640 8412 32646 8424
rect 35069 8415 35127 8421
rect 35069 8412 35081 8415
rect 32640 8384 35081 8412
rect 32640 8372 32646 8384
rect 35069 8381 35081 8384
rect 35115 8381 35127 8415
rect 35069 8375 35127 8381
rect 35529 8415 35587 8421
rect 35529 8381 35541 8415
rect 35575 8381 35587 8415
rect 35894 8412 35900 8424
rect 35855 8384 35900 8412
rect 35529 8375 35587 8381
rect 34330 8344 34336 8356
rect 33428 8316 34336 8344
rect 33428 8276 33456 8316
rect 34330 8304 34336 8316
rect 34388 8304 34394 8356
rect 35544 8344 35572 8375
rect 35894 8372 35900 8384
rect 35952 8372 35958 8424
rect 36538 8412 36544 8424
rect 36499 8384 36544 8412
rect 36538 8372 36544 8384
rect 36596 8372 36602 8424
rect 36630 8372 36636 8424
rect 36688 8412 36694 8424
rect 36924 8412 36952 8452
rect 38749 8449 38761 8452
rect 38795 8449 38807 8483
rect 38749 8443 38807 8449
rect 36688 8384 36952 8412
rect 36688 8372 36694 8384
rect 38102 8372 38108 8424
rect 38160 8412 38166 8424
rect 38657 8415 38715 8421
rect 38657 8412 38669 8415
rect 38160 8384 38669 8412
rect 38160 8372 38166 8384
rect 38657 8381 38669 8384
rect 38703 8381 38715 8415
rect 38657 8375 38715 8381
rect 35986 8344 35992 8356
rect 35544 8316 35992 8344
rect 35986 8304 35992 8316
rect 36044 8304 36050 8356
rect 33870 8276 33876 8288
rect 32508 8248 33456 8276
rect 33831 8248 33876 8276
rect 33870 8236 33876 8248
rect 33928 8236 33934 8288
rect 1104 8186 39836 8208
rect 1104 8134 19606 8186
rect 19658 8134 19670 8186
rect 19722 8134 19734 8186
rect 19786 8134 19798 8186
rect 19850 8134 39836 8186
rect 1104 8112 39836 8134
rect 3234 8072 3240 8084
rect 3195 8044 3240 8072
rect 3234 8032 3240 8044
rect 3292 8032 3298 8084
rect 6454 8072 6460 8084
rect 6415 8044 6460 8072
rect 6454 8032 6460 8044
rect 6512 8032 6518 8084
rect 11330 8032 11336 8084
rect 11388 8072 11394 8084
rect 11609 8075 11667 8081
rect 11609 8072 11621 8075
rect 11388 8044 11621 8072
rect 11388 8032 11394 8044
rect 11609 8041 11621 8044
rect 11655 8041 11667 8075
rect 14550 8072 14556 8084
rect 11609 8035 11667 8041
rect 12084 8044 14556 8072
rect 2133 7939 2191 7945
rect 2133 7905 2145 7939
rect 2179 7936 2191 7939
rect 2866 7936 2872 7948
rect 2179 7908 2872 7936
rect 2179 7905 2191 7908
rect 2133 7899 2191 7905
rect 2866 7896 2872 7908
rect 2924 7896 2930 7948
rect 4157 7939 4215 7945
rect 4157 7905 4169 7939
rect 4203 7936 4215 7939
rect 4614 7936 4620 7948
rect 4203 7908 4620 7936
rect 4203 7905 4215 7908
rect 4157 7899 4215 7905
rect 4614 7896 4620 7908
rect 4672 7896 4678 7948
rect 4706 7896 4712 7948
rect 4764 7936 4770 7948
rect 5077 7939 5135 7945
rect 5077 7936 5089 7939
rect 4764 7908 5089 7936
rect 4764 7896 4770 7908
rect 5077 7905 5089 7908
rect 5123 7905 5135 7939
rect 5077 7899 5135 7905
rect 5353 7939 5411 7945
rect 5353 7905 5365 7939
rect 5399 7936 5411 7939
rect 5626 7936 5632 7948
rect 5399 7908 5632 7936
rect 5399 7905 5411 7908
rect 5353 7899 5411 7905
rect 5626 7896 5632 7908
rect 5684 7896 5690 7948
rect 7469 7939 7527 7945
rect 7469 7905 7481 7939
rect 7515 7905 7527 7939
rect 8018 7936 8024 7948
rect 7979 7908 8024 7936
rect 7469 7899 7527 7905
rect 1857 7871 1915 7877
rect 1857 7837 1869 7871
rect 1903 7868 1915 7871
rect 3050 7868 3056 7880
rect 1903 7840 3056 7868
rect 1903 7837 1915 7840
rect 1857 7831 1915 7837
rect 3050 7828 3056 7840
rect 3108 7868 3114 7880
rect 3786 7868 3792 7880
rect 3108 7840 3792 7868
rect 3108 7828 3114 7840
rect 3786 7828 3792 7840
rect 3844 7828 3850 7880
rect 4062 7692 4068 7744
rect 4120 7732 4126 7744
rect 4249 7735 4307 7741
rect 4249 7732 4261 7735
rect 4120 7704 4261 7732
rect 4120 7692 4126 7704
rect 4249 7701 4261 7704
rect 4295 7701 4307 7735
rect 7484 7732 7512 7899
rect 8018 7896 8024 7908
rect 8076 7896 8082 7948
rect 8386 7936 8392 7948
rect 8347 7908 8392 7936
rect 8386 7896 8392 7908
rect 8444 7936 8450 7948
rect 9306 7936 9312 7948
rect 8444 7908 9312 7936
rect 8444 7896 8450 7908
rect 9306 7896 9312 7908
rect 9364 7896 9370 7948
rect 9858 7936 9864 7948
rect 9819 7908 9864 7936
rect 9858 7896 9864 7908
rect 9916 7896 9922 7948
rect 10042 7936 10048 7948
rect 10003 7908 10048 7936
rect 10042 7896 10048 7908
rect 10100 7896 10106 7948
rect 10502 7936 10508 7948
rect 10463 7908 10508 7936
rect 10502 7896 10508 7908
rect 10560 7896 10566 7948
rect 10686 7896 10692 7948
rect 10744 7936 10750 7948
rect 11790 7936 11796 7948
rect 10744 7908 11796 7936
rect 10744 7896 10750 7908
rect 11790 7896 11796 7908
rect 11848 7896 11854 7948
rect 12084 7945 12112 8044
rect 14550 8032 14556 8044
rect 14608 8032 14614 8084
rect 17678 8072 17684 8084
rect 16592 8044 17684 8072
rect 12526 7964 12532 8016
rect 12584 7964 12590 8016
rect 12069 7939 12127 7945
rect 12069 7905 12081 7939
rect 12115 7905 12127 7939
rect 12544 7936 12572 7964
rect 12989 7939 13047 7945
rect 12069 7899 12127 7905
rect 12176 7908 12572 7936
rect 12636 7908 12940 7936
rect 7650 7868 7656 7880
rect 7611 7840 7656 7868
rect 7650 7828 7656 7840
rect 7708 7828 7714 7880
rect 12176 7868 12204 7908
rect 9600 7840 12204 7868
rect 7834 7732 7840 7744
rect 7484 7704 7840 7732
rect 4249 7695 4307 7701
rect 7834 7692 7840 7704
rect 7892 7732 7898 7744
rect 9600 7732 9628 7840
rect 12526 7828 12532 7880
rect 12584 7868 12590 7880
rect 12636 7868 12664 7908
rect 12584 7840 12664 7868
rect 12713 7871 12771 7877
rect 12584 7828 12590 7840
rect 12713 7837 12725 7871
rect 12759 7837 12771 7871
rect 12912 7868 12940 7908
rect 12989 7905 13001 7939
rect 13035 7936 13047 7939
rect 13814 7936 13820 7948
rect 13035 7908 13820 7936
rect 13035 7905 13047 7908
rect 12989 7899 13047 7905
rect 13814 7896 13820 7908
rect 13872 7896 13878 7948
rect 15289 7939 15347 7945
rect 15289 7905 15301 7939
rect 15335 7936 15347 7939
rect 15470 7936 15476 7948
rect 15335 7908 15476 7936
rect 15335 7905 15347 7908
rect 15289 7899 15347 7905
rect 15470 7896 15476 7908
rect 15528 7896 15534 7948
rect 16206 7936 16212 7948
rect 16167 7908 16212 7936
rect 16206 7896 16212 7908
rect 16264 7896 16270 7948
rect 16592 7945 16620 8044
rect 17678 8032 17684 8044
rect 17736 8032 17742 8084
rect 21269 8075 21327 8081
rect 21269 8041 21281 8075
rect 21315 8072 21327 8075
rect 22094 8072 22100 8084
rect 21315 8044 22100 8072
rect 21315 8041 21327 8044
rect 21269 8035 21327 8041
rect 22094 8032 22100 8044
rect 22152 8072 22158 8084
rect 22554 8072 22560 8084
rect 22152 8044 22560 8072
rect 22152 8032 22158 8044
rect 22554 8032 22560 8044
rect 22612 8032 22618 8084
rect 23750 8032 23756 8084
rect 23808 8072 23814 8084
rect 24026 8072 24032 8084
rect 23808 8044 24032 8072
rect 23808 8032 23814 8044
rect 24026 8032 24032 8044
rect 24084 8032 24090 8084
rect 27614 8032 27620 8084
rect 27672 8072 27678 8084
rect 27893 8075 27951 8081
rect 27893 8072 27905 8075
rect 27672 8044 27905 8072
rect 27672 8032 27678 8044
rect 27893 8041 27905 8044
rect 27939 8041 27951 8075
rect 27893 8035 27951 8041
rect 31018 8032 31024 8084
rect 31076 8072 31082 8084
rect 32217 8075 32275 8081
rect 32217 8072 32229 8075
rect 31076 8044 32229 8072
rect 31076 8032 31082 8044
rect 32217 8041 32229 8044
rect 32263 8041 32275 8075
rect 34514 8072 34520 8084
rect 32217 8035 32275 8041
rect 33336 8044 34520 8072
rect 16850 7964 16856 8016
rect 16908 7964 16914 8016
rect 23474 7964 23480 8016
rect 23532 8004 23538 8016
rect 25869 8007 25927 8013
rect 23532 7976 24808 8004
rect 23532 7964 23538 7976
rect 16577 7939 16635 7945
rect 16577 7905 16589 7939
rect 16623 7905 16635 7939
rect 16868 7936 16896 7964
rect 17129 7939 17187 7945
rect 17129 7936 17141 7939
rect 16868 7908 17141 7936
rect 16577 7899 16635 7905
rect 17129 7905 17141 7908
rect 17175 7905 17187 7939
rect 17129 7899 17187 7905
rect 17313 7939 17371 7945
rect 17313 7905 17325 7939
rect 17359 7936 17371 7939
rect 17954 7936 17960 7948
rect 17359 7908 17960 7936
rect 17359 7905 17371 7908
rect 17313 7899 17371 7905
rect 17954 7896 17960 7908
rect 18012 7896 18018 7948
rect 18138 7896 18144 7948
rect 18196 7936 18202 7948
rect 18233 7939 18291 7945
rect 18233 7936 18245 7939
rect 18196 7908 18245 7936
rect 18196 7896 18202 7908
rect 18233 7905 18245 7908
rect 18279 7905 18291 7939
rect 18598 7936 18604 7948
rect 18559 7908 18604 7936
rect 18233 7899 18291 7905
rect 18598 7896 18604 7908
rect 18656 7896 18662 7948
rect 19242 7936 19248 7948
rect 19203 7908 19248 7936
rect 19242 7896 19248 7908
rect 19300 7896 19306 7948
rect 19889 7939 19947 7945
rect 19889 7905 19901 7939
rect 19935 7936 19947 7939
rect 21082 7936 21088 7948
rect 19935 7908 21088 7936
rect 19935 7905 19947 7908
rect 19889 7899 19947 7905
rect 21082 7896 21088 7908
rect 21140 7896 21146 7948
rect 21177 7939 21235 7945
rect 21177 7905 21189 7939
rect 21223 7936 21235 7939
rect 23106 7936 23112 7948
rect 21223 7908 23112 7936
rect 21223 7905 21235 7908
rect 21177 7899 21235 7905
rect 23106 7896 23112 7908
rect 23164 7896 23170 7948
rect 23934 7936 23940 7948
rect 23895 7908 23940 7936
rect 23934 7896 23940 7908
rect 23992 7896 23998 7948
rect 24780 7945 24808 7976
rect 25869 7973 25881 8007
rect 25915 7973 25927 8007
rect 25869 7967 25927 7973
rect 29457 8007 29515 8013
rect 29457 7973 29469 8007
rect 29503 8004 29515 8007
rect 29546 8004 29552 8016
rect 29503 7976 29552 8004
rect 29503 7973 29515 7976
rect 29457 7967 29515 7973
rect 24765 7939 24823 7945
rect 24765 7905 24777 7939
rect 24811 7905 24823 7939
rect 25314 7936 25320 7948
rect 25275 7908 25320 7936
rect 24765 7899 24823 7905
rect 25314 7896 25320 7908
rect 25372 7896 25378 7948
rect 25498 7936 25504 7948
rect 25459 7908 25504 7936
rect 25498 7896 25504 7908
rect 25556 7896 25562 7948
rect 25884 7936 25912 7967
rect 29546 7964 29552 7976
rect 29604 7964 29610 8016
rect 29822 7964 29828 8016
rect 29880 8004 29886 8016
rect 33336 8013 33364 8044
rect 34514 8032 34520 8044
rect 34572 8032 34578 8084
rect 33321 8007 33379 8013
rect 29880 7976 30512 8004
rect 29880 7964 29886 7976
rect 26789 7939 26847 7945
rect 26789 7936 26801 7939
rect 25884 7908 26801 7936
rect 26789 7905 26801 7908
rect 26835 7905 26847 7939
rect 26789 7899 26847 7905
rect 28629 7939 28687 7945
rect 28629 7905 28641 7939
rect 28675 7936 28687 7939
rect 29270 7936 29276 7948
rect 28675 7908 29276 7936
rect 28675 7905 28687 7908
rect 28629 7899 28687 7905
rect 29270 7896 29276 7908
rect 29328 7896 29334 7948
rect 29914 7896 29920 7948
rect 29972 7936 29978 7948
rect 30009 7939 30067 7945
rect 30009 7936 30021 7939
rect 29972 7908 30021 7936
rect 29972 7896 29978 7908
rect 30009 7905 30021 7908
rect 30055 7905 30067 7939
rect 30009 7899 30067 7905
rect 30285 7939 30343 7945
rect 30285 7905 30297 7939
rect 30331 7936 30343 7939
rect 30374 7936 30380 7948
rect 30331 7908 30380 7936
rect 30331 7905 30343 7908
rect 30285 7899 30343 7905
rect 30374 7896 30380 7908
rect 30432 7896 30438 7948
rect 30484 7945 30512 7976
rect 33321 7973 33333 8007
rect 33367 7973 33379 8007
rect 33321 7967 33379 7973
rect 37090 7964 37096 8016
rect 37148 8004 37154 8016
rect 38286 8004 38292 8016
rect 37148 7976 38292 8004
rect 37148 7964 37154 7976
rect 38286 7964 38292 7976
rect 38344 8004 38350 8016
rect 38344 7976 38516 8004
rect 38344 7964 38350 7976
rect 30469 7939 30527 7945
rect 30469 7905 30481 7939
rect 30515 7905 30527 7939
rect 31110 7936 31116 7948
rect 31071 7908 31116 7936
rect 30469 7899 30527 7905
rect 31110 7896 31116 7908
rect 31168 7896 31174 7948
rect 32125 7939 32183 7945
rect 32125 7905 32137 7939
rect 32171 7936 32183 7939
rect 32490 7936 32496 7948
rect 32171 7908 32496 7936
rect 32171 7905 32183 7908
rect 32125 7899 32183 7905
rect 32490 7896 32496 7908
rect 32548 7896 32554 7948
rect 32861 7939 32919 7945
rect 32861 7905 32873 7939
rect 32907 7936 32919 7939
rect 33870 7936 33876 7948
rect 32907 7908 33876 7936
rect 32907 7905 32919 7908
rect 32861 7899 32919 7905
rect 33870 7896 33876 7908
rect 33928 7896 33934 7948
rect 34330 7936 34336 7948
rect 33980 7908 34336 7936
rect 16485 7871 16543 7877
rect 12912 7840 16436 7868
rect 12713 7831 12771 7837
rect 9674 7760 9680 7812
rect 9732 7800 9738 7812
rect 10505 7803 10563 7809
rect 10505 7800 10517 7803
rect 9732 7772 10517 7800
rect 9732 7760 9738 7772
rect 10505 7769 10517 7772
rect 10551 7769 10563 7803
rect 10505 7763 10563 7769
rect 12434 7760 12440 7812
rect 12492 7800 12498 7812
rect 12618 7800 12624 7812
rect 12492 7772 12624 7800
rect 12492 7760 12498 7772
rect 12618 7760 12624 7772
rect 12676 7800 12682 7812
rect 12728 7800 12756 7831
rect 12676 7772 12756 7800
rect 12676 7760 12682 7772
rect 7892 7704 9628 7732
rect 7892 7692 7898 7704
rect 13814 7692 13820 7744
rect 13872 7732 13878 7744
rect 14093 7735 14151 7741
rect 14093 7732 14105 7735
rect 13872 7704 14105 7732
rect 13872 7692 13878 7704
rect 14093 7701 14105 7704
rect 14139 7701 14151 7735
rect 14093 7695 14151 7701
rect 14642 7692 14648 7744
rect 14700 7732 14706 7744
rect 15473 7735 15531 7741
rect 15473 7732 15485 7735
rect 14700 7704 15485 7732
rect 14700 7692 14706 7704
rect 15473 7701 15485 7704
rect 15519 7701 15531 7735
rect 16022 7732 16028 7744
rect 15983 7704 16028 7732
rect 15473 7695 15531 7701
rect 16022 7692 16028 7704
rect 16080 7692 16086 7744
rect 16408 7732 16436 7840
rect 16485 7837 16497 7871
rect 16531 7868 16543 7871
rect 16531 7840 16620 7868
rect 16531 7837 16543 7840
rect 16485 7831 16543 7837
rect 16592 7812 16620 7840
rect 20990 7828 20996 7880
rect 21048 7868 21054 7880
rect 21818 7868 21824 7880
rect 21048 7840 21824 7868
rect 21048 7828 21054 7840
rect 21818 7828 21824 7840
rect 21876 7828 21882 7880
rect 22097 7871 22155 7877
rect 22097 7837 22109 7871
rect 22143 7868 22155 7871
rect 22278 7868 22284 7880
rect 22143 7840 22284 7868
rect 22143 7837 22155 7840
rect 22097 7831 22155 7837
rect 22278 7828 22284 7840
rect 22336 7828 22342 7880
rect 24670 7868 24676 7880
rect 24631 7840 24676 7868
rect 24670 7828 24676 7840
rect 24728 7828 24734 7880
rect 25774 7828 25780 7880
rect 25832 7868 25838 7880
rect 26513 7871 26571 7877
rect 26513 7868 26525 7871
rect 25832 7840 26525 7868
rect 25832 7828 25838 7840
rect 26513 7837 26525 7840
rect 26559 7837 26571 7871
rect 26513 7831 26571 7837
rect 28166 7828 28172 7880
rect 28224 7868 28230 7880
rect 31021 7871 31079 7877
rect 31021 7868 31033 7871
rect 28224 7840 31033 7868
rect 28224 7828 28230 7840
rect 31021 7837 31033 7840
rect 31067 7868 31079 7871
rect 31386 7868 31392 7880
rect 31067 7840 31392 7868
rect 31067 7837 31079 7840
rect 31021 7831 31079 7837
rect 31386 7828 31392 7840
rect 31444 7828 31450 7880
rect 32306 7828 32312 7880
rect 32364 7868 32370 7880
rect 32769 7871 32827 7877
rect 32769 7868 32781 7871
rect 32364 7840 32781 7868
rect 32364 7828 32370 7840
rect 32769 7837 32781 7840
rect 32815 7868 32827 7871
rect 32950 7868 32956 7880
rect 32815 7840 32956 7868
rect 32815 7837 32827 7840
rect 32769 7831 32827 7837
rect 32950 7828 32956 7840
rect 33008 7828 33014 7880
rect 33781 7871 33839 7877
rect 33781 7837 33793 7871
rect 33827 7868 33839 7871
rect 33980 7868 34008 7908
rect 34330 7896 34336 7908
rect 34388 7896 34394 7948
rect 35894 7896 35900 7948
rect 35952 7936 35958 7948
rect 36081 7939 36139 7945
rect 36081 7936 36093 7939
rect 35952 7908 36093 7936
rect 35952 7896 35958 7908
rect 36081 7905 36093 7908
rect 36127 7905 36139 7939
rect 36630 7936 36636 7948
rect 36591 7908 36636 7936
rect 36081 7899 36139 7905
rect 33827 7840 34008 7868
rect 34057 7871 34115 7877
rect 33827 7837 33839 7840
rect 33781 7831 33839 7837
rect 34057 7837 34069 7871
rect 34103 7868 34115 7871
rect 34790 7868 34796 7880
rect 34103 7840 34796 7868
rect 34103 7837 34115 7840
rect 34057 7831 34115 7837
rect 34790 7828 34796 7840
rect 34848 7828 34854 7880
rect 36096 7868 36124 7899
rect 36630 7896 36636 7908
rect 36688 7896 36694 7948
rect 37001 7939 37059 7945
rect 37001 7905 37013 7939
rect 37047 7936 37059 7939
rect 37642 7936 37648 7948
rect 37047 7908 37648 7936
rect 37047 7905 37059 7908
rect 37001 7899 37059 7905
rect 37642 7896 37648 7908
rect 37700 7896 37706 7948
rect 37734 7896 37740 7948
rect 37792 7936 37798 7948
rect 37918 7936 37924 7948
rect 37792 7908 37924 7936
rect 37792 7896 37798 7908
rect 37918 7896 37924 7908
rect 37976 7896 37982 7948
rect 38488 7945 38516 7976
rect 38105 7939 38163 7945
rect 38105 7905 38117 7939
rect 38151 7905 38163 7939
rect 38105 7899 38163 7905
rect 38473 7939 38531 7945
rect 38473 7905 38485 7939
rect 38519 7905 38531 7939
rect 38473 7899 38531 7905
rect 38120 7868 38148 7899
rect 36096 7840 38148 7868
rect 38381 7871 38439 7877
rect 38381 7837 38393 7871
rect 38427 7868 38439 7871
rect 38427 7840 38516 7868
rect 38427 7837 38439 7840
rect 38381 7831 38439 7837
rect 16574 7760 16580 7812
rect 16632 7760 16638 7812
rect 17494 7800 17500 7812
rect 17455 7772 17500 7800
rect 17494 7760 17500 7772
rect 17552 7760 17558 7812
rect 20622 7800 20628 7812
rect 18248 7772 20628 7800
rect 18248 7732 18276 7772
rect 20622 7760 20628 7772
rect 20680 7760 20686 7812
rect 31754 7800 31760 7812
rect 27448 7772 31760 7800
rect 16408 7704 18276 7732
rect 18325 7735 18383 7741
rect 18325 7701 18337 7735
rect 18371 7732 18383 7735
rect 18414 7732 18420 7744
rect 18371 7704 18420 7732
rect 18371 7701 18383 7704
rect 18325 7695 18383 7701
rect 18414 7692 18420 7704
rect 18472 7692 18478 7744
rect 19978 7692 19984 7744
rect 20036 7732 20042 7744
rect 20073 7735 20131 7741
rect 20073 7732 20085 7735
rect 20036 7704 20085 7732
rect 20036 7692 20042 7704
rect 20073 7701 20085 7704
rect 20119 7701 20131 7735
rect 20073 7695 20131 7701
rect 22002 7692 22008 7744
rect 22060 7732 22066 7744
rect 23201 7735 23259 7741
rect 23201 7732 23213 7735
rect 22060 7704 23213 7732
rect 22060 7692 22066 7704
rect 23201 7701 23213 7704
rect 23247 7701 23259 7735
rect 23201 7695 23259 7701
rect 23842 7692 23848 7744
rect 23900 7732 23906 7744
rect 24394 7732 24400 7744
rect 23900 7704 24400 7732
rect 23900 7692 23906 7704
rect 24394 7692 24400 7704
rect 24452 7732 24458 7744
rect 27448 7732 27476 7772
rect 31754 7760 31760 7772
rect 31812 7760 31818 7812
rect 24452 7704 27476 7732
rect 24452 7692 24458 7704
rect 28534 7692 28540 7744
rect 28592 7732 28598 7744
rect 28813 7735 28871 7741
rect 28813 7732 28825 7735
rect 28592 7704 28825 7732
rect 28592 7692 28598 7704
rect 28813 7701 28825 7704
rect 28859 7701 28871 7735
rect 28813 7695 28871 7701
rect 30926 7692 30932 7744
rect 30984 7732 30990 7744
rect 31297 7735 31355 7741
rect 31297 7732 31309 7735
rect 30984 7704 31309 7732
rect 30984 7692 30990 7704
rect 31297 7701 31309 7704
rect 31343 7701 31355 7735
rect 32968 7732 32996 7828
rect 38488 7812 38516 7840
rect 35986 7760 35992 7812
rect 36044 7800 36050 7812
rect 36909 7803 36967 7809
rect 36909 7800 36921 7803
rect 36044 7772 36921 7800
rect 36044 7760 36050 7772
rect 36909 7769 36921 7772
rect 36955 7769 36967 7803
rect 36909 7763 36967 7769
rect 38470 7760 38476 7812
rect 38528 7760 38534 7812
rect 34514 7732 34520 7744
rect 32968 7704 34520 7732
rect 31297 7695 31355 7701
rect 34514 7692 34520 7704
rect 34572 7692 34578 7744
rect 35345 7735 35403 7741
rect 35345 7701 35357 7735
rect 35391 7732 35403 7735
rect 36722 7732 36728 7744
rect 35391 7704 36728 7732
rect 35391 7701 35403 7704
rect 35345 7695 35403 7701
rect 36722 7692 36728 7704
rect 36780 7692 36786 7744
rect 1104 7642 39836 7664
rect 1104 7590 4246 7642
rect 4298 7590 4310 7642
rect 4362 7590 4374 7642
rect 4426 7590 4438 7642
rect 4490 7590 34966 7642
rect 35018 7590 35030 7642
rect 35082 7590 35094 7642
rect 35146 7590 35158 7642
rect 35210 7590 39836 7642
rect 1104 7568 39836 7590
rect 2958 7488 2964 7540
rect 3016 7528 3022 7540
rect 3145 7531 3203 7537
rect 3145 7528 3157 7531
rect 3016 7500 3157 7528
rect 3016 7488 3022 7500
rect 3145 7497 3157 7500
rect 3191 7497 3203 7531
rect 5166 7528 5172 7540
rect 5127 7500 5172 7528
rect 3145 7491 3203 7497
rect 5166 7488 5172 7500
rect 5224 7488 5230 7540
rect 7190 7528 7196 7540
rect 7024 7500 7196 7528
rect 1854 7352 1860 7404
rect 1912 7392 1918 7404
rect 2133 7395 2191 7401
rect 2133 7392 2145 7395
rect 1912 7364 2145 7392
rect 1912 7352 1918 7364
rect 2133 7361 2145 7364
rect 2179 7361 2191 7395
rect 2133 7355 2191 7361
rect 2593 7395 2651 7401
rect 2593 7361 2605 7395
rect 2639 7392 2651 7395
rect 3234 7392 3240 7404
rect 2639 7364 3240 7392
rect 2639 7361 2651 7364
rect 2593 7355 2651 7361
rect 3234 7352 3240 7364
rect 3292 7352 3298 7404
rect 4062 7392 4068 7404
rect 4023 7364 4068 7392
rect 4062 7352 4068 7364
rect 4120 7352 4126 7404
rect 7024 7401 7052 7500
rect 7190 7488 7196 7500
rect 7248 7528 7254 7540
rect 12526 7528 12532 7540
rect 7248 7500 12532 7528
rect 7248 7488 7254 7500
rect 12526 7488 12532 7500
rect 12584 7488 12590 7540
rect 14366 7488 14372 7540
rect 14424 7528 14430 7540
rect 19978 7528 19984 7540
rect 14424 7500 19984 7528
rect 14424 7488 14430 7500
rect 19978 7488 19984 7500
rect 20036 7488 20042 7540
rect 21082 7488 21088 7540
rect 21140 7528 21146 7540
rect 23842 7528 23848 7540
rect 21140 7500 23848 7528
rect 21140 7488 21146 7500
rect 23842 7488 23848 7500
rect 23900 7488 23906 7540
rect 23934 7488 23940 7540
rect 23992 7528 23998 7540
rect 25041 7531 25099 7537
rect 25041 7528 25053 7531
rect 23992 7500 25053 7528
rect 23992 7488 23998 7500
rect 25041 7497 25053 7500
rect 25087 7497 25099 7531
rect 26234 7528 26240 7540
rect 26195 7500 26240 7528
rect 25041 7491 25099 7497
rect 26234 7488 26240 7500
rect 26292 7528 26298 7540
rect 26292 7500 30880 7528
rect 26292 7488 26298 7500
rect 7282 7420 7288 7472
rect 7340 7460 7346 7472
rect 7653 7463 7711 7469
rect 7653 7460 7665 7463
rect 7340 7432 7665 7460
rect 7340 7420 7346 7432
rect 7653 7429 7665 7432
rect 7699 7429 7711 7463
rect 7653 7423 7711 7429
rect 9950 7420 9956 7472
rect 10008 7460 10014 7472
rect 18138 7460 18144 7472
rect 10008 7432 18144 7460
rect 10008 7420 10014 7432
rect 18138 7420 18144 7432
rect 18196 7420 18202 7472
rect 22278 7460 22284 7472
rect 22239 7432 22284 7460
rect 22278 7420 22284 7432
rect 22336 7420 22342 7472
rect 27430 7420 27436 7472
rect 27488 7460 27494 7472
rect 29365 7463 29423 7469
rect 29365 7460 29377 7463
rect 27488 7432 29377 7460
rect 27488 7420 27494 7432
rect 29365 7429 29377 7432
rect 29411 7429 29423 7463
rect 30852 7460 30880 7500
rect 31110 7488 31116 7540
rect 31168 7528 31174 7540
rect 31297 7531 31355 7537
rect 31297 7528 31309 7531
rect 31168 7500 31309 7528
rect 31168 7488 31174 7500
rect 31297 7497 31309 7500
rect 31343 7497 31355 7531
rect 31297 7491 31355 7497
rect 31386 7488 31392 7540
rect 31444 7528 31450 7540
rect 35802 7528 35808 7540
rect 31444 7500 35808 7528
rect 31444 7488 31450 7500
rect 35802 7488 35808 7500
rect 35860 7488 35866 7540
rect 35894 7488 35900 7540
rect 35952 7528 35958 7540
rect 36541 7531 36599 7537
rect 36541 7528 36553 7531
rect 35952 7500 36553 7528
rect 35952 7488 35958 7500
rect 36541 7497 36553 7500
rect 36587 7497 36599 7531
rect 36541 7491 36599 7497
rect 32122 7460 32128 7472
rect 30852 7432 32128 7460
rect 29365 7423 29423 7429
rect 32122 7420 32128 7432
rect 32180 7420 32186 7472
rect 36556 7460 36584 7491
rect 36556 7432 37964 7460
rect 7009 7395 7067 7401
rect 7009 7361 7021 7395
rect 7055 7361 7067 7395
rect 9766 7392 9772 7404
rect 7009 7355 7067 7361
rect 8956 7364 9772 7392
rect 2409 7327 2467 7333
rect 2409 7293 2421 7327
rect 2455 7324 2467 7327
rect 2774 7324 2780 7336
rect 2455 7296 2780 7324
rect 2455 7293 2467 7296
rect 2409 7287 2467 7293
rect 2774 7284 2780 7296
rect 2832 7284 2838 7336
rect 3053 7327 3111 7333
rect 3053 7293 3065 7327
rect 3099 7293 3111 7327
rect 3786 7324 3792 7336
rect 3747 7296 3792 7324
rect 3053 7287 3111 7293
rect 1578 7256 1584 7268
rect 1539 7228 1584 7256
rect 1578 7216 1584 7228
rect 1636 7216 1642 7268
rect 1762 7216 1768 7268
rect 1820 7256 1826 7268
rect 3068 7256 3096 7287
rect 3786 7284 3792 7296
rect 3844 7284 3850 7336
rect 7374 7324 7380 7336
rect 7335 7296 7380 7324
rect 7374 7284 7380 7296
rect 7432 7284 7438 7336
rect 7650 7324 7656 7336
rect 7611 7296 7656 7324
rect 7650 7284 7656 7296
rect 7708 7284 7714 7336
rect 8956 7333 8984 7364
rect 9766 7352 9772 7364
rect 9824 7352 9830 7404
rect 9861 7395 9919 7401
rect 9861 7361 9873 7395
rect 9907 7392 9919 7395
rect 10502 7392 10508 7404
rect 9907 7364 10508 7392
rect 9907 7361 9919 7364
rect 9861 7355 9919 7361
rect 10502 7352 10508 7364
rect 10560 7352 10566 7404
rect 12986 7392 12992 7404
rect 12947 7364 12992 7392
rect 12986 7352 12992 7364
rect 13044 7352 13050 7404
rect 13998 7392 14004 7404
rect 13959 7364 14004 7392
rect 13998 7352 14004 7364
rect 14056 7352 14062 7404
rect 18966 7392 18972 7404
rect 15304 7364 18460 7392
rect 18927 7364 18972 7392
rect 8941 7327 8999 7333
rect 8941 7293 8953 7327
rect 8987 7293 8999 7327
rect 8941 7287 8999 7293
rect 9217 7327 9275 7333
rect 9217 7293 9229 7327
rect 9263 7293 9275 7327
rect 9217 7287 9275 7293
rect 1820 7228 3096 7256
rect 1820 7216 1826 7228
rect 8018 7216 8024 7268
rect 8076 7256 8082 7268
rect 9232 7256 9260 7287
rect 9306 7284 9312 7336
rect 9364 7324 9370 7336
rect 9493 7327 9551 7333
rect 9493 7324 9505 7327
rect 9364 7296 9505 7324
rect 9364 7284 9370 7296
rect 9493 7293 9505 7296
rect 9539 7293 9551 7327
rect 9493 7287 9551 7293
rect 10597 7327 10655 7333
rect 10597 7293 10609 7327
rect 10643 7324 10655 7327
rect 10686 7324 10692 7336
rect 10643 7296 10692 7324
rect 10643 7293 10655 7296
rect 10597 7287 10655 7293
rect 10686 7284 10692 7296
rect 10744 7284 10750 7336
rect 10870 7324 10876 7336
rect 10831 7296 10876 7324
rect 10870 7284 10876 7296
rect 10928 7284 10934 7336
rect 11517 7327 11575 7333
rect 11517 7293 11529 7327
rect 11563 7324 11575 7327
rect 11606 7324 11612 7336
rect 11563 7296 11612 7324
rect 11563 7293 11575 7296
rect 11517 7287 11575 7293
rect 11606 7284 11612 7296
rect 11664 7284 11670 7336
rect 12434 7324 12440 7336
rect 12395 7296 12440 7324
rect 12434 7284 12440 7296
rect 12492 7284 12498 7336
rect 12894 7324 12900 7336
rect 12855 7296 12900 7324
rect 12894 7284 12900 7296
rect 12952 7284 12958 7336
rect 13170 7284 13176 7336
rect 13228 7324 13234 7336
rect 13817 7327 13875 7333
rect 13817 7324 13829 7327
rect 13228 7296 13829 7324
rect 13228 7284 13234 7296
rect 13817 7293 13829 7296
rect 13863 7293 13875 7327
rect 13817 7287 13875 7293
rect 13906 7284 13912 7336
rect 13964 7324 13970 7336
rect 14458 7324 14464 7336
rect 13964 7296 14009 7324
rect 14419 7296 14464 7324
rect 13964 7284 13970 7296
rect 14458 7284 14464 7296
rect 14516 7284 14522 7336
rect 14642 7324 14648 7336
rect 14603 7296 14648 7324
rect 14642 7284 14648 7296
rect 14700 7284 14706 7336
rect 15304 7333 15332 7364
rect 18432 7336 18460 7364
rect 18966 7352 18972 7364
rect 19024 7352 19030 7404
rect 20809 7395 20867 7401
rect 19812 7364 20484 7392
rect 15289 7327 15347 7333
rect 15289 7293 15301 7327
rect 15335 7293 15347 7327
rect 15562 7324 15568 7336
rect 15523 7296 15568 7324
rect 15289 7287 15347 7293
rect 15562 7284 15568 7296
rect 15620 7284 15626 7336
rect 16666 7324 16672 7336
rect 16627 7296 16672 7324
rect 16666 7284 16672 7296
rect 16724 7284 16730 7336
rect 16853 7327 16911 7333
rect 16853 7293 16865 7327
rect 16899 7293 16911 7327
rect 16853 7287 16911 7293
rect 14366 7256 14372 7268
rect 8076 7228 14372 7256
rect 8076 7216 8082 7228
rect 14366 7216 14372 7228
rect 14424 7216 14430 7268
rect 16868 7256 16896 7287
rect 16942 7284 16948 7336
rect 17000 7324 17006 7336
rect 17129 7327 17187 7333
rect 17129 7324 17141 7327
rect 17000 7296 17141 7324
rect 17000 7284 17006 7296
rect 17129 7293 17141 7296
rect 17175 7293 17187 7327
rect 17129 7287 17187 7293
rect 18233 7327 18291 7333
rect 18233 7293 18245 7327
rect 18279 7293 18291 7327
rect 18414 7324 18420 7336
rect 18375 7296 18420 7324
rect 18233 7287 18291 7293
rect 17954 7256 17960 7268
rect 16868 7228 17960 7256
rect 17954 7216 17960 7228
rect 18012 7216 18018 7268
rect 18248 7256 18276 7287
rect 18414 7284 18420 7296
rect 18472 7284 18478 7336
rect 18877 7327 18935 7333
rect 18877 7293 18889 7327
rect 18923 7324 18935 7327
rect 19334 7324 19340 7336
rect 18923 7296 19340 7324
rect 18923 7293 18935 7296
rect 18877 7287 18935 7293
rect 19334 7284 19340 7296
rect 19392 7284 19398 7336
rect 19812 7256 19840 7364
rect 20456 7336 20484 7364
rect 20809 7361 20821 7395
rect 20855 7392 20867 7395
rect 21726 7392 21732 7404
rect 20855 7364 21732 7392
rect 20855 7361 20867 7364
rect 20809 7355 20867 7361
rect 21726 7352 21732 7364
rect 21784 7352 21790 7404
rect 23658 7352 23664 7404
rect 23716 7392 23722 7404
rect 27614 7392 27620 7404
rect 23716 7364 23761 7392
rect 27575 7364 27620 7392
rect 23716 7352 23722 7364
rect 27614 7352 27620 7364
rect 27672 7352 27678 7404
rect 28166 7392 28172 7404
rect 28127 7364 28172 7392
rect 28166 7352 28172 7364
rect 28224 7352 28230 7404
rect 28721 7395 28779 7401
rect 28721 7361 28733 7395
rect 28767 7392 28779 7395
rect 30193 7395 30251 7401
rect 30193 7392 30205 7395
rect 28767 7364 30205 7392
rect 28767 7361 28779 7364
rect 28721 7355 28779 7361
rect 30193 7361 30205 7364
rect 30239 7361 30251 7395
rect 30193 7355 30251 7361
rect 32398 7352 32404 7404
rect 32456 7392 32462 7404
rect 32493 7395 32551 7401
rect 32493 7392 32505 7395
rect 32456 7364 32505 7392
rect 32456 7352 32462 7364
rect 32493 7361 32505 7364
rect 32539 7361 32551 7395
rect 32493 7355 32551 7361
rect 33134 7352 33140 7404
rect 33192 7392 33198 7404
rect 35437 7395 35495 7401
rect 35437 7392 35449 7395
rect 33192 7364 35449 7392
rect 33192 7352 33198 7364
rect 35437 7361 35449 7364
rect 35483 7361 35495 7395
rect 37826 7392 37832 7404
rect 37787 7364 37832 7392
rect 35437 7355 35495 7361
rect 37826 7352 37832 7364
rect 37884 7352 37890 7404
rect 19889 7327 19947 7333
rect 19889 7293 19901 7327
rect 19935 7293 19947 7327
rect 19889 7287 19947 7293
rect 18248 7228 19840 7256
rect 19904 7256 19932 7287
rect 19978 7284 19984 7336
rect 20036 7324 20042 7336
rect 20438 7324 20444 7336
rect 20036 7296 20081 7324
rect 20399 7296 20444 7324
rect 20036 7284 20042 7296
rect 20438 7284 20444 7296
rect 20496 7284 20502 7336
rect 20622 7284 20628 7336
rect 20680 7324 20686 7336
rect 21545 7327 21603 7333
rect 21545 7324 21557 7327
rect 20680 7296 21557 7324
rect 20680 7284 20686 7296
rect 21545 7293 21557 7296
rect 21591 7293 21603 7327
rect 21545 7287 21603 7293
rect 22005 7327 22063 7333
rect 22005 7293 22017 7327
rect 22051 7324 22063 7327
rect 22094 7324 22100 7336
rect 22051 7296 22100 7324
rect 22051 7293 22063 7296
rect 22005 7287 22063 7293
rect 22094 7284 22100 7296
rect 22152 7284 22158 7336
rect 22370 7324 22376 7336
rect 22331 7296 22376 7324
rect 22370 7284 22376 7296
rect 22428 7284 22434 7336
rect 23198 7324 23204 7336
rect 23159 7296 23204 7324
rect 23198 7284 23204 7296
rect 23256 7284 23262 7336
rect 23937 7327 23995 7333
rect 23937 7293 23949 7327
rect 23983 7324 23995 7327
rect 24210 7324 24216 7336
rect 23983 7296 24216 7324
rect 23983 7293 23995 7296
rect 23937 7287 23995 7293
rect 24210 7284 24216 7296
rect 24268 7284 24274 7336
rect 26145 7327 26203 7333
rect 26145 7293 26157 7327
rect 26191 7324 26203 7327
rect 26694 7324 26700 7336
rect 26191 7296 26700 7324
rect 26191 7293 26203 7296
rect 26145 7287 26203 7293
rect 26694 7284 26700 7296
rect 26752 7324 26758 7336
rect 26789 7327 26847 7333
rect 26789 7324 26801 7327
rect 26752 7296 26801 7324
rect 26752 7284 26758 7296
rect 26789 7293 26801 7296
rect 26835 7293 26847 7327
rect 26789 7287 26847 7293
rect 27246 7284 27252 7336
rect 27304 7324 27310 7336
rect 27525 7327 27583 7333
rect 27525 7324 27537 7327
rect 27304 7296 27537 7324
rect 27304 7284 27310 7296
rect 27525 7293 27537 7296
rect 27571 7293 27583 7327
rect 27525 7287 27583 7293
rect 28074 7284 28080 7336
rect 28132 7324 28138 7336
rect 28261 7327 28319 7333
rect 28261 7324 28273 7327
rect 28132 7296 28273 7324
rect 28132 7284 28138 7296
rect 28261 7293 28273 7296
rect 28307 7293 28319 7327
rect 29270 7324 29276 7336
rect 29231 7296 29276 7324
rect 28261 7287 28319 7293
rect 29270 7284 29276 7296
rect 29328 7284 29334 7336
rect 29917 7327 29975 7333
rect 29917 7293 29929 7327
rect 29963 7324 29975 7327
rect 30282 7324 30288 7336
rect 29963 7296 30288 7324
rect 29963 7293 29975 7296
rect 29917 7287 29975 7293
rect 30282 7284 30288 7296
rect 30340 7284 30346 7336
rect 32217 7327 32275 7333
rect 32217 7293 32229 7327
rect 32263 7324 32275 7327
rect 34330 7324 34336 7336
rect 32263 7296 34336 7324
rect 32263 7293 32275 7296
rect 32217 7287 32275 7293
rect 34330 7284 34336 7296
rect 34388 7324 34394 7336
rect 35161 7327 35219 7333
rect 35161 7324 35173 7327
rect 34388 7296 35173 7324
rect 34388 7284 34394 7296
rect 35161 7293 35173 7296
rect 35207 7293 35219 7327
rect 37734 7324 37740 7336
rect 37695 7296 37740 7324
rect 35161 7287 35219 7293
rect 37734 7284 37740 7296
rect 37792 7284 37798 7336
rect 37936 7333 37964 7432
rect 37921 7327 37979 7333
rect 37921 7293 37933 7327
rect 37967 7293 37979 7327
rect 38286 7324 38292 7336
rect 38247 7296 38292 7324
rect 37921 7287 37979 7293
rect 38286 7284 38292 7296
rect 38344 7284 38350 7336
rect 38838 7324 38844 7336
rect 38799 7296 38844 7324
rect 38838 7284 38844 7296
rect 38896 7284 38902 7336
rect 21450 7256 21456 7268
rect 19904 7228 21456 7256
rect 21450 7216 21456 7228
rect 21508 7216 21514 7268
rect 33873 7259 33931 7265
rect 33873 7225 33885 7259
rect 33919 7256 33931 7259
rect 34698 7256 34704 7268
rect 33919 7228 34704 7256
rect 33919 7225 33931 7228
rect 33873 7219 33931 7225
rect 34698 7216 34704 7228
rect 34756 7216 34762 7268
rect 10318 7148 10324 7200
rect 10376 7188 10382 7200
rect 10413 7191 10471 7197
rect 10413 7188 10425 7191
rect 10376 7160 10425 7188
rect 10376 7148 10382 7160
rect 10413 7157 10425 7160
rect 10459 7157 10471 7191
rect 10413 7151 10471 7157
rect 10502 7148 10508 7200
rect 10560 7188 10566 7200
rect 11701 7191 11759 7197
rect 11701 7188 11713 7191
rect 10560 7160 11713 7188
rect 10560 7148 10566 7160
rect 11701 7157 11713 7160
rect 11747 7188 11759 7191
rect 12434 7188 12440 7200
rect 11747 7160 12440 7188
rect 11747 7157 11759 7160
rect 11701 7151 11759 7157
rect 12434 7148 12440 7160
rect 12492 7148 12498 7200
rect 12618 7148 12624 7200
rect 12676 7188 12682 7200
rect 13078 7188 13084 7200
rect 12676 7160 13084 7188
rect 12676 7148 12682 7160
rect 13078 7148 13084 7160
rect 13136 7188 13142 7200
rect 13633 7191 13691 7197
rect 13633 7188 13645 7191
rect 13136 7160 13645 7188
rect 13136 7148 13142 7160
rect 13633 7157 13645 7160
rect 13679 7188 13691 7191
rect 15286 7188 15292 7200
rect 13679 7160 15292 7188
rect 13679 7157 13691 7160
rect 13633 7151 13691 7157
rect 15286 7148 15292 7160
rect 15344 7188 15350 7200
rect 15470 7188 15476 7200
rect 15344 7160 15476 7188
rect 15344 7148 15350 7160
rect 15470 7148 15476 7160
rect 15528 7148 15534 7200
rect 16574 7148 16580 7200
rect 16632 7188 16638 7200
rect 21082 7188 21088 7200
rect 16632 7160 21088 7188
rect 16632 7148 16638 7160
rect 21082 7148 21088 7160
rect 21140 7148 21146 7200
rect 22922 7148 22928 7200
rect 22980 7188 22986 7200
rect 23017 7191 23075 7197
rect 23017 7188 23029 7191
rect 22980 7160 23029 7188
rect 22980 7148 22986 7160
rect 23017 7157 23029 7160
rect 23063 7157 23075 7191
rect 23017 7151 23075 7157
rect 23198 7148 23204 7200
rect 23256 7188 23262 7200
rect 26973 7191 27031 7197
rect 26973 7188 26985 7191
rect 23256 7160 26985 7188
rect 23256 7148 23262 7160
rect 26973 7157 26985 7160
rect 27019 7188 27031 7191
rect 27154 7188 27160 7200
rect 27019 7160 27160 7188
rect 27019 7157 27031 7160
rect 26973 7151 27031 7157
rect 27154 7148 27160 7160
rect 27212 7188 27218 7200
rect 29086 7188 29092 7200
rect 27212 7160 29092 7188
rect 27212 7148 27218 7160
rect 29086 7148 29092 7160
rect 29144 7148 29150 7200
rect 1104 7098 39836 7120
rect 1104 7046 19606 7098
rect 19658 7046 19670 7098
rect 19722 7046 19734 7098
rect 19786 7046 19798 7098
rect 19850 7046 39836 7098
rect 1104 7024 39836 7046
rect 7834 6984 7840 6996
rect 7795 6956 7840 6984
rect 7834 6944 7840 6956
rect 7892 6944 7898 6996
rect 9953 6987 10011 6993
rect 9953 6953 9965 6987
rect 9999 6984 10011 6987
rect 10226 6984 10232 6996
rect 9999 6956 10232 6984
rect 9999 6953 10011 6956
rect 9953 6947 10011 6953
rect 10226 6944 10232 6956
rect 10284 6944 10290 6996
rect 18138 6944 18144 6996
rect 18196 6944 18202 6996
rect 18230 6944 18236 6996
rect 18288 6984 18294 6996
rect 29270 6984 29276 6996
rect 18288 6956 24532 6984
rect 29231 6956 29276 6984
rect 18288 6944 18294 6956
rect 5166 6876 5172 6928
rect 5224 6916 5230 6928
rect 5224 6888 5488 6916
rect 5224 6876 5230 6888
rect 2406 6848 2412 6860
rect 2367 6820 2412 6848
rect 2406 6808 2412 6820
rect 2464 6808 2470 6860
rect 2498 6808 2504 6860
rect 2556 6848 2562 6860
rect 2961 6851 3019 6857
rect 2961 6848 2973 6851
rect 2556 6820 2973 6848
rect 2556 6808 2562 6820
rect 2961 6817 2973 6820
rect 3007 6817 3019 6851
rect 2961 6811 3019 6817
rect 3145 6851 3203 6857
rect 3145 6817 3157 6851
rect 3191 6848 3203 6851
rect 3602 6848 3608 6860
rect 3191 6820 3608 6848
rect 3191 6817 3203 6820
rect 3145 6811 3203 6817
rect 3602 6808 3608 6820
rect 3660 6808 3666 6860
rect 5074 6848 5080 6860
rect 5035 6820 5080 6848
rect 5074 6808 5080 6820
rect 5132 6808 5138 6860
rect 5261 6851 5319 6857
rect 5261 6817 5273 6851
rect 5307 6848 5319 6851
rect 5350 6848 5356 6860
rect 5307 6820 5356 6848
rect 5307 6817 5319 6820
rect 5261 6811 5319 6817
rect 5350 6808 5356 6820
rect 5408 6808 5414 6860
rect 5460 6857 5488 6888
rect 11900 6888 13032 6916
rect 5445 6851 5503 6857
rect 5445 6817 5457 6851
rect 5491 6817 5503 6851
rect 5445 6811 5503 6817
rect 6549 6851 6607 6857
rect 6549 6817 6561 6851
rect 6595 6848 6607 6851
rect 7282 6848 7288 6860
rect 6595 6820 7288 6848
rect 6595 6817 6607 6820
rect 6549 6811 6607 6817
rect 7282 6808 7288 6820
rect 7340 6808 7346 6860
rect 8941 6851 8999 6857
rect 8941 6817 8953 6851
rect 8987 6848 8999 6851
rect 9490 6848 9496 6860
rect 8987 6820 9496 6848
rect 8987 6817 8999 6820
rect 8941 6811 8999 6817
rect 9490 6808 9496 6820
rect 9548 6808 9554 6860
rect 9953 6851 10011 6857
rect 9953 6817 9965 6851
rect 9999 6848 10011 6851
rect 10134 6848 10140 6860
rect 9999 6820 10140 6848
rect 9999 6817 10011 6820
rect 9953 6811 10011 6817
rect 10134 6808 10140 6820
rect 10192 6808 10198 6860
rect 10229 6851 10287 6857
rect 10229 6817 10241 6851
rect 10275 6848 10287 6851
rect 10275 6820 10364 6848
rect 10275 6817 10287 6820
rect 10229 6811 10287 6817
rect 4614 6780 4620 6792
rect 4575 6752 4620 6780
rect 4614 6740 4620 6752
rect 4672 6740 4678 6792
rect 4706 6740 4712 6792
rect 4764 6780 4770 6792
rect 6270 6780 6276 6792
rect 4764 6752 6276 6780
rect 4764 6740 4770 6752
rect 6270 6740 6276 6752
rect 6328 6740 6334 6792
rect 10336 6724 10364 6820
rect 10502 6808 10508 6860
rect 10560 6848 10566 6860
rect 11425 6851 11483 6857
rect 11425 6848 11437 6851
rect 10560 6820 11437 6848
rect 10560 6808 10566 6820
rect 11425 6817 11437 6820
rect 11471 6817 11483 6851
rect 11425 6811 11483 6817
rect 11517 6851 11575 6857
rect 11517 6817 11529 6851
rect 11563 6848 11575 6851
rect 11900 6848 11928 6888
rect 11563 6820 11928 6848
rect 11977 6851 12035 6857
rect 11563 6817 11575 6820
rect 11517 6811 11575 6817
rect 11977 6817 11989 6851
rect 12023 6848 12035 6851
rect 12066 6848 12072 6860
rect 12023 6820 12072 6848
rect 12023 6817 12035 6820
rect 11977 6811 12035 6817
rect 12066 6808 12072 6820
rect 12124 6808 12130 6860
rect 12161 6851 12219 6857
rect 12161 6817 12173 6851
rect 12207 6848 12219 6851
rect 12894 6848 12900 6860
rect 12207 6820 12900 6848
rect 12207 6817 12219 6820
rect 12161 6811 12219 6817
rect 12894 6808 12900 6820
rect 12952 6808 12958 6860
rect 13004 6848 13032 6888
rect 14458 6876 14464 6928
rect 14516 6916 14522 6928
rect 15381 6919 15439 6925
rect 15381 6916 15393 6919
rect 14516 6888 15393 6916
rect 14516 6876 14522 6888
rect 15381 6885 15393 6888
rect 15427 6885 15439 6919
rect 18156 6916 18184 6944
rect 24504 6928 24532 6956
rect 29270 6944 29276 6956
rect 29328 6944 29334 6996
rect 23198 6916 23204 6928
rect 18156 6888 23204 6916
rect 15381 6879 15439 6885
rect 13357 6851 13415 6857
rect 13004 6820 13308 6848
rect 13078 6780 13084 6792
rect 13039 6752 13084 6780
rect 13078 6740 13084 6752
rect 13136 6740 13142 6792
rect 13280 6780 13308 6820
rect 13357 6817 13369 6851
rect 13403 6848 13415 6851
rect 13998 6848 14004 6860
rect 13403 6820 14004 6848
rect 13403 6817 13415 6820
rect 13357 6811 13415 6817
rect 13998 6808 14004 6820
rect 14056 6808 14062 6860
rect 14737 6851 14795 6857
rect 14737 6817 14749 6851
rect 14783 6848 14795 6851
rect 15289 6851 15347 6857
rect 15289 6848 15301 6851
rect 14783 6820 15301 6848
rect 14783 6817 14795 6820
rect 14737 6811 14795 6817
rect 15289 6817 15301 6820
rect 15335 6817 15347 6851
rect 15289 6811 15347 6817
rect 15470 6808 15476 6860
rect 15528 6848 15534 6860
rect 16485 6851 16543 6857
rect 16485 6848 16497 6851
rect 15528 6820 16497 6848
rect 15528 6808 15534 6820
rect 16485 6817 16497 6820
rect 16531 6817 16543 6851
rect 16485 6811 16543 6817
rect 16761 6851 16819 6857
rect 16761 6817 16773 6851
rect 16807 6848 16819 6851
rect 17494 6848 17500 6860
rect 16807 6820 17500 6848
rect 16807 6817 16819 6820
rect 16761 6811 16819 6817
rect 17494 6808 17500 6820
rect 17552 6808 17558 6860
rect 18141 6851 18199 6857
rect 18141 6817 18153 6851
rect 18187 6848 18199 6851
rect 18322 6848 18328 6860
rect 18187 6820 18328 6848
rect 18187 6817 18199 6820
rect 18141 6811 18199 6817
rect 18322 6808 18328 6820
rect 18380 6808 18386 6860
rect 19429 6851 19487 6857
rect 19429 6817 19441 6851
rect 19475 6817 19487 6851
rect 19429 6811 19487 6817
rect 19797 6851 19855 6857
rect 19797 6817 19809 6851
rect 19843 6848 19855 6851
rect 19978 6848 19984 6860
rect 19843 6820 19984 6848
rect 19843 6817 19855 6820
rect 19797 6811 19855 6817
rect 18230 6780 18236 6792
rect 13280 6752 14320 6780
rect 2958 6712 2964 6724
rect 2919 6684 2964 6712
rect 2958 6672 2964 6684
rect 3016 6672 3022 6724
rect 9033 6715 9091 6721
rect 9033 6681 9045 6715
rect 9079 6712 9091 6715
rect 10318 6712 10324 6724
rect 9079 6684 10324 6712
rect 9079 6681 9091 6684
rect 9033 6675 9091 6681
rect 10318 6672 10324 6684
rect 10376 6672 10382 6724
rect 12066 6672 12072 6724
rect 12124 6712 12130 6724
rect 14292 6712 14320 6752
rect 16500 6752 18236 6780
rect 16500 6712 16528 6752
rect 18230 6740 18236 6752
rect 18288 6740 18294 6792
rect 19334 6780 19340 6792
rect 19295 6752 19340 6780
rect 19334 6740 19340 6752
rect 19392 6740 19398 6792
rect 19444 6780 19472 6811
rect 19978 6808 19984 6820
rect 20036 6808 20042 6860
rect 20165 6851 20223 6857
rect 20165 6817 20177 6851
rect 20211 6848 20223 6851
rect 20438 6848 20444 6860
rect 20211 6820 20444 6848
rect 20211 6817 20223 6820
rect 20165 6811 20223 6817
rect 20438 6808 20444 6820
rect 20496 6808 20502 6860
rect 21082 6848 21088 6860
rect 21043 6820 21088 6848
rect 21082 6808 21088 6820
rect 21140 6808 21146 6860
rect 21453 6851 21511 6857
rect 21453 6848 21465 6851
rect 21376 6820 21465 6848
rect 20070 6780 20076 6792
rect 19444 6752 20076 6780
rect 20070 6740 20076 6752
rect 20128 6740 20134 6792
rect 21266 6780 21272 6792
rect 21227 6752 21272 6780
rect 21266 6740 21272 6752
rect 21324 6740 21330 6792
rect 12124 6684 12572 6712
rect 14292 6684 16528 6712
rect 12124 6672 12130 6684
rect 11974 6604 11980 6656
rect 12032 6644 12038 6656
rect 12437 6647 12495 6653
rect 12437 6644 12449 6647
rect 12032 6616 12449 6644
rect 12032 6604 12038 6616
rect 12437 6613 12449 6616
rect 12483 6613 12495 6647
rect 12544 6644 12572 6684
rect 20898 6672 20904 6724
rect 20956 6712 20962 6724
rect 21376 6712 21404 6820
rect 21453 6817 21465 6820
rect 21499 6817 21511 6851
rect 21453 6811 21511 6817
rect 22005 6851 22063 6857
rect 22005 6817 22017 6851
rect 22051 6848 22063 6851
rect 22094 6848 22100 6860
rect 22051 6820 22100 6848
rect 22051 6817 22063 6820
rect 22005 6811 22063 6817
rect 22094 6808 22100 6820
rect 22152 6808 22158 6860
rect 22848 6857 22876 6888
rect 23198 6876 23204 6888
rect 23256 6876 23262 6928
rect 24121 6919 24179 6925
rect 23676 6888 23980 6916
rect 22833 6851 22891 6857
rect 22833 6817 22845 6851
rect 22879 6817 22891 6851
rect 22833 6811 22891 6817
rect 23017 6851 23075 6857
rect 23017 6817 23029 6851
rect 23063 6848 23075 6851
rect 23474 6848 23480 6860
rect 23063 6820 23480 6848
rect 23063 6817 23075 6820
rect 23017 6811 23075 6817
rect 23474 6808 23480 6820
rect 23532 6808 23538 6860
rect 23569 6851 23627 6857
rect 23569 6817 23581 6851
rect 23615 6848 23627 6851
rect 23676 6848 23704 6888
rect 23615 6820 23704 6848
rect 23615 6817 23627 6820
rect 23569 6811 23627 6817
rect 23750 6808 23756 6860
rect 23808 6848 23814 6860
rect 23808 6820 23853 6848
rect 23808 6808 23814 6820
rect 23952 6780 23980 6888
rect 24121 6885 24133 6919
rect 24167 6916 24179 6919
rect 24210 6916 24216 6928
rect 24167 6888 24216 6916
rect 24167 6885 24179 6888
rect 24121 6879 24179 6885
rect 24210 6876 24216 6888
rect 24268 6876 24274 6928
rect 24486 6876 24492 6928
rect 24544 6916 24550 6928
rect 26786 6916 26792 6928
rect 24544 6888 26792 6916
rect 24544 6876 24550 6888
rect 26786 6876 26792 6888
rect 26844 6876 26850 6928
rect 30668 6888 35204 6916
rect 24578 6808 24584 6860
rect 24636 6848 24642 6860
rect 24673 6851 24731 6857
rect 24673 6848 24685 6851
rect 24636 6820 24685 6848
rect 24636 6808 24642 6820
rect 24673 6817 24685 6820
rect 24719 6817 24731 6851
rect 24673 6811 24731 6817
rect 24762 6808 24768 6860
rect 24820 6848 24826 6860
rect 25409 6851 25467 6857
rect 25409 6848 25421 6851
rect 24820 6820 25421 6848
rect 24820 6808 24826 6820
rect 25409 6817 25421 6820
rect 25455 6817 25467 6851
rect 25409 6811 25467 6817
rect 26973 6851 27031 6857
rect 26973 6817 26985 6851
rect 27019 6848 27031 6851
rect 27246 6848 27252 6860
rect 27019 6820 27252 6848
rect 27019 6817 27031 6820
rect 26973 6811 27031 6817
rect 27246 6808 27252 6820
rect 27304 6808 27310 6860
rect 30668 6857 30696 6888
rect 30653 6851 30711 6857
rect 30653 6817 30665 6851
rect 30699 6817 30711 6851
rect 31478 6848 31484 6860
rect 31439 6820 31484 6848
rect 30653 6811 30711 6817
rect 31478 6808 31484 6820
rect 31536 6808 31542 6860
rect 32309 6851 32367 6857
rect 32309 6817 32321 6851
rect 32355 6848 32367 6851
rect 32582 6848 32588 6860
rect 32355 6820 32588 6848
rect 32355 6817 32367 6820
rect 32309 6811 32367 6817
rect 32582 6808 32588 6820
rect 32640 6808 32646 6860
rect 33226 6808 33232 6860
rect 33284 6848 33290 6860
rect 33505 6851 33563 6857
rect 33505 6848 33517 6851
rect 33284 6820 33517 6848
rect 33284 6808 33290 6820
rect 33505 6817 33517 6820
rect 33551 6817 33563 6851
rect 33505 6811 33563 6817
rect 33781 6851 33839 6857
rect 33781 6817 33793 6851
rect 33827 6848 33839 6851
rect 34606 6848 34612 6860
rect 33827 6820 34612 6848
rect 33827 6817 33839 6820
rect 33781 6811 33839 6817
rect 34606 6808 34612 6820
rect 34664 6808 34670 6860
rect 25314 6780 25320 6792
rect 23952 6752 25320 6780
rect 25314 6740 25320 6752
rect 25372 6740 25378 6792
rect 27430 6740 27436 6792
rect 27488 6780 27494 6792
rect 27709 6783 27767 6789
rect 27709 6780 27721 6783
rect 27488 6752 27721 6780
rect 27488 6740 27494 6752
rect 27709 6749 27721 6752
rect 27755 6780 27767 6783
rect 27890 6780 27896 6792
rect 27755 6752 27896 6780
rect 27755 6749 27767 6752
rect 27709 6743 27767 6749
rect 27890 6740 27896 6752
rect 27948 6740 27954 6792
rect 27985 6783 28043 6789
rect 27985 6749 27997 6783
rect 28031 6780 28043 6783
rect 29825 6783 29883 6789
rect 29825 6780 29837 6783
rect 28031 6752 29837 6780
rect 28031 6749 28043 6752
rect 27985 6743 28043 6749
rect 29825 6749 29837 6752
rect 29871 6749 29883 6783
rect 29825 6743 29883 6749
rect 29914 6740 29920 6792
rect 29972 6780 29978 6792
rect 30377 6783 30435 6789
rect 30377 6780 30389 6783
rect 29972 6752 30389 6780
rect 29972 6740 29978 6752
rect 30377 6749 30389 6752
rect 30423 6749 30435 6783
rect 30834 6780 30840 6792
rect 30795 6752 30840 6780
rect 30377 6743 30435 6749
rect 30834 6740 30840 6752
rect 30892 6740 30898 6792
rect 32953 6783 33011 6789
rect 32953 6749 32965 6783
rect 32999 6780 33011 6783
rect 33962 6780 33968 6792
rect 32999 6752 33456 6780
rect 33923 6752 33968 6780
rect 32999 6749 33011 6752
rect 32953 6743 33011 6749
rect 20956 6684 21404 6712
rect 20956 6672 20962 6684
rect 24670 6672 24676 6724
rect 24728 6712 24734 6724
rect 32401 6715 32459 6721
rect 24728 6684 27200 6712
rect 24728 6672 24734 6684
rect 16758 6644 16764 6656
rect 12544 6616 16764 6644
rect 12437 6607 12495 6613
rect 16758 6604 16764 6616
rect 16816 6604 16822 6656
rect 22186 6604 22192 6656
rect 22244 6644 22250 6656
rect 24762 6644 24768 6656
rect 22244 6616 24768 6644
rect 22244 6604 22250 6616
rect 24762 6604 24768 6616
rect 24820 6604 24826 6656
rect 24857 6647 24915 6653
rect 24857 6613 24869 6647
rect 24903 6644 24915 6647
rect 25038 6644 25044 6656
rect 24903 6616 25044 6644
rect 24903 6613 24915 6616
rect 24857 6607 24915 6613
rect 25038 6604 25044 6616
rect 25096 6604 25102 6656
rect 25593 6647 25651 6653
rect 25593 6613 25605 6647
rect 25639 6644 25651 6647
rect 26234 6644 26240 6656
rect 25639 6616 26240 6644
rect 25639 6613 25651 6616
rect 25593 6607 25651 6613
rect 26234 6604 26240 6616
rect 26292 6604 26298 6656
rect 27172 6653 27200 6684
rect 32401 6681 32413 6715
rect 32447 6712 32459 6715
rect 33134 6712 33140 6724
rect 32447 6684 33140 6712
rect 32447 6681 32459 6684
rect 32401 6675 32459 6681
rect 33134 6672 33140 6684
rect 33192 6672 33198 6724
rect 33428 6712 33456 6752
rect 33962 6740 33968 6752
rect 34020 6740 34026 6792
rect 34422 6780 34428 6792
rect 34383 6752 34428 6780
rect 34422 6740 34428 6752
rect 34480 6740 34486 6792
rect 34977 6783 35035 6789
rect 34977 6749 34989 6783
rect 35023 6749 35035 6783
rect 35176 6780 35204 6888
rect 35253 6851 35311 6857
rect 35253 6817 35265 6851
rect 35299 6848 35311 6851
rect 36262 6848 36268 6860
rect 35299 6820 36268 6848
rect 35299 6817 35311 6820
rect 35253 6811 35311 6817
rect 36262 6808 36268 6820
rect 36320 6848 36326 6860
rect 36722 6848 36728 6860
rect 36320 6820 36584 6848
rect 36683 6820 36728 6848
rect 36320 6808 36326 6820
rect 35434 6780 35440 6792
rect 35176 6752 35440 6780
rect 34977 6743 35035 6749
rect 34992 6712 35020 6743
rect 35434 6740 35440 6752
rect 35492 6740 35498 6792
rect 35894 6780 35900 6792
rect 35855 6752 35900 6780
rect 35894 6740 35900 6752
rect 35952 6740 35958 6792
rect 36170 6740 36176 6792
rect 36228 6780 36234 6792
rect 36449 6783 36507 6789
rect 36449 6780 36461 6783
rect 36228 6752 36461 6780
rect 36228 6740 36234 6752
rect 36449 6749 36461 6752
rect 36495 6749 36507 6783
rect 36556 6780 36584 6820
rect 36722 6808 36728 6820
rect 36780 6808 36786 6860
rect 38010 6848 38016 6860
rect 37971 6820 38016 6848
rect 38010 6808 38016 6820
rect 38068 6808 38074 6860
rect 38378 6848 38384 6860
rect 38339 6820 38384 6848
rect 38378 6808 38384 6820
rect 38436 6808 38442 6860
rect 38470 6808 38476 6860
rect 38528 6848 38534 6860
rect 38657 6851 38715 6857
rect 38657 6848 38669 6851
rect 38528 6820 38669 6848
rect 38528 6808 38534 6820
rect 38657 6817 38669 6820
rect 38703 6817 38715 6851
rect 38657 6811 38715 6817
rect 36909 6783 36967 6789
rect 36909 6780 36921 6783
rect 36556 6752 36921 6780
rect 36449 6743 36507 6749
rect 36909 6749 36921 6752
rect 36955 6749 36967 6783
rect 36909 6743 36967 6749
rect 33428 6684 35020 6712
rect 37734 6672 37740 6724
rect 37792 6712 37798 6724
rect 37921 6715 37979 6721
rect 37921 6712 37933 6715
rect 37792 6684 37933 6712
rect 37792 6672 37798 6684
rect 37921 6681 37933 6684
rect 37967 6681 37979 6715
rect 37921 6675 37979 6681
rect 27157 6647 27215 6653
rect 27157 6613 27169 6647
rect 27203 6644 27215 6647
rect 27338 6644 27344 6656
rect 27203 6616 27344 6644
rect 27203 6613 27215 6616
rect 27157 6607 27215 6613
rect 27338 6604 27344 6616
rect 27396 6604 27402 6656
rect 28166 6604 28172 6656
rect 28224 6644 28230 6656
rect 31202 6644 31208 6656
rect 28224 6616 31208 6644
rect 28224 6604 28230 6616
rect 31202 6604 31208 6616
rect 31260 6604 31266 6656
rect 31297 6647 31355 6653
rect 31297 6613 31309 6647
rect 31343 6644 31355 6647
rect 31386 6644 31392 6656
rect 31343 6616 31392 6644
rect 31343 6613 31355 6616
rect 31297 6607 31355 6613
rect 31386 6604 31392 6616
rect 31444 6644 31450 6656
rect 32306 6644 32312 6656
rect 31444 6616 32312 6644
rect 31444 6604 31450 6616
rect 32306 6604 32312 6616
rect 32364 6604 32370 6656
rect 1104 6554 39836 6576
rect 1104 6502 4246 6554
rect 4298 6502 4310 6554
rect 4362 6502 4374 6554
rect 4426 6502 4438 6554
rect 4490 6502 34966 6554
rect 35018 6502 35030 6554
rect 35082 6502 35094 6554
rect 35146 6502 35158 6554
rect 35210 6502 39836 6554
rect 1104 6480 39836 6502
rect 5074 6440 5080 6452
rect 4632 6412 5080 6440
rect 3602 6332 3608 6384
rect 3660 6372 3666 6384
rect 3789 6375 3847 6381
rect 3789 6372 3801 6375
rect 3660 6344 3801 6372
rect 3660 6332 3666 6344
rect 3789 6341 3801 6344
rect 3835 6341 3847 6375
rect 3789 6335 3847 6341
rect 2406 6304 2412 6316
rect 2148 6276 2412 6304
rect 2148 6245 2176 6276
rect 2406 6264 2412 6276
rect 2464 6264 2470 6316
rect 2593 6307 2651 6313
rect 2593 6273 2605 6307
rect 2639 6304 2651 6307
rect 3973 6307 4031 6313
rect 2639 6276 3832 6304
rect 2639 6273 2651 6276
rect 2593 6267 2651 6273
rect 2133 6239 2191 6245
rect 2133 6205 2145 6239
rect 2179 6205 2191 6239
rect 2133 6199 2191 6205
rect 2317 6239 2375 6245
rect 2317 6205 2329 6239
rect 2363 6205 2375 6239
rect 3326 6236 3332 6248
rect 3287 6208 3332 6236
rect 2317 6199 2375 6205
rect 2332 6168 2360 6199
rect 3326 6196 3332 6208
rect 3384 6196 3390 6248
rect 3602 6168 3608 6180
rect 2332 6140 3608 6168
rect 3602 6128 3608 6140
rect 3660 6128 3666 6180
rect 3804 6168 3832 6276
rect 3973 6273 3985 6307
rect 4019 6304 4031 6307
rect 4632 6304 4660 6412
rect 5074 6400 5080 6412
rect 5132 6440 5138 6452
rect 5997 6443 6055 6449
rect 5997 6440 6009 6443
rect 5132 6412 6009 6440
rect 5132 6400 5138 6412
rect 5997 6409 6009 6412
rect 6043 6409 6055 6443
rect 9490 6440 9496 6452
rect 9451 6412 9496 6440
rect 5997 6403 6055 6409
rect 9490 6400 9496 6412
rect 9548 6400 9554 6452
rect 13538 6440 13544 6452
rect 13499 6412 13544 6440
rect 13538 6400 13544 6412
rect 13596 6400 13602 6452
rect 14090 6400 14096 6452
rect 14148 6440 14154 6452
rect 14918 6440 14924 6452
rect 14148 6412 14924 6440
rect 14148 6400 14154 6412
rect 14918 6400 14924 6412
rect 14976 6400 14982 6452
rect 15838 6400 15844 6452
rect 15896 6440 15902 6452
rect 20070 6440 20076 6452
rect 15896 6412 19932 6440
rect 20031 6412 20076 6440
rect 15896 6400 15902 6412
rect 11606 6332 11612 6384
rect 11664 6372 11670 6384
rect 16666 6372 16672 6384
rect 11664 6344 16528 6372
rect 16627 6344 16672 6372
rect 11664 6332 11670 6344
rect 4019 6276 4660 6304
rect 4019 6273 4031 6276
rect 3973 6267 4031 6273
rect 6270 6264 6276 6316
rect 6328 6304 6334 6316
rect 7929 6307 7987 6313
rect 7929 6304 7941 6307
rect 6328 6276 7941 6304
rect 6328 6264 6334 6276
rect 7929 6273 7941 6276
rect 7975 6304 7987 6307
rect 8294 6304 8300 6316
rect 7975 6276 8300 6304
rect 7975 6273 7987 6276
rect 7929 6267 7987 6273
rect 8294 6264 8300 6276
rect 8352 6304 8358 6316
rect 8570 6304 8576 6316
rect 8352 6276 8576 6304
rect 8352 6264 8358 6276
rect 8570 6264 8576 6276
rect 8628 6304 8634 6316
rect 10229 6307 10287 6313
rect 10229 6304 10241 6307
rect 8628 6276 10241 6304
rect 8628 6264 8634 6276
rect 10229 6273 10241 6276
rect 10275 6273 10287 6307
rect 14274 6304 14280 6316
rect 14235 6276 14280 6304
rect 10229 6267 10287 6273
rect 14274 6264 14280 6276
rect 14332 6264 14338 6316
rect 3881 6239 3939 6245
rect 3881 6205 3893 6239
rect 3927 6236 3939 6239
rect 4154 6236 4160 6248
rect 3927 6208 4160 6236
rect 3927 6205 3939 6208
rect 3881 6199 3939 6205
rect 4154 6196 4160 6208
rect 4212 6196 4218 6248
rect 4617 6239 4675 6245
rect 4617 6205 4629 6239
rect 4663 6205 4675 6239
rect 4890 6236 4896 6248
rect 4851 6208 4896 6236
rect 4617 6199 4675 6205
rect 4522 6168 4528 6180
rect 3804 6140 4528 6168
rect 4522 6128 4528 6140
rect 4580 6128 4586 6180
rect 3142 6060 3148 6112
rect 3200 6100 3206 6112
rect 3786 6100 3792 6112
rect 3200 6072 3792 6100
rect 3200 6060 3206 6072
rect 3786 6060 3792 6072
rect 3844 6100 3850 6112
rect 4632 6100 4660 6199
rect 4890 6196 4896 6208
rect 4948 6196 4954 6248
rect 8202 6236 8208 6248
rect 8163 6208 8208 6236
rect 8202 6196 8208 6208
rect 8260 6196 8266 6248
rect 10505 6239 10563 6245
rect 10505 6205 10517 6239
rect 10551 6236 10563 6239
rect 11422 6236 11428 6248
rect 10551 6208 11428 6236
rect 10551 6205 10563 6208
rect 10505 6199 10563 6205
rect 11422 6196 11428 6208
rect 11480 6196 11486 6248
rect 11885 6239 11943 6245
rect 11885 6205 11897 6239
rect 11931 6236 11943 6239
rect 12437 6239 12495 6245
rect 12437 6236 12449 6239
rect 11931 6208 12449 6236
rect 11931 6205 11943 6208
rect 11885 6199 11943 6205
rect 12437 6205 12449 6208
rect 12483 6236 12495 6239
rect 13262 6236 13268 6248
rect 12483 6208 13268 6236
rect 12483 6205 12495 6208
rect 12437 6199 12495 6205
rect 13262 6196 13268 6208
rect 13320 6196 13326 6248
rect 13449 6239 13507 6245
rect 13449 6205 13461 6239
rect 13495 6236 13507 6239
rect 13814 6236 13820 6248
rect 13495 6208 13820 6236
rect 13495 6205 13507 6208
rect 13449 6199 13507 6205
rect 13814 6196 13820 6208
rect 13872 6196 13878 6248
rect 13906 6196 13912 6248
rect 13964 6236 13970 6248
rect 14093 6239 14151 6245
rect 14093 6236 14105 6239
rect 13964 6208 14105 6236
rect 13964 6196 13970 6208
rect 14093 6205 14105 6208
rect 14139 6205 14151 6239
rect 14550 6236 14556 6248
rect 14511 6208 14556 6236
rect 14093 6199 14151 6205
rect 14550 6196 14556 6208
rect 14608 6196 14614 6248
rect 14642 6196 14648 6248
rect 14700 6236 14706 6248
rect 14829 6239 14887 6245
rect 14829 6236 14841 6239
rect 14700 6208 14841 6236
rect 14700 6196 14706 6208
rect 14829 6205 14841 6208
rect 14875 6205 14887 6239
rect 14829 6199 14887 6205
rect 15473 6239 15531 6245
rect 15473 6205 15485 6239
rect 15519 6205 15531 6239
rect 15473 6199 15531 6205
rect 15488 6168 15516 6199
rect 15562 6196 15568 6248
rect 15620 6236 15626 6248
rect 16500 6245 16528 6344
rect 16666 6332 16672 6344
rect 16724 6332 16730 6384
rect 18966 6304 18972 6316
rect 16592 6276 17356 6304
rect 15749 6239 15807 6245
rect 15749 6236 15761 6239
rect 15620 6208 15761 6236
rect 15620 6196 15626 6208
rect 15749 6205 15761 6208
rect 15795 6205 15807 6239
rect 15749 6199 15807 6205
rect 16485 6239 16543 6245
rect 16485 6205 16497 6239
rect 16531 6205 16543 6239
rect 16485 6199 16543 6205
rect 16592 6168 16620 6276
rect 16850 6196 16856 6248
rect 16908 6236 16914 6248
rect 17221 6239 17279 6245
rect 17221 6236 17233 6239
rect 16908 6208 17233 6236
rect 16908 6196 16914 6208
rect 17221 6205 17233 6208
rect 17267 6205 17279 6239
rect 17328 6236 17356 6276
rect 17512 6276 18828 6304
rect 18927 6276 18972 6304
rect 17512 6236 17540 6276
rect 18046 6236 18052 6248
rect 17328 6208 17540 6236
rect 18007 6208 18052 6236
rect 17221 6199 17279 6205
rect 18046 6196 18052 6208
rect 18104 6196 18110 6248
rect 18506 6196 18512 6248
rect 18564 6236 18570 6248
rect 18693 6239 18751 6245
rect 18693 6236 18705 6239
rect 18564 6208 18705 6236
rect 18564 6196 18570 6208
rect 18693 6205 18705 6208
rect 18739 6205 18751 6239
rect 18800 6236 18828 6276
rect 18966 6264 18972 6276
rect 19024 6264 19030 6316
rect 19904 6304 19932 6412
rect 20070 6400 20076 6412
rect 20128 6400 20134 6452
rect 20714 6400 20720 6452
rect 20772 6440 20778 6452
rect 20901 6443 20959 6449
rect 20901 6440 20913 6443
rect 20772 6412 20913 6440
rect 20772 6400 20778 6412
rect 20901 6409 20913 6412
rect 20947 6409 20959 6443
rect 20901 6403 20959 6409
rect 23017 6443 23075 6449
rect 23017 6409 23029 6443
rect 23063 6440 23075 6443
rect 23382 6440 23388 6452
rect 23063 6412 23388 6440
rect 23063 6409 23075 6412
rect 23017 6403 23075 6409
rect 23382 6400 23388 6412
rect 23440 6400 23446 6452
rect 23658 6400 23664 6452
rect 23716 6440 23722 6452
rect 26694 6440 26700 6452
rect 23716 6412 25176 6440
rect 26655 6412 26700 6440
rect 23716 6400 23722 6412
rect 24670 6372 24676 6384
rect 20824 6344 24676 6372
rect 20824 6304 20852 6344
rect 24670 6332 24676 6344
rect 24728 6332 24734 6384
rect 24578 6304 24584 6316
rect 19904 6276 20852 6304
rect 20346 6236 20352 6248
rect 18800 6208 20352 6236
rect 18693 6199 18751 6205
rect 20346 6196 20352 6208
rect 20404 6196 20410 6248
rect 20824 6245 20852 6276
rect 22940 6276 24584 6304
rect 20809 6239 20867 6245
rect 20809 6205 20821 6239
rect 20855 6205 20867 6239
rect 20809 6199 20867 6205
rect 20898 6196 20904 6248
rect 20956 6236 20962 6248
rect 21177 6239 21235 6245
rect 21177 6236 21189 6239
rect 20956 6208 21189 6236
rect 20956 6196 20962 6208
rect 21177 6205 21189 6208
rect 21223 6236 21235 6239
rect 21266 6236 21272 6248
rect 21223 6208 21272 6236
rect 21223 6205 21235 6208
rect 21177 6199 21235 6205
rect 21266 6196 21272 6208
rect 21324 6196 21330 6248
rect 21821 6239 21879 6245
rect 21821 6205 21833 6239
rect 21867 6236 21879 6239
rect 22186 6236 22192 6248
rect 21867 6208 22192 6236
rect 21867 6205 21879 6208
rect 21821 6199 21879 6205
rect 22186 6196 22192 6208
rect 22244 6196 22250 6248
rect 22940 6245 22968 6276
rect 24578 6264 24584 6276
rect 24636 6264 24642 6316
rect 25038 6304 25044 6316
rect 24688 6276 25044 6304
rect 22925 6239 22983 6245
rect 22925 6205 22937 6239
rect 22971 6205 22983 6239
rect 24394 6236 24400 6248
rect 24355 6208 24400 6236
rect 22925 6199 22983 6205
rect 24394 6196 24400 6208
rect 24452 6196 24458 6248
rect 24688 6245 24716 6276
rect 25038 6264 25044 6276
rect 25096 6264 25102 6316
rect 25148 6304 25176 6412
rect 26694 6400 26700 6412
rect 26752 6400 26758 6452
rect 31478 6440 31484 6452
rect 30024 6412 31484 6440
rect 27430 6372 27436 6384
rect 27343 6344 27436 6372
rect 27430 6332 27436 6344
rect 27488 6332 27494 6384
rect 30024 6381 30052 6412
rect 31478 6400 31484 6412
rect 31536 6400 31542 6452
rect 31665 6443 31723 6449
rect 31665 6440 31677 6443
rect 31588 6412 31677 6440
rect 30009 6375 30067 6381
rect 30009 6372 30021 6375
rect 27632 6344 30021 6372
rect 25317 6307 25375 6313
rect 25317 6304 25329 6307
rect 25148 6276 25329 6304
rect 25317 6273 25329 6276
rect 25363 6304 25375 6307
rect 25774 6304 25780 6316
rect 25363 6276 25780 6304
rect 25363 6273 25375 6276
rect 25317 6267 25375 6273
rect 25774 6264 25780 6276
rect 25832 6304 25838 6316
rect 27448 6304 27476 6332
rect 25832 6276 27476 6304
rect 25832 6264 25838 6276
rect 24673 6239 24731 6245
rect 24673 6205 24685 6239
rect 24719 6205 24731 6239
rect 24673 6199 24731 6205
rect 24762 6196 24768 6248
rect 24820 6236 24826 6248
rect 24857 6239 24915 6245
rect 24857 6236 24869 6239
rect 24820 6208 24869 6236
rect 24820 6196 24826 6208
rect 24857 6205 24869 6208
rect 24903 6205 24915 6239
rect 25590 6236 25596 6248
rect 25551 6208 25596 6236
rect 24857 6199 24915 6205
rect 25590 6196 25596 6208
rect 25648 6196 25654 6248
rect 26234 6196 26240 6248
rect 26292 6196 26298 6248
rect 27632 6245 27660 6344
rect 30009 6341 30021 6344
rect 30055 6341 30067 6375
rect 30009 6335 30067 6341
rect 31294 6332 31300 6384
rect 31352 6372 31358 6384
rect 31588 6372 31616 6412
rect 31665 6409 31677 6412
rect 31711 6409 31723 6443
rect 31665 6403 31723 6409
rect 32306 6400 32312 6452
rect 32364 6440 32370 6452
rect 33134 6440 33140 6452
rect 32364 6412 33140 6440
rect 32364 6400 32370 6412
rect 33134 6400 33140 6412
rect 33192 6400 33198 6452
rect 35253 6443 35311 6449
rect 35253 6409 35265 6443
rect 35299 6440 35311 6443
rect 35986 6440 35992 6452
rect 35299 6412 35992 6440
rect 35299 6409 35311 6412
rect 35253 6403 35311 6409
rect 35986 6400 35992 6412
rect 36044 6440 36050 6452
rect 38838 6440 38844 6452
rect 36044 6412 37504 6440
rect 38799 6412 38844 6440
rect 36044 6400 36050 6412
rect 31352 6344 31616 6372
rect 31352 6332 31358 6344
rect 27709 6307 27767 6313
rect 27709 6273 27721 6307
rect 27755 6304 27767 6307
rect 29914 6304 29920 6316
rect 27755 6276 29920 6304
rect 27755 6273 27767 6276
rect 27709 6267 27767 6273
rect 29914 6264 29920 6276
rect 29972 6264 29978 6316
rect 31386 6304 31392 6316
rect 30484 6276 31392 6304
rect 27617 6239 27675 6245
rect 27617 6205 27629 6239
rect 27663 6205 27675 6239
rect 27617 6199 27675 6205
rect 28261 6239 28319 6245
rect 28261 6205 28273 6239
rect 28307 6205 28319 6239
rect 28534 6236 28540 6248
rect 28495 6208 28540 6236
rect 28261 6199 28319 6205
rect 15488 6140 16620 6168
rect 16758 6128 16764 6180
rect 16816 6168 16822 6180
rect 23845 6171 23903 6177
rect 16816 6140 17448 6168
rect 16816 6128 16822 6140
rect 5258 6100 5264 6112
rect 3844 6072 5264 6100
rect 3844 6060 3850 6072
rect 5258 6060 5264 6072
rect 5316 6060 5322 6112
rect 12526 6100 12532 6112
rect 12487 6072 12532 6100
rect 12526 6060 12532 6072
rect 12584 6060 12590 6112
rect 17420 6109 17448 6140
rect 23845 6137 23857 6171
rect 23891 6168 23903 6171
rect 25406 6168 25412 6180
rect 23891 6140 25412 6168
rect 23891 6137 23903 6140
rect 23845 6131 23903 6137
rect 25406 6128 25412 6140
rect 25464 6128 25470 6180
rect 26252 6168 26280 6196
rect 28276 6168 28304 6199
rect 28534 6196 28540 6208
rect 28592 6196 28598 6248
rect 28721 6239 28779 6245
rect 28721 6205 28733 6239
rect 28767 6236 28779 6239
rect 29086 6236 29092 6248
rect 28767 6208 29092 6236
rect 28767 6205 28779 6208
rect 28721 6199 28779 6205
rect 29086 6196 29092 6208
rect 29144 6196 29150 6248
rect 29178 6196 29184 6248
rect 29236 6236 29242 6248
rect 29273 6239 29331 6245
rect 29273 6236 29285 6239
rect 29236 6208 29285 6236
rect 29236 6196 29242 6208
rect 29273 6205 29285 6208
rect 29319 6205 29331 6239
rect 30190 6236 30196 6248
rect 30151 6208 30196 6236
rect 29273 6199 29331 6205
rect 30190 6196 30196 6208
rect 30248 6196 30254 6248
rect 30282 6196 30288 6248
rect 30340 6236 30346 6248
rect 30484 6236 30512 6276
rect 31386 6264 31392 6276
rect 31444 6264 31450 6316
rect 32677 6307 32735 6313
rect 32677 6273 32689 6307
rect 32723 6304 32735 6307
rect 34422 6304 34428 6316
rect 32723 6276 34428 6304
rect 32723 6273 32735 6276
rect 32677 6267 32735 6273
rect 34422 6264 34428 6276
rect 34480 6264 34486 6316
rect 36078 6304 36084 6316
rect 34532 6276 36084 6304
rect 30340 6208 30512 6236
rect 30561 6239 30619 6245
rect 30340 6196 30346 6208
rect 30561 6205 30573 6239
rect 30607 6236 30619 6239
rect 32122 6236 32128 6248
rect 30607 6208 32128 6236
rect 30607 6205 30619 6208
rect 30561 6199 30619 6205
rect 32122 6196 32128 6208
rect 32180 6196 32186 6248
rect 32398 6236 32404 6248
rect 32359 6208 32404 6236
rect 32398 6196 32404 6208
rect 32456 6196 32462 6248
rect 32950 6196 32956 6248
rect 33008 6236 33014 6248
rect 33962 6236 33968 6248
rect 33008 6208 33968 6236
rect 33008 6196 33014 6208
rect 33962 6196 33968 6208
rect 34020 6236 34026 6248
rect 34057 6239 34115 6245
rect 34057 6236 34069 6239
rect 34020 6208 34069 6236
rect 34020 6196 34026 6208
rect 34057 6205 34069 6208
rect 34103 6236 34115 6239
rect 34532 6236 34560 6276
rect 36078 6264 36084 6276
rect 36136 6264 36142 6316
rect 37476 6313 37504 6412
rect 38838 6400 38844 6412
rect 38896 6400 38902 6452
rect 37461 6307 37519 6313
rect 37461 6273 37473 6307
rect 37507 6273 37519 6307
rect 37734 6304 37740 6316
rect 37695 6276 37740 6304
rect 37461 6267 37519 6273
rect 37734 6264 37740 6276
rect 37792 6264 37798 6316
rect 34103 6208 34560 6236
rect 35253 6239 35311 6245
rect 34103 6205 34115 6208
rect 34057 6199 34115 6205
rect 35253 6205 35265 6239
rect 35299 6236 35311 6239
rect 35345 6239 35403 6245
rect 35345 6236 35357 6239
rect 35299 6208 35357 6236
rect 35299 6205 35311 6208
rect 35253 6199 35311 6205
rect 35345 6205 35357 6208
rect 35391 6205 35403 6239
rect 35345 6199 35403 6205
rect 35621 6239 35679 6245
rect 35621 6205 35633 6239
rect 35667 6236 35679 6239
rect 37366 6236 37372 6248
rect 35667 6208 37372 6236
rect 35667 6205 35679 6208
rect 35621 6199 35679 6205
rect 37366 6196 37372 6208
rect 37424 6196 37430 6248
rect 30374 6168 30380 6180
rect 26252 6140 30380 6168
rect 30374 6128 30380 6140
rect 30432 6128 30438 6180
rect 32306 6168 32312 6180
rect 31220 6140 32312 6168
rect 17405 6103 17463 6109
rect 17405 6069 17417 6103
rect 17451 6069 17463 6103
rect 17405 6063 17463 6069
rect 17770 6060 17776 6112
rect 17828 6100 17834 6112
rect 18141 6103 18199 6109
rect 18141 6100 18153 6103
rect 17828 6072 18153 6100
rect 17828 6060 17834 6072
rect 18141 6069 18153 6072
rect 18187 6069 18199 6103
rect 18141 6063 18199 6069
rect 20898 6060 20904 6112
rect 20956 6100 20962 6112
rect 25038 6100 25044 6112
rect 20956 6072 25044 6100
rect 20956 6060 20962 6072
rect 25038 6060 25044 6072
rect 25096 6060 25102 6112
rect 29457 6103 29515 6109
rect 29457 6069 29469 6103
rect 29503 6100 29515 6103
rect 29822 6100 29828 6112
rect 29503 6072 29828 6100
rect 29503 6069 29515 6072
rect 29457 6063 29515 6069
rect 29822 6060 29828 6072
rect 29880 6100 29886 6112
rect 31220 6100 31248 6140
rect 32306 6128 32312 6140
rect 32364 6128 32370 6180
rect 29880 6072 31248 6100
rect 29880 6060 29886 6072
rect 33962 6060 33968 6112
rect 34020 6100 34026 6112
rect 36725 6103 36783 6109
rect 36725 6100 36737 6103
rect 34020 6072 36737 6100
rect 34020 6060 34026 6072
rect 36725 6069 36737 6072
rect 36771 6069 36783 6103
rect 36725 6063 36783 6069
rect 1104 6010 39836 6032
rect 1104 5958 19606 6010
rect 19658 5958 19670 6010
rect 19722 5958 19734 6010
rect 19786 5958 19798 6010
rect 19850 5958 39836 6010
rect 1104 5936 39836 5958
rect 2498 5896 2504 5908
rect 2459 5868 2504 5896
rect 2498 5856 2504 5868
rect 2556 5856 2562 5908
rect 4157 5899 4215 5905
rect 4157 5896 4169 5899
rect 2608 5868 4169 5896
rect 2608 5769 2636 5868
rect 4157 5865 4169 5868
rect 4203 5865 4215 5899
rect 4157 5859 4215 5865
rect 4264 5868 6316 5896
rect 3970 5788 3976 5840
rect 4028 5828 4034 5840
rect 4264 5828 4292 5868
rect 4028 5800 4292 5828
rect 6288 5828 6316 5868
rect 8202 5856 8208 5908
rect 8260 5896 8266 5908
rect 10873 5899 10931 5905
rect 10873 5896 10885 5899
rect 8260 5868 10885 5896
rect 8260 5856 8266 5868
rect 10873 5865 10885 5868
rect 10919 5865 10931 5899
rect 10873 5859 10931 5865
rect 10980 5868 12848 5896
rect 10980 5828 11008 5868
rect 6288 5800 11008 5828
rect 12820 5828 12848 5868
rect 12894 5856 12900 5908
rect 12952 5896 12958 5908
rect 13909 5899 13967 5905
rect 13909 5896 13921 5899
rect 12952 5868 13921 5896
rect 12952 5856 12958 5868
rect 13909 5865 13921 5868
rect 13955 5865 13967 5899
rect 13909 5859 13967 5865
rect 14550 5856 14556 5908
rect 14608 5896 14614 5908
rect 15381 5899 15439 5905
rect 15381 5896 15393 5899
rect 14608 5868 15393 5896
rect 14608 5856 14614 5868
rect 15381 5865 15393 5868
rect 15427 5865 15439 5899
rect 15381 5859 15439 5865
rect 16850 5856 16856 5908
rect 16908 5856 16914 5908
rect 17954 5856 17960 5908
rect 18012 5896 18018 5908
rect 19705 5899 19763 5905
rect 19705 5896 19717 5899
rect 18012 5868 19717 5896
rect 18012 5856 18018 5868
rect 19705 5865 19717 5868
rect 19751 5865 19763 5899
rect 24578 5896 24584 5908
rect 24539 5868 24584 5896
rect 19705 5859 19763 5865
rect 24578 5856 24584 5868
rect 24636 5856 24642 5908
rect 28626 5896 28632 5908
rect 24688 5868 28632 5896
rect 16868 5828 16896 5856
rect 12820 5800 13952 5828
rect 4028 5788 4034 5800
rect 2593 5763 2651 5769
rect 2593 5729 2605 5763
rect 2639 5729 2651 5763
rect 2593 5723 2651 5729
rect 3145 5763 3203 5769
rect 3145 5729 3157 5763
rect 3191 5729 3203 5763
rect 3145 5723 3203 5729
rect 3160 5692 3188 5723
rect 3326 5720 3332 5772
rect 3384 5760 3390 5772
rect 3421 5763 3479 5769
rect 3421 5760 3433 5763
rect 3384 5732 3433 5760
rect 3384 5720 3390 5732
rect 3421 5729 3433 5732
rect 3467 5760 3479 5763
rect 4065 5763 4123 5769
rect 4065 5760 4077 5763
rect 3467 5732 4077 5760
rect 3467 5729 3479 5732
rect 3421 5723 3479 5729
rect 4065 5729 4077 5732
rect 4111 5729 4123 5763
rect 4065 5723 4123 5729
rect 4154 5720 4160 5772
rect 4212 5760 4218 5772
rect 4617 5763 4675 5769
rect 4617 5760 4629 5763
rect 4212 5732 4629 5760
rect 4212 5720 4218 5732
rect 4617 5729 4629 5732
rect 4663 5760 4675 5763
rect 4982 5760 4988 5772
rect 4663 5732 4988 5760
rect 4663 5729 4675 5732
rect 4617 5723 4675 5729
rect 4982 5720 4988 5732
rect 5040 5720 5046 5772
rect 5258 5720 5264 5772
rect 5316 5760 5322 5772
rect 5353 5763 5411 5769
rect 5353 5760 5365 5763
rect 5316 5732 5365 5760
rect 5316 5720 5322 5732
rect 5353 5729 5365 5732
rect 5399 5729 5411 5763
rect 5353 5723 5411 5729
rect 8941 5763 8999 5769
rect 8941 5729 8953 5763
rect 8987 5760 8999 5763
rect 9674 5760 9680 5772
rect 8987 5732 9680 5760
rect 8987 5729 8999 5732
rect 8941 5723 8999 5729
rect 9674 5720 9680 5732
rect 9732 5720 9738 5772
rect 9861 5763 9919 5769
rect 9861 5729 9873 5763
rect 9907 5729 9919 5763
rect 9861 5723 9919 5729
rect 4706 5692 4712 5704
rect 3160 5664 4712 5692
rect 4706 5652 4712 5664
rect 4764 5652 4770 5704
rect 5629 5695 5687 5701
rect 5629 5661 5641 5695
rect 5675 5692 5687 5695
rect 6270 5692 6276 5704
rect 5675 5664 6276 5692
rect 5675 5661 5687 5664
rect 5629 5655 5687 5661
rect 6270 5652 6276 5664
rect 6328 5652 6334 5704
rect 4522 5584 4528 5636
rect 4580 5624 4586 5636
rect 4798 5624 4804 5636
rect 4580 5596 4804 5624
rect 4580 5584 4586 5596
rect 4798 5584 4804 5596
rect 4856 5584 4862 5636
rect 9876 5624 9904 5723
rect 9950 5720 9956 5772
rect 10008 5760 10014 5772
rect 10318 5760 10324 5772
rect 10008 5732 10053 5760
rect 10279 5732 10324 5760
rect 10008 5720 10014 5732
rect 10318 5720 10324 5732
rect 10376 5720 10382 5772
rect 10413 5763 10471 5769
rect 10413 5729 10425 5763
rect 10459 5760 10471 5763
rect 10962 5760 10968 5772
rect 10459 5732 10968 5760
rect 10459 5729 10471 5732
rect 10413 5723 10471 5729
rect 10962 5720 10968 5732
rect 11020 5720 11026 5772
rect 11974 5760 11980 5772
rect 11935 5732 11980 5760
rect 11974 5720 11980 5732
rect 12032 5720 12038 5772
rect 13817 5763 13875 5769
rect 13817 5760 13829 5763
rect 13096 5732 13829 5760
rect 11701 5695 11759 5701
rect 11701 5661 11713 5695
rect 11747 5692 11759 5695
rect 11882 5692 11888 5704
rect 11747 5664 11888 5692
rect 11747 5661 11759 5664
rect 11701 5655 11759 5661
rect 11882 5652 11888 5664
rect 11940 5692 11946 5704
rect 12618 5692 12624 5704
rect 11940 5664 12624 5692
rect 11940 5652 11946 5664
rect 12618 5652 12624 5664
rect 12676 5652 12682 5704
rect 12802 5652 12808 5704
rect 12860 5692 12866 5704
rect 13096 5701 13124 5732
rect 13817 5729 13829 5732
rect 13863 5729 13875 5763
rect 13817 5723 13875 5729
rect 13081 5695 13139 5701
rect 13081 5692 13093 5695
rect 12860 5664 13093 5692
rect 12860 5652 12866 5664
rect 13081 5661 13093 5664
rect 13127 5661 13139 5695
rect 13081 5655 13139 5661
rect 10410 5624 10416 5636
rect 9876 5596 10416 5624
rect 10410 5584 10416 5596
rect 10468 5584 10474 5636
rect 12636 5624 12664 5652
rect 13722 5624 13728 5636
rect 12636 5596 13728 5624
rect 13722 5584 13728 5596
rect 13780 5584 13786 5636
rect 5350 5516 5356 5568
rect 5408 5556 5414 5568
rect 6733 5559 6791 5565
rect 6733 5556 6745 5559
rect 5408 5528 6745 5556
rect 5408 5516 5414 5528
rect 6733 5525 6745 5528
rect 6779 5525 6791 5559
rect 6733 5519 6791 5525
rect 9033 5559 9091 5565
rect 9033 5525 9045 5559
rect 9079 5556 9091 5559
rect 10778 5556 10784 5568
rect 9079 5528 10784 5556
rect 9079 5525 9091 5528
rect 9033 5519 9091 5525
rect 10778 5516 10784 5528
rect 10836 5516 10842 5568
rect 13924 5556 13952 5800
rect 16684 5800 18092 5828
rect 15286 5760 15292 5772
rect 15247 5732 15292 5760
rect 15286 5720 15292 5732
rect 15344 5720 15350 5772
rect 16117 5763 16175 5769
rect 16117 5729 16129 5763
rect 16163 5729 16175 5763
rect 16117 5723 16175 5729
rect 16209 5763 16267 5769
rect 16209 5729 16221 5763
rect 16255 5760 16267 5763
rect 16298 5760 16304 5772
rect 16255 5732 16304 5760
rect 16255 5729 16267 5732
rect 16209 5723 16267 5729
rect 15654 5584 15660 5636
rect 15712 5624 15718 5636
rect 16132 5624 16160 5723
rect 16298 5720 16304 5732
rect 16356 5720 16362 5772
rect 16684 5769 16712 5800
rect 16669 5763 16727 5769
rect 16669 5729 16681 5763
rect 16715 5729 16727 5763
rect 16669 5723 16727 5729
rect 16853 5763 16911 5769
rect 16853 5729 16865 5763
rect 16899 5760 16911 5763
rect 17034 5760 17040 5772
rect 16899 5732 17040 5760
rect 16899 5729 16911 5732
rect 16853 5723 16911 5729
rect 17034 5720 17040 5732
rect 17092 5720 17098 5772
rect 17678 5720 17684 5772
rect 17736 5760 17742 5772
rect 17957 5763 18015 5769
rect 17957 5760 17969 5763
rect 17736 5732 17969 5760
rect 17736 5720 17742 5732
rect 17957 5729 17969 5732
rect 18003 5729 18015 5763
rect 18064 5760 18092 5800
rect 18322 5788 18328 5840
rect 18380 5828 18386 5840
rect 18380 5800 19656 5828
rect 18380 5788 18386 5800
rect 18509 5763 18567 5769
rect 18509 5760 18521 5763
rect 18064 5732 18521 5760
rect 17957 5723 18015 5729
rect 18509 5729 18521 5732
rect 18555 5729 18567 5763
rect 18509 5723 18567 5729
rect 18693 5763 18751 5769
rect 18693 5729 18705 5763
rect 18739 5760 18751 5763
rect 19334 5760 19340 5772
rect 18739 5732 19340 5760
rect 18739 5729 18751 5732
rect 18693 5723 18751 5729
rect 19334 5720 19340 5732
rect 19392 5720 19398 5772
rect 19628 5769 19656 5800
rect 19613 5763 19671 5769
rect 19613 5729 19625 5763
rect 19659 5729 19671 5763
rect 20898 5760 20904 5772
rect 20859 5732 20904 5760
rect 19613 5723 19671 5729
rect 20898 5720 20904 5732
rect 20956 5720 20962 5772
rect 21266 5760 21272 5772
rect 21227 5732 21272 5760
rect 21266 5720 21272 5732
rect 21324 5720 21330 5772
rect 21913 5763 21971 5769
rect 21913 5729 21925 5763
rect 21959 5760 21971 5763
rect 22186 5760 22192 5772
rect 21959 5732 22192 5760
rect 21959 5729 21971 5732
rect 21913 5723 21971 5729
rect 22186 5720 22192 5732
rect 22244 5760 22250 5772
rect 22738 5760 22744 5772
rect 22244 5732 22744 5760
rect 22244 5720 22250 5732
rect 22738 5720 22744 5732
rect 22796 5760 22802 5772
rect 24688 5760 24716 5868
rect 28626 5856 28632 5868
rect 28684 5896 28690 5908
rect 28684 5868 30328 5896
rect 28684 5856 28690 5868
rect 28077 5831 28135 5837
rect 28077 5797 28089 5831
rect 28123 5828 28135 5831
rect 29730 5828 29736 5840
rect 28123 5800 29736 5828
rect 28123 5797 28135 5800
rect 28077 5791 28135 5797
rect 29730 5788 29736 5800
rect 29788 5788 29794 5840
rect 30300 5828 30328 5868
rect 30484 5868 36768 5896
rect 30484 5828 30512 5868
rect 30300 5800 30512 5828
rect 30561 5831 30619 5837
rect 30561 5797 30573 5831
rect 30607 5828 30619 5831
rect 36170 5828 36176 5840
rect 30607 5800 33088 5828
rect 36131 5800 36176 5828
rect 30607 5797 30619 5800
rect 30561 5791 30619 5797
rect 22796 5732 24716 5760
rect 22796 5720 22802 5732
rect 24854 5720 24860 5772
rect 24912 5760 24918 5772
rect 25133 5763 25191 5769
rect 25133 5760 25145 5763
rect 24912 5732 25145 5760
rect 24912 5720 24918 5732
rect 25133 5729 25145 5732
rect 25179 5729 25191 5763
rect 27062 5760 27068 5772
rect 25133 5723 25191 5729
rect 25332 5732 27068 5760
rect 17218 5692 17224 5704
rect 17179 5664 17224 5692
rect 17218 5652 17224 5664
rect 17276 5652 17282 5704
rect 17696 5624 17724 5720
rect 17862 5692 17868 5704
rect 17823 5664 17868 5692
rect 17862 5652 17868 5664
rect 17920 5652 17926 5704
rect 20346 5652 20352 5704
rect 20404 5692 20410 5704
rect 20993 5695 21051 5701
rect 20993 5692 21005 5695
rect 20404 5664 21005 5692
rect 20404 5652 20410 5664
rect 20993 5661 21005 5664
rect 21039 5661 21051 5695
rect 21284 5692 21312 5720
rect 22094 5692 22100 5704
rect 21284 5664 22100 5692
rect 20993 5655 21051 5661
rect 22094 5652 22100 5664
rect 22152 5652 22158 5704
rect 23014 5692 23020 5704
rect 22975 5664 23020 5692
rect 23014 5652 23020 5664
rect 23072 5652 23078 5704
rect 23293 5695 23351 5701
rect 23293 5661 23305 5695
rect 23339 5692 23351 5695
rect 25038 5692 25044 5704
rect 23339 5664 25044 5692
rect 23339 5661 23351 5664
rect 23293 5655 23351 5661
rect 25038 5652 25044 5664
rect 25096 5652 25102 5704
rect 18874 5624 18880 5636
rect 15712 5596 17724 5624
rect 18835 5596 18880 5624
rect 15712 5584 15718 5596
rect 18874 5584 18880 5596
rect 18932 5584 18938 5636
rect 21266 5584 21272 5636
rect 21324 5624 21330 5636
rect 23032 5624 23060 5652
rect 21324 5596 23060 5624
rect 21324 5584 21330 5596
rect 24394 5584 24400 5636
rect 24452 5624 24458 5636
rect 25332 5633 25360 5732
rect 27062 5720 27068 5732
rect 27120 5720 27126 5772
rect 27154 5720 27160 5772
rect 27212 5760 27218 5772
rect 27341 5763 27399 5769
rect 27341 5760 27353 5763
rect 27212 5732 27353 5760
rect 27212 5720 27218 5732
rect 27341 5729 27353 5732
rect 27387 5729 27399 5763
rect 27341 5723 27399 5729
rect 28905 5763 28963 5769
rect 28905 5729 28917 5763
rect 28951 5760 28963 5763
rect 29270 5760 29276 5772
rect 28951 5732 29276 5760
rect 28951 5729 28963 5732
rect 28905 5723 28963 5729
rect 29270 5720 29276 5732
rect 29328 5720 29334 5772
rect 29549 5763 29607 5769
rect 29549 5729 29561 5763
rect 29595 5760 29607 5763
rect 30374 5760 30380 5772
rect 29595 5732 30380 5760
rect 29595 5729 29607 5732
rect 29549 5723 29607 5729
rect 30374 5720 30380 5732
rect 30432 5760 30438 5772
rect 30834 5760 30840 5772
rect 30432 5732 30840 5760
rect 30432 5720 30438 5732
rect 30834 5720 30840 5732
rect 30892 5720 30898 5772
rect 31294 5720 31300 5772
rect 31352 5760 31358 5772
rect 31389 5763 31447 5769
rect 31389 5760 31401 5763
rect 31352 5732 31401 5760
rect 31352 5720 31358 5732
rect 31389 5729 31401 5732
rect 31435 5729 31447 5763
rect 31389 5723 31447 5729
rect 31573 5763 31631 5769
rect 31573 5729 31585 5763
rect 31619 5760 31631 5763
rect 31846 5760 31852 5772
rect 31619 5732 31852 5760
rect 31619 5729 31631 5732
rect 31573 5723 31631 5729
rect 31846 5720 31852 5732
rect 31904 5720 31910 5772
rect 32815 5763 32873 5769
rect 32815 5760 32827 5763
rect 32048 5732 32827 5760
rect 26510 5692 26516 5704
rect 26471 5664 26516 5692
rect 26510 5652 26516 5664
rect 26568 5652 26574 5704
rect 27525 5695 27583 5701
rect 27525 5661 27537 5695
rect 27571 5692 27583 5695
rect 28258 5692 28264 5704
rect 27571 5664 28264 5692
rect 27571 5661 27583 5664
rect 27525 5655 27583 5661
rect 28258 5652 28264 5664
rect 28316 5652 28322 5704
rect 28629 5695 28687 5701
rect 28629 5661 28641 5695
rect 28675 5661 28687 5695
rect 28629 5655 28687 5661
rect 25317 5627 25375 5633
rect 25317 5624 25329 5627
rect 24452 5596 25329 5624
rect 24452 5584 24458 5596
rect 25317 5593 25329 5596
rect 25363 5593 25375 5627
rect 25317 5587 25375 5593
rect 27062 5584 27068 5636
rect 27120 5624 27126 5636
rect 28644 5624 28672 5655
rect 28810 5652 28816 5704
rect 28868 5692 28874 5704
rect 29089 5695 29147 5701
rect 29089 5692 29101 5695
rect 28868 5664 29101 5692
rect 28868 5652 28874 5664
rect 29089 5661 29101 5664
rect 29135 5661 29147 5695
rect 29089 5655 29147 5661
rect 30558 5652 30564 5704
rect 30616 5692 30622 5704
rect 31113 5695 31171 5701
rect 31113 5692 31125 5695
rect 30616 5664 31125 5692
rect 30616 5652 30622 5664
rect 31113 5661 31125 5664
rect 31159 5692 31171 5695
rect 31478 5692 31484 5704
rect 31159 5664 31484 5692
rect 31159 5661 31171 5664
rect 31113 5655 31171 5661
rect 31478 5652 31484 5664
rect 31536 5652 31542 5704
rect 31662 5652 31668 5704
rect 31720 5692 31726 5704
rect 32048 5692 32076 5732
rect 32815 5729 32827 5732
rect 32861 5729 32873 5763
rect 32950 5760 32956 5772
rect 32911 5732 32956 5760
rect 32815 5723 32873 5729
rect 32950 5720 32956 5732
rect 33008 5720 33014 5772
rect 31720 5664 32076 5692
rect 31720 5652 31726 5664
rect 32122 5652 32128 5704
rect 32180 5692 32186 5704
rect 32677 5695 32735 5701
rect 32180 5664 32225 5692
rect 32180 5652 32186 5664
rect 32677 5661 32689 5695
rect 32723 5692 32735 5695
rect 33060 5692 33088 5800
rect 36170 5788 36176 5800
rect 36228 5788 36234 5840
rect 34333 5763 34391 5769
rect 34333 5729 34345 5763
rect 34379 5760 34391 5763
rect 35894 5760 35900 5772
rect 34379 5732 35900 5760
rect 34379 5729 34391 5732
rect 34333 5723 34391 5729
rect 35894 5720 35900 5732
rect 35952 5720 35958 5772
rect 36740 5769 36768 5868
rect 37366 5856 37372 5908
rect 37424 5896 37430 5908
rect 37829 5899 37887 5905
rect 37829 5896 37841 5899
rect 37424 5868 37841 5896
rect 37424 5856 37430 5868
rect 37829 5865 37841 5868
rect 37875 5865 37887 5899
rect 37829 5859 37887 5865
rect 38378 5856 38384 5908
rect 38436 5896 38442 5908
rect 39025 5899 39083 5905
rect 39025 5896 39037 5899
rect 38436 5868 39037 5896
rect 38436 5856 38442 5868
rect 39025 5865 39037 5868
rect 39071 5865 39083 5899
rect 39025 5859 39083 5865
rect 36725 5763 36783 5769
rect 36725 5729 36737 5763
rect 36771 5729 36783 5763
rect 36998 5760 37004 5772
rect 36959 5732 37004 5760
rect 36725 5723 36783 5729
rect 36998 5720 37004 5732
rect 37056 5720 37062 5772
rect 37826 5760 37832 5772
rect 37787 5732 37832 5760
rect 37826 5720 37832 5732
rect 37884 5720 37890 5772
rect 38194 5760 38200 5772
rect 38155 5732 38200 5760
rect 38194 5720 38200 5732
rect 38252 5720 38258 5772
rect 38838 5720 38844 5772
rect 38896 5760 38902 5772
rect 38933 5763 38991 5769
rect 38933 5760 38945 5763
rect 38896 5732 38945 5760
rect 38896 5720 38902 5732
rect 38933 5729 38945 5732
rect 38979 5729 38991 5763
rect 38933 5723 38991 5729
rect 32723 5664 33088 5692
rect 34057 5695 34115 5701
rect 32723 5661 32735 5664
rect 32677 5655 32735 5661
rect 34057 5661 34069 5695
rect 34103 5692 34115 5695
rect 35986 5692 35992 5704
rect 34103 5664 35992 5692
rect 34103 5661 34115 5664
rect 34057 5655 34115 5661
rect 27120 5596 28672 5624
rect 27120 5584 27126 5596
rect 32398 5584 32404 5636
rect 32456 5624 32462 5636
rect 32950 5624 32956 5636
rect 32456 5596 32956 5624
rect 32456 5584 32462 5596
rect 32950 5584 32956 5596
rect 33008 5624 33014 5636
rect 34072 5624 34100 5655
rect 35986 5652 35992 5664
rect 36044 5652 36050 5704
rect 37185 5695 37243 5701
rect 37185 5661 37197 5695
rect 37231 5661 37243 5695
rect 37185 5655 37243 5661
rect 35434 5624 35440 5636
rect 33008 5596 34100 5624
rect 35395 5596 35440 5624
rect 33008 5584 33014 5596
rect 35434 5584 35440 5596
rect 35492 5624 35498 5636
rect 37200 5624 37228 5655
rect 35492 5596 37228 5624
rect 35492 5584 35498 5596
rect 19242 5556 19248 5568
rect 13924 5528 19248 5556
rect 19242 5516 19248 5528
rect 19300 5516 19306 5568
rect 23290 5516 23296 5568
rect 23348 5556 23354 5568
rect 28166 5556 28172 5568
rect 23348 5528 28172 5556
rect 23348 5516 23354 5528
rect 28166 5516 28172 5528
rect 28224 5516 28230 5568
rect 28350 5516 28356 5568
rect 28408 5556 28414 5568
rect 29733 5559 29791 5565
rect 29733 5556 29745 5559
rect 28408 5528 29745 5556
rect 28408 5516 28414 5528
rect 29733 5525 29745 5528
rect 29779 5525 29791 5559
rect 29733 5519 29791 5525
rect 1104 5466 39836 5488
rect 1104 5414 4246 5466
rect 4298 5414 4310 5466
rect 4362 5414 4374 5466
rect 4426 5414 4438 5466
rect 4490 5414 34966 5466
rect 35018 5414 35030 5466
rect 35082 5414 35094 5466
rect 35146 5414 35158 5466
rect 35210 5414 39836 5466
rect 1104 5392 39836 5414
rect 3053 5355 3111 5361
rect 3053 5321 3065 5355
rect 3099 5352 3111 5355
rect 3326 5352 3332 5364
rect 3099 5324 3332 5352
rect 3099 5321 3111 5324
rect 3053 5315 3111 5321
rect 3326 5312 3332 5324
rect 3384 5312 3390 5364
rect 9674 5352 9680 5364
rect 9587 5324 9680 5352
rect 9674 5312 9680 5324
rect 9732 5352 9738 5364
rect 10594 5352 10600 5364
rect 9732 5324 10600 5352
rect 9732 5312 9738 5324
rect 10594 5312 10600 5324
rect 10652 5312 10658 5364
rect 10778 5312 10784 5364
rect 10836 5352 10842 5364
rect 10836 5324 17356 5352
rect 10836 5312 10842 5324
rect 5074 5284 5080 5296
rect 4448 5256 5080 5284
rect 1765 5219 1823 5225
rect 1765 5185 1777 5219
rect 1811 5216 1823 5219
rect 2958 5216 2964 5228
rect 1811 5188 2964 5216
rect 1811 5185 1823 5188
rect 1765 5179 1823 5185
rect 2958 5176 2964 5188
rect 3016 5176 3022 5228
rect 1489 5151 1547 5157
rect 1489 5117 1501 5151
rect 1535 5148 1547 5151
rect 3142 5148 3148 5160
rect 1535 5120 3148 5148
rect 1535 5117 1547 5120
rect 1489 5111 1547 5117
rect 3142 5108 3148 5120
rect 3200 5108 3206 5160
rect 4341 5151 4399 5157
rect 4341 5117 4353 5151
rect 4387 5148 4399 5151
rect 4448 5148 4476 5256
rect 5074 5244 5080 5256
rect 5132 5244 5138 5296
rect 11333 5287 11391 5293
rect 11333 5284 11345 5287
rect 9876 5256 11345 5284
rect 4706 5216 4712 5228
rect 4667 5188 4712 5216
rect 4706 5176 4712 5188
rect 4764 5176 4770 5228
rect 5166 5216 5172 5228
rect 5092 5188 5172 5216
rect 5092 5157 5120 5188
rect 5166 5176 5172 5188
rect 5224 5176 5230 5228
rect 8113 5219 8171 5225
rect 8113 5185 8125 5219
rect 8159 5216 8171 5219
rect 8294 5216 8300 5228
rect 8159 5188 8300 5216
rect 8159 5185 8171 5188
rect 8113 5179 8171 5185
rect 8294 5176 8300 5188
rect 8352 5176 8358 5228
rect 8389 5219 8447 5225
rect 8389 5185 8401 5219
rect 8435 5216 8447 5219
rect 9876 5216 9904 5256
rect 11333 5253 11345 5256
rect 11379 5253 11391 5287
rect 11333 5247 11391 5253
rect 11422 5244 11428 5296
rect 11480 5284 11486 5296
rect 13725 5287 13783 5293
rect 13725 5284 13737 5287
rect 11480 5256 13737 5284
rect 11480 5244 11486 5256
rect 13725 5253 13737 5256
rect 13771 5253 13783 5287
rect 13725 5247 13783 5253
rect 8435 5188 9904 5216
rect 8435 5185 8447 5188
rect 8389 5179 8447 5185
rect 12526 5176 12532 5228
rect 12584 5216 12590 5228
rect 12584 5188 14136 5216
rect 12584 5176 12590 5188
rect 4387 5120 4476 5148
rect 4617 5151 4675 5157
rect 4387 5117 4399 5120
rect 4341 5111 4399 5117
rect 4617 5117 4629 5151
rect 4663 5117 4675 5151
rect 4617 5111 4675 5117
rect 5077 5151 5135 5157
rect 5077 5117 5089 5151
rect 5123 5117 5135 5151
rect 5077 5111 5135 5117
rect 4522 4972 4528 5024
rect 4580 5012 4586 5024
rect 4632 5012 4660 5111
rect 5350 5108 5356 5160
rect 5408 5148 5414 5160
rect 5721 5151 5779 5157
rect 5721 5148 5733 5151
rect 5408 5120 5733 5148
rect 5408 5108 5414 5120
rect 5721 5117 5733 5120
rect 5767 5117 5779 5151
rect 5721 5111 5779 5117
rect 5905 5151 5963 5157
rect 5905 5117 5917 5151
rect 5951 5117 5963 5151
rect 10410 5148 10416 5160
rect 10371 5120 10416 5148
rect 5905 5111 5963 5117
rect 5166 5040 5172 5092
rect 5224 5080 5230 5092
rect 5920 5080 5948 5111
rect 10410 5108 10416 5120
rect 10468 5108 10474 5160
rect 10505 5151 10563 5157
rect 10505 5117 10517 5151
rect 10551 5148 10563 5151
rect 10594 5148 10600 5160
rect 10551 5120 10600 5148
rect 10551 5117 10563 5120
rect 10505 5111 10563 5117
rect 10594 5108 10600 5120
rect 10652 5108 10658 5160
rect 10778 5108 10784 5160
rect 10836 5148 10842 5160
rect 10873 5151 10931 5157
rect 10873 5148 10885 5151
rect 10836 5120 10885 5148
rect 10836 5108 10842 5120
rect 10873 5117 10885 5120
rect 10919 5117 10931 5151
rect 10873 5111 10931 5117
rect 10962 5108 10968 5160
rect 11020 5148 11026 5160
rect 12066 5148 12072 5160
rect 11020 5120 12072 5148
rect 11020 5108 11026 5120
rect 12066 5108 12072 5120
rect 12124 5108 12130 5160
rect 12434 5108 12440 5160
rect 12492 5148 12498 5160
rect 12618 5148 12624 5160
rect 12492 5120 12624 5148
rect 12492 5108 12498 5120
rect 12618 5108 12624 5120
rect 12676 5108 12682 5160
rect 12897 5151 12955 5157
rect 12897 5117 12909 5151
rect 12943 5117 12955 5151
rect 12897 5111 12955 5117
rect 13725 5151 13783 5157
rect 13725 5117 13737 5151
rect 13771 5148 13783 5151
rect 13906 5148 13912 5160
rect 13771 5120 13912 5148
rect 13771 5117 13783 5120
rect 13725 5111 13783 5117
rect 5224 5052 5948 5080
rect 5224 5040 5230 5052
rect 11054 5040 11060 5092
rect 11112 5080 11118 5092
rect 12912 5080 12940 5111
rect 13906 5108 13912 5120
rect 13964 5108 13970 5160
rect 14108 5157 14136 5188
rect 15194 5176 15200 5228
rect 15252 5216 15258 5228
rect 15252 5188 16436 5216
rect 15252 5176 15258 5188
rect 16408 5160 16436 5188
rect 14093 5151 14151 5157
rect 14093 5117 14105 5151
rect 14139 5117 14151 5151
rect 14642 5148 14648 5160
rect 14603 5120 14648 5148
rect 14093 5111 14151 5117
rect 14642 5108 14648 5120
rect 14700 5108 14706 5160
rect 15010 5148 15016 5160
rect 14971 5120 15016 5148
rect 15010 5108 15016 5120
rect 15068 5108 15074 5160
rect 15562 5148 15568 5160
rect 15523 5120 15568 5148
rect 15562 5108 15568 5120
rect 15620 5108 15626 5160
rect 15838 5108 15844 5160
rect 15896 5148 15902 5160
rect 16025 5151 16083 5157
rect 16025 5148 16037 5151
rect 15896 5120 16037 5148
rect 15896 5108 15902 5120
rect 16025 5117 16037 5120
rect 16071 5117 16083 5151
rect 16206 5148 16212 5160
rect 16167 5120 16212 5148
rect 16025 5111 16083 5117
rect 16206 5108 16212 5120
rect 16264 5108 16270 5160
rect 16390 5108 16396 5160
rect 16448 5148 16454 5160
rect 16669 5151 16727 5157
rect 16669 5148 16681 5151
rect 16448 5120 16681 5148
rect 16448 5108 16454 5120
rect 16669 5117 16681 5120
rect 16715 5117 16727 5151
rect 16669 5111 16727 5117
rect 16758 5108 16764 5160
rect 16816 5148 16822 5160
rect 16816 5120 16861 5148
rect 16816 5108 16822 5120
rect 11112 5052 12940 5080
rect 11112 5040 11118 5052
rect 5350 5012 5356 5024
rect 4580 4984 5356 5012
rect 4580 4972 4586 4984
rect 5350 4972 5356 4984
rect 5408 4972 5414 5024
rect 5810 4972 5816 5024
rect 5868 5012 5874 5024
rect 5997 5015 6055 5021
rect 5997 5012 6009 5015
rect 5868 4984 6009 5012
rect 5868 4972 5874 4984
rect 5997 4981 6009 4984
rect 6043 4981 6055 5015
rect 12710 5012 12716 5024
rect 12671 4984 12716 5012
rect 5997 4975 6055 4981
rect 12710 4972 12716 4984
rect 12768 4972 12774 5024
rect 16574 4972 16580 5024
rect 16632 5012 16638 5024
rect 17221 5015 17279 5021
rect 17221 5012 17233 5015
rect 16632 4984 17233 5012
rect 16632 4972 16638 4984
rect 17221 4981 17233 4984
rect 17267 4981 17279 5015
rect 17328 5012 17356 5324
rect 18782 5312 18788 5364
rect 18840 5352 18846 5364
rect 19889 5355 19947 5361
rect 19889 5352 19901 5355
rect 18840 5324 19901 5352
rect 18840 5312 18846 5324
rect 19889 5321 19901 5324
rect 19935 5321 19947 5355
rect 19889 5315 19947 5321
rect 23845 5355 23903 5361
rect 23845 5321 23857 5355
rect 23891 5352 23903 5355
rect 24486 5352 24492 5364
rect 23891 5324 24492 5352
rect 23891 5321 23903 5324
rect 23845 5315 23903 5321
rect 18785 5219 18843 5225
rect 18785 5185 18797 5219
rect 18831 5216 18843 5219
rect 18874 5216 18880 5228
rect 18831 5188 18880 5216
rect 18831 5185 18843 5188
rect 18785 5179 18843 5185
rect 18874 5176 18880 5188
rect 18932 5176 18938 5228
rect 17954 5108 17960 5160
rect 18012 5148 18018 5160
rect 18506 5148 18512 5160
rect 18012 5120 18512 5148
rect 18012 5108 18018 5120
rect 18506 5108 18512 5120
rect 18564 5108 18570 5160
rect 19426 5108 19432 5160
rect 19484 5108 19490 5160
rect 19904 5148 19932 5315
rect 24486 5312 24492 5324
rect 24544 5312 24550 5364
rect 27246 5352 27252 5364
rect 27207 5324 27252 5352
rect 27246 5312 27252 5324
rect 27304 5312 27310 5364
rect 28258 5312 28264 5364
rect 28316 5352 28322 5364
rect 28629 5355 28687 5361
rect 28629 5352 28641 5355
rect 28316 5324 28641 5352
rect 28316 5312 28322 5324
rect 28629 5321 28641 5324
rect 28675 5352 28687 5355
rect 28810 5352 28816 5364
rect 28675 5324 28816 5352
rect 28675 5321 28687 5324
rect 28629 5315 28687 5321
rect 28810 5312 28816 5324
rect 28868 5312 28874 5364
rect 29362 5312 29368 5364
rect 29420 5352 29426 5364
rect 29457 5355 29515 5361
rect 29457 5352 29469 5355
rect 29420 5324 29469 5352
rect 29420 5312 29426 5324
rect 29457 5321 29469 5324
rect 29503 5321 29515 5355
rect 29457 5315 29515 5321
rect 31754 5312 31760 5364
rect 31812 5352 31818 5364
rect 31812 5324 31857 5352
rect 31812 5312 31818 5324
rect 34790 5312 34796 5364
rect 34848 5352 34854 5364
rect 35161 5355 35219 5361
rect 35161 5352 35173 5355
rect 34848 5324 35173 5352
rect 34848 5312 34854 5324
rect 35161 5321 35173 5324
rect 35207 5321 35219 5355
rect 36998 5352 37004 5364
rect 35161 5315 35219 5321
rect 36096 5324 37004 5352
rect 22462 5284 22468 5296
rect 22388 5256 22468 5284
rect 22388 5225 22416 5256
rect 22462 5244 22468 5256
rect 22520 5244 22526 5296
rect 22373 5219 22431 5225
rect 22373 5185 22385 5219
rect 22419 5185 22431 5219
rect 22373 5179 22431 5185
rect 24949 5219 25007 5225
rect 24949 5185 24961 5219
rect 24995 5216 25007 5219
rect 26510 5216 26516 5228
rect 24995 5188 26516 5216
rect 24995 5185 25007 5188
rect 24949 5179 25007 5185
rect 26510 5176 26516 5188
rect 26568 5176 26574 5228
rect 30377 5219 30435 5225
rect 30377 5185 30389 5219
rect 30423 5216 30435 5219
rect 30558 5216 30564 5228
rect 30423 5188 30564 5216
rect 30423 5185 30435 5188
rect 30377 5179 30435 5185
rect 30558 5176 30564 5188
rect 30616 5216 30622 5228
rect 31386 5216 31392 5228
rect 30616 5188 31392 5216
rect 30616 5176 30622 5188
rect 31386 5176 31392 5188
rect 31444 5176 31450 5228
rect 31772 5216 31800 5312
rect 31846 5244 31852 5296
rect 31904 5284 31910 5296
rect 31904 5256 33548 5284
rect 31904 5244 31910 5256
rect 33520 5225 33548 5256
rect 34606 5244 34612 5296
rect 34664 5284 34670 5296
rect 36096 5284 36124 5324
rect 36998 5312 37004 5324
rect 37056 5352 37062 5364
rect 37461 5355 37519 5361
rect 37461 5352 37473 5355
rect 37056 5324 37473 5352
rect 37056 5312 37062 5324
rect 37461 5321 37473 5324
rect 37507 5321 37519 5355
rect 37461 5315 37519 5321
rect 38010 5312 38016 5364
rect 38068 5352 38074 5364
rect 38289 5355 38347 5361
rect 38289 5352 38301 5355
rect 38068 5324 38301 5352
rect 38068 5312 38074 5324
rect 38289 5321 38301 5324
rect 38335 5321 38347 5355
rect 38289 5315 38347 5321
rect 34664 5256 36124 5284
rect 34664 5244 34670 5256
rect 33505 5219 33563 5225
rect 31772 5188 33364 5216
rect 20625 5151 20683 5157
rect 20625 5148 20637 5151
rect 19904 5120 20637 5148
rect 20625 5117 20637 5120
rect 20671 5117 20683 5151
rect 20625 5111 20683 5117
rect 22005 5151 22063 5157
rect 22005 5117 22017 5151
rect 22051 5117 22063 5151
rect 22005 5111 22063 5117
rect 19444 5080 19472 5108
rect 20717 5083 20775 5089
rect 20717 5080 20729 5083
rect 19444 5052 20729 5080
rect 20717 5049 20729 5052
rect 20763 5049 20775 5083
rect 22020 5080 22048 5111
rect 22094 5108 22100 5160
rect 22152 5148 22158 5160
rect 22738 5148 22744 5160
rect 22152 5120 22197 5148
rect 22699 5120 22744 5148
rect 22152 5108 22158 5120
rect 22738 5108 22744 5120
rect 22796 5108 22802 5160
rect 22830 5108 22836 5160
rect 22888 5148 22894 5160
rect 23661 5151 23719 5157
rect 23661 5148 23673 5151
rect 22888 5120 23673 5148
rect 22888 5108 22894 5120
rect 23661 5117 23673 5120
rect 23707 5117 23719 5151
rect 25222 5148 25228 5160
rect 25183 5120 25228 5148
rect 23661 5111 23719 5117
rect 25222 5108 25228 5120
rect 25280 5108 25286 5160
rect 25409 5151 25467 5157
rect 25409 5117 25421 5151
rect 25455 5148 25467 5151
rect 25498 5148 25504 5160
rect 25455 5120 25504 5148
rect 25455 5117 25467 5120
rect 25409 5111 25467 5117
rect 25498 5108 25504 5120
rect 25556 5108 25562 5160
rect 25774 5108 25780 5160
rect 25832 5148 25838 5160
rect 25869 5151 25927 5157
rect 25869 5148 25881 5151
rect 25832 5120 25881 5148
rect 25832 5108 25838 5120
rect 25869 5117 25881 5120
rect 25915 5117 25927 5151
rect 25869 5111 25927 5117
rect 26145 5151 26203 5157
rect 26145 5117 26157 5151
rect 26191 5148 26203 5151
rect 26602 5148 26608 5160
rect 26191 5120 26608 5148
rect 26191 5117 26203 5120
rect 26145 5111 26203 5117
rect 26602 5108 26608 5120
rect 26660 5108 26666 5160
rect 28445 5151 28503 5157
rect 28445 5117 28457 5151
rect 28491 5148 28503 5151
rect 29086 5148 29092 5160
rect 28491 5120 29092 5148
rect 28491 5117 28503 5120
rect 28445 5111 28503 5117
rect 29086 5108 29092 5120
rect 29144 5108 29150 5160
rect 29270 5148 29276 5160
rect 29231 5120 29276 5148
rect 29270 5108 29276 5120
rect 29328 5108 29334 5160
rect 30653 5151 30711 5157
rect 30653 5117 30665 5151
rect 30699 5148 30711 5151
rect 32122 5148 32128 5160
rect 30699 5120 32128 5148
rect 30699 5117 30711 5120
rect 30653 5111 30711 5117
rect 32122 5108 32128 5120
rect 32180 5108 32186 5160
rect 33336 5157 33364 5188
rect 33505 5185 33517 5219
rect 33551 5216 33563 5219
rect 33962 5216 33968 5228
rect 33551 5188 33968 5216
rect 33551 5185 33563 5188
rect 33505 5179 33563 5185
rect 33962 5176 33968 5188
rect 34020 5176 34026 5228
rect 34698 5176 34704 5228
rect 34756 5216 34762 5228
rect 34756 5188 35020 5216
rect 34756 5176 34762 5188
rect 33045 5151 33103 5157
rect 33045 5148 33057 5151
rect 32416 5120 33057 5148
rect 23106 5080 23112 5092
rect 22020 5052 23112 5080
rect 20717 5043 20775 5049
rect 23106 5040 23112 5052
rect 23164 5040 23170 5092
rect 24397 5083 24455 5089
rect 24397 5049 24409 5083
rect 24443 5080 24455 5083
rect 25590 5080 25596 5092
rect 24443 5052 25596 5080
rect 24443 5049 24455 5052
rect 24397 5043 24455 5049
rect 25590 5040 25596 5052
rect 25648 5040 25654 5092
rect 31478 5040 31484 5092
rect 31536 5080 31542 5092
rect 32416 5080 32444 5120
rect 33045 5117 33057 5120
rect 33091 5117 33103 5151
rect 33045 5111 33103 5117
rect 33321 5151 33379 5157
rect 33321 5117 33333 5151
rect 33367 5117 33379 5151
rect 33321 5111 33379 5117
rect 34514 5108 34520 5160
rect 34572 5148 34578 5160
rect 34992 5157 35020 5188
rect 35986 5176 35992 5228
rect 36044 5216 36050 5228
rect 36081 5219 36139 5225
rect 36081 5216 36093 5219
rect 36044 5188 36093 5216
rect 36044 5176 36050 5188
rect 36081 5185 36093 5188
rect 36127 5185 36139 5219
rect 36354 5216 36360 5228
rect 36315 5188 36360 5216
rect 36081 5179 36139 5185
rect 36354 5176 36360 5188
rect 36412 5176 36418 5228
rect 37826 5176 37832 5228
rect 37884 5216 37890 5228
rect 37884 5188 38792 5216
rect 37884 5176 37890 5188
rect 34885 5151 34943 5157
rect 34885 5148 34897 5151
rect 34572 5120 34897 5148
rect 34572 5108 34578 5120
rect 34885 5117 34897 5120
rect 34931 5117 34943 5151
rect 34885 5111 34943 5117
rect 34977 5151 35035 5157
rect 34977 5117 34989 5151
rect 35023 5117 35035 5151
rect 34977 5111 35035 5117
rect 37642 5108 37648 5160
rect 37700 5148 37706 5160
rect 38764 5157 38792 5188
rect 38197 5151 38255 5157
rect 38197 5148 38209 5151
rect 37700 5120 38209 5148
rect 37700 5108 37706 5120
rect 38197 5117 38209 5120
rect 38243 5117 38255 5151
rect 38197 5111 38255 5117
rect 38749 5151 38807 5157
rect 38749 5117 38761 5151
rect 38795 5117 38807 5151
rect 38749 5111 38807 5117
rect 31536 5052 32444 5080
rect 32493 5083 32551 5089
rect 31536 5040 31542 5052
rect 32493 5049 32505 5083
rect 32539 5080 32551 5083
rect 32674 5080 32680 5092
rect 32539 5052 32680 5080
rect 32539 5049 32551 5052
rect 32493 5043 32551 5049
rect 32674 5040 32680 5052
rect 32732 5040 32738 5092
rect 19426 5012 19432 5024
rect 17328 4984 19432 5012
rect 17221 4975 17279 4981
rect 19426 4972 19432 4984
rect 19484 4972 19490 5024
rect 1104 4922 39836 4944
rect 1104 4870 19606 4922
rect 19658 4870 19670 4922
rect 19722 4870 19734 4922
rect 19786 4870 19798 4922
rect 19850 4870 39836 4922
rect 1104 4848 39836 4870
rect 10410 4808 10416 4820
rect 10323 4780 10416 4808
rect 4522 4672 4528 4684
rect 4483 4644 4528 4672
rect 4522 4632 4528 4644
rect 4580 4632 4586 4684
rect 5166 4672 5172 4684
rect 5127 4644 5172 4672
rect 5166 4632 5172 4644
rect 5224 4632 5230 4684
rect 10336 4681 10364 4780
rect 10410 4768 10416 4780
rect 10468 4808 10474 4820
rect 10468 4780 14596 4808
rect 10468 4768 10474 4780
rect 10962 4740 10968 4752
rect 10888 4712 10968 4740
rect 10321 4675 10379 4681
rect 10321 4641 10333 4675
rect 10367 4641 10379 4675
rect 10321 4635 10379 4641
rect 10410 4632 10416 4684
rect 10468 4672 10474 4684
rect 10888 4681 10916 4712
rect 10962 4700 10968 4712
rect 11020 4700 11026 4752
rect 11425 4743 11483 4749
rect 11425 4709 11437 4743
rect 11471 4709 11483 4743
rect 11425 4703 11483 4709
rect 10873 4675 10931 4681
rect 10468 4644 10513 4672
rect 10468 4632 10474 4644
rect 10873 4641 10885 4675
rect 10919 4641 10931 4675
rect 11054 4672 11060 4684
rect 11015 4644 11060 4672
rect 10873 4635 10931 4641
rect 11054 4632 11060 4644
rect 11112 4632 11118 4684
rect 11440 4672 11468 4703
rect 12253 4675 12311 4681
rect 12253 4672 12265 4675
rect 11440 4644 12265 4672
rect 12253 4641 12265 4644
rect 12299 4641 12311 4675
rect 14182 4672 14188 4684
rect 14143 4644 14188 4672
rect 12253 4635 12311 4641
rect 14182 4632 14188 4644
rect 14240 4632 14246 4684
rect 4893 4607 4951 4613
rect 4893 4573 4905 4607
rect 4939 4604 4951 4607
rect 4982 4604 4988 4616
rect 4939 4576 4988 4604
rect 4939 4573 4951 4576
rect 4893 4567 4951 4573
rect 4982 4564 4988 4576
rect 5040 4564 5046 4616
rect 6822 4604 6828 4616
rect 6783 4576 6828 4604
rect 6822 4564 6828 4576
rect 6880 4564 6886 4616
rect 7101 4607 7159 4613
rect 7101 4573 7113 4607
rect 7147 4604 7159 4607
rect 9582 4604 9588 4616
rect 7147 4576 9588 4604
rect 7147 4573 7159 4576
rect 7101 4567 7159 4573
rect 9582 4564 9588 4576
rect 9640 4564 9646 4616
rect 11882 4564 11888 4616
rect 11940 4604 11946 4616
rect 11977 4607 12035 4613
rect 11977 4604 11989 4607
rect 11940 4576 11989 4604
rect 11940 4564 11946 4576
rect 11977 4573 11989 4576
rect 12023 4573 12035 4607
rect 11977 4567 12035 4573
rect 13906 4564 13912 4616
rect 13964 4604 13970 4616
rect 14090 4604 14096 4616
rect 13964 4576 14096 4604
rect 13964 4564 13970 4576
rect 14090 4564 14096 4576
rect 14148 4564 14154 4616
rect 14568 4536 14596 4780
rect 15010 4768 15016 4820
rect 15068 4808 15074 4820
rect 22462 4808 22468 4820
rect 15068 4780 22468 4808
rect 15068 4768 15074 4780
rect 22462 4768 22468 4780
rect 22520 4768 22526 4820
rect 22830 4808 22836 4820
rect 22791 4780 22836 4808
rect 22830 4768 22836 4780
rect 22888 4768 22894 4820
rect 29641 4811 29699 4817
rect 29641 4808 29653 4811
rect 29564 4780 29653 4808
rect 14645 4743 14703 4749
rect 14645 4709 14657 4743
rect 14691 4740 14703 4743
rect 20257 4743 20315 4749
rect 14691 4712 16436 4740
rect 14691 4709 14703 4712
rect 14645 4703 14703 4709
rect 15565 4675 15623 4681
rect 15565 4641 15577 4675
rect 15611 4672 15623 4675
rect 15654 4672 15660 4684
rect 15611 4644 15660 4672
rect 15611 4641 15623 4644
rect 15565 4635 15623 4641
rect 15654 4632 15660 4644
rect 15712 4632 15718 4684
rect 16298 4604 16304 4616
rect 16259 4576 16304 4604
rect 16298 4564 16304 4576
rect 16356 4564 16362 4616
rect 16408 4604 16436 4712
rect 20257 4709 20269 4743
rect 20303 4740 20315 4743
rect 20622 4740 20628 4752
rect 20303 4712 20628 4740
rect 20303 4709 20315 4712
rect 20257 4703 20315 4709
rect 20622 4700 20628 4712
rect 20680 4700 20686 4752
rect 16574 4672 16580 4684
rect 16535 4644 16580 4672
rect 16574 4632 16580 4644
rect 16632 4632 16638 4684
rect 18966 4672 18972 4684
rect 18927 4644 18972 4672
rect 18966 4632 18972 4644
rect 19024 4632 19030 4684
rect 19150 4632 19156 4684
rect 19208 4672 19214 4684
rect 19429 4675 19487 4681
rect 19429 4672 19441 4675
rect 19208 4644 19441 4672
rect 19208 4632 19214 4644
rect 19429 4641 19441 4644
rect 19475 4641 19487 4675
rect 19429 4635 19487 4641
rect 20165 4675 20223 4681
rect 20165 4641 20177 4675
rect 20211 4672 20223 4675
rect 22848 4672 22876 4768
rect 23106 4700 23112 4752
rect 23164 4740 23170 4752
rect 23164 4712 28212 4740
rect 23164 4700 23170 4712
rect 24394 4672 24400 4684
rect 20211 4644 22876 4672
rect 24355 4644 24400 4672
rect 20211 4641 20223 4644
rect 20165 4635 20223 4641
rect 24394 4632 24400 4644
rect 24452 4632 24458 4684
rect 24486 4632 24492 4684
rect 24544 4672 24550 4684
rect 24673 4675 24731 4681
rect 24673 4672 24685 4675
rect 24544 4644 24685 4672
rect 24544 4632 24550 4644
rect 24673 4641 24685 4644
rect 24719 4641 24731 4675
rect 24673 4635 24731 4641
rect 24762 4632 24768 4684
rect 24820 4672 24826 4684
rect 24857 4675 24915 4681
rect 24857 4672 24869 4675
rect 24820 4644 24869 4672
rect 24820 4632 24826 4644
rect 24857 4641 24869 4644
rect 24903 4672 24915 4675
rect 24903 4644 27292 4672
rect 24903 4641 24915 4644
rect 24857 4635 24915 4641
rect 19702 4604 19708 4616
rect 16408 4576 18092 4604
rect 19663 4576 19708 4604
rect 15749 4539 15807 4545
rect 15749 4536 15761 4539
rect 14568 4508 15761 4536
rect 15749 4505 15761 4508
rect 15795 4536 15807 4539
rect 16206 4536 16212 4548
rect 15795 4508 16212 4536
rect 15795 4505 15807 4508
rect 15749 4499 15807 4505
rect 16206 4496 16212 4508
rect 16264 4496 16270 4548
rect 18064 4536 18092 4576
rect 19702 4564 19708 4576
rect 19760 4564 19766 4616
rect 21266 4604 21272 4616
rect 21227 4576 21272 4604
rect 21266 4564 21272 4576
rect 21324 4564 21330 4616
rect 21545 4607 21603 4613
rect 21545 4573 21557 4607
rect 21591 4604 21603 4607
rect 22830 4604 22836 4616
rect 21591 4576 22836 4604
rect 21591 4573 21603 4576
rect 21545 4567 21603 4573
rect 22830 4564 22836 4576
rect 22888 4564 22894 4616
rect 23842 4604 23848 4616
rect 23803 4576 23848 4604
rect 23842 4564 23848 4576
rect 23900 4564 23906 4616
rect 26510 4604 26516 4616
rect 26471 4576 26516 4604
rect 26510 4564 26516 4576
rect 26568 4564 26574 4616
rect 27062 4604 27068 4616
rect 27023 4576 27068 4604
rect 27062 4564 27068 4576
rect 27120 4564 27126 4616
rect 27264 4604 27292 4644
rect 27338 4632 27344 4684
rect 27396 4672 27402 4684
rect 27396 4644 27441 4672
rect 27396 4632 27402 4644
rect 27890 4632 27896 4684
rect 27948 4672 27954 4684
rect 28077 4675 28135 4681
rect 28077 4672 28089 4675
rect 27948 4644 28089 4672
rect 27948 4632 27954 4644
rect 28077 4641 28089 4644
rect 28123 4641 28135 4675
rect 28184 4672 28212 4712
rect 29270 4672 29276 4684
rect 28184 4644 29276 4672
rect 28077 4635 28135 4641
rect 29270 4632 29276 4644
rect 29328 4672 29334 4684
rect 29564 4672 29592 4780
rect 29641 4777 29653 4780
rect 29687 4777 29699 4811
rect 29641 4771 29699 4777
rect 37001 4811 37059 4817
rect 37001 4777 37013 4811
rect 37047 4808 37059 4811
rect 38194 4808 38200 4820
rect 37047 4780 38200 4808
rect 37047 4777 37059 4780
rect 37001 4771 37059 4777
rect 38194 4768 38200 4780
rect 38252 4768 38258 4820
rect 32122 4740 32128 4752
rect 32083 4712 32128 4740
rect 32122 4700 32128 4712
rect 32180 4700 32186 4752
rect 33410 4700 33416 4752
rect 33468 4740 33474 4752
rect 33468 4712 34468 4740
rect 33468 4700 33474 4712
rect 29328 4644 29592 4672
rect 29328 4632 29334 4644
rect 29730 4632 29736 4684
rect 29788 4672 29794 4684
rect 30745 4675 30803 4681
rect 30745 4672 30757 4675
rect 29788 4644 30757 4672
rect 29788 4632 29794 4644
rect 30745 4641 30757 4644
rect 30791 4641 30803 4675
rect 30745 4635 30803 4641
rect 31021 4675 31079 4681
rect 31021 4641 31033 4675
rect 31067 4672 31079 4675
rect 32030 4672 32036 4684
rect 31067 4644 32036 4672
rect 31067 4641 31079 4644
rect 31021 4635 31079 4641
rect 32030 4632 32036 4644
rect 32088 4632 32094 4684
rect 32674 4672 32680 4684
rect 32635 4644 32680 4672
rect 32674 4632 32680 4644
rect 32732 4632 32738 4684
rect 34330 4681 34336 4684
rect 32953 4675 33011 4681
rect 32953 4641 32965 4675
rect 32999 4672 33011 4675
rect 34287 4675 34336 4681
rect 34287 4672 34299 4675
rect 32999 4644 34299 4672
rect 32999 4641 33011 4644
rect 32953 4635 33011 4641
rect 34287 4641 34299 4644
rect 34333 4641 34336 4675
rect 34287 4635 34336 4641
rect 34330 4632 34336 4635
rect 34388 4632 34394 4684
rect 34440 4681 34468 4712
rect 34425 4675 34483 4681
rect 34425 4641 34437 4675
rect 34471 4641 34483 4675
rect 34425 4635 34483 4641
rect 35897 4675 35955 4681
rect 35897 4641 35909 4675
rect 35943 4641 35955 4675
rect 36078 4672 36084 4684
rect 36039 4644 36084 4672
rect 35897 4635 35955 4641
rect 27525 4607 27583 4613
rect 27525 4604 27537 4607
rect 27264 4576 27537 4604
rect 27525 4573 27537 4576
rect 27571 4604 27583 4607
rect 28258 4604 28264 4616
rect 27571 4576 28264 4604
rect 27571 4573 27583 4576
rect 27525 4567 27583 4573
rect 28258 4564 28264 4576
rect 28316 4564 28322 4616
rect 28353 4607 28411 4613
rect 28353 4573 28365 4607
rect 28399 4604 28411 4607
rect 30193 4607 30251 4613
rect 30193 4604 30205 4607
rect 28399 4576 30205 4604
rect 28399 4573 28411 4576
rect 28353 4567 28411 4573
rect 30193 4573 30205 4576
rect 30239 4573 30251 4607
rect 30193 4567 30251 4573
rect 30374 4564 30380 4616
rect 30432 4604 30438 4616
rect 31205 4607 31263 4613
rect 31205 4604 31217 4607
rect 30432 4576 31217 4604
rect 30432 4564 30438 4576
rect 31205 4573 31217 4576
rect 31251 4604 31263 4607
rect 31662 4604 31668 4616
rect 31251 4576 31668 4604
rect 31251 4573 31263 4576
rect 31205 4567 31263 4573
rect 31662 4564 31668 4576
rect 31720 4604 31726 4616
rect 32815 4607 32873 4613
rect 32815 4604 32827 4607
rect 31720 4576 31800 4604
rect 31720 4564 31726 4576
rect 31772 4536 31800 4576
rect 32416 4576 32827 4604
rect 32416 4536 32444 4576
rect 32815 4573 32827 4576
rect 32861 4573 32873 4607
rect 32815 4567 32873 4573
rect 33597 4607 33655 4613
rect 33597 4573 33609 4607
rect 33643 4573 33655 4607
rect 33597 4567 33655 4573
rect 34149 4607 34207 4613
rect 34149 4573 34161 4607
rect 34195 4604 34207 4607
rect 34514 4604 34520 4616
rect 34195 4576 34520 4604
rect 34195 4573 34207 4576
rect 34149 4567 34207 4573
rect 18064 4508 20392 4536
rect 31772 4508 32444 4536
rect 7558 4428 7564 4480
rect 7616 4468 7622 4480
rect 8205 4471 8263 4477
rect 8205 4468 8217 4471
rect 7616 4440 8217 4468
rect 7616 4428 7622 4440
rect 8205 4437 8217 4440
rect 8251 4437 8263 4471
rect 8205 4431 8263 4437
rect 12342 4428 12348 4480
rect 12400 4468 12406 4480
rect 13357 4471 13415 4477
rect 13357 4468 13369 4471
rect 12400 4440 13369 4468
rect 12400 4428 12406 4440
rect 13357 4437 13369 4440
rect 13403 4437 13415 4471
rect 13357 4431 13415 4437
rect 15562 4428 15568 4480
rect 15620 4468 15626 4480
rect 16482 4468 16488 4480
rect 15620 4440 16488 4468
rect 15620 4428 15626 4440
rect 16482 4428 16488 4440
rect 16540 4468 16546 4480
rect 17770 4468 17776 4480
rect 16540 4440 17776 4468
rect 16540 4428 16546 4440
rect 17770 4428 17776 4440
rect 17828 4428 17834 4480
rect 17865 4471 17923 4477
rect 17865 4437 17877 4471
rect 17911 4468 17923 4471
rect 18046 4468 18052 4480
rect 17911 4440 18052 4468
rect 17911 4437 17923 4440
rect 17865 4431 17923 4437
rect 18046 4428 18052 4440
rect 18104 4428 18110 4480
rect 20364 4468 20392 4508
rect 30006 4468 30012 4480
rect 20364 4440 30012 4468
rect 30006 4428 30012 4440
rect 30064 4428 30070 4480
rect 30834 4428 30840 4480
rect 30892 4468 30898 4480
rect 33612 4468 33640 4567
rect 34514 4564 34520 4576
rect 34572 4564 34578 4616
rect 34698 4564 34704 4616
rect 34756 4604 34762 4616
rect 35069 4607 35127 4613
rect 35069 4604 35081 4607
rect 34756 4576 35081 4604
rect 34756 4564 34762 4576
rect 35069 4573 35081 4576
rect 35115 4573 35127 4607
rect 35618 4604 35624 4616
rect 35579 4576 35624 4604
rect 35069 4567 35127 4573
rect 35618 4564 35624 4576
rect 35676 4564 35682 4616
rect 35912 4604 35940 4635
rect 36078 4632 36084 4644
rect 36136 4632 36142 4684
rect 36909 4675 36967 4681
rect 36909 4641 36921 4675
rect 36955 4672 36967 4675
rect 37642 4672 37648 4684
rect 36955 4644 37648 4672
rect 36955 4641 36967 4644
rect 36909 4635 36967 4641
rect 37642 4632 37648 4644
rect 37700 4632 37706 4684
rect 35986 4604 35992 4616
rect 35912 4576 35992 4604
rect 35986 4564 35992 4576
rect 36044 4604 36050 4616
rect 36262 4604 36268 4616
rect 36044 4576 36268 4604
rect 36044 4564 36050 4576
rect 36262 4564 36268 4576
rect 36320 4564 36326 4616
rect 30892 4440 33640 4468
rect 30892 4428 30898 4440
rect 1104 4378 39836 4400
rect 1104 4326 4246 4378
rect 4298 4326 4310 4378
rect 4362 4326 4374 4378
rect 4426 4326 4438 4378
rect 4490 4326 34966 4378
rect 35018 4326 35030 4378
rect 35082 4326 35094 4378
rect 35146 4326 35158 4378
rect 35210 4326 39836 4378
rect 1104 4304 39836 4326
rect 10410 4224 10416 4276
rect 10468 4264 10474 4276
rect 20898 4264 20904 4276
rect 10468 4236 20904 4264
rect 10468 4224 10474 4236
rect 20898 4224 20904 4236
rect 20956 4224 20962 4276
rect 35986 4264 35992 4276
rect 34256 4236 35992 4264
rect 16390 4156 16396 4208
rect 16448 4196 16454 4208
rect 18141 4199 18199 4205
rect 18141 4196 18153 4199
rect 16448 4168 18153 4196
rect 16448 4156 16454 4168
rect 18141 4165 18153 4168
rect 18187 4196 18199 4199
rect 19150 4196 19156 4208
rect 18187 4168 19156 4196
rect 18187 4165 18199 4168
rect 18141 4159 18199 4165
rect 19150 4156 19156 4168
rect 19208 4156 19214 4208
rect 24854 4156 24860 4208
rect 24912 4196 24918 4208
rect 25498 4196 25504 4208
rect 24912 4168 25504 4196
rect 24912 4156 24918 4168
rect 25498 4156 25504 4168
rect 25556 4196 25562 4208
rect 28350 4196 28356 4208
rect 25556 4168 28356 4196
rect 25556 4156 25562 4168
rect 4341 4131 4399 4137
rect 4341 4097 4353 4131
rect 4387 4128 4399 4131
rect 4798 4128 4804 4140
rect 4387 4100 4804 4128
rect 4387 4097 4399 4100
rect 4341 4091 4399 4097
rect 4798 4088 4804 4100
rect 4856 4088 4862 4140
rect 4890 4088 4896 4140
rect 4948 4128 4954 4140
rect 5077 4131 5135 4137
rect 5077 4128 5089 4131
rect 4948 4100 5089 4128
rect 4948 4088 4954 4100
rect 5077 4097 5089 4100
rect 5123 4097 5135 4131
rect 6270 4128 6276 4140
rect 6231 4100 6276 4128
rect 5077 4091 5135 4097
rect 6270 4088 6276 4100
rect 6328 4088 6334 4140
rect 7469 4131 7527 4137
rect 7469 4097 7481 4131
rect 7515 4128 7527 4131
rect 9674 4128 9680 4140
rect 7515 4100 9680 4128
rect 7515 4097 7527 4100
rect 7469 4091 7527 4097
rect 9674 4088 9680 4100
rect 9732 4088 9738 4140
rect 11072 4100 12848 4128
rect 4614 4060 4620 4072
rect 4575 4032 4620 4060
rect 4614 4020 4620 4032
rect 4672 4020 4678 4072
rect 4816 4060 4844 4088
rect 5537 4063 5595 4069
rect 5537 4060 5549 4063
rect 4816 4032 5549 4060
rect 5537 4029 5549 4032
rect 5583 4029 5595 4063
rect 5810 4060 5816 4072
rect 5771 4032 5816 4060
rect 5537 4023 5595 4029
rect 5810 4020 5816 4032
rect 5868 4020 5874 4072
rect 7558 4060 7564 4072
rect 7519 4032 7564 4060
rect 7558 4020 7564 4032
rect 7616 4020 7622 4072
rect 8478 4060 8484 4072
rect 7668 4032 8484 4060
rect 4525 3995 4583 4001
rect 4525 3961 4537 3995
rect 4571 3992 4583 3995
rect 4706 3992 4712 4004
rect 4571 3964 4712 3992
rect 4571 3961 4583 3964
rect 4525 3955 4583 3961
rect 4706 3952 4712 3964
rect 4764 3952 4770 4004
rect 4982 3952 4988 4004
rect 5040 3992 5046 4004
rect 5721 3995 5779 4001
rect 5721 3992 5733 3995
rect 5040 3964 5733 3992
rect 5040 3952 5046 3964
rect 5721 3961 5733 3964
rect 5767 3961 5779 3995
rect 5721 3955 5779 3961
rect 6822 3952 6828 4004
rect 6880 3992 6886 4004
rect 7668 3992 7696 4032
rect 8478 4020 8484 4032
rect 8536 4020 8542 4072
rect 8754 4060 8760 4072
rect 8715 4032 8760 4060
rect 8754 4020 8760 4032
rect 8812 4020 8818 4072
rect 10962 4020 10968 4072
rect 11020 4060 11026 4072
rect 11072 4069 11100 4100
rect 12820 4072 12848 4100
rect 13814 4088 13820 4140
rect 13872 4128 13878 4140
rect 14001 4131 14059 4137
rect 14001 4128 14013 4131
rect 13872 4100 14013 4128
rect 13872 4088 13878 4100
rect 14001 4097 14013 4100
rect 14047 4097 14059 4131
rect 14274 4128 14280 4140
rect 14235 4100 14280 4128
rect 14001 4091 14059 4097
rect 11057 4063 11115 4069
rect 11057 4060 11069 4063
rect 11020 4032 11069 4060
rect 11020 4020 11026 4032
rect 11057 4029 11069 4032
rect 11103 4029 11115 4063
rect 11238 4060 11244 4072
rect 11199 4032 11244 4060
rect 11057 4023 11115 4029
rect 11238 4020 11244 4032
rect 11296 4020 11302 4072
rect 12802 4060 12808 4072
rect 12763 4032 12808 4060
rect 12802 4020 12808 4032
rect 12860 4020 12866 4072
rect 13357 4063 13415 4069
rect 13357 4029 13369 4063
rect 13403 4029 13415 4063
rect 14016 4060 14044 4091
rect 14274 4088 14280 4100
rect 14332 4088 14338 4140
rect 15286 4088 15292 4140
rect 15344 4128 15350 4140
rect 15381 4131 15439 4137
rect 15381 4128 15393 4131
rect 15344 4100 15393 4128
rect 15344 4088 15350 4100
rect 15381 4097 15393 4100
rect 15427 4097 15439 4131
rect 18966 4128 18972 4140
rect 15381 4091 15439 4097
rect 16684 4100 18972 4128
rect 16684 4072 16712 4100
rect 16298 4060 16304 4072
rect 14016 4032 16304 4060
rect 13357 4023 13415 4029
rect 6880 3964 7696 3992
rect 6880 3952 6886 3964
rect 7742 3952 7748 4004
rect 7800 3992 7806 4004
rect 8021 3995 8079 4001
rect 8021 3992 8033 3995
rect 7800 3964 8033 3992
rect 7800 3952 7806 3964
rect 8021 3961 8033 3964
rect 8067 3961 8079 3995
rect 10134 3992 10140 4004
rect 10095 3964 10140 3992
rect 8021 3955 8079 3961
rect 10134 3952 10140 3964
rect 10192 3952 10198 4004
rect 7466 3884 7472 3936
rect 7524 3924 7530 3936
rect 10873 3927 10931 3933
rect 10873 3924 10885 3927
rect 7524 3896 10885 3924
rect 7524 3884 7530 3896
rect 10873 3893 10885 3896
rect 10919 3893 10931 3927
rect 13372 3924 13400 4023
rect 16298 4020 16304 4032
rect 16356 4020 16362 4072
rect 16666 4060 16672 4072
rect 16627 4032 16672 4060
rect 16666 4020 16672 4032
rect 16724 4020 16730 4072
rect 17034 4060 17040 4072
rect 16995 4032 17040 4060
rect 17034 4020 17040 4032
rect 17092 4020 17098 4072
rect 18046 4060 18052 4072
rect 18007 4032 18052 4060
rect 18046 4020 18052 4032
rect 18104 4020 18110 4072
rect 18800 4069 18828 4100
rect 18966 4088 18972 4100
rect 19024 4088 19030 4140
rect 19702 4088 19708 4140
rect 19760 4128 19766 4140
rect 20257 4131 20315 4137
rect 20257 4128 20269 4131
rect 19760 4100 20269 4128
rect 19760 4088 19766 4100
rect 20257 4097 20269 4100
rect 20303 4097 20315 4131
rect 20257 4091 20315 4097
rect 20714 4088 20720 4140
rect 20772 4128 20778 4140
rect 20772 4100 22784 4128
rect 20772 4088 20778 4100
rect 18785 4063 18843 4069
rect 18785 4029 18797 4063
rect 18831 4029 18843 4063
rect 19334 4060 19340 4072
rect 19295 4032 19340 4060
rect 18785 4023 18843 4029
rect 19334 4020 19340 4032
rect 19392 4020 19398 4072
rect 19981 4063 20039 4069
rect 19981 4029 19993 4063
rect 20027 4060 20039 4063
rect 20346 4060 20352 4072
rect 20027 4032 20352 4060
rect 20027 4029 20039 4032
rect 19981 4023 20039 4029
rect 20346 4020 20352 4032
rect 20404 4020 20410 4072
rect 22094 4060 22100 4072
rect 22055 4032 22100 4060
rect 22094 4020 22100 4032
rect 22152 4020 22158 4072
rect 22189 4063 22247 4069
rect 22189 4029 22201 4063
rect 22235 4029 22247 4063
rect 22189 4023 22247 4029
rect 13538 3992 13544 4004
rect 13499 3964 13544 3992
rect 13538 3952 13544 3964
rect 13596 3952 13602 4004
rect 19521 3995 19579 4001
rect 19521 3961 19533 3995
rect 19567 3961 19579 3995
rect 19521 3955 19579 3961
rect 14550 3924 14556 3936
rect 13372 3896 14556 3924
rect 10873 3887 10931 3893
rect 14550 3884 14556 3896
rect 14608 3884 14614 3936
rect 16114 3884 16120 3936
rect 16172 3924 16178 3936
rect 16577 3927 16635 3933
rect 16577 3924 16589 3927
rect 16172 3896 16589 3924
rect 16172 3884 16178 3896
rect 16577 3893 16589 3896
rect 16623 3893 16635 3927
rect 19536 3924 19564 3955
rect 20622 3924 20628 3936
rect 19536 3896 20628 3924
rect 16577 3887 16635 3893
rect 20622 3884 20628 3896
rect 20680 3884 20686 3936
rect 21545 3927 21603 3933
rect 21545 3893 21557 3927
rect 21591 3924 21603 3927
rect 22204 3924 22232 4023
rect 22649 3995 22707 4001
rect 22649 3961 22661 3995
rect 22695 3961 22707 3995
rect 22756 3992 22784 4100
rect 22830 4088 22836 4140
rect 22888 4128 22894 4140
rect 23661 4131 23719 4137
rect 23661 4128 23673 4131
rect 22888 4100 23673 4128
rect 22888 4088 22894 4100
rect 23661 4097 23673 4100
rect 23707 4097 23719 4131
rect 23661 4091 23719 4097
rect 23842 4088 23848 4140
rect 23900 4128 23906 4140
rect 24213 4131 24271 4137
rect 24213 4128 24225 4131
rect 23900 4100 24225 4128
rect 23900 4088 23906 4100
rect 24213 4097 24225 4100
rect 24259 4097 24271 4131
rect 24213 4091 24271 4097
rect 24320 4100 24992 4128
rect 23474 4020 23480 4072
rect 23532 4060 23538 4072
rect 24320 4060 24348 4100
rect 24486 4060 24492 4072
rect 23532 4032 24348 4060
rect 24447 4032 24492 4060
rect 23532 4020 23538 4032
rect 24486 4020 24492 4032
rect 24544 4020 24550 4072
rect 24673 4063 24731 4069
rect 24673 4029 24685 4063
rect 24719 4060 24731 4063
rect 24854 4060 24860 4072
rect 24719 4032 24860 4060
rect 24719 4029 24731 4032
rect 24673 4023 24731 4029
rect 24854 4020 24860 4032
rect 24912 4020 24918 4072
rect 24964 4060 24992 4100
rect 25038 4088 25044 4140
rect 25096 4128 25102 4140
rect 25133 4131 25191 4137
rect 25133 4128 25145 4131
rect 25096 4100 25145 4128
rect 25096 4088 25102 4100
rect 25133 4097 25145 4100
rect 25179 4097 25191 4131
rect 25133 4091 25191 4097
rect 25406 4088 25412 4140
rect 25464 4128 25470 4140
rect 26160 4137 26188 4168
rect 25685 4131 25743 4137
rect 25685 4128 25697 4131
rect 25464 4100 25697 4128
rect 25464 4088 25470 4100
rect 25685 4097 25697 4100
rect 25731 4097 25743 4131
rect 25685 4091 25743 4097
rect 26145 4131 26203 4137
rect 26145 4097 26157 4131
rect 26191 4097 26203 4131
rect 26145 4091 26203 4097
rect 26510 4088 26516 4140
rect 26568 4128 26574 4140
rect 27632 4137 27660 4168
rect 28350 4156 28356 4168
rect 28408 4156 28414 4208
rect 34256 4205 34284 4236
rect 35986 4224 35992 4236
rect 36044 4224 36050 4276
rect 34241 4199 34299 4205
rect 34241 4196 34253 4199
rect 34072 4168 34253 4196
rect 27157 4131 27215 4137
rect 27157 4128 27169 4131
rect 26568 4100 27169 4128
rect 26568 4088 26574 4100
rect 27157 4097 27169 4100
rect 27203 4097 27215 4131
rect 27157 4091 27215 4097
rect 27617 4131 27675 4137
rect 27617 4097 27629 4131
rect 27663 4097 27675 4131
rect 27617 4091 27675 4097
rect 29549 4131 29607 4137
rect 29549 4097 29561 4131
rect 29595 4128 29607 4131
rect 30374 4128 30380 4140
rect 29595 4100 30380 4128
rect 29595 4097 29607 4100
rect 29549 4091 29607 4097
rect 30374 4088 30380 4100
rect 30432 4088 30438 4140
rect 30558 4128 30564 4140
rect 30519 4100 30564 4128
rect 30558 4088 30564 4100
rect 30616 4088 30622 4140
rect 30834 4128 30840 4140
rect 30795 4100 30840 4128
rect 30834 4088 30840 4100
rect 30892 4088 30898 4140
rect 33594 4088 33600 4140
rect 33652 4128 33658 4140
rect 34072 4128 34100 4168
rect 34241 4165 34253 4168
rect 34287 4165 34299 4199
rect 34241 4159 34299 4165
rect 34624 4168 35756 4196
rect 34624 4140 34652 4168
rect 34606 4128 34612 4140
rect 33652 4100 34100 4128
rect 34164 4100 34612 4128
rect 33652 4088 33658 4100
rect 25961 4063 26019 4069
rect 25961 4060 25973 4063
rect 24964 4032 25973 4060
rect 25961 4029 25973 4032
rect 26007 4029 26019 4063
rect 26602 4060 26608 4072
rect 26563 4032 26608 4060
rect 25961 4023 26019 4029
rect 26602 4020 26608 4032
rect 26660 4020 26666 4072
rect 27430 4060 27436 4072
rect 27391 4032 27436 4060
rect 27430 4020 27436 4032
rect 27488 4020 27494 4072
rect 29086 4020 29092 4072
rect 29144 4060 29150 4072
rect 29457 4063 29515 4069
rect 29457 4060 29469 4063
rect 29144 4032 29469 4060
rect 29144 4020 29150 4032
rect 29457 4029 29469 4032
rect 29503 4029 29515 4063
rect 32582 4060 32588 4072
rect 29457 4023 29515 4029
rect 30668 4032 32588 4060
rect 22756 3964 27292 3992
rect 22649 3955 22707 3961
rect 21591 3896 22232 3924
rect 22664 3924 22692 3955
rect 27154 3924 27160 3936
rect 22664 3896 27160 3924
rect 21591 3893 21603 3896
rect 21545 3887 21603 3893
rect 27154 3884 27160 3896
rect 27212 3884 27218 3936
rect 27264 3924 27292 3964
rect 27522 3952 27528 4004
rect 27580 3992 27586 4004
rect 30668 3992 30696 4032
rect 32582 4020 32588 4032
rect 32640 4020 32646 4072
rect 33226 4060 33232 4072
rect 33187 4032 33232 4060
rect 33226 4020 33232 4032
rect 33284 4020 33290 4072
rect 33410 4020 33416 4072
rect 33468 4060 33474 4072
rect 33505 4063 33563 4069
rect 33505 4060 33517 4063
rect 33468 4032 33517 4060
rect 33468 4020 33474 4032
rect 33505 4029 33517 4032
rect 33551 4029 33563 4063
rect 33686 4060 33692 4072
rect 33647 4032 33692 4060
rect 33505 4023 33563 4029
rect 33686 4020 33692 4032
rect 33744 4020 33750 4072
rect 33870 4020 33876 4072
rect 33928 4060 33934 4072
rect 34164 4069 34192 4100
rect 34606 4088 34612 4100
rect 34664 4088 34670 4140
rect 34885 4131 34943 4137
rect 34885 4097 34897 4131
rect 34931 4128 34943 4131
rect 35618 4128 35624 4140
rect 34931 4100 35624 4128
rect 34931 4097 34943 4100
rect 34885 4091 34943 4097
rect 35618 4088 35624 4100
rect 35676 4088 35682 4140
rect 34149 4063 34207 4069
rect 34149 4060 34161 4063
rect 33928 4032 34161 4060
rect 33928 4020 33934 4032
rect 34149 4029 34161 4032
rect 34195 4029 34207 4063
rect 34149 4023 34207 4029
rect 34422 4020 34428 4072
rect 34480 4060 34486 4072
rect 35728 4069 35756 4168
rect 38930 4128 38936 4140
rect 38891 4100 38936 4128
rect 38930 4088 38936 4100
rect 38988 4088 38994 4140
rect 35437 4063 35495 4069
rect 35437 4060 35449 4063
rect 34480 4032 35449 4060
rect 34480 4020 34486 4032
rect 35437 4029 35449 4032
rect 35483 4029 35495 4063
rect 35437 4023 35495 4029
rect 35713 4063 35771 4069
rect 35713 4029 35725 4063
rect 35759 4029 35771 4063
rect 35897 4063 35955 4069
rect 35897 4060 35909 4063
rect 35713 4023 35771 4029
rect 35820 4032 35909 4060
rect 32674 3992 32680 4004
rect 27580 3964 30696 3992
rect 32635 3964 32680 3992
rect 27580 3952 27586 3964
rect 32674 3952 32680 3964
rect 32732 3952 32738 4004
rect 34330 3952 34336 4004
rect 34388 3992 34394 4004
rect 35820 3992 35848 4032
rect 35897 4029 35909 4032
rect 35943 4029 35955 4063
rect 37461 4063 37519 4069
rect 37461 4060 37473 4063
rect 35897 4023 35955 4029
rect 36004 4032 37473 4060
rect 34388 3964 35848 3992
rect 34388 3952 34394 3964
rect 31294 3924 31300 3936
rect 27264 3896 31300 3924
rect 31294 3884 31300 3896
rect 31352 3884 31358 3936
rect 32030 3884 32036 3936
rect 32088 3924 32094 3936
rect 32125 3927 32183 3933
rect 32125 3924 32137 3927
rect 32088 3896 32137 3924
rect 32088 3884 32094 3896
rect 32125 3893 32137 3896
rect 32171 3924 32183 3927
rect 33686 3924 33692 3936
rect 32171 3896 33692 3924
rect 32171 3893 32183 3896
rect 32125 3887 32183 3893
rect 33686 3884 33692 3896
rect 33744 3884 33750 3936
rect 35434 3884 35440 3936
rect 35492 3924 35498 3936
rect 36004 3924 36032 4032
rect 37461 4029 37473 4032
rect 37507 4029 37519 4063
rect 37734 4060 37740 4072
rect 37695 4032 37740 4060
rect 37461 4023 37519 4029
rect 37734 4020 37740 4032
rect 37792 4020 37798 4072
rect 35492 3896 36032 3924
rect 35492 3884 35498 3896
rect 1104 3834 39836 3856
rect 1104 3782 19606 3834
rect 19658 3782 19670 3834
rect 19722 3782 19734 3834
rect 19786 3782 19798 3834
rect 19850 3782 39836 3834
rect 1104 3760 39836 3782
rect 9674 3680 9680 3732
rect 9732 3720 9738 3732
rect 14826 3720 14832 3732
rect 9732 3692 14832 3720
rect 9732 3680 9738 3692
rect 14826 3680 14832 3692
rect 14884 3680 14890 3732
rect 17034 3680 17040 3732
rect 17092 3720 17098 3732
rect 19797 3723 19855 3729
rect 19797 3720 19809 3723
rect 17092 3692 19809 3720
rect 17092 3680 17098 3692
rect 19797 3689 19809 3692
rect 19843 3689 19855 3723
rect 19797 3683 19855 3689
rect 23566 3680 23572 3732
rect 23624 3720 23630 3732
rect 25130 3720 25136 3732
rect 23624 3692 25136 3720
rect 23624 3680 23630 3692
rect 25130 3680 25136 3692
rect 25188 3680 25194 3732
rect 27430 3680 27436 3732
rect 27488 3720 27494 3732
rect 29641 3723 29699 3729
rect 29641 3720 29653 3723
rect 27488 3692 29653 3720
rect 27488 3680 27494 3692
rect 29641 3689 29653 3692
rect 29687 3720 29699 3723
rect 31202 3720 31208 3732
rect 29687 3692 31208 3720
rect 29687 3689 29699 3692
rect 29641 3683 29699 3689
rect 31202 3680 31208 3692
rect 31260 3680 31266 3732
rect 31294 3680 31300 3732
rect 31352 3720 31358 3732
rect 31352 3692 33916 3720
rect 31352 3680 31358 3692
rect 8754 3612 8760 3664
rect 8812 3652 8818 3664
rect 10229 3655 10287 3661
rect 10229 3652 10241 3655
rect 8812 3624 10241 3652
rect 8812 3612 8818 3624
rect 10229 3621 10241 3624
rect 10275 3621 10287 3655
rect 10229 3615 10287 3621
rect 24486 3612 24492 3664
rect 24544 3652 24550 3664
rect 24673 3655 24731 3661
rect 24673 3652 24685 3655
rect 24544 3624 24685 3652
rect 24544 3612 24550 3624
rect 24673 3621 24685 3624
rect 24719 3652 24731 3655
rect 24719 3624 27568 3652
rect 24719 3621 24731 3624
rect 24673 3615 24731 3621
rect 6822 3544 6828 3596
rect 6880 3584 6886 3596
rect 7193 3587 7251 3593
rect 7193 3584 7205 3587
rect 6880 3556 7205 3584
rect 6880 3544 6886 3556
rect 7193 3553 7205 3556
rect 7239 3553 7251 3587
rect 7466 3584 7472 3596
rect 7427 3556 7472 3584
rect 7193 3547 7251 3553
rect 7466 3544 7472 3556
rect 7524 3544 7530 3596
rect 8849 3587 8907 3593
rect 8849 3553 8861 3587
rect 8895 3584 8907 3587
rect 9769 3587 9827 3593
rect 9769 3584 9781 3587
rect 8895 3556 9781 3584
rect 8895 3553 8907 3556
rect 8849 3547 8907 3553
rect 9769 3553 9781 3556
rect 9815 3553 9827 3587
rect 10962 3584 10968 3596
rect 10923 3556 10968 3584
rect 9769 3547 9827 3553
rect 10962 3544 10968 3556
rect 11020 3544 11026 3596
rect 11333 3587 11391 3593
rect 11333 3553 11345 3587
rect 11379 3584 11391 3587
rect 12526 3584 12532 3596
rect 11379 3556 12532 3584
rect 11379 3553 11391 3556
rect 11333 3547 11391 3553
rect 12526 3544 12532 3556
rect 12584 3544 12590 3596
rect 13538 3544 13544 3596
rect 13596 3584 13602 3596
rect 15565 3587 15623 3593
rect 15565 3584 15577 3587
rect 13596 3556 15577 3584
rect 13596 3544 13602 3556
rect 15565 3553 15577 3556
rect 15611 3553 15623 3587
rect 15565 3547 15623 3553
rect 17218 3544 17224 3596
rect 17276 3584 17282 3596
rect 17865 3587 17923 3593
rect 17865 3584 17877 3587
rect 17276 3556 17877 3584
rect 17276 3544 17282 3556
rect 17865 3553 17877 3556
rect 17911 3553 17923 3587
rect 17865 3547 17923 3553
rect 19245 3587 19303 3593
rect 19245 3553 19257 3587
rect 19291 3584 19303 3587
rect 19705 3587 19763 3593
rect 19705 3584 19717 3587
rect 19291 3556 19717 3584
rect 19291 3553 19303 3556
rect 19245 3547 19303 3553
rect 19705 3553 19717 3556
rect 19751 3553 19763 3587
rect 22922 3584 22928 3596
rect 19705 3547 19763 3553
rect 20916 3556 22928 3584
rect 566 3476 572 3528
rect 624 3516 630 3528
rect 1762 3516 1768 3528
rect 624 3488 1768 3516
rect 624 3476 630 3488
rect 1762 3476 1768 3488
rect 1820 3476 1826 3528
rect 9674 3516 9680 3528
rect 9635 3488 9680 3516
rect 9674 3476 9680 3488
rect 9732 3476 9738 3528
rect 11241 3519 11299 3525
rect 11241 3516 11253 3519
rect 9784 3488 11253 3516
rect 9784 3460 9812 3488
rect 11241 3485 11253 3488
rect 11287 3485 11299 3519
rect 12434 3516 12440 3528
rect 12395 3488 12440 3516
rect 11241 3479 11299 3485
rect 12434 3476 12440 3488
rect 12492 3476 12498 3528
rect 12713 3519 12771 3525
rect 12713 3485 12725 3519
rect 12759 3516 12771 3519
rect 13170 3516 13176 3528
rect 12759 3488 13176 3516
rect 12759 3485 12771 3488
rect 12713 3479 12771 3485
rect 13170 3476 13176 3488
rect 13228 3476 13234 3528
rect 15286 3516 15292 3528
rect 15247 3488 15292 3516
rect 15286 3476 15292 3488
rect 15344 3476 15350 3528
rect 16298 3476 16304 3528
rect 16356 3516 16362 3528
rect 17589 3519 17647 3525
rect 17589 3516 17601 3519
rect 16356 3488 17601 3516
rect 16356 3476 16362 3488
rect 17589 3485 17601 3488
rect 17635 3516 17647 3519
rect 17954 3516 17960 3528
rect 17635 3488 17960 3516
rect 17635 3485 17647 3488
rect 17589 3479 17647 3485
rect 17954 3476 17960 3488
rect 18012 3476 18018 3528
rect 20346 3476 20352 3528
rect 20404 3516 20410 3528
rect 20916 3525 20944 3556
rect 22922 3544 22928 3556
rect 22980 3544 22986 3596
rect 23014 3544 23020 3596
rect 23072 3584 23078 3596
rect 25133 3587 25191 3593
rect 23072 3556 23117 3584
rect 23072 3544 23078 3556
rect 25133 3553 25145 3587
rect 25179 3584 25191 3587
rect 25590 3584 25596 3596
rect 25179 3556 25596 3584
rect 25179 3553 25191 3556
rect 25133 3547 25191 3553
rect 25590 3544 25596 3556
rect 25648 3544 25654 3596
rect 27341 3587 27399 3593
rect 27341 3584 27353 3587
rect 27264 3556 27353 3584
rect 20901 3519 20959 3525
rect 20901 3516 20913 3519
rect 20404 3488 20913 3516
rect 20404 3476 20410 3488
rect 20901 3485 20913 3488
rect 20947 3485 20959 3519
rect 20901 3479 20959 3485
rect 21082 3476 21088 3528
rect 21140 3516 21146 3528
rect 21177 3519 21235 3525
rect 21177 3516 21189 3519
rect 21140 3488 21189 3516
rect 21140 3476 21146 3488
rect 21177 3485 21189 3488
rect 21223 3485 21235 3519
rect 21177 3479 21235 3485
rect 23198 3476 23204 3528
rect 23256 3516 23262 3528
rect 23293 3519 23351 3525
rect 23293 3516 23305 3519
rect 23256 3488 23305 3516
rect 23256 3476 23262 3488
rect 23293 3485 23305 3488
rect 23339 3485 23351 3519
rect 23293 3479 23351 3485
rect 24578 3476 24584 3528
rect 24636 3516 24642 3528
rect 26513 3519 26571 3525
rect 26513 3516 26525 3519
rect 24636 3488 26525 3516
rect 24636 3476 24642 3488
rect 26513 3485 26525 3488
rect 26559 3485 26571 3519
rect 27062 3516 27068 3528
rect 27023 3488 27068 3516
rect 26513 3479 26571 3485
rect 27062 3476 27068 3488
rect 27120 3476 27126 3528
rect 8662 3408 8668 3460
rect 8720 3448 8726 3460
rect 8720 3420 9720 3448
rect 8720 3408 8726 3420
rect 9692 3380 9720 3420
rect 9766 3408 9772 3460
rect 9824 3408 9830 3460
rect 25225 3451 25283 3457
rect 25225 3448 25237 3451
rect 23952 3420 25237 3448
rect 12618 3380 12624 3392
rect 9692 3352 12624 3380
rect 12618 3340 12624 3352
rect 12676 3340 12682 3392
rect 14001 3383 14059 3389
rect 14001 3349 14013 3383
rect 14047 3380 14059 3383
rect 14090 3380 14096 3392
rect 14047 3352 14096 3380
rect 14047 3349 14059 3352
rect 14001 3343 14059 3349
rect 14090 3340 14096 3352
rect 14148 3340 14154 3392
rect 14918 3340 14924 3392
rect 14976 3380 14982 3392
rect 16669 3383 16727 3389
rect 16669 3380 16681 3383
rect 14976 3352 16681 3380
rect 14976 3340 14982 3352
rect 16669 3349 16681 3352
rect 16715 3349 16727 3383
rect 16669 3343 16727 3349
rect 22465 3383 22523 3389
rect 22465 3349 22477 3383
rect 22511 3380 22523 3383
rect 22554 3380 22560 3392
rect 22511 3352 22560 3380
rect 22511 3349 22523 3352
rect 22465 3343 22523 3349
rect 22554 3340 22560 3352
rect 22612 3340 22618 3392
rect 22646 3340 22652 3392
rect 22704 3380 22710 3392
rect 23952 3380 23980 3420
rect 25225 3417 25237 3420
rect 25271 3417 25283 3451
rect 25225 3411 25283 3417
rect 22704 3352 23980 3380
rect 22704 3340 22710 3352
rect 24394 3340 24400 3392
rect 24452 3380 24458 3392
rect 27264 3380 27292 3556
rect 27341 3553 27353 3556
rect 27387 3553 27399 3587
rect 27341 3547 27399 3553
rect 27540 3525 27568 3624
rect 27614 3612 27620 3664
rect 27672 3652 27678 3664
rect 27890 3652 27896 3664
rect 27672 3624 27896 3652
rect 27672 3612 27678 3624
rect 27890 3612 27896 3624
rect 27948 3652 27954 3664
rect 32674 3652 32680 3664
rect 27948 3624 28120 3652
rect 27948 3612 27954 3624
rect 28092 3593 28120 3624
rect 30852 3624 32680 3652
rect 28077 3587 28135 3593
rect 28077 3553 28089 3587
rect 28123 3553 28135 3587
rect 28077 3547 28135 3553
rect 28353 3587 28411 3593
rect 28353 3553 28365 3587
rect 28399 3584 28411 3587
rect 30852 3584 30880 3624
rect 32674 3612 32680 3624
rect 32732 3612 32738 3664
rect 28399 3556 30880 3584
rect 28399 3553 28411 3556
rect 28353 3547 28411 3553
rect 31018 3544 31024 3596
rect 31076 3584 31082 3596
rect 32217 3587 32275 3593
rect 31076 3556 31121 3584
rect 31076 3544 31082 3556
rect 32217 3553 32229 3587
rect 32263 3584 32275 3587
rect 33594 3584 33600 3596
rect 32263 3556 33600 3584
rect 32263 3553 32275 3556
rect 32217 3547 32275 3553
rect 33594 3544 33600 3556
rect 33652 3544 33658 3596
rect 33888 3584 33916 3692
rect 34330 3680 34336 3732
rect 34388 3720 34394 3732
rect 34517 3723 34575 3729
rect 34517 3720 34529 3723
rect 34388 3692 34529 3720
rect 34388 3680 34394 3692
rect 34517 3689 34529 3692
rect 34563 3689 34575 3723
rect 34517 3683 34575 3689
rect 35805 3587 35863 3593
rect 35805 3584 35817 3587
rect 33888 3556 35817 3584
rect 35805 3553 35817 3556
rect 35851 3553 35863 3587
rect 35805 3547 35863 3553
rect 27525 3519 27583 3525
rect 27525 3485 27537 3519
rect 27571 3516 27583 3519
rect 27890 3516 27896 3528
rect 27571 3488 27896 3516
rect 27571 3485 27583 3488
rect 27525 3479 27583 3485
rect 27890 3476 27896 3488
rect 27948 3476 27954 3528
rect 28258 3476 28264 3528
rect 28316 3516 28322 3528
rect 30193 3519 30251 3525
rect 30193 3516 30205 3519
rect 28316 3488 30205 3516
rect 28316 3476 28322 3488
rect 30193 3485 30205 3488
rect 30239 3485 30251 3519
rect 30193 3479 30251 3485
rect 30745 3519 30803 3525
rect 30745 3485 30757 3519
rect 30791 3485 30803 3519
rect 31202 3516 31208 3528
rect 31115 3488 31208 3516
rect 30745 3479 30803 3485
rect 29270 3408 29276 3460
rect 29328 3448 29334 3460
rect 30760 3448 30788 3479
rect 31202 3476 31208 3488
rect 31260 3516 31266 3528
rect 31662 3516 31668 3528
rect 31260 3488 31668 3516
rect 31260 3476 31266 3488
rect 31662 3476 31668 3488
rect 31720 3476 31726 3528
rect 32950 3516 32956 3528
rect 32911 3488 32956 3516
rect 32950 3476 32956 3488
rect 33008 3476 33014 3528
rect 33229 3519 33287 3525
rect 33229 3485 33241 3519
rect 33275 3516 33287 3519
rect 34698 3516 34704 3528
rect 33275 3488 34704 3516
rect 33275 3485 33287 3488
rect 33229 3479 33287 3485
rect 34698 3476 34704 3488
rect 34756 3476 34762 3528
rect 35529 3519 35587 3525
rect 35529 3516 35541 3519
rect 35452 3488 35541 3516
rect 29328 3420 30788 3448
rect 29328 3408 29334 3420
rect 35452 3392 35480 3488
rect 35529 3485 35541 3488
rect 35575 3485 35587 3519
rect 35529 3479 35587 3485
rect 31018 3380 31024 3392
rect 24452 3352 31024 3380
rect 24452 3340 24458 3352
rect 31018 3340 31024 3352
rect 31076 3380 31082 3392
rect 32401 3383 32459 3389
rect 32401 3380 32413 3383
rect 31076 3352 32413 3380
rect 31076 3340 31082 3352
rect 32401 3349 32413 3352
rect 32447 3380 32459 3383
rect 33410 3380 33416 3392
rect 32447 3352 33416 3380
rect 32447 3349 32459 3352
rect 32401 3343 32459 3349
rect 33410 3340 33416 3352
rect 33468 3340 33474 3392
rect 33594 3340 33600 3392
rect 33652 3380 33658 3392
rect 35434 3380 35440 3392
rect 33652 3352 35440 3380
rect 33652 3340 33658 3352
rect 35434 3340 35440 3352
rect 35492 3340 35498 3392
rect 37090 3380 37096 3392
rect 37051 3352 37096 3380
rect 37090 3340 37096 3352
rect 37148 3340 37154 3392
rect 1104 3290 39836 3312
rect 1104 3238 4246 3290
rect 4298 3238 4310 3290
rect 4362 3238 4374 3290
rect 4426 3238 4438 3290
rect 4490 3238 34966 3290
rect 35018 3238 35030 3290
rect 35082 3238 35094 3290
rect 35146 3238 35158 3290
rect 35210 3238 39836 3290
rect 1104 3216 39836 3238
rect 8018 3136 8024 3188
rect 8076 3176 8082 3188
rect 14001 3179 14059 3185
rect 8076 3148 13952 3176
rect 8076 3136 8082 3148
rect 8478 3068 8484 3120
rect 8536 3108 8542 3120
rect 9398 3108 9404 3120
rect 8536 3080 9404 3108
rect 8536 3068 8542 3080
rect 9398 3068 9404 3080
rect 9456 3068 9462 3120
rect 11054 3068 11060 3120
rect 11112 3108 11118 3120
rect 11793 3111 11851 3117
rect 11793 3108 11805 3111
rect 11112 3080 11805 3108
rect 11112 3068 11118 3080
rect 11793 3077 11805 3080
rect 11839 3077 11851 3111
rect 13924 3108 13952 3148
rect 14001 3145 14013 3179
rect 14047 3176 14059 3179
rect 14182 3176 14188 3188
rect 14047 3148 14188 3176
rect 14047 3145 14059 3148
rect 14001 3139 14059 3145
rect 14182 3136 14188 3148
rect 14240 3136 14246 3188
rect 18325 3179 18383 3185
rect 18325 3176 18337 3179
rect 14292 3148 18337 3176
rect 14292 3108 14320 3148
rect 18325 3145 18337 3148
rect 18371 3145 18383 3179
rect 20714 3176 20720 3188
rect 18325 3139 18383 3145
rect 20364 3148 20720 3176
rect 20364 3108 20392 3148
rect 20714 3136 20720 3148
rect 20772 3136 20778 3188
rect 25222 3136 25228 3188
rect 25280 3176 25286 3188
rect 25685 3179 25743 3185
rect 25685 3176 25697 3179
rect 25280 3148 25697 3176
rect 25280 3136 25286 3148
rect 25685 3145 25697 3148
rect 25731 3176 25743 3179
rect 25774 3176 25780 3188
rect 25731 3148 25780 3176
rect 25731 3145 25743 3148
rect 25685 3139 25743 3145
rect 25774 3136 25780 3148
rect 25832 3136 25838 3188
rect 25884 3148 27384 3176
rect 13924 3080 14320 3108
rect 17972 3080 20392 3108
rect 11793 3071 11851 3077
rect 3421 3043 3479 3049
rect 3421 3009 3433 3043
rect 3467 3040 3479 3043
rect 8018 3040 8024 3052
rect 3467 3012 8024 3040
rect 3467 3009 3479 3012
rect 3421 3003 3479 3009
rect 8018 3000 8024 3012
rect 8076 3000 8082 3052
rect 9033 3043 9091 3049
rect 9033 3009 9045 3043
rect 9079 3040 9091 3043
rect 9769 3043 9827 3049
rect 9769 3040 9781 3043
rect 9079 3012 9781 3040
rect 9079 3009 9091 3012
rect 9033 3003 9091 3009
rect 9769 3009 9781 3012
rect 9815 3009 9827 3043
rect 12710 3040 12716 3052
rect 12671 3012 12716 3040
rect 9769 3003 9827 3009
rect 12710 3000 12716 3012
rect 12768 3000 12774 3052
rect 14826 3040 14832 3052
rect 14787 3012 14832 3040
rect 14826 3000 14832 3012
rect 14884 3000 14890 3052
rect 15381 3043 15439 3049
rect 15381 3009 15393 3043
rect 15427 3040 15439 3043
rect 16114 3040 16120 3052
rect 15427 3012 15976 3040
rect 16075 3012 16120 3040
rect 15427 3009 15439 3012
rect 15381 3003 15439 3009
rect 3142 2972 3148 2984
rect 3103 2944 3148 2972
rect 3142 2932 3148 2944
rect 3200 2932 3206 2984
rect 7282 2972 7288 2984
rect 7243 2944 7288 2972
rect 7282 2932 7288 2944
rect 7340 2932 7346 2984
rect 7377 2975 7435 2981
rect 7377 2941 7389 2975
rect 7423 2941 7435 2975
rect 7377 2935 7435 2941
rect 8573 2975 8631 2981
rect 8573 2941 8585 2975
rect 8619 2972 8631 2975
rect 8662 2972 8668 2984
rect 8619 2944 8668 2972
rect 8619 2941 8631 2944
rect 8573 2935 8631 2941
rect 4525 2839 4583 2845
rect 4525 2805 4537 2839
rect 4571 2836 4583 2839
rect 4614 2836 4620 2848
rect 4571 2808 4620 2836
rect 4571 2805 4583 2808
rect 4525 2799 4583 2805
rect 4614 2796 4620 2808
rect 4672 2796 4678 2848
rect 7392 2836 7420 2935
rect 8662 2932 8668 2944
rect 8720 2932 8726 2984
rect 8846 2972 8852 2984
rect 8807 2944 8852 2972
rect 8846 2932 8852 2944
rect 8904 2932 8910 2984
rect 9398 2932 9404 2984
rect 9456 2972 9462 2984
rect 9493 2975 9551 2981
rect 9493 2972 9505 2975
rect 9456 2944 9505 2972
rect 9456 2932 9462 2944
rect 9493 2941 9505 2944
rect 9539 2941 9551 2975
rect 11701 2975 11759 2981
rect 9493 2935 9551 2941
rect 9600 2944 11652 2972
rect 9600 2916 9628 2944
rect 7837 2907 7895 2913
rect 7837 2873 7849 2907
rect 7883 2904 7895 2907
rect 9214 2904 9220 2916
rect 7883 2876 9220 2904
rect 7883 2873 7895 2876
rect 7837 2867 7895 2873
rect 9214 2864 9220 2876
rect 9272 2864 9278 2916
rect 9582 2864 9588 2916
rect 9640 2864 9646 2916
rect 10873 2839 10931 2845
rect 10873 2836 10885 2839
rect 7392 2808 10885 2836
rect 10873 2805 10885 2808
rect 10919 2805 10931 2839
rect 11624 2836 11652 2944
rect 11701 2941 11713 2975
rect 11747 2972 11759 2975
rect 12342 2972 12348 2984
rect 11747 2944 12348 2972
rect 11747 2941 11759 2944
rect 11701 2935 11759 2941
rect 12342 2932 12348 2944
rect 12400 2932 12406 2984
rect 12434 2932 12440 2984
rect 12492 2972 12498 2984
rect 14182 2972 14188 2984
rect 12492 2944 14188 2972
rect 12492 2932 12498 2944
rect 14182 2932 14188 2944
rect 14240 2932 14246 2984
rect 14918 2972 14924 2984
rect 14879 2944 14924 2972
rect 14918 2932 14924 2944
rect 14976 2932 14982 2984
rect 15286 2932 15292 2984
rect 15344 2972 15350 2984
rect 15841 2975 15899 2981
rect 15841 2972 15853 2975
rect 15344 2944 15853 2972
rect 15344 2932 15350 2944
rect 15841 2941 15853 2944
rect 15887 2941 15899 2975
rect 15948 2972 15976 3012
rect 16114 3000 16120 3012
rect 16172 3000 16178 3052
rect 17972 2972 18000 3080
rect 22922 3068 22928 3120
rect 22980 3108 22986 3120
rect 22980 3080 24164 3108
rect 22980 3068 22986 3080
rect 18049 3043 18107 3049
rect 18049 3009 18061 3043
rect 18095 3040 18107 3043
rect 19797 3043 19855 3049
rect 18095 3012 18276 3040
rect 18095 3009 18107 3012
rect 18049 3003 18107 3009
rect 15948 2944 18000 2972
rect 18141 2975 18199 2981
rect 15841 2935 15899 2941
rect 18141 2941 18153 2975
rect 18187 2941 18199 2975
rect 18141 2935 18199 2941
rect 17497 2907 17555 2913
rect 17497 2873 17509 2907
rect 17543 2904 17555 2907
rect 18156 2904 18184 2935
rect 17543 2876 18184 2904
rect 17543 2873 17555 2876
rect 17497 2867 17555 2873
rect 13906 2836 13912 2848
rect 11624 2808 13912 2836
rect 10873 2799 10931 2805
rect 13906 2796 13912 2808
rect 13964 2796 13970 2848
rect 15930 2796 15936 2848
rect 15988 2836 15994 2848
rect 18248 2836 18276 3012
rect 19797 3009 19809 3043
rect 19843 3040 19855 3043
rect 21082 3040 21088 3052
rect 19843 3012 21088 3040
rect 19843 3009 19855 3012
rect 19797 3003 19855 3009
rect 21082 3000 21088 3012
rect 21140 3000 21146 3052
rect 24136 3040 24164 3080
rect 24578 3040 24584 3052
rect 24136 3012 24440 3040
rect 24539 3012 24584 3040
rect 18966 2932 18972 2984
rect 19024 2972 19030 2984
rect 19061 2975 19119 2981
rect 19061 2972 19073 2975
rect 19024 2944 19073 2972
rect 19024 2932 19030 2944
rect 19061 2941 19073 2944
rect 19107 2941 19119 2975
rect 19061 2935 19119 2941
rect 19426 2932 19432 2984
rect 19484 2972 19490 2984
rect 19521 2975 19579 2981
rect 19521 2972 19533 2975
rect 19484 2944 19533 2972
rect 19484 2932 19490 2944
rect 19521 2941 19533 2944
rect 19567 2941 19579 2975
rect 20346 2972 20352 2984
rect 20307 2944 20352 2972
rect 19521 2935 19579 2941
rect 20346 2932 20352 2944
rect 20404 2932 20410 2984
rect 20622 2972 20628 2984
rect 20583 2944 20628 2972
rect 20622 2932 20628 2944
rect 20680 2932 20686 2984
rect 22094 2932 22100 2984
rect 22152 2972 22158 2984
rect 22465 2975 22523 2981
rect 22465 2972 22477 2975
rect 22152 2944 22477 2972
rect 22152 2932 22158 2944
rect 22465 2941 22477 2944
rect 22511 2941 22523 2975
rect 22465 2935 22523 2941
rect 22112 2904 22140 2932
rect 21284 2876 22140 2904
rect 22480 2904 22508 2935
rect 22554 2932 22560 2984
rect 22612 2972 22618 2984
rect 22612 2944 22657 2972
rect 22612 2932 22618 2944
rect 23106 2932 23112 2984
rect 23164 2972 23170 2984
rect 24305 2975 24363 2981
rect 24305 2972 24317 2975
rect 23164 2944 24317 2972
rect 23164 2932 23170 2944
rect 24305 2941 24317 2944
rect 24351 2941 24363 2975
rect 24412 2972 24440 3012
rect 24578 3000 24584 3012
rect 24636 3000 24642 3052
rect 25884 2972 25912 3148
rect 27356 3108 27384 3148
rect 27430 3136 27436 3188
rect 27488 3176 27494 3188
rect 37734 3176 37740 3188
rect 27488 3148 37740 3176
rect 27488 3136 27494 3148
rect 37734 3136 37740 3148
rect 37792 3136 37798 3188
rect 29638 3108 29644 3120
rect 27356 3080 29644 3108
rect 29638 3068 29644 3080
rect 29696 3068 29702 3120
rect 32582 3068 32588 3120
rect 32640 3108 32646 3120
rect 32640 3080 35020 3108
rect 32640 3068 32646 3080
rect 26697 3043 26755 3049
rect 26697 3009 26709 3043
rect 26743 3040 26755 3043
rect 28258 3040 28264 3052
rect 26743 3012 28264 3040
rect 26743 3009 26755 3012
rect 26697 3003 26755 3009
rect 28258 3000 28264 3012
rect 28316 3000 28322 3052
rect 29270 3040 29276 3052
rect 29231 3012 29276 3040
rect 29270 3000 29276 3012
rect 29328 3000 29334 3052
rect 29822 3040 29828 3052
rect 29783 3012 29828 3040
rect 29822 3000 29828 3012
rect 29880 3000 29886 3052
rect 30190 3000 30196 3052
rect 30248 3040 30254 3052
rect 31573 3043 31631 3049
rect 31573 3040 31585 3043
rect 30248 3012 31585 3040
rect 30248 3000 30254 3012
rect 31573 3009 31585 3012
rect 31619 3040 31631 3043
rect 31619 3012 31984 3040
rect 31619 3009 31631 3012
rect 31573 3003 31631 3009
rect 24412 2944 25912 2972
rect 26421 2975 26479 2981
rect 24305 2935 24363 2941
rect 26421 2941 26433 2975
rect 26467 2972 26479 2975
rect 27614 2972 27620 2984
rect 26467 2944 27620 2972
rect 26467 2941 26479 2944
rect 26421 2935 26479 2941
rect 27614 2932 27620 2944
rect 27672 2932 27678 2984
rect 29963 2975 30021 2981
rect 29963 2972 29975 2975
rect 29196 2944 29975 2972
rect 22738 2904 22744 2916
rect 22480 2876 22744 2904
rect 21284 2836 21312 2876
rect 22738 2864 22744 2876
rect 22796 2864 22802 2916
rect 23014 2904 23020 2916
rect 22975 2876 23020 2904
rect 23014 2864 23020 2876
rect 23072 2864 23078 2916
rect 15988 2808 21312 2836
rect 21913 2839 21971 2845
rect 15988 2796 15994 2808
rect 21913 2805 21925 2839
rect 21959 2836 21971 2839
rect 23382 2836 23388 2848
rect 21959 2808 23388 2836
rect 21959 2805 21971 2808
rect 21913 2799 21971 2805
rect 23382 2796 23388 2808
rect 23440 2796 23446 2848
rect 23474 2796 23480 2848
rect 23532 2836 23538 2848
rect 27801 2839 27859 2845
rect 27801 2836 27813 2839
rect 23532 2808 27813 2836
rect 23532 2796 23538 2808
rect 27801 2805 27813 2808
rect 27847 2836 27859 2839
rect 29196 2836 29224 2944
rect 29963 2941 29975 2944
rect 30009 2941 30021 2975
rect 29963 2935 30021 2941
rect 30101 2975 30159 2981
rect 30101 2941 30113 2975
rect 30147 2941 30159 2975
rect 31846 2972 31852 2984
rect 31807 2944 31852 2972
rect 30101 2935 30159 2941
rect 29822 2864 29828 2916
rect 29880 2904 29886 2916
rect 30116 2904 30144 2935
rect 31846 2932 31852 2944
rect 31904 2932 31910 2984
rect 31956 2972 31984 3012
rect 34514 3000 34520 3052
rect 34572 3040 34578 3052
rect 34885 3043 34943 3049
rect 34885 3040 34897 3043
rect 34572 3012 34897 3040
rect 34572 3000 34578 3012
rect 34885 3009 34897 3012
rect 34931 3009 34943 3043
rect 34992 3040 35020 3080
rect 35434 3068 35440 3120
rect 35492 3108 35498 3120
rect 36725 3111 36783 3117
rect 36725 3108 36737 3111
rect 35492 3080 36737 3108
rect 35492 3068 35498 3080
rect 36725 3077 36737 3080
rect 36771 3077 36783 3111
rect 36725 3071 36783 3077
rect 37093 3043 37151 3049
rect 37093 3040 37105 3043
rect 34992 3012 37105 3040
rect 34885 3003 34943 3009
rect 37093 3009 37105 3012
rect 37139 3009 37151 3043
rect 37093 3003 37151 3009
rect 33594 2972 33600 2984
rect 31956 2944 33600 2972
rect 33594 2932 33600 2944
rect 33652 2932 33658 2984
rect 33689 2975 33747 2981
rect 33689 2941 33701 2975
rect 33735 2972 33747 2975
rect 33870 2972 33876 2984
rect 33735 2944 33876 2972
rect 33735 2941 33747 2944
rect 33689 2935 33747 2941
rect 33870 2932 33876 2944
rect 33928 2932 33934 2984
rect 34422 2932 34428 2984
rect 34480 2972 34486 2984
rect 35437 2975 35495 2981
rect 35437 2972 35449 2975
rect 34480 2944 35449 2972
rect 34480 2932 34486 2944
rect 35437 2941 35449 2944
rect 35483 2941 35495 2975
rect 35437 2935 35495 2941
rect 35713 2975 35771 2981
rect 35713 2941 35725 2975
rect 35759 2941 35771 2975
rect 35894 2972 35900 2984
rect 35855 2944 35900 2972
rect 35713 2935 35771 2941
rect 29880 2876 30144 2904
rect 29880 2864 29886 2876
rect 27847 2808 29224 2836
rect 30116 2836 30144 2876
rect 33229 2907 33287 2913
rect 33229 2873 33241 2907
rect 33275 2904 33287 2907
rect 33318 2904 33324 2916
rect 33275 2876 33324 2904
rect 33275 2873 33287 2876
rect 33229 2867 33287 2873
rect 33318 2864 33324 2876
rect 33376 2864 33382 2916
rect 35728 2904 35756 2935
rect 35894 2932 35900 2944
rect 35952 2932 35958 2984
rect 36725 2975 36783 2981
rect 36725 2941 36737 2975
rect 36771 2972 36783 2975
rect 36817 2975 36875 2981
rect 36817 2972 36829 2975
rect 36771 2944 36829 2972
rect 36771 2941 36783 2944
rect 36725 2935 36783 2941
rect 36817 2941 36829 2944
rect 36863 2941 36875 2975
rect 36817 2935 36875 2941
rect 33888 2876 35756 2904
rect 38473 2907 38531 2913
rect 33502 2836 33508 2848
rect 30116 2808 33508 2836
rect 27847 2805 27859 2808
rect 27801 2799 27859 2805
rect 33502 2796 33508 2808
rect 33560 2836 33566 2848
rect 33888 2845 33916 2876
rect 38473 2873 38485 2907
rect 38519 2904 38531 2907
rect 39022 2904 39028 2916
rect 38519 2876 39028 2904
rect 38519 2873 38531 2876
rect 38473 2867 38531 2873
rect 39022 2864 39028 2876
rect 39080 2864 39086 2916
rect 33873 2839 33931 2845
rect 33873 2836 33885 2839
rect 33560 2808 33885 2836
rect 33560 2796 33566 2808
rect 33873 2805 33885 2808
rect 33919 2805 33931 2839
rect 33873 2799 33931 2805
rect 1104 2746 39836 2768
rect 1104 2694 19606 2746
rect 19658 2694 19670 2746
rect 19722 2694 19734 2746
rect 19786 2694 19798 2746
rect 19850 2694 39836 2746
rect 1104 2672 39836 2694
rect 3418 2592 3424 2644
rect 3476 2632 3482 2644
rect 24394 2632 24400 2644
rect 3476 2604 19564 2632
rect 3476 2592 3482 2604
rect 15562 2564 15568 2576
rect 13096 2536 15568 2564
rect 3142 2456 3148 2508
rect 3200 2496 3206 2508
rect 7193 2499 7251 2505
rect 7193 2496 7205 2499
rect 3200 2468 7205 2496
rect 3200 2456 3206 2468
rect 7193 2465 7205 2468
rect 7239 2465 7251 2499
rect 7193 2459 7251 2465
rect 7469 2499 7527 2505
rect 7469 2465 7481 2499
rect 7515 2496 7527 2499
rect 7742 2496 7748 2508
rect 7515 2468 7748 2496
rect 7515 2465 7527 2468
rect 7469 2459 7527 2465
rect 7742 2456 7748 2468
rect 7800 2456 7806 2508
rect 9214 2456 9220 2508
rect 9272 2496 9278 2508
rect 10689 2499 10747 2505
rect 10689 2496 10701 2499
rect 9272 2468 10701 2496
rect 9272 2456 9278 2468
rect 10689 2465 10701 2468
rect 10735 2465 10747 2499
rect 12618 2496 12624 2508
rect 12579 2468 12624 2496
rect 10689 2459 10747 2465
rect 12618 2456 12624 2468
rect 12676 2456 12682 2508
rect 13096 2505 13124 2536
rect 15562 2524 15568 2536
rect 15620 2524 15626 2576
rect 18877 2567 18935 2573
rect 18877 2533 18889 2567
rect 18923 2564 18935 2567
rect 19242 2564 19248 2576
rect 18923 2536 19248 2564
rect 18923 2533 18935 2536
rect 18877 2527 18935 2533
rect 19242 2524 19248 2536
rect 19300 2524 19306 2576
rect 13081 2499 13139 2505
rect 13081 2465 13093 2499
rect 13127 2465 13139 2499
rect 14090 2496 14096 2508
rect 14051 2468 14096 2496
rect 13081 2459 13139 2465
rect 14090 2456 14096 2468
rect 14148 2456 14154 2508
rect 14553 2499 14611 2505
rect 14553 2465 14565 2499
rect 14599 2496 14611 2499
rect 15749 2499 15807 2505
rect 15749 2496 15761 2499
rect 14599 2468 15761 2496
rect 14599 2465 14611 2468
rect 14553 2459 14611 2465
rect 15749 2465 15761 2468
rect 15795 2465 15807 2499
rect 15749 2459 15807 2465
rect 16022 2456 16028 2508
rect 16080 2456 16086 2508
rect 9674 2388 9680 2440
rect 9732 2428 9738 2440
rect 10413 2431 10471 2437
rect 10413 2428 10425 2431
rect 9732 2400 10425 2428
rect 9732 2388 9738 2400
rect 10413 2397 10425 2400
rect 10459 2428 10471 2431
rect 12434 2428 12440 2440
rect 10459 2400 12440 2428
rect 10459 2397 10471 2400
rect 10413 2391 10471 2397
rect 12434 2388 12440 2400
rect 12492 2388 12498 2440
rect 13170 2428 13176 2440
rect 13131 2400 13176 2428
rect 13170 2388 13176 2400
rect 13228 2388 13234 2440
rect 13906 2388 13912 2440
rect 13964 2428 13970 2440
rect 14001 2431 14059 2437
rect 14001 2428 14013 2431
rect 13964 2400 14013 2428
rect 13964 2388 13970 2400
rect 14001 2397 14013 2400
rect 14047 2397 14059 2431
rect 14001 2391 14059 2397
rect 14182 2388 14188 2440
rect 14240 2428 14246 2440
rect 15473 2431 15531 2437
rect 15473 2428 15485 2431
rect 14240 2400 15485 2428
rect 14240 2388 14246 2400
rect 15473 2397 15485 2400
rect 15519 2428 15531 2431
rect 16040 2428 16068 2456
rect 15519 2400 16068 2428
rect 19429 2431 19487 2437
rect 15519 2397 15531 2400
rect 15473 2391 15531 2397
rect 19429 2397 19441 2431
rect 19475 2397 19487 2431
rect 19536 2428 19564 2604
rect 23308 2604 24400 2632
rect 22465 2567 22523 2573
rect 22465 2533 22477 2567
rect 22511 2564 22523 2567
rect 23198 2564 23204 2576
rect 22511 2536 23204 2564
rect 22511 2533 22523 2536
rect 22465 2527 22523 2533
rect 23198 2524 23204 2536
rect 23256 2524 23262 2576
rect 19702 2496 19708 2508
rect 19663 2468 19708 2496
rect 19702 2456 19708 2468
rect 19760 2496 19766 2508
rect 21177 2499 21235 2505
rect 21177 2496 21189 2499
rect 19760 2468 21189 2496
rect 19760 2456 19766 2468
rect 21177 2465 21189 2468
rect 21223 2465 21235 2499
rect 21177 2459 21235 2465
rect 21913 2499 21971 2505
rect 21913 2465 21925 2499
rect 21959 2496 21971 2499
rect 22646 2496 22652 2508
rect 21959 2468 22652 2496
rect 21959 2465 21971 2468
rect 21913 2459 21971 2465
rect 22646 2456 22652 2468
rect 22704 2456 22710 2508
rect 22738 2456 22744 2508
rect 22796 2496 22802 2508
rect 23308 2505 23336 2604
rect 24394 2592 24400 2604
rect 24452 2592 24458 2644
rect 27062 2632 27068 2644
rect 25148 2604 27068 2632
rect 23382 2524 23388 2576
rect 23440 2564 23446 2576
rect 25148 2573 25176 2604
rect 27062 2592 27068 2604
rect 27120 2592 27126 2644
rect 31588 2604 35572 2632
rect 25133 2567 25191 2573
rect 23440 2536 24164 2564
rect 23440 2524 23446 2536
rect 23293 2499 23351 2505
rect 22796 2468 23152 2496
rect 22796 2456 22802 2468
rect 19889 2431 19947 2437
rect 19889 2428 19901 2431
rect 19536 2400 19901 2428
rect 19429 2391 19487 2397
rect 19889 2397 19901 2400
rect 19935 2397 19947 2431
rect 19889 2391 19947 2397
rect 23017 2431 23075 2437
rect 23017 2397 23029 2431
rect 23063 2397 23075 2431
rect 23124 2428 23152 2468
rect 23293 2465 23305 2499
rect 23339 2465 23351 2499
rect 23474 2496 23480 2508
rect 23435 2468 23480 2496
rect 23293 2459 23351 2465
rect 23474 2456 23480 2468
rect 23532 2456 23538 2508
rect 24136 2505 24164 2536
rect 25133 2533 25145 2567
rect 25179 2533 25191 2567
rect 26234 2564 26240 2576
rect 25133 2527 25191 2533
rect 25700 2536 26240 2564
rect 25700 2505 25728 2536
rect 26234 2524 26240 2536
rect 26292 2564 26298 2576
rect 29822 2564 29828 2576
rect 26292 2536 27476 2564
rect 26292 2524 26298 2536
rect 27448 2505 27476 2536
rect 27724 2536 29828 2564
rect 27724 2505 27752 2536
rect 29822 2524 29828 2536
rect 29880 2524 29886 2576
rect 24121 2499 24179 2505
rect 24121 2465 24133 2499
rect 24167 2465 24179 2499
rect 24121 2459 24179 2465
rect 25685 2499 25743 2505
rect 25685 2465 25697 2499
rect 25731 2465 25743 2499
rect 25685 2459 25743 2465
rect 25961 2499 26019 2505
rect 25961 2465 25973 2499
rect 26007 2496 26019 2499
rect 27433 2499 27491 2505
rect 26007 2468 27384 2496
rect 26007 2465 26019 2468
rect 25961 2459 26019 2465
rect 24029 2431 24087 2437
rect 24029 2428 24041 2431
rect 23124 2400 24041 2428
rect 23017 2391 23075 2397
rect 24029 2397 24041 2400
rect 24075 2397 24087 2431
rect 24578 2428 24584 2440
rect 24539 2400 24584 2428
rect 24029 2391 24087 2397
rect 19444 2360 19472 2391
rect 21269 2363 21327 2369
rect 21269 2360 21281 2363
rect 19444 2332 21281 2360
rect 21269 2329 21281 2332
rect 21315 2329 21327 2363
rect 23032 2360 23060 2391
rect 24578 2388 24584 2400
rect 24636 2388 24642 2440
rect 25774 2388 25780 2440
rect 25832 2428 25838 2440
rect 26145 2431 26203 2437
rect 26145 2428 26157 2431
rect 25832 2400 26157 2428
rect 25832 2388 25838 2400
rect 26145 2397 26157 2400
rect 26191 2397 26203 2431
rect 26145 2391 26203 2397
rect 26881 2431 26939 2437
rect 26881 2397 26893 2431
rect 26927 2397 26939 2431
rect 27356 2428 27384 2468
rect 27433 2465 27445 2499
rect 27479 2465 27491 2499
rect 27433 2459 27491 2465
rect 27709 2499 27767 2505
rect 27709 2465 27721 2499
rect 27755 2465 27767 2499
rect 27890 2496 27896 2508
rect 27851 2468 27896 2496
rect 27709 2459 27767 2465
rect 27724 2428 27752 2459
rect 27890 2456 27896 2468
rect 27948 2456 27954 2508
rect 28353 2499 28411 2505
rect 28353 2465 28365 2499
rect 28399 2496 28411 2499
rect 28902 2496 28908 2508
rect 28399 2468 28908 2496
rect 28399 2465 28411 2468
rect 28353 2459 28411 2465
rect 28902 2456 28908 2468
rect 28960 2456 28966 2508
rect 29638 2456 29644 2508
rect 29696 2496 29702 2508
rect 29733 2499 29791 2505
rect 29733 2496 29745 2499
rect 29696 2468 29745 2496
rect 29696 2456 29702 2468
rect 29733 2465 29745 2468
rect 29779 2465 29791 2499
rect 30006 2496 30012 2508
rect 29919 2468 30012 2496
rect 29733 2459 29791 2465
rect 27356 2400 27752 2428
rect 29748 2428 29776 2459
rect 30006 2456 30012 2468
rect 30064 2496 30070 2508
rect 31481 2499 31539 2505
rect 31481 2496 31493 2499
rect 30064 2468 31493 2496
rect 30064 2456 30070 2468
rect 31481 2465 31493 2468
rect 31527 2465 31539 2499
rect 31481 2459 31539 2465
rect 30190 2428 30196 2440
rect 29748 2400 30196 2428
rect 26881 2391 26939 2397
rect 26896 2360 26924 2391
rect 30190 2388 30196 2400
rect 30248 2388 30254 2440
rect 31588 2360 31616 2604
rect 32585 2567 32643 2573
rect 32585 2533 32597 2567
rect 32631 2564 32643 2567
rect 33226 2564 33232 2576
rect 32631 2536 33232 2564
rect 32631 2533 32643 2536
rect 32585 2527 32643 2533
rect 33226 2524 33232 2536
rect 33284 2524 33290 2576
rect 33502 2505 33508 2508
rect 33459 2499 33508 2505
rect 33459 2465 33471 2499
rect 33505 2465 33508 2499
rect 33459 2459 33508 2465
rect 33502 2456 33508 2459
rect 33560 2456 33566 2508
rect 35434 2496 35440 2508
rect 35395 2468 35440 2496
rect 35434 2456 35440 2468
rect 35492 2456 35498 2508
rect 35544 2496 35572 2604
rect 35713 2499 35771 2505
rect 35713 2496 35725 2499
rect 35544 2468 35725 2496
rect 35713 2465 35725 2468
rect 35759 2465 35771 2499
rect 35713 2459 35771 2465
rect 33134 2428 33140 2440
rect 33095 2400 33140 2428
rect 33134 2388 33140 2400
rect 33192 2388 33198 2440
rect 33597 2431 33655 2437
rect 33597 2397 33609 2431
rect 33643 2397 33655 2431
rect 33597 2391 33655 2397
rect 23032 2332 26924 2360
rect 26988 2332 28672 2360
rect 21269 2323 21327 2329
rect 2406 2252 2412 2304
rect 2464 2292 2470 2304
rect 8573 2295 8631 2301
rect 8573 2292 8585 2295
rect 2464 2264 8585 2292
rect 2464 2252 2470 2264
rect 8573 2261 8585 2264
rect 8619 2261 8631 2295
rect 11974 2292 11980 2304
rect 11935 2264 11980 2292
rect 8573 2255 8631 2261
rect 11974 2252 11980 2264
rect 12032 2252 12038 2304
rect 15838 2252 15844 2304
rect 15896 2292 15902 2304
rect 16853 2295 16911 2301
rect 16853 2292 16865 2295
rect 15896 2264 16865 2292
rect 15896 2252 15902 2264
rect 16853 2261 16865 2264
rect 16899 2261 16911 2295
rect 16853 2255 16911 2261
rect 23014 2252 23020 2304
rect 23072 2292 23078 2304
rect 26988 2292 27016 2332
rect 23072 2264 27016 2292
rect 23072 2252 23078 2264
rect 27430 2252 27436 2304
rect 27488 2292 27494 2304
rect 28537 2295 28595 2301
rect 28537 2292 28549 2295
rect 27488 2264 28549 2292
rect 27488 2252 27494 2264
rect 28537 2261 28549 2264
rect 28583 2261 28595 2295
rect 28644 2292 28672 2332
rect 30668 2332 31616 2360
rect 30668 2292 30696 2332
rect 31662 2320 31668 2372
rect 31720 2360 31726 2372
rect 33612 2360 33640 2391
rect 31720 2332 33640 2360
rect 31720 2320 31726 2332
rect 31294 2292 31300 2304
rect 28644 2264 30696 2292
rect 31255 2264 31300 2292
rect 28537 2255 28595 2261
rect 31294 2252 31300 2264
rect 31352 2252 31358 2304
rect 33134 2252 33140 2304
rect 33192 2292 33198 2304
rect 34422 2292 34428 2304
rect 33192 2264 34428 2292
rect 33192 2252 33198 2264
rect 34422 2252 34428 2264
rect 34480 2252 34486 2304
rect 37001 2295 37059 2301
rect 37001 2261 37013 2295
rect 37047 2292 37059 2295
rect 37182 2292 37188 2304
rect 37047 2264 37188 2292
rect 37047 2261 37059 2264
rect 37001 2255 37059 2261
rect 37182 2252 37188 2264
rect 37240 2252 37246 2304
rect 1104 2202 39836 2224
rect 1104 2150 4246 2202
rect 4298 2150 4310 2202
rect 4362 2150 4374 2202
rect 4426 2150 4438 2202
rect 4490 2150 34966 2202
rect 35018 2150 35030 2202
rect 35082 2150 35094 2202
rect 35146 2150 35158 2202
rect 35210 2150 39836 2202
rect 1104 2128 39836 2150
rect 24578 2048 24584 2100
rect 24636 2088 24642 2100
rect 31846 2088 31852 2100
rect 24636 2060 31852 2088
rect 24636 2048 24642 2060
rect 31846 2048 31852 2060
rect 31904 2048 31910 2100
rect 29730 1096 29736 1148
rect 29788 1136 29794 1148
rect 35158 1136 35164 1148
rect 29788 1108 35164 1136
rect 29788 1096 29794 1108
rect 35158 1096 35164 1108
rect 35216 1096 35222 1148
<< via1 >>
rect 19606 38598 19658 38650
rect 19670 38598 19722 38650
rect 19734 38598 19786 38650
rect 19798 38598 19850 38650
rect 10508 38496 10560 38548
rect 14372 38496 14424 38548
rect 17316 38496 17368 38548
rect 6000 38428 6052 38480
rect 8300 38403 8352 38412
rect 8300 38369 8309 38403
rect 8309 38369 8343 38403
rect 8343 38369 8352 38403
rect 8300 38360 8352 38369
rect 8668 38428 8720 38480
rect 9588 38428 9640 38480
rect 16580 38428 16632 38480
rect 12900 38360 12952 38412
rect 14188 38403 14240 38412
rect 14188 38369 14197 38403
rect 14197 38369 14231 38403
rect 14231 38369 14240 38403
rect 14188 38360 14240 38369
rect 14740 38403 14792 38412
rect 14740 38369 14749 38403
rect 14749 38369 14783 38403
rect 14783 38369 14792 38403
rect 14740 38360 14792 38369
rect 8668 38292 8720 38344
rect 9312 38292 9364 38344
rect 10876 38292 10928 38344
rect 20996 38360 21048 38412
rect 21548 38360 21600 38412
rect 26240 38428 26292 38480
rect 22284 38360 22336 38412
rect 35900 38496 35952 38548
rect 29920 38360 29972 38412
rect 20720 38292 20772 38344
rect 24952 38335 25004 38344
rect 14096 38224 14148 38276
rect 21824 38224 21876 38276
rect 12716 38156 12768 38208
rect 15568 38199 15620 38208
rect 15568 38165 15577 38199
rect 15577 38165 15611 38199
rect 15611 38165 15620 38199
rect 15568 38156 15620 38165
rect 20536 38156 20588 38208
rect 21640 38156 21692 38208
rect 24952 38301 24961 38335
rect 24961 38301 24995 38335
rect 24995 38301 25004 38335
rect 24952 38292 25004 38301
rect 27436 38292 27488 38344
rect 28632 38292 28684 38344
rect 24860 38156 24912 38208
rect 26424 38156 26476 38208
rect 27620 38156 27672 38208
rect 30012 38199 30064 38208
rect 30012 38165 30021 38199
rect 30021 38165 30055 38199
rect 30055 38165 30064 38199
rect 30012 38156 30064 38165
rect 31024 38199 31076 38208
rect 31024 38165 31033 38199
rect 31033 38165 31067 38199
rect 31067 38165 31076 38199
rect 31024 38156 31076 38165
rect 4246 38054 4298 38106
rect 4310 38054 4362 38106
rect 4374 38054 4426 38106
rect 4438 38054 4490 38106
rect 34966 38054 35018 38106
rect 35030 38054 35082 38106
rect 35094 38054 35146 38106
rect 35158 38054 35210 38106
rect 4620 37952 4672 38004
rect 10876 37995 10928 38004
rect 10876 37961 10885 37995
rect 10885 37961 10919 37995
rect 10919 37961 10928 37995
rect 10876 37952 10928 37961
rect 9680 37884 9732 37936
rect 12348 37884 12400 37936
rect 3608 37859 3660 37868
rect 3608 37825 3617 37859
rect 3617 37825 3651 37859
rect 3651 37825 3660 37859
rect 3608 37816 3660 37825
rect 5632 37816 5684 37868
rect 6644 37816 6696 37868
rect 12440 37859 12492 37868
rect 12440 37825 12449 37859
rect 12449 37825 12483 37859
rect 12483 37825 12492 37859
rect 12440 37816 12492 37825
rect 12716 37859 12768 37868
rect 12716 37825 12725 37859
rect 12725 37825 12759 37859
rect 12759 37825 12768 37859
rect 12716 37816 12768 37825
rect 16212 37952 16264 38004
rect 17224 37952 17276 38004
rect 22100 37952 22152 38004
rect 16212 37816 16264 37868
rect 22468 37816 22520 37868
rect 24308 37952 24360 38004
rect 27804 37952 27856 38004
rect 31668 37952 31720 38004
rect 39396 37952 39448 38004
rect 3976 37748 4028 37800
rect 8392 37748 8444 37800
rect 9220 37748 9272 37800
rect 10600 37791 10652 37800
rect 10600 37757 10609 37791
rect 10609 37757 10643 37791
rect 10643 37757 10652 37791
rect 10600 37748 10652 37757
rect 11060 37748 11112 37800
rect 13820 37748 13872 37800
rect 15016 37748 15068 37800
rect 15752 37791 15804 37800
rect 15752 37757 15761 37791
rect 15761 37757 15795 37791
rect 15795 37757 15804 37791
rect 15752 37748 15804 37757
rect 18512 37748 18564 37800
rect 18696 37791 18748 37800
rect 18696 37757 18705 37791
rect 18705 37757 18739 37791
rect 18739 37757 18748 37791
rect 18696 37748 18748 37757
rect 19156 37791 19208 37800
rect 19156 37757 19165 37791
rect 19165 37757 19199 37791
rect 19199 37757 19208 37791
rect 19156 37748 19208 37757
rect 19432 37791 19484 37800
rect 19432 37757 19441 37791
rect 19441 37757 19475 37791
rect 19475 37757 19484 37791
rect 19432 37748 19484 37757
rect 20536 37791 20588 37800
rect 20536 37757 20545 37791
rect 20545 37757 20579 37791
rect 20579 37757 20588 37791
rect 20536 37748 20588 37757
rect 22652 37791 22704 37800
rect 22652 37757 22661 37791
rect 22661 37757 22695 37791
rect 22695 37757 22704 37791
rect 22652 37748 22704 37757
rect 19340 37680 19392 37732
rect 21732 37680 21784 37732
rect 26424 37859 26476 37868
rect 23388 37748 23440 37800
rect 24860 37748 24912 37800
rect 25780 37748 25832 37800
rect 26424 37825 26433 37859
rect 26433 37825 26467 37859
rect 26467 37825 26476 37859
rect 26424 37816 26476 37825
rect 29000 37816 29052 37868
rect 23756 37680 23808 37732
rect 28080 37748 28132 37800
rect 30104 37748 30156 37800
rect 32036 37748 32088 37800
rect 32772 37748 32824 37800
rect 14924 37612 14976 37664
rect 18880 37612 18932 37664
rect 21180 37612 21232 37664
rect 22468 37612 22520 37664
rect 23388 37612 23440 37664
rect 23480 37612 23532 37664
rect 27528 37655 27580 37664
rect 27528 37621 27537 37655
rect 27537 37621 27571 37655
rect 27571 37621 27580 37655
rect 27528 37612 27580 37621
rect 29828 37655 29880 37664
rect 29828 37621 29837 37655
rect 29837 37621 29871 37655
rect 29871 37621 29880 37655
rect 29828 37612 29880 37621
rect 32128 37612 32180 37664
rect 38292 37612 38344 37664
rect 19606 37510 19658 37562
rect 19670 37510 19722 37562
rect 19734 37510 19786 37562
rect 19798 37510 19850 37562
rect 7656 37408 7708 37460
rect 8300 37408 8352 37460
rect 8116 37315 8168 37324
rect 8116 37281 8125 37315
rect 8125 37281 8159 37315
rect 8159 37281 8168 37315
rect 8116 37272 8168 37281
rect 10140 37340 10192 37392
rect 17224 37408 17276 37460
rect 18788 37451 18840 37460
rect 18788 37417 18797 37451
rect 18797 37417 18831 37451
rect 18831 37417 18840 37451
rect 18788 37408 18840 37417
rect 20996 37451 21048 37460
rect 20996 37417 21005 37451
rect 21005 37417 21039 37451
rect 21039 37417 21048 37451
rect 20996 37408 21048 37417
rect 21732 37451 21784 37460
rect 21732 37417 21741 37451
rect 21741 37417 21775 37451
rect 21775 37417 21784 37451
rect 21732 37408 21784 37417
rect 21824 37408 21876 37460
rect 29828 37408 29880 37460
rect 30104 37408 30156 37460
rect 33692 37451 33744 37460
rect 33692 37417 33701 37451
rect 33701 37417 33735 37451
rect 33735 37417 33744 37451
rect 33692 37408 33744 37417
rect 35532 37408 35584 37460
rect 12808 37340 12860 37392
rect 12992 37340 13044 37392
rect 8668 37315 8720 37324
rect 8668 37281 8677 37315
rect 8677 37281 8711 37315
rect 8711 37281 8720 37315
rect 8668 37272 8720 37281
rect 9680 37315 9732 37324
rect 9680 37281 9689 37315
rect 9689 37281 9723 37315
rect 9723 37281 9732 37315
rect 9680 37272 9732 37281
rect 10692 37272 10744 37324
rect 13084 37272 13136 37324
rect 13820 37315 13872 37324
rect 13820 37281 13829 37315
rect 13829 37281 13863 37315
rect 13863 37281 13872 37315
rect 13820 37272 13872 37281
rect 5632 37247 5684 37256
rect 5632 37213 5641 37247
rect 5641 37213 5675 37247
rect 5675 37213 5684 37247
rect 5632 37204 5684 37213
rect 8392 37247 8444 37256
rect 8392 37213 8401 37247
rect 8401 37213 8435 37247
rect 8435 37213 8444 37247
rect 8392 37204 8444 37213
rect 12440 37204 12492 37256
rect 14188 37247 14240 37256
rect 14188 37213 14197 37247
rect 14197 37213 14231 37247
rect 14231 37213 14240 37247
rect 14188 37204 14240 37213
rect 4804 37068 4856 37120
rect 9588 37136 9640 37188
rect 18236 37340 18288 37392
rect 19340 37340 19392 37392
rect 22284 37383 22336 37392
rect 15844 37272 15896 37324
rect 16488 37315 16540 37324
rect 16212 37247 16264 37256
rect 16212 37213 16221 37247
rect 16221 37213 16255 37247
rect 16255 37213 16264 37247
rect 16212 37204 16264 37213
rect 16488 37281 16497 37315
rect 16497 37281 16531 37315
rect 16531 37281 16540 37315
rect 16488 37272 16540 37281
rect 18512 37315 18564 37324
rect 18512 37281 18521 37315
rect 18521 37281 18555 37315
rect 18555 37281 18564 37315
rect 18512 37272 18564 37281
rect 22284 37349 22293 37383
rect 22293 37349 22327 37383
rect 22327 37349 22336 37383
rect 22284 37340 22336 37349
rect 19892 37315 19944 37324
rect 18696 37204 18748 37256
rect 19892 37281 19901 37315
rect 19901 37281 19935 37315
rect 19935 37281 19944 37315
rect 19892 37272 19944 37281
rect 20904 37315 20956 37324
rect 20904 37281 20913 37315
rect 20913 37281 20947 37315
rect 20947 37281 20956 37315
rect 20904 37272 20956 37281
rect 21640 37315 21692 37324
rect 21640 37281 21649 37315
rect 21649 37281 21683 37315
rect 21683 37281 21692 37315
rect 21640 37272 21692 37281
rect 19432 37204 19484 37256
rect 21916 37204 21968 37256
rect 22928 37315 22980 37324
rect 22928 37281 22937 37315
rect 22937 37281 22971 37315
rect 22971 37281 22980 37315
rect 23204 37315 23256 37324
rect 22928 37272 22980 37281
rect 23204 37281 23213 37315
rect 23213 37281 23247 37315
rect 23247 37281 23256 37315
rect 23204 37272 23256 37281
rect 23388 37315 23440 37324
rect 23388 37281 23397 37315
rect 23397 37281 23431 37315
rect 23431 37281 23440 37315
rect 23388 37272 23440 37281
rect 23572 37315 23624 37324
rect 23572 37281 23581 37315
rect 23581 37281 23615 37315
rect 23615 37281 23624 37315
rect 23572 37272 23624 37281
rect 23756 37272 23808 37324
rect 6000 37068 6052 37120
rect 7196 37111 7248 37120
rect 7196 37077 7205 37111
rect 7205 37077 7239 37111
rect 7239 37077 7248 37111
rect 7196 37068 7248 37077
rect 13176 37068 13228 37120
rect 15108 37136 15160 37188
rect 17316 37136 17368 37188
rect 22652 37136 22704 37188
rect 23480 37204 23532 37256
rect 24860 37272 24912 37324
rect 26608 37272 26660 37324
rect 27620 37315 27672 37324
rect 27620 37281 27629 37315
rect 27629 37281 27663 37315
rect 27663 37281 27672 37315
rect 27620 37272 27672 37281
rect 25780 37204 25832 37256
rect 29276 37272 29328 37324
rect 31024 37272 31076 37324
rect 31944 37272 31996 37324
rect 32128 37315 32180 37324
rect 32128 37281 32137 37315
rect 32137 37281 32171 37315
rect 32171 37281 32180 37315
rect 32128 37272 32180 37281
rect 35532 37272 35584 37324
rect 31852 37204 31904 37256
rect 23204 37136 23256 37188
rect 27988 37068 28040 37120
rect 28724 37111 28776 37120
rect 28724 37077 28733 37111
rect 28733 37077 28767 37111
rect 28767 37077 28776 37111
rect 28724 37068 28776 37077
rect 4246 36966 4298 37018
rect 4310 36966 4362 37018
rect 4374 36966 4426 37018
rect 4438 36966 4490 37018
rect 34966 36966 35018 37018
rect 35030 36966 35082 37018
rect 35094 36966 35146 37018
rect 35158 36966 35210 37018
rect 2780 36907 2832 36916
rect 2780 36873 2789 36907
rect 2789 36873 2823 36907
rect 2823 36873 2832 36907
rect 2780 36864 2832 36873
rect 2964 36864 3016 36916
rect 11152 36864 11204 36916
rect 3608 36728 3660 36780
rect 4804 36771 4856 36780
rect 4804 36737 4813 36771
rect 4813 36737 4847 36771
rect 4847 36737 4856 36771
rect 4804 36728 4856 36737
rect 1952 36660 2004 36712
rect 5356 36703 5408 36712
rect 5356 36669 5365 36703
rect 5365 36669 5399 36703
rect 5399 36669 5408 36703
rect 5356 36660 5408 36669
rect 6460 36728 6512 36780
rect 6920 36660 6972 36712
rect 9680 36796 9732 36848
rect 7288 36728 7340 36780
rect 8116 36771 8168 36780
rect 7196 36660 7248 36712
rect 7840 36703 7892 36712
rect 7840 36669 7849 36703
rect 7849 36669 7883 36703
rect 7883 36669 7892 36703
rect 7840 36660 7892 36669
rect 8116 36737 8125 36771
rect 8125 36737 8159 36771
rect 8159 36737 8168 36771
rect 8116 36728 8168 36737
rect 8576 36592 8628 36644
rect 7380 36524 7432 36576
rect 9956 36524 10008 36576
rect 10324 36660 10376 36712
rect 11428 36703 11480 36712
rect 11428 36669 11437 36703
rect 11437 36669 11471 36703
rect 11471 36669 11480 36703
rect 11428 36660 11480 36669
rect 12900 36771 12952 36780
rect 12900 36737 12909 36771
rect 12909 36737 12943 36771
rect 12943 36737 12952 36771
rect 16212 36864 16264 36916
rect 18788 36864 18840 36916
rect 21548 36907 21600 36916
rect 16304 36796 16356 36848
rect 19892 36796 19944 36848
rect 21272 36796 21324 36848
rect 21548 36873 21557 36907
rect 21557 36873 21591 36907
rect 21591 36873 21600 36907
rect 21548 36864 21600 36873
rect 24952 36864 25004 36916
rect 27804 36864 27856 36916
rect 32772 36907 32824 36916
rect 32772 36873 32781 36907
rect 32781 36873 32815 36907
rect 32815 36873 32824 36907
rect 32772 36864 32824 36873
rect 12900 36728 12952 36737
rect 15568 36728 15620 36780
rect 16212 36728 16264 36780
rect 18236 36728 18288 36780
rect 18420 36728 18472 36780
rect 12808 36703 12860 36712
rect 12808 36669 12817 36703
rect 12817 36669 12851 36703
rect 12851 36669 12860 36703
rect 12808 36660 12860 36669
rect 13176 36703 13228 36712
rect 13176 36669 13185 36703
rect 13185 36669 13219 36703
rect 13219 36669 13228 36703
rect 13176 36660 13228 36669
rect 15016 36660 15068 36712
rect 12992 36592 13044 36644
rect 19800 36660 19852 36712
rect 21180 36660 21232 36712
rect 21916 36703 21968 36712
rect 12164 36524 12216 36576
rect 12808 36524 12860 36576
rect 14924 36524 14976 36576
rect 15016 36524 15068 36576
rect 20076 36592 20128 36644
rect 21916 36669 21925 36703
rect 21925 36669 21959 36703
rect 21959 36669 21968 36703
rect 21916 36660 21968 36669
rect 23940 36728 23992 36780
rect 25780 36771 25832 36780
rect 23480 36660 23532 36712
rect 24124 36660 24176 36712
rect 24308 36703 24360 36712
rect 24308 36669 24317 36703
rect 24317 36669 24351 36703
rect 24351 36669 24360 36703
rect 24308 36660 24360 36669
rect 25780 36737 25789 36771
rect 25789 36737 25823 36771
rect 25823 36737 25832 36771
rect 25780 36728 25832 36737
rect 29276 36771 29328 36780
rect 29276 36737 29285 36771
rect 29285 36737 29319 36771
rect 29319 36737 29328 36771
rect 29276 36728 29328 36737
rect 30012 36728 30064 36780
rect 26056 36703 26108 36712
rect 26056 36669 26065 36703
rect 26065 36669 26099 36703
rect 26099 36669 26108 36703
rect 26056 36660 26108 36669
rect 28172 36703 28224 36712
rect 28172 36669 28181 36703
rect 28181 36669 28215 36703
rect 28215 36669 28224 36703
rect 28172 36660 28224 36669
rect 29000 36660 29052 36712
rect 32496 36703 32548 36712
rect 18144 36524 18196 36576
rect 20260 36524 20312 36576
rect 20444 36567 20496 36576
rect 20444 36533 20453 36567
rect 20453 36533 20487 36567
rect 20487 36533 20496 36567
rect 20444 36524 20496 36533
rect 23572 36592 23624 36644
rect 27436 36592 27488 36644
rect 32496 36669 32505 36703
rect 32505 36669 32539 36703
rect 32539 36669 32548 36703
rect 32496 36660 32548 36669
rect 37556 36660 37608 36712
rect 25136 36524 25188 36576
rect 26424 36524 26476 36576
rect 30656 36567 30708 36576
rect 30656 36533 30665 36567
rect 30665 36533 30699 36567
rect 30699 36533 30708 36567
rect 30656 36524 30708 36533
rect 19606 36422 19658 36474
rect 19670 36422 19722 36474
rect 19734 36422 19786 36474
rect 19798 36422 19850 36474
rect 7196 36320 7248 36372
rect 8576 36363 8628 36372
rect 8576 36329 8585 36363
rect 8585 36329 8619 36363
rect 8619 36329 8628 36363
rect 8576 36320 8628 36329
rect 11060 36363 11112 36372
rect 11060 36329 11069 36363
rect 11069 36329 11103 36363
rect 11103 36329 11112 36363
rect 11060 36320 11112 36329
rect 11152 36320 11204 36372
rect 5356 36252 5408 36304
rect 4804 36227 4856 36236
rect 4804 36193 4813 36227
rect 4813 36193 4847 36227
rect 4847 36193 4856 36227
rect 4804 36184 4856 36193
rect 7656 36252 7708 36304
rect 9680 36252 9732 36304
rect 14740 36252 14792 36304
rect 14924 36252 14976 36304
rect 17040 36252 17092 36304
rect 18512 36252 18564 36304
rect 6644 36227 6696 36236
rect 4712 36116 4764 36168
rect 5080 36159 5132 36168
rect 5080 36125 5089 36159
rect 5089 36125 5123 36159
rect 5123 36125 5132 36159
rect 5080 36116 5132 36125
rect 4620 36048 4672 36100
rect 6000 36091 6052 36100
rect 6000 36057 6009 36091
rect 6009 36057 6043 36091
rect 6043 36057 6052 36091
rect 6000 36048 6052 36057
rect 20 35980 72 36032
rect 756 35980 808 36032
rect 6644 36193 6653 36227
rect 6653 36193 6687 36227
rect 6687 36193 6696 36227
rect 6644 36184 6696 36193
rect 7380 36227 7432 36236
rect 7380 36193 7389 36227
rect 7389 36193 7423 36227
rect 7423 36193 7432 36227
rect 7380 36184 7432 36193
rect 9956 36227 10008 36236
rect 6460 36116 6512 36168
rect 6736 36048 6788 36100
rect 9956 36193 9965 36227
rect 9965 36193 9999 36227
rect 9999 36193 10008 36227
rect 9956 36184 10008 36193
rect 11428 36184 11480 36236
rect 12808 36227 12860 36236
rect 12808 36193 12817 36227
rect 12817 36193 12851 36227
rect 12851 36193 12860 36227
rect 12808 36184 12860 36193
rect 12992 36227 13044 36236
rect 12992 36193 13001 36227
rect 13001 36193 13035 36227
rect 13035 36193 13044 36227
rect 12992 36184 13044 36193
rect 9312 36116 9364 36168
rect 13084 36159 13136 36168
rect 13084 36125 13093 36159
rect 13093 36125 13127 36159
rect 13127 36125 13136 36159
rect 13084 36116 13136 36125
rect 15108 36184 15160 36236
rect 16304 36184 16356 36236
rect 16580 36227 16632 36236
rect 15016 36116 15068 36168
rect 16580 36193 16589 36227
rect 16589 36193 16623 36227
rect 16623 36193 16632 36227
rect 16580 36184 16632 36193
rect 16856 36227 16908 36236
rect 16856 36193 16865 36227
rect 16865 36193 16899 36227
rect 16899 36193 16908 36227
rect 16856 36184 16908 36193
rect 18144 36227 18196 36236
rect 18144 36193 18153 36227
rect 18153 36193 18187 36227
rect 18187 36193 18196 36227
rect 18144 36184 18196 36193
rect 19432 36252 19484 36304
rect 20444 36252 20496 36304
rect 19156 36184 19208 36236
rect 19340 36184 19392 36236
rect 16672 36116 16724 36168
rect 17316 36159 17368 36168
rect 17316 36125 17325 36159
rect 17325 36125 17359 36159
rect 17359 36125 17368 36159
rect 17316 36116 17368 36125
rect 18696 36116 18748 36168
rect 20536 36184 20588 36236
rect 20904 36184 20956 36236
rect 21272 36227 21324 36236
rect 21272 36193 21281 36227
rect 21281 36193 21315 36227
rect 21315 36193 21324 36227
rect 21272 36184 21324 36193
rect 26056 36252 26108 36304
rect 20628 36116 20680 36168
rect 22836 36227 22888 36236
rect 22836 36193 22845 36227
rect 22845 36193 22879 36227
rect 22879 36193 22888 36227
rect 22836 36184 22888 36193
rect 26608 36227 26660 36236
rect 26608 36193 26617 36227
rect 26617 36193 26651 36227
rect 26651 36193 26660 36227
rect 26608 36184 26660 36193
rect 27804 36227 27856 36236
rect 23756 36159 23808 36168
rect 6920 35980 6972 36032
rect 7196 35980 7248 36032
rect 7932 36023 7984 36032
rect 7932 35989 7941 36023
rect 7941 35989 7975 36023
rect 7975 35989 7984 36023
rect 7932 35980 7984 35989
rect 9680 35980 9732 36032
rect 14924 35980 14976 36032
rect 19156 36048 19208 36100
rect 20720 36048 20772 36100
rect 23756 36125 23765 36159
rect 23765 36125 23799 36159
rect 23799 36125 23808 36159
rect 23756 36116 23808 36125
rect 25412 36116 25464 36168
rect 27804 36193 27813 36227
rect 27813 36193 27847 36227
rect 27847 36193 27856 36227
rect 27804 36184 27856 36193
rect 31208 36320 31260 36372
rect 34520 36252 34572 36304
rect 32496 36184 32548 36236
rect 27252 36048 27304 36100
rect 28172 36116 28224 36168
rect 32312 36116 32364 36168
rect 33140 36184 33192 36236
rect 33968 36227 34020 36236
rect 33968 36193 33977 36227
rect 33977 36193 34011 36227
rect 34011 36193 34020 36227
rect 33968 36184 34020 36193
rect 35900 36184 35952 36236
rect 31208 36048 31260 36100
rect 22560 36023 22612 36032
rect 22560 35989 22569 36023
rect 22569 35989 22603 36023
rect 22603 35989 22612 36023
rect 22560 35980 22612 35989
rect 25872 35980 25924 36032
rect 27804 35980 27856 36032
rect 34152 36023 34204 36032
rect 34152 35989 34161 36023
rect 34161 35989 34195 36023
rect 34195 35989 34204 36023
rect 34152 35980 34204 35989
rect 35256 36023 35308 36032
rect 35256 35989 35265 36023
rect 35265 35989 35299 36023
rect 35299 35989 35308 36023
rect 35256 35980 35308 35989
rect 4246 35878 4298 35930
rect 4310 35878 4362 35930
rect 4374 35878 4426 35930
rect 4438 35878 4490 35930
rect 34966 35878 35018 35930
rect 35030 35878 35082 35930
rect 35094 35878 35146 35930
rect 35158 35878 35210 35930
rect 7380 35776 7432 35828
rect 8024 35776 8076 35828
rect 16672 35819 16724 35828
rect 16672 35785 16681 35819
rect 16681 35785 16715 35819
rect 16715 35785 16724 35819
rect 16672 35776 16724 35785
rect 23388 35776 23440 35828
rect 25780 35776 25832 35828
rect 26332 35776 26384 35828
rect 27252 35819 27304 35828
rect 27252 35785 27261 35819
rect 27261 35785 27295 35819
rect 27295 35785 27304 35819
rect 27252 35776 27304 35785
rect 33968 35776 34020 35828
rect 4712 35751 4764 35760
rect 4712 35717 4721 35751
rect 4721 35717 4755 35751
rect 4755 35717 4764 35751
rect 4712 35708 4764 35717
rect 4804 35640 4856 35692
rect 6644 35640 6696 35692
rect 9312 35640 9364 35692
rect 12164 35708 12216 35760
rect 5080 35504 5132 35556
rect 6092 35615 6144 35624
rect 6092 35581 6101 35615
rect 6101 35581 6135 35615
rect 6135 35581 6144 35615
rect 6092 35572 6144 35581
rect 6736 35572 6788 35624
rect 10416 35572 10468 35624
rect 15108 35640 15160 35692
rect 16856 35640 16908 35692
rect 11152 35615 11204 35624
rect 11152 35581 11161 35615
rect 11161 35581 11195 35615
rect 11195 35581 11204 35615
rect 11152 35572 11204 35581
rect 13268 35615 13320 35624
rect 13268 35581 13277 35615
rect 13277 35581 13311 35615
rect 13311 35581 13320 35615
rect 13268 35572 13320 35581
rect 13636 35572 13688 35624
rect 14924 35615 14976 35624
rect 14924 35581 14933 35615
rect 14933 35581 14967 35615
rect 14967 35581 14976 35615
rect 14924 35572 14976 35581
rect 15568 35615 15620 35624
rect 15568 35581 15577 35615
rect 15577 35581 15611 35615
rect 15611 35581 15620 35615
rect 15568 35572 15620 35581
rect 15844 35615 15896 35624
rect 15844 35581 15853 35615
rect 15853 35581 15887 35615
rect 15887 35581 15896 35615
rect 15844 35572 15896 35581
rect 16764 35615 16816 35624
rect 16764 35581 16773 35615
rect 16773 35581 16807 35615
rect 16807 35581 16816 35615
rect 16764 35572 16816 35581
rect 16948 35572 17000 35624
rect 6184 35504 6236 35556
rect 7932 35504 7984 35556
rect 20260 35708 20312 35760
rect 21364 35708 21416 35760
rect 21824 35708 21876 35760
rect 18788 35683 18840 35692
rect 18788 35649 18797 35683
rect 18797 35649 18831 35683
rect 18831 35649 18840 35683
rect 18788 35640 18840 35649
rect 18328 35572 18380 35624
rect 18880 35615 18932 35624
rect 18880 35581 18889 35615
rect 18889 35581 18923 35615
rect 18923 35581 18932 35615
rect 18880 35572 18932 35581
rect 19340 35572 19392 35624
rect 20628 35640 20680 35692
rect 21916 35640 21968 35692
rect 19892 35504 19944 35556
rect 21640 35615 21692 35624
rect 21640 35581 21649 35615
rect 21649 35581 21683 35615
rect 21683 35581 21692 35615
rect 21824 35615 21876 35624
rect 21640 35572 21692 35581
rect 21824 35581 21833 35615
rect 21833 35581 21867 35615
rect 21867 35581 21876 35615
rect 21824 35572 21876 35581
rect 22008 35615 22060 35624
rect 22008 35581 22017 35615
rect 22017 35581 22051 35615
rect 22051 35581 22060 35615
rect 22008 35572 22060 35581
rect 22652 35572 22704 35624
rect 26240 35708 26292 35760
rect 33140 35708 33192 35760
rect 29368 35640 29420 35692
rect 32036 35683 32088 35692
rect 32036 35649 32045 35683
rect 32045 35649 32079 35683
rect 32079 35649 32088 35683
rect 32312 35683 32364 35692
rect 32036 35640 32088 35649
rect 24860 35572 24912 35624
rect 25044 35615 25096 35624
rect 25044 35581 25053 35615
rect 25053 35581 25087 35615
rect 25087 35581 25096 35615
rect 25044 35572 25096 35581
rect 20904 35504 20956 35556
rect 22560 35504 22612 35556
rect 27620 35572 27672 35624
rect 28448 35572 28500 35624
rect 30196 35615 30248 35624
rect 6644 35436 6696 35488
rect 7748 35436 7800 35488
rect 11244 35436 11296 35488
rect 18420 35436 18472 35488
rect 25504 35436 25556 35488
rect 28172 35436 28224 35488
rect 29736 35436 29788 35488
rect 30196 35581 30205 35615
rect 30205 35581 30239 35615
rect 30239 35581 30248 35615
rect 30196 35572 30248 35581
rect 32312 35649 32321 35683
rect 32321 35649 32355 35683
rect 32355 35649 32364 35683
rect 32312 35640 32364 35649
rect 35256 35640 35308 35692
rect 35440 35572 35492 35624
rect 30840 35436 30892 35488
rect 31300 35479 31352 35488
rect 31300 35445 31309 35479
rect 31309 35445 31343 35479
rect 31343 35445 31352 35479
rect 31300 35436 31352 35445
rect 32036 35436 32088 35488
rect 19606 35334 19658 35386
rect 19670 35334 19722 35386
rect 19734 35334 19786 35386
rect 19798 35334 19850 35386
rect 4068 35232 4120 35284
rect 10416 35275 10468 35284
rect 3608 35096 3660 35148
rect 4620 35096 4672 35148
rect 6184 35139 6236 35148
rect 6184 35105 6193 35139
rect 6193 35105 6227 35139
rect 6227 35105 6236 35139
rect 6184 35096 6236 35105
rect 6276 35096 6328 35148
rect 7656 35096 7708 35148
rect 10416 35241 10425 35275
rect 10425 35241 10459 35275
rect 10459 35241 10468 35275
rect 10416 35232 10468 35241
rect 19432 35232 19484 35284
rect 4804 35028 4856 35080
rect 7840 35028 7892 35080
rect 11244 35139 11296 35148
rect 11244 35105 11253 35139
rect 11253 35105 11287 35139
rect 11287 35105 11296 35139
rect 11244 35096 11296 35105
rect 11336 35096 11388 35148
rect 13636 35139 13688 35148
rect 13636 35105 13645 35139
rect 13645 35105 13679 35139
rect 13679 35105 13688 35139
rect 13636 35096 13688 35105
rect 16764 35164 16816 35216
rect 20904 35207 20956 35216
rect 20904 35173 20913 35207
rect 20913 35173 20947 35207
rect 20947 35173 20956 35207
rect 21640 35232 21692 35284
rect 22468 35232 22520 35284
rect 27436 35232 27488 35284
rect 30288 35232 30340 35284
rect 21272 35207 21324 35216
rect 20904 35164 20956 35173
rect 21272 35173 21281 35207
rect 21281 35173 21315 35207
rect 21315 35173 21324 35207
rect 21272 35164 21324 35173
rect 22008 35164 22060 35216
rect 16120 35139 16172 35148
rect 10968 35071 11020 35080
rect 10968 35037 10977 35071
rect 10977 35037 11011 35071
rect 11011 35037 11020 35071
rect 10968 35028 11020 35037
rect 6828 34960 6880 35012
rect 6460 34892 6512 34944
rect 12532 34935 12584 34944
rect 12532 34901 12541 34935
rect 12541 34901 12575 34935
rect 12575 34901 12584 34935
rect 12532 34892 12584 34901
rect 12624 34892 12676 34944
rect 16120 35105 16129 35139
rect 16129 35105 16163 35139
rect 16163 35105 16172 35139
rect 16120 35096 16172 35105
rect 16948 35096 17000 35148
rect 18972 35139 19024 35148
rect 18972 35105 18981 35139
rect 18981 35105 19015 35139
rect 19015 35105 19024 35139
rect 18972 35096 19024 35105
rect 19340 35139 19392 35148
rect 19340 35105 19349 35139
rect 19349 35105 19383 35139
rect 19383 35105 19392 35139
rect 19340 35096 19392 35105
rect 20260 35096 20312 35148
rect 20720 35096 20772 35148
rect 21456 35096 21508 35148
rect 22560 35096 22612 35148
rect 22652 35139 22704 35148
rect 22652 35105 22661 35139
rect 22661 35105 22695 35139
rect 22695 35105 22704 35139
rect 22652 35096 22704 35105
rect 23112 35139 23164 35148
rect 16304 35071 16356 35080
rect 16304 35037 16313 35071
rect 16313 35037 16347 35071
rect 16347 35037 16356 35071
rect 16304 35028 16356 35037
rect 16396 35028 16448 35080
rect 17132 35071 17184 35080
rect 17132 35037 17141 35071
rect 17141 35037 17175 35071
rect 17175 35037 17184 35071
rect 17132 35028 17184 35037
rect 20996 35028 21048 35080
rect 16580 34960 16632 35012
rect 22836 35071 22888 35080
rect 22836 35037 22845 35071
rect 22845 35037 22879 35071
rect 22879 35037 22888 35071
rect 22836 35028 22888 35037
rect 23112 35105 23121 35139
rect 23121 35105 23155 35139
rect 23155 35105 23164 35139
rect 23112 35096 23164 35105
rect 23204 35096 23256 35148
rect 25872 35164 25924 35216
rect 23756 35096 23808 35148
rect 25504 35139 25556 35148
rect 25504 35105 25513 35139
rect 25513 35105 25547 35139
rect 25547 35105 25556 35139
rect 25504 35096 25556 35105
rect 26608 35139 26660 35148
rect 26608 35105 26617 35139
rect 26617 35105 26651 35139
rect 26651 35105 26660 35139
rect 26608 35096 26660 35105
rect 27620 35139 27672 35148
rect 27620 35105 27629 35139
rect 27629 35105 27663 35139
rect 27663 35105 27672 35139
rect 27620 35096 27672 35105
rect 28724 35096 28776 35148
rect 29736 35096 29788 35148
rect 34152 35096 34204 35148
rect 34520 35139 34572 35148
rect 34520 35105 34529 35139
rect 34529 35105 34563 35139
rect 34563 35105 34572 35139
rect 34520 35096 34572 35105
rect 37924 35096 37976 35148
rect 38200 35139 38252 35148
rect 38200 35105 38209 35139
rect 38209 35105 38243 35139
rect 38243 35105 38252 35139
rect 38200 35096 38252 35105
rect 23388 35028 23440 35080
rect 25412 35071 25464 35080
rect 25412 35037 25421 35071
rect 25421 35037 25455 35071
rect 25455 35037 25464 35071
rect 25412 35028 25464 35037
rect 25964 35071 26016 35080
rect 25964 35037 25973 35071
rect 25973 35037 26007 35071
rect 26007 35037 26016 35071
rect 25964 35028 26016 35037
rect 27436 35028 27488 35080
rect 29276 35028 29328 35080
rect 29368 35071 29420 35080
rect 29368 35037 29377 35071
rect 29377 35037 29411 35071
rect 29411 35037 29420 35071
rect 29368 35028 29420 35037
rect 23572 34960 23624 35012
rect 32036 35028 32088 35080
rect 32864 35028 32916 35080
rect 35440 35028 35492 35080
rect 16212 34892 16264 34944
rect 26792 34935 26844 34944
rect 26792 34901 26801 34935
rect 26801 34901 26835 34935
rect 26835 34901 26844 34935
rect 26792 34892 26844 34901
rect 30932 34935 30984 34944
rect 30932 34901 30941 34935
rect 30941 34901 30975 34935
rect 30975 34901 30984 34935
rect 30932 34892 30984 34901
rect 33232 34892 33284 34944
rect 38108 34892 38160 34944
rect 4246 34790 4298 34842
rect 4310 34790 4362 34842
rect 4374 34790 4426 34842
rect 4438 34790 4490 34842
rect 34966 34790 35018 34842
rect 35030 34790 35082 34842
rect 35094 34790 35146 34842
rect 35158 34790 35210 34842
rect 16120 34688 16172 34740
rect 16764 34688 16816 34740
rect 19432 34688 19484 34740
rect 5080 34620 5132 34672
rect 5264 34620 5316 34672
rect 4712 34484 4764 34536
rect 4804 34484 4856 34536
rect 7748 34620 7800 34672
rect 16028 34620 16080 34672
rect 16488 34620 16540 34672
rect 6276 34595 6328 34604
rect 6276 34561 6285 34595
rect 6285 34561 6319 34595
rect 6319 34561 6328 34595
rect 6276 34552 6328 34561
rect 7104 34552 7156 34604
rect 6828 34527 6880 34536
rect 6828 34493 6837 34527
rect 6837 34493 6871 34527
rect 6871 34493 6880 34527
rect 6828 34484 6880 34493
rect 10968 34552 11020 34604
rect 7656 34527 7708 34536
rect 7656 34493 7665 34527
rect 7665 34493 7699 34527
rect 7699 34493 7708 34527
rect 7656 34484 7708 34493
rect 7748 34484 7800 34536
rect 9496 34527 9548 34536
rect 9496 34493 9505 34527
rect 9505 34493 9539 34527
rect 9539 34493 9548 34527
rect 9496 34484 9548 34493
rect 11336 34527 11388 34536
rect 11336 34493 11345 34527
rect 11345 34493 11379 34527
rect 11379 34493 11388 34527
rect 11336 34484 11388 34493
rect 12624 34484 12676 34536
rect 14924 34552 14976 34604
rect 15292 34595 15344 34604
rect 13820 34527 13872 34536
rect 12716 34416 12768 34468
rect 13820 34493 13829 34527
rect 13829 34493 13863 34527
rect 13863 34493 13872 34527
rect 13820 34484 13872 34493
rect 14372 34527 14424 34536
rect 14372 34493 14381 34527
rect 14381 34493 14415 34527
rect 14415 34493 14424 34527
rect 14372 34484 14424 34493
rect 15292 34561 15301 34595
rect 15301 34561 15335 34595
rect 15335 34561 15344 34595
rect 15292 34552 15344 34561
rect 15568 34552 15620 34604
rect 15844 34527 15896 34536
rect 15844 34493 15853 34527
rect 15853 34493 15887 34527
rect 15887 34493 15896 34527
rect 15844 34484 15896 34493
rect 16488 34527 16540 34536
rect 16488 34493 16497 34527
rect 16497 34493 16531 34527
rect 16531 34493 16540 34527
rect 16488 34484 16540 34493
rect 18972 34552 19024 34604
rect 20996 34552 21048 34604
rect 18328 34527 18380 34536
rect 18328 34493 18337 34527
rect 18337 34493 18371 34527
rect 18371 34493 18380 34527
rect 18328 34484 18380 34493
rect 3332 34348 3384 34400
rect 6920 34391 6972 34400
rect 6920 34357 6929 34391
rect 6929 34357 6963 34391
rect 6963 34357 6972 34391
rect 6920 34348 6972 34357
rect 11704 34348 11756 34400
rect 18696 34348 18748 34400
rect 20536 34527 20588 34536
rect 20536 34493 20545 34527
rect 20545 34493 20579 34527
rect 20579 34493 20588 34527
rect 20536 34484 20588 34493
rect 21456 34484 21508 34536
rect 23388 34620 23440 34672
rect 20168 34416 20220 34468
rect 20628 34416 20680 34468
rect 22100 34416 22152 34468
rect 21548 34348 21600 34400
rect 24308 34552 24360 34604
rect 22836 34527 22888 34536
rect 22836 34493 22845 34527
rect 22845 34493 22879 34527
rect 22879 34493 22888 34527
rect 22836 34484 22888 34493
rect 23480 34484 23532 34536
rect 23664 34527 23716 34536
rect 23664 34493 23673 34527
rect 23673 34493 23707 34527
rect 23707 34493 23716 34527
rect 23664 34484 23716 34493
rect 23020 34416 23072 34468
rect 25688 34688 25740 34740
rect 30196 34688 30248 34740
rect 28448 34620 28500 34672
rect 25044 34552 25096 34604
rect 25964 34552 26016 34604
rect 29276 34552 29328 34604
rect 29828 34595 29880 34604
rect 29828 34561 29837 34595
rect 29837 34561 29871 34595
rect 29871 34561 29880 34595
rect 29828 34552 29880 34561
rect 26332 34527 26384 34536
rect 26332 34493 26341 34527
rect 26341 34493 26375 34527
rect 26375 34493 26384 34527
rect 26332 34484 26384 34493
rect 28724 34484 28776 34536
rect 30656 34484 30708 34536
rect 31208 34620 31260 34672
rect 32496 34552 32548 34604
rect 26240 34416 26292 34468
rect 30196 34416 30248 34468
rect 32220 34527 32272 34536
rect 32220 34493 32229 34527
rect 32229 34493 32263 34527
rect 32263 34493 32272 34527
rect 32220 34484 32272 34493
rect 34060 34552 34112 34604
rect 35440 34552 35492 34604
rect 38016 34552 38068 34604
rect 38200 34552 38252 34604
rect 33140 34527 33192 34536
rect 33140 34493 33149 34527
rect 33149 34493 33183 34527
rect 33183 34493 33192 34527
rect 33140 34484 33192 34493
rect 33324 34527 33376 34536
rect 33324 34493 33333 34527
rect 33333 34493 33367 34527
rect 33367 34493 33376 34527
rect 33324 34484 33376 34493
rect 36084 34527 36136 34536
rect 36084 34493 36093 34527
rect 36093 34493 36127 34527
rect 36127 34493 36136 34527
rect 36084 34484 36136 34493
rect 36360 34527 36412 34536
rect 36360 34493 36369 34527
rect 36369 34493 36403 34527
rect 36403 34493 36412 34527
rect 36360 34484 36412 34493
rect 37372 34527 37424 34536
rect 37372 34493 37381 34527
rect 37381 34493 37415 34527
rect 37415 34493 37424 34527
rect 37372 34484 37424 34493
rect 35348 34348 35400 34400
rect 35716 34348 35768 34400
rect 19606 34246 19658 34298
rect 19670 34246 19722 34298
rect 19734 34246 19786 34298
rect 19798 34246 19850 34298
rect 7840 34144 7892 34196
rect 9496 34144 9548 34196
rect 17132 34144 17184 34196
rect 23848 34144 23900 34196
rect 28908 34144 28960 34196
rect 37372 34144 37424 34196
rect 2688 34008 2740 34060
rect 3608 34008 3660 34060
rect 6828 34008 6880 34060
rect 7104 34051 7156 34060
rect 7104 34017 7113 34051
rect 7113 34017 7147 34051
rect 7147 34017 7156 34051
rect 7104 34008 7156 34017
rect 8024 34051 8076 34060
rect 1860 33983 1912 33992
rect 1860 33949 1869 33983
rect 1869 33949 1903 33983
rect 1903 33949 1912 33983
rect 1860 33940 1912 33949
rect 5448 33940 5500 33992
rect 6184 33940 6236 33992
rect 8024 34017 8033 34051
rect 8033 34017 8067 34051
rect 8067 34017 8076 34051
rect 8024 34008 8076 34017
rect 8944 34051 8996 34060
rect 8944 34017 8953 34051
rect 8953 34017 8987 34051
rect 8987 34017 8996 34051
rect 8944 34008 8996 34017
rect 9864 34051 9916 34060
rect 9864 34017 9873 34051
rect 9873 34017 9907 34051
rect 9907 34017 9916 34051
rect 9864 34008 9916 34017
rect 11152 33983 11204 33992
rect 11152 33949 11161 33983
rect 11161 33949 11195 33983
rect 11195 33949 11204 33983
rect 11152 33940 11204 33949
rect 11888 34008 11940 34060
rect 12716 34051 12768 34060
rect 11704 33940 11756 33992
rect 12716 34017 12725 34051
rect 12725 34017 12759 34051
rect 12759 34017 12768 34051
rect 12716 34008 12768 34017
rect 13912 34076 13964 34128
rect 22652 34076 22704 34128
rect 12900 34008 12952 34060
rect 12532 33940 12584 33992
rect 13636 33940 13688 33992
rect 11060 33872 11112 33924
rect 12348 33872 12400 33924
rect 15108 34008 15160 34060
rect 16304 34051 16356 34060
rect 16304 34017 16313 34051
rect 16313 34017 16347 34051
rect 16347 34017 16356 34051
rect 16304 34008 16356 34017
rect 16948 34051 17000 34060
rect 16948 34017 16957 34051
rect 16957 34017 16991 34051
rect 16991 34017 17000 34051
rect 16948 34008 17000 34017
rect 17316 34008 17368 34060
rect 18236 34008 18288 34060
rect 18696 34051 18748 34060
rect 18696 34017 18705 34051
rect 18705 34017 18739 34051
rect 18739 34017 18748 34051
rect 18696 34008 18748 34017
rect 21180 34051 21232 34060
rect 21180 34017 21189 34051
rect 21189 34017 21223 34051
rect 21223 34017 21232 34051
rect 21180 34008 21232 34017
rect 21364 34051 21416 34060
rect 21364 34017 21373 34051
rect 21373 34017 21407 34051
rect 21407 34017 21416 34051
rect 21364 34008 21416 34017
rect 21640 34051 21692 34060
rect 21640 34017 21649 34051
rect 21649 34017 21683 34051
rect 21683 34017 21692 34051
rect 21640 34008 21692 34017
rect 22100 34008 22152 34060
rect 23480 34051 23532 34060
rect 23480 34017 23489 34051
rect 23489 34017 23523 34051
rect 23523 34017 23532 34051
rect 23480 34008 23532 34017
rect 26608 34076 26660 34128
rect 26332 34008 26384 34060
rect 26792 34051 26844 34060
rect 15200 33940 15252 33992
rect 16488 33983 16540 33992
rect 16488 33949 16497 33983
rect 16497 33949 16531 33983
rect 16531 33949 16540 33983
rect 16488 33940 16540 33949
rect 17224 33940 17276 33992
rect 23756 33940 23808 33992
rect 24584 33983 24636 33992
rect 24584 33949 24593 33983
rect 24593 33949 24627 33983
rect 24627 33949 24636 33983
rect 24584 33940 24636 33949
rect 26792 34017 26801 34051
rect 26801 34017 26835 34051
rect 26835 34017 26844 34051
rect 26792 34008 26844 34017
rect 29644 34008 29696 34060
rect 32864 34008 32916 34060
rect 33140 34008 33192 34060
rect 34796 34051 34848 34060
rect 34796 34017 34805 34051
rect 34805 34017 34839 34051
rect 34839 34017 34848 34051
rect 34796 34008 34848 34017
rect 35440 34051 35492 34060
rect 35440 34017 35449 34051
rect 35449 34017 35483 34051
rect 35483 34017 35492 34051
rect 35440 34008 35492 34017
rect 35716 34051 35768 34060
rect 35716 34017 35725 34051
rect 35725 34017 35759 34051
rect 35759 34017 35768 34051
rect 35716 34008 35768 34017
rect 35808 34008 35860 34060
rect 38292 34051 38344 34060
rect 38292 34017 38301 34051
rect 38301 34017 38335 34051
rect 38335 34017 38344 34051
rect 38292 34008 38344 34017
rect 29552 33940 29604 33992
rect 29828 33940 29880 33992
rect 32404 33983 32456 33992
rect 32404 33949 32413 33983
rect 32413 33949 32447 33983
rect 32447 33949 32456 33983
rect 32404 33940 32456 33949
rect 37648 33940 37700 33992
rect 29736 33872 29788 33924
rect 3240 33804 3292 33856
rect 5632 33847 5684 33856
rect 5632 33813 5641 33847
rect 5641 33813 5675 33847
rect 5675 33813 5684 33847
rect 5632 33804 5684 33813
rect 9680 33804 9732 33856
rect 12992 33804 13044 33856
rect 15936 33804 15988 33856
rect 19984 33847 20036 33856
rect 19984 33813 19993 33847
rect 19993 33813 20027 33847
rect 20027 33813 20036 33847
rect 19984 33804 20036 33813
rect 22376 33804 22428 33856
rect 26700 33804 26752 33856
rect 30380 33804 30432 33856
rect 33508 33847 33560 33856
rect 33508 33813 33517 33847
rect 33517 33813 33551 33847
rect 33551 33813 33560 33847
rect 33508 33804 33560 33813
rect 34336 33847 34388 33856
rect 34336 33813 34345 33847
rect 34345 33813 34379 33847
rect 34379 33813 34388 33847
rect 34336 33804 34388 33813
rect 36636 33804 36688 33856
rect 4246 33702 4298 33754
rect 4310 33702 4362 33754
rect 4374 33702 4426 33754
rect 4438 33702 4490 33754
rect 34966 33702 35018 33754
rect 35030 33702 35082 33754
rect 35094 33702 35146 33754
rect 35158 33702 35210 33754
rect 5448 33643 5500 33652
rect 5448 33609 5457 33643
rect 5457 33609 5491 33643
rect 5491 33609 5500 33643
rect 5448 33600 5500 33609
rect 7656 33600 7708 33652
rect 9864 33600 9916 33652
rect 13820 33643 13872 33652
rect 13820 33609 13829 33643
rect 13829 33609 13863 33643
rect 13863 33609 13872 33643
rect 13820 33600 13872 33609
rect 16948 33600 17000 33652
rect 17224 33643 17276 33652
rect 17224 33609 17233 33643
rect 17233 33609 17267 33643
rect 17267 33609 17276 33643
rect 17224 33600 17276 33609
rect 20260 33600 20312 33652
rect 22652 33600 22704 33652
rect 24584 33600 24636 33652
rect 28632 33643 28684 33652
rect 28632 33609 28641 33643
rect 28641 33609 28675 33643
rect 28675 33609 28684 33643
rect 28632 33600 28684 33609
rect 28908 33600 28960 33652
rect 29184 33600 29236 33652
rect 29552 33643 29604 33652
rect 29552 33609 29561 33643
rect 29561 33609 29595 33643
rect 29595 33609 29604 33643
rect 29552 33600 29604 33609
rect 30564 33643 30616 33652
rect 30564 33609 30573 33643
rect 30573 33609 30607 33643
rect 30607 33609 30616 33643
rect 30564 33600 30616 33609
rect 34060 33643 34112 33652
rect 34060 33609 34069 33643
rect 34069 33609 34103 33643
rect 34103 33609 34112 33643
rect 34060 33600 34112 33609
rect 1584 33532 1636 33584
rect 8944 33532 8996 33584
rect 11520 33532 11572 33584
rect 19064 33532 19116 33584
rect 3240 33464 3292 33516
rect 2136 33439 2188 33448
rect 2136 33405 2145 33439
rect 2145 33405 2179 33439
rect 2179 33405 2188 33439
rect 2136 33396 2188 33405
rect 3332 33439 3384 33448
rect 2780 33328 2832 33380
rect 2872 33328 2924 33380
rect 3332 33405 3341 33439
rect 3341 33405 3375 33439
rect 3375 33405 3384 33439
rect 3332 33396 3384 33405
rect 5080 33464 5132 33516
rect 10416 33464 10468 33516
rect 3608 33328 3660 33380
rect 4620 33396 4672 33448
rect 5264 33439 5316 33448
rect 5264 33405 5273 33439
rect 5273 33405 5307 33439
rect 5307 33405 5316 33439
rect 5264 33396 5316 33405
rect 7196 33439 7248 33448
rect 7196 33405 7205 33439
rect 7205 33405 7239 33439
rect 7239 33405 7248 33439
rect 7196 33396 7248 33405
rect 8208 33396 8260 33448
rect 9680 33439 9732 33448
rect 4896 33328 4948 33380
rect 9680 33405 9689 33439
rect 9689 33405 9723 33439
rect 9723 33405 9732 33439
rect 9680 33396 9732 33405
rect 10048 33439 10100 33448
rect 10048 33405 10057 33439
rect 10057 33405 10091 33439
rect 10091 33405 10100 33439
rect 10048 33396 10100 33405
rect 11152 33439 11204 33448
rect 2044 33260 2096 33312
rect 9772 33328 9824 33380
rect 11152 33405 11161 33439
rect 11161 33405 11195 33439
rect 11195 33405 11204 33439
rect 11152 33396 11204 33405
rect 12348 33464 12400 33516
rect 13268 33464 13320 33516
rect 12900 33396 12952 33448
rect 13912 33396 13964 33448
rect 15292 33464 15344 33516
rect 15936 33507 15988 33516
rect 15936 33473 15945 33507
rect 15945 33473 15979 33507
rect 15979 33473 15988 33507
rect 15936 33464 15988 33473
rect 23480 33532 23532 33584
rect 23572 33532 23624 33584
rect 35808 33575 35860 33584
rect 35808 33541 35817 33575
rect 35817 33541 35851 33575
rect 35851 33541 35860 33575
rect 35808 33532 35860 33541
rect 15200 33439 15252 33448
rect 15200 33405 15209 33439
rect 15209 33405 15243 33439
rect 15243 33405 15252 33439
rect 15200 33396 15252 33405
rect 15660 33439 15712 33448
rect 15660 33405 15669 33439
rect 15669 33405 15703 33439
rect 15703 33405 15712 33439
rect 15660 33396 15712 33405
rect 16396 33396 16448 33448
rect 18328 33396 18380 33448
rect 18972 33439 19024 33448
rect 11060 33328 11112 33380
rect 11612 33328 11664 33380
rect 13820 33328 13872 33380
rect 18972 33405 18981 33439
rect 18981 33405 19015 33439
rect 19015 33405 19024 33439
rect 18972 33396 19024 33405
rect 19892 33396 19944 33448
rect 21548 33464 21600 33516
rect 24400 33464 24452 33516
rect 26240 33464 26292 33516
rect 21364 33396 21416 33448
rect 19064 33328 19116 33380
rect 21824 33439 21876 33448
rect 21824 33405 21833 33439
rect 21833 33405 21867 33439
rect 21867 33405 21876 33439
rect 22376 33439 22428 33448
rect 21824 33396 21876 33405
rect 22376 33405 22385 33439
rect 22385 33405 22419 33439
rect 22419 33405 22428 33439
rect 22376 33396 22428 33405
rect 23572 33396 23624 33448
rect 23756 33396 23808 33448
rect 23940 33439 23992 33448
rect 23940 33405 23949 33439
rect 23949 33405 23983 33439
rect 23983 33405 23992 33439
rect 23940 33396 23992 33405
rect 25044 33396 25096 33448
rect 27160 33396 27212 33448
rect 27344 33396 27396 33448
rect 27804 33439 27856 33448
rect 27804 33405 27813 33439
rect 27813 33405 27847 33439
rect 27847 33405 27856 33439
rect 27804 33396 27856 33405
rect 27896 33439 27948 33448
rect 27896 33405 27905 33439
rect 27905 33405 27939 33439
rect 27939 33405 27948 33439
rect 27896 33396 27948 33405
rect 26792 33371 26844 33380
rect 8576 33303 8628 33312
rect 8576 33269 8585 33303
rect 8585 33269 8619 33303
rect 8619 33269 8628 33303
rect 8576 33260 8628 33269
rect 10416 33260 10468 33312
rect 11704 33260 11756 33312
rect 17684 33260 17736 33312
rect 18144 33303 18196 33312
rect 18144 33269 18153 33303
rect 18153 33269 18187 33303
rect 18187 33269 18196 33303
rect 18144 33260 18196 33269
rect 19248 33260 19300 33312
rect 26792 33337 26801 33371
rect 26801 33337 26835 33371
rect 26835 33337 26844 33371
rect 26792 33328 26844 33337
rect 28172 33464 28224 33516
rect 32404 33464 32456 33516
rect 32864 33464 32916 33516
rect 34336 33464 34388 33516
rect 28448 33439 28500 33448
rect 28448 33405 28457 33439
rect 28457 33405 28491 33439
rect 28491 33405 28500 33439
rect 28448 33396 28500 33405
rect 30380 33439 30432 33448
rect 20076 33303 20128 33312
rect 20076 33269 20085 33303
rect 20085 33269 20119 33303
rect 20119 33269 20128 33303
rect 20076 33260 20128 33269
rect 30380 33405 30389 33439
rect 30389 33405 30423 33439
rect 30423 33405 30432 33439
rect 30380 33396 30432 33405
rect 31944 33439 31996 33448
rect 31944 33405 31953 33439
rect 31953 33405 31987 33439
rect 31987 33405 31996 33439
rect 31944 33396 31996 33405
rect 33600 33396 33652 33448
rect 35808 33439 35860 33448
rect 32312 33328 32364 33380
rect 35808 33405 35817 33439
rect 35817 33405 35851 33439
rect 35851 33405 35860 33439
rect 35808 33396 35860 33405
rect 36636 33396 36688 33448
rect 38476 33532 38528 33584
rect 38292 33507 38344 33516
rect 38292 33473 38301 33507
rect 38301 33473 38335 33507
rect 38335 33473 38344 33507
rect 38292 33464 38344 33473
rect 38108 33439 38160 33448
rect 38108 33405 38117 33439
rect 38117 33405 38151 33439
rect 38151 33405 38160 33439
rect 38108 33396 38160 33405
rect 29920 33303 29972 33312
rect 29920 33269 29929 33303
rect 29929 33269 29963 33303
rect 29963 33269 29972 33303
rect 29920 33260 29972 33269
rect 34520 33260 34572 33312
rect 36728 33328 36780 33380
rect 36360 33260 36412 33312
rect 37648 33260 37700 33312
rect 19606 33158 19658 33210
rect 19670 33158 19722 33210
rect 19734 33158 19786 33210
rect 19798 33158 19850 33210
rect 4804 33056 4856 33108
rect 5172 33056 5224 33108
rect 13912 33056 13964 33108
rect 1860 32988 1912 33040
rect 5080 33031 5132 33040
rect 5080 32997 5089 33031
rect 5089 32997 5123 33031
rect 5123 32997 5132 33031
rect 5080 32988 5132 32997
rect 5632 32988 5684 33040
rect 2872 32963 2924 32972
rect 2872 32929 2881 32963
rect 2881 32929 2915 32963
rect 2915 32929 2924 32963
rect 2872 32920 2924 32929
rect 3148 32963 3200 32972
rect 3148 32929 3157 32963
rect 3157 32929 3191 32963
rect 3191 32929 3200 32963
rect 3148 32920 3200 32929
rect 3240 32920 3292 32972
rect 5264 32920 5316 32972
rect 6276 32963 6328 32972
rect 6276 32929 6285 32963
rect 6285 32929 6319 32963
rect 6319 32929 6328 32963
rect 6276 32920 6328 32929
rect 6460 32988 6512 33040
rect 10048 33031 10100 33040
rect 10048 32997 10057 33031
rect 10057 32997 10091 33031
rect 10091 32997 10100 33031
rect 10048 32988 10100 32997
rect 12440 33031 12492 33040
rect 12440 32997 12449 33031
rect 12449 32997 12483 33031
rect 12483 32997 12492 33031
rect 12440 32988 12492 32997
rect 12624 32988 12676 33040
rect 16580 33056 16632 33108
rect 17316 33056 17368 33108
rect 20168 33056 20220 33108
rect 24492 33056 24544 33108
rect 4896 32852 4948 32904
rect 8024 32920 8076 32972
rect 8668 32920 8720 32972
rect 10416 32963 10468 32972
rect 10416 32929 10425 32963
rect 10425 32929 10459 32963
rect 10459 32929 10468 32963
rect 10416 32920 10468 32929
rect 11060 32963 11112 32972
rect 11060 32929 11069 32963
rect 11069 32929 11103 32963
rect 11103 32929 11112 32963
rect 11060 32920 11112 32929
rect 11612 32963 11664 32972
rect 11612 32929 11621 32963
rect 11621 32929 11655 32963
rect 11655 32929 11664 32963
rect 11612 32920 11664 32929
rect 12256 32963 12308 32972
rect 12256 32929 12265 32963
rect 12265 32929 12299 32963
rect 12299 32929 12308 32963
rect 12256 32920 12308 32929
rect 15476 32963 15528 32972
rect 11796 32852 11848 32904
rect 15476 32929 15485 32963
rect 15485 32929 15519 32963
rect 15519 32929 15528 32963
rect 15476 32920 15528 32929
rect 15568 32963 15620 32972
rect 15568 32929 15577 32963
rect 15577 32929 15611 32963
rect 15611 32929 15620 32963
rect 17224 32988 17276 33040
rect 15568 32920 15620 32929
rect 16948 32963 17000 32972
rect 7196 32784 7248 32836
rect 11980 32784 12032 32836
rect 13820 32895 13872 32904
rect 13820 32861 13829 32895
rect 13829 32861 13863 32895
rect 13863 32861 13872 32895
rect 13820 32852 13872 32861
rect 14280 32895 14332 32904
rect 14280 32861 14289 32895
rect 14289 32861 14323 32895
rect 14323 32861 14332 32895
rect 14280 32852 14332 32861
rect 15292 32895 15344 32904
rect 15292 32861 15301 32895
rect 15301 32861 15335 32895
rect 15335 32861 15344 32895
rect 15292 32852 15344 32861
rect 16948 32929 16957 32963
rect 16957 32929 16991 32963
rect 16991 32929 17000 32963
rect 16948 32920 17000 32929
rect 17500 32963 17552 32972
rect 17500 32929 17509 32963
rect 17509 32929 17543 32963
rect 17543 32929 17552 32963
rect 17500 32920 17552 32929
rect 18144 32920 18196 32972
rect 18328 32963 18380 32972
rect 18328 32929 18337 32963
rect 18337 32929 18371 32963
rect 18371 32929 18380 32963
rect 18328 32920 18380 32929
rect 19064 32963 19116 32972
rect 19064 32929 19073 32963
rect 19073 32929 19107 32963
rect 19107 32929 19116 32963
rect 19064 32920 19116 32929
rect 19984 32920 20036 32972
rect 22192 32988 22244 33040
rect 22100 32963 22152 32972
rect 22100 32929 22109 32963
rect 22109 32929 22143 32963
rect 22143 32929 22152 32963
rect 22100 32920 22152 32929
rect 22836 32920 22888 32972
rect 23480 32963 23532 32972
rect 23480 32929 23489 32963
rect 23489 32929 23523 32963
rect 23523 32929 23532 32963
rect 23480 32920 23532 32929
rect 30840 33056 30892 33108
rect 31116 33056 31168 33108
rect 33232 33056 33284 33108
rect 25504 32920 25556 32972
rect 27160 32920 27212 32972
rect 19248 32852 19300 32904
rect 20260 32852 20312 32904
rect 24860 32852 24912 32904
rect 26332 32852 26384 32904
rect 27712 32895 27764 32904
rect 27712 32861 27721 32895
rect 27721 32861 27755 32895
rect 27755 32861 27764 32895
rect 27712 32852 27764 32861
rect 29552 32852 29604 32904
rect 30564 32920 30616 32972
rect 33508 32988 33560 33040
rect 35348 33031 35400 33040
rect 35348 32997 35357 33031
rect 35357 32997 35391 33031
rect 35391 32997 35400 33031
rect 35348 32988 35400 32997
rect 37924 32988 37976 33040
rect 31668 32852 31720 32904
rect 33324 32920 33376 32972
rect 34060 32920 34112 32972
rect 34520 32920 34572 32972
rect 35808 32920 35860 32972
rect 36452 32920 36504 32972
rect 36728 32920 36780 32972
rect 36912 32963 36964 32972
rect 36912 32929 36921 32963
rect 36921 32929 36955 32963
rect 36955 32929 36964 32963
rect 36912 32920 36964 32929
rect 38568 32920 38620 32972
rect 36268 32895 36320 32904
rect 36268 32861 36277 32895
rect 36277 32861 36311 32895
rect 36311 32861 36320 32895
rect 36268 32852 36320 32861
rect 38752 32895 38804 32904
rect 38752 32861 38761 32895
rect 38761 32861 38795 32895
rect 38795 32861 38804 32895
rect 38752 32852 38804 32861
rect 15936 32784 15988 32836
rect 16856 32827 16908 32836
rect 16856 32793 16865 32827
rect 16865 32793 16899 32827
rect 16899 32793 16908 32827
rect 16856 32784 16908 32793
rect 19064 32784 19116 32836
rect 19156 32784 19208 32836
rect 21824 32784 21876 32836
rect 32312 32827 32364 32836
rect 32312 32793 32321 32827
rect 32321 32793 32355 32827
rect 32355 32793 32364 32827
rect 32312 32784 32364 32793
rect 32772 32784 32824 32836
rect 36084 32784 36136 32836
rect 3608 32716 3660 32768
rect 10416 32716 10468 32768
rect 17868 32716 17920 32768
rect 21732 32716 21784 32768
rect 22468 32716 22520 32768
rect 23480 32716 23532 32768
rect 24584 32716 24636 32768
rect 29092 32716 29144 32768
rect 4246 32614 4298 32666
rect 4310 32614 4362 32666
rect 4374 32614 4426 32666
rect 4438 32614 4490 32666
rect 34966 32614 35018 32666
rect 35030 32614 35082 32666
rect 35094 32614 35146 32666
rect 35158 32614 35210 32666
rect 6184 32555 6236 32564
rect 6184 32521 6193 32555
rect 6193 32521 6227 32555
rect 6227 32521 6236 32555
rect 6184 32512 6236 32521
rect 8208 32555 8260 32564
rect 8208 32521 8217 32555
rect 8217 32521 8251 32555
rect 8251 32521 8260 32555
rect 8208 32512 8260 32521
rect 15476 32512 15528 32564
rect 3424 32444 3476 32496
rect 11060 32444 11112 32496
rect 12440 32444 12492 32496
rect 12716 32487 12768 32496
rect 12716 32453 12725 32487
rect 12725 32453 12759 32487
rect 12759 32453 12768 32487
rect 12716 32444 12768 32453
rect 3148 32376 3200 32428
rect 1860 32240 1912 32292
rect 2780 32308 2832 32360
rect 3056 32308 3108 32360
rect 5080 32308 5132 32360
rect 5632 32376 5684 32428
rect 8576 32376 8628 32428
rect 9680 32376 9732 32428
rect 12624 32376 12676 32428
rect 3332 32172 3384 32224
rect 4712 32172 4764 32224
rect 5540 32351 5592 32360
rect 5540 32317 5549 32351
rect 5549 32317 5583 32351
rect 5583 32317 5592 32351
rect 5540 32308 5592 32317
rect 5264 32240 5316 32292
rect 6736 32308 6788 32360
rect 7104 32351 7156 32360
rect 7104 32317 7113 32351
rect 7113 32317 7147 32351
rect 7147 32317 7156 32351
rect 7104 32308 7156 32317
rect 9312 32308 9364 32360
rect 11520 32308 11572 32360
rect 12532 32351 12584 32360
rect 12532 32317 12541 32351
rect 12541 32317 12575 32351
rect 12575 32317 12584 32351
rect 12532 32308 12584 32317
rect 12900 32308 12952 32360
rect 10416 32240 10468 32292
rect 13820 32376 13872 32428
rect 14280 32376 14332 32428
rect 14832 32376 14884 32428
rect 14372 32351 14424 32360
rect 14372 32317 14381 32351
rect 14381 32317 14415 32351
rect 14415 32317 14424 32351
rect 14372 32308 14424 32317
rect 14556 32351 14608 32360
rect 14556 32317 14565 32351
rect 14565 32317 14599 32351
rect 14599 32317 14608 32351
rect 14556 32308 14608 32317
rect 15384 32376 15436 32428
rect 15660 32419 15712 32428
rect 15660 32385 15669 32419
rect 15669 32385 15703 32419
rect 15703 32385 15712 32419
rect 15660 32376 15712 32385
rect 15936 32419 15988 32428
rect 15936 32385 15945 32419
rect 15945 32385 15979 32419
rect 15979 32385 15988 32419
rect 15936 32376 15988 32385
rect 16396 32376 16448 32428
rect 19984 32512 20036 32564
rect 21732 32512 21784 32564
rect 23480 32512 23532 32564
rect 23572 32512 23624 32564
rect 29368 32512 29420 32564
rect 39028 32555 39080 32564
rect 17500 32444 17552 32496
rect 19156 32444 19208 32496
rect 18604 32351 18656 32360
rect 14464 32240 14516 32292
rect 6644 32172 6696 32224
rect 9496 32172 9548 32224
rect 11796 32215 11848 32224
rect 11796 32181 11805 32215
rect 11805 32181 11839 32215
rect 11839 32181 11848 32215
rect 11796 32172 11848 32181
rect 18604 32317 18613 32351
rect 18613 32317 18647 32351
rect 18647 32317 18656 32351
rect 18604 32308 18656 32317
rect 26792 32444 26844 32496
rect 20076 32376 20128 32428
rect 21180 32376 21232 32428
rect 29092 32444 29144 32496
rect 19340 32308 19392 32360
rect 21824 32308 21876 32360
rect 20260 32240 20312 32292
rect 22100 32308 22152 32360
rect 23572 32308 23624 32360
rect 22192 32240 22244 32292
rect 23848 32308 23900 32360
rect 24400 32351 24452 32360
rect 24400 32317 24409 32351
rect 24409 32317 24443 32351
rect 24443 32317 24452 32351
rect 24400 32308 24452 32317
rect 25320 32351 25372 32360
rect 25320 32317 25329 32351
rect 25329 32317 25363 32351
rect 25363 32317 25372 32351
rect 25320 32308 25372 32317
rect 27160 32351 27212 32360
rect 23756 32240 23808 32292
rect 27160 32317 27169 32351
rect 27169 32317 27203 32351
rect 27203 32317 27212 32351
rect 27160 32308 27212 32317
rect 27344 32351 27396 32360
rect 27344 32317 27353 32351
rect 27353 32317 27387 32351
rect 27387 32317 27396 32351
rect 27344 32308 27396 32317
rect 30380 32376 30432 32428
rect 39028 32521 39037 32555
rect 39037 32521 39071 32555
rect 39071 32521 39080 32555
rect 39028 32512 39080 32521
rect 35348 32444 35400 32496
rect 36912 32419 36964 32428
rect 36912 32385 36921 32419
rect 36921 32385 36955 32419
rect 36955 32385 36964 32419
rect 36912 32376 36964 32385
rect 27896 32351 27948 32360
rect 27896 32317 27905 32351
rect 27905 32317 27939 32351
rect 27939 32317 27948 32351
rect 27896 32308 27948 32317
rect 20076 32172 20128 32224
rect 22284 32172 22336 32224
rect 22560 32172 22612 32224
rect 26056 32240 26108 32292
rect 29000 32240 29052 32292
rect 29552 32308 29604 32360
rect 31668 32351 31720 32360
rect 31668 32317 31677 32351
rect 31677 32317 31711 32351
rect 31711 32317 31720 32351
rect 31668 32308 31720 32317
rect 32956 32351 33008 32360
rect 32956 32317 32965 32351
rect 32965 32317 32999 32351
rect 32999 32317 33008 32351
rect 32956 32308 33008 32317
rect 33324 32351 33376 32360
rect 33324 32317 33333 32351
rect 33333 32317 33367 32351
rect 33367 32317 33376 32351
rect 33324 32308 33376 32317
rect 33784 32308 33836 32360
rect 35808 32351 35860 32360
rect 33232 32240 33284 32292
rect 34520 32240 34572 32292
rect 35808 32317 35817 32351
rect 35817 32317 35851 32351
rect 35851 32317 35860 32351
rect 35808 32308 35860 32317
rect 36636 32351 36688 32360
rect 36636 32317 36645 32351
rect 36645 32317 36679 32351
rect 36679 32317 36688 32351
rect 36636 32308 36688 32317
rect 36544 32240 36596 32292
rect 37924 32376 37976 32428
rect 37464 32351 37516 32360
rect 37464 32317 37473 32351
rect 37473 32317 37507 32351
rect 37507 32317 37516 32351
rect 37464 32308 37516 32317
rect 37740 32351 37792 32360
rect 37740 32317 37749 32351
rect 37749 32317 37783 32351
rect 37783 32317 37792 32351
rect 37740 32308 37792 32317
rect 25228 32172 25280 32224
rect 27344 32172 27396 32224
rect 30012 32172 30064 32224
rect 33508 32172 33560 32224
rect 19606 32070 19658 32122
rect 19670 32070 19722 32122
rect 19734 32070 19786 32122
rect 19798 32070 19850 32122
rect 2688 31968 2740 32020
rect 1400 31875 1452 31884
rect 1400 31841 1409 31875
rect 1409 31841 1443 31875
rect 1443 31841 1452 31875
rect 1400 31832 1452 31841
rect 1676 31807 1728 31816
rect 1676 31773 1685 31807
rect 1685 31773 1719 31807
rect 1719 31773 1728 31807
rect 1676 31764 1728 31773
rect 5080 31968 5132 32020
rect 4620 31900 4672 31952
rect 3884 31875 3936 31884
rect 3884 31841 3893 31875
rect 3893 31841 3927 31875
rect 3927 31841 3936 31875
rect 3884 31832 3936 31841
rect 4712 31832 4764 31884
rect 4988 31875 5040 31884
rect 4988 31841 4997 31875
rect 4997 31841 5031 31875
rect 5031 31841 5040 31875
rect 4988 31832 5040 31841
rect 5172 31875 5224 31884
rect 5172 31841 5181 31875
rect 5181 31841 5215 31875
rect 5215 31841 5224 31875
rect 5172 31832 5224 31841
rect 5264 31832 5316 31884
rect 7104 31968 7156 32020
rect 6276 31900 6328 31952
rect 6920 31875 6972 31884
rect 5448 31764 5500 31816
rect 6920 31841 6929 31875
rect 6929 31841 6963 31875
rect 6963 31841 6972 31875
rect 6920 31832 6972 31841
rect 9496 31900 9548 31952
rect 8760 31832 8812 31884
rect 9588 31832 9640 31884
rect 11796 31968 11848 32020
rect 10508 31875 10560 31884
rect 7012 31764 7064 31816
rect 10508 31841 10517 31875
rect 10517 31841 10551 31875
rect 10551 31841 10560 31875
rect 10508 31832 10560 31841
rect 10876 31832 10928 31884
rect 12256 31875 12308 31884
rect 12256 31841 12265 31875
rect 12265 31841 12299 31875
rect 12299 31841 12308 31875
rect 12256 31832 12308 31841
rect 12716 31900 12768 31952
rect 15660 31900 15712 31952
rect 10416 31764 10468 31816
rect 11980 31764 12032 31816
rect 12440 31764 12492 31816
rect 15476 31832 15528 31884
rect 17868 31968 17920 32020
rect 17132 31900 17184 31952
rect 18420 31943 18472 31952
rect 17224 31875 17276 31884
rect 4804 31696 4856 31748
rect 9772 31739 9824 31748
rect 9772 31705 9781 31739
rect 9781 31705 9815 31739
rect 9815 31705 9824 31739
rect 9772 31696 9824 31705
rect 14464 31764 14516 31816
rect 15200 31764 15252 31816
rect 16948 31764 17000 31816
rect 17224 31841 17233 31875
rect 17233 31841 17267 31875
rect 17267 31841 17276 31875
rect 17224 31832 17276 31841
rect 18420 31909 18429 31943
rect 18429 31909 18463 31943
rect 18463 31909 18472 31943
rect 18420 31900 18472 31909
rect 18788 31968 18840 32020
rect 19432 31968 19484 32020
rect 23940 31968 23992 32020
rect 33784 32011 33836 32020
rect 18604 31900 18656 31952
rect 19248 31900 19300 31952
rect 17592 31764 17644 31816
rect 18880 31832 18932 31884
rect 18972 31875 19024 31884
rect 18972 31841 18981 31875
rect 18981 31841 19015 31875
rect 19015 31841 19024 31875
rect 18972 31832 19024 31841
rect 19340 31832 19392 31884
rect 19432 31875 19484 31884
rect 19432 31841 19441 31875
rect 19441 31841 19475 31875
rect 19475 31841 19484 31875
rect 19432 31832 19484 31841
rect 19984 31832 20036 31884
rect 20352 31875 20404 31884
rect 20352 31841 20361 31875
rect 20361 31841 20395 31875
rect 20395 31841 20404 31875
rect 20352 31832 20404 31841
rect 20996 31832 21048 31884
rect 21272 31875 21324 31884
rect 21272 31841 21281 31875
rect 21281 31841 21315 31875
rect 21315 31841 21324 31875
rect 21272 31832 21324 31841
rect 24308 31900 24360 31952
rect 24768 31900 24820 31952
rect 22468 31875 22520 31884
rect 22468 31841 22477 31875
rect 22477 31841 22511 31875
rect 22511 31841 22520 31875
rect 22468 31832 22520 31841
rect 23664 31875 23716 31884
rect 23664 31841 23673 31875
rect 23673 31841 23707 31875
rect 23707 31841 23716 31875
rect 23664 31832 23716 31841
rect 25228 31832 25280 31884
rect 22008 31764 22060 31816
rect 23296 31807 23348 31816
rect 23296 31773 23305 31807
rect 23305 31773 23339 31807
rect 23339 31773 23348 31807
rect 23296 31764 23348 31773
rect 23572 31764 23624 31816
rect 17224 31696 17276 31748
rect 18972 31696 19024 31748
rect 19800 31696 19852 31748
rect 2504 31628 2556 31680
rect 2780 31628 2832 31680
rect 3516 31628 3568 31680
rect 14832 31628 14884 31680
rect 20352 31628 20404 31680
rect 21824 31696 21876 31748
rect 23848 31628 23900 31680
rect 25688 31832 25740 31884
rect 26332 31832 26384 31884
rect 26148 31764 26200 31816
rect 25688 31696 25740 31748
rect 27528 31875 27580 31884
rect 27528 31841 27537 31875
rect 27537 31841 27571 31875
rect 27571 31841 27580 31875
rect 27528 31832 27580 31841
rect 28172 31875 28224 31884
rect 28172 31841 28181 31875
rect 28181 31841 28215 31875
rect 28215 31841 28224 31875
rect 28172 31832 28224 31841
rect 28816 31832 28868 31884
rect 33784 31977 33793 32011
rect 33793 31977 33827 32011
rect 33827 31977 33836 32011
rect 33784 31968 33836 31977
rect 36268 31968 36320 32020
rect 30840 31943 30892 31952
rect 30840 31909 30849 31943
rect 30849 31909 30883 31943
rect 30883 31909 30892 31943
rect 30840 31900 30892 31909
rect 30012 31875 30064 31884
rect 30012 31841 30021 31875
rect 30021 31841 30055 31875
rect 30055 31841 30064 31875
rect 30012 31832 30064 31841
rect 30104 31832 30156 31884
rect 27896 31764 27948 31816
rect 28448 31764 28500 31816
rect 28632 31764 28684 31816
rect 28908 31764 28960 31816
rect 30196 31764 30248 31816
rect 30932 31832 30984 31884
rect 31024 31764 31076 31816
rect 31760 31764 31812 31816
rect 32496 31807 32548 31816
rect 27252 31628 27304 31680
rect 27712 31628 27764 31680
rect 32496 31773 32505 31807
rect 32505 31773 32539 31807
rect 32539 31773 32548 31807
rect 32496 31764 32548 31773
rect 35532 31832 35584 31884
rect 38016 31875 38068 31884
rect 38016 31841 38025 31875
rect 38025 31841 38059 31875
rect 38059 31841 38068 31875
rect 38016 31832 38068 31841
rect 38292 31832 38344 31884
rect 38476 31900 38528 31952
rect 38752 31875 38804 31884
rect 38752 31841 38761 31875
rect 38761 31841 38795 31875
rect 38795 31841 38804 31875
rect 38752 31832 38804 31841
rect 34704 31764 34756 31816
rect 35256 31807 35308 31816
rect 35256 31773 35265 31807
rect 35265 31773 35299 31807
rect 35299 31773 35308 31807
rect 35256 31764 35308 31773
rect 38476 31764 38528 31816
rect 32680 31628 32732 31680
rect 35440 31628 35492 31680
rect 4246 31526 4298 31578
rect 4310 31526 4362 31578
rect 4374 31526 4426 31578
rect 4438 31526 4490 31578
rect 34966 31526 35018 31578
rect 35030 31526 35082 31578
rect 35094 31526 35146 31578
rect 35158 31526 35210 31578
rect 1676 31467 1728 31476
rect 1676 31433 1685 31467
rect 1685 31433 1719 31467
rect 1719 31433 1728 31467
rect 1676 31424 1728 31433
rect 4804 31424 4856 31476
rect 5632 31424 5684 31476
rect 6736 31424 6788 31476
rect 13084 31424 13136 31476
rect 2872 31331 2924 31340
rect 2872 31297 2881 31331
rect 2881 31297 2915 31331
rect 2915 31297 2924 31331
rect 2872 31288 2924 31297
rect 12256 31356 12308 31408
rect 1584 31263 1636 31272
rect 1584 31229 1593 31263
rect 1593 31229 1627 31263
rect 1627 31229 1636 31263
rect 1584 31220 1636 31229
rect 2504 31263 2556 31272
rect 2504 31229 2513 31263
rect 2513 31229 2547 31263
rect 2547 31229 2556 31263
rect 2504 31220 2556 31229
rect 2780 31220 2832 31272
rect 3056 31220 3108 31272
rect 3332 31220 3384 31272
rect 4068 31220 4120 31272
rect 4988 31263 5040 31272
rect 4988 31229 4997 31263
rect 4997 31229 5031 31263
rect 5031 31229 5040 31263
rect 4988 31220 5040 31229
rect 5356 31263 5408 31272
rect 5356 31229 5365 31263
rect 5365 31229 5399 31263
rect 5399 31229 5408 31263
rect 5356 31220 5408 31229
rect 6828 31263 6880 31272
rect 6828 31229 6837 31263
rect 6837 31229 6871 31263
rect 6871 31229 6880 31263
rect 6828 31220 6880 31229
rect 7748 31263 7800 31272
rect 7748 31229 7757 31263
rect 7757 31229 7791 31263
rect 7791 31229 7800 31263
rect 7748 31220 7800 31229
rect 11520 31288 11572 31340
rect 12440 31288 12492 31340
rect 13820 31288 13872 31340
rect 14556 31424 14608 31476
rect 15384 31424 15436 31476
rect 19892 31424 19944 31476
rect 20628 31424 20680 31476
rect 22376 31356 22428 31408
rect 15200 31288 15252 31340
rect 21640 31288 21692 31340
rect 21732 31288 21784 31340
rect 23296 31288 23348 31340
rect 26332 31356 26384 31408
rect 4804 31152 4856 31204
rect 9220 31152 9272 31204
rect 10692 31220 10744 31272
rect 11152 31220 11204 31272
rect 11520 31152 11572 31204
rect 11704 31220 11756 31272
rect 14188 31263 14240 31272
rect 12716 31152 12768 31204
rect 14188 31229 14197 31263
rect 14197 31229 14231 31263
rect 14231 31229 14240 31263
rect 14188 31220 14240 31229
rect 14004 31152 14056 31204
rect 15384 31220 15436 31272
rect 17316 31263 17368 31272
rect 17316 31229 17325 31263
rect 17325 31229 17359 31263
rect 17359 31229 17368 31263
rect 17316 31220 17368 31229
rect 18880 31220 18932 31272
rect 19340 31263 19392 31272
rect 19340 31229 19349 31263
rect 19349 31229 19383 31263
rect 19383 31229 19392 31263
rect 19800 31263 19852 31272
rect 19340 31220 19392 31229
rect 19800 31229 19809 31263
rect 19809 31229 19843 31263
rect 19843 31229 19852 31263
rect 19800 31220 19852 31229
rect 19892 31220 19944 31272
rect 20352 31263 20404 31272
rect 20352 31229 20361 31263
rect 20361 31229 20395 31263
rect 20395 31229 20404 31263
rect 20352 31220 20404 31229
rect 21088 31263 21140 31272
rect 21088 31229 21097 31263
rect 21097 31229 21131 31263
rect 21131 31229 21140 31263
rect 21088 31220 21140 31229
rect 20168 31152 20220 31204
rect 23572 31220 23624 31272
rect 23112 31152 23164 31204
rect 4896 31084 4948 31136
rect 5448 31084 5500 31136
rect 6920 31127 6972 31136
rect 6920 31093 6929 31127
rect 6929 31093 6963 31127
rect 6963 31093 6972 31127
rect 6920 31084 6972 31093
rect 11888 31127 11940 31136
rect 11888 31093 11897 31127
rect 11897 31093 11931 31127
rect 11931 31093 11940 31127
rect 11888 31084 11940 31093
rect 14372 31084 14424 31136
rect 16396 31127 16448 31136
rect 16396 31093 16405 31127
rect 16405 31093 16439 31127
rect 16439 31093 16448 31127
rect 16396 31084 16448 31093
rect 22008 31084 22060 31136
rect 22468 31084 22520 31136
rect 23572 31084 23624 31136
rect 23756 31220 23808 31272
rect 25136 31220 25188 31272
rect 25780 31263 25832 31272
rect 25780 31229 25789 31263
rect 25789 31229 25823 31263
rect 25823 31229 25832 31263
rect 25780 31220 25832 31229
rect 26516 31263 26568 31272
rect 26516 31229 26525 31263
rect 26525 31229 26559 31263
rect 26559 31229 26568 31263
rect 26516 31220 26568 31229
rect 26700 31263 26752 31272
rect 26700 31229 26709 31263
rect 26709 31229 26743 31263
rect 26743 31229 26752 31263
rect 26700 31220 26752 31229
rect 27160 31263 27212 31272
rect 27160 31229 27169 31263
rect 27169 31229 27203 31263
rect 27203 31229 27212 31263
rect 27160 31220 27212 31229
rect 27252 31263 27304 31272
rect 27252 31229 27261 31263
rect 27261 31229 27295 31263
rect 27295 31229 27304 31263
rect 29736 31331 29788 31340
rect 29736 31297 29745 31331
rect 29745 31297 29779 31331
rect 29779 31297 29788 31331
rect 29736 31288 29788 31297
rect 31760 31331 31812 31340
rect 31760 31297 31769 31331
rect 31769 31297 31803 31331
rect 31803 31297 31812 31331
rect 31760 31288 31812 31297
rect 32220 31356 32272 31408
rect 27252 31220 27304 31229
rect 25688 31152 25740 31204
rect 32036 31220 32088 31272
rect 33416 31263 33468 31272
rect 33416 31229 33425 31263
rect 33425 31229 33459 31263
rect 33459 31229 33468 31263
rect 33416 31220 33468 31229
rect 34520 31288 34572 31340
rect 35808 31424 35860 31476
rect 35716 31288 35768 31340
rect 35164 31220 35216 31272
rect 35992 31263 36044 31272
rect 35992 31229 36001 31263
rect 36001 31229 36035 31263
rect 36035 31229 36044 31263
rect 35992 31220 36044 31229
rect 36452 31263 36504 31272
rect 36452 31229 36461 31263
rect 36461 31229 36495 31263
rect 36495 31229 36504 31263
rect 36452 31220 36504 31229
rect 36636 31220 36688 31272
rect 36820 31263 36872 31272
rect 36820 31229 36829 31263
rect 36829 31229 36863 31263
rect 36863 31229 36872 31263
rect 36820 31220 36872 31229
rect 37740 31263 37792 31272
rect 32680 31152 32732 31204
rect 35440 31152 35492 31204
rect 35532 31152 35584 31204
rect 37740 31229 37749 31263
rect 37749 31229 37783 31263
rect 37783 31229 37792 31263
rect 37740 31220 37792 31229
rect 27988 31084 28040 31136
rect 28448 31084 28500 31136
rect 29460 31084 29512 31136
rect 30380 31084 30432 31136
rect 38108 31084 38160 31136
rect 38568 31084 38620 31136
rect 19606 30982 19658 31034
rect 19670 30982 19722 31034
rect 19734 30982 19786 31034
rect 19798 30982 19850 31034
rect 2136 30812 2188 30864
rect 3332 30787 3384 30796
rect 3332 30753 3341 30787
rect 3341 30753 3375 30787
rect 3375 30753 3384 30787
rect 3332 30744 3384 30753
rect 3516 30787 3568 30796
rect 3516 30753 3525 30787
rect 3525 30753 3559 30787
rect 3559 30753 3568 30787
rect 3516 30744 3568 30753
rect 4896 30787 4948 30796
rect 4896 30753 4905 30787
rect 4905 30753 4939 30787
rect 4939 30753 4948 30787
rect 4896 30744 4948 30753
rect 6828 30880 6880 30932
rect 8760 30880 8812 30932
rect 11704 30880 11756 30932
rect 12532 30880 12584 30932
rect 7012 30744 7064 30796
rect 8944 30812 8996 30864
rect 8300 30744 8352 30796
rect 4712 30676 4764 30728
rect 5632 30719 5684 30728
rect 5632 30685 5641 30719
rect 5641 30685 5675 30719
rect 5675 30685 5684 30719
rect 5632 30676 5684 30685
rect 8484 30719 8536 30728
rect 8484 30685 8493 30719
rect 8493 30685 8527 30719
rect 8527 30685 8536 30719
rect 8484 30676 8536 30685
rect 9680 30787 9732 30796
rect 9680 30753 9689 30787
rect 9689 30753 9723 30787
rect 9723 30753 9732 30787
rect 9680 30744 9732 30753
rect 10692 30744 10744 30796
rect 11152 30787 11204 30796
rect 11152 30753 11161 30787
rect 11161 30753 11195 30787
rect 11195 30753 11204 30787
rect 11152 30744 11204 30753
rect 11520 30787 11572 30796
rect 11520 30753 11529 30787
rect 11529 30753 11563 30787
rect 11563 30753 11572 30787
rect 11520 30744 11572 30753
rect 13728 30744 13780 30796
rect 14832 30812 14884 30864
rect 15292 30812 15344 30864
rect 14004 30787 14056 30796
rect 14004 30753 14013 30787
rect 14013 30753 14047 30787
rect 14047 30753 14056 30787
rect 14004 30744 14056 30753
rect 17868 30812 17920 30864
rect 16120 30787 16172 30796
rect 10968 30676 11020 30728
rect 12808 30676 12860 30728
rect 15384 30676 15436 30728
rect 16120 30753 16129 30787
rect 16129 30753 16163 30787
rect 16163 30753 16172 30787
rect 16120 30744 16172 30753
rect 17132 30744 17184 30796
rect 17224 30787 17276 30796
rect 17224 30753 17233 30787
rect 17233 30753 17267 30787
rect 17267 30753 17276 30787
rect 17592 30787 17644 30796
rect 17224 30744 17276 30753
rect 17592 30753 17601 30787
rect 17601 30753 17635 30787
rect 17635 30753 17644 30787
rect 17592 30744 17644 30753
rect 17684 30744 17736 30796
rect 18880 30744 18932 30796
rect 20260 30880 20312 30932
rect 21732 30880 21784 30932
rect 26148 30812 26200 30864
rect 29644 30855 29696 30864
rect 29644 30821 29653 30855
rect 29653 30821 29687 30855
rect 29687 30821 29696 30855
rect 29644 30812 29696 30821
rect 21640 30787 21692 30796
rect 5540 30608 5592 30660
rect 8760 30608 8812 30660
rect 15108 30608 15160 30660
rect 16396 30676 16448 30728
rect 21640 30753 21649 30787
rect 21649 30753 21683 30787
rect 21683 30753 21692 30787
rect 21640 30744 21692 30753
rect 22376 30787 22428 30796
rect 22376 30753 22385 30787
rect 22385 30753 22419 30787
rect 22419 30753 22428 30787
rect 22376 30744 22428 30753
rect 23572 30744 23624 30796
rect 24216 30787 24268 30796
rect 24216 30753 24225 30787
rect 24225 30753 24259 30787
rect 24259 30753 24268 30787
rect 24216 30744 24268 30753
rect 25228 30787 25280 30796
rect 25228 30753 25237 30787
rect 25237 30753 25271 30787
rect 25271 30753 25280 30787
rect 25228 30744 25280 30753
rect 25412 30744 25464 30796
rect 25780 30787 25832 30796
rect 25780 30753 25789 30787
rect 25789 30753 25823 30787
rect 25823 30753 25832 30787
rect 25780 30744 25832 30753
rect 27068 30787 27120 30796
rect 27068 30753 27077 30787
rect 27077 30753 27111 30787
rect 27111 30753 27120 30787
rect 27068 30744 27120 30753
rect 20352 30676 20404 30728
rect 22284 30676 22336 30728
rect 28632 30744 28684 30796
rect 33416 30880 33468 30932
rect 35256 30880 35308 30932
rect 36820 30880 36872 30932
rect 37740 30880 37792 30932
rect 36268 30812 36320 30864
rect 18236 30608 18288 30660
rect 19984 30651 20036 30660
rect 19984 30617 19993 30651
rect 19993 30617 20027 30651
rect 20027 30617 20036 30651
rect 19984 30608 20036 30617
rect 22100 30608 22152 30660
rect 27620 30676 27672 30728
rect 27252 30608 27304 30660
rect 29736 30676 29788 30728
rect 30564 30719 30616 30728
rect 30564 30685 30573 30719
rect 30573 30685 30607 30719
rect 30607 30685 30616 30719
rect 30564 30676 30616 30685
rect 32956 30787 33008 30796
rect 31116 30676 31168 30728
rect 9312 30583 9364 30592
rect 9312 30549 9321 30583
rect 9321 30549 9355 30583
rect 9355 30549 9364 30583
rect 9312 30540 9364 30549
rect 15292 30540 15344 30592
rect 29000 30540 29052 30592
rect 29184 30540 29236 30592
rect 30748 30540 30800 30592
rect 32680 30719 32732 30728
rect 32680 30685 32689 30719
rect 32689 30685 32723 30719
rect 32723 30685 32732 30719
rect 32680 30676 32732 30685
rect 32956 30753 32965 30787
rect 32965 30753 32999 30787
rect 32999 30753 33008 30787
rect 32956 30744 33008 30753
rect 35348 30744 35400 30796
rect 35716 30787 35768 30796
rect 35716 30753 35725 30787
rect 35725 30753 35759 30787
rect 35759 30753 35768 30787
rect 35716 30744 35768 30753
rect 36452 30744 36504 30796
rect 36912 30744 36964 30796
rect 38476 30787 38528 30796
rect 38476 30753 38485 30787
rect 38485 30753 38519 30787
rect 38519 30753 38528 30787
rect 38476 30744 38528 30753
rect 34796 30676 34848 30728
rect 36360 30676 36412 30728
rect 37648 30676 37700 30728
rect 37832 30676 37884 30728
rect 32036 30540 32088 30592
rect 4246 30438 4298 30490
rect 4310 30438 4362 30490
rect 4374 30438 4426 30490
rect 4438 30438 4490 30490
rect 34966 30438 35018 30490
rect 35030 30438 35082 30490
rect 35094 30438 35146 30490
rect 35158 30438 35210 30490
rect 1768 30200 1820 30252
rect 7748 30336 7800 30388
rect 4068 30268 4120 30320
rect 2780 30175 2832 30184
rect 2780 30141 2789 30175
rect 2789 30141 2823 30175
rect 2823 30141 2832 30175
rect 2964 30175 3016 30184
rect 2780 30132 2832 30141
rect 2964 30141 2973 30175
rect 2973 30141 3007 30175
rect 3007 30141 3016 30175
rect 2964 30132 3016 30141
rect 3240 30175 3292 30184
rect 3240 30141 3249 30175
rect 3249 30141 3283 30175
rect 3283 30141 3292 30175
rect 3240 30132 3292 30141
rect 3424 30175 3476 30184
rect 3424 30141 3433 30175
rect 3433 30141 3467 30175
rect 3467 30141 3476 30175
rect 3424 30132 3476 30141
rect 3516 30132 3568 30184
rect 5816 30268 5868 30320
rect 7564 30268 7616 30320
rect 8484 30336 8536 30388
rect 8944 30379 8996 30388
rect 8944 30345 8953 30379
rect 8953 30345 8987 30379
rect 8987 30345 8996 30379
rect 8944 30336 8996 30345
rect 19524 30336 19576 30388
rect 20260 30336 20312 30388
rect 4988 30175 5040 30184
rect 1492 30064 1544 30116
rect 4988 30141 4997 30175
rect 4997 30141 5031 30175
rect 5031 30141 5040 30175
rect 4988 30132 5040 30141
rect 5356 30132 5408 30184
rect 11152 30268 11204 30320
rect 23756 30336 23808 30388
rect 25504 30336 25556 30388
rect 33048 30336 33100 30388
rect 34520 30336 34572 30388
rect 24216 30268 24268 30320
rect 31944 30311 31996 30320
rect 10508 30243 10560 30252
rect 10508 30209 10517 30243
rect 10517 30209 10551 30243
rect 10551 30209 10560 30243
rect 10508 30200 10560 30209
rect 12716 30243 12768 30252
rect 12716 30209 12725 30243
rect 12725 30209 12759 30243
rect 12759 30209 12768 30243
rect 12716 30200 12768 30209
rect 14372 30200 14424 30252
rect 16120 30200 16172 30252
rect 18512 30200 18564 30252
rect 24492 30243 24544 30252
rect 4712 30064 4764 30116
rect 3884 29996 3936 30048
rect 7840 30064 7892 30116
rect 9036 30175 9088 30184
rect 9036 30141 9045 30175
rect 9045 30141 9079 30175
rect 9079 30141 9088 30175
rect 9220 30175 9272 30184
rect 9036 30132 9088 30141
rect 9220 30141 9229 30175
rect 9229 30141 9263 30175
rect 9263 30141 9272 30175
rect 9220 30132 9272 30141
rect 10876 30132 10928 30184
rect 11060 30132 11112 30184
rect 11796 30132 11848 30184
rect 13084 30132 13136 30184
rect 14464 30132 14516 30184
rect 14832 30107 14884 30116
rect 14832 30073 14841 30107
rect 14841 30073 14875 30107
rect 14875 30073 14884 30107
rect 14832 30064 14884 30073
rect 7656 29996 7708 30048
rect 14188 29996 14240 30048
rect 15200 29996 15252 30048
rect 15568 29996 15620 30048
rect 19156 30132 19208 30184
rect 19524 30175 19576 30184
rect 19524 30141 19533 30175
rect 19533 30141 19567 30175
rect 19567 30141 19576 30175
rect 19524 30132 19576 30141
rect 19800 30175 19852 30184
rect 19800 30141 19809 30175
rect 19809 30141 19843 30175
rect 19843 30141 19852 30175
rect 19800 30132 19852 30141
rect 19892 30132 19944 30184
rect 20536 30175 20588 30184
rect 20536 30141 20545 30175
rect 20545 30141 20579 30175
rect 20579 30141 20588 30175
rect 20536 30132 20588 30141
rect 21088 30132 21140 30184
rect 21640 30132 21692 30184
rect 19340 30064 19392 30116
rect 22100 30175 22152 30184
rect 22100 30141 22109 30175
rect 22109 30141 22143 30175
rect 22143 30141 22152 30175
rect 24492 30209 24501 30243
rect 24501 30209 24535 30243
rect 24535 30209 24544 30243
rect 24492 30200 24544 30209
rect 25320 30200 25372 30252
rect 25504 30200 25556 30252
rect 26332 30243 26384 30252
rect 26332 30209 26341 30243
rect 26341 30209 26375 30243
rect 26375 30209 26384 30243
rect 26332 30200 26384 30209
rect 22100 30132 22152 30141
rect 21824 30064 21876 30116
rect 23848 30132 23900 30184
rect 24308 30132 24360 30184
rect 26056 30175 26108 30184
rect 26056 30141 26065 30175
rect 26065 30141 26099 30175
rect 26099 30141 26108 30175
rect 26056 30132 26108 30141
rect 26424 30175 26476 30184
rect 26424 30141 26433 30175
rect 26433 30141 26467 30175
rect 26467 30141 26476 30175
rect 26424 30132 26476 30141
rect 31944 30277 31953 30311
rect 31953 30277 31987 30311
rect 31987 30277 31996 30311
rect 31944 30268 31996 30277
rect 32036 30268 32088 30320
rect 34152 30268 34204 30320
rect 36912 30268 36964 30320
rect 30288 30200 30340 30252
rect 30564 30243 30616 30252
rect 30564 30209 30573 30243
rect 30573 30209 30607 30243
rect 30607 30209 30616 30243
rect 30564 30200 30616 30209
rect 30748 30200 30800 30252
rect 37464 30243 37516 30252
rect 28540 30132 28592 30184
rect 29828 30175 29880 30184
rect 29828 30141 29837 30175
rect 29837 30141 29871 30175
rect 29871 30141 29880 30175
rect 29828 30132 29880 30141
rect 30104 30132 30156 30184
rect 31208 30175 31260 30184
rect 31208 30141 31217 30175
rect 31217 30141 31251 30175
rect 31251 30141 31260 30175
rect 31208 30132 31260 30141
rect 29644 30064 29696 30116
rect 30472 30064 30524 30116
rect 37464 30209 37473 30243
rect 37473 30209 37507 30243
rect 37507 30209 37516 30243
rect 37464 30200 37516 30209
rect 39120 30243 39172 30252
rect 39120 30209 39129 30243
rect 39129 30209 39163 30243
rect 39163 30209 39172 30243
rect 39120 30200 39172 30209
rect 33324 30132 33376 30184
rect 33508 30175 33560 30184
rect 33508 30141 33517 30175
rect 33517 30141 33551 30175
rect 33551 30141 33560 30175
rect 33508 30132 33560 30141
rect 34428 30132 34480 30184
rect 34520 30132 34572 30184
rect 35624 30132 35676 30184
rect 35808 30175 35860 30184
rect 35808 30141 35817 30175
rect 35817 30141 35851 30175
rect 35851 30141 35860 30175
rect 35808 30132 35860 30141
rect 36912 30132 36964 30184
rect 37372 30132 37424 30184
rect 36452 30107 36504 30116
rect 36452 30073 36461 30107
rect 36461 30073 36495 30107
rect 36495 30073 36504 30107
rect 36452 30064 36504 30073
rect 27160 30039 27212 30048
rect 27160 30005 27169 30039
rect 27169 30005 27203 30039
rect 27203 30005 27212 30039
rect 27160 29996 27212 30005
rect 27712 30039 27764 30048
rect 27712 30005 27721 30039
rect 27721 30005 27755 30039
rect 27755 30005 27764 30039
rect 27712 29996 27764 30005
rect 28448 29996 28500 30048
rect 30012 30039 30064 30048
rect 30012 30005 30021 30039
rect 30021 30005 30055 30039
rect 30055 30005 30064 30039
rect 30012 29996 30064 30005
rect 30104 30039 30156 30048
rect 30104 30005 30113 30039
rect 30113 30005 30147 30039
rect 30147 30005 30156 30039
rect 30104 29996 30156 30005
rect 32680 29996 32732 30048
rect 33048 29996 33100 30048
rect 38568 29996 38620 30048
rect 19606 29894 19658 29946
rect 19670 29894 19722 29946
rect 19734 29894 19786 29946
rect 19798 29894 19850 29946
rect 2780 29835 2832 29844
rect 2780 29801 2789 29835
rect 2789 29801 2823 29835
rect 2823 29801 2832 29835
rect 2780 29792 2832 29801
rect 3516 29792 3568 29844
rect 5448 29792 5500 29844
rect 5540 29792 5592 29844
rect 3148 29724 3200 29776
rect 3424 29724 3476 29776
rect 5356 29724 5408 29776
rect 1400 29699 1452 29708
rect 1400 29665 1409 29699
rect 1409 29665 1443 29699
rect 1443 29665 1452 29699
rect 1400 29656 1452 29665
rect 2872 29656 2924 29708
rect 6920 29724 6972 29776
rect 8300 29724 8352 29776
rect 6000 29699 6052 29708
rect 1676 29631 1728 29640
rect 1676 29597 1685 29631
rect 1685 29597 1719 29631
rect 1719 29597 1728 29631
rect 1676 29588 1728 29597
rect 5448 29588 5500 29640
rect 6000 29665 6009 29699
rect 6009 29665 6043 29699
rect 6043 29665 6052 29699
rect 6000 29656 6052 29665
rect 7012 29656 7064 29708
rect 4804 29520 4856 29572
rect 8760 29656 8812 29708
rect 8944 29699 8996 29708
rect 8944 29665 8953 29699
rect 8953 29665 8987 29699
rect 8987 29665 8996 29699
rect 8944 29656 8996 29665
rect 9404 29656 9456 29708
rect 11428 29724 11480 29776
rect 10232 29656 10284 29708
rect 10508 29699 10560 29708
rect 10508 29665 10517 29699
rect 10517 29665 10551 29699
rect 10551 29665 10560 29699
rect 10508 29656 10560 29665
rect 10692 29699 10744 29708
rect 10692 29665 10701 29699
rect 10701 29665 10735 29699
rect 10735 29665 10744 29699
rect 10692 29656 10744 29665
rect 11244 29699 11296 29708
rect 11244 29665 11253 29699
rect 11253 29665 11287 29699
rect 11287 29665 11296 29699
rect 11244 29656 11296 29665
rect 11796 29699 11848 29708
rect 11796 29665 11805 29699
rect 11805 29665 11839 29699
rect 11839 29665 11848 29699
rect 11796 29656 11848 29665
rect 12624 29724 12676 29776
rect 12440 29656 12492 29708
rect 13728 29656 13780 29708
rect 14280 29699 14332 29708
rect 14280 29665 14289 29699
rect 14289 29665 14323 29699
rect 14323 29665 14332 29699
rect 14280 29656 14332 29665
rect 15292 29699 15344 29708
rect 15292 29665 15301 29699
rect 15301 29665 15335 29699
rect 15335 29665 15344 29699
rect 15292 29656 15344 29665
rect 15384 29656 15436 29708
rect 15936 29656 15988 29708
rect 17592 29656 17644 29708
rect 18236 29699 18288 29708
rect 18236 29665 18245 29699
rect 18245 29665 18279 29699
rect 18279 29665 18288 29699
rect 18236 29656 18288 29665
rect 19984 29724 20036 29776
rect 19064 29699 19116 29708
rect 19064 29665 19073 29699
rect 19073 29665 19107 29699
rect 19107 29665 19116 29699
rect 19064 29656 19116 29665
rect 19800 29699 19852 29708
rect 19800 29665 19809 29699
rect 19809 29665 19843 29699
rect 19843 29665 19852 29699
rect 19800 29656 19852 29665
rect 9220 29588 9272 29640
rect 13544 29588 13596 29640
rect 15660 29631 15712 29640
rect 15660 29597 15669 29631
rect 15669 29597 15703 29631
rect 15703 29597 15712 29631
rect 15660 29588 15712 29597
rect 11336 29563 11388 29572
rect 11336 29529 11345 29563
rect 11345 29529 11379 29563
rect 11379 29529 11388 29563
rect 11336 29520 11388 29529
rect 12900 29563 12952 29572
rect 12900 29529 12909 29563
rect 12909 29529 12943 29563
rect 12943 29529 12952 29563
rect 12900 29520 12952 29529
rect 13636 29520 13688 29572
rect 19616 29588 19668 29640
rect 20536 29724 20588 29776
rect 21180 29724 21232 29776
rect 21824 29724 21876 29776
rect 24492 29724 24544 29776
rect 25320 29724 25372 29776
rect 20720 29656 20772 29708
rect 20904 29699 20956 29708
rect 20904 29665 20913 29699
rect 20913 29665 20947 29699
rect 20947 29665 20956 29699
rect 20904 29656 20956 29665
rect 21088 29656 21140 29708
rect 21548 29656 21600 29708
rect 22560 29699 22612 29708
rect 22560 29665 22569 29699
rect 22569 29665 22603 29699
rect 22603 29665 22612 29699
rect 22560 29656 22612 29665
rect 22928 29699 22980 29708
rect 22928 29665 22937 29699
rect 22937 29665 22971 29699
rect 22971 29665 22980 29699
rect 22928 29656 22980 29665
rect 23204 29699 23256 29708
rect 23204 29665 23213 29699
rect 23213 29665 23247 29699
rect 23247 29665 23256 29699
rect 23204 29656 23256 29665
rect 24400 29656 24452 29708
rect 18420 29563 18472 29572
rect 18420 29529 18429 29563
rect 18429 29529 18463 29563
rect 18463 29529 18472 29563
rect 18420 29520 18472 29529
rect 18788 29520 18840 29572
rect 4620 29452 4672 29504
rect 7472 29495 7524 29504
rect 7472 29461 7481 29495
rect 7481 29461 7515 29495
rect 7515 29461 7524 29495
rect 7472 29452 7524 29461
rect 15200 29452 15252 29504
rect 20996 29588 21048 29640
rect 25504 29699 25556 29708
rect 25504 29665 25513 29699
rect 25513 29665 25547 29699
rect 25547 29665 25556 29699
rect 25504 29656 25556 29665
rect 26608 29656 26660 29708
rect 27620 29699 27672 29708
rect 20168 29520 20220 29572
rect 23296 29563 23348 29572
rect 23296 29529 23305 29563
rect 23305 29529 23339 29563
rect 23339 29529 23348 29563
rect 23296 29520 23348 29529
rect 24216 29563 24268 29572
rect 24216 29529 24225 29563
rect 24225 29529 24259 29563
rect 24259 29529 24268 29563
rect 24216 29520 24268 29529
rect 26700 29588 26752 29640
rect 27252 29588 27304 29640
rect 27620 29665 27629 29699
rect 27629 29665 27663 29699
rect 27663 29665 27672 29699
rect 27620 29656 27672 29665
rect 28908 29656 28960 29708
rect 30104 29792 30156 29844
rect 30472 29792 30524 29844
rect 30656 29792 30708 29844
rect 31300 29792 31352 29844
rect 36268 29792 36320 29844
rect 29644 29724 29696 29776
rect 30840 29767 30892 29776
rect 30840 29733 30849 29767
rect 30849 29733 30883 29767
rect 30883 29733 30892 29767
rect 30840 29724 30892 29733
rect 31208 29767 31260 29776
rect 31208 29733 31217 29767
rect 31217 29733 31251 29767
rect 31251 29733 31260 29767
rect 31208 29724 31260 29733
rect 36636 29724 36688 29776
rect 30012 29656 30064 29708
rect 31024 29656 31076 29708
rect 29828 29588 29880 29640
rect 25688 29563 25740 29572
rect 25688 29529 25697 29563
rect 25697 29529 25731 29563
rect 25731 29529 25740 29563
rect 25688 29520 25740 29529
rect 26516 29452 26568 29504
rect 27804 29452 27856 29504
rect 28540 29452 28592 29504
rect 29368 29452 29420 29504
rect 29736 29495 29788 29504
rect 29736 29461 29745 29495
rect 29745 29461 29779 29495
rect 29779 29461 29788 29495
rect 29736 29452 29788 29461
rect 33048 29656 33100 29708
rect 35532 29699 35584 29708
rect 35532 29665 35541 29699
rect 35541 29665 35575 29699
rect 35575 29665 35584 29699
rect 35532 29656 35584 29665
rect 37740 29699 37792 29708
rect 37740 29665 37749 29699
rect 37749 29665 37783 29699
rect 37783 29665 37792 29699
rect 37740 29656 37792 29665
rect 37924 29656 37976 29708
rect 38568 29699 38620 29708
rect 38568 29665 38577 29699
rect 38577 29665 38611 29699
rect 38611 29665 38620 29699
rect 38568 29656 38620 29665
rect 33232 29631 33284 29640
rect 33232 29597 33241 29631
rect 33241 29597 33275 29631
rect 33275 29597 33284 29631
rect 33232 29588 33284 29597
rect 35716 29588 35768 29640
rect 34428 29520 34480 29572
rect 34520 29495 34572 29504
rect 34520 29461 34529 29495
rect 34529 29461 34563 29495
rect 34563 29461 34572 29495
rect 34520 29452 34572 29461
rect 36176 29452 36228 29504
rect 36912 29495 36964 29504
rect 36912 29461 36921 29495
rect 36921 29461 36955 29495
rect 36955 29461 36964 29495
rect 36912 29452 36964 29461
rect 4246 29350 4298 29402
rect 4310 29350 4362 29402
rect 4374 29350 4426 29402
rect 4438 29350 4490 29402
rect 34966 29350 35018 29402
rect 35030 29350 35082 29402
rect 35094 29350 35146 29402
rect 35158 29350 35210 29402
rect 1492 29291 1544 29300
rect 1492 29257 1501 29291
rect 1501 29257 1535 29291
rect 1535 29257 1544 29291
rect 1492 29248 1544 29257
rect 1676 29248 1728 29300
rect 5356 29248 5408 29300
rect 10876 29248 10928 29300
rect 11244 29248 11296 29300
rect 11428 29291 11480 29300
rect 11428 29257 11437 29291
rect 11437 29257 11471 29291
rect 11471 29257 11480 29291
rect 11428 29248 11480 29257
rect 11796 29248 11848 29300
rect 14280 29248 14332 29300
rect 17592 29248 17644 29300
rect 18328 29248 18380 29300
rect 20996 29248 21048 29300
rect 23204 29248 23256 29300
rect 25320 29248 25372 29300
rect 26332 29248 26384 29300
rect 1860 29112 1912 29164
rect 1768 29087 1820 29096
rect 1768 29053 1777 29087
rect 1777 29053 1811 29087
rect 1811 29053 1820 29087
rect 1768 29044 1820 29053
rect 3148 29112 3200 29164
rect 3332 29112 3384 29164
rect 9220 29180 9272 29232
rect 4988 29112 5040 29164
rect 5724 29155 5776 29164
rect 5724 29121 5733 29155
rect 5733 29121 5767 29155
rect 5767 29121 5776 29155
rect 5724 29112 5776 29121
rect 3516 29044 3568 29096
rect 5264 29087 5316 29096
rect 2044 28976 2096 29028
rect 2780 28976 2832 29028
rect 4620 28976 4672 29028
rect 5264 29053 5273 29087
rect 5273 29053 5307 29087
rect 5307 29053 5316 29087
rect 5264 29044 5316 29053
rect 5816 29044 5868 29096
rect 7472 29112 7524 29164
rect 7012 29044 7064 29096
rect 8300 29044 8352 29096
rect 8484 29112 8536 29164
rect 12440 29112 12492 29164
rect 9312 29044 9364 29096
rect 9956 29087 10008 29096
rect 9956 29053 9965 29087
rect 9965 29053 9999 29087
rect 9999 29053 10008 29087
rect 9956 29044 10008 29053
rect 10140 29087 10192 29096
rect 10140 29053 10149 29087
rect 10149 29053 10183 29087
rect 10183 29053 10192 29087
rect 10140 29044 10192 29053
rect 10416 29087 10468 29096
rect 10416 29053 10425 29087
rect 10425 29053 10459 29087
rect 10459 29053 10468 29087
rect 10416 29044 10468 29053
rect 5632 28976 5684 29028
rect 6000 28976 6052 29028
rect 9036 28976 9088 29028
rect 13360 29044 13412 29096
rect 13544 29087 13596 29096
rect 13544 29053 13553 29087
rect 13553 29053 13587 29087
rect 13587 29053 13596 29087
rect 13544 29044 13596 29053
rect 13728 29087 13780 29096
rect 13728 29053 13737 29087
rect 13737 29053 13771 29087
rect 13771 29053 13780 29087
rect 13728 29044 13780 29053
rect 14280 29087 14332 29096
rect 14280 29053 14289 29087
rect 14289 29053 14323 29087
rect 14323 29053 14332 29087
rect 14280 29044 14332 29053
rect 14648 29044 14700 29096
rect 17316 29180 17368 29232
rect 18788 29180 18840 29232
rect 15660 29044 15712 29096
rect 15936 29044 15988 29096
rect 16396 29044 16448 29096
rect 16948 29044 17000 29096
rect 17224 29087 17276 29096
rect 17224 29053 17233 29087
rect 17233 29053 17267 29087
rect 17267 29053 17276 29087
rect 17224 29044 17276 29053
rect 17960 29044 18012 29096
rect 18420 29087 18472 29096
rect 18420 29053 18429 29087
rect 18429 29053 18463 29087
rect 18463 29053 18472 29087
rect 18420 29044 18472 29053
rect 14556 28976 14608 29028
rect 17500 28976 17552 29028
rect 19432 29044 19484 29096
rect 23940 29180 23992 29232
rect 24400 29223 24452 29232
rect 24400 29189 24409 29223
rect 24409 29189 24443 29223
rect 24443 29189 24452 29223
rect 24400 29180 24452 29189
rect 20536 29044 20588 29096
rect 21364 29044 21416 29096
rect 21824 29087 21876 29096
rect 21824 29053 21833 29087
rect 21833 29053 21867 29087
rect 21867 29053 21876 29087
rect 21824 29044 21876 29053
rect 22008 29044 22060 29096
rect 22836 29044 22888 29096
rect 23848 29044 23900 29096
rect 24032 29044 24084 29096
rect 24492 29087 24544 29096
rect 24492 29053 24501 29087
rect 24501 29053 24535 29087
rect 24535 29053 24544 29087
rect 24492 29044 24544 29053
rect 24584 29044 24636 29096
rect 24952 28976 25004 29028
rect 9864 28908 9916 28960
rect 10140 28908 10192 28960
rect 20260 28908 20312 28960
rect 22836 28908 22888 28960
rect 25964 29044 26016 29096
rect 26056 29087 26108 29096
rect 26056 29053 26065 29087
rect 26065 29053 26099 29087
rect 26099 29053 26108 29087
rect 26056 29044 26108 29053
rect 26608 29087 26660 29096
rect 26608 29053 26617 29087
rect 26617 29053 26651 29087
rect 26651 29053 26660 29087
rect 26608 29044 26660 29053
rect 26976 29112 27028 29164
rect 30012 29248 30064 29300
rect 36452 29248 36504 29300
rect 28172 29180 28224 29232
rect 29000 29180 29052 29232
rect 30288 29180 30340 29232
rect 33232 29180 33284 29232
rect 35716 29223 35768 29232
rect 35716 29189 35725 29223
rect 35725 29189 35759 29223
rect 35759 29189 35768 29223
rect 35716 29180 35768 29189
rect 37556 29180 37608 29232
rect 36452 29155 36504 29164
rect 27804 29044 27856 29096
rect 28172 29087 28224 29096
rect 28172 29053 28181 29087
rect 28181 29053 28215 29087
rect 28215 29053 28224 29087
rect 28172 29044 28224 29053
rect 29092 29044 29144 29096
rect 29184 29044 29236 29096
rect 29552 29087 29604 29096
rect 29552 29053 29561 29087
rect 29561 29053 29595 29087
rect 29595 29053 29604 29087
rect 29552 29044 29604 29053
rect 32036 29044 32088 29096
rect 36452 29121 36461 29155
rect 36461 29121 36495 29155
rect 36495 29121 36504 29155
rect 36452 29112 36504 29121
rect 34152 29044 34204 29096
rect 35440 29087 35492 29096
rect 35440 29053 35449 29087
rect 35449 29053 35483 29087
rect 35483 29053 35492 29087
rect 35440 29044 35492 29053
rect 36176 29087 36228 29096
rect 36176 29053 36185 29087
rect 36185 29053 36219 29087
rect 36219 29053 36228 29087
rect 36176 29044 36228 29053
rect 36360 29044 36412 29096
rect 34520 28976 34572 29028
rect 37832 29087 37884 29096
rect 37832 29053 37841 29087
rect 37841 29053 37875 29087
rect 37875 29053 37884 29087
rect 37832 29044 37884 29053
rect 38476 29044 38528 29096
rect 38660 28976 38712 29028
rect 25964 28908 26016 28960
rect 26240 28908 26292 28960
rect 33140 28908 33192 28960
rect 19606 28806 19658 28858
rect 19670 28806 19722 28858
rect 19734 28806 19786 28858
rect 19798 28806 19850 28858
rect 2872 28704 2924 28756
rect 3240 28747 3292 28756
rect 3240 28713 3249 28747
rect 3249 28713 3283 28747
rect 3283 28713 3292 28747
rect 3240 28704 3292 28713
rect 4804 28747 4856 28756
rect 4804 28713 4813 28747
rect 4813 28713 4847 28747
rect 4847 28713 4856 28747
rect 4804 28704 4856 28713
rect 7012 28704 7064 28756
rect 8300 28747 8352 28756
rect 8300 28713 8309 28747
rect 8309 28713 8343 28747
rect 8343 28713 8352 28747
rect 8300 28704 8352 28713
rect 10416 28704 10468 28756
rect 13452 28704 13504 28756
rect 16672 28704 16724 28756
rect 17132 28704 17184 28756
rect 4620 28611 4672 28620
rect 4620 28577 4629 28611
rect 4629 28577 4663 28611
rect 4663 28577 4672 28611
rect 4620 28568 4672 28577
rect 5632 28636 5684 28688
rect 12440 28636 12492 28688
rect 17408 28636 17460 28688
rect 17960 28679 18012 28688
rect 17960 28645 17969 28679
rect 17969 28645 18003 28679
rect 18003 28645 18012 28679
rect 17960 28636 18012 28645
rect 19156 28704 19208 28756
rect 20260 28704 20312 28756
rect 21456 28704 21508 28756
rect 22468 28704 22520 28756
rect 5540 28568 5592 28620
rect 8484 28568 8536 28620
rect 8944 28611 8996 28620
rect 8944 28577 8953 28611
rect 8953 28577 8987 28611
rect 8987 28577 8996 28611
rect 8944 28568 8996 28577
rect 9128 28568 9180 28620
rect 11336 28568 11388 28620
rect 11520 28568 11572 28620
rect 15660 28611 15712 28620
rect 15660 28577 15669 28611
rect 15669 28577 15703 28611
rect 15703 28577 15712 28611
rect 15660 28568 15712 28577
rect 16396 28568 16448 28620
rect 16948 28611 17000 28620
rect 16948 28577 16957 28611
rect 16957 28577 16991 28611
rect 16991 28577 17000 28611
rect 16948 28568 17000 28577
rect 1400 28500 1452 28552
rect 4068 28500 4120 28552
rect 5448 28543 5500 28552
rect 5448 28509 5457 28543
rect 5457 28509 5491 28543
rect 5491 28509 5500 28543
rect 5448 28500 5500 28509
rect 6552 28500 6604 28552
rect 9312 28500 9364 28552
rect 13084 28543 13136 28552
rect 13084 28509 13093 28543
rect 13093 28509 13127 28543
rect 13127 28509 13136 28543
rect 13084 28500 13136 28509
rect 15200 28500 15252 28552
rect 16672 28432 16724 28484
rect 18236 28611 18288 28620
rect 18236 28577 18245 28611
rect 18245 28577 18279 28611
rect 18279 28577 18288 28611
rect 18236 28568 18288 28577
rect 18972 28568 19024 28620
rect 18328 28500 18380 28552
rect 19340 28568 19392 28620
rect 19432 28568 19484 28620
rect 7656 28364 7708 28416
rect 13360 28364 13412 28416
rect 13728 28364 13780 28416
rect 14648 28364 14700 28416
rect 20168 28500 20220 28552
rect 20996 28500 21048 28552
rect 21364 28568 21416 28620
rect 22100 28611 22152 28620
rect 22100 28577 22109 28611
rect 22109 28577 22143 28611
rect 22143 28577 22152 28611
rect 22100 28568 22152 28577
rect 22836 28611 22888 28620
rect 21824 28500 21876 28552
rect 22836 28577 22845 28611
rect 22845 28577 22879 28611
rect 22879 28577 22888 28611
rect 22836 28568 22888 28577
rect 23480 28611 23532 28620
rect 23480 28577 23489 28611
rect 23489 28577 23523 28611
rect 23523 28577 23532 28611
rect 23480 28568 23532 28577
rect 23756 28568 23808 28620
rect 24584 28568 24636 28620
rect 24952 28611 25004 28620
rect 24952 28577 24961 28611
rect 24961 28577 24995 28611
rect 24995 28577 25004 28611
rect 24952 28568 25004 28577
rect 22928 28500 22980 28552
rect 20720 28432 20772 28484
rect 24400 28500 24452 28552
rect 26516 28704 26568 28756
rect 29000 28704 29052 28756
rect 27620 28636 27672 28688
rect 26332 28568 26384 28620
rect 27712 28568 27764 28620
rect 28264 28611 28316 28620
rect 28264 28577 28273 28611
rect 28273 28577 28307 28611
rect 28307 28577 28316 28611
rect 28264 28568 28316 28577
rect 29092 28636 29144 28688
rect 32128 28636 32180 28688
rect 34428 28636 34480 28688
rect 36360 28679 36412 28688
rect 30288 28568 30340 28620
rect 26240 28500 26292 28552
rect 26608 28543 26660 28552
rect 26608 28509 26617 28543
rect 26617 28509 26651 28543
rect 26651 28509 26660 28543
rect 26608 28500 26660 28509
rect 26700 28500 26752 28552
rect 30472 28568 30524 28620
rect 31392 28611 31444 28620
rect 31392 28577 31401 28611
rect 31401 28577 31435 28611
rect 31435 28577 31444 28611
rect 31392 28568 31444 28577
rect 33048 28568 33100 28620
rect 30012 28432 30064 28484
rect 19616 28364 19668 28416
rect 22376 28364 22428 28416
rect 22836 28364 22888 28416
rect 24124 28364 24176 28416
rect 24768 28364 24820 28416
rect 26608 28364 26660 28416
rect 27436 28364 27488 28416
rect 27528 28364 27580 28416
rect 29092 28364 29144 28416
rect 34796 28568 34848 28620
rect 35716 28611 35768 28620
rect 35716 28577 35725 28611
rect 35725 28577 35759 28611
rect 35759 28577 35768 28611
rect 35716 28568 35768 28577
rect 35808 28568 35860 28620
rect 36360 28645 36369 28679
rect 36369 28645 36403 28679
rect 36403 28645 36412 28679
rect 36360 28636 36412 28645
rect 38108 28611 38160 28620
rect 38108 28577 38117 28611
rect 38117 28577 38151 28611
rect 38151 28577 38160 28611
rect 38108 28568 38160 28577
rect 38292 28611 38344 28620
rect 38292 28577 38301 28611
rect 38301 28577 38335 28611
rect 38335 28577 38344 28611
rect 38292 28568 38344 28577
rect 38384 28568 38436 28620
rect 33416 28543 33468 28552
rect 33416 28509 33425 28543
rect 33425 28509 33459 28543
rect 33459 28509 33468 28543
rect 33416 28500 33468 28509
rect 38660 28432 38712 28484
rect 32404 28407 32456 28416
rect 32404 28373 32413 28407
rect 32413 28373 32447 28407
rect 32447 28373 32456 28407
rect 32404 28364 32456 28373
rect 34520 28407 34572 28416
rect 34520 28373 34529 28407
rect 34529 28373 34563 28407
rect 34563 28373 34572 28407
rect 34520 28364 34572 28373
rect 35716 28364 35768 28416
rect 4246 28262 4298 28314
rect 4310 28262 4362 28314
rect 4374 28262 4426 28314
rect 4438 28262 4490 28314
rect 34966 28262 35018 28314
rect 35030 28262 35082 28314
rect 35094 28262 35146 28314
rect 35158 28262 35210 28314
rect 2964 28160 3016 28212
rect 2780 28092 2832 28144
rect 2872 28024 2924 28076
rect 7840 28160 7892 28212
rect 4436 28092 4488 28144
rect 4620 28092 4672 28144
rect 5264 28135 5316 28144
rect 5264 28101 5273 28135
rect 5273 28101 5307 28135
rect 5307 28101 5316 28135
rect 5264 28092 5316 28101
rect 6920 28135 6972 28144
rect 6920 28101 6929 28135
rect 6929 28101 6963 28135
rect 6963 28101 6972 28135
rect 6920 28092 6972 28101
rect 3424 27999 3476 28008
rect 3424 27965 3433 27999
rect 3433 27965 3467 27999
rect 3467 27965 3476 27999
rect 3424 27956 3476 27965
rect 4436 27999 4488 28008
rect 4068 27888 4120 27940
rect 4436 27965 4445 27999
rect 4445 27965 4479 27999
rect 4479 27965 4488 27999
rect 4436 27956 4488 27965
rect 4988 27999 5040 28008
rect 4988 27965 4997 27999
rect 4997 27965 5031 27999
rect 5031 27965 5040 27999
rect 4988 27956 5040 27965
rect 5448 27956 5500 28008
rect 5632 27956 5684 28008
rect 7196 27956 7248 28008
rect 7380 27999 7432 28008
rect 7380 27965 7389 27999
rect 7389 27965 7423 27999
rect 7423 27965 7432 27999
rect 7380 27956 7432 27965
rect 6644 27888 6696 27940
rect 8760 28160 8812 28212
rect 10508 28160 10560 28212
rect 10968 28160 11020 28212
rect 12624 28203 12676 28212
rect 12624 28169 12633 28203
rect 12633 28169 12667 28203
rect 12667 28169 12676 28203
rect 12624 28160 12676 28169
rect 15200 28203 15252 28212
rect 15200 28169 15209 28203
rect 15209 28169 15243 28203
rect 15243 28169 15252 28203
rect 15200 28160 15252 28169
rect 13820 28135 13872 28144
rect 13820 28101 13829 28135
rect 13829 28101 13863 28135
rect 13863 28101 13872 28135
rect 13820 28092 13872 28101
rect 14924 28092 14976 28144
rect 20628 28160 20680 28212
rect 21732 28160 21784 28212
rect 22284 28160 22336 28212
rect 25504 28203 25556 28212
rect 9956 28024 10008 28076
rect 10968 28024 11020 28076
rect 8300 27999 8352 28008
rect 8300 27965 8309 27999
rect 8309 27965 8343 27999
rect 8343 27965 8352 27999
rect 8300 27956 8352 27965
rect 9128 27956 9180 28008
rect 10048 27956 10100 28008
rect 10232 27999 10284 28008
rect 10232 27965 10241 27999
rect 10241 27965 10275 27999
rect 10275 27965 10284 27999
rect 10232 27956 10284 27965
rect 11428 27956 11480 28008
rect 12808 27956 12860 28008
rect 16672 28067 16724 28076
rect 13176 27888 13228 27940
rect 14464 27956 14516 28008
rect 15844 27999 15896 28008
rect 15844 27965 15853 27999
rect 15853 27965 15887 27999
rect 15887 27965 15896 27999
rect 15844 27956 15896 27965
rect 15384 27888 15436 27940
rect 16672 28033 16681 28067
rect 16681 28033 16715 28067
rect 16715 28033 16724 28067
rect 16672 28024 16724 28033
rect 18236 28024 18288 28076
rect 19708 28092 19760 28144
rect 17868 27956 17920 28008
rect 18328 27999 18380 28008
rect 18328 27965 18337 27999
rect 18337 27965 18371 27999
rect 18371 27965 18380 27999
rect 18328 27956 18380 27965
rect 19432 28024 19484 28076
rect 19156 27999 19208 28008
rect 19156 27965 19165 27999
rect 19165 27965 19199 27999
rect 19199 27965 19208 27999
rect 19156 27956 19208 27965
rect 19340 27999 19392 28008
rect 19340 27965 19349 27999
rect 19349 27965 19383 27999
rect 19383 27965 19392 27999
rect 19340 27956 19392 27965
rect 19616 27956 19668 28008
rect 17592 27888 17644 27940
rect 20812 27956 20864 28008
rect 21548 28024 21600 28076
rect 21364 27999 21416 28008
rect 21364 27965 21373 27999
rect 21373 27965 21407 27999
rect 21407 27965 21416 27999
rect 21364 27956 21416 27965
rect 21916 27999 21968 28008
rect 21916 27965 21925 27999
rect 21925 27965 21959 27999
rect 21959 27965 21968 27999
rect 21916 27956 21968 27965
rect 22284 27999 22336 28008
rect 22284 27965 22293 27999
rect 22293 27965 22327 27999
rect 22327 27965 22336 27999
rect 22284 27956 22336 27965
rect 25504 28169 25513 28203
rect 25513 28169 25547 28203
rect 25547 28169 25556 28203
rect 25504 28160 25556 28169
rect 29552 28203 29604 28212
rect 29552 28169 29561 28203
rect 29561 28169 29595 28203
rect 29595 28169 29604 28203
rect 29552 28160 29604 28169
rect 30012 28160 30064 28212
rect 24124 28135 24176 28144
rect 24124 28101 24133 28135
rect 24133 28101 24167 28135
rect 24167 28101 24176 28135
rect 24124 28092 24176 28101
rect 24032 28024 24084 28076
rect 24308 28024 24360 28076
rect 27804 28067 27856 28076
rect 25412 27999 25464 28008
rect 21732 27888 21784 27940
rect 2596 27820 2648 27872
rect 9864 27820 9916 27872
rect 10784 27820 10836 27872
rect 12072 27820 12124 27872
rect 15936 27863 15988 27872
rect 15936 27829 15945 27863
rect 15945 27829 15979 27863
rect 15979 27829 15988 27863
rect 15936 27820 15988 27829
rect 21640 27820 21692 27872
rect 22744 27820 22796 27872
rect 25412 27965 25421 27999
rect 25421 27965 25455 27999
rect 25455 27965 25464 27999
rect 25412 27956 25464 27965
rect 25780 27956 25832 28008
rect 25964 27999 26016 28008
rect 25964 27965 25973 27999
rect 25973 27965 26007 27999
rect 26007 27965 26016 27999
rect 25964 27956 26016 27965
rect 26424 27999 26476 28008
rect 26424 27965 26433 27999
rect 26433 27965 26467 27999
rect 26467 27965 26476 27999
rect 26424 27956 26476 27965
rect 26884 27956 26936 28008
rect 27804 28033 27813 28067
rect 27813 28033 27847 28067
rect 27847 28033 27856 28067
rect 27804 28024 27856 28033
rect 29184 28092 29236 28144
rect 29276 28067 29328 28076
rect 29276 28033 29285 28067
rect 29285 28033 29319 28067
rect 29319 28033 29328 28067
rect 29276 28024 29328 28033
rect 30012 28024 30064 28076
rect 32404 28024 32456 28076
rect 24768 27888 24820 27940
rect 26516 27888 26568 27940
rect 27068 27931 27120 27940
rect 27068 27897 27077 27931
rect 27077 27897 27111 27931
rect 27111 27897 27120 27931
rect 27068 27888 27120 27897
rect 27528 27888 27580 27940
rect 29368 27999 29420 28008
rect 29368 27965 29377 27999
rect 29377 27965 29411 27999
rect 29411 27965 29420 27999
rect 33508 28160 33560 28212
rect 37740 28160 37792 28212
rect 33416 28067 33468 28076
rect 33416 28033 33425 28067
rect 33425 28033 33459 28067
rect 33459 28033 33468 28067
rect 33416 28024 33468 28033
rect 37556 28067 37608 28076
rect 37556 28033 37565 28067
rect 37565 28033 37599 28067
rect 37599 28033 37608 28067
rect 37556 28024 37608 28033
rect 29368 27956 29420 27965
rect 24032 27820 24084 27872
rect 25688 27820 25740 27872
rect 25872 27820 25924 27872
rect 29460 27820 29512 27872
rect 31392 27820 31444 27872
rect 31852 27863 31904 27872
rect 31852 27829 31861 27863
rect 31861 27829 31895 27863
rect 31895 27829 31904 27863
rect 31852 27820 31904 27829
rect 33324 27999 33376 28008
rect 33324 27965 33333 27999
rect 33333 27965 33367 27999
rect 33367 27965 33376 27999
rect 33324 27956 33376 27965
rect 33968 27999 34020 28008
rect 33968 27965 33977 27999
rect 33977 27965 34011 27999
rect 34011 27965 34020 27999
rect 33968 27956 34020 27965
rect 36084 27956 36136 28008
rect 37280 27999 37332 28008
rect 37280 27965 37289 27999
rect 37289 27965 37323 27999
rect 37323 27965 37332 27999
rect 37280 27956 37332 27965
rect 33508 27888 33560 27940
rect 34060 27820 34112 27872
rect 38016 27820 38068 27872
rect 19606 27718 19658 27770
rect 19670 27718 19722 27770
rect 19734 27718 19786 27770
rect 19798 27718 19850 27770
rect 4160 27659 4212 27668
rect 4160 27625 4169 27659
rect 4169 27625 4203 27659
rect 4203 27625 4212 27659
rect 4160 27616 4212 27625
rect 15936 27616 15988 27668
rect 5540 27548 5592 27600
rect 2044 27480 2096 27532
rect 2504 27523 2556 27532
rect 2504 27489 2513 27523
rect 2513 27489 2547 27523
rect 2547 27489 2556 27523
rect 2504 27480 2556 27489
rect 2596 27523 2648 27532
rect 2596 27489 2605 27523
rect 2605 27489 2639 27523
rect 2639 27489 2648 27523
rect 2596 27480 2648 27489
rect 3424 27480 3476 27532
rect 3884 27523 3936 27532
rect 3884 27489 3893 27523
rect 3893 27489 3927 27523
rect 3927 27489 3936 27523
rect 3884 27480 3936 27489
rect 4068 27523 4120 27532
rect 4068 27489 4077 27523
rect 4077 27489 4111 27523
rect 4111 27489 4120 27523
rect 4068 27480 4120 27489
rect 4620 27523 4672 27532
rect 4620 27489 4629 27523
rect 4629 27489 4663 27523
rect 4663 27489 4672 27523
rect 4620 27480 4672 27489
rect 4988 27523 5040 27532
rect 4988 27489 4997 27523
rect 4997 27489 5031 27523
rect 5031 27489 5040 27523
rect 4988 27480 5040 27489
rect 6920 27548 6972 27600
rect 7380 27548 7432 27600
rect 6000 27480 6052 27532
rect 8300 27548 8352 27600
rect 10876 27591 10928 27600
rect 7656 27523 7708 27532
rect 7656 27489 7665 27523
rect 7665 27489 7699 27523
rect 7699 27489 7708 27523
rect 7932 27523 7984 27532
rect 7656 27480 7708 27489
rect 7932 27489 7941 27523
rect 7941 27489 7975 27523
rect 7975 27489 7984 27523
rect 7932 27480 7984 27489
rect 5724 27412 5776 27464
rect 6644 27412 6696 27464
rect 9128 27480 9180 27532
rect 10232 27523 10284 27532
rect 10232 27489 10241 27523
rect 10241 27489 10275 27523
rect 10275 27489 10284 27523
rect 10232 27480 10284 27489
rect 10876 27557 10885 27591
rect 10885 27557 10919 27591
rect 10919 27557 10928 27591
rect 10876 27548 10928 27557
rect 11336 27523 11388 27532
rect 11336 27489 11345 27523
rect 11345 27489 11379 27523
rect 11379 27489 11388 27523
rect 11336 27480 11388 27489
rect 12072 27523 12124 27532
rect 12072 27489 12081 27523
rect 12081 27489 12115 27523
rect 12115 27489 12124 27523
rect 12072 27480 12124 27489
rect 12440 27523 12492 27532
rect 12440 27489 12449 27523
rect 12449 27489 12483 27523
rect 12483 27489 12492 27523
rect 14280 27548 14332 27600
rect 15384 27591 15436 27600
rect 12440 27480 12492 27489
rect 8576 27412 8628 27464
rect 11796 27412 11848 27464
rect 1400 27344 1452 27396
rect 3976 27344 4028 27396
rect 6552 27344 6604 27396
rect 2044 27276 2096 27328
rect 2780 27319 2832 27328
rect 2780 27285 2789 27319
rect 2789 27285 2823 27319
rect 2823 27285 2832 27319
rect 5724 27319 5776 27328
rect 2780 27276 2832 27285
rect 5724 27285 5733 27319
rect 5733 27285 5767 27319
rect 5767 27285 5776 27319
rect 5724 27276 5776 27285
rect 5816 27276 5868 27328
rect 11980 27344 12032 27396
rect 14464 27480 14516 27532
rect 14556 27523 14608 27532
rect 14556 27489 14565 27523
rect 14565 27489 14599 27523
rect 14599 27489 14608 27523
rect 15384 27557 15393 27591
rect 15393 27557 15427 27591
rect 15427 27557 15436 27591
rect 15384 27548 15436 27557
rect 14556 27480 14608 27489
rect 13728 27344 13780 27396
rect 8300 27276 8352 27328
rect 9036 27319 9088 27328
rect 9036 27285 9045 27319
rect 9045 27285 9079 27319
rect 9079 27285 9088 27319
rect 9036 27276 9088 27285
rect 11060 27276 11112 27328
rect 17040 27480 17092 27532
rect 17960 27548 18012 27600
rect 21824 27548 21876 27600
rect 23572 27548 23624 27600
rect 19432 27480 19484 27532
rect 19892 27480 19944 27532
rect 19984 27480 20036 27532
rect 17224 27455 17276 27464
rect 17224 27421 17233 27455
rect 17233 27421 17267 27455
rect 17267 27421 17276 27455
rect 17224 27412 17276 27421
rect 17408 27412 17460 27464
rect 17040 27344 17092 27396
rect 17316 27344 17368 27396
rect 17868 27387 17920 27396
rect 17868 27353 17877 27387
rect 17877 27353 17911 27387
rect 17911 27353 17920 27387
rect 17868 27344 17920 27353
rect 20720 27480 20772 27532
rect 21088 27523 21140 27532
rect 21088 27489 21097 27523
rect 21097 27489 21131 27523
rect 21131 27489 21140 27523
rect 21088 27480 21140 27489
rect 21548 27523 21600 27532
rect 21548 27489 21557 27523
rect 21557 27489 21591 27523
rect 21591 27489 21600 27523
rect 21548 27480 21600 27489
rect 22284 27480 22336 27532
rect 24032 27616 24084 27668
rect 25412 27616 25464 27668
rect 25688 27616 25740 27668
rect 27528 27616 27580 27668
rect 24768 27548 24820 27600
rect 20352 27455 20404 27464
rect 20352 27421 20361 27455
rect 20361 27421 20395 27455
rect 20395 27421 20404 27455
rect 20352 27412 20404 27421
rect 20812 27344 20864 27396
rect 18604 27276 18656 27328
rect 21364 27276 21416 27328
rect 21732 27344 21784 27396
rect 22468 27276 22520 27328
rect 23940 27412 23992 27464
rect 24492 27480 24544 27532
rect 24032 27344 24084 27396
rect 25412 27480 25464 27532
rect 25596 27523 25648 27532
rect 25596 27489 25605 27523
rect 25605 27489 25639 27523
rect 25639 27489 25648 27523
rect 25596 27480 25648 27489
rect 27068 27548 27120 27600
rect 29644 27616 29696 27668
rect 28264 27548 28316 27600
rect 29092 27523 29144 27532
rect 29092 27489 29101 27523
rect 29101 27489 29135 27523
rect 29135 27489 29144 27523
rect 29092 27480 29144 27489
rect 29184 27480 29236 27532
rect 30472 27480 30524 27532
rect 30656 27523 30708 27532
rect 30656 27489 30665 27523
rect 30665 27489 30699 27523
rect 30699 27489 30708 27523
rect 30656 27480 30708 27489
rect 29000 27344 29052 27396
rect 29460 27387 29512 27396
rect 29460 27353 29469 27387
rect 29469 27353 29503 27387
rect 29503 27353 29512 27387
rect 29460 27344 29512 27353
rect 30380 27412 30432 27464
rect 32036 27480 32088 27532
rect 34520 27548 34572 27600
rect 37096 27548 37148 27600
rect 38384 27548 38436 27600
rect 33324 27480 33376 27532
rect 33968 27480 34020 27532
rect 34244 27523 34296 27532
rect 34244 27489 34253 27523
rect 34253 27489 34287 27523
rect 34287 27489 34296 27523
rect 34244 27480 34296 27489
rect 35716 27480 35768 27532
rect 35808 27523 35860 27532
rect 35808 27489 35817 27523
rect 35817 27489 35851 27523
rect 35851 27489 35860 27523
rect 35808 27480 35860 27489
rect 38016 27523 38068 27532
rect 38016 27489 38025 27523
rect 38025 27489 38059 27523
rect 38059 27489 38068 27523
rect 38016 27480 38068 27489
rect 38292 27523 38344 27532
rect 38292 27489 38301 27523
rect 38301 27489 38335 27523
rect 38335 27489 38344 27523
rect 38292 27480 38344 27489
rect 38568 27480 38620 27532
rect 31852 27412 31904 27464
rect 33048 27412 33100 27464
rect 30932 27387 30984 27396
rect 30932 27353 30941 27387
rect 30941 27353 30975 27387
rect 30975 27353 30984 27387
rect 30932 27344 30984 27353
rect 31484 27344 31536 27396
rect 32496 27387 32548 27396
rect 24860 27276 24912 27328
rect 26976 27276 27028 27328
rect 29736 27276 29788 27328
rect 30564 27276 30616 27328
rect 31024 27276 31076 27328
rect 32496 27353 32505 27387
rect 32505 27353 32539 27387
rect 32539 27353 32548 27387
rect 32496 27344 32548 27353
rect 33968 27344 34020 27396
rect 35900 27387 35952 27396
rect 34152 27276 34204 27328
rect 35900 27353 35909 27387
rect 35909 27353 35943 27387
rect 35943 27353 35952 27387
rect 35900 27344 35952 27353
rect 36636 27344 36688 27396
rect 38844 27276 38896 27328
rect 39948 27251 40000 27260
rect 4246 27174 4298 27226
rect 4310 27174 4362 27226
rect 4374 27174 4426 27226
rect 4438 27174 4490 27226
rect 34966 27174 35018 27226
rect 35030 27174 35082 27226
rect 35094 27174 35146 27226
rect 35158 27174 35210 27226
rect 39948 27217 39957 27251
rect 39957 27217 39991 27251
rect 39991 27217 40000 27251
rect 39948 27208 40000 27217
rect 5632 27072 5684 27124
rect 6644 27072 6696 27124
rect 13452 27072 13504 27124
rect 13728 27072 13780 27124
rect 2780 26936 2832 26988
rect 5724 26936 5776 26988
rect 1400 26868 1452 26920
rect 2596 26868 2648 26920
rect 4252 26911 4304 26920
rect 4252 26877 4261 26911
rect 4261 26877 4295 26911
rect 4295 26877 4304 26911
rect 4252 26868 4304 26877
rect 4804 26868 4856 26920
rect 5632 26868 5684 26920
rect 6000 26911 6052 26920
rect 6000 26877 6009 26911
rect 6009 26877 6043 26911
rect 6043 26877 6052 26911
rect 6000 26868 6052 26877
rect 6552 26868 6604 26920
rect 9036 26868 9088 26920
rect 10508 26936 10560 26988
rect 10600 26936 10652 26988
rect 10876 26936 10928 26988
rect 11060 26868 11112 26920
rect 11428 26911 11480 26920
rect 11428 26877 11437 26911
rect 11437 26877 11471 26911
rect 11471 26877 11480 26911
rect 11428 26868 11480 26877
rect 11888 26911 11940 26920
rect 11888 26877 11897 26911
rect 11897 26877 11931 26911
rect 11931 26877 11940 26911
rect 11888 26868 11940 26877
rect 13544 26911 13596 26920
rect 13544 26877 13553 26911
rect 13553 26877 13587 26911
rect 13587 26877 13596 26911
rect 13544 26868 13596 26877
rect 13820 26911 13872 26920
rect 13820 26877 13829 26911
rect 13829 26877 13863 26911
rect 13863 26877 13872 26911
rect 17960 26936 18012 26988
rect 13820 26868 13872 26877
rect 16580 26911 16632 26920
rect 16580 26877 16589 26911
rect 16589 26877 16623 26911
rect 16623 26877 16632 26911
rect 16580 26868 16632 26877
rect 16856 26911 16908 26920
rect 16856 26877 16865 26911
rect 16865 26877 16899 26911
rect 16899 26877 16908 26911
rect 16856 26868 16908 26877
rect 17408 26868 17460 26920
rect 23572 27072 23624 27124
rect 34796 27072 34848 27124
rect 35624 27072 35676 27124
rect 8576 26800 8628 26852
rect 11980 26800 12032 26852
rect 13636 26800 13688 26852
rect 2504 26732 2556 26784
rect 5724 26732 5776 26784
rect 9680 26732 9732 26784
rect 10600 26775 10652 26784
rect 10600 26741 10609 26775
rect 10609 26741 10643 26775
rect 10643 26741 10652 26775
rect 10600 26732 10652 26741
rect 12440 26732 12492 26784
rect 13820 26732 13872 26784
rect 15476 26800 15528 26852
rect 19156 26936 19208 26988
rect 18604 26868 18656 26920
rect 18788 26911 18840 26920
rect 18788 26877 18797 26911
rect 18797 26877 18831 26911
rect 18831 26877 18840 26911
rect 18788 26868 18840 26877
rect 22192 27004 22244 27056
rect 20536 26936 20588 26988
rect 20352 26868 20404 26920
rect 22100 26936 22152 26988
rect 25320 27004 25372 27056
rect 29736 27047 29788 27056
rect 24032 26979 24084 26988
rect 24032 26945 24041 26979
rect 24041 26945 24075 26979
rect 24075 26945 24084 26979
rect 24032 26936 24084 26945
rect 24768 26936 24820 26988
rect 22192 26911 22244 26920
rect 22192 26877 22201 26911
rect 22201 26877 22235 26911
rect 22235 26877 22244 26911
rect 22192 26868 22244 26877
rect 22744 26868 22796 26920
rect 23572 26868 23624 26920
rect 25964 26936 26016 26988
rect 17868 26732 17920 26784
rect 19156 26732 19208 26784
rect 22560 26732 22612 26784
rect 23020 26775 23072 26784
rect 23020 26741 23029 26775
rect 23029 26741 23063 26775
rect 23063 26741 23072 26775
rect 23020 26732 23072 26741
rect 26884 26911 26936 26920
rect 26884 26877 26893 26911
rect 26893 26877 26927 26911
rect 26927 26877 26936 26911
rect 26884 26868 26936 26877
rect 29460 26936 29512 26988
rect 29736 27013 29745 27047
rect 29745 27013 29779 27047
rect 29779 27013 29788 27047
rect 29736 27004 29788 27013
rect 30288 27004 30340 27056
rect 36084 27047 36136 27056
rect 36084 27013 36093 27047
rect 36093 27013 36127 27047
rect 36127 27013 36136 27047
rect 36084 27004 36136 27013
rect 25412 26843 25464 26852
rect 25412 26809 25421 26843
rect 25421 26809 25455 26843
rect 25455 26809 25464 26843
rect 25412 26800 25464 26809
rect 28356 26800 28408 26852
rect 28632 26911 28684 26920
rect 28632 26877 28641 26911
rect 28641 26877 28675 26911
rect 28675 26877 28684 26911
rect 34152 26979 34204 26988
rect 28632 26868 28684 26877
rect 30012 26868 30064 26920
rect 30932 26911 30984 26920
rect 30932 26877 30941 26911
rect 30941 26877 30975 26911
rect 30975 26877 30984 26911
rect 30932 26868 30984 26877
rect 33140 26911 33192 26920
rect 33140 26877 33149 26911
rect 33149 26877 33183 26911
rect 33183 26877 33192 26911
rect 33140 26868 33192 26877
rect 34152 26945 34161 26979
rect 34161 26945 34195 26979
rect 34195 26945 34204 26979
rect 34152 26936 34204 26945
rect 37832 26936 37884 26988
rect 38568 26979 38620 26988
rect 38568 26945 38577 26979
rect 38577 26945 38611 26979
rect 38611 26945 38620 26979
rect 38568 26936 38620 26945
rect 34060 26868 34112 26920
rect 35256 26868 35308 26920
rect 35900 26911 35952 26920
rect 35900 26877 35909 26911
rect 35909 26877 35943 26911
rect 35943 26877 35952 26911
rect 35900 26868 35952 26877
rect 36636 26911 36688 26920
rect 36636 26877 36645 26911
rect 36645 26877 36679 26911
rect 36679 26877 36688 26911
rect 36636 26868 36688 26877
rect 37740 26868 37792 26920
rect 30564 26800 30616 26852
rect 37096 26800 37148 26852
rect 31024 26732 31076 26784
rect 31208 26732 31260 26784
rect 33048 26732 33100 26784
rect 33784 26732 33836 26784
rect 19606 26630 19658 26682
rect 19670 26630 19722 26682
rect 19734 26630 19786 26682
rect 19798 26630 19850 26682
rect 2044 26503 2096 26512
rect 2044 26469 2053 26503
rect 2053 26469 2087 26503
rect 2087 26469 2096 26503
rect 2044 26460 2096 26469
rect 2596 26435 2648 26444
rect 2596 26401 2605 26435
rect 2605 26401 2639 26435
rect 2639 26401 2648 26435
rect 2596 26392 2648 26401
rect 2688 26435 2740 26444
rect 2688 26401 2697 26435
rect 2697 26401 2731 26435
rect 2731 26401 2740 26435
rect 4068 26528 4120 26580
rect 5632 26571 5684 26580
rect 5632 26537 5641 26571
rect 5641 26537 5675 26571
rect 5675 26537 5684 26571
rect 5632 26528 5684 26537
rect 5724 26528 5776 26580
rect 11888 26528 11940 26580
rect 18512 26571 18564 26580
rect 2688 26392 2740 26401
rect 3148 26435 3200 26444
rect 3148 26401 3157 26435
rect 3157 26401 3191 26435
rect 3191 26401 3200 26435
rect 3148 26392 3200 26401
rect 3976 26392 4028 26444
rect 6000 26392 6052 26444
rect 7380 26435 7432 26444
rect 7380 26401 7389 26435
rect 7389 26401 7423 26435
rect 7423 26401 7432 26435
rect 7380 26392 7432 26401
rect 7748 26435 7800 26444
rect 7748 26401 7757 26435
rect 7757 26401 7791 26435
rect 7791 26401 7800 26435
rect 7748 26392 7800 26401
rect 8116 26435 8168 26444
rect 8116 26401 8125 26435
rect 8125 26401 8159 26435
rect 8159 26401 8168 26435
rect 8116 26392 8168 26401
rect 8576 26435 8628 26444
rect 8576 26401 8585 26435
rect 8585 26401 8619 26435
rect 8619 26401 8628 26435
rect 8576 26392 8628 26401
rect 12072 26435 12124 26444
rect 12072 26401 12081 26435
rect 12081 26401 12115 26435
rect 12115 26401 12124 26435
rect 12072 26392 12124 26401
rect 12440 26460 12492 26512
rect 12624 26460 12676 26512
rect 12348 26392 12400 26444
rect 2780 26256 2832 26308
rect 4252 26324 4304 26376
rect 4712 26324 4764 26376
rect 7196 26367 7248 26376
rect 7196 26333 7205 26367
rect 7205 26333 7239 26367
rect 7239 26333 7248 26367
rect 7196 26324 7248 26333
rect 9680 26367 9732 26376
rect 9680 26333 9689 26367
rect 9689 26333 9723 26367
rect 9723 26333 9732 26367
rect 9680 26324 9732 26333
rect 9864 26324 9916 26376
rect 11336 26367 11388 26376
rect 11336 26333 11345 26367
rect 11345 26333 11379 26367
rect 11379 26333 11388 26367
rect 13268 26392 13320 26444
rect 13728 26435 13780 26444
rect 13728 26401 13737 26435
rect 13737 26401 13771 26435
rect 13771 26401 13780 26435
rect 13728 26392 13780 26401
rect 13820 26392 13872 26444
rect 15108 26435 15160 26444
rect 15108 26401 15117 26435
rect 15117 26401 15151 26435
rect 15151 26401 15160 26435
rect 15108 26392 15160 26401
rect 16120 26435 16172 26444
rect 16120 26401 16129 26435
rect 16129 26401 16163 26435
rect 16163 26401 16172 26435
rect 16120 26392 16172 26401
rect 11336 26324 11388 26333
rect 12808 26367 12860 26376
rect 12808 26333 12817 26367
rect 12817 26333 12851 26367
rect 12851 26333 12860 26367
rect 12808 26324 12860 26333
rect 13176 26324 13228 26376
rect 18512 26537 18521 26571
rect 18521 26537 18555 26571
rect 18555 26537 18564 26571
rect 18512 26528 18564 26537
rect 22100 26528 22152 26580
rect 25596 26528 25648 26580
rect 16396 26392 16448 26444
rect 17132 26392 17184 26444
rect 17868 26392 17920 26444
rect 18144 26392 18196 26444
rect 18788 26392 18840 26444
rect 19156 26435 19208 26444
rect 19156 26401 19165 26435
rect 19165 26401 19199 26435
rect 19199 26401 19208 26435
rect 19156 26392 19208 26401
rect 22192 26460 22244 26512
rect 20812 26392 20864 26444
rect 21640 26435 21692 26444
rect 21640 26401 21649 26435
rect 21649 26401 21683 26435
rect 21683 26401 21692 26435
rect 21640 26392 21692 26401
rect 22376 26435 22428 26444
rect 22376 26401 22385 26435
rect 22385 26401 22419 26435
rect 22419 26401 22428 26435
rect 22376 26392 22428 26401
rect 22928 26435 22980 26444
rect 22928 26401 22937 26435
rect 22937 26401 22971 26435
rect 22971 26401 22980 26435
rect 22928 26392 22980 26401
rect 23848 26435 23900 26444
rect 23848 26401 23857 26435
rect 23857 26401 23891 26435
rect 23891 26401 23900 26435
rect 23848 26392 23900 26401
rect 24492 26435 24544 26444
rect 24492 26401 24501 26435
rect 24501 26401 24535 26435
rect 24535 26401 24544 26435
rect 24492 26392 24544 26401
rect 23112 26367 23164 26376
rect 23112 26333 23121 26367
rect 23121 26333 23155 26367
rect 23155 26333 23164 26367
rect 23112 26324 23164 26333
rect 23572 26324 23624 26376
rect 25320 26392 25372 26444
rect 26884 26460 26936 26512
rect 25780 26435 25832 26444
rect 25780 26401 25789 26435
rect 25789 26401 25823 26435
rect 25823 26401 25832 26435
rect 25780 26392 25832 26401
rect 28172 26392 28224 26444
rect 12624 26256 12676 26308
rect 13636 26256 13688 26308
rect 15200 26256 15252 26308
rect 5356 26188 5408 26240
rect 11060 26188 11112 26240
rect 14924 26231 14976 26240
rect 14924 26197 14933 26231
rect 14933 26197 14967 26231
rect 14967 26197 14976 26231
rect 14924 26188 14976 26197
rect 21088 26231 21140 26240
rect 21088 26197 21097 26231
rect 21097 26197 21131 26231
rect 21131 26197 21140 26231
rect 21088 26188 21140 26197
rect 23940 26299 23992 26308
rect 23296 26188 23348 26240
rect 23940 26265 23949 26299
rect 23949 26265 23983 26299
rect 23983 26265 23992 26299
rect 23940 26256 23992 26265
rect 27252 26367 27304 26376
rect 27252 26333 27261 26367
rect 27261 26333 27295 26367
rect 27295 26333 27304 26367
rect 27252 26324 27304 26333
rect 27620 26324 27672 26376
rect 26608 26256 26660 26308
rect 28632 26528 28684 26580
rect 31484 26571 31536 26580
rect 31484 26537 31493 26571
rect 31493 26537 31527 26571
rect 31527 26537 31536 26571
rect 31484 26528 31536 26537
rect 28356 26460 28408 26512
rect 31208 26460 31260 26512
rect 29552 26392 29604 26444
rect 33140 26460 33192 26512
rect 37924 26528 37976 26580
rect 38476 26571 38528 26580
rect 38476 26537 38485 26571
rect 38485 26537 38519 26571
rect 38519 26537 38528 26571
rect 38476 26528 38528 26537
rect 38660 26460 38712 26512
rect 29368 26324 29420 26376
rect 32036 26392 32088 26444
rect 33784 26435 33836 26444
rect 30748 26324 30800 26376
rect 33324 26324 33376 26376
rect 33508 26367 33560 26376
rect 33508 26333 33517 26367
rect 33517 26333 33551 26367
rect 33551 26333 33560 26367
rect 33508 26324 33560 26333
rect 33784 26401 33793 26435
rect 33793 26401 33827 26435
rect 33827 26401 33836 26435
rect 33784 26392 33836 26401
rect 35992 26435 36044 26444
rect 35992 26401 36001 26435
rect 36001 26401 36035 26435
rect 36035 26401 36044 26435
rect 35992 26392 36044 26401
rect 36268 26392 36320 26444
rect 37740 26435 37792 26444
rect 35348 26324 35400 26376
rect 35716 26324 35768 26376
rect 37740 26401 37749 26435
rect 37749 26401 37783 26435
rect 37783 26401 37792 26435
rect 37740 26392 37792 26401
rect 38384 26392 38436 26444
rect 38752 26392 38804 26444
rect 38292 26324 38344 26376
rect 24584 26188 24636 26240
rect 32496 26256 32548 26308
rect 27712 26188 27764 26240
rect 28172 26188 28224 26240
rect 36084 26231 36136 26240
rect 36084 26197 36093 26231
rect 36093 26197 36127 26231
rect 36127 26197 36136 26231
rect 36084 26188 36136 26197
rect 4246 26086 4298 26138
rect 4310 26086 4362 26138
rect 4374 26086 4426 26138
rect 4438 26086 4490 26138
rect 34966 26086 35018 26138
rect 35030 26086 35082 26138
rect 35094 26086 35146 26138
rect 35158 26086 35210 26138
rect 2688 25984 2740 26036
rect 5448 25984 5500 26036
rect 9404 25984 9456 26036
rect 3608 25916 3660 25968
rect 4068 25916 4120 25968
rect 5908 25916 5960 25968
rect 2412 25891 2464 25900
rect 2412 25857 2421 25891
rect 2421 25857 2455 25891
rect 2455 25857 2464 25891
rect 2412 25848 2464 25857
rect 5448 25891 5500 25900
rect 5448 25857 5457 25891
rect 5457 25857 5491 25891
rect 5491 25857 5500 25891
rect 5448 25848 5500 25857
rect 7380 25848 7432 25900
rect 9956 25916 10008 25968
rect 9864 25848 9916 25900
rect 1768 25823 1820 25832
rect 1768 25789 1777 25823
rect 1777 25789 1811 25823
rect 1811 25789 1820 25823
rect 1768 25780 1820 25789
rect 2320 25780 2372 25832
rect 2964 25780 3016 25832
rect 3608 25780 3660 25832
rect 4068 25780 4120 25832
rect 5724 25823 5776 25832
rect 4620 25712 4672 25764
rect 1676 25644 1728 25696
rect 3148 25644 3200 25696
rect 4068 25644 4120 25696
rect 5724 25789 5733 25823
rect 5733 25789 5767 25823
rect 5767 25789 5776 25823
rect 5724 25780 5776 25789
rect 6184 25823 6236 25832
rect 6184 25789 6193 25823
rect 6193 25789 6227 25823
rect 6227 25789 6236 25823
rect 6184 25780 6236 25789
rect 7748 25780 7800 25832
rect 8116 25823 8168 25832
rect 8116 25789 8125 25823
rect 8125 25789 8159 25823
rect 8159 25789 8168 25823
rect 8116 25780 8168 25789
rect 9496 25823 9548 25832
rect 9496 25789 9505 25823
rect 9505 25789 9539 25823
rect 9539 25789 9548 25823
rect 9496 25780 9548 25789
rect 9956 25823 10008 25832
rect 5356 25644 5408 25696
rect 9036 25712 9088 25764
rect 9956 25789 9965 25823
rect 9965 25789 9999 25823
rect 9999 25789 10008 25823
rect 9956 25780 10008 25789
rect 10692 25984 10744 26036
rect 11428 25984 11480 26036
rect 14280 25984 14332 26036
rect 16580 25984 16632 26036
rect 18328 26027 18380 26036
rect 18328 25993 18337 26027
rect 18337 25993 18371 26027
rect 18371 25993 18380 26027
rect 18328 25984 18380 25993
rect 22560 25984 22612 26036
rect 23572 25984 23624 26036
rect 25596 25984 25648 26036
rect 33324 26027 33376 26036
rect 33324 25993 33333 26027
rect 33333 25993 33367 26027
rect 33367 25993 33376 26027
rect 33324 25984 33376 25993
rect 34244 25984 34296 26036
rect 36268 25984 36320 26036
rect 38660 26027 38712 26036
rect 38660 25993 38669 26027
rect 38669 25993 38703 26027
rect 38703 25993 38712 26027
rect 38660 25984 38712 25993
rect 10600 25848 10652 25900
rect 11336 25823 11388 25832
rect 10968 25712 11020 25764
rect 5908 25644 5960 25696
rect 7656 25644 7708 25696
rect 8852 25644 8904 25696
rect 11336 25789 11345 25823
rect 11345 25789 11379 25823
rect 11379 25789 11388 25823
rect 11336 25780 11388 25789
rect 12440 25780 12492 25832
rect 13360 25823 13412 25832
rect 13360 25789 13369 25823
rect 13369 25789 13403 25823
rect 13403 25789 13412 25823
rect 13360 25780 13412 25789
rect 13636 25823 13688 25832
rect 13636 25789 13645 25823
rect 13645 25789 13679 25823
rect 13679 25789 13688 25823
rect 13636 25780 13688 25789
rect 13820 25823 13872 25832
rect 13820 25789 13829 25823
rect 13829 25789 13863 25823
rect 13863 25789 13872 25823
rect 13820 25780 13872 25789
rect 14280 25823 14332 25832
rect 14280 25789 14289 25823
rect 14289 25789 14323 25823
rect 14323 25789 14332 25823
rect 14280 25780 14332 25789
rect 13912 25712 13964 25764
rect 16120 25780 16172 25832
rect 16396 25780 16448 25832
rect 25228 25959 25280 25968
rect 17132 25823 17184 25832
rect 17132 25789 17141 25823
rect 17141 25789 17175 25823
rect 17175 25789 17184 25823
rect 17132 25780 17184 25789
rect 17960 25780 18012 25832
rect 18144 25780 18196 25832
rect 18328 25780 18380 25832
rect 20076 25848 20128 25900
rect 25228 25925 25237 25959
rect 25237 25925 25271 25959
rect 25271 25925 25280 25959
rect 25228 25916 25280 25925
rect 30104 25916 30156 25968
rect 19984 25823 20036 25832
rect 19984 25789 19993 25823
rect 19993 25789 20027 25823
rect 20027 25789 20036 25823
rect 19984 25780 20036 25789
rect 20720 25823 20772 25832
rect 20720 25789 20729 25823
rect 20729 25789 20763 25823
rect 20763 25789 20772 25823
rect 20720 25780 20772 25789
rect 22008 25823 22060 25832
rect 22008 25789 22017 25823
rect 22017 25789 22051 25823
rect 22051 25789 22060 25823
rect 22008 25780 22060 25789
rect 22284 25823 22336 25832
rect 22284 25789 22293 25823
rect 22293 25789 22327 25823
rect 22327 25789 22336 25823
rect 22284 25780 22336 25789
rect 22652 25780 22704 25832
rect 23572 25780 23624 25832
rect 15660 25712 15712 25764
rect 22560 25712 22612 25764
rect 11980 25644 12032 25696
rect 12256 25644 12308 25696
rect 17316 25687 17368 25696
rect 17316 25653 17325 25687
rect 17325 25653 17359 25687
rect 17359 25653 17368 25687
rect 17316 25644 17368 25653
rect 23848 25644 23900 25696
rect 24584 25780 24636 25832
rect 25412 25823 25464 25832
rect 25412 25789 25421 25823
rect 25421 25789 25455 25823
rect 25455 25789 25464 25823
rect 25412 25780 25464 25789
rect 26976 25848 27028 25900
rect 25964 25780 26016 25832
rect 33508 25848 33560 25900
rect 37280 25891 37332 25900
rect 37280 25857 37289 25891
rect 37289 25857 37323 25891
rect 37323 25857 37332 25891
rect 37280 25848 37332 25857
rect 27252 25823 27304 25832
rect 27252 25789 27261 25823
rect 27261 25789 27295 25823
rect 27295 25789 27304 25823
rect 27252 25780 27304 25789
rect 28172 25823 28224 25832
rect 28172 25789 28181 25823
rect 28181 25789 28215 25823
rect 28215 25789 28224 25823
rect 28172 25780 28224 25789
rect 28264 25780 28316 25832
rect 29552 25780 29604 25832
rect 30564 25823 30616 25832
rect 25044 25712 25096 25764
rect 30564 25789 30573 25823
rect 30573 25789 30607 25823
rect 30607 25789 30616 25823
rect 30564 25780 30616 25789
rect 33876 25780 33928 25832
rect 34060 25823 34112 25832
rect 34060 25789 34069 25823
rect 34069 25789 34103 25823
rect 34103 25789 34112 25823
rect 34060 25780 34112 25789
rect 35440 25823 35492 25832
rect 35440 25789 35449 25823
rect 35449 25789 35483 25823
rect 35483 25789 35492 25823
rect 35440 25780 35492 25789
rect 37556 25823 37608 25832
rect 37556 25789 37565 25823
rect 37565 25789 37599 25823
rect 37599 25789 37608 25823
rect 37556 25780 37608 25789
rect 26884 25644 26936 25696
rect 33968 25644 34020 25696
rect 35808 25644 35860 25696
rect 37924 25644 37976 25696
rect 19606 25542 19658 25594
rect 19670 25542 19722 25594
rect 19734 25542 19786 25594
rect 19798 25542 19850 25594
rect 5724 25483 5776 25492
rect 5724 25449 5733 25483
rect 5733 25449 5767 25483
rect 5767 25449 5776 25483
rect 5724 25440 5776 25449
rect 8116 25440 8168 25492
rect 9036 25483 9088 25492
rect 9036 25449 9045 25483
rect 9045 25449 9079 25483
rect 9079 25449 9088 25483
rect 9036 25440 9088 25449
rect 9496 25440 9548 25492
rect 9956 25440 10008 25492
rect 10600 25440 10652 25492
rect 11060 25440 11112 25492
rect 11244 25440 11296 25492
rect 4712 25372 4764 25424
rect 1492 25304 1544 25356
rect 1676 25347 1728 25356
rect 1676 25313 1685 25347
rect 1685 25313 1719 25347
rect 1719 25313 1728 25347
rect 1676 25304 1728 25313
rect 4620 25347 4672 25356
rect 4620 25313 4629 25347
rect 4629 25313 4663 25347
rect 4663 25313 4672 25347
rect 4620 25304 4672 25313
rect 4804 25304 4856 25356
rect 5632 25304 5684 25356
rect 6552 25347 6604 25356
rect 6552 25313 6561 25347
rect 6561 25313 6595 25347
rect 6595 25313 6604 25347
rect 6552 25304 6604 25313
rect 8852 25347 8904 25356
rect 8852 25313 8861 25347
rect 8861 25313 8895 25347
rect 8895 25313 8904 25347
rect 8852 25304 8904 25313
rect 9864 25347 9916 25356
rect 9864 25313 9873 25347
rect 9873 25313 9907 25347
rect 9907 25313 9916 25347
rect 9864 25304 9916 25313
rect 11152 25372 11204 25424
rect 10600 25347 10652 25356
rect 10600 25313 10609 25347
rect 10609 25313 10643 25347
rect 10643 25313 10652 25347
rect 10600 25304 10652 25313
rect 14280 25372 14332 25424
rect 12440 25304 12492 25356
rect 12808 25304 12860 25356
rect 13268 25347 13320 25356
rect 13268 25313 13277 25347
rect 13277 25313 13311 25347
rect 13311 25313 13320 25347
rect 13268 25304 13320 25313
rect 6920 25236 6972 25288
rect 7748 25236 7800 25288
rect 10692 25236 10744 25288
rect 11060 25236 11112 25288
rect 13452 25279 13504 25288
rect 13452 25245 13461 25279
rect 13461 25245 13495 25279
rect 13495 25245 13504 25279
rect 13452 25236 13504 25245
rect 14188 25304 14240 25356
rect 18052 25440 18104 25492
rect 18328 25415 18380 25424
rect 18328 25381 18337 25415
rect 18337 25381 18371 25415
rect 18371 25381 18380 25415
rect 18328 25372 18380 25381
rect 16120 25304 16172 25356
rect 17316 25304 17368 25356
rect 17868 25304 17920 25356
rect 18144 25304 18196 25356
rect 19156 25347 19208 25356
rect 19156 25313 19165 25347
rect 19165 25313 19199 25347
rect 19199 25313 19208 25347
rect 19156 25304 19208 25313
rect 20720 25372 20772 25424
rect 22008 25415 22060 25424
rect 22008 25381 22017 25415
rect 22017 25381 22051 25415
rect 22051 25381 22060 25415
rect 22008 25372 22060 25381
rect 20904 25347 20956 25356
rect 13820 25236 13872 25288
rect 15660 25236 15712 25288
rect 20904 25313 20913 25347
rect 20913 25313 20947 25347
rect 20947 25313 20956 25347
rect 20904 25304 20956 25313
rect 21088 25304 21140 25356
rect 21824 25347 21876 25356
rect 21824 25313 21833 25347
rect 21833 25313 21867 25347
rect 21867 25313 21876 25347
rect 21824 25304 21876 25313
rect 23940 25372 23992 25424
rect 28264 25415 28316 25424
rect 28264 25381 28273 25415
rect 28273 25381 28307 25415
rect 28307 25381 28316 25415
rect 28264 25372 28316 25381
rect 32404 25372 32456 25424
rect 23296 25347 23348 25356
rect 23296 25313 23305 25347
rect 23305 25313 23339 25347
rect 23339 25313 23348 25347
rect 23296 25304 23348 25313
rect 23756 25347 23808 25356
rect 23756 25313 23765 25347
rect 23765 25313 23799 25347
rect 23799 25313 23808 25347
rect 23756 25304 23808 25313
rect 23848 25304 23900 25356
rect 25044 25347 25096 25356
rect 25044 25313 25053 25347
rect 25053 25313 25087 25347
rect 25087 25313 25096 25347
rect 25044 25304 25096 25313
rect 25228 25304 25280 25356
rect 26608 25347 26660 25356
rect 26608 25313 26617 25347
rect 26617 25313 26651 25347
rect 26651 25313 26660 25347
rect 26608 25304 26660 25313
rect 27252 25304 27304 25356
rect 29552 25347 29604 25356
rect 29552 25313 29561 25347
rect 29561 25313 29595 25347
rect 29595 25313 29604 25347
rect 29552 25304 29604 25313
rect 30564 25347 30616 25356
rect 20812 25236 20864 25288
rect 22008 25236 22060 25288
rect 25872 25279 25924 25288
rect 25872 25245 25881 25279
rect 25881 25245 25915 25279
rect 25915 25245 25924 25279
rect 25872 25236 25924 25245
rect 28172 25236 28224 25288
rect 28356 25236 28408 25288
rect 29644 25279 29696 25288
rect 29644 25245 29653 25279
rect 29653 25245 29687 25279
rect 29687 25245 29696 25279
rect 29644 25236 29696 25245
rect 2780 25143 2832 25152
rect 2780 25109 2789 25143
rect 2789 25109 2823 25143
rect 2823 25109 2832 25143
rect 18880 25168 18932 25220
rect 22560 25168 22612 25220
rect 24952 25211 25004 25220
rect 2780 25100 2832 25109
rect 16672 25100 16724 25152
rect 16948 25100 17000 25152
rect 17040 25100 17092 25152
rect 17316 25100 17368 25152
rect 22192 25100 22244 25152
rect 24492 25100 24544 25152
rect 24952 25177 24961 25211
rect 24961 25177 24995 25211
rect 24995 25177 25004 25211
rect 24952 25168 25004 25177
rect 30564 25313 30573 25347
rect 30573 25313 30607 25347
rect 30607 25313 30616 25347
rect 30564 25304 30616 25313
rect 30748 25347 30800 25356
rect 30748 25313 30757 25347
rect 30757 25313 30791 25347
rect 30791 25313 30800 25347
rect 30748 25304 30800 25313
rect 31852 25304 31904 25356
rect 34060 25440 34112 25492
rect 35440 25483 35492 25492
rect 35440 25449 35449 25483
rect 35449 25449 35483 25483
rect 35483 25449 35492 25483
rect 35440 25440 35492 25449
rect 32680 25347 32732 25356
rect 32680 25313 32689 25347
rect 32689 25313 32723 25347
rect 32723 25313 32732 25347
rect 32680 25304 32732 25313
rect 32496 25236 32548 25288
rect 33140 25304 33192 25356
rect 35532 25347 35584 25356
rect 35532 25313 35541 25347
rect 35541 25313 35575 25347
rect 35575 25313 35584 25347
rect 35532 25304 35584 25313
rect 36084 25347 36136 25356
rect 36084 25313 36093 25347
rect 36093 25313 36127 25347
rect 36127 25313 36136 25347
rect 36084 25304 36136 25313
rect 25504 25100 25556 25152
rect 30748 25100 30800 25152
rect 35900 25236 35952 25288
rect 38476 25304 38528 25356
rect 38752 25347 38804 25356
rect 38752 25313 38761 25347
rect 38761 25313 38795 25347
rect 38795 25313 38804 25347
rect 38752 25304 38804 25313
rect 39120 25304 39172 25356
rect 37740 25236 37792 25288
rect 38384 25236 38436 25288
rect 38844 25279 38896 25288
rect 38844 25245 38853 25279
rect 38853 25245 38887 25279
rect 38887 25245 38896 25279
rect 38844 25236 38896 25245
rect 33968 25168 34020 25220
rect 38292 25211 38344 25220
rect 38292 25177 38301 25211
rect 38301 25177 38335 25211
rect 38335 25177 38344 25211
rect 38292 25168 38344 25177
rect 36084 25100 36136 25152
rect 37096 25143 37148 25152
rect 37096 25109 37105 25143
rect 37105 25109 37139 25143
rect 37139 25109 37148 25143
rect 37096 25100 37148 25109
rect 4246 24998 4298 25050
rect 4310 24998 4362 25050
rect 4374 24998 4426 25050
rect 4438 24998 4490 25050
rect 34966 24998 35018 25050
rect 35030 24998 35082 25050
rect 35094 24998 35146 25050
rect 35158 24998 35210 25050
rect 22744 24896 22796 24948
rect 23848 24939 23900 24948
rect 23848 24905 23857 24939
rect 23857 24905 23891 24939
rect 23891 24905 23900 24939
rect 23848 24896 23900 24905
rect 23940 24896 23992 24948
rect 27988 24896 28040 24948
rect 2412 24828 2464 24880
rect 5724 24828 5776 24880
rect 20352 24871 20404 24880
rect 20352 24837 20361 24871
rect 20361 24837 20395 24871
rect 20395 24837 20404 24871
rect 20352 24828 20404 24837
rect 3976 24760 4028 24812
rect 2780 24692 2832 24744
rect 2964 24735 3016 24744
rect 2964 24701 2973 24735
rect 2973 24701 3007 24735
rect 3007 24701 3016 24735
rect 2964 24692 3016 24701
rect 3240 24735 3292 24744
rect 3240 24701 3249 24735
rect 3249 24701 3283 24735
rect 3283 24701 3292 24735
rect 3240 24692 3292 24701
rect 3608 24692 3660 24744
rect 3700 24735 3752 24744
rect 3700 24701 3709 24735
rect 3709 24701 3743 24735
rect 3743 24701 3752 24735
rect 4068 24735 4120 24744
rect 3700 24692 3752 24701
rect 4068 24701 4077 24735
rect 4077 24701 4111 24735
rect 4111 24701 4120 24735
rect 4068 24692 4120 24701
rect 5632 24692 5684 24744
rect 7564 24760 7616 24812
rect 7932 24760 7984 24812
rect 13636 24760 13688 24812
rect 15660 24803 15712 24812
rect 15660 24769 15669 24803
rect 15669 24769 15703 24803
rect 15703 24769 15712 24803
rect 15660 24760 15712 24769
rect 19156 24760 19208 24812
rect 7104 24735 7156 24744
rect 7104 24701 7113 24735
rect 7113 24701 7147 24735
rect 7147 24701 7156 24735
rect 7104 24692 7156 24701
rect 7656 24735 7708 24744
rect 7656 24701 7665 24735
rect 7665 24701 7699 24735
rect 7699 24701 7708 24735
rect 7656 24692 7708 24701
rect 8760 24735 8812 24744
rect 6184 24624 6236 24676
rect 6920 24599 6972 24608
rect 6920 24565 6929 24599
rect 6929 24565 6963 24599
rect 6963 24565 6972 24599
rect 6920 24556 6972 24565
rect 8760 24701 8769 24735
rect 8769 24701 8803 24735
rect 8803 24701 8812 24735
rect 8760 24692 8812 24701
rect 11060 24692 11112 24744
rect 11244 24692 11296 24744
rect 13544 24692 13596 24744
rect 14004 24735 14056 24744
rect 14004 24701 14013 24735
rect 14013 24701 14047 24735
rect 14047 24701 14056 24735
rect 14004 24692 14056 24701
rect 15384 24692 15436 24744
rect 18328 24692 18380 24744
rect 20536 24760 20588 24812
rect 21916 24828 21968 24880
rect 22836 24828 22888 24880
rect 29460 24828 29512 24880
rect 21824 24760 21876 24812
rect 20168 24735 20220 24744
rect 11152 24624 11204 24676
rect 11980 24624 12032 24676
rect 12808 24667 12860 24676
rect 12808 24633 12817 24667
rect 12817 24633 12851 24667
rect 12851 24633 12860 24667
rect 12808 24624 12860 24633
rect 16580 24624 16632 24676
rect 20168 24701 20177 24735
rect 20177 24701 20211 24735
rect 20211 24701 20220 24735
rect 20168 24692 20220 24701
rect 19156 24624 19208 24676
rect 21732 24692 21784 24744
rect 22652 24692 22704 24744
rect 23480 24760 23532 24812
rect 24952 24760 25004 24812
rect 25780 24760 25832 24812
rect 26516 24760 26568 24812
rect 27252 24760 27304 24812
rect 24400 24692 24452 24744
rect 24584 24692 24636 24744
rect 30564 24760 30616 24812
rect 31024 24760 31076 24812
rect 33140 24760 33192 24812
rect 35900 24760 35952 24812
rect 37556 24760 37608 24812
rect 9680 24556 9732 24608
rect 9956 24556 10008 24608
rect 10692 24556 10744 24608
rect 11244 24556 11296 24608
rect 11336 24556 11388 24608
rect 13268 24556 13320 24608
rect 16120 24556 16172 24608
rect 18788 24599 18840 24608
rect 18788 24565 18797 24599
rect 18797 24565 18831 24599
rect 18831 24565 18840 24599
rect 18788 24556 18840 24565
rect 26884 24624 26936 24676
rect 27436 24556 27488 24608
rect 29276 24692 29328 24744
rect 30012 24692 30064 24744
rect 30840 24692 30892 24744
rect 31116 24735 31168 24744
rect 31116 24701 31125 24735
rect 31125 24701 31159 24735
rect 31159 24701 31168 24735
rect 31116 24692 31168 24701
rect 31852 24692 31904 24744
rect 28540 24624 28592 24676
rect 30104 24667 30156 24676
rect 30104 24633 30113 24667
rect 30113 24633 30147 24667
rect 30147 24633 30156 24667
rect 30104 24624 30156 24633
rect 31576 24624 31628 24676
rect 33324 24692 33376 24744
rect 34060 24735 34112 24744
rect 34060 24701 34069 24735
rect 34069 24701 34103 24735
rect 34103 24701 34112 24735
rect 34060 24692 34112 24701
rect 35348 24692 35400 24744
rect 35624 24692 35676 24744
rect 35808 24692 35860 24744
rect 36912 24692 36964 24744
rect 37280 24692 37332 24744
rect 37464 24735 37516 24744
rect 37464 24701 37473 24735
rect 37473 24701 37507 24735
rect 37507 24701 37516 24735
rect 37464 24692 37516 24701
rect 35256 24624 35308 24676
rect 32772 24556 32824 24608
rect 33048 24556 33100 24608
rect 35440 24556 35492 24608
rect 38568 24599 38620 24608
rect 38568 24565 38577 24599
rect 38577 24565 38611 24599
rect 38611 24565 38620 24599
rect 38568 24556 38620 24565
rect 19606 24454 19658 24506
rect 19670 24454 19722 24506
rect 19734 24454 19786 24506
rect 19798 24454 19850 24506
rect 1860 24395 1912 24404
rect 1860 24361 1869 24395
rect 1869 24361 1903 24395
rect 1903 24361 1912 24395
rect 1860 24352 1912 24361
rect 7104 24352 7156 24404
rect 8760 24352 8812 24404
rect 7748 24284 7800 24336
rect 11152 24352 11204 24404
rect 15384 24395 15436 24404
rect 1768 24259 1820 24268
rect 1768 24225 1777 24259
rect 1777 24225 1811 24259
rect 1811 24225 1820 24259
rect 1768 24216 1820 24225
rect 2596 24259 2648 24268
rect 2596 24225 2605 24259
rect 2605 24225 2639 24259
rect 2639 24225 2648 24259
rect 2596 24216 2648 24225
rect 3332 24259 3384 24268
rect 3332 24225 3341 24259
rect 3341 24225 3375 24259
rect 3375 24225 3384 24259
rect 3332 24216 3384 24225
rect 3976 24216 4028 24268
rect 7104 24259 7156 24268
rect 7104 24225 7113 24259
rect 7113 24225 7147 24259
rect 7147 24225 7156 24259
rect 7104 24216 7156 24225
rect 9036 24259 9088 24268
rect 9036 24225 9045 24259
rect 9045 24225 9079 24259
rect 9079 24225 9088 24259
rect 9036 24216 9088 24225
rect 11980 24284 12032 24336
rect 11060 24216 11112 24268
rect 4804 24148 4856 24200
rect 4988 24191 5040 24200
rect 4988 24157 4997 24191
rect 4997 24157 5031 24191
rect 5031 24157 5040 24191
rect 4988 24148 5040 24157
rect 11244 24216 11296 24268
rect 11888 24259 11940 24268
rect 11888 24225 11897 24259
rect 11897 24225 11931 24259
rect 11931 24225 11940 24259
rect 11888 24216 11940 24225
rect 12256 24259 12308 24268
rect 12256 24225 12265 24259
rect 12265 24225 12299 24259
rect 12299 24225 12308 24259
rect 12256 24216 12308 24225
rect 13452 24259 13504 24268
rect 13452 24225 13461 24259
rect 13461 24225 13495 24259
rect 13495 24225 13504 24259
rect 13452 24216 13504 24225
rect 13912 24259 13964 24268
rect 13912 24225 13921 24259
rect 13921 24225 13955 24259
rect 13955 24225 13964 24259
rect 13912 24216 13964 24225
rect 15384 24361 15393 24395
rect 15393 24361 15427 24395
rect 15427 24361 15436 24395
rect 15384 24352 15436 24361
rect 15844 24284 15896 24336
rect 20352 24352 20404 24404
rect 20904 24352 20956 24404
rect 22100 24352 22152 24404
rect 18972 24284 19024 24336
rect 19156 24284 19208 24336
rect 22192 24284 22244 24336
rect 23848 24352 23900 24404
rect 24308 24395 24360 24404
rect 24308 24361 24317 24395
rect 24317 24361 24351 24395
rect 24351 24361 24360 24395
rect 24308 24352 24360 24361
rect 27620 24352 27672 24404
rect 31024 24352 31076 24404
rect 17776 24259 17828 24268
rect 16672 24148 16724 24200
rect 17776 24225 17785 24259
rect 17785 24225 17819 24259
rect 17819 24225 17828 24259
rect 17776 24216 17828 24225
rect 18328 24259 18380 24268
rect 18328 24225 18337 24259
rect 18337 24225 18371 24259
rect 18371 24225 18380 24259
rect 18328 24216 18380 24225
rect 18788 24216 18840 24268
rect 19064 24259 19116 24268
rect 19064 24225 19073 24259
rect 19073 24225 19107 24259
rect 19107 24225 19116 24259
rect 19064 24216 19116 24225
rect 19524 24216 19576 24268
rect 20260 24216 20312 24268
rect 20904 24259 20956 24268
rect 20904 24225 20913 24259
rect 20913 24225 20947 24259
rect 20947 24225 20956 24259
rect 20904 24216 20956 24225
rect 21732 24259 21784 24268
rect 21732 24225 21741 24259
rect 21741 24225 21775 24259
rect 21775 24225 21784 24259
rect 21732 24216 21784 24225
rect 22652 24216 22704 24268
rect 23848 24259 23900 24268
rect 18696 24148 18748 24200
rect 20168 24148 20220 24200
rect 23848 24225 23857 24259
rect 23857 24225 23891 24259
rect 23891 24225 23900 24259
rect 23848 24216 23900 24225
rect 25596 24284 25648 24336
rect 25964 24284 26016 24336
rect 26516 24216 26568 24268
rect 27160 24191 27212 24200
rect 27160 24157 27169 24191
rect 27169 24157 27203 24191
rect 27203 24157 27212 24191
rect 27160 24148 27212 24157
rect 28356 24259 28408 24268
rect 28356 24225 28365 24259
rect 28365 24225 28399 24259
rect 28399 24225 28408 24259
rect 28356 24216 28408 24225
rect 28540 24259 28592 24268
rect 28540 24225 28549 24259
rect 28549 24225 28583 24259
rect 28583 24225 28592 24259
rect 28540 24216 28592 24225
rect 27896 24148 27948 24200
rect 29460 24148 29512 24200
rect 36268 24284 36320 24336
rect 36452 24284 36504 24336
rect 30104 24259 30156 24268
rect 30104 24225 30113 24259
rect 30113 24225 30147 24259
rect 30147 24225 30156 24259
rect 30104 24216 30156 24225
rect 31852 24216 31904 24268
rect 32128 24216 32180 24268
rect 32588 24216 32640 24268
rect 33324 24259 33376 24268
rect 33324 24225 33333 24259
rect 33333 24225 33367 24259
rect 33367 24225 33376 24259
rect 36360 24259 36412 24268
rect 33324 24216 33376 24225
rect 30288 24148 30340 24200
rect 32496 24148 32548 24200
rect 33968 24191 34020 24200
rect 33968 24157 33977 24191
rect 33977 24157 34011 24191
rect 34011 24157 34020 24191
rect 33968 24148 34020 24157
rect 34244 24191 34296 24200
rect 34244 24157 34253 24191
rect 34253 24157 34287 24191
rect 34287 24157 34296 24191
rect 34244 24148 34296 24157
rect 36360 24225 36369 24259
rect 36369 24225 36403 24259
rect 36403 24225 36412 24259
rect 36360 24216 36412 24225
rect 38292 24259 38344 24268
rect 36452 24191 36504 24200
rect 36452 24157 36461 24191
rect 36461 24157 36495 24191
rect 36495 24157 36504 24191
rect 36452 24148 36504 24157
rect 38292 24225 38301 24259
rect 38301 24225 38335 24259
rect 38335 24225 38344 24259
rect 38292 24216 38344 24225
rect 38936 24259 38988 24268
rect 38936 24225 38945 24259
rect 38945 24225 38979 24259
rect 38979 24225 38988 24259
rect 38936 24216 38988 24225
rect 38108 24148 38160 24200
rect 18328 24080 18380 24132
rect 22284 24080 22336 24132
rect 27528 24080 27580 24132
rect 33140 24123 33192 24132
rect 33140 24089 33149 24123
rect 33149 24089 33183 24123
rect 33183 24089 33192 24123
rect 33140 24080 33192 24089
rect 37464 24080 37516 24132
rect 3424 24055 3476 24064
rect 3424 24021 3433 24055
rect 3433 24021 3467 24055
rect 3467 24021 3476 24055
rect 3424 24012 3476 24021
rect 4620 24012 4672 24064
rect 5632 24012 5684 24064
rect 6828 24012 6880 24064
rect 9956 24012 10008 24064
rect 14004 24012 14056 24064
rect 22468 24012 22520 24064
rect 23112 24012 23164 24064
rect 31484 24012 31536 24064
rect 4246 23910 4298 23962
rect 4310 23910 4362 23962
rect 4374 23910 4426 23962
rect 4438 23910 4490 23962
rect 34966 23910 35018 23962
rect 35030 23910 35082 23962
rect 35094 23910 35146 23962
rect 35158 23910 35210 23962
rect 7748 23851 7800 23860
rect 7748 23817 7757 23851
rect 7757 23817 7791 23851
rect 7791 23817 7800 23851
rect 7748 23808 7800 23817
rect 8024 23808 8076 23860
rect 15476 23808 15528 23860
rect 2596 23783 2648 23792
rect 2596 23749 2605 23783
rect 2605 23749 2639 23783
rect 2639 23749 2648 23783
rect 2596 23740 2648 23749
rect 3700 23740 3752 23792
rect 7104 23740 7156 23792
rect 11888 23740 11940 23792
rect 15292 23740 15344 23792
rect 2964 23672 3016 23724
rect 9680 23715 9732 23724
rect 9680 23681 9689 23715
rect 9689 23681 9723 23715
rect 9723 23681 9732 23715
rect 9680 23672 9732 23681
rect 3240 23647 3292 23656
rect 3240 23613 3249 23647
rect 3249 23613 3283 23647
rect 3283 23613 3292 23647
rect 3240 23604 3292 23613
rect 3976 23604 4028 23656
rect 5724 23647 5776 23656
rect 5724 23613 5733 23647
rect 5733 23613 5767 23647
rect 5767 23613 5776 23647
rect 5724 23604 5776 23613
rect 6184 23647 6236 23656
rect 6184 23613 6193 23647
rect 6193 23613 6227 23647
rect 6227 23613 6236 23647
rect 6184 23604 6236 23613
rect 7840 23604 7892 23656
rect 6828 23536 6880 23588
rect 9036 23604 9088 23656
rect 9772 23604 9824 23656
rect 11152 23604 11204 23656
rect 14004 23715 14056 23724
rect 10508 23536 10560 23588
rect 12072 23604 12124 23656
rect 12624 23647 12676 23656
rect 12624 23613 12633 23647
rect 12633 23613 12667 23647
rect 12667 23613 12676 23647
rect 12624 23604 12676 23613
rect 14004 23681 14013 23715
rect 14013 23681 14047 23715
rect 14047 23681 14056 23715
rect 14004 23672 14056 23681
rect 13728 23604 13780 23656
rect 14556 23604 14608 23656
rect 12256 23536 12308 23588
rect 15200 23536 15252 23588
rect 1492 23468 1544 23520
rect 4988 23468 5040 23520
rect 11060 23511 11112 23520
rect 11060 23477 11069 23511
rect 11069 23477 11103 23511
rect 11103 23477 11112 23511
rect 11060 23468 11112 23477
rect 12992 23468 13044 23520
rect 17592 23808 17644 23860
rect 18880 23808 18932 23860
rect 18328 23715 18380 23724
rect 18328 23681 18337 23715
rect 18337 23681 18371 23715
rect 18371 23681 18380 23715
rect 18328 23672 18380 23681
rect 19524 23808 19576 23860
rect 21180 23808 21232 23860
rect 29552 23808 29604 23860
rect 32680 23808 32732 23860
rect 34520 23808 34572 23860
rect 34704 23808 34756 23860
rect 38936 23808 38988 23860
rect 20168 23740 20220 23792
rect 18696 23647 18748 23656
rect 18696 23613 18705 23647
rect 18705 23613 18739 23647
rect 18739 23613 18748 23647
rect 18696 23604 18748 23613
rect 18788 23604 18840 23656
rect 19156 23604 19208 23656
rect 20536 23647 20588 23656
rect 20536 23613 20545 23647
rect 20545 23613 20579 23647
rect 20579 23613 20588 23647
rect 20536 23604 20588 23613
rect 20812 23647 20864 23656
rect 20812 23613 20821 23647
rect 20821 23613 20855 23647
rect 20855 23613 20864 23647
rect 20812 23604 20864 23613
rect 20904 23604 20956 23656
rect 21732 23604 21784 23656
rect 22100 23672 22152 23724
rect 22744 23672 22796 23724
rect 22652 23647 22704 23656
rect 22652 23613 22661 23647
rect 22661 23613 22695 23647
rect 22695 23613 22704 23647
rect 22652 23604 22704 23613
rect 23664 23672 23716 23724
rect 27896 23740 27948 23792
rect 27344 23672 27396 23724
rect 23848 23647 23900 23656
rect 23848 23613 23857 23647
rect 23857 23613 23891 23647
rect 23891 23613 23900 23647
rect 23848 23604 23900 23613
rect 24400 23647 24452 23656
rect 22284 23536 22336 23588
rect 24400 23613 24409 23647
rect 24409 23613 24443 23647
rect 24443 23613 24452 23647
rect 24400 23604 24452 23613
rect 25780 23604 25832 23656
rect 26240 23647 26292 23656
rect 26240 23613 26249 23647
rect 26249 23613 26283 23647
rect 26283 23613 26292 23647
rect 26240 23604 26292 23613
rect 26700 23604 26752 23656
rect 26884 23604 26936 23656
rect 27896 23647 27948 23656
rect 27896 23613 27905 23647
rect 27905 23613 27939 23647
rect 27939 23613 27948 23647
rect 27896 23604 27948 23613
rect 28448 23604 28500 23656
rect 31116 23672 31168 23724
rect 32496 23740 32548 23792
rect 32588 23740 32640 23792
rect 31576 23672 31628 23724
rect 33140 23672 33192 23724
rect 31668 23647 31720 23656
rect 28356 23536 28408 23588
rect 31668 23613 31677 23647
rect 31677 23613 31711 23647
rect 31711 23613 31720 23647
rect 31668 23604 31720 23613
rect 33232 23604 33284 23656
rect 33968 23740 34020 23792
rect 37280 23672 37332 23724
rect 27712 23468 27764 23520
rect 28448 23468 28500 23520
rect 30288 23511 30340 23520
rect 30288 23477 30297 23511
rect 30297 23477 30331 23511
rect 30331 23477 30340 23511
rect 30288 23468 30340 23477
rect 31484 23536 31536 23588
rect 32588 23536 32640 23588
rect 32772 23536 32824 23588
rect 34152 23604 34204 23656
rect 35992 23604 36044 23656
rect 37740 23647 37792 23656
rect 37740 23613 37749 23647
rect 37749 23613 37783 23647
rect 37783 23613 37792 23647
rect 37740 23604 37792 23613
rect 32036 23468 32088 23520
rect 34060 23468 34112 23520
rect 36360 23468 36412 23520
rect 19606 23366 19658 23418
rect 19670 23366 19722 23418
rect 19734 23366 19786 23418
rect 19798 23366 19850 23418
rect 5448 23264 5500 23316
rect 7840 23264 7892 23316
rect 9772 23307 9824 23316
rect 3976 23196 4028 23248
rect 1492 23171 1544 23180
rect 1492 23137 1501 23171
rect 1501 23137 1535 23171
rect 1535 23137 1544 23171
rect 1492 23128 1544 23137
rect 1860 23128 1912 23180
rect 3424 23128 3476 23180
rect 4896 23171 4948 23180
rect 4896 23137 4905 23171
rect 4905 23137 4939 23171
rect 4939 23137 4948 23171
rect 4896 23128 4948 23137
rect 5080 23171 5132 23180
rect 5080 23137 5089 23171
rect 5089 23137 5123 23171
rect 5123 23137 5132 23171
rect 5080 23128 5132 23137
rect 6000 23171 6052 23180
rect 6000 23137 6009 23171
rect 6009 23137 6043 23171
rect 6043 23137 6052 23171
rect 6000 23128 6052 23137
rect 6644 23128 6696 23180
rect 7380 23128 7432 23180
rect 7840 23171 7892 23180
rect 7840 23137 7849 23171
rect 7849 23137 7883 23171
rect 7883 23137 7892 23171
rect 7840 23128 7892 23137
rect 8668 23128 8720 23180
rect 9772 23273 9781 23307
rect 9781 23273 9815 23307
rect 9815 23273 9824 23307
rect 9772 23264 9824 23273
rect 10600 23264 10652 23316
rect 9036 23196 9088 23248
rect 19432 23264 19484 23316
rect 21456 23264 21508 23316
rect 21732 23264 21784 23316
rect 22560 23264 22612 23316
rect 24400 23264 24452 23316
rect 26240 23264 26292 23316
rect 28172 23307 28224 23316
rect 28172 23273 28181 23307
rect 28181 23273 28215 23307
rect 28215 23273 28224 23307
rect 28172 23264 28224 23273
rect 30840 23307 30892 23316
rect 30840 23273 30849 23307
rect 30849 23273 30883 23307
rect 30883 23273 30892 23307
rect 30840 23264 30892 23273
rect 32220 23307 32272 23316
rect 32220 23273 32229 23307
rect 32229 23273 32263 23307
rect 32263 23273 32272 23307
rect 32220 23264 32272 23273
rect 33692 23307 33744 23316
rect 33692 23273 33701 23307
rect 33701 23273 33735 23307
rect 33735 23273 33744 23307
rect 33692 23264 33744 23273
rect 33968 23264 34020 23316
rect 35992 23264 36044 23316
rect 9404 23128 9456 23180
rect 10508 23171 10560 23180
rect 10508 23137 10517 23171
rect 10517 23137 10551 23171
rect 10551 23137 10560 23171
rect 10508 23128 10560 23137
rect 11428 23128 11480 23180
rect 12072 23171 12124 23180
rect 12072 23137 12081 23171
rect 12081 23137 12115 23171
rect 12115 23137 12124 23171
rect 12072 23128 12124 23137
rect 12348 23171 12400 23180
rect 12348 23137 12357 23171
rect 12357 23137 12391 23171
rect 12391 23137 12400 23171
rect 12348 23128 12400 23137
rect 13728 23171 13780 23180
rect 13728 23137 13737 23171
rect 13737 23137 13771 23171
rect 13771 23137 13780 23171
rect 13728 23128 13780 23137
rect 6736 23103 6788 23112
rect 6736 23069 6745 23103
rect 6745 23069 6779 23103
rect 6779 23069 6788 23103
rect 6736 23060 6788 23069
rect 12440 23103 12492 23112
rect 12440 23069 12449 23103
rect 12449 23069 12483 23103
rect 12483 23069 12492 23103
rect 12440 23060 12492 23069
rect 13176 23103 13228 23112
rect 13176 23069 13185 23103
rect 13185 23069 13219 23103
rect 13219 23069 13228 23103
rect 13176 23060 13228 23069
rect 14188 23128 14240 23180
rect 15292 23128 15344 23180
rect 16488 23171 16540 23180
rect 15200 23060 15252 23112
rect 16120 23103 16172 23112
rect 16120 23069 16129 23103
rect 16129 23069 16163 23103
rect 16163 23069 16172 23103
rect 16120 23060 16172 23069
rect 16488 23137 16497 23171
rect 16497 23137 16531 23171
rect 16531 23137 16540 23171
rect 16488 23128 16540 23137
rect 16580 23128 16632 23180
rect 16672 23171 16724 23180
rect 16672 23137 16681 23171
rect 16681 23137 16715 23171
rect 16715 23137 16724 23171
rect 16672 23128 16724 23137
rect 17224 23128 17276 23180
rect 17868 23128 17920 23180
rect 18604 23171 18656 23180
rect 18604 23137 18613 23171
rect 18613 23137 18647 23171
rect 18647 23137 18656 23171
rect 18604 23128 18656 23137
rect 18788 23171 18840 23180
rect 18788 23137 18797 23171
rect 18797 23137 18831 23171
rect 18831 23137 18840 23171
rect 18788 23128 18840 23137
rect 19984 23196 20036 23248
rect 19156 23171 19208 23180
rect 19156 23137 19165 23171
rect 19165 23137 19199 23171
rect 19199 23137 19208 23171
rect 19156 23128 19208 23137
rect 22652 23196 22704 23248
rect 20904 23128 20956 23180
rect 18144 23060 18196 23112
rect 20720 23060 20772 23112
rect 21640 23103 21692 23112
rect 21640 23069 21649 23103
rect 21649 23069 21683 23103
rect 21683 23069 21692 23103
rect 21640 23060 21692 23069
rect 7196 22992 7248 23044
rect 21824 23128 21876 23180
rect 22284 23171 22336 23180
rect 22284 23137 22293 23171
rect 22293 23137 22327 23171
rect 22327 23137 22336 23171
rect 22284 23128 22336 23137
rect 5908 22924 5960 22976
rect 7472 22924 7524 22976
rect 11428 22924 11480 22976
rect 14188 22924 14240 22976
rect 16672 22924 16724 22976
rect 21364 22924 21416 22976
rect 23480 23128 23532 23180
rect 24216 23128 24268 23180
rect 27620 23196 27672 23248
rect 31760 23196 31812 23248
rect 25412 23128 25464 23180
rect 26424 23128 26476 23180
rect 27068 23128 27120 23180
rect 23572 23060 23624 23112
rect 23664 23060 23716 23112
rect 27528 23128 27580 23180
rect 28356 23128 28408 23180
rect 27252 23103 27304 23112
rect 27252 23069 27261 23103
rect 27261 23069 27295 23103
rect 27295 23069 27304 23103
rect 27252 23060 27304 23069
rect 30288 23128 30340 23180
rect 31668 23128 31720 23180
rect 31852 23128 31904 23180
rect 32128 23171 32180 23180
rect 32128 23137 32137 23171
rect 32137 23137 32171 23171
rect 32171 23137 32180 23171
rect 32128 23128 32180 23137
rect 32588 23171 32640 23180
rect 32588 23137 32597 23171
rect 32597 23137 32631 23171
rect 32631 23137 32640 23171
rect 32588 23128 32640 23137
rect 30472 23060 30524 23112
rect 32036 23060 32088 23112
rect 33508 23128 33560 23180
rect 34244 23196 34296 23248
rect 33232 23060 33284 23112
rect 35256 23128 35308 23180
rect 36360 23196 36412 23248
rect 36452 23171 36504 23180
rect 35440 23060 35492 23112
rect 28356 22992 28408 23044
rect 33324 22992 33376 23044
rect 36452 23137 36461 23171
rect 36461 23137 36495 23171
rect 36495 23137 36504 23171
rect 36452 23128 36504 23137
rect 38016 23171 38068 23180
rect 38016 23137 38025 23171
rect 38025 23137 38059 23171
rect 38059 23137 38068 23171
rect 38016 23128 38068 23137
rect 38292 23171 38344 23180
rect 38292 23137 38301 23171
rect 38301 23137 38335 23171
rect 38335 23137 38344 23171
rect 38292 23128 38344 23137
rect 36636 23103 36688 23112
rect 36636 23069 36645 23103
rect 36645 23069 36679 23103
rect 36679 23069 36688 23103
rect 36636 23060 36688 23069
rect 36820 23060 36872 23112
rect 37740 22992 37792 23044
rect 31760 22967 31812 22976
rect 31760 22933 31769 22967
rect 31769 22933 31803 22967
rect 31803 22933 31812 22967
rect 31760 22924 31812 22933
rect 35440 22924 35492 22976
rect 36544 22924 36596 22976
rect 39028 22967 39080 22976
rect 39028 22933 39037 22967
rect 39037 22933 39071 22967
rect 39071 22933 39080 22967
rect 39028 22924 39080 22933
rect 4246 22822 4298 22874
rect 4310 22822 4362 22874
rect 4374 22822 4426 22874
rect 4438 22822 4490 22874
rect 34966 22822 35018 22874
rect 35030 22822 35082 22874
rect 35094 22822 35146 22874
rect 35158 22822 35210 22874
rect 5080 22720 5132 22772
rect 12624 22720 12676 22772
rect 17224 22720 17276 22772
rect 18972 22763 19024 22772
rect 18972 22729 18981 22763
rect 18981 22729 19015 22763
rect 19015 22729 19024 22763
rect 18972 22720 19024 22729
rect 22284 22720 22336 22772
rect 26700 22720 26752 22772
rect 29000 22720 29052 22772
rect 29460 22720 29512 22772
rect 30472 22720 30524 22772
rect 32128 22720 32180 22772
rect 32404 22720 32456 22772
rect 36636 22720 36688 22772
rect 37004 22720 37056 22772
rect 4804 22652 4856 22704
rect 2320 22584 2372 22636
rect 2964 22627 3016 22636
rect 2964 22593 2973 22627
rect 2973 22593 3007 22627
rect 3007 22593 3016 22627
rect 2964 22584 3016 22593
rect 2688 22559 2740 22568
rect 2688 22525 2697 22559
rect 2697 22525 2731 22559
rect 2731 22525 2740 22559
rect 2688 22516 2740 22525
rect 3240 22516 3292 22568
rect 3424 22516 3476 22568
rect 4620 22584 4672 22636
rect 19892 22695 19944 22704
rect 19892 22661 19901 22695
rect 19901 22661 19935 22695
rect 19935 22661 19944 22695
rect 19892 22652 19944 22661
rect 4528 22559 4580 22568
rect 4528 22525 4537 22559
rect 4537 22525 4571 22559
rect 4571 22525 4580 22559
rect 4896 22559 4948 22568
rect 4528 22516 4580 22525
rect 4896 22525 4905 22559
rect 4905 22525 4939 22559
rect 4939 22525 4948 22559
rect 4896 22516 4948 22525
rect 5908 22584 5960 22636
rect 6184 22627 6236 22636
rect 6184 22593 6193 22627
rect 6193 22593 6227 22627
rect 6227 22593 6236 22627
rect 6184 22584 6236 22593
rect 5632 22516 5684 22568
rect 6000 22559 6052 22568
rect 6000 22525 6009 22559
rect 6009 22525 6043 22559
rect 6043 22525 6052 22559
rect 6000 22516 6052 22525
rect 6828 22559 6880 22568
rect 6828 22525 6837 22559
rect 6837 22525 6871 22559
rect 6871 22525 6880 22559
rect 6828 22516 6880 22525
rect 7380 22559 7432 22568
rect 7380 22525 7389 22559
rect 7389 22525 7423 22559
rect 7423 22525 7432 22559
rect 7380 22516 7432 22525
rect 8300 22559 8352 22568
rect 8300 22525 8309 22559
rect 8309 22525 8343 22559
rect 8343 22525 8352 22559
rect 8300 22516 8352 22525
rect 10600 22584 10652 22636
rect 13820 22627 13872 22636
rect 13820 22593 13829 22627
rect 13829 22593 13863 22627
rect 13863 22593 13872 22627
rect 13820 22584 13872 22593
rect 14004 22584 14056 22636
rect 14188 22584 14240 22636
rect 17500 22627 17552 22636
rect 9956 22516 10008 22568
rect 10416 22559 10468 22568
rect 10416 22525 10425 22559
rect 10425 22525 10459 22559
rect 10459 22525 10468 22559
rect 10416 22516 10468 22525
rect 11060 22516 11112 22568
rect 12992 22559 13044 22568
rect 12992 22525 13001 22559
rect 13001 22525 13035 22559
rect 13035 22525 13044 22559
rect 12992 22516 13044 22525
rect 15384 22516 15436 22568
rect 16120 22516 16172 22568
rect 16488 22516 16540 22568
rect 16672 22516 16724 22568
rect 17500 22593 17509 22627
rect 17509 22593 17543 22627
rect 17543 22593 17552 22627
rect 17500 22584 17552 22593
rect 17224 22516 17276 22568
rect 18052 22559 18104 22568
rect 18052 22525 18061 22559
rect 18061 22525 18095 22559
rect 18095 22525 18104 22559
rect 18052 22516 18104 22525
rect 18788 22559 18840 22568
rect 18788 22525 18797 22559
rect 18797 22525 18831 22559
rect 18831 22525 18840 22559
rect 18788 22516 18840 22525
rect 23940 22584 23992 22636
rect 25412 22584 25464 22636
rect 31576 22652 31628 22704
rect 35532 22652 35584 22704
rect 36360 22652 36412 22704
rect 27252 22584 27304 22636
rect 20260 22516 20312 22568
rect 20628 22559 20680 22568
rect 20628 22525 20637 22559
rect 20637 22525 20671 22559
rect 20671 22525 20680 22559
rect 20628 22516 20680 22525
rect 21364 22559 21416 22568
rect 21364 22525 21373 22559
rect 21373 22525 21407 22559
rect 21407 22525 21416 22559
rect 21364 22516 21416 22525
rect 21640 22559 21692 22568
rect 21640 22525 21649 22559
rect 21649 22525 21683 22559
rect 21683 22525 21692 22559
rect 21640 22516 21692 22525
rect 23664 22559 23716 22568
rect 23664 22525 23673 22559
rect 23673 22525 23707 22559
rect 23707 22525 23716 22559
rect 23664 22516 23716 22525
rect 24860 22559 24912 22568
rect 24860 22525 24869 22559
rect 24869 22525 24903 22559
rect 24903 22525 24912 22559
rect 24860 22516 24912 22525
rect 26424 22559 26476 22568
rect 7840 22448 7892 22500
rect 2964 22380 3016 22432
rect 12348 22380 12400 22432
rect 13728 22380 13780 22432
rect 17132 22448 17184 22500
rect 20076 22448 20128 22500
rect 24308 22448 24360 22500
rect 24584 22448 24636 22500
rect 26424 22525 26433 22559
rect 26433 22525 26467 22559
rect 26467 22525 26476 22559
rect 26424 22516 26476 22525
rect 24216 22380 24268 22432
rect 26792 22559 26844 22568
rect 26792 22525 26801 22559
rect 26801 22525 26835 22559
rect 26835 22525 26844 22559
rect 27068 22559 27120 22568
rect 26792 22516 26844 22525
rect 27068 22525 27077 22559
rect 27077 22525 27111 22559
rect 27111 22525 27120 22559
rect 27068 22516 27120 22525
rect 27160 22559 27212 22568
rect 27160 22525 27169 22559
rect 27169 22525 27203 22559
rect 27203 22525 27212 22559
rect 27160 22516 27212 22525
rect 28264 22516 28316 22568
rect 31760 22584 31812 22636
rect 32312 22627 32364 22636
rect 32312 22593 32321 22627
rect 32321 22593 32355 22627
rect 32355 22593 32364 22627
rect 32312 22584 32364 22593
rect 34060 22584 34112 22636
rect 34428 22584 34480 22636
rect 29460 22516 29512 22568
rect 29828 22559 29880 22568
rect 29828 22525 29837 22559
rect 29837 22525 29871 22559
rect 29871 22525 29880 22559
rect 29828 22516 29880 22525
rect 30288 22516 30340 22568
rect 32036 22559 32088 22568
rect 32036 22525 32045 22559
rect 32045 22525 32079 22559
rect 32079 22525 32088 22559
rect 32036 22516 32088 22525
rect 32404 22559 32456 22568
rect 32404 22525 32413 22559
rect 32413 22525 32447 22559
rect 32447 22525 32456 22559
rect 32404 22516 32456 22525
rect 32496 22516 32548 22568
rect 33600 22559 33652 22568
rect 33600 22525 33609 22559
rect 33609 22525 33643 22559
rect 33643 22525 33652 22559
rect 33600 22516 33652 22525
rect 35256 22516 35308 22568
rect 26976 22448 27028 22500
rect 33968 22448 34020 22500
rect 37280 22584 37332 22636
rect 37924 22627 37976 22636
rect 37924 22593 37933 22627
rect 37933 22593 37967 22627
rect 37967 22593 37976 22627
rect 37924 22584 37976 22593
rect 38292 22584 38344 22636
rect 36176 22559 36228 22568
rect 36176 22525 36185 22559
rect 36185 22525 36219 22559
rect 36219 22525 36228 22559
rect 36176 22516 36228 22525
rect 27620 22380 27672 22432
rect 27896 22380 27948 22432
rect 28540 22380 28592 22432
rect 31024 22380 31076 22432
rect 31668 22380 31720 22432
rect 33784 22380 33836 22432
rect 35532 22380 35584 22432
rect 38108 22559 38160 22568
rect 38108 22525 38117 22559
rect 38117 22525 38151 22559
rect 38151 22525 38160 22559
rect 38108 22516 38160 22525
rect 38568 22516 38620 22568
rect 37188 22448 37240 22500
rect 37372 22380 37424 22432
rect 19606 22278 19658 22330
rect 19670 22278 19722 22330
rect 19734 22278 19786 22330
rect 19798 22278 19850 22330
rect 2320 22176 2372 22228
rect 3240 22176 3292 22228
rect 7380 22219 7432 22228
rect 7380 22185 7389 22219
rect 7389 22185 7423 22219
rect 7423 22185 7432 22219
rect 7380 22176 7432 22185
rect 8300 22219 8352 22228
rect 8300 22185 8309 22219
rect 8309 22185 8343 22219
rect 8343 22185 8352 22219
rect 8300 22176 8352 22185
rect 10416 22176 10468 22228
rect 11428 22219 11480 22228
rect 11428 22185 11437 22219
rect 11437 22185 11471 22219
rect 11471 22185 11480 22219
rect 11428 22176 11480 22185
rect 14188 22176 14240 22228
rect 15292 22176 15344 22228
rect 18972 22176 19024 22228
rect 19156 22176 19208 22228
rect 25320 22219 25372 22228
rect 25320 22185 25329 22219
rect 25329 22185 25363 22219
rect 25363 22185 25372 22219
rect 25320 22176 25372 22185
rect 27528 22176 27580 22228
rect 29828 22219 29880 22228
rect 29828 22185 29837 22219
rect 29837 22185 29871 22219
rect 29871 22185 29880 22219
rect 29828 22176 29880 22185
rect 33232 22176 33284 22228
rect 37832 22219 37884 22228
rect 37832 22185 37841 22219
rect 37841 22185 37875 22219
rect 37875 22185 37884 22219
rect 37832 22176 37884 22185
rect 2320 22083 2372 22092
rect 2320 22049 2329 22083
rect 2329 22049 2363 22083
rect 2363 22049 2372 22083
rect 2320 22040 2372 22049
rect 2688 22083 2740 22092
rect 2688 22049 2697 22083
rect 2697 22049 2731 22083
rect 2731 22049 2740 22083
rect 2688 22040 2740 22049
rect 2964 22083 3016 22092
rect 2964 22049 2973 22083
rect 2973 22049 3007 22083
rect 3007 22049 3016 22083
rect 2964 22040 3016 22049
rect 4528 22083 4580 22092
rect 4528 22049 4537 22083
rect 4537 22049 4571 22083
rect 4571 22049 4580 22083
rect 4528 22040 4580 22049
rect 4988 22040 5040 22092
rect 8024 22083 8076 22092
rect 8024 22049 8033 22083
rect 8033 22049 8067 22083
rect 8067 22049 8076 22083
rect 8024 22040 8076 22049
rect 8852 22083 8904 22092
rect 8852 22049 8861 22083
rect 8861 22049 8895 22083
rect 8895 22049 8904 22083
rect 8852 22040 8904 22049
rect 9036 22083 9088 22092
rect 9036 22049 9045 22083
rect 9045 22049 9079 22083
rect 9079 22049 9088 22083
rect 9036 22040 9088 22049
rect 9680 22083 9732 22092
rect 9680 22049 9689 22083
rect 9689 22049 9723 22083
rect 9723 22049 9732 22083
rect 9680 22040 9732 22049
rect 9956 22040 10008 22092
rect 10600 22083 10652 22092
rect 10600 22049 10609 22083
rect 10609 22049 10643 22083
rect 10643 22049 10652 22083
rect 10600 22040 10652 22049
rect 11060 22040 11112 22092
rect 12624 22108 12676 22160
rect 15200 22108 15252 22160
rect 12440 22083 12492 22092
rect 12440 22049 12449 22083
rect 12449 22049 12483 22083
rect 12483 22049 12492 22083
rect 12440 22040 12492 22049
rect 12532 22040 12584 22092
rect 13176 22083 13228 22092
rect 13176 22049 13185 22083
rect 13185 22049 13219 22083
rect 13219 22049 13228 22083
rect 13176 22040 13228 22049
rect 14188 22083 14240 22092
rect 14188 22049 14197 22083
rect 14197 22049 14231 22083
rect 14231 22049 14240 22083
rect 14188 22040 14240 22049
rect 14556 22083 14608 22092
rect 14556 22049 14565 22083
rect 14565 22049 14599 22083
rect 14599 22049 14608 22083
rect 14556 22040 14608 22049
rect 5540 21972 5592 22024
rect 6920 21972 6972 22024
rect 7196 21972 7248 22024
rect 1860 21904 1912 21956
rect 12164 21904 12216 21956
rect 13728 21972 13780 22024
rect 17868 22108 17920 22160
rect 18696 22108 18748 22160
rect 16764 22040 16816 22092
rect 16948 22083 17000 22092
rect 16948 22049 16957 22083
rect 16957 22049 16991 22083
rect 16991 22049 17000 22083
rect 16948 22040 17000 22049
rect 16580 21972 16632 22024
rect 17224 22040 17276 22092
rect 17592 22040 17644 22092
rect 17408 22015 17460 22024
rect 17408 21981 17417 22015
rect 17417 21981 17451 22015
rect 17451 21981 17460 22015
rect 17408 21972 17460 21981
rect 18972 21972 19024 22024
rect 19340 22040 19392 22092
rect 19892 22040 19944 22092
rect 26792 22108 26844 22160
rect 22652 22040 22704 22092
rect 23664 22083 23716 22092
rect 23664 22049 23673 22083
rect 23673 22049 23707 22083
rect 23707 22049 23716 22083
rect 23664 22040 23716 22049
rect 24308 22083 24360 22092
rect 24308 22049 24317 22083
rect 24317 22049 24351 22083
rect 24351 22049 24360 22083
rect 24308 22040 24360 22049
rect 25504 22083 25556 22092
rect 25504 22049 25513 22083
rect 25513 22049 25547 22083
rect 25547 22049 25556 22083
rect 25504 22040 25556 22049
rect 25688 22083 25740 22092
rect 25688 22049 25697 22083
rect 25697 22049 25731 22083
rect 25731 22049 25740 22083
rect 25688 22040 25740 22049
rect 26976 22083 27028 22092
rect 26976 22049 26985 22083
rect 26985 22049 27019 22083
rect 27019 22049 27028 22083
rect 26976 22040 27028 22049
rect 27068 22040 27120 22092
rect 27620 22108 27672 22160
rect 27712 22083 27764 22092
rect 27712 22049 27721 22083
rect 27721 22049 27755 22083
rect 27755 22049 27764 22083
rect 27712 22040 27764 22049
rect 28172 22040 28224 22092
rect 29092 22083 29144 22092
rect 29092 22049 29101 22083
rect 29101 22049 29135 22083
rect 29135 22049 29144 22083
rect 29092 22040 29144 22049
rect 29552 22040 29604 22092
rect 21180 22015 21232 22024
rect 15292 21904 15344 21956
rect 16488 21904 16540 21956
rect 21180 21981 21189 22015
rect 21189 21981 21223 22015
rect 21223 21981 21232 22015
rect 21180 21972 21232 21981
rect 21364 21972 21416 22024
rect 24124 21972 24176 22024
rect 30288 22040 30340 22092
rect 30840 22040 30892 22092
rect 32220 22108 32272 22160
rect 33692 22108 33744 22160
rect 34428 22108 34480 22160
rect 31392 22083 31444 22092
rect 31392 22049 31401 22083
rect 31401 22049 31435 22083
rect 31435 22049 31444 22083
rect 31392 22040 31444 22049
rect 32128 22040 32180 22092
rect 32772 22040 32824 22092
rect 33508 22040 33560 22092
rect 36820 22083 36872 22092
rect 33784 22015 33836 22024
rect 23848 21947 23900 21956
rect 23848 21913 23857 21947
rect 23857 21913 23891 21947
rect 23891 21913 23900 21947
rect 23848 21904 23900 21913
rect 3332 21836 3384 21888
rect 19340 21879 19392 21888
rect 19340 21845 19349 21879
rect 19349 21845 19383 21879
rect 19383 21845 19392 21879
rect 19340 21836 19392 21845
rect 20168 21836 20220 21888
rect 20536 21836 20588 21888
rect 23664 21836 23716 21888
rect 29184 21836 29236 21888
rect 33784 21981 33793 22015
rect 33793 21981 33827 22015
rect 33827 21981 33836 22015
rect 33784 21972 33836 21981
rect 31484 21904 31536 21956
rect 33600 21904 33652 21956
rect 36820 22049 36829 22083
rect 36829 22049 36863 22083
rect 36863 22049 36872 22083
rect 36820 22040 36872 22049
rect 37372 22040 37424 22092
rect 38108 22040 38160 22092
rect 34428 21972 34480 22024
rect 35440 22015 35492 22024
rect 35440 21981 35449 22015
rect 35449 21981 35483 22015
rect 35483 21981 35492 22015
rect 35440 21972 35492 21981
rect 38476 22015 38528 22024
rect 38476 21981 38485 22015
rect 38485 21981 38519 22015
rect 38519 21981 38528 22015
rect 38476 21972 38528 21981
rect 31760 21836 31812 21888
rect 4246 21734 4298 21786
rect 4310 21734 4362 21786
rect 4374 21734 4426 21786
rect 4438 21734 4490 21786
rect 34966 21734 35018 21786
rect 35030 21734 35082 21786
rect 35094 21734 35146 21786
rect 35158 21734 35210 21786
rect 3332 21632 3384 21684
rect 5540 21564 5592 21616
rect 6920 21607 6972 21616
rect 1768 21496 1820 21548
rect 3976 21496 4028 21548
rect 4896 21496 4948 21548
rect 6920 21573 6929 21607
rect 6929 21573 6963 21607
rect 6963 21573 6972 21607
rect 6920 21564 6972 21573
rect 1492 21428 1544 21480
rect 1952 21428 2004 21480
rect 4068 21471 4120 21480
rect 4068 21437 4077 21471
rect 4077 21437 4111 21471
rect 4111 21437 4120 21471
rect 4068 21428 4120 21437
rect 4988 21471 5040 21480
rect 2964 21360 3016 21412
rect 4988 21437 4997 21471
rect 4997 21437 5031 21471
rect 5031 21437 5040 21471
rect 4988 21428 5040 21437
rect 10784 21496 10836 21548
rect 6736 21428 6788 21480
rect 7472 21471 7524 21480
rect 7472 21437 7481 21471
rect 7481 21437 7515 21471
rect 7515 21437 7524 21471
rect 7472 21428 7524 21437
rect 10692 21471 10744 21480
rect 10692 21437 10701 21471
rect 10701 21437 10735 21471
rect 10735 21437 10744 21471
rect 10692 21428 10744 21437
rect 12532 21496 12584 21548
rect 12440 21428 12492 21480
rect 12716 21428 12768 21480
rect 16948 21632 17000 21684
rect 18144 21675 18196 21684
rect 18144 21641 18153 21675
rect 18153 21641 18187 21675
rect 18187 21641 18196 21675
rect 18144 21632 18196 21641
rect 20352 21564 20404 21616
rect 13728 21539 13780 21548
rect 13728 21505 13737 21539
rect 13737 21505 13771 21539
rect 13771 21505 13780 21539
rect 13728 21496 13780 21505
rect 13820 21496 13872 21548
rect 21456 21564 21508 21616
rect 22560 21564 22612 21616
rect 13176 21471 13228 21480
rect 13176 21437 13185 21471
rect 13185 21437 13219 21471
rect 13219 21437 13228 21471
rect 13176 21428 13228 21437
rect 14464 21471 14516 21480
rect 5540 21360 5592 21412
rect 11704 21360 11756 21412
rect 14464 21437 14473 21471
rect 14473 21437 14507 21471
rect 14507 21437 14516 21471
rect 14464 21428 14516 21437
rect 16580 21471 16632 21480
rect 16580 21437 16589 21471
rect 16589 21437 16623 21471
rect 16623 21437 16632 21471
rect 16580 21428 16632 21437
rect 13728 21360 13780 21412
rect 16120 21360 16172 21412
rect 16488 21360 16540 21412
rect 17132 21428 17184 21480
rect 19156 21471 19208 21480
rect 13084 21292 13136 21344
rect 19156 21437 19165 21471
rect 19165 21437 19199 21471
rect 19199 21437 19208 21471
rect 19156 21428 19208 21437
rect 20904 21360 20956 21412
rect 21456 21471 21508 21480
rect 21456 21437 21465 21471
rect 21465 21437 21499 21471
rect 21499 21437 21508 21471
rect 21456 21428 21508 21437
rect 21916 21360 21968 21412
rect 22560 21471 22612 21480
rect 22560 21437 22569 21471
rect 22569 21437 22603 21471
rect 22603 21437 22612 21471
rect 22560 21428 22612 21437
rect 22836 21428 22888 21480
rect 25688 21632 25740 21684
rect 25780 21632 25832 21684
rect 34152 21632 34204 21684
rect 26792 21564 26844 21616
rect 23480 21496 23532 21548
rect 23848 21496 23900 21548
rect 26148 21471 26200 21480
rect 26148 21437 26157 21471
rect 26157 21437 26191 21471
rect 26191 21437 26200 21471
rect 26148 21428 26200 21437
rect 29000 21496 29052 21548
rect 34336 21564 34388 21616
rect 32312 21539 32364 21548
rect 32312 21505 32321 21539
rect 32321 21505 32355 21539
rect 32355 21505 32364 21539
rect 32312 21496 32364 21505
rect 32956 21496 33008 21548
rect 26976 21471 27028 21480
rect 26424 21360 26476 21412
rect 26976 21437 26985 21471
rect 26985 21437 27019 21471
rect 27019 21437 27028 21471
rect 26976 21428 27028 21437
rect 27712 21471 27764 21480
rect 27712 21437 27721 21471
rect 27721 21437 27755 21471
rect 27755 21437 27764 21471
rect 27712 21428 27764 21437
rect 28172 21471 28224 21480
rect 28172 21437 28181 21471
rect 28181 21437 28215 21471
rect 28215 21437 28224 21471
rect 28172 21428 28224 21437
rect 29184 21428 29236 21480
rect 27988 21360 28040 21412
rect 31484 21428 31536 21480
rect 33232 21471 33284 21480
rect 33232 21437 33241 21471
rect 33241 21437 33275 21471
rect 33275 21437 33284 21471
rect 33232 21428 33284 21437
rect 33968 21496 34020 21548
rect 34152 21471 34204 21480
rect 34152 21437 34161 21471
rect 34161 21437 34195 21471
rect 34195 21437 34204 21471
rect 34152 21428 34204 21437
rect 36176 21632 36228 21684
rect 35624 21564 35676 21616
rect 35808 21564 35860 21616
rect 35440 21539 35492 21548
rect 35440 21505 35449 21539
rect 35449 21505 35483 21539
rect 35483 21505 35492 21539
rect 35440 21496 35492 21505
rect 36452 21496 36504 21548
rect 37832 21496 37884 21548
rect 35808 21471 35860 21480
rect 22560 21292 22612 21344
rect 23296 21335 23348 21344
rect 23296 21301 23305 21335
rect 23305 21301 23339 21335
rect 23339 21301 23348 21335
rect 23296 21292 23348 21301
rect 23388 21292 23440 21344
rect 25780 21292 25832 21344
rect 26240 21335 26292 21344
rect 26240 21301 26249 21335
rect 26249 21301 26283 21335
rect 26283 21301 26292 21335
rect 26240 21292 26292 21301
rect 27620 21292 27672 21344
rect 29368 21292 29420 21344
rect 30012 21292 30064 21344
rect 31852 21292 31904 21344
rect 33048 21335 33100 21344
rect 33048 21301 33057 21335
rect 33057 21301 33091 21335
rect 33091 21301 33100 21335
rect 33048 21292 33100 21301
rect 34060 21292 34112 21344
rect 35808 21437 35817 21471
rect 35817 21437 35851 21471
rect 35851 21437 35860 21471
rect 35808 21428 35860 21437
rect 35992 21428 36044 21480
rect 36268 21428 36320 21480
rect 36544 21428 36596 21480
rect 36912 21428 36964 21480
rect 39028 21360 39080 21412
rect 38660 21292 38712 21344
rect 19606 21190 19658 21242
rect 19670 21190 19722 21242
rect 19734 21190 19786 21242
rect 19798 21190 19850 21242
rect 1952 21131 2004 21140
rect 1952 21097 1961 21131
rect 1961 21097 1995 21131
rect 1995 21097 2004 21131
rect 1952 21088 2004 21097
rect 5540 21088 5592 21140
rect 5908 21088 5960 21140
rect 1768 21020 1820 21072
rect 2504 21020 2556 21072
rect 1860 20995 1912 21004
rect 1860 20961 1869 20995
rect 1869 20961 1903 20995
rect 1903 20961 1912 20995
rect 1860 20952 1912 20961
rect 2964 20995 3016 21004
rect 2964 20961 2973 20995
rect 2973 20961 3007 20995
rect 3007 20961 3016 20995
rect 2964 20952 3016 20961
rect 3332 20995 3384 21004
rect 3332 20961 3341 20995
rect 3341 20961 3375 20995
rect 3375 20961 3384 20995
rect 3332 20952 3384 20961
rect 5632 20952 5684 21004
rect 9864 21088 9916 21140
rect 15384 21131 15436 21140
rect 8852 21020 8904 21072
rect 1676 20884 1728 20936
rect 4988 20884 5040 20936
rect 3976 20816 4028 20868
rect 9956 20995 10008 21004
rect 5816 20927 5868 20936
rect 5816 20893 5825 20927
rect 5825 20893 5859 20927
rect 5859 20893 5868 20927
rect 5816 20884 5868 20893
rect 6920 20884 6972 20936
rect 9128 20884 9180 20936
rect 8668 20816 8720 20868
rect 9956 20961 9965 20995
rect 9965 20961 9999 20995
rect 9999 20961 10008 20995
rect 9956 20952 10008 20961
rect 10416 20995 10468 21004
rect 10416 20961 10425 20995
rect 10425 20961 10459 20995
rect 10459 20961 10468 20995
rect 10416 20952 10468 20961
rect 13176 21020 13228 21072
rect 15384 21097 15393 21131
rect 15393 21097 15427 21131
rect 15427 21097 15436 21131
rect 15384 21088 15436 21097
rect 17592 21088 17644 21140
rect 21640 21088 21692 21140
rect 24860 21088 24912 21140
rect 26516 21088 26568 21140
rect 28264 21088 28316 21140
rect 32220 21088 32272 21140
rect 34152 21088 34204 21140
rect 35440 21088 35492 21140
rect 35808 21088 35860 21140
rect 11152 20995 11204 21004
rect 11152 20961 11161 20995
rect 11161 20961 11195 20995
rect 11195 20961 11204 20995
rect 11152 20952 11204 20961
rect 11612 20995 11664 21004
rect 11612 20961 11621 20995
rect 11621 20961 11655 20995
rect 11655 20961 11664 20995
rect 11612 20952 11664 20961
rect 12716 20995 12768 21004
rect 12716 20961 12725 20995
rect 12725 20961 12759 20995
rect 12759 20961 12768 20995
rect 12716 20952 12768 20961
rect 14188 21020 14240 21072
rect 14280 21020 14332 21072
rect 13728 20995 13780 21004
rect 13728 20961 13737 20995
rect 13737 20961 13771 20995
rect 13771 20961 13780 20995
rect 13728 20952 13780 20961
rect 15292 20995 15344 21004
rect 13084 20884 13136 20936
rect 15292 20961 15301 20995
rect 15301 20961 15335 20995
rect 15335 20961 15344 20995
rect 15292 20952 15344 20961
rect 16672 20995 16724 21004
rect 16672 20961 16681 20995
rect 16681 20961 16715 20995
rect 16715 20961 16724 20995
rect 16672 20952 16724 20961
rect 16856 20995 16908 21004
rect 16856 20961 16865 20995
rect 16865 20961 16899 20995
rect 16899 20961 16908 20995
rect 16856 20952 16908 20961
rect 17132 20995 17184 21004
rect 17132 20961 17141 20995
rect 17141 20961 17175 20995
rect 17175 20961 17184 20995
rect 17132 20952 17184 20961
rect 17316 20995 17368 21004
rect 17316 20961 17325 20995
rect 17325 20961 17359 20995
rect 17359 20961 17368 20995
rect 17316 20952 17368 20961
rect 17592 20995 17644 21004
rect 17592 20961 17601 20995
rect 17601 20961 17635 20995
rect 17635 20961 17644 20995
rect 17592 20952 17644 20961
rect 19156 21020 19208 21072
rect 19432 21020 19484 21072
rect 19984 21063 20036 21072
rect 19984 21029 19993 21063
rect 19993 21029 20027 21063
rect 20027 21029 20036 21063
rect 19984 21020 20036 21029
rect 19892 20995 19944 21004
rect 10416 20816 10468 20868
rect 12164 20816 12216 20868
rect 18880 20884 18932 20936
rect 19892 20961 19901 20995
rect 19901 20961 19935 20995
rect 19935 20961 19944 20995
rect 19892 20952 19944 20961
rect 20168 20952 20220 21004
rect 22836 21020 22888 21072
rect 20904 20952 20956 21004
rect 21272 20952 21324 21004
rect 22560 20995 22612 21004
rect 22560 20961 22569 20995
rect 22569 20961 22603 20995
rect 22603 20961 22612 20995
rect 22560 20952 22612 20961
rect 23388 20952 23440 21004
rect 25688 21020 25740 21072
rect 23756 20995 23808 21004
rect 23756 20961 23765 20995
rect 23765 20961 23799 20995
rect 23799 20961 23808 20995
rect 23756 20952 23808 20961
rect 24124 20995 24176 21004
rect 24124 20961 24133 20995
rect 24133 20961 24167 20995
rect 24167 20961 24176 20995
rect 24124 20952 24176 20961
rect 24584 20952 24636 21004
rect 4620 20791 4672 20800
rect 4620 20757 4629 20791
rect 4629 20757 4663 20791
rect 4663 20757 4672 20791
rect 4620 20748 4672 20757
rect 5080 20791 5132 20800
rect 5080 20757 5089 20791
rect 5089 20757 5123 20791
rect 5123 20757 5132 20791
rect 5080 20748 5132 20757
rect 12992 20748 13044 20800
rect 13176 20748 13228 20800
rect 19064 20748 19116 20800
rect 21824 20884 21876 20936
rect 22376 20884 22428 20936
rect 22652 20884 22704 20936
rect 25596 20952 25648 21004
rect 28448 21020 28500 21072
rect 28908 21020 28960 21072
rect 26792 20995 26844 21004
rect 26792 20961 26801 20995
rect 26801 20961 26835 20995
rect 26835 20961 26844 20995
rect 26792 20952 26844 20961
rect 23112 20816 23164 20868
rect 25964 20884 26016 20936
rect 27068 20884 27120 20936
rect 26148 20816 26200 20868
rect 22100 20748 22152 20800
rect 22744 20791 22796 20800
rect 22744 20757 22753 20791
rect 22753 20757 22787 20791
rect 22787 20757 22796 20791
rect 22744 20748 22796 20757
rect 24768 20748 24820 20800
rect 27620 20952 27672 21004
rect 27712 20884 27764 20936
rect 30288 21020 30340 21072
rect 32956 21020 33008 21072
rect 34796 21063 34848 21072
rect 34796 21029 34805 21063
rect 34805 21029 34839 21063
rect 34839 21029 34848 21063
rect 34796 21020 34848 21029
rect 35256 21020 35308 21072
rect 29828 20927 29880 20936
rect 29828 20893 29837 20927
rect 29837 20893 29871 20927
rect 29871 20893 29880 20927
rect 29828 20884 29880 20893
rect 32312 20952 32364 21004
rect 32128 20884 32180 20936
rect 33692 20952 33744 21004
rect 37004 20952 37056 21004
rect 38660 20995 38712 21004
rect 33416 20927 33468 20936
rect 33416 20893 33425 20927
rect 33425 20893 33459 20927
rect 33459 20893 33468 20927
rect 33416 20884 33468 20893
rect 36452 20884 36504 20936
rect 37280 20884 37332 20936
rect 27896 20816 27948 20868
rect 29552 20816 29604 20868
rect 33140 20816 33192 20868
rect 36544 20816 36596 20868
rect 38660 20961 38669 20995
rect 38669 20961 38703 20995
rect 38703 20961 38712 20995
rect 38660 20952 38712 20961
rect 31208 20748 31260 20800
rect 34244 20748 34296 20800
rect 36636 20748 36688 20800
rect 36820 20748 36872 20800
rect 4246 20646 4298 20698
rect 4310 20646 4362 20698
rect 4374 20646 4426 20698
rect 4438 20646 4490 20698
rect 34966 20646 35018 20698
rect 35030 20646 35082 20698
rect 35094 20646 35146 20698
rect 35158 20646 35210 20698
rect 2964 20587 3016 20596
rect 2964 20553 2973 20587
rect 2973 20553 3007 20587
rect 3007 20553 3016 20587
rect 2964 20544 3016 20553
rect 4620 20544 4672 20596
rect 9956 20544 10008 20596
rect 12716 20544 12768 20596
rect 16304 20587 16356 20596
rect 16304 20553 16313 20587
rect 16313 20553 16347 20587
rect 16347 20553 16356 20587
rect 16304 20544 16356 20553
rect 18604 20544 18656 20596
rect 30288 20544 30340 20596
rect 10416 20476 10468 20528
rect 5080 20408 5132 20460
rect 6828 20408 6880 20460
rect 10232 20408 10284 20460
rect 10692 20451 10744 20460
rect 10692 20417 10701 20451
rect 10701 20417 10735 20451
rect 10735 20417 10744 20451
rect 10692 20408 10744 20417
rect 15108 20476 15160 20528
rect 23756 20519 23808 20528
rect 23756 20485 23765 20519
rect 23765 20485 23799 20519
rect 23799 20485 23808 20519
rect 23756 20476 23808 20485
rect 12440 20451 12492 20460
rect 12440 20417 12449 20451
rect 12449 20417 12483 20451
rect 12483 20417 12492 20451
rect 12440 20408 12492 20417
rect 1400 20383 1452 20392
rect 1400 20349 1409 20383
rect 1409 20349 1443 20383
rect 1443 20349 1452 20383
rect 1400 20340 1452 20349
rect 2044 20340 2096 20392
rect 4068 20340 4120 20392
rect 4160 20272 4212 20324
rect 5816 20340 5868 20392
rect 8208 20383 8260 20392
rect 8208 20349 8217 20383
rect 8217 20349 8251 20383
rect 8251 20349 8260 20383
rect 8208 20340 8260 20349
rect 10876 20383 10928 20392
rect 9128 20204 9180 20256
rect 10140 20204 10192 20256
rect 10876 20349 10885 20383
rect 10885 20349 10919 20383
rect 10919 20349 10928 20383
rect 10876 20340 10928 20349
rect 11704 20383 11756 20392
rect 11704 20349 11713 20383
rect 11713 20349 11747 20383
rect 11747 20349 11756 20383
rect 11704 20340 11756 20349
rect 13176 20408 13228 20460
rect 13452 20408 13504 20460
rect 19064 20408 19116 20460
rect 19432 20408 19484 20460
rect 26240 20408 26292 20460
rect 26792 20408 26844 20460
rect 13268 20383 13320 20392
rect 11152 20272 11204 20324
rect 11612 20272 11664 20324
rect 13268 20349 13277 20383
rect 13277 20349 13311 20383
rect 13311 20349 13320 20383
rect 13268 20340 13320 20349
rect 13728 20340 13780 20392
rect 13820 20340 13872 20392
rect 15016 20340 15068 20392
rect 16120 20383 16172 20392
rect 16120 20349 16129 20383
rect 16129 20349 16163 20383
rect 16163 20349 16172 20383
rect 16120 20340 16172 20349
rect 17500 20340 17552 20392
rect 22928 20340 22980 20392
rect 18512 20272 18564 20324
rect 18788 20272 18840 20324
rect 19432 20315 19484 20324
rect 19432 20281 19441 20315
rect 19441 20281 19475 20315
rect 19475 20281 19484 20315
rect 19432 20272 19484 20281
rect 21640 20315 21692 20324
rect 21640 20281 21649 20315
rect 21649 20281 21683 20315
rect 21683 20281 21692 20315
rect 21640 20272 21692 20281
rect 24216 20340 24268 20392
rect 24860 20383 24912 20392
rect 24860 20349 24869 20383
rect 24869 20349 24903 20383
rect 24903 20349 24912 20383
rect 24860 20340 24912 20349
rect 25688 20340 25740 20392
rect 26424 20383 26476 20392
rect 26424 20349 26433 20383
rect 26433 20349 26467 20383
rect 26467 20349 26476 20383
rect 26424 20340 26476 20349
rect 30104 20408 30156 20460
rect 38108 20544 38160 20596
rect 31392 20519 31444 20528
rect 31392 20485 31401 20519
rect 31401 20485 31435 20519
rect 31435 20485 31444 20519
rect 31392 20476 31444 20485
rect 32128 20451 32180 20460
rect 32128 20417 32137 20451
rect 32137 20417 32171 20451
rect 32171 20417 32180 20451
rect 32128 20408 32180 20417
rect 29184 20340 29236 20392
rect 29552 20383 29604 20392
rect 29552 20349 29561 20383
rect 29561 20349 29595 20383
rect 29595 20349 29604 20383
rect 29552 20340 29604 20349
rect 30472 20383 30524 20392
rect 30472 20349 30481 20383
rect 30481 20349 30515 20383
rect 30515 20349 30524 20383
rect 30472 20340 30524 20349
rect 30564 20340 30616 20392
rect 31024 20383 31076 20392
rect 31024 20349 31033 20383
rect 31033 20349 31067 20383
rect 31067 20349 31076 20383
rect 31024 20340 31076 20349
rect 31484 20340 31536 20392
rect 33140 20408 33192 20460
rect 34244 20408 34296 20460
rect 36452 20451 36504 20460
rect 36452 20417 36461 20451
rect 36461 20417 36495 20451
rect 36495 20417 36504 20451
rect 36452 20408 36504 20417
rect 32864 20340 32916 20392
rect 11796 20247 11848 20256
rect 11796 20213 11805 20247
rect 11805 20213 11839 20247
rect 11839 20213 11848 20247
rect 11796 20204 11848 20213
rect 15292 20247 15344 20256
rect 15292 20213 15301 20247
rect 15301 20213 15335 20247
rect 15335 20213 15344 20247
rect 15292 20204 15344 20213
rect 18696 20204 18748 20256
rect 22836 20204 22888 20256
rect 24492 20272 24544 20324
rect 24400 20204 24452 20256
rect 29276 20272 29328 20324
rect 32312 20272 32364 20324
rect 33508 20340 33560 20392
rect 34796 20340 34848 20392
rect 35256 20340 35308 20392
rect 36176 20340 36228 20392
rect 37740 20340 37792 20392
rect 38292 20340 38344 20392
rect 27712 20204 27764 20256
rect 29184 20204 29236 20256
rect 30012 20204 30064 20256
rect 34704 20204 34756 20256
rect 37004 20204 37056 20256
rect 38752 20204 38804 20256
rect 19606 20102 19658 20154
rect 19670 20102 19722 20154
rect 19734 20102 19786 20154
rect 19798 20102 19850 20154
rect 10140 20043 10192 20052
rect 10140 20009 10149 20043
rect 10149 20009 10183 20043
rect 10183 20009 10192 20043
rect 10140 20000 10192 20009
rect 11428 20000 11480 20052
rect 2964 19932 3016 19984
rect 8208 19932 8260 19984
rect 9128 19932 9180 19984
rect 13084 19932 13136 19984
rect 17224 20000 17276 20052
rect 17776 20000 17828 20052
rect 17316 19932 17368 19984
rect 19984 20000 20036 20052
rect 3332 19907 3384 19916
rect 3332 19873 3341 19907
rect 3341 19873 3375 19907
rect 3375 19873 3384 19907
rect 4068 19907 4120 19916
rect 3332 19864 3384 19873
rect 3516 19839 3568 19848
rect 3516 19805 3525 19839
rect 3525 19805 3559 19839
rect 3559 19805 3568 19839
rect 3516 19796 3568 19805
rect 4068 19873 4077 19907
rect 4077 19873 4111 19907
rect 4111 19873 4120 19907
rect 4068 19864 4120 19873
rect 4804 19907 4856 19916
rect 4804 19873 4813 19907
rect 4813 19873 4847 19907
rect 4847 19873 4856 19907
rect 4804 19864 4856 19873
rect 4988 19907 5040 19916
rect 4988 19873 4997 19907
rect 4997 19873 5031 19907
rect 5031 19873 5040 19907
rect 4988 19864 5040 19873
rect 5816 19864 5868 19916
rect 6828 19864 6880 19916
rect 8668 19907 8720 19916
rect 8668 19873 8677 19907
rect 8677 19873 8711 19907
rect 8711 19873 8720 19907
rect 8668 19864 8720 19873
rect 9956 19907 10008 19916
rect 9956 19873 9965 19907
rect 9965 19873 9999 19907
rect 9999 19873 10008 19907
rect 9956 19864 10008 19873
rect 10692 19907 10744 19916
rect 10692 19873 10701 19907
rect 10701 19873 10735 19907
rect 10735 19873 10744 19907
rect 10692 19864 10744 19873
rect 11796 19907 11848 19916
rect 11796 19873 11805 19907
rect 11805 19873 11839 19907
rect 11839 19873 11848 19907
rect 11796 19864 11848 19873
rect 14188 19907 14240 19916
rect 14188 19873 14197 19907
rect 14197 19873 14231 19907
rect 14231 19873 14240 19907
rect 14188 19864 14240 19873
rect 15200 19864 15252 19916
rect 16212 19864 16264 19916
rect 16856 19907 16908 19916
rect 3976 19796 4028 19848
rect 6000 19839 6052 19848
rect 6000 19805 6009 19839
rect 6009 19805 6043 19839
rect 6043 19805 6052 19839
rect 6000 19796 6052 19805
rect 10876 19796 10928 19848
rect 4712 19728 4764 19780
rect 10232 19728 10284 19780
rect 12440 19796 12492 19848
rect 14740 19796 14792 19848
rect 16856 19873 16865 19907
rect 16865 19873 16899 19907
rect 16899 19873 16908 19907
rect 16856 19864 16908 19873
rect 16948 19907 17000 19916
rect 16948 19873 16957 19907
rect 16957 19873 16991 19907
rect 16991 19873 17000 19907
rect 17132 19907 17184 19916
rect 16948 19864 17000 19873
rect 17132 19873 17141 19907
rect 17141 19873 17175 19907
rect 17175 19873 17184 19907
rect 17132 19864 17184 19873
rect 17500 19907 17552 19916
rect 17500 19873 17509 19907
rect 17509 19873 17543 19907
rect 17543 19873 17552 19907
rect 17500 19864 17552 19873
rect 17684 19907 17736 19916
rect 7104 19703 7156 19712
rect 7104 19669 7113 19703
rect 7113 19669 7147 19703
rect 7147 19669 7156 19703
rect 7104 19660 7156 19669
rect 14832 19728 14884 19780
rect 16672 19796 16724 19848
rect 17684 19873 17693 19907
rect 17693 19873 17727 19907
rect 17727 19873 17736 19907
rect 17684 19864 17736 19873
rect 18604 19907 18656 19916
rect 18604 19873 18613 19907
rect 18613 19873 18647 19907
rect 18647 19873 18656 19907
rect 18604 19864 18656 19873
rect 19708 19932 19760 19984
rect 18144 19796 18196 19848
rect 18512 19796 18564 19848
rect 18788 19796 18840 19848
rect 20352 19864 20404 19916
rect 19800 19796 19852 19848
rect 20812 19796 20864 19848
rect 21916 19839 21968 19848
rect 21916 19805 21925 19839
rect 21925 19805 21959 19839
rect 21959 19805 21968 19839
rect 21916 19796 21968 19805
rect 22284 19796 22336 19848
rect 17500 19728 17552 19780
rect 20352 19728 20404 19780
rect 24768 20000 24820 20052
rect 25964 20000 26016 20052
rect 22836 19932 22888 19984
rect 29368 20000 29420 20052
rect 23020 19907 23072 19916
rect 23020 19873 23029 19907
rect 23029 19873 23063 19907
rect 23063 19873 23072 19907
rect 23020 19864 23072 19873
rect 22836 19796 22888 19848
rect 24584 19907 24636 19916
rect 24584 19873 24593 19907
rect 24593 19873 24627 19907
rect 24627 19873 24636 19907
rect 24584 19864 24636 19873
rect 25504 19864 25556 19916
rect 27712 19932 27764 19984
rect 27620 19907 27672 19916
rect 27620 19873 27629 19907
rect 27629 19873 27663 19907
rect 27663 19873 27672 19907
rect 27620 19864 27672 19873
rect 27896 19907 27948 19916
rect 27896 19873 27905 19907
rect 27905 19873 27939 19907
rect 27939 19873 27948 19907
rect 27896 19864 27948 19873
rect 31668 20000 31720 20052
rect 30104 19932 30156 19984
rect 29736 19864 29788 19916
rect 30656 19907 30708 19916
rect 30656 19873 30665 19907
rect 30665 19873 30699 19907
rect 30699 19873 30708 19907
rect 30656 19864 30708 19873
rect 30748 19864 30800 19916
rect 32220 19907 32272 19916
rect 32220 19873 32229 19907
rect 32229 19873 32263 19907
rect 32263 19873 32272 19907
rect 32220 19864 32272 19873
rect 34336 20000 34388 20052
rect 36912 20000 36964 20052
rect 36544 19932 36596 19984
rect 34428 19907 34480 19916
rect 27988 19839 28040 19848
rect 24032 19771 24084 19780
rect 24032 19737 24041 19771
rect 24041 19737 24075 19771
rect 24075 19737 24084 19771
rect 24032 19728 24084 19737
rect 24124 19728 24176 19780
rect 27988 19805 27997 19839
rect 27997 19805 28031 19839
rect 28031 19805 28040 19839
rect 27988 19796 28040 19805
rect 30472 19796 30524 19848
rect 32128 19839 32180 19848
rect 32128 19805 32137 19839
rect 32137 19805 32171 19839
rect 32171 19805 32180 19839
rect 32128 19796 32180 19805
rect 33416 19839 33468 19848
rect 33416 19805 33425 19839
rect 33425 19805 33459 19839
rect 33459 19805 33468 19839
rect 33416 19796 33468 19805
rect 32036 19728 32088 19780
rect 34428 19873 34437 19907
rect 34437 19873 34471 19907
rect 34471 19873 34480 19907
rect 34428 19864 34480 19873
rect 35808 19864 35860 19916
rect 36820 19932 36872 19984
rect 37740 19975 37792 19984
rect 35900 19796 35952 19848
rect 36728 19796 36780 19848
rect 36268 19728 36320 19780
rect 37004 19864 37056 19916
rect 37740 19941 37749 19975
rect 37749 19941 37783 19975
rect 37783 19941 37792 19975
rect 37740 19932 37792 19941
rect 37188 19864 37240 19916
rect 38752 19907 38804 19916
rect 38752 19873 38761 19907
rect 38761 19873 38795 19907
rect 38795 19873 38804 19907
rect 38752 19864 38804 19873
rect 38292 19796 38344 19848
rect 38936 19728 38988 19780
rect 14096 19660 14148 19712
rect 19340 19660 19392 19712
rect 19708 19660 19760 19712
rect 20168 19660 20220 19712
rect 20812 19660 20864 19712
rect 22192 19660 22244 19712
rect 29000 19660 29052 19712
rect 29736 19660 29788 19712
rect 4246 19558 4298 19610
rect 4310 19558 4362 19610
rect 4374 19558 4426 19610
rect 4438 19558 4490 19610
rect 34966 19558 35018 19610
rect 35030 19558 35082 19610
rect 35094 19558 35146 19610
rect 35158 19558 35210 19610
rect 2044 19499 2096 19508
rect 2044 19465 2053 19499
rect 2053 19465 2087 19499
rect 2087 19465 2096 19499
rect 2044 19456 2096 19465
rect 4620 19456 4672 19508
rect 4988 19456 5040 19508
rect 10692 19456 10744 19508
rect 1676 19295 1728 19304
rect 1676 19261 1685 19295
rect 1685 19261 1719 19295
rect 1719 19261 1728 19295
rect 1676 19252 1728 19261
rect 1768 19295 1820 19304
rect 1768 19261 1777 19295
rect 1777 19261 1811 19295
rect 1811 19261 1820 19295
rect 1768 19252 1820 19261
rect 3516 19320 3568 19372
rect 3056 19295 3108 19304
rect 1400 19116 1452 19168
rect 3056 19261 3065 19295
rect 3065 19261 3099 19295
rect 3099 19261 3108 19295
rect 3056 19252 3108 19261
rect 3884 19252 3936 19304
rect 5908 19295 5960 19304
rect 5908 19261 5917 19295
rect 5917 19261 5951 19295
rect 5951 19261 5960 19295
rect 5908 19252 5960 19261
rect 7196 19252 7248 19304
rect 4804 19184 4856 19236
rect 8576 19252 8628 19304
rect 9036 19252 9088 19304
rect 11244 19252 11296 19304
rect 12440 19388 12492 19440
rect 14188 19456 14240 19508
rect 15200 19388 15252 19440
rect 12992 19252 13044 19304
rect 14740 19320 14792 19372
rect 14924 19320 14976 19372
rect 13820 19252 13872 19304
rect 15016 19295 15068 19304
rect 15016 19261 15025 19295
rect 15025 19261 15059 19295
rect 15059 19261 15068 19295
rect 15016 19252 15068 19261
rect 15292 19252 15344 19304
rect 6920 19159 6972 19168
rect 6920 19125 6929 19159
rect 6929 19125 6963 19159
rect 6963 19125 6972 19159
rect 6920 19116 6972 19125
rect 9864 19116 9916 19168
rect 13544 19184 13596 19236
rect 15936 19252 15988 19304
rect 16212 19252 16264 19304
rect 17040 19456 17092 19508
rect 18512 19456 18564 19508
rect 19156 19456 19208 19508
rect 20720 19456 20772 19508
rect 29552 19456 29604 19508
rect 32220 19456 32272 19508
rect 34244 19499 34296 19508
rect 34244 19465 34253 19499
rect 34253 19465 34287 19499
rect 34287 19465 34296 19499
rect 34244 19456 34296 19465
rect 16948 19388 17000 19440
rect 19616 19388 19668 19440
rect 20444 19388 20496 19440
rect 21088 19388 21140 19440
rect 21732 19388 21784 19440
rect 22192 19388 22244 19440
rect 32496 19388 32548 19440
rect 35256 19456 35308 19508
rect 19340 19320 19392 19372
rect 17224 19252 17276 19304
rect 17500 19252 17552 19304
rect 17684 19252 17736 19304
rect 18788 19252 18840 19304
rect 23388 19320 23440 19372
rect 25872 19363 25924 19372
rect 25872 19329 25881 19363
rect 25881 19329 25915 19363
rect 25915 19329 25924 19363
rect 25872 19320 25924 19329
rect 19616 19295 19668 19304
rect 19616 19261 19625 19295
rect 19625 19261 19659 19295
rect 19659 19261 19668 19295
rect 19616 19252 19668 19261
rect 19708 19295 19760 19304
rect 19708 19261 19717 19295
rect 19717 19261 19751 19295
rect 19751 19261 19760 19295
rect 19708 19252 19760 19261
rect 19984 19295 20036 19304
rect 19984 19261 19993 19295
rect 19993 19261 20027 19295
rect 20027 19261 20036 19295
rect 19984 19252 20036 19261
rect 20352 19252 20404 19304
rect 20904 19252 20956 19304
rect 21272 19252 21324 19304
rect 21824 19295 21876 19304
rect 21824 19261 21833 19295
rect 21833 19261 21867 19295
rect 21867 19261 21876 19295
rect 21824 19252 21876 19261
rect 22100 19252 22152 19304
rect 22836 19295 22888 19304
rect 11704 19159 11756 19168
rect 11704 19125 11713 19159
rect 11713 19125 11747 19159
rect 11747 19125 11756 19159
rect 11704 19116 11756 19125
rect 14556 19116 14608 19168
rect 15844 19116 15896 19168
rect 16856 19116 16908 19168
rect 16948 19116 17000 19168
rect 22836 19261 22845 19295
rect 22845 19261 22879 19295
rect 22879 19261 22888 19295
rect 22836 19252 22888 19261
rect 22928 19295 22980 19304
rect 22928 19261 22937 19295
rect 22937 19261 22971 19295
rect 22971 19261 22980 19295
rect 23664 19295 23716 19304
rect 22928 19252 22980 19261
rect 23664 19261 23673 19295
rect 23673 19261 23707 19295
rect 23707 19261 23716 19295
rect 23664 19252 23716 19261
rect 24032 19252 24084 19304
rect 24676 19295 24728 19304
rect 24676 19261 24685 19295
rect 24685 19261 24719 19295
rect 24719 19261 24728 19295
rect 24676 19252 24728 19261
rect 24124 19184 24176 19236
rect 23480 19116 23532 19168
rect 23572 19116 23624 19168
rect 26608 19295 26660 19304
rect 26608 19261 26617 19295
rect 26617 19261 26651 19295
rect 26651 19261 26660 19295
rect 26608 19252 26660 19261
rect 27712 19252 27764 19304
rect 27160 19184 27212 19236
rect 26792 19116 26844 19168
rect 27068 19116 27120 19168
rect 28448 19295 28500 19304
rect 28448 19261 28457 19295
rect 28457 19261 28491 19295
rect 28491 19261 28500 19295
rect 28448 19252 28500 19261
rect 29736 19320 29788 19372
rect 30748 19320 30800 19372
rect 29092 19252 29144 19304
rect 29644 19295 29696 19304
rect 29368 19184 29420 19236
rect 29644 19261 29653 19295
rect 29653 19261 29687 19295
rect 29687 19261 29696 19295
rect 29644 19252 29696 19261
rect 30104 19295 30156 19304
rect 30104 19261 30113 19295
rect 30113 19261 30147 19295
rect 30147 19261 30156 19295
rect 30104 19252 30156 19261
rect 31392 19295 31444 19304
rect 31392 19261 31401 19295
rect 31401 19261 31435 19295
rect 31435 19261 31444 19295
rect 31392 19252 31444 19261
rect 30656 19184 30708 19236
rect 31300 19184 31352 19236
rect 31668 19252 31720 19304
rect 32864 19320 32916 19372
rect 32220 19295 32272 19304
rect 32220 19261 32229 19295
rect 32229 19261 32263 19295
rect 32263 19261 32272 19295
rect 32220 19252 32272 19261
rect 33140 19295 33192 19304
rect 33140 19261 33149 19295
rect 33149 19261 33183 19295
rect 33183 19261 33192 19295
rect 33140 19252 33192 19261
rect 33324 19295 33376 19304
rect 33324 19261 33333 19295
rect 33333 19261 33367 19295
rect 33367 19261 33376 19295
rect 33324 19252 33376 19261
rect 33968 19252 34020 19304
rect 34796 19320 34848 19372
rect 34152 19295 34204 19304
rect 34152 19261 34161 19295
rect 34161 19261 34195 19295
rect 34195 19261 34204 19295
rect 36452 19320 36504 19372
rect 34152 19252 34204 19261
rect 36360 19295 36412 19304
rect 36360 19261 36369 19295
rect 36369 19261 36403 19295
rect 36403 19261 36412 19295
rect 36360 19252 36412 19261
rect 36728 19295 36780 19304
rect 36728 19261 36737 19295
rect 36737 19261 36771 19295
rect 36771 19261 36780 19295
rect 36728 19252 36780 19261
rect 36912 19252 36964 19304
rect 30380 19116 30432 19168
rect 32128 19116 32180 19168
rect 34520 19116 34572 19168
rect 36544 19116 36596 19168
rect 36728 19116 36780 19168
rect 19606 19014 19658 19066
rect 19670 19014 19722 19066
rect 19734 19014 19786 19066
rect 19798 19014 19850 19066
rect 2780 18955 2832 18964
rect 2780 18921 2789 18955
rect 2789 18921 2823 18955
rect 2823 18921 2832 18955
rect 4160 18955 4212 18964
rect 2780 18912 2832 18921
rect 4160 18921 4169 18955
rect 4169 18921 4203 18955
rect 4203 18921 4212 18955
rect 4160 18912 4212 18921
rect 6000 18912 6052 18964
rect 9036 18955 9088 18964
rect 9036 18921 9045 18955
rect 9045 18921 9079 18955
rect 9079 18921 9088 18955
rect 9036 18912 9088 18921
rect 14372 18912 14424 18964
rect 1400 18819 1452 18828
rect 1400 18785 1409 18819
rect 1409 18785 1443 18819
rect 1443 18785 1452 18819
rect 1400 18776 1452 18785
rect 3516 18776 3568 18828
rect 5172 18819 5224 18828
rect 5172 18785 5181 18819
rect 5181 18785 5215 18819
rect 5215 18785 5224 18819
rect 5172 18776 5224 18785
rect 6276 18819 6328 18828
rect 6276 18785 6285 18819
rect 6285 18785 6319 18819
rect 6319 18785 6328 18819
rect 6276 18776 6328 18785
rect 6828 18819 6880 18828
rect 6828 18785 6837 18819
rect 6837 18785 6871 18819
rect 6871 18785 6880 18819
rect 6828 18776 6880 18785
rect 7104 18819 7156 18828
rect 7104 18785 7113 18819
rect 7113 18785 7147 18819
rect 7147 18785 7156 18819
rect 7104 18776 7156 18785
rect 5080 18751 5132 18760
rect 5080 18717 5089 18751
rect 5089 18717 5123 18751
rect 5123 18717 5132 18751
rect 5080 18708 5132 18717
rect 7932 18572 7984 18624
rect 15384 18844 15436 18896
rect 14556 18819 14608 18828
rect 14556 18785 14565 18819
rect 14565 18785 14599 18819
rect 14599 18785 14608 18819
rect 14556 18776 14608 18785
rect 15844 18776 15896 18828
rect 16948 18776 17000 18828
rect 10232 18708 10284 18760
rect 10600 18751 10652 18760
rect 10600 18717 10609 18751
rect 10609 18717 10643 18751
rect 10643 18717 10652 18751
rect 10600 18708 10652 18717
rect 12440 18751 12492 18760
rect 12440 18717 12449 18751
rect 12449 18717 12483 18751
rect 12483 18717 12492 18751
rect 12440 18708 12492 18717
rect 13544 18708 13596 18760
rect 16764 18708 16816 18760
rect 19064 18912 19116 18964
rect 20076 18912 20128 18964
rect 21180 18912 21232 18964
rect 21456 18912 21508 18964
rect 17316 18776 17368 18828
rect 18420 18819 18472 18828
rect 18420 18785 18429 18819
rect 18429 18785 18463 18819
rect 18463 18785 18472 18819
rect 18420 18776 18472 18785
rect 18788 18776 18840 18828
rect 19524 18844 19576 18896
rect 19616 18887 19668 18896
rect 19616 18853 19625 18887
rect 19625 18853 19659 18887
rect 19659 18853 19668 18887
rect 19616 18844 19668 18853
rect 20168 18844 20220 18896
rect 21364 18844 21416 18896
rect 22008 18844 22060 18896
rect 22836 18844 22888 18896
rect 25136 18844 25188 18896
rect 21272 18776 21324 18828
rect 21916 18819 21968 18828
rect 21916 18785 21925 18819
rect 21925 18785 21959 18819
rect 21959 18785 21968 18819
rect 21916 18776 21968 18785
rect 22468 18819 22520 18828
rect 22468 18785 22477 18819
rect 22477 18785 22511 18819
rect 22511 18785 22520 18819
rect 22468 18776 22520 18785
rect 24032 18819 24084 18828
rect 21824 18708 21876 18760
rect 24032 18785 24041 18819
rect 24041 18785 24075 18819
rect 24075 18785 24084 18819
rect 24032 18776 24084 18785
rect 25504 18776 25556 18828
rect 25688 18819 25740 18828
rect 25688 18785 25697 18819
rect 25697 18785 25731 18819
rect 25731 18785 25740 18819
rect 25688 18776 25740 18785
rect 26792 18819 26844 18828
rect 26792 18785 26801 18819
rect 26801 18785 26835 18819
rect 26835 18785 26844 18819
rect 26792 18776 26844 18785
rect 11980 18640 12032 18692
rect 11888 18615 11940 18624
rect 11888 18581 11897 18615
rect 11897 18581 11931 18615
rect 11931 18581 11940 18615
rect 11888 18572 11940 18581
rect 12624 18572 12676 18624
rect 17500 18640 17552 18692
rect 18972 18640 19024 18692
rect 13728 18572 13780 18624
rect 14372 18572 14424 18624
rect 20352 18572 20404 18624
rect 20536 18572 20588 18624
rect 21180 18572 21232 18624
rect 22376 18572 22428 18624
rect 23848 18640 23900 18692
rect 24676 18708 24728 18760
rect 26240 18708 26292 18760
rect 26976 18776 27028 18828
rect 27160 18819 27212 18828
rect 27160 18785 27169 18819
rect 27169 18785 27203 18819
rect 27203 18785 27212 18819
rect 27160 18776 27212 18785
rect 27436 18819 27488 18828
rect 27436 18785 27445 18819
rect 27445 18785 27479 18819
rect 27479 18785 27488 18819
rect 27436 18776 27488 18785
rect 27712 18819 27764 18828
rect 27712 18785 27721 18819
rect 27721 18785 27755 18819
rect 27755 18785 27764 18819
rect 27712 18776 27764 18785
rect 29368 18819 29420 18828
rect 29092 18751 29144 18760
rect 29092 18717 29101 18751
rect 29101 18717 29135 18751
rect 29135 18717 29144 18751
rect 29092 18708 29144 18717
rect 29368 18785 29377 18819
rect 29377 18785 29411 18819
rect 29411 18785 29420 18819
rect 29368 18776 29420 18785
rect 30656 18912 30708 18964
rect 30748 18887 30800 18896
rect 30748 18853 30757 18887
rect 30757 18853 30791 18887
rect 30791 18853 30800 18887
rect 30748 18844 30800 18853
rect 31576 18844 31628 18896
rect 31300 18776 31352 18828
rect 35716 18912 35768 18964
rect 37372 18912 37424 18964
rect 37740 18912 37792 18964
rect 32864 18887 32916 18896
rect 32864 18853 32873 18887
rect 32873 18853 32907 18887
rect 32907 18853 32916 18887
rect 32864 18844 32916 18853
rect 32956 18844 33008 18896
rect 32588 18819 32640 18828
rect 32588 18785 32597 18819
rect 32597 18785 32631 18819
rect 32631 18785 32640 18819
rect 32588 18776 32640 18785
rect 33048 18776 33100 18828
rect 27068 18640 27120 18692
rect 28264 18640 28316 18692
rect 33508 18708 33560 18760
rect 33784 18844 33836 18896
rect 33968 18819 34020 18828
rect 33968 18785 33977 18819
rect 33977 18785 34011 18819
rect 34011 18785 34020 18819
rect 33968 18776 34020 18785
rect 34520 18776 34572 18828
rect 35256 18819 35308 18828
rect 35256 18785 35265 18819
rect 35265 18785 35299 18819
rect 35299 18785 35308 18819
rect 35256 18776 35308 18785
rect 35440 18819 35492 18828
rect 35440 18785 35449 18819
rect 35449 18785 35483 18819
rect 35483 18785 35492 18819
rect 35440 18776 35492 18785
rect 36544 18776 36596 18828
rect 36636 18776 36688 18828
rect 38292 18819 38344 18828
rect 38292 18785 38301 18819
rect 38301 18785 38335 18819
rect 38335 18785 38344 18819
rect 38292 18776 38344 18785
rect 38936 18819 38988 18828
rect 38936 18785 38945 18819
rect 38945 18785 38979 18819
rect 38979 18785 38988 18819
rect 38936 18776 38988 18785
rect 32496 18640 32548 18692
rect 37188 18640 37240 18692
rect 27712 18572 27764 18624
rect 28908 18572 28960 18624
rect 31208 18572 31260 18624
rect 36544 18572 36596 18624
rect 36636 18572 36688 18624
rect 4246 18470 4298 18522
rect 4310 18470 4362 18522
rect 4374 18470 4426 18522
rect 4438 18470 4490 18522
rect 34966 18470 35018 18522
rect 35030 18470 35082 18522
rect 35094 18470 35146 18522
rect 35158 18470 35210 18522
rect 5172 18368 5224 18420
rect 3056 18232 3108 18284
rect 4712 18232 4764 18284
rect 3976 18207 4028 18216
rect 3976 18173 3985 18207
rect 3985 18173 4019 18207
rect 4019 18173 4028 18207
rect 3976 18164 4028 18173
rect 5448 18164 5500 18216
rect 8392 18232 8444 18284
rect 10232 18368 10284 18420
rect 11244 18411 11296 18420
rect 11244 18377 11253 18411
rect 11253 18377 11287 18411
rect 11287 18377 11296 18411
rect 11244 18368 11296 18377
rect 15384 18368 15436 18420
rect 16212 18343 16264 18352
rect 16212 18309 16221 18343
rect 16221 18309 16255 18343
rect 16255 18309 16264 18343
rect 16212 18300 16264 18309
rect 19156 18300 19208 18352
rect 21456 18300 21508 18352
rect 26792 18368 26844 18420
rect 27436 18368 27488 18420
rect 28540 18368 28592 18420
rect 22836 18300 22888 18352
rect 25688 18300 25740 18352
rect 30288 18368 30340 18420
rect 32312 18343 32364 18352
rect 11888 18232 11940 18284
rect 8024 18207 8076 18216
rect 4620 18096 4672 18148
rect 6092 18096 6144 18148
rect 8024 18173 8033 18207
rect 8033 18173 8067 18207
rect 8067 18173 8076 18207
rect 8024 18164 8076 18173
rect 10232 18164 10284 18216
rect 11704 18164 11756 18216
rect 6828 18028 6880 18080
rect 7380 18028 7432 18080
rect 9404 18096 9456 18148
rect 13820 18207 13872 18216
rect 13820 18173 13829 18207
rect 13829 18173 13863 18207
rect 13863 18173 13872 18207
rect 13820 18164 13872 18173
rect 16120 18232 16172 18284
rect 17316 18232 17368 18284
rect 19616 18275 19668 18284
rect 16948 18207 17000 18216
rect 16948 18173 16957 18207
rect 16957 18173 16991 18207
rect 16991 18173 17000 18207
rect 16948 18164 17000 18173
rect 17040 18207 17092 18216
rect 17040 18173 17049 18207
rect 17049 18173 17083 18207
rect 17083 18173 17092 18207
rect 17040 18164 17092 18173
rect 19616 18241 19625 18275
rect 19625 18241 19659 18275
rect 19659 18241 19668 18275
rect 19616 18232 19668 18241
rect 19708 18232 19760 18284
rect 21916 18232 21968 18284
rect 18420 18164 18472 18216
rect 19156 18164 19208 18216
rect 17684 18096 17736 18148
rect 17776 18096 17828 18148
rect 20536 18164 20588 18216
rect 21364 18164 21416 18216
rect 21824 18164 21876 18216
rect 25872 18232 25924 18284
rect 28356 18232 28408 18284
rect 15200 18071 15252 18080
rect 15200 18037 15209 18071
rect 15209 18037 15243 18071
rect 15243 18037 15252 18071
rect 15200 18028 15252 18037
rect 15936 18028 15988 18080
rect 20352 18028 20404 18080
rect 21180 18028 21232 18080
rect 24768 18164 24820 18216
rect 24952 18164 25004 18216
rect 25136 18207 25188 18216
rect 25136 18173 25156 18207
rect 25156 18173 25188 18207
rect 25136 18164 25188 18173
rect 26424 18164 26476 18216
rect 26792 18164 26844 18216
rect 27160 18207 27212 18216
rect 27160 18173 27169 18207
rect 27169 18173 27203 18207
rect 27203 18173 27212 18207
rect 27160 18164 27212 18173
rect 27712 18207 27764 18216
rect 26884 18096 26936 18148
rect 27068 18096 27120 18148
rect 27712 18173 27721 18207
rect 27721 18173 27755 18207
rect 27755 18173 27764 18207
rect 27712 18164 27764 18173
rect 28632 18164 28684 18216
rect 29552 18232 29604 18284
rect 29644 18207 29696 18216
rect 29644 18173 29653 18207
rect 29653 18173 29687 18207
rect 29687 18173 29696 18207
rect 29644 18164 29696 18173
rect 32312 18309 32321 18343
rect 32321 18309 32355 18343
rect 32355 18309 32364 18343
rect 32312 18300 32364 18309
rect 30012 18232 30064 18284
rect 36912 18368 36964 18420
rect 37372 18368 37424 18420
rect 32680 18343 32732 18352
rect 32680 18309 32689 18343
rect 32689 18309 32723 18343
rect 32723 18309 32732 18343
rect 32680 18300 32732 18309
rect 31208 18207 31260 18216
rect 31208 18173 31217 18207
rect 31217 18173 31251 18207
rect 31251 18173 31260 18207
rect 32496 18207 32548 18216
rect 31208 18164 31260 18173
rect 32496 18173 32505 18207
rect 32505 18173 32539 18207
rect 32539 18173 32548 18207
rect 32496 18164 32548 18173
rect 33324 18232 33376 18284
rect 36084 18275 36136 18284
rect 36084 18241 36093 18275
rect 36093 18241 36127 18275
rect 36127 18241 36136 18275
rect 36084 18232 36136 18241
rect 36176 18232 36228 18284
rect 33048 18164 33100 18216
rect 33232 18207 33284 18216
rect 33232 18173 33241 18207
rect 33241 18173 33275 18207
rect 33275 18173 33284 18207
rect 33232 18164 33284 18173
rect 33508 18164 33560 18216
rect 35256 18207 35308 18216
rect 35256 18173 35265 18207
rect 35265 18173 35299 18207
rect 35299 18173 35308 18207
rect 35256 18164 35308 18173
rect 35440 18207 35492 18216
rect 35440 18173 35449 18207
rect 35449 18173 35483 18207
rect 35483 18173 35492 18207
rect 35440 18164 35492 18173
rect 35808 18164 35860 18216
rect 36452 18207 36504 18216
rect 36452 18173 36461 18207
rect 36461 18173 36495 18207
rect 36495 18173 36504 18207
rect 36452 18164 36504 18173
rect 37188 18207 37240 18216
rect 37188 18173 37197 18207
rect 37197 18173 37231 18207
rect 37231 18173 37240 18207
rect 37188 18164 37240 18173
rect 37648 18207 37700 18216
rect 37648 18173 37657 18207
rect 37657 18173 37691 18207
rect 37691 18173 37700 18207
rect 37648 18164 37700 18173
rect 29000 18028 29052 18080
rect 30564 18028 30616 18080
rect 32956 18096 33008 18148
rect 34520 18096 34572 18148
rect 33876 18028 33928 18080
rect 38292 18028 38344 18080
rect 19606 17926 19658 17978
rect 19670 17926 19722 17978
rect 19734 17926 19786 17978
rect 19798 17926 19850 17978
rect 9588 17824 9640 17876
rect 3148 17756 3200 17808
rect 8024 17756 8076 17808
rect 10784 17756 10836 17808
rect 1400 17731 1452 17740
rect 1400 17697 1409 17731
rect 1409 17697 1443 17731
rect 1443 17697 1452 17731
rect 1400 17688 1452 17697
rect 5264 17688 5316 17740
rect 7380 17688 7432 17740
rect 7932 17688 7984 17740
rect 8852 17688 8904 17740
rect 11428 17731 11480 17740
rect 11428 17697 11437 17731
rect 11437 17697 11471 17731
rect 11471 17697 11480 17731
rect 11428 17688 11480 17697
rect 11796 17731 11848 17740
rect 11796 17697 11805 17731
rect 11805 17697 11839 17731
rect 11839 17697 11848 17731
rect 11796 17688 11848 17697
rect 11980 17731 12032 17740
rect 11980 17697 11989 17731
rect 11989 17697 12023 17731
rect 12023 17697 12032 17731
rect 11980 17688 12032 17697
rect 12624 17731 12676 17740
rect 12624 17697 12633 17731
rect 12633 17697 12667 17731
rect 12667 17697 12676 17731
rect 12624 17688 12676 17697
rect 13176 17731 13228 17740
rect 13176 17697 13185 17731
rect 13185 17697 13219 17731
rect 13219 17697 13228 17731
rect 13176 17688 13228 17697
rect 15200 17688 15252 17740
rect 15844 17731 15896 17740
rect 15844 17697 15853 17731
rect 15853 17697 15887 17731
rect 15887 17697 15896 17731
rect 15844 17688 15896 17697
rect 4068 17620 4120 17672
rect 5448 17663 5500 17672
rect 5448 17629 5457 17663
rect 5457 17629 5491 17663
rect 5491 17629 5500 17663
rect 5448 17620 5500 17629
rect 6092 17663 6144 17672
rect 6092 17629 6101 17663
rect 6101 17629 6135 17663
rect 6135 17629 6144 17663
rect 6092 17620 6144 17629
rect 7196 17620 7248 17672
rect 8576 17595 8628 17604
rect 8576 17561 8585 17595
rect 8585 17561 8619 17595
rect 8619 17561 8628 17595
rect 8576 17552 8628 17561
rect 5080 17484 5132 17536
rect 11704 17620 11756 17672
rect 12716 17620 12768 17672
rect 11336 17552 11388 17604
rect 13268 17552 13320 17604
rect 15660 17620 15712 17672
rect 16212 17552 16264 17604
rect 17040 17552 17092 17604
rect 18052 17688 18104 17740
rect 22468 17824 22520 17876
rect 25872 17867 25924 17876
rect 25872 17833 25881 17867
rect 25881 17833 25915 17867
rect 25915 17833 25924 17867
rect 25872 17824 25924 17833
rect 19340 17756 19392 17808
rect 18788 17688 18840 17740
rect 19708 17688 19760 17740
rect 20168 17756 20220 17808
rect 26240 17756 26292 17808
rect 27068 17756 27120 17808
rect 28632 17756 28684 17808
rect 18696 17620 18748 17672
rect 22560 17688 22612 17740
rect 23848 17731 23900 17740
rect 23848 17697 23857 17731
rect 23857 17697 23891 17731
rect 23891 17697 23900 17731
rect 23848 17688 23900 17697
rect 24584 17688 24636 17740
rect 20536 17620 20588 17672
rect 21824 17620 21876 17672
rect 24768 17620 24820 17672
rect 19156 17552 19208 17604
rect 26884 17688 26936 17740
rect 27160 17688 27212 17740
rect 27436 17731 27488 17740
rect 27436 17697 27445 17731
rect 27445 17697 27479 17731
rect 27479 17697 27488 17731
rect 28540 17731 28592 17740
rect 27436 17688 27488 17697
rect 28540 17697 28549 17731
rect 28549 17697 28583 17731
rect 28583 17697 28592 17731
rect 28540 17688 28592 17697
rect 29000 17824 29052 17876
rect 29368 17824 29420 17876
rect 32588 17824 32640 17876
rect 29184 17756 29236 17808
rect 30656 17756 30708 17808
rect 33508 17824 33560 17876
rect 35900 17824 35952 17876
rect 37648 17824 37700 17876
rect 38016 17824 38068 17876
rect 28632 17663 28684 17672
rect 28632 17629 28641 17663
rect 28641 17629 28675 17663
rect 28675 17629 28684 17663
rect 28632 17620 28684 17629
rect 29368 17731 29420 17740
rect 29368 17697 29377 17731
rect 29377 17697 29411 17731
rect 29411 17697 29420 17731
rect 29368 17688 29420 17697
rect 29552 17731 29604 17740
rect 29552 17697 29561 17731
rect 29561 17697 29595 17731
rect 29595 17697 29604 17731
rect 29552 17688 29604 17697
rect 29644 17688 29696 17740
rect 30840 17731 30892 17740
rect 30840 17697 30849 17731
rect 30849 17697 30883 17731
rect 30883 17697 30892 17731
rect 30840 17688 30892 17697
rect 29276 17552 29328 17604
rect 30104 17552 30156 17604
rect 10324 17484 10376 17536
rect 15752 17484 15804 17536
rect 19064 17484 19116 17536
rect 22836 17484 22888 17536
rect 23388 17484 23440 17536
rect 23848 17484 23900 17536
rect 25412 17484 25464 17536
rect 26608 17484 26660 17536
rect 32312 17731 32364 17740
rect 32312 17697 32321 17731
rect 32321 17697 32355 17731
rect 32355 17697 32364 17731
rect 32312 17688 32364 17697
rect 32680 17688 32732 17740
rect 34796 17688 34848 17740
rect 35532 17688 35584 17740
rect 35900 17688 35952 17740
rect 36636 17688 36688 17740
rect 36728 17731 36780 17740
rect 36728 17697 36737 17731
rect 36737 17697 36771 17731
rect 36771 17697 36780 17731
rect 36728 17688 36780 17697
rect 31760 17620 31812 17672
rect 34152 17620 34204 17672
rect 34704 17620 34756 17672
rect 38660 17688 38712 17740
rect 38936 17731 38988 17740
rect 38936 17697 38945 17731
rect 38945 17697 38979 17731
rect 38979 17697 38988 17731
rect 38936 17688 38988 17697
rect 36360 17552 36412 17604
rect 32772 17484 32824 17536
rect 37464 17484 37516 17536
rect 4246 17382 4298 17434
rect 4310 17382 4362 17434
rect 4374 17382 4426 17434
rect 4438 17382 4490 17434
rect 34966 17382 35018 17434
rect 35030 17382 35082 17434
rect 35094 17382 35146 17434
rect 35158 17382 35210 17434
rect 2872 17280 2924 17332
rect 1400 17187 1452 17196
rect 1400 17153 1409 17187
rect 1409 17153 1443 17187
rect 1443 17153 1452 17187
rect 1400 17144 1452 17153
rect 8852 17323 8904 17332
rect 8852 17289 8861 17323
rect 8861 17289 8895 17323
rect 8895 17289 8904 17323
rect 8852 17280 8904 17289
rect 9036 17280 9088 17332
rect 15844 17280 15896 17332
rect 16212 17280 16264 17332
rect 26148 17280 26200 17332
rect 32772 17280 32824 17332
rect 32956 17280 33008 17332
rect 35440 17280 35492 17332
rect 4712 17144 4764 17196
rect 5080 17144 5132 17196
rect 6828 17144 6880 17196
rect 12440 17187 12492 17196
rect 12440 17153 12449 17187
rect 12449 17153 12483 17187
rect 12483 17153 12492 17187
rect 12440 17144 12492 17153
rect 12716 17187 12768 17196
rect 12716 17153 12725 17187
rect 12725 17153 12759 17187
rect 12759 17153 12768 17187
rect 12716 17144 12768 17153
rect 13820 17144 13872 17196
rect 15476 17144 15528 17196
rect 2504 17076 2556 17128
rect 5540 17076 5592 17128
rect 7564 17119 7616 17128
rect 7564 17085 7573 17119
rect 7573 17085 7607 17119
rect 7607 17085 7616 17119
rect 7564 17076 7616 17085
rect 8576 17076 8628 17128
rect 11520 17076 11572 17128
rect 11796 17076 11848 17128
rect 10600 16940 10652 16992
rect 10692 16940 10744 16992
rect 13820 16983 13872 16992
rect 13820 16949 13829 16983
rect 13829 16949 13863 16983
rect 13863 16949 13872 16983
rect 13820 16940 13872 16949
rect 19064 17212 19116 17264
rect 19432 17212 19484 17264
rect 19708 17212 19760 17264
rect 16120 17144 16172 17196
rect 29000 17212 29052 17264
rect 26148 17187 26200 17196
rect 17316 17119 17368 17128
rect 17316 17085 17325 17119
rect 17325 17085 17359 17119
rect 17359 17085 17368 17119
rect 17316 17076 17368 17085
rect 18328 17119 18380 17128
rect 18328 17085 18337 17119
rect 18337 17085 18371 17119
rect 18371 17085 18380 17119
rect 18328 17076 18380 17085
rect 19340 17076 19392 17128
rect 19984 17076 20036 17128
rect 20076 17076 20128 17128
rect 20720 17119 20772 17128
rect 20720 17085 20729 17119
rect 20729 17085 20763 17119
rect 20763 17085 20772 17119
rect 20720 17076 20772 17085
rect 21272 17119 21324 17128
rect 21272 17085 21281 17119
rect 21281 17085 21315 17119
rect 21315 17085 21324 17119
rect 21272 17076 21324 17085
rect 26148 17153 26157 17187
rect 26157 17153 26191 17187
rect 26191 17153 26200 17187
rect 26148 17144 26200 17153
rect 27252 17144 27304 17196
rect 22836 17119 22888 17128
rect 22836 17085 22845 17119
rect 22845 17085 22879 17119
rect 22879 17085 22888 17119
rect 22836 17076 22888 17085
rect 24032 17119 24084 17128
rect 24032 17085 24041 17119
rect 24041 17085 24075 17119
rect 24075 17085 24084 17119
rect 24032 17076 24084 17085
rect 24308 17119 24360 17128
rect 24308 17085 24317 17119
rect 24317 17085 24351 17119
rect 24351 17085 24360 17119
rect 24308 17076 24360 17085
rect 27620 17119 27672 17128
rect 17224 16940 17276 16992
rect 21272 16940 21324 16992
rect 22192 16983 22244 16992
rect 22192 16949 22201 16983
rect 22201 16949 22235 16983
rect 22235 16949 22244 16983
rect 22192 16940 22244 16949
rect 22560 16940 22612 16992
rect 27620 17085 27629 17119
rect 27629 17085 27663 17119
rect 27663 17085 27672 17119
rect 27620 17076 27672 17085
rect 27804 17144 27856 17196
rect 32588 17212 32640 17264
rect 29552 17144 29604 17196
rect 30380 17076 30432 17128
rect 30656 17119 30708 17128
rect 30656 17085 30665 17119
rect 30665 17085 30699 17119
rect 30699 17085 30708 17119
rect 30656 17076 30708 17085
rect 31300 17119 31352 17128
rect 31300 17085 31309 17119
rect 31309 17085 31343 17119
rect 31343 17085 31352 17119
rect 31300 17076 31352 17085
rect 32036 17144 32088 17196
rect 33048 17144 33100 17196
rect 31760 17119 31812 17128
rect 31760 17085 31769 17119
rect 31769 17085 31803 17119
rect 31803 17085 31812 17119
rect 31760 17076 31812 17085
rect 33784 17119 33836 17128
rect 33784 17085 33793 17119
rect 33793 17085 33827 17119
rect 33827 17085 33836 17119
rect 33784 17076 33836 17085
rect 34152 17119 34204 17128
rect 34152 17085 34161 17119
rect 34161 17085 34195 17119
rect 34195 17085 34204 17119
rect 34152 17076 34204 17085
rect 34796 17076 34848 17128
rect 35716 17144 35768 17196
rect 38936 17280 38988 17332
rect 38476 17212 38528 17264
rect 38200 17144 38252 17196
rect 27896 17008 27948 17060
rect 30288 17008 30340 17060
rect 30472 17051 30524 17060
rect 30472 17017 30481 17051
rect 30481 17017 30515 17051
rect 30515 17017 30524 17051
rect 30472 17008 30524 17017
rect 36268 17008 36320 17060
rect 24952 16940 25004 16992
rect 26424 16940 26476 16992
rect 26792 16940 26844 16992
rect 28264 16940 28316 16992
rect 28816 16940 28868 16992
rect 32128 16940 32180 16992
rect 34060 16940 34112 16992
rect 36176 16940 36228 16992
rect 36360 16940 36412 16992
rect 37464 17119 37516 17128
rect 37464 17085 37473 17119
rect 37473 17085 37507 17119
rect 37507 17085 37516 17119
rect 37464 17076 37516 17085
rect 38568 17076 38620 17128
rect 38660 16940 38712 16992
rect 19606 16838 19658 16890
rect 19670 16838 19722 16890
rect 19734 16838 19786 16890
rect 19798 16838 19850 16890
rect 1952 16779 2004 16788
rect 1952 16745 1961 16779
rect 1961 16745 1995 16779
rect 1995 16745 2004 16779
rect 1952 16736 2004 16745
rect 2504 16779 2556 16788
rect 2504 16745 2513 16779
rect 2513 16745 2547 16779
rect 2547 16745 2556 16779
rect 2504 16736 2556 16745
rect 5264 16779 5316 16788
rect 1768 16643 1820 16652
rect 1768 16609 1777 16643
rect 1777 16609 1811 16643
rect 1811 16609 1820 16643
rect 1768 16600 1820 16609
rect 5264 16745 5273 16779
rect 5273 16745 5307 16779
rect 5307 16745 5316 16779
rect 5264 16736 5316 16745
rect 6276 16668 6328 16720
rect 4620 16600 4672 16652
rect 4712 16600 4764 16652
rect 5724 16643 5776 16652
rect 5724 16609 5733 16643
rect 5733 16609 5767 16643
rect 5767 16609 5776 16643
rect 5724 16600 5776 16609
rect 6552 16643 6604 16652
rect 6552 16609 6561 16643
rect 6561 16609 6595 16643
rect 6595 16609 6604 16643
rect 6552 16600 6604 16609
rect 10692 16736 10744 16788
rect 7564 16668 7616 16720
rect 5356 16464 5408 16516
rect 7288 16600 7340 16652
rect 9036 16668 9088 16720
rect 10876 16668 10928 16720
rect 11796 16736 11848 16788
rect 15660 16736 15712 16788
rect 15844 16736 15896 16788
rect 16212 16779 16264 16788
rect 16212 16745 16221 16779
rect 16221 16745 16255 16779
rect 16255 16745 16264 16779
rect 16212 16736 16264 16745
rect 19984 16736 20036 16788
rect 13820 16668 13872 16720
rect 23572 16736 23624 16788
rect 26792 16736 26844 16788
rect 30840 16736 30892 16788
rect 31760 16736 31812 16788
rect 8116 16532 8168 16584
rect 9128 16575 9180 16584
rect 9128 16541 9137 16575
rect 9137 16541 9171 16575
rect 9171 16541 9180 16575
rect 9128 16532 9180 16541
rect 10048 16643 10100 16652
rect 10048 16609 10057 16643
rect 10057 16609 10091 16643
rect 10091 16609 10100 16643
rect 10416 16643 10468 16652
rect 10048 16600 10100 16609
rect 10416 16609 10425 16643
rect 10425 16609 10459 16643
rect 10459 16609 10468 16643
rect 10416 16600 10468 16609
rect 11336 16643 11388 16652
rect 11336 16609 11345 16643
rect 11345 16609 11379 16643
rect 11379 16609 11388 16643
rect 11336 16600 11388 16609
rect 12440 16643 12492 16652
rect 12440 16609 12449 16643
rect 12449 16609 12483 16643
rect 12483 16609 12492 16643
rect 12440 16600 12492 16609
rect 14004 16600 14056 16652
rect 15292 16643 15344 16652
rect 15292 16609 15301 16643
rect 15301 16609 15335 16643
rect 15335 16609 15344 16643
rect 15292 16600 15344 16609
rect 17040 16643 17092 16652
rect 17040 16609 17049 16643
rect 17049 16609 17083 16643
rect 17083 16609 17092 16643
rect 17040 16600 17092 16609
rect 19156 16643 19208 16652
rect 19156 16609 19165 16643
rect 19165 16609 19199 16643
rect 19199 16609 19208 16643
rect 19156 16600 19208 16609
rect 20352 16600 20404 16652
rect 20536 16600 20588 16652
rect 22192 16668 22244 16720
rect 21916 16643 21968 16652
rect 21916 16609 21925 16643
rect 21925 16609 21959 16643
rect 21959 16609 21968 16643
rect 21916 16600 21968 16609
rect 22376 16643 22428 16652
rect 22376 16609 22385 16643
rect 22385 16609 22419 16643
rect 22419 16609 22428 16643
rect 22376 16600 22428 16609
rect 22652 16643 22704 16652
rect 22652 16609 22661 16643
rect 22661 16609 22695 16643
rect 22695 16609 22704 16643
rect 22652 16600 22704 16609
rect 23388 16643 23440 16652
rect 23388 16609 23397 16643
rect 23397 16609 23431 16643
rect 23431 16609 23440 16643
rect 23388 16600 23440 16609
rect 23480 16600 23532 16652
rect 26608 16600 26660 16652
rect 26792 16643 26844 16652
rect 26792 16609 26801 16643
rect 26801 16609 26835 16643
rect 26835 16609 26844 16643
rect 26792 16600 26844 16609
rect 27344 16668 27396 16720
rect 33416 16736 33468 16788
rect 27252 16600 27304 16652
rect 27804 16643 27856 16652
rect 27804 16609 27813 16643
rect 27813 16609 27847 16643
rect 27847 16609 27856 16643
rect 27804 16600 27856 16609
rect 28264 16643 28316 16652
rect 28264 16609 28273 16643
rect 28273 16609 28307 16643
rect 28307 16609 28316 16643
rect 28264 16600 28316 16609
rect 28632 16600 28684 16652
rect 30288 16600 30340 16652
rect 32220 16600 32272 16652
rect 32404 16600 32456 16652
rect 33692 16643 33744 16652
rect 33692 16609 33701 16643
rect 33701 16609 33735 16643
rect 33735 16609 33744 16643
rect 33692 16600 33744 16609
rect 34612 16600 34664 16652
rect 36176 16736 36228 16788
rect 38016 16736 38068 16788
rect 38292 16668 38344 16720
rect 38568 16711 38620 16720
rect 38568 16677 38577 16711
rect 38577 16677 38611 16711
rect 38611 16677 38620 16711
rect 38568 16668 38620 16677
rect 35900 16600 35952 16652
rect 36636 16643 36688 16652
rect 36636 16609 36645 16643
rect 36645 16609 36679 16643
rect 36679 16609 36688 16643
rect 36636 16600 36688 16609
rect 36820 16643 36872 16652
rect 36820 16609 36829 16643
rect 36829 16609 36863 16643
rect 36863 16609 36872 16643
rect 36820 16600 36872 16609
rect 38660 16600 38712 16652
rect 16764 16575 16816 16584
rect 16764 16541 16773 16575
rect 16773 16541 16807 16575
rect 16807 16541 16816 16575
rect 16764 16532 16816 16541
rect 17776 16532 17828 16584
rect 21824 16575 21876 16584
rect 21824 16541 21833 16575
rect 21833 16541 21867 16575
rect 21867 16541 21876 16575
rect 21824 16532 21876 16541
rect 22468 16532 22520 16584
rect 23296 16532 23348 16584
rect 24032 16575 24084 16584
rect 24032 16541 24041 16575
rect 24041 16541 24075 16575
rect 24075 16541 24084 16575
rect 24032 16532 24084 16541
rect 26884 16575 26936 16584
rect 26884 16541 26893 16575
rect 26893 16541 26927 16575
rect 26927 16541 26936 16575
rect 26884 16532 26936 16541
rect 29092 16532 29144 16584
rect 30104 16532 30156 16584
rect 37556 16532 37608 16584
rect 38384 16532 38436 16584
rect 4068 16396 4120 16448
rect 10048 16396 10100 16448
rect 13912 16396 13964 16448
rect 23388 16464 23440 16516
rect 17960 16396 18012 16448
rect 19340 16439 19392 16448
rect 19340 16405 19349 16439
rect 19349 16405 19383 16439
rect 19383 16405 19392 16439
rect 19340 16396 19392 16405
rect 19432 16396 19484 16448
rect 21640 16396 21692 16448
rect 23572 16396 23624 16448
rect 24216 16396 24268 16448
rect 30288 16439 30340 16448
rect 30288 16405 30297 16439
rect 30297 16405 30331 16439
rect 30331 16405 30340 16439
rect 30288 16396 30340 16405
rect 34796 16396 34848 16448
rect 4246 16294 4298 16346
rect 4310 16294 4362 16346
rect 4374 16294 4426 16346
rect 4438 16294 4490 16346
rect 34966 16294 35018 16346
rect 35030 16294 35082 16346
rect 35094 16294 35146 16346
rect 35158 16294 35210 16346
rect 4620 16192 4672 16244
rect 11336 16192 11388 16244
rect 18328 16192 18380 16244
rect 7104 16167 7156 16176
rect 7104 16133 7113 16167
rect 7113 16133 7147 16167
rect 7147 16133 7156 16167
rect 7104 16124 7156 16133
rect 14004 16167 14056 16176
rect 2504 16056 2556 16108
rect 5264 16056 5316 16108
rect 5540 16056 5592 16108
rect 9128 16056 9180 16108
rect 14004 16133 14013 16167
rect 14013 16133 14047 16167
rect 14047 16133 14056 16167
rect 14004 16124 14056 16133
rect 5356 16031 5408 16040
rect 5356 15997 5365 16031
rect 5365 15997 5399 16031
rect 5399 15997 5408 16031
rect 5356 15988 5408 15997
rect 6184 15988 6236 16040
rect 7380 16031 7432 16040
rect 6000 15920 6052 15972
rect 7380 15997 7389 16031
rect 7389 15997 7423 16031
rect 7423 15997 7432 16031
rect 7380 15988 7432 15997
rect 7564 16031 7616 16040
rect 7564 15997 7573 16031
rect 7573 15997 7607 16031
rect 7607 15997 7616 16031
rect 7564 15988 7616 15997
rect 8208 16031 8260 16040
rect 8208 15997 8217 16031
rect 8217 15997 8251 16031
rect 8251 15997 8260 16031
rect 8208 15988 8260 15997
rect 9036 15988 9088 16040
rect 9404 16031 9456 16040
rect 9404 15997 9413 16031
rect 9413 15997 9447 16031
rect 9447 15997 9456 16031
rect 9404 15988 9456 15997
rect 11520 16031 11572 16040
rect 11520 15997 11529 16031
rect 11529 15997 11563 16031
rect 11563 15997 11572 16031
rect 11520 15988 11572 15997
rect 12808 16031 12860 16040
rect 12808 15997 12817 16031
rect 12817 15997 12851 16031
rect 12851 15997 12860 16031
rect 12808 15988 12860 15997
rect 13452 16031 13504 16040
rect 13452 15997 13461 16031
rect 13461 15997 13495 16031
rect 13495 15997 13504 16031
rect 13452 15988 13504 15997
rect 14280 15988 14332 16040
rect 14556 16031 14608 16040
rect 14556 15997 14565 16031
rect 14565 15997 14599 16031
rect 14599 15997 14608 16031
rect 14556 15988 14608 15997
rect 16120 16124 16172 16176
rect 18052 16124 18104 16176
rect 21364 16124 21416 16176
rect 21916 16124 21968 16176
rect 19984 16099 20036 16108
rect 19984 16065 19993 16099
rect 19993 16065 20027 16099
rect 20027 16065 20036 16099
rect 19984 16056 20036 16065
rect 22376 16056 22428 16108
rect 34612 16192 34664 16244
rect 38936 16192 38988 16244
rect 15936 15988 15988 16040
rect 17960 15988 18012 16040
rect 18420 15988 18472 16040
rect 19340 15988 19392 16040
rect 20260 16031 20312 16040
rect 11428 15852 11480 15904
rect 13176 15852 13228 15904
rect 19432 15920 19484 15972
rect 18788 15895 18840 15904
rect 18788 15861 18797 15895
rect 18797 15861 18831 15895
rect 18831 15861 18840 15895
rect 18788 15852 18840 15861
rect 20260 15997 20269 16031
rect 20269 15997 20303 16031
rect 20303 15997 20312 16031
rect 20260 15988 20312 15997
rect 20720 16031 20772 16040
rect 20720 15997 20729 16031
rect 20729 15997 20763 16031
rect 20763 15997 20772 16031
rect 20720 15988 20772 15997
rect 20996 15988 21048 16040
rect 21180 15988 21232 16040
rect 22468 15988 22520 16040
rect 23480 16056 23532 16108
rect 24308 16099 24360 16108
rect 24308 16065 24317 16099
rect 24317 16065 24351 16099
rect 24351 16065 24360 16099
rect 24308 16056 24360 16065
rect 28908 16124 28960 16176
rect 26884 16056 26936 16108
rect 30472 16056 30524 16108
rect 23664 16031 23716 16040
rect 21824 15920 21876 15972
rect 23664 15997 23673 16031
rect 23673 15997 23707 16031
rect 23707 15997 23716 16031
rect 23664 15988 23716 15997
rect 24216 16031 24268 16040
rect 24216 15997 24225 16031
rect 24225 15997 24259 16031
rect 24259 15997 24268 16031
rect 24216 15988 24268 15997
rect 26516 15920 26568 15972
rect 27620 15988 27672 16040
rect 28080 16031 28132 16040
rect 28080 15997 28089 16031
rect 28089 15997 28123 16031
rect 28123 15997 28132 16031
rect 28080 15988 28132 15997
rect 28264 16031 28316 16040
rect 28264 15997 28273 16031
rect 28273 15997 28307 16031
rect 28307 15997 28316 16031
rect 28264 15988 28316 15997
rect 30104 15988 30156 16040
rect 32312 16056 32364 16108
rect 32404 16031 32456 16040
rect 32404 15997 32413 16031
rect 32413 15997 32447 16031
rect 32447 15997 32456 16031
rect 32404 15988 32456 15997
rect 34796 16056 34848 16108
rect 35900 16056 35952 16108
rect 37556 16099 37608 16108
rect 33508 16031 33560 16040
rect 33508 15997 33517 16031
rect 33517 15997 33551 16031
rect 33551 15997 33560 16031
rect 33508 15988 33560 15997
rect 35808 15988 35860 16040
rect 35992 16031 36044 16040
rect 35992 15997 36001 16031
rect 36001 15997 36035 16031
rect 36035 15997 36044 16031
rect 35992 15988 36044 15997
rect 37556 16065 37565 16099
rect 37565 16065 37599 16099
rect 37599 16065 37608 16099
rect 37556 16056 37608 16065
rect 34704 15920 34756 15972
rect 20536 15852 20588 15904
rect 20996 15852 21048 15904
rect 21272 15852 21324 15904
rect 21640 15852 21692 15904
rect 22928 15852 22980 15904
rect 23388 15852 23440 15904
rect 30104 15852 30156 15904
rect 31668 15895 31720 15904
rect 31668 15861 31677 15895
rect 31677 15861 31711 15895
rect 31711 15861 31720 15895
rect 31668 15852 31720 15861
rect 32220 15852 32272 15904
rect 34336 15852 34388 15904
rect 37372 15988 37424 16040
rect 19606 15750 19658 15802
rect 19670 15750 19722 15802
rect 19734 15750 19786 15802
rect 19798 15750 19850 15802
rect 1400 15555 1452 15564
rect 1400 15521 1409 15555
rect 1409 15521 1443 15555
rect 1443 15521 1452 15555
rect 1400 15512 1452 15521
rect 7196 15648 7248 15700
rect 13912 15648 13964 15700
rect 7932 15580 7984 15632
rect 8208 15580 8260 15632
rect 2504 15512 2556 15564
rect 2688 15512 2740 15564
rect 12624 15580 12676 15632
rect 12808 15580 12860 15632
rect 14464 15648 14516 15700
rect 14556 15648 14608 15700
rect 16120 15648 16172 15700
rect 21180 15648 21232 15700
rect 28724 15648 28776 15700
rect 18420 15623 18472 15632
rect 8392 15512 8444 15564
rect 10876 15555 10928 15564
rect 10876 15521 10885 15555
rect 10885 15521 10919 15555
rect 10919 15521 10928 15555
rect 10876 15512 10928 15521
rect 11428 15555 11480 15564
rect 11428 15521 11437 15555
rect 11437 15521 11471 15555
rect 11471 15521 11480 15555
rect 11428 15512 11480 15521
rect 11796 15555 11848 15564
rect 11796 15521 11805 15555
rect 11805 15521 11839 15555
rect 11839 15521 11848 15555
rect 11796 15512 11848 15521
rect 11980 15512 12032 15564
rect 5172 15444 5224 15496
rect 6828 15444 6880 15496
rect 7564 15444 7616 15496
rect 2872 15308 2924 15360
rect 8208 15308 8260 15360
rect 11888 15444 11940 15496
rect 11612 15419 11664 15428
rect 11612 15385 11621 15419
rect 11621 15385 11655 15419
rect 11655 15385 11664 15419
rect 11612 15376 11664 15385
rect 13636 15308 13688 15360
rect 14648 15512 14700 15564
rect 18420 15589 18429 15623
rect 18429 15589 18463 15623
rect 18463 15589 18472 15623
rect 18420 15580 18472 15589
rect 18788 15580 18840 15632
rect 16764 15555 16816 15564
rect 16764 15521 16773 15555
rect 16773 15521 16807 15555
rect 16807 15521 16816 15555
rect 16764 15512 16816 15521
rect 16304 15444 16356 15496
rect 18972 15512 19024 15564
rect 19156 15512 19208 15564
rect 20536 15512 20588 15564
rect 22100 15512 22152 15564
rect 22376 15512 22428 15564
rect 22468 15555 22520 15564
rect 22468 15521 22477 15555
rect 22477 15521 22511 15555
rect 22511 15521 22520 15555
rect 22468 15512 22520 15521
rect 22652 15512 22704 15564
rect 23664 15555 23716 15564
rect 23664 15521 23673 15555
rect 23673 15521 23707 15555
rect 23707 15521 23716 15555
rect 23664 15512 23716 15521
rect 26608 15555 26660 15564
rect 15108 15376 15160 15428
rect 15476 15376 15528 15428
rect 18880 15487 18932 15496
rect 18880 15453 18889 15487
rect 18889 15453 18923 15487
rect 18923 15453 18932 15487
rect 18880 15444 18932 15453
rect 22192 15487 22244 15496
rect 22192 15453 22201 15487
rect 22201 15453 22235 15487
rect 22235 15453 22244 15487
rect 22192 15444 22244 15453
rect 23020 15444 23072 15496
rect 26608 15521 26617 15555
rect 26617 15521 26651 15555
rect 26651 15521 26660 15555
rect 26608 15512 26660 15521
rect 28724 15512 28776 15564
rect 29184 15512 29236 15564
rect 24400 15487 24452 15496
rect 24400 15453 24409 15487
rect 24409 15453 24443 15487
rect 24443 15453 24452 15487
rect 24400 15444 24452 15453
rect 26148 15444 26200 15496
rect 29000 15444 29052 15496
rect 30104 15648 30156 15700
rect 33508 15648 33560 15700
rect 33600 15648 33652 15700
rect 34428 15648 34480 15700
rect 30104 15512 30156 15564
rect 31852 15512 31904 15564
rect 32036 15512 32088 15564
rect 32772 15555 32824 15564
rect 32772 15521 32781 15555
rect 32781 15521 32815 15555
rect 32815 15521 32824 15555
rect 32772 15512 32824 15521
rect 34336 15512 34388 15564
rect 34520 15555 34572 15564
rect 34520 15521 34529 15555
rect 34529 15521 34563 15555
rect 34563 15521 34572 15555
rect 34520 15512 34572 15521
rect 35900 15648 35952 15700
rect 36636 15648 36688 15700
rect 37924 15555 37976 15564
rect 37924 15521 37933 15555
rect 37933 15521 37967 15555
rect 37967 15521 37976 15555
rect 37924 15512 37976 15521
rect 38476 15555 38528 15564
rect 38476 15521 38485 15555
rect 38485 15521 38519 15555
rect 38519 15521 38528 15555
rect 38476 15512 38528 15521
rect 28540 15376 28592 15428
rect 22284 15308 22336 15360
rect 27160 15308 27212 15360
rect 31944 15444 31996 15496
rect 32312 15444 32364 15496
rect 37372 15444 37424 15496
rect 38384 15487 38436 15496
rect 38384 15453 38393 15487
rect 38393 15453 38427 15487
rect 38427 15453 38436 15487
rect 38384 15444 38436 15453
rect 30380 15376 30432 15428
rect 32220 15376 32272 15428
rect 33324 15376 33376 15428
rect 31392 15308 31444 15360
rect 31484 15351 31536 15360
rect 31484 15317 31493 15351
rect 31493 15317 31527 15351
rect 31527 15317 31536 15351
rect 31484 15308 31536 15317
rect 37924 15308 37976 15360
rect 4246 15206 4298 15258
rect 4310 15206 4362 15258
rect 4374 15206 4426 15258
rect 4438 15206 4490 15258
rect 34966 15206 35018 15258
rect 35030 15206 35082 15258
rect 35094 15206 35146 15258
rect 35158 15206 35210 15258
rect 4068 15104 4120 15156
rect 5172 15147 5224 15156
rect 5172 15113 5181 15147
rect 5181 15113 5215 15147
rect 5215 15113 5224 15147
rect 5172 15104 5224 15113
rect 8392 15147 8444 15156
rect 8392 15113 8401 15147
rect 8401 15113 8435 15147
rect 8435 15113 8444 15147
rect 8392 15104 8444 15113
rect 9220 15104 9272 15156
rect 9404 15104 9456 15156
rect 11428 15104 11480 15156
rect 12440 15104 12492 15156
rect 12900 15104 12952 15156
rect 17500 15104 17552 15156
rect 19432 15104 19484 15156
rect 19892 15104 19944 15156
rect 20168 15104 20220 15156
rect 20536 15104 20588 15156
rect 21824 15147 21876 15156
rect 21824 15113 21833 15147
rect 21833 15113 21867 15147
rect 21867 15113 21876 15147
rect 21824 15104 21876 15113
rect 29000 15104 29052 15156
rect 30288 15104 30340 15156
rect 31392 15104 31444 15156
rect 33232 15104 33284 15156
rect 38108 15104 38160 15156
rect 12164 15036 12216 15088
rect 7104 15011 7156 15020
rect 7104 14977 7113 15011
rect 7113 14977 7147 15011
rect 7147 14977 7156 15011
rect 7104 14968 7156 14977
rect 13176 14968 13228 15020
rect 1400 14900 1452 14952
rect 1952 14943 2004 14952
rect 1952 14909 1961 14943
rect 1961 14909 1995 14943
rect 1995 14909 2004 14943
rect 1952 14900 2004 14909
rect 2688 14900 2740 14952
rect 6828 14943 6880 14952
rect 6828 14909 6837 14943
rect 6837 14909 6871 14943
rect 6871 14909 6880 14943
rect 6828 14900 6880 14909
rect 7564 14900 7616 14952
rect 8852 14900 8904 14952
rect 9772 14943 9824 14952
rect 6736 14764 6788 14816
rect 6920 14764 6972 14816
rect 9220 14764 9272 14816
rect 9772 14909 9781 14943
rect 9781 14909 9815 14943
rect 9815 14909 9824 14943
rect 9772 14900 9824 14909
rect 10692 14943 10744 14952
rect 10692 14909 10701 14943
rect 10701 14909 10735 14943
rect 10735 14909 10744 14943
rect 10692 14900 10744 14909
rect 11060 14943 11112 14952
rect 11060 14909 11069 14943
rect 11069 14909 11103 14943
rect 11103 14909 11112 14943
rect 11060 14900 11112 14909
rect 11336 14943 11388 14952
rect 11336 14909 11345 14943
rect 11345 14909 11379 14943
rect 11379 14909 11388 14943
rect 11336 14900 11388 14909
rect 12072 14943 12124 14952
rect 12072 14909 12081 14943
rect 12081 14909 12115 14943
rect 12115 14909 12124 14943
rect 12072 14900 12124 14909
rect 12440 14943 12492 14952
rect 12440 14909 12449 14943
rect 12449 14909 12483 14943
rect 12483 14909 12492 14943
rect 13820 15036 13872 15088
rect 30012 15036 30064 15088
rect 14096 14968 14148 15020
rect 12440 14900 12492 14909
rect 14004 14900 14056 14952
rect 14556 14943 14608 14952
rect 14556 14909 14565 14943
rect 14565 14909 14599 14943
rect 14599 14909 14608 14943
rect 14556 14900 14608 14909
rect 17040 14968 17092 15020
rect 18328 14968 18380 15020
rect 15292 14900 15344 14952
rect 16764 14900 16816 14952
rect 16948 14943 17000 14952
rect 16948 14909 16957 14943
rect 16957 14909 16991 14943
rect 16991 14909 17000 14943
rect 16948 14900 17000 14909
rect 18236 14943 18288 14952
rect 9404 14832 9456 14884
rect 18236 14909 18245 14943
rect 18245 14909 18279 14943
rect 18279 14909 18288 14943
rect 18236 14900 18288 14909
rect 19340 14943 19392 14952
rect 11244 14764 11296 14816
rect 11336 14764 11388 14816
rect 11796 14764 11848 14816
rect 13544 14764 13596 14816
rect 18052 14832 18104 14884
rect 19340 14909 19349 14943
rect 19349 14909 19383 14943
rect 19383 14909 19392 14943
rect 19340 14900 19392 14909
rect 20168 14968 20220 15020
rect 21272 14968 21324 15020
rect 24308 14968 24360 15020
rect 24492 14968 24544 15020
rect 24768 14968 24820 15020
rect 26516 15011 26568 15020
rect 26516 14977 26525 15011
rect 26525 14977 26559 15011
rect 26559 14977 26568 15011
rect 26516 14968 26568 14977
rect 28908 14968 28960 15020
rect 31576 14968 31628 15020
rect 33048 15011 33100 15020
rect 33048 14977 33057 15011
rect 33057 14977 33091 15011
rect 33091 14977 33100 15011
rect 33048 14968 33100 14977
rect 37372 14968 37424 15020
rect 20720 14943 20772 14952
rect 20720 14909 20729 14943
rect 20729 14909 20763 14943
rect 20763 14909 20772 14943
rect 20720 14900 20772 14909
rect 20996 14943 21048 14952
rect 20996 14909 21005 14943
rect 21005 14909 21039 14943
rect 21039 14909 21048 14943
rect 20996 14900 21048 14909
rect 21088 14900 21140 14952
rect 22928 14943 22980 14952
rect 22928 14909 22937 14943
rect 22937 14909 22971 14943
rect 22971 14909 22980 14943
rect 22928 14900 22980 14909
rect 24124 14943 24176 14952
rect 24124 14909 24133 14943
rect 24133 14909 24167 14943
rect 24167 14909 24176 14943
rect 24124 14900 24176 14909
rect 24860 14900 24912 14952
rect 22836 14832 22888 14884
rect 27896 14875 27948 14884
rect 27896 14841 27905 14875
rect 27905 14841 27939 14875
rect 27939 14841 27948 14875
rect 27896 14832 27948 14841
rect 28356 14832 28408 14884
rect 17132 14764 17184 14816
rect 17408 14764 17460 14816
rect 22100 14764 22152 14816
rect 23020 14807 23072 14816
rect 23020 14773 23029 14807
rect 23029 14773 23063 14807
rect 23063 14773 23072 14807
rect 23020 14764 23072 14773
rect 26608 14764 26660 14816
rect 28908 14764 28960 14816
rect 29184 14900 29236 14952
rect 30104 14900 30156 14952
rect 30564 14900 30616 14952
rect 30748 14900 30800 14952
rect 31668 14900 31720 14952
rect 32312 14943 32364 14952
rect 32312 14909 32321 14943
rect 32321 14909 32355 14943
rect 32355 14909 32364 14943
rect 32312 14900 32364 14909
rect 32772 14943 32824 14952
rect 32220 14832 32272 14884
rect 32772 14909 32781 14943
rect 32781 14909 32815 14943
rect 32815 14909 32824 14943
rect 32772 14900 32824 14909
rect 33600 14900 33652 14952
rect 33784 14900 33836 14952
rect 36084 14943 36136 14952
rect 35808 14832 35860 14884
rect 34520 14764 34572 14816
rect 36084 14909 36093 14943
rect 36093 14909 36127 14943
rect 36127 14909 36136 14943
rect 36084 14900 36136 14909
rect 36268 14943 36320 14952
rect 36268 14909 36277 14943
rect 36277 14909 36311 14943
rect 36311 14909 36320 14943
rect 36268 14900 36320 14909
rect 37740 14943 37792 14952
rect 37740 14909 37749 14943
rect 37749 14909 37783 14943
rect 37783 14909 37792 14943
rect 37740 14900 37792 14909
rect 38476 14764 38528 14816
rect 19606 14662 19658 14714
rect 19670 14662 19722 14714
rect 19734 14662 19786 14714
rect 19798 14662 19850 14714
rect 1952 14560 2004 14612
rect 9496 14560 9548 14612
rect 13544 14603 13596 14612
rect 1676 14467 1728 14476
rect 1676 14433 1685 14467
rect 1685 14433 1719 14467
rect 1719 14433 1728 14467
rect 1676 14424 1728 14433
rect 3884 14467 3936 14476
rect 3884 14433 3893 14467
rect 3893 14433 3927 14467
rect 3927 14433 3936 14467
rect 3884 14424 3936 14433
rect 6920 14424 6972 14476
rect 10692 14492 10744 14544
rect 9956 14467 10008 14476
rect 9956 14433 9965 14467
rect 9965 14433 9999 14467
rect 9999 14433 10008 14467
rect 9956 14424 10008 14433
rect 10048 14467 10100 14476
rect 10048 14433 10057 14467
rect 10057 14433 10091 14467
rect 10091 14433 10100 14467
rect 10416 14467 10468 14476
rect 10048 14424 10100 14433
rect 10416 14433 10425 14467
rect 10425 14433 10459 14467
rect 10459 14433 10468 14467
rect 10416 14424 10468 14433
rect 11428 14424 11480 14476
rect 11612 14467 11664 14476
rect 11612 14433 11621 14467
rect 11621 14433 11655 14467
rect 11655 14433 11664 14467
rect 11612 14424 11664 14433
rect 13544 14569 13553 14603
rect 13553 14569 13587 14603
rect 13587 14569 13596 14603
rect 13544 14560 13596 14569
rect 14556 14560 14608 14612
rect 22928 14560 22980 14612
rect 24676 14560 24728 14612
rect 27804 14560 27856 14612
rect 29828 14560 29880 14612
rect 28080 14492 28132 14544
rect 31208 14492 31260 14544
rect 13544 14424 13596 14476
rect 13728 14424 13780 14476
rect 13912 14424 13964 14476
rect 15384 14424 15436 14476
rect 15660 14424 15712 14476
rect 15936 14467 15988 14476
rect 15936 14433 15945 14467
rect 15945 14433 15979 14467
rect 15979 14433 15988 14467
rect 15936 14424 15988 14433
rect 17132 14467 17184 14476
rect 1400 14399 1452 14408
rect 1400 14365 1409 14399
rect 1409 14365 1443 14399
rect 1443 14365 1452 14399
rect 1400 14356 1452 14365
rect 4068 14399 4120 14408
rect 4068 14365 4077 14399
rect 4077 14365 4111 14399
rect 4111 14365 4120 14399
rect 4068 14356 4120 14365
rect 5632 14356 5684 14408
rect 6460 14399 6512 14408
rect 6460 14365 6469 14399
rect 6469 14365 6503 14399
rect 6503 14365 6512 14399
rect 6460 14356 6512 14365
rect 5080 14288 5132 14340
rect 9036 14356 9088 14408
rect 9772 14399 9824 14408
rect 9772 14365 9781 14399
rect 9781 14365 9815 14399
rect 9815 14365 9824 14399
rect 9772 14356 9824 14365
rect 12440 14356 12492 14408
rect 17132 14433 17141 14467
rect 17141 14433 17175 14467
rect 17175 14433 17184 14467
rect 17132 14424 17184 14433
rect 18144 14424 18196 14476
rect 18328 14467 18380 14476
rect 18328 14433 18337 14467
rect 18337 14433 18371 14467
rect 18371 14433 18380 14467
rect 18328 14424 18380 14433
rect 19432 14424 19484 14476
rect 22192 14467 22244 14476
rect 22192 14433 22201 14467
rect 22201 14433 22235 14467
rect 22235 14433 22244 14467
rect 22192 14424 22244 14433
rect 24400 14467 24452 14476
rect 24400 14433 24409 14467
rect 24409 14433 24443 14467
rect 24443 14433 24452 14467
rect 24400 14424 24452 14433
rect 26608 14467 26660 14476
rect 26608 14433 26617 14467
rect 26617 14433 26651 14467
rect 26651 14433 26660 14467
rect 26608 14424 26660 14433
rect 27712 14424 27764 14476
rect 28264 14424 28316 14476
rect 28540 14467 28592 14476
rect 11152 14288 11204 14340
rect 16212 14288 16264 14340
rect 16764 14288 16816 14340
rect 19156 14356 19208 14408
rect 23480 14356 23532 14408
rect 24124 14399 24176 14408
rect 24124 14365 24133 14399
rect 24133 14365 24167 14399
rect 24167 14365 24176 14399
rect 24124 14356 24176 14365
rect 26148 14356 26200 14408
rect 27620 14356 27672 14408
rect 28080 14356 28132 14408
rect 4712 14220 4764 14272
rect 6552 14220 6604 14272
rect 7748 14263 7800 14272
rect 7748 14229 7757 14263
rect 7757 14229 7791 14263
rect 7791 14229 7800 14263
rect 7748 14220 7800 14229
rect 8760 14220 8812 14272
rect 19156 14220 19208 14272
rect 19432 14263 19484 14272
rect 19432 14229 19441 14263
rect 19441 14229 19475 14263
rect 19475 14229 19484 14263
rect 19432 14220 19484 14229
rect 20168 14220 20220 14272
rect 24124 14220 24176 14272
rect 25044 14220 25096 14272
rect 26792 14263 26844 14272
rect 26792 14229 26801 14263
rect 26801 14229 26835 14263
rect 26835 14229 26844 14263
rect 26792 14220 26844 14229
rect 26884 14220 26936 14272
rect 28540 14433 28549 14467
rect 28549 14433 28583 14467
rect 28583 14433 28592 14467
rect 28540 14424 28592 14433
rect 29092 14467 29144 14476
rect 29092 14433 29101 14467
rect 29101 14433 29135 14467
rect 29135 14433 29144 14467
rect 29092 14424 29144 14433
rect 30012 14424 30064 14476
rect 34336 14560 34388 14612
rect 37740 14560 37792 14612
rect 31576 14492 31628 14544
rect 32128 14467 32180 14476
rect 30288 14356 30340 14408
rect 32128 14433 32137 14467
rect 32137 14433 32171 14467
rect 32171 14433 32180 14467
rect 32128 14424 32180 14433
rect 34612 14424 34664 14476
rect 35532 14424 35584 14476
rect 33324 14356 33376 14408
rect 33876 14399 33928 14408
rect 33876 14365 33885 14399
rect 33885 14365 33919 14399
rect 33919 14365 33928 14399
rect 33876 14356 33928 14365
rect 34060 14356 34112 14408
rect 35808 14424 35860 14476
rect 36544 14467 36596 14476
rect 36544 14433 36553 14467
rect 36553 14433 36587 14467
rect 36587 14433 36596 14467
rect 36544 14424 36596 14433
rect 37740 14467 37792 14476
rect 37740 14433 37749 14467
rect 37749 14433 37783 14467
rect 37783 14433 37792 14467
rect 37740 14424 37792 14433
rect 37832 14424 37884 14476
rect 38568 14399 38620 14408
rect 38568 14365 38577 14399
rect 38577 14365 38611 14399
rect 38611 14365 38620 14399
rect 38568 14356 38620 14365
rect 29368 14288 29420 14340
rect 31208 14288 31260 14340
rect 32772 14288 32824 14340
rect 35808 14331 35860 14340
rect 35808 14297 35817 14331
rect 35817 14297 35851 14331
rect 35851 14297 35860 14331
rect 35808 14288 35860 14297
rect 30104 14220 30156 14272
rect 32588 14220 32640 14272
rect 33232 14220 33284 14272
rect 4246 14118 4298 14170
rect 4310 14118 4362 14170
rect 4374 14118 4426 14170
rect 4438 14118 4490 14170
rect 34966 14118 35018 14170
rect 35030 14118 35082 14170
rect 35094 14118 35146 14170
rect 35158 14118 35210 14170
rect 9956 14016 10008 14068
rect 11244 14016 11296 14068
rect 12072 14059 12124 14068
rect 12072 14025 12081 14059
rect 12081 14025 12115 14059
rect 12115 14025 12124 14059
rect 12072 14016 12124 14025
rect 12164 14016 12216 14068
rect 24860 14016 24912 14068
rect 5540 13948 5592 14000
rect 2688 13855 2740 13864
rect 2688 13821 2689 13855
rect 2689 13821 2723 13855
rect 2723 13821 2740 13855
rect 2688 13812 2740 13821
rect 4896 13812 4948 13864
rect 6000 13855 6052 13864
rect 6000 13821 6009 13855
rect 6009 13821 6043 13855
rect 6043 13821 6052 13855
rect 6000 13812 6052 13821
rect 6460 13948 6512 14000
rect 6736 13880 6788 13932
rect 7288 13855 7340 13864
rect 7288 13821 7297 13855
rect 7297 13821 7331 13855
rect 7331 13821 7340 13855
rect 7288 13812 7340 13821
rect 7748 13880 7800 13932
rect 8208 13855 8260 13864
rect 8208 13821 8217 13855
rect 8217 13821 8251 13855
rect 8251 13821 8260 13855
rect 8208 13812 8260 13821
rect 8760 13855 8812 13864
rect 8760 13821 8769 13855
rect 8769 13821 8803 13855
rect 8803 13821 8812 13855
rect 8760 13812 8812 13821
rect 9220 13855 9272 13864
rect 9220 13821 9229 13855
rect 9229 13821 9263 13855
rect 9263 13821 9272 13855
rect 9220 13812 9272 13821
rect 9404 13880 9456 13932
rect 10416 13812 10468 13864
rect 12440 13812 12492 13864
rect 13268 13812 13320 13864
rect 13360 13855 13412 13864
rect 13360 13821 13369 13855
rect 13369 13821 13403 13855
rect 13403 13821 13412 13855
rect 13360 13812 13412 13821
rect 13728 13812 13780 13864
rect 13912 13855 13964 13864
rect 13912 13821 13921 13855
rect 13921 13821 13955 13855
rect 13955 13821 13964 13855
rect 13912 13812 13964 13821
rect 15568 13948 15620 14000
rect 16120 13948 16172 14000
rect 16580 13948 16632 14000
rect 12900 13744 12952 13796
rect 15200 13855 15252 13864
rect 15200 13821 15209 13855
rect 15209 13821 15243 13855
rect 15243 13821 15252 13855
rect 15200 13812 15252 13821
rect 18512 13880 18564 13932
rect 16764 13812 16816 13864
rect 18052 13855 18104 13864
rect 18052 13821 18061 13855
rect 18061 13821 18095 13855
rect 18095 13821 18104 13855
rect 18052 13812 18104 13821
rect 18420 13855 18472 13864
rect 18420 13821 18429 13855
rect 18429 13821 18463 13855
rect 18463 13821 18472 13855
rect 18420 13812 18472 13821
rect 23204 13948 23256 14000
rect 19156 13880 19208 13932
rect 21088 13923 21140 13932
rect 21088 13889 21097 13923
rect 21097 13889 21131 13923
rect 21131 13889 21140 13923
rect 21088 13880 21140 13889
rect 22192 13880 22244 13932
rect 22284 13880 22336 13932
rect 24308 13923 24360 13932
rect 24308 13889 24317 13923
rect 24317 13889 24351 13923
rect 24351 13889 24360 13923
rect 24308 13880 24360 13889
rect 26148 14016 26200 14068
rect 19984 13812 20036 13864
rect 22560 13855 22612 13864
rect 22560 13821 22569 13855
rect 22569 13821 22603 13855
rect 22603 13821 22612 13855
rect 22560 13812 22612 13821
rect 23664 13855 23716 13864
rect 23664 13821 23673 13855
rect 23673 13821 23707 13855
rect 23707 13821 23716 13855
rect 23664 13812 23716 13821
rect 24124 13855 24176 13864
rect 24124 13821 24133 13855
rect 24133 13821 24167 13855
rect 24167 13821 24176 13855
rect 24124 13812 24176 13821
rect 25044 13855 25096 13864
rect 25044 13821 25053 13855
rect 25053 13821 25087 13855
rect 25087 13821 25096 13855
rect 31484 14016 31536 14068
rect 33416 14016 33468 14068
rect 37740 14016 37792 14068
rect 27252 13948 27304 14000
rect 34704 13948 34756 14000
rect 25044 13812 25096 13821
rect 27620 13880 27672 13932
rect 28080 13923 28132 13932
rect 28080 13889 28089 13923
rect 28089 13889 28123 13923
rect 28123 13889 28132 13923
rect 28080 13880 28132 13889
rect 28540 13880 28592 13932
rect 30012 13923 30064 13932
rect 30012 13889 30021 13923
rect 30021 13889 30055 13923
rect 30055 13889 30064 13923
rect 30012 13880 30064 13889
rect 30840 13923 30892 13932
rect 30840 13889 30849 13923
rect 30849 13889 30883 13923
rect 30883 13889 30892 13923
rect 30840 13880 30892 13889
rect 34152 13923 34204 13932
rect 34152 13889 34161 13923
rect 34161 13889 34195 13923
rect 34195 13889 34204 13923
rect 34152 13880 34204 13889
rect 35532 13923 35584 13932
rect 35532 13889 35541 13923
rect 35541 13889 35575 13923
rect 35575 13889 35584 13923
rect 35532 13880 35584 13889
rect 35808 13923 35860 13932
rect 35808 13889 35817 13923
rect 35817 13889 35851 13923
rect 35851 13889 35860 13923
rect 35808 13880 35860 13889
rect 38568 13880 38620 13932
rect 26884 13812 26936 13864
rect 27160 13855 27212 13864
rect 27160 13821 27169 13855
rect 27169 13821 27203 13855
rect 27203 13821 27212 13855
rect 27160 13812 27212 13821
rect 27436 13812 27488 13864
rect 27896 13812 27948 13864
rect 28724 13812 28776 13864
rect 28908 13812 28960 13864
rect 29092 13812 29144 13864
rect 29368 13812 29420 13864
rect 31392 13855 31444 13864
rect 31392 13821 31401 13855
rect 31401 13821 31435 13855
rect 31435 13821 31444 13855
rect 31392 13812 31444 13821
rect 31760 13855 31812 13864
rect 31760 13821 31769 13855
rect 31769 13821 31803 13855
rect 31803 13821 31812 13855
rect 31760 13812 31812 13821
rect 32496 13855 32548 13864
rect 4068 13676 4120 13728
rect 4344 13676 4396 13728
rect 16948 13744 17000 13796
rect 27252 13744 27304 13796
rect 28540 13744 28592 13796
rect 15292 13676 15344 13728
rect 16672 13676 16724 13728
rect 28724 13676 28776 13728
rect 28908 13676 28960 13728
rect 31208 13787 31260 13796
rect 31208 13753 31217 13787
rect 31217 13753 31251 13787
rect 31251 13753 31260 13787
rect 31208 13744 31260 13753
rect 31668 13744 31720 13796
rect 32496 13821 32505 13855
rect 32505 13821 32539 13855
rect 32539 13821 32548 13855
rect 32496 13812 32548 13821
rect 33232 13855 33284 13864
rect 33232 13821 33241 13855
rect 33241 13821 33275 13855
rect 33275 13821 33284 13855
rect 33232 13812 33284 13821
rect 33324 13812 33376 13864
rect 34336 13812 34388 13864
rect 38108 13855 38160 13864
rect 38108 13821 38117 13855
rect 38117 13821 38151 13855
rect 38151 13821 38160 13855
rect 38108 13812 38160 13821
rect 38476 13855 38528 13864
rect 38476 13821 38485 13855
rect 38485 13821 38519 13855
rect 38519 13821 38528 13855
rect 38476 13812 38528 13821
rect 29552 13719 29604 13728
rect 29552 13685 29561 13719
rect 29561 13685 29595 13719
rect 29595 13685 29604 13719
rect 29552 13676 29604 13685
rect 36544 13676 36596 13728
rect 19606 13574 19658 13626
rect 19670 13574 19722 13626
rect 19734 13574 19786 13626
rect 19798 13574 19850 13626
rect 5632 13515 5684 13524
rect 5632 13481 5641 13515
rect 5641 13481 5675 13515
rect 5675 13481 5684 13515
rect 5632 13472 5684 13481
rect 7288 13472 7340 13524
rect 8116 13472 8168 13524
rect 4068 13379 4120 13388
rect 4068 13345 4077 13379
rect 4077 13345 4111 13379
rect 4111 13345 4120 13379
rect 4068 13336 4120 13345
rect 4344 13379 4396 13388
rect 4344 13345 4353 13379
rect 4353 13345 4387 13379
rect 4387 13345 4396 13379
rect 4344 13336 4396 13345
rect 7748 13404 7800 13456
rect 1400 13311 1452 13320
rect 1400 13277 1409 13311
rect 1409 13277 1443 13311
rect 1443 13277 1452 13311
rect 1400 13268 1452 13277
rect 1676 13311 1728 13320
rect 1676 13277 1685 13311
rect 1685 13277 1719 13311
rect 1719 13277 1728 13311
rect 1676 13268 1728 13277
rect 7104 13311 7156 13320
rect 7104 13277 7113 13311
rect 7113 13277 7147 13311
rect 7147 13277 7156 13311
rect 7104 13268 7156 13277
rect 7380 13268 7432 13320
rect 8300 13336 8352 13388
rect 9680 13472 9732 13524
rect 10416 13472 10468 13524
rect 16948 13472 17000 13524
rect 17224 13472 17276 13524
rect 20628 13472 20680 13524
rect 22192 13472 22244 13524
rect 10140 13379 10192 13388
rect 10140 13345 10149 13379
rect 10149 13345 10183 13379
rect 10183 13345 10192 13379
rect 10140 13336 10192 13345
rect 10784 13379 10836 13388
rect 10784 13345 10793 13379
rect 10793 13345 10827 13379
rect 10827 13345 10836 13379
rect 10784 13336 10836 13345
rect 11060 13336 11112 13388
rect 11980 13379 12032 13388
rect 11980 13345 11989 13379
rect 11989 13345 12023 13379
rect 12023 13345 12032 13379
rect 11980 13336 12032 13345
rect 8116 13268 8168 13320
rect 13728 13379 13780 13388
rect 13728 13345 13737 13379
rect 13737 13345 13771 13379
rect 13771 13345 13780 13379
rect 13728 13336 13780 13345
rect 15752 13379 15804 13388
rect 7288 13200 7340 13252
rect 3792 13132 3844 13184
rect 13820 13268 13872 13320
rect 13268 13200 13320 13252
rect 14004 13200 14056 13252
rect 15752 13345 15761 13379
rect 15761 13345 15795 13379
rect 15795 13345 15804 13379
rect 15752 13336 15804 13345
rect 16120 13379 16172 13388
rect 16120 13345 16129 13379
rect 16129 13345 16163 13379
rect 16163 13345 16172 13379
rect 16120 13336 16172 13345
rect 16764 13336 16816 13388
rect 15936 13268 15988 13320
rect 18512 13336 18564 13388
rect 18236 13268 18288 13320
rect 13544 13132 13596 13184
rect 15108 13132 15160 13184
rect 15752 13132 15804 13184
rect 17132 13132 17184 13184
rect 19340 13336 19392 13388
rect 19892 13379 19944 13388
rect 19892 13345 19901 13379
rect 19901 13345 19935 13379
rect 19935 13345 19944 13379
rect 19892 13336 19944 13345
rect 20352 13379 20404 13388
rect 20352 13345 20361 13379
rect 20361 13345 20395 13379
rect 20395 13345 20404 13379
rect 20352 13336 20404 13345
rect 20444 13336 20496 13388
rect 20628 13336 20680 13388
rect 21180 13336 21232 13388
rect 21456 13379 21508 13388
rect 21456 13345 21465 13379
rect 21465 13345 21499 13379
rect 21499 13345 21508 13379
rect 21456 13336 21508 13345
rect 22652 13268 22704 13320
rect 23940 13404 23992 13456
rect 26424 13472 26476 13524
rect 29368 13515 29420 13524
rect 29368 13481 29377 13515
rect 29377 13481 29411 13515
rect 29411 13481 29420 13515
rect 29368 13472 29420 13481
rect 32312 13515 32364 13524
rect 26976 13404 27028 13456
rect 27344 13404 27396 13456
rect 19156 13200 19208 13252
rect 22284 13200 22336 13252
rect 21916 13132 21968 13184
rect 23572 13336 23624 13388
rect 24216 13268 24268 13320
rect 23664 13200 23716 13252
rect 27528 13336 27580 13388
rect 28080 13379 28132 13388
rect 28080 13345 28089 13379
rect 28089 13345 28123 13379
rect 28123 13345 28132 13379
rect 28080 13336 28132 13345
rect 29552 13404 29604 13456
rect 29000 13336 29052 13388
rect 30288 13336 30340 13388
rect 30840 13379 30892 13388
rect 30840 13345 30849 13379
rect 30849 13345 30883 13379
rect 30883 13345 30892 13379
rect 30840 13336 30892 13345
rect 31208 13336 31260 13388
rect 32312 13481 32321 13515
rect 32321 13481 32355 13515
rect 32355 13481 32364 13515
rect 32312 13472 32364 13481
rect 33876 13472 33928 13524
rect 33968 13472 34020 13524
rect 34060 13404 34112 13456
rect 33692 13379 33744 13388
rect 33692 13345 33701 13379
rect 33701 13345 33735 13379
rect 33735 13345 33744 13379
rect 33692 13336 33744 13345
rect 34152 13379 34204 13388
rect 34152 13345 34161 13379
rect 34161 13345 34195 13379
rect 34195 13345 34204 13379
rect 34152 13336 34204 13345
rect 37832 13404 37884 13456
rect 36084 13379 36136 13388
rect 36084 13345 36093 13379
rect 36093 13345 36127 13379
rect 36127 13345 36136 13379
rect 36084 13336 36136 13345
rect 36544 13379 36596 13388
rect 36544 13345 36553 13379
rect 36553 13345 36587 13379
rect 36587 13345 36596 13379
rect 36544 13336 36596 13345
rect 36728 13379 36780 13388
rect 36728 13345 36737 13379
rect 36737 13345 36771 13379
rect 36771 13345 36780 13379
rect 36728 13336 36780 13345
rect 37740 13379 37792 13388
rect 37740 13345 37749 13379
rect 37749 13345 37783 13379
rect 37783 13345 37792 13379
rect 37740 13336 37792 13345
rect 38200 13336 38252 13388
rect 27712 13268 27764 13320
rect 28908 13268 28960 13320
rect 30656 13311 30708 13320
rect 30656 13277 30665 13311
rect 30665 13277 30699 13311
rect 30699 13277 30708 13311
rect 30656 13268 30708 13277
rect 31392 13268 31444 13320
rect 32036 13268 32088 13320
rect 32312 13268 32364 13320
rect 38568 13311 38620 13320
rect 38568 13277 38577 13311
rect 38577 13277 38611 13311
rect 38611 13277 38620 13311
rect 38568 13268 38620 13277
rect 29736 13200 29788 13252
rect 31300 13243 31352 13252
rect 31300 13209 31309 13243
rect 31309 13209 31343 13243
rect 31343 13209 31352 13243
rect 31300 13200 31352 13209
rect 37740 13200 37792 13252
rect 35808 13132 35860 13184
rect 4246 13030 4298 13082
rect 4310 13030 4362 13082
rect 4374 13030 4426 13082
rect 4438 13030 4490 13082
rect 34966 13030 35018 13082
rect 35030 13030 35082 13082
rect 35094 13030 35146 13082
rect 35158 13030 35210 13082
rect 1676 12928 1728 12980
rect 4896 12971 4948 12980
rect 4896 12937 4905 12971
rect 4905 12937 4939 12971
rect 4939 12937 4948 12971
rect 4896 12928 4948 12937
rect 6184 12971 6236 12980
rect 6184 12937 6193 12971
rect 6193 12937 6227 12971
rect 6227 12937 6236 12971
rect 6184 12928 6236 12937
rect 16764 12928 16816 12980
rect 11060 12860 11112 12912
rect 13728 12860 13780 12912
rect 1400 12835 1452 12844
rect 1400 12801 1409 12835
rect 1409 12801 1443 12835
rect 1443 12801 1452 12835
rect 1400 12792 1452 12801
rect 1860 12792 1912 12844
rect 3792 12835 3844 12844
rect 3240 12724 3292 12776
rect 3792 12801 3801 12835
rect 3801 12801 3835 12835
rect 3835 12801 3844 12835
rect 3792 12792 3844 12801
rect 6920 12792 6972 12844
rect 7288 12835 7340 12844
rect 7288 12801 7297 12835
rect 7297 12801 7331 12835
rect 7331 12801 7340 12835
rect 7288 12792 7340 12801
rect 9864 12792 9916 12844
rect 13820 12792 13872 12844
rect 4068 12724 4120 12776
rect 9128 12767 9180 12776
rect 9128 12733 9137 12767
rect 9137 12733 9171 12767
rect 9171 12733 9180 12767
rect 9128 12724 9180 12733
rect 10692 12767 10744 12776
rect 8024 12656 8076 12708
rect 8484 12588 8536 12640
rect 10692 12733 10701 12767
rect 10701 12733 10735 12767
rect 10735 12733 10744 12767
rect 10692 12724 10744 12733
rect 10876 12767 10928 12776
rect 10876 12733 10885 12767
rect 10885 12733 10919 12767
rect 10919 12733 10928 12767
rect 10876 12724 10928 12733
rect 11796 12724 11848 12776
rect 12440 12588 12492 12640
rect 13728 12724 13780 12776
rect 14004 12724 14056 12776
rect 14188 12724 14240 12776
rect 15108 12767 15160 12776
rect 15108 12733 15117 12767
rect 15117 12733 15151 12767
rect 15151 12733 15160 12767
rect 15108 12724 15160 12733
rect 13268 12656 13320 12708
rect 13360 12588 13412 12640
rect 14004 12588 14056 12640
rect 14280 12588 14332 12640
rect 16580 12792 16632 12844
rect 15844 12724 15896 12776
rect 19248 12860 19300 12912
rect 18144 12792 18196 12844
rect 19156 12835 19208 12844
rect 19156 12801 19165 12835
rect 19165 12801 19199 12835
rect 19199 12801 19208 12835
rect 19156 12792 19208 12801
rect 20996 12928 21048 12980
rect 22284 12928 22336 12980
rect 22468 12928 22520 12980
rect 22836 12928 22888 12980
rect 20904 12860 20956 12912
rect 22652 12903 22704 12912
rect 22652 12869 22661 12903
rect 22661 12869 22695 12903
rect 22695 12869 22704 12903
rect 22652 12860 22704 12869
rect 18052 12767 18104 12776
rect 18052 12733 18061 12767
rect 18061 12733 18095 12767
rect 18095 12733 18104 12767
rect 18052 12724 18104 12733
rect 18420 12724 18472 12776
rect 17132 12656 17184 12708
rect 22100 12792 22152 12844
rect 19984 12767 20036 12776
rect 19984 12733 19993 12767
rect 19993 12733 20027 12767
rect 20027 12733 20036 12767
rect 19984 12724 20036 12733
rect 20076 12724 20128 12776
rect 20352 12724 20404 12776
rect 20536 12767 20588 12776
rect 20536 12733 20545 12767
rect 20545 12733 20579 12767
rect 20579 12733 20588 12767
rect 20536 12724 20588 12733
rect 20904 12767 20956 12776
rect 20904 12733 20913 12767
rect 20913 12733 20947 12767
rect 20947 12733 20956 12767
rect 20904 12724 20956 12733
rect 21916 12724 21968 12776
rect 22652 12767 22704 12776
rect 22652 12733 22661 12767
rect 22661 12733 22695 12767
rect 22695 12733 22704 12767
rect 22652 12724 22704 12733
rect 25780 12767 25832 12776
rect 25780 12733 25789 12767
rect 25789 12733 25823 12767
rect 25823 12733 25832 12767
rect 25780 12724 25832 12733
rect 28356 12860 28408 12912
rect 27344 12792 27396 12844
rect 27528 12792 27580 12844
rect 29828 12792 29880 12844
rect 30840 12835 30892 12844
rect 30840 12801 30849 12835
rect 30849 12801 30883 12835
rect 30883 12801 30892 12835
rect 30840 12792 30892 12801
rect 32036 12928 32088 12980
rect 32496 12928 32548 12980
rect 38200 12928 38252 12980
rect 31208 12860 31260 12912
rect 31392 12792 31444 12844
rect 18788 12588 18840 12640
rect 19340 12588 19392 12640
rect 27344 12656 27396 12708
rect 27712 12656 27764 12708
rect 28356 12699 28408 12708
rect 28356 12665 28365 12699
rect 28365 12665 28399 12699
rect 28399 12665 28408 12699
rect 28356 12656 28408 12665
rect 29092 12656 29144 12708
rect 30104 12656 30156 12708
rect 31760 12724 31812 12776
rect 32496 12724 32548 12776
rect 32680 12835 32732 12844
rect 32680 12801 32689 12835
rect 32689 12801 32723 12835
rect 32723 12801 32732 12835
rect 32680 12792 32732 12801
rect 33232 12767 33284 12776
rect 33232 12733 33241 12767
rect 33241 12733 33275 12767
rect 33275 12733 33284 12767
rect 33232 12724 33284 12733
rect 37740 12835 37792 12844
rect 37740 12801 37749 12835
rect 37749 12801 37783 12835
rect 37783 12801 37792 12835
rect 37740 12792 37792 12801
rect 39120 12835 39172 12844
rect 39120 12801 39129 12835
rect 39129 12801 39163 12835
rect 39163 12801 39172 12835
rect 39120 12792 39172 12801
rect 34060 12767 34112 12776
rect 34060 12733 34069 12767
rect 34069 12733 34103 12767
rect 34103 12733 34112 12767
rect 34060 12724 34112 12733
rect 31852 12656 31904 12708
rect 35256 12724 35308 12776
rect 36084 12767 36136 12776
rect 36084 12733 36093 12767
rect 36093 12733 36127 12767
rect 36127 12733 36136 12767
rect 36084 12724 36136 12733
rect 34244 12656 34296 12708
rect 36176 12656 36228 12708
rect 36544 12724 36596 12776
rect 37188 12724 37240 12776
rect 20628 12588 20680 12640
rect 23572 12588 23624 12640
rect 29552 12588 29604 12640
rect 31668 12588 31720 12640
rect 19606 12486 19658 12538
rect 19670 12486 19722 12538
rect 19734 12486 19786 12538
rect 19798 12486 19850 12538
rect 3240 12427 3292 12436
rect 3240 12393 3249 12427
rect 3249 12393 3283 12427
rect 3283 12393 3292 12427
rect 3240 12384 3292 12393
rect 10048 12384 10100 12436
rect 11980 12384 12032 12436
rect 1860 12291 1912 12300
rect 1860 12257 1869 12291
rect 1869 12257 1903 12291
rect 1903 12257 1912 12291
rect 1860 12248 1912 12257
rect 4712 12248 4764 12300
rect 5540 12291 5592 12300
rect 5540 12257 5549 12291
rect 5549 12257 5583 12291
rect 5583 12257 5592 12291
rect 5540 12248 5592 12257
rect 6184 12316 6236 12368
rect 6736 12316 6788 12368
rect 6276 12291 6328 12300
rect 6276 12257 6285 12291
rect 6285 12257 6319 12291
rect 6319 12257 6328 12291
rect 6276 12248 6328 12257
rect 7012 12316 7064 12368
rect 8208 12316 8260 12368
rect 7196 12248 7248 12300
rect 7840 12248 7892 12300
rect 8024 12291 8076 12300
rect 8024 12257 8033 12291
rect 8033 12257 8067 12291
rect 8067 12257 8076 12291
rect 8024 12248 8076 12257
rect 11152 12316 11204 12368
rect 8760 12291 8812 12300
rect 8760 12257 8769 12291
rect 8769 12257 8803 12291
rect 8803 12257 8812 12291
rect 8760 12248 8812 12257
rect 2136 12223 2188 12232
rect 2136 12189 2145 12223
rect 2145 12189 2179 12223
rect 2179 12189 2188 12223
rect 2136 12180 2188 12189
rect 7104 12180 7156 12232
rect 8300 12223 8352 12232
rect 8300 12189 8309 12223
rect 8309 12189 8343 12223
rect 8343 12189 8352 12223
rect 8300 12180 8352 12189
rect 10416 12248 10468 12300
rect 10692 12291 10744 12300
rect 10692 12257 10701 12291
rect 10701 12257 10735 12291
rect 10735 12257 10744 12291
rect 10692 12248 10744 12257
rect 11520 12291 11572 12300
rect 11520 12257 11529 12291
rect 11529 12257 11563 12291
rect 11563 12257 11572 12291
rect 11520 12248 11572 12257
rect 10140 12223 10192 12232
rect 10140 12189 10149 12223
rect 10149 12189 10183 12223
rect 10183 12189 10192 12223
rect 10140 12180 10192 12189
rect 11888 12248 11940 12300
rect 13636 12384 13688 12436
rect 17132 12384 17184 12436
rect 18880 12384 18932 12436
rect 13912 12316 13964 12368
rect 14372 12316 14424 12368
rect 12348 12180 12400 12232
rect 12532 12223 12584 12232
rect 12532 12189 12541 12223
rect 12541 12189 12575 12223
rect 12575 12189 12584 12223
rect 12532 12180 12584 12189
rect 14280 12248 14332 12300
rect 14556 12248 14608 12300
rect 18052 12316 18104 12368
rect 18236 12316 18288 12368
rect 19524 12316 19576 12368
rect 20260 12316 20312 12368
rect 17408 12291 17460 12300
rect 17408 12257 17417 12291
rect 17417 12257 17451 12291
rect 17451 12257 17460 12291
rect 17408 12248 17460 12257
rect 17960 12248 18012 12300
rect 19064 12291 19116 12300
rect 19064 12257 19073 12291
rect 19073 12257 19107 12291
rect 19107 12257 19116 12291
rect 19064 12248 19116 12257
rect 19432 12291 19484 12300
rect 19432 12257 19441 12291
rect 19441 12257 19475 12291
rect 19475 12257 19484 12291
rect 19432 12248 19484 12257
rect 20076 12291 20128 12300
rect 20076 12257 20085 12291
rect 20085 12257 20119 12291
rect 20119 12257 20128 12291
rect 20076 12248 20128 12257
rect 11520 12112 11572 12164
rect 17224 12180 17276 12232
rect 18236 12180 18288 12232
rect 19248 12180 19300 12232
rect 19892 12180 19944 12232
rect 20168 12180 20220 12232
rect 21088 12248 21140 12300
rect 23020 12384 23072 12436
rect 26792 12384 26844 12436
rect 27528 12384 27580 12436
rect 27712 12384 27764 12436
rect 28080 12384 28132 12436
rect 22836 12248 22888 12300
rect 23756 12316 23808 12368
rect 25780 12359 25832 12368
rect 25780 12325 25789 12359
rect 25789 12325 25823 12359
rect 25823 12325 25832 12359
rect 25780 12316 25832 12325
rect 28356 12316 28408 12368
rect 29092 12384 29144 12436
rect 29828 12384 29880 12436
rect 30748 12384 30800 12436
rect 32312 12384 32364 12436
rect 27620 12291 27672 12300
rect 27620 12257 27629 12291
rect 27629 12257 27663 12291
rect 27663 12257 27672 12291
rect 27620 12248 27672 12257
rect 28264 12291 28316 12300
rect 28264 12257 28273 12291
rect 28273 12257 28307 12291
rect 28307 12257 28316 12291
rect 28264 12248 28316 12257
rect 29552 12248 29604 12300
rect 30288 12291 30340 12300
rect 30288 12257 30297 12291
rect 30297 12257 30331 12291
rect 30331 12257 30340 12291
rect 30288 12248 30340 12257
rect 31392 12248 31444 12300
rect 32128 12291 32180 12300
rect 32128 12257 32137 12291
rect 32137 12257 32171 12291
rect 32171 12257 32180 12291
rect 32128 12248 32180 12257
rect 24124 12223 24176 12232
rect 2780 12044 2832 12096
rect 3700 12044 3752 12096
rect 13636 12044 13688 12096
rect 19248 12044 19300 12096
rect 20260 12087 20312 12096
rect 20260 12053 20269 12087
rect 20269 12053 20303 12087
rect 20303 12053 20312 12087
rect 20260 12044 20312 12053
rect 20904 12112 20956 12164
rect 24124 12189 24133 12223
rect 24133 12189 24167 12223
rect 24167 12189 24176 12223
rect 24124 12180 24176 12189
rect 24492 12180 24544 12232
rect 30564 12180 30616 12232
rect 32680 12248 32732 12300
rect 34060 12291 34112 12300
rect 34060 12257 34069 12291
rect 34069 12257 34103 12291
rect 34103 12257 34112 12291
rect 34060 12248 34112 12257
rect 22836 12112 22888 12164
rect 28080 12112 28132 12164
rect 28908 12112 28960 12164
rect 22560 12044 22612 12096
rect 27804 12044 27856 12096
rect 33232 12180 33284 12232
rect 34520 12223 34572 12232
rect 34520 12189 34529 12223
rect 34529 12189 34563 12223
rect 34563 12189 34572 12223
rect 34520 12180 34572 12189
rect 34796 12223 34848 12232
rect 34796 12189 34805 12223
rect 34805 12189 34839 12223
rect 34839 12189 34848 12223
rect 34796 12180 34848 12189
rect 36544 12248 36596 12300
rect 39120 12316 39172 12368
rect 38568 12291 38620 12300
rect 38568 12257 38577 12291
rect 38577 12257 38611 12291
rect 38611 12257 38620 12291
rect 38568 12248 38620 12257
rect 38476 12180 38528 12232
rect 31300 12087 31352 12096
rect 31300 12053 31309 12087
rect 31309 12053 31343 12087
rect 31343 12053 31352 12087
rect 31300 12044 31352 12053
rect 4246 11942 4298 11994
rect 4310 11942 4362 11994
rect 4374 11942 4426 11994
rect 4438 11942 4490 11994
rect 34966 11942 35018 11994
rect 35030 11942 35082 11994
rect 35094 11942 35146 11994
rect 35158 11942 35210 11994
rect 2136 11840 2188 11892
rect 8484 11840 8536 11892
rect 9680 11840 9732 11892
rect 12348 11840 12400 11892
rect 15384 11840 15436 11892
rect 18236 11883 18288 11892
rect 18236 11849 18245 11883
rect 18245 11849 18279 11883
rect 18279 11849 18288 11883
rect 18236 11840 18288 11849
rect 3516 11704 3568 11756
rect 7104 11747 7156 11756
rect 7104 11713 7113 11747
rect 7113 11713 7147 11747
rect 7147 11713 7156 11747
rect 7104 11704 7156 11713
rect 2688 11679 2740 11688
rect 2688 11645 2697 11679
rect 2697 11645 2731 11679
rect 2731 11645 2740 11679
rect 2688 11636 2740 11645
rect 4896 11636 4948 11688
rect 6920 11636 6972 11688
rect 16120 11772 16172 11824
rect 16580 11772 16632 11824
rect 19616 11840 19668 11892
rect 20628 11840 20680 11892
rect 19340 11772 19392 11824
rect 23664 11840 23716 11892
rect 22652 11772 22704 11824
rect 10784 11747 10836 11756
rect 10784 11713 10793 11747
rect 10793 11713 10827 11747
rect 10827 11713 10836 11747
rect 10784 11704 10836 11713
rect 13820 11747 13872 11756
rect 13820 11713 13829 11747
rect 13829 11713 13863 11747
rect 13863 11713 13872 11747
rect 13820 11704 13872 11713
rect 14096 11704 14148 11756
rect 9864 11679 9916 11688
rect 9864 11645 9873 11679
rect 9873 11645 9907 11679
rect 9907 11645 9916 11679
rect 9864 11636 9916 11645
rect 10140 11636 10192 11688
rect 11060 11636 11112 11688
rect 12440 11679 12492 11688
rect 12440 11645 12449 11679
rect 12449 11645 12483 11679
rect 12483 11645 12492 11679
rect 12440 11636 12492 11645
rect 12900 11568 12952 11620
rect 2780 11543 2832 11552
rect 2780 11509 2789 11543
rect 2789 11509 2823 11543
rect 2823 11509 2832 11543
rect 2780 11500 2832 11509
rect 8392 11500 8444 11552
rect 9128 11500 9180 11552
rect 11888 11500 11940 11552
rect 13912 11679 13964 11688
rect 13912 11645 13921 11679
rect 13921 11645 13955 11679
rect 13955 11645 13964 11679
rect 13912 11636 13964 11645
rect 15844 11636 15896 11688
rect 16304 11679 16356 11688
rect 16304 11645 16313 11679
rect 16313 11645 16347 11679
rect 16347 11645 16356 11679
rect 17224 11679 17276 11688
rect 16304 11636 16356 11645
rect 17224 11645 17233 11679
rect 17233 11645 17267 11679
rect 17267 11645 17276 11679
rect 17224 11636 17276 11645
rect 17960 11636 18012 11688
rect 19984 11704 20036 11756
rect 20260 11704 20312 11756
rect 26884 11840 26936 11892
rect 27620 11840 27672 11892
rect 27804 11840 27856 11892
rect 31852 11840 31904 11892
rect 33692 11840 33744 11892
rect 24308 11772 24360 11824
rect 19616 11679 19668 11688
rect 19616 11645 19625 11679
rect 19625 11645 19659 11679
rect 19659 11645 19668 11679
rect 19616 11636 19668 11645
rect 20628 11679 20680 11688
rect 17776 11568 17828 11620
rect 20628 11645 20637 11679
rect 20637 11645 20671 11679
rect 20671 11645 20680 11679
rect 20628 11636 20680 11645
rect 20996 11679 21048 11688
rect 20996 11645 21005 11679
rect 21005 11645 21039 11679
rect 21039 11645 21048 11679
rect 20996 11636 21048 11645
rect 22008 11636 22060 11688
rect 21548 11568 21600 11620
rect 22652 11636 22704 11688
rect 22928 11679 22980 11688
rect 22928 11645 22937 11679
rect 22937 11645 22971 11679
rect 22971 11645 22980 11679
rect 22928 11636 22980 11645
rect 23204 11636 23256 11688
rect 23848 11636 23900 11688
rect 29000 11704 29052 11756
rect 30472 11772 30524 11824
rect 31668 11772 31720 11824
rect 34796 11772 34848 11824
rect 36728 11772 36780 11824
rect 29460 11747 29512 11756
rect 29460 11713 29469 11747
rect 29469 11713 29503 11747
rect 29503 11713 29512 11747
rect 29460 11704 29512 11713
rect 27344 11679 27396 11688
rect 13912 11500 13964 11552
rect 19156 11500 19208 11552
rect 20628 11500 20680 11552
rect 22192 11568 22244 11620
rect 23940 11568 23992 11620
rect 22008 11500 22060 11552
rect 27344 11645 27353 11679
rect 27353 11645 27387 11679
rect 27387 11645 27396 11679
rect 27344 11636 27396 11645
rect 27712 11679 27764 11688
rect 27712 11645 27721 11679
rect 27721 11645 27755 11679
rect 27755 11645 27764 11679
rect 27712 11636 27764 11645
rect 27804 11636 27856 11688
rect 27988 11636 28040 11688
rect 29276 11636 29328 11688
rect 30656 11704 30708 11756
rect 30564 11679 30616 11688
rect 30564 11645 30573 11679
rect 30573 11645 30607 11679
rect 30607 11645 30616 11679
rect 34060 11704 34112 11756
rect 34244 11747 34296 11756
rect 34244 11713 34253 11747
rect 34253 11713 34287 11747
rect 34287 11713 34296 11747
rect 34244 11704 34296 11713
rect 35256 11704 35308 11756
rect 35716 11704 35768 11756
rect 30564 11636 30616 11645
rect 31484 11636 31536 11688
rect 32312 11679 32364 11688
rect 32312 11645 32321 11679
rect 32321 11645 32355 11679
rect 32355 11645 32364 11679
rect 32312 11636 32364 11645
rect 32772 11679 32824 11688
rect 32772 11645 32781 11679
rect 32781 11645 32815 11679
rect 32815 11645 32824 11679
rect 32772 11636 32824 11645
rect 33416 11679 33468 11688
rect 33416 11645 33425 11679
rect 33425 11645 33459 11679
rect 33459 11645 33468 11679
rect 33416 11636 33468 11645
rect 33692 11636 33744 11688
rect 34796 11636 34848 11688
rect 37188 11704 37240 11756
rect 37924 11704 37976 11756
rect 36176 11679 36228 11688
rect 25504 11500 25556 11552
rect 32404 11568 32456 11620
rect 36176 11645 36185 11679
rect 36185 11645 36219 11679
rect 36219 11645 36228 11679
rect 36176 11636 36228 11645
rect 30840 11500 30892 11552
rect 37832 11500 37884 11552
rect 19606 11398 19658 11450
rect 19670 11398 19722 11450
rect 19734 11398 19786 11450
rect 19798 11398 19850 11450
rect 7840 11339 7892 11348
rect 7840 11305 7849 11339
rect 7849 11305 7883 11339
rect 7883 11305 7892 11339
rect 7840 11296 7892 11305
rect 12716 11296 12768 11348
rect 13360 11296 13412 11348
rect 14372 11339 14424 11348
rect 14372 11305 14381 11339
rect 14381 11305 14415 11339
rect 14415 11305 14424 11339
rect 14372 11296 14424 11305
rect 1676 11160 1728 11212
rect 2780 11203 2832 11212
rect 2780 11169 2789 11203
rect 2789 11169 2823 11203
rect 2823 11169 2832 11203
rect 2964 11203 3016 11212
rect 2780 11160 2832 11169
rect 2964 11169 2973 11203
rect 2973 11169 3007 11203
rect 3007 11169 3016 11203
rect 2964 11160 3016 11169
rect 5540 11160 5592 11212
rect 5724 11160 5776 11212
rect 6368 11160 6420 11212
rect 7012 11228 7064 11280
rect 7196 11203 7248 11212
rect 7196 11169 7205 11203
rect 7205 11169 7239 11203
rect 7239 11169 7248 11203
rect 7196 11160 7248 11169
rect 6000 11092 6052 11144
rect 8392 11203 8444 11212
rect 2596 11024 2648 11076
rect 5540 11067 5592 11076
rect 5540 11033 5549 11067
rect 5549 11033 5583 11067
rect 5583 11033 5592 11067
rect 5540 11024 5592 11033
rect 8392 11169 8401 11203
rect 8401 11169 8435 11203
rect 8435 11169 8444 11203
rect 8392 11160 8444 11169
rect 8484 11160 8536 11212
rect 9680 11203 9732 11212
rect 9680 11169 9689 11203
rect 9689 11169 9723 11203
rect 9723 11169 9732 11203
rect 9680 11160 9732 11169
rect 11244 11203 11296 11212
rect 11244 11169 11253 11203
rect 11253 11169 11287 11203
rect 11287 11169 11296 11203
rect 11244 11160 11296 11169
rect 12072 11228 12124 11280
rect 16304 11296 16356 11348
rect 18236 11296 18288 11348
rect 19064 11296 19116 11348
rect 20076 11296 20128 11348
rect 12348 11203 12400 11212
rect 12348 11169 12357 11203
rect 12357 11169 12391 11203
rect 12391 11169 12400 11203
rect 12348 11160 12400 11169
rect 18328 11228 18380 11280
rect 21456 11296 21508 11348
rect 21548 11296 21600 11348
rect 25136 11296 25188 11348
rect 12532 11160 12584 11212
rect 13544 11203 13596 11212
rect 13544 11169 13553 11203
rect 13553 11169 13587 11203
rect 13587 11169 13596 11203
rect 13544 11160 13596 11169
rect 14188 11203 14240 11212
rect 14188 11169 14197 11203
rect 14197 11169 14231 11203
rect 14231 11169 14240 11203
rect 14188 11160 14240 11169
rect 15108 11160 15160 11212
rect 17960 11203 18012 11212
rect 17960 11169 17969 11203
rect 17969 11169 18003 11203
rect 18003 11169 18012 11203
rect 17960 11160 18012 11169
rect 18788 11160 18840 11212
rect 19064 11203 19116 11212
rect 19064 11169 19073 11203
rect 19073 11169 19107 11203
rect 19107 11169 19116 11203
rect 19064 11160 19116 11169
rect 19800 11160 19852 11212
rect 20076 11203 20128 11212
rect 20076 11169 20085 11203
rect 20085 11169 20119 11203
rect 20119 11169 20128 11203
rect 20076 11160 20128 11169
rect 20996 11203 21048 11212
rect 10876 11092 10928 11144
rect 10140 11024 10192 11076
rect 11428 11067 11480 11076
rect 11428 11033 11437 11067
rect 11437 11033 11471 11067
rect 11471 11033 11480 11067
rect 11428 11024 11480 11033
rect 13636 11092 13688 11144
rect 16212 11092 16264 11144
rect 11980 11024 12032 11076
rect 17776 11067 17828 11076
rect 17776 11033 17785 11067
rect 17785 11033 17819 11067
rect 17819 11033 17828 11067
rect 17776 11024 17828 11033
rect 19984 11024 20036 11076
rect 20996 11169 21005 11203
rect 21005 11169 21039 11203
rect 21039 11169 21048 11203
rect 20996 11160 21048 11169
rect 21916 11092 21968 11144
rect 22192 11160 22244 11212
rect 23204 11228 23256 11280
rect 27988 11296 28040 11348
rect 30564 11296 30616 11348
rect 32312 11296 32364 11348
rect 33600 11296 33652 11348
rect 23020 11160 23072 11212
rect 23848 11160 23900 11212
rect 25136 11203 25188 11212
rect 25136 11169 25145 11203
rect 25145 11169 25179 11203
rect 25179 11169 25188 11203
rect 25136 11160 25188 11169
rect 25688 11160 25740 11212
rect 23296 11135 23348 11144
rect 23296 11101 23305 11135
rect 23305 11101 23339 11135
rect 23339 11101 23348 11135
rect 23296 11092 23348 11101
rect 26424 11160 26476 11212
rect 26608 11160 26660 11212
rect 27712 11228 27764 11280
rect 27344 11160 27396 11212
rect 28264 11092 28316 11144
rect 29276 11203 29328 11212
rect 29276 11169 29285 11203
rect 29285 11169 29319 11203
rect 29319 11169 29328 11203
rect 29276 11160 29328 11169
rect 29828 11160 29880 11212
rect 30564 11203 30616 11212
rect 30564 11169 30573 11203
rect 30573 11169 30607 11203
rect 30607 11169 30616 11203
rect 30564 11160 30616 11169
rect 30840 11160 30892 11212
rect 32956 11228 33008 11280
rect 35808 11296 35860 11348
rect 36084 11296 36136 11348
rect 38660 11296 38712 11348
rect 32128 11203 32180 11212
rect 32128 11169 32137 11203
rect 32137 11169 32171 11203
rect 32171 11169 32180 11203
rect 32128 11160 32180 11169
rect 32312 11160 32364 11212
rect 32588 11160 32640 11212
rect 33048 11203 33100 11212
rect 33048 11169 33057 11203
rect 33057 11169 33091 11203
rect 33091 11169 33100 11203
rect 33048 11160 33100 11169
rect 33692 11203 33744 11212
rect 33692 11169 33701 11203
rect 33701 11169 33735 11203
rect 33735 11169 33744 11203
rect 33692 11160 33744 11169
rect 33784 11160 33836 11212
rect 37832 11203 37884 11212
rect 37832 11169 37841 11203
rect 37841 11169 37875 11203
rect 37875 11169 37884 11203
rect 37832 11160 37884 11169
rect 37924 11160 37976 11212
rect 22560 11024 22612 11076
rect 26976 11024 27028 11076
rect 10508 10956 10560 11008
rect 18052 10956 18104 11008
rect 20720 10956 20772 11008
rect 21272 10956 21324 11008
rect 24492 10999 24544 11008
rect 24492 10965 24501 10999
rect 24501 10965 24535 10999
rect 24535 10965 24544 10999
rect 24492 10956 24544 10965
rect 29000 11024 29052 11076
rect 30288 11092 30340 11144
rect 31484 11092 31536 11144
rect 32772 11092 32824 11144
rect 30840 11024 30892 11076
rect 32588 11024 32640 11076
rect 34612 11092 34664 11144
rect 36176 11092 36228 11144
rect 33968 11067 34020 11076
rect 33968 11033 33977 11067
rect 33977 11033 34011 11067
rect 34011 11033 34020 11067
rect 33968 11024 34020 11033
rect 28908 10956 28960 11008
rect 29092 10956 29144 11008
rect 33140 10956 33192 11008
rect 34336 10956 34388 11008
rect 35808 10956 35860 11008
rect 4246 10854 4298 10906
rect 4310 10854 4362 10906
rect 4374 10854 4426 10906
rect 4438 10854 4490 10906
rect 34966 10854 35018 10906
rect 35030 10854 35082 10906
rect 35094 10854 35146 10906
rect 35158 10854 35210 10906
rect 2688 10752 2740 10804
rect 4896 10795 4948 10804
rect 4896 10761 4905 10795
rect 4905 10761 4939 10795
rect 4939 10761 4948 10795
rect 4896 10752 4948 10761
rect 6000 10795 6052 10804
rect 6000 10761 6009 10795
rect 6009 10761 6043 10795
rect 6043 10761 6052 10795
rect 6000 10752 6052 10761
rect 16764 10795 16816 10804
rect 4620 10616 4672 10668
rect 11520 10684 11572 10736
rect 16764 10761 16773 10795
rect 16773 10761 16807 10795
rect 16807 10761 16816 10795
rect 16764 10752 16816 10761
rect 17132 10752 17184 10804
rect 20812 10752 20864 10804
rect 13176 10616 13228 10668
rect 1400 10591 1452 10600
rect 1400 10557 1409 10591
rect 1409 10557 1443 10591
rect 1443 10557 1452 10591
rect 1400 10548 1452 10557
rect 1676 10591 1728 10600
rect 1676 10557 1685 10591
rect 1685 10557 1719 10591
rect 1719 10557 1728 10591
rect 1676 10548 1728 10557
rect 3516 10591 3568 10600
rect 3516 10557 3525 10591
rect 3525 10557 3559 10591
rect 3559 10557 3568 10591
rect 3516 10548 3568 10557
rect 3792 10591 3844 10600
rect 3792 10557 3801 10591
rect 3801 10557 3835 10591
rect 3835 10557 3844 10591
rect 3792 10548 3844 10557
rect 5908 10591 5960 10600
rect 5908 10557 5917 10591
rect 5917 10557 5951 10591
rect 5951 10557 5960 10591
rect 5908 10548 5960 10557
rect 7104 10591 7156 10600
rect 7104 10557 7113 10591
rect 7113 10557 7147 10591
rect 7147 10557 7156 10591
rect 7104 10548 7156 10557
rect 9312 10591 9364 10600
rect 9312 10557 9321 10591
rect 9321 10557 9355 10591
rect 9355 10557 9364 10591
rect 9312 10548 9364 10557
rect 9864 10591 9916 10600
rect 9864 10557 9873 10591
rect 9873 10557 9907 10591
rect 9907 10557 9916 10591
rect 9864 10548 9916 10557
rect 11244 10548 11296 10600
rect 11520 10591 11572 10600
rect 11520 10557 11529 10591
rect 11529 10557 11563 10591
rect 11563 10557 11572 10591
rect 11520 10548 11572 10557
rect 11704 10591 11756 10600
rect 11704 10557 11713 10591
rect 11713 10557 11747 10591
rect 11747 10557 11756 10591
rect 11704 10548 11756 10557
rect 11888 10548 11940 10600
rect 14004 10591 14056 10600
rect 8944 10480 8996 10532
rect 10600 10480 10652 10532
rect 14004 10557 14013 10591
rect 14013 10557 14047 10591
rect 14047 10557 14056 10591
rect 14004 10548 14056 10557
rect 15568 10616 15620 10668
rect 8852 10412 8904 10464
rect 15292 10548 15344 10600
rect 16028 10616 16080 10668
rect 17224 10684 17276 10736
rect 26240 10752 26292 10804
rect 26424 10752 26476 10804
rect 27160 10795 27212 10804
rect 27160 10761 27169 10795
rect 27169 10761 27203 10795
rect 27203 10761 27212 10795
rect 27160 10752 27212 10761
rect 31484 10752 31536 10804
rect 33324 10752 33376 10804
rect 34796 10752 34848 10804
rect 37924 10752 37976 10804
rect 24860 10684 24912 10736
rect 25044 10684 25096 10736
rect 25320 10684 25372 10736
rect 26148 10684 26200 10736
rect 17408 10616 17460 10668
rect 22008 10659 22060 10668
rect 16212 10548 16264 10600
rect 17316 10591 17368 10600
rect 17316 10557 17325 10591
rect 17325 10557 17359 10591
rect 17359 10557 17368 10591
rect 17316 10548 17368 10557
rect 17500 10548 17552 10600
rect 18972 10548 19024 10600
rect 22008 10625 22017 10659
rect 22017 10625 22051 10659
rect 22051 10625 22060 10659
rect 22008 10616 22060 10625
rect 24308 10616 24360 10668
rect 20812 10591 20864 10600
rect 15476 10412 15528 10464
rect 17132 10480 17184 10532
rect 17960 10480 18012 10532
rect 19156 10480 19208 10532
rect 20812 10557 20821 10591
rect 20821 10557 20855 10591
rect 20855 10557 20864 10591
rect 20812 10548 20864 10557
rect 20996 10591 21048 10600
rect 20996 10557 21005 10591
rect 21005 10557 21039 10591
rect 21039 10557 21048 10591
rect 20996 10548 21048 10557
rect 21916 10548 21968 10600
rect 22928 10591 22980 10600
rect 22928 10557 22937 10591
rect 22937 10557 22971 10591
rect 22971 10557 22980 10591
rect 23756 10591 23808 10600
rect 22928 10548 22980 10557
rect 23756 10557 23765 10591
rect 23765 10557 23799 10591
rect 23799 10557 23808 10591
rect 23756 10548 23808 10557
rect 24584 10548 24636 10600
rect 23204 10480 23256 10532
rect 23848 10480 23900 10532
rect 25044 10591 25096 10600
rect 25044 10557 25053 10591
rect 25053 10557 25087 10591
rect 25087 10557 25096 10591
rect 25044 10548 25096 10557
rect 27160 10616 27212 10668
rect 26608 10548 26660 10600
rect 26976 10591 27028 10600
rect 26976 10557 26985 10591
rect 26985 10557 27019 10591
rect 27019 10557 27028 10591
rect 26976 10548 27028 10557
rect 28540 10591 28592 10600
rect 25780 10480 25832 10532
rect 17224 10412 17276 10464
rect 18236 10455 18288 10464
rect 18236 10421 18245 10455
rect 18245 10421 18279 10455
rect 18279 10421 18288 10455
rect 18236 10412 18288 10421
rect 19340 10412 19392 10464
rect 20628 10455 20680 10464
rect 20628 10421 20637 10455
rect 20637 10421 20671 10455
rect 20671 10421 20680 10455
rect 20628 10412 20680 10421
rect 21088 10455 21140 10464
rect 21088 10421 21097 10455
rect 21097 10421 21131 10455
rect 21131 10421 21140 10455
rect 21088 10412 21140 10421
rect 23480 10412 23532 10464
rect 24400 10412 24452 10464
rect 24584 10412 24636 10464
rect 25964 10455 26016 10464
rect 25964 10421 25973 10455
rect 25973 10421 26007 10455
rect 26007 10421 26016 10455
rect 25964 10412 26016 10421
rect 27804 10480 27856 10532
rect 28540 10557 28549 10591
rect 28549 10557 28583 10591
rect 28583 10557 28592 10591
rect 28540 10548 28592 10557
rect 29828 10684 29880 10736
rect 35716 10684 35768 10736
rect 29368 10616 29420 10668
rect 30564 10616 30616 10668
rect 30472 10548 30524 10600
rect 31300 10616 31352 10668
rect 32772 10659 32824 10668
rect 29184 10480 29236 10532
rect 32220 10548 32272 10600
rect 32496 10591 32548 10600
rect 32496 10557 32505 10591
rect 32505 10557 32539 10591
rect 32539 10557 32548 10591
rect 32496 10548 32548 10557
rect 32772 10625 32781 10659
rect 32781 10625 32815 10659
rect 32815 10625 32824 10659
rect 32772 10616 32824 10625
rect 33232 10616 33284 10668
rect 36176 10659 36228 10668
rect 32680 10548 32732 10600
rect 32864 10548 32916 10600
rect 36176 10625 36185 10659
rect 36185 10625 36219 10659
rect 36219 10625 36228 10659
rect 36176 10616 36228 10625
rect 36544 10616 36596 10668
rect 37188 10616 37240 10668
rect 31576 10480 31628 10532
rect 33600 10412 33652 10464
rect 36452 10591 36504 10600
rect 36452 10557 36461 10591
rect 36461 10557 36495 10591
rect 36495 10557 36504 10591
rect 36452 10548 36504 10557
rect 19606 10310 19658 10362
rect 19670 10310 19722 10362
rect 19734 10310 19786 10362
rect 19798 10310 19850 10362
rect 1676 10208 1728 10260
rect 5908 10208 5960 10260
rect 7012 10208 7064 10260
rect 9772 10251 9824 10260
rect 6368 10140 6420 10192
rect 2872 10072 2924 10124
rect 3700 10072 3752 10124
rect 5540 10072 5592 10124
rect 5632 10072 5684 10124
rect 9772 10217 9781 10251
rect 9781 10217 9815 10251
rect 9815 10217 9824 10251
rect 9772 10208 9824 10217
rect 17224 10208 17276 10260
rect 22560 10208 22612 10260
rect 22928 10208 22980 10260
rect 25688 10251 25740 10260
rect 25688 10217 25697 10251
rect 25697 10217 25731 10251
rect 25731 10217 25740 10251
rect 25688 10208 25740 10217
rect 26976 10208 27028 10260
rect 29092 10208 29144 10260
rect 29460 10208 29512 10260
rect 33140 10251 33192 10260
rect 33140 10217 33149 10251
rect 33149 10217 33183 10251
rect 33183 10217 33192 10251
rect 33140 10208 33192 10217
rect 33324 10208 33376 10260
rect 9956 10140 10008 10192
rect 11520 10140 11572 10192
rect 14556 10183 14608 10192
rect 14556 10149 14565 10183
rect 14565 10149 14599 10183
rect 14599 10149 14608 10183
rect 14556 10140 14608 10149
rect 15568 10140 15620 10192
rect 8944 10115 8996 10124
rect 1400 10047 1452 10056
rect 1400 10013 1409 10047
rect 1409 10013 1443 10047
rect 1443 10013 1452 10047
rect 1400 10004 1452 10013
rect 4620 10004 4672 10056
rect 5356 10004 5408 10056
rect 7104 10047 7156 10056
rect 7104 10013 7113 10047
rect 7113 10013 7147 10047
rect 7147 10013 7156 10047
rect 7104 10004 7156 10013
rect 8944 10081 8953 10115
rect 8953 10081 8987 10115
rect 8987 10081 8996 10115
rect 8944 10072 8996 10081
rect 9680 10115 9732 10124
rect 9680 10081 9689 10115
rect 9689 10081 9723 10115
rect 9723 10081 9732 10115
rect 9680 10072 9732 10081
rect 10048 10072 10100 10124
rect 10876 10072 10928 10124
rect 12808 10072 12860 10124
rect 13176 10115 13228 10124
rect 13176 10081 13185 10115
rect 13185 10081 13219 10115
rect 13219 10081 13228 10115
rect 13176 10072 13228 10081
rect 14004 10072 14056 10124
rect 16488 10115 16540 10124
rect 11796 10047 11848 10056
rect 11796 10013 11805 10047
rect 11805 10013 11839 10047
rect 11839 10013 11848 10047
rect 11796 10004 11848 10013
rect 12624 10004 12676 10056
rect 12440 9936 12492 9988
rect 2964 9868 3016 9920
rect 3516 9868 3568 9920
rect 16488 10081 16497 10115
rect 16497 10081 16531 10115
rect 16531 10081 16540 10115
rect 16488 10072 16540 10081
rect 18696 10140 18748 10192
rect 18972 10183 19024 10192
rect 18972 10149 18981 10183
rect 18981 10149 19015 10183
rect 19015 10149 19024 10183
rect 18972 10140 19024 10149
rect 18236 10115 18288 10124
rect 16028 10004 16080 10056
rect 18236 10081 18245 10115
rect 18245 10081 18279 10115
rect 18279 10081 18288 10115
rect 18236 10072 18288 10081
rect 19432 10072 19484 10124
rect 19984 10115 20036 10124
rect 19984 10081 19993 10115
rect 19993 10081 20027 10115
rect 20027 10081 20036 10115
rect 19984 10072 20036 10081
rect 21456 10115 21508 10124
rect 21456 10081 21465 10115
rect 21465 10081 21499 10115
rect 21499 10081 21508 10115
rect 21456 10072 21508 10081
rect 24124 10140 24176 10192
rect 29000 10183 29052 10192
rect 29000 10149 29009 10183
rect 29009 10149 29043 10183
rect 29043 10149 29052 10183
rect 29000 10140 29052 10149
rect 29368 10183 29420 10192
rect 29368 10149 29377 10183
rect 29377 10149 29411 10183
rect 29411 10149 29420 10183
rect 29368 10140 29420 10149
rect 29828 10140 29880 10192
rect 23480 10072 23532 10124
rect 19892 10004 19944 10056
rect 20076 10047 20128 10056
rect 20076 10013 20085 10047
rect 20085 10013 20119 10047
rect 20119 10013 20128 10047
rect 20076 10004 20128 10013
rect 21272 10047 21324 10056
rect 21272 10013 21281 10047
rect 21281 10013 21315 10047
rect 21315 10013 21324 10047
rect 21272 10004 21324 10013
rect 24216 10004 24268 10056
rect 16120 9979 16172 9988
rect 16120 9945 16129 9979
rect 16129 9945 16163 9979
rect 16163 9945 16172 9979
rect 16120 9936 16172 9945
rect 17408 9936 17460 9988
rect 22192 9936 22244 9988
rect 24124 9936 24176 9988
rect 24492 10004 24544 10056
rect 27160 10047 27212 10056
rect 16764 9868 16816 9920
rect 17316 9868 17368 9920
rect 18328 9868 18380 9920
rect 20076 9868 20128 9920
rect 25688 9868 25740 9920
rect 27160 10013 27169 10047
rect 27169 10013 27203 10047
rect 27203 10013 27212 10047
rect 27160 10004 27212 10013
rect 29736 10004 29788 10056
rect 31024 10072 31076 10124
rect 31300 10072 31352 10124
rect 32220 10115 32272 10124
rect 32220 10081 32249 10115
rect 32249 10081 32272 10115
rect 32220 10072 32272 10081
rect 32956 10004 33008 10056
rect 28908 9936 28960 9988
rect 30380 9979 30432 9988
rect 30380 9945 30389 9979
rect 30389 9945 30423 9979
rect 30423 9945 30432 9979
rect 30380 9936 30432 9945
rect 30840 9936 30892 9988
rect 33416 10047 33468 10056
rect 33416 10013 33425 10047
rect 33425 10013 33459 10047
rect 33459 10013 33468 10047
rect 33968 10072 34020 10124
rect 34704 10072 34756 10124
rect 37188 10115 37240 10124
rect 37188 10081 37197 10115
rect 37197 10081 37231 10115
rect 37231 10081 37240 10115
rect 37188 10072 37240 10081
rect 37924 10115 37976 10124
rect 37924 10081 37933 10115
rect 37933 10081 37967 10115
rect 37967 10081 37976 10115
rect 37924 10072 37976 10081
rect 38108 10115 38160 10124
rect 38108 10081 38117 10115
rect 38117 10081 38151 10115
rect 38151 10081 38160 10115
rect 38108 10072 38160 10081
rect 38384 10115 38436 10124
rect 38384 10081 38393 10115
rect 38393 10081 38427 10115
rect 38427 10081 38436 10115
rect 38384 10072 38436 10081
rect 33416 10004 33468 10013
rect 37004 10004 37056 10056
rect 37464 9936 37516 9988
rect 28172 9868 28224 9920
rect 32220 9868 32272 9920
rect 32404 9911 32456 9920
rect 32404 9877 32413 9911
rect 32413 9877 32447 9911
rect 32447 9877 32456 9911
rect 32404 9868 32456 9877
rect 38292 9868 38344 9920
rect 4246 9766 4298 9818
rect 4310 9766 4362 9818
rect 4374 9766 4426 9818
rect 4438 9766 4490 9818
rect 34966 9766 35018 9818
rect 35030 9766 35082 9818
rect 35094 9766 35146 9818
rect 35158 9766 35210 9818
rect 3792 9664 3844 9716
rect 9312 9707 9364 9716
rect 9312 9673 9321 9707
rect 9321 9673 9355 9707
rect 9355 9673 9364 9707
rect 9312 9664 9364 9673
rect 2688 9528 2740 9580
rect 4068 9528 4120 9580
rect 8024 9596 8076 9648
rect 5632 9528 5684 9580
rect 12532 9596 12584 9648
rect 15292 9664 15344 9716
rect 19524 9664 19576 9716
rect 20168 9596 20220 9648
rect 2964 9460 3016 9512
rect 4620 9503 4672 9512
rect 4620 9469 4629 9503
rect 4629 9469 4663 9503
rect 4663 9469 4672 9503
rect 4620 9460 4672 9469
rect 4896 9503 4948 9512
rect 4896 9469 4905 9503
rect 4905 9469 4939 9503
rect 4939 9469 4948 9503
rect 4896 9460 4948 9469
rect 7380 9503 7432 9512
rect 7380 9469 7389 9503
rect 7389 9469 7423 9503
rect 7423 9469 7432 9503
rect 7380 9460 7432 9469
rect 7840 9460 7892 9512
rect 7196 9392 7248 9444
rect 11152 9528 11204 9580
rect 8576 9503 8628 9512
rect 8576 9469 8585 9503
rect 8585 9469 8619 9503
rect 8619 9469 8628 9503
rect 8576 9460 8628 9469
rect 9772 9460 9824 9512
rect 10140 9460 10192 9512
rect 9496 9392 9548 9444
rect 11060 9460 11112 9512
rect 11244 9460 11296 9512
rect 11428 9460 11480 9512
rect 11796 9528 11848 9580
rect 15108 9571 15160 9580
rect 12532 9460 12584 9512
rect 15108 9537 15117 9571
rect 15117 9537 15151 9571
rect 15151 9537 15160 9571
rect 15108 9528 15160 9537
rect 14372 9503 14424 9512
rect 14372 9469 14381 9503
rect 14381 9469 14415 9503
rect 14415 9469 14424 9503
rect 14372 9460 14424 9469
rect 14648 9503 14700 9512
rect 14648 9469 14657 9503
rect 14657 9469 14691 9503
rect 14691 9469 14700 9503
rect 14648 9460 14700 9469
rect 14740 9460 14792 9512
rect 18052 9528 18104 9580
rect 15568 9460 15620 9512
rect 16580 9503 16632 9512
rect 16580 9469 16589 9503
rect 16589 9469 16623 9503
rect 16623 9469 16632 9503
rect 16580 9460 16632 9469
rect 16672 9503 16724 9512
rect 16672 9469 16681 9503
rect 16681 9469 16715 9503
rect 16715 9469 16724 9503
rect 16672 9460 16724 9469
rect 17132 9460 17184 9512
rect 17868 9460 17920 9512
rect 18604 9503 18656 9512
rect 18604 9469 18613 9503
rect 18613 9469 18647 9503
rect 18647 9469 18656 9503
rect 18604 9460 18656 9469
rect 18972 9503 19024 9512
rect 18972 9469 18981 9503
rect 18981 9469 19015 9503
rect 19015 9469 19024 9503
rect 18972 9460 19024 9469
rect 21180 9528 21232 9580
rect 21272 9528 21324 9580
rect 21088 9503 21140 9512
rect 21088 9469 21097 9503
rect 21097 9469 21131 9503
rect 21131 9469 21140 9503
rect 21088 9460 21140 9469
rect 24584 9664 24636 9716
rect 29000 9664 29052 9716
rect 21640 9596 21692 9648
rect 23296 9528 23348 9580
rect 7748 9324 7800 9376
rect 8852 9324 8904 9376
rect 10140 9324 10192 9376
rect 15844 9324 15896 9376
rect 19064 9324 19116 9376
rect 21640 9392 21692 9444
rect 21824 9392 21876 9444
rect 22560 9460 22612 9512
rect 23664 9503 23716 9512
rect 23664 9469 23673 9503
rect 23673 9469 23707 9503
rect 23707 9469 23716 9503
rect 23664 9460 23716 9469
rect 23848 9503 23900 9512
rect 23848 9469 23857 9503
rect 23857 9469 23891 9503
rect 23891 9469 23900 9503
rect 23848 9460 23900 9469
rect 24216 9596 24268 9648
rect 26884 9639 26936 9648
rect 26884 9605 26893 9639
rect 26893 9605 26927 9639
rect 26927 9605 26936 9639
rect 26884 9596 26936 9605
rect 28448 9596 28500 9648
rect 28908 9596 28960 9648
rect 33416 9664 33468 9716
rect 30840 9639 30892 9648
rect 25688 9528 25740 9580
rect 25964 9528 26016 9580
rect 24308 9503 24360 9512
rect 24308 9469 24317 9503
rect 24317 9469 24351 9503
rect 24351 9469 24360 9503
rect 24308 9460 24360 9469
rect 24860 9460 24912 9512
rect 25320 9460 25372 9512
rect 27344 9460 27396 9512
rect 20260 9324 20312 9376
rect 20628 9324 20680 9376
rect 23204 9324 23256 9376
rect 23388 9324 23440 9376
rect 27896 9460 27948 9512
rect 29092 9528 29144 9580
rect 29828 9528 29880 9580
rect 30840 9605 30849 9639
rect 30849 9605 30883 9639
rect 30883 9605 30892 9639
rect 30840 9596 30892 9605
rect 32036 9596 32088 9648
rect 32680 9596 32732 9648
rect 30288 9460 30340 9512
rect 31116 9503 31168 9512
rect 31116 9469 31125 9503
rect 31125 9469 31159 9503
rect 31159 9469 31168 9503
rect 31116 9460 31168 9469
rect 31576 9460 31628 9512
rect 31852 9503 31904 9512
rect 31852 9469 31861 9503
rect 31861 9469 31895 9503
rect 31895 9469 31904 9503
rect 31852 9460 31904 9469
rect 32312 9528 32364 9580
rect 32772 9503 32824 9512
rect 32772 9469 32781 9503
rect 32781 9469 32815 9503
rect 32815 9469 32824 9503
rect 32772 9460 32824 9469
rect 33600 9460 33652 9512
rect 33784 9503 33836 9512
rect 33784 9469 33793 9503
rect 33793 9469 33827 9503
rect 33827 9469 33836 9503
rect 33784 9460 33836 9469
rect 38752 9596 38804 9648
rect 37004 9571 37056 9580
rect 37004 9537 37013 9571
rect 37013 9537 37047 9571
rect 37047 9537 37056 9571
rect 37004 9528 37056 9537
rect 36176 9503 36228 9512
rect 28540 9324 28592 9376
rect 31300 9367 31352 9376
rect 31300 9333 31309 9367
rect 31309 9333 31343 9367
rect 31343 9333 31352 9367
rect 31300 9324 31352 9333
rect 31392 9324 31444 9376
rect 36176 9469 36185 9503
rect 36185 9469 36219 9503
rect 36219 9469 36228 9503
rect 36176 9460 36228 9469
rect 38108 9528 38160 9580
rect 37464 9503 37516 9512
rect 37464 9469 37473 9503
rect 37473 9469 37507 9503
rect 37507 9469 37516 9503
rect 37740 9503 37792 9512
rect 37464 9460 37516 9469
rect 37740 9469 37749 9503
rect 37749 9469 37783 9503
rect 37783 9469 37792 9503
rect 37740 9460 37792 9469
rect 37280 9367 37332 9376
rect 37280 9333 37289 9367
rect 37289 9333 37323 9367
rect 37323 9333 37332 9367
rect 37280 9324 37332 9333
rect 37740 9324 37792 9376
rect 38568 9324 38620 9376
rect 19606 9222 19658 9274
rect 19670 9222 19722 9274
rect 19734 9222 19786 9274
rect 19798 9222 19850 9274
rect 2872 9163 2924 9172
rect 2872 9129 2881 9163
rect 2881 9129 2915 9163
rect 2915 9129 2924 9163
rect 2872 9120 2924 9129
rect 3056 9120 3108 9172
rect 2780 9052 2832 9104
rect 8484 9120 8536 9172
rect 8576 9120 8628 9172
rect 14556 9120 14608 9172
rect 18144 9120 18196 9172
rect 19432 9120 19484 9172
rect 22284 9120 22336 9172
rect 23112 9120 23164 9172
rect 23480 9120 23532 9172
rect 23848 9120 23900 9172
rect 1860 8959 1912 8968
rect 1860 8925 1869 8959
rect 1869 8925 1903 8959
rect 1903 8925 1912 8959
rect 1860 8916 1912 8925
rect 2596 8984 2648 9036
rect 3332 9027 3384 9036
rect 2964 8916 3016 8968
rect 3332 8993 3341 9027
rect 3341 8993 3375 9027
rect 3375 8993 3384 9027
rect 3332 8984 3384 8993
rect 4068 9027 4120 9036
rect 4068 8993 4077 9027
rect 4077 8993 4111 9027
rect 4111 8993 4120 9027
rect 4068 8984 4120 8993
rect 5172 8984 5224 9036
rect 5356 9027 5408 9036
rect 5356 8993 5365 9027
rect 5365 8993 5399 9027
rect 5399 8993 5408 9027
rect 5356 8984 5408 8993
rect 9864 9052 9916 9104
rect 10968 9052 11020 9104
rect 6368 9027 6420 9036
rect 6368 8993 6377 9027
rect 6377 8993 6411 9027
rect 6411 8993 6420 9027
rect 6368 8984 6420 8993
rect 6920 8984 6972 9036
rect 7196 9027 7248 9036
rect 7196 8993 7205 9027
rect 7205 8993 7239 9027
rect 7239 8993 7248 9027
rect 7196 8984 7248 8993
rect 7748 9027 7800 9036
rect 7748 8993 7757 9027
rect 7757 8993 7791 9027
rect 7791 8993 7800 9027
rect 7748 8984 7800 8993
rect 10324 9027 10376 9036
rect 4620 8959 4672 8968
rect 4620 8925 4629 8959
rect 4629 8925 4663 8959
rect 4663 8925 4672 8959
rect 4620 8916 4672 8925
rect 4896 8916 4948 8968
rect 1768 8848 1820 8900
rect 10324 8993 10333 9027
rect 10333 8993 10367 9027
rect 10367 8993 10376 9027
rect 10324 8984 10376 8993
rect 10416 9027 10468 9036
rect 10416 8993 10425 9027
rect 10425 8993 10459 9027
rect 10459 8993 10468 9027
rect 10416 8984 10468 8993
rect 11704 9052 11756 9104
rect 12164 9027 12216 9036
rect 9864 8916 9916 8968
rect 12164 8993 12173 9027
rect 12173 8993 12207 9027
rect 12207 8993 12216 9027
rect 12164 8984 12216 8993
rect 15844 9052 15896 9104
rect 17224 9052 17276 9104
rect 19892 9052 19944 9104
rect 12532 9027 12584 9036
rect 12532 8993 12541 9027
rect 12541 8993 12575 9027
rect 12575 8993 12584 9027
rect 12532 8984 12584 8993
rect 12624 9027 12676 9036
rect 12624 8993 12633 9027
rect 12633 8993 12667 9027
rect 12667 8993 12676 9027
rect 12624 8984 12676 8993
rect 11060 8916 11112 8968
rect 12072 8916 12124 8968
rect 13176 8984 13228 9036
rect 13360 9027 13412 9036
rect 13360 8993 13369 9027
rect 13369 8993 13403 9027
rect 13403 8993 13412 9027
rect 13360 8984 13412 8993
rect 13820 9027 13872 9036
rect 13820 8993 13829 9027
rect 13829 8993 13863 9027
rect 13863 8993 13872 9027
rect 13820 8984 13872 8993
rect 14280 9027 14332 9036
rect 14280 8993 14289 9027
rect 14289 8993 14323 9027
rect 14323 8993 14332 9027
rect 14280 8984 14332 8993
rect 16120 9027 16172 9036
rect 16120 8993 16129 9027
rect 16129 8993 16163 9027
rect 16163 8993 16172 9027
rect 16120 8984 16172 8993
rect 18604 9027 18656 9036
rect 15292 8916 15344 8968
rect 16304 8916 16356 8968
rect 18604 8993 18613 9027
rect 18613 8993 18647 9027
rect 18647 8993 18656 9027
rect 18604 8984 18656 8993
rect 19064 8984 19116 9036
rect 21916 9052 21968 9104
rect 26148 9120 26200 9172
rect 26608 9163 26660 9172
rect 26608 9129 26617 9163
rect 26617 9129 26651 9163
rect 26651 9129 26660 9163
rect 26608 9120 26660 9129
rect 29184 9120 29236 9172
rect 30288 9120 30340 9172
rect 37280 9120 37332 9172
rect 18880 8916 18932 8968
rect 8576 8780 8628 8832
rect 14096 8848 14148 8900
rect 15108 8848 15160 8900
rect 18696 8848 18748 8900
rect 19156 8848 19208 8900
rect 20260 8984 20312 9036
rect 20536 8984 20588 9036
rect 19708 8916 19760 8968
rect 21732 9027 21784 9036
rect 21732 8993 21741 9027
rect 21741 8993 21775 9027
rect 21775 8993 21784 9027
rect 21732 8984 21784 8993
rect 22192 8984 22244 9036
rect 23112 8984 23164 9036
rect 23848 8984 23900 9036
rect 24400 9027 24452 9036
rect 24400 8993 24409 9027
rect 24409 8993 24443 9027
rect 24443 8993 24452 9027
rect 24400 8984 24452 8993
rect 24676 8984 24728 9036
rect 25320 9052 25372 9104
rect 27160 9052 27212 9104
rect 27344 9052 27396 9104
rect 29092 9052 29144 9104
rect 26884 8984 26936 9036
rect 27804 9027 27856 9036
rect 27804 8993 27813 9027
rect 27813 8993 27847 9027
rect 27847 8993 27856 9027
rect 27804 8984 27856 8993
rect 28080 9027 28132 9036
rect 28080 8993 28089 9027
rect 28089 8993 28123 9027
rect 28123 8993 28132 9027
rect 28080 8984 28132 8993
rect 28448 8984 28500 9036
rect 28816 8984 28868 9036
rect 29000 8984 29052 9036
rect 30656 9052 30708 9104
rect 20444 8848 20496 8900
rect 25412 8916 25464 8968
rect 29368 8916 29420 8968
rect 29920 8959 29972 8968
rect 29920 8925 29929 8959
rect 29929 8925 29963 8959
rect 29963 8925 29972 8959
rect 29920 8916 29972 8925
rect 31116 8984 31168 9036
rect 37924 9052 37976 9104
rect 32864 8984 32916 9036
rect 33140 9027 33192 9036
rect 32036 8916 32088 8968
rect 21180 8848 21232 8900
rect 22744 8848 22796 8900
rect 13176 8823 13228 8832
rect 13176 8789 13185 8823
rect 13185 8789 13219 8823
rect 13219 8789 13228 8823
rect 13176 8780 13228 8789
rect 20260 8780 20312 8832
rect 24952 8848 25004 8900
rect 29460 8848 29512 8900
rect 29644 8848 29696 8900
rect 32588 8891 32640 8900
rect 32588 8857 32597 8891
rect 32597 8857 32631 8891
rect 32631 8857 32640 8891
rect 32588 8848 32640 8857
rect 31300 8780 31352 8832
rect 33140 8993 33149 9027
rect 33149 8993 33183 9027
rect 33183 8993 33192 9027
rect 33140 8984 33192 8993
rect 34336 9027 34388 9036
rect 34336 8993 34345 9027
rect 34345 8993 34379 9027
rect 34379 8993 34388 9027
rect 34336 8984 34388 8993
rect 37096 8984 37148 9036
rect 38292 9027 38344 9036
rect 34520 8916 34572 8968
rect 35808 8916 35860 8968
rect 36820 8916 36872 8968
rect 38292 8993 38301 9027
rect 38301 8993 38335 9027
rect 38335 8993 38344 9027
rect 38292 8984 38344 8993
rect 36452 8780 36504 8832
rect 4246 8678 4298 8730
rect 4310 8678 4362 8730
rect 4374 8678 4426 8730
rect 4438 8678 4490 8730
rect 34966 8678 35018 8730
rect 35030 8678 35082 8730
rect 35094 8678 35146 8730
rect 35158 8678 35210 8730
rect 3332 8508 3384 8560
rect 3240 8415 3292 8424
rect 3240 8381 3249 8415
rect 3249 8381 3283 8415
rect 3283 8381 3292 8415
rect 3240 8372 3292 8381
rect 3608 8415 3660 8424
rect 3608 8381 3617 8415
rect 3617 8381 3651 8415
rect 3651 8381 3660 8415
rect 3608 8372 3660 8381
rect 4068 8372 4120 8424
rect 7840 8483 7892 8492
rect 7840 8449 7849 8483
rect 7849 8449 7883 8483
rect 7883 8449 7892 8483
rect 7840 8440 7892 8449
rect 8392 8440 8444 8492
rect 8760 8440 8812 8492
rect 8576 8415 8628 8424
rect 3424 8304 3476 8356
rect 6460 8304 6512 8356
rect 8576 8381 8585 8415
rect 8585 8381 8619 8415
rect 8619 8381 8628 8415
rect 8576 8372 8628 8381
rect 9680 8372 9732 8424
rect 8024 8304 8076 8356
rect 11152 8576 11204 8628
rect 16212 8576 16264 8628
rect 21456 8576 21508 8628
rect 22652 8576 22704 8628
rect 36176 8576 36228 8628
rect 37924 8619 37976 8628
rect 37924 8585 37933 8619
rect 37933 8585 37967 8619
rect 37967 8585 37976 8619
rect 37924 8576 37976 8585
rect 10508 8508 10560 8560
rect 17224 8508 17276 8560
rect 9864 8440 9916 8492
rect 10784 8440 10836 8492
rect 10968 8440 11020 8492
rect 12164 8440 12216 8492
rect 13820 8483 13872 8492
rect 13820 8449 13829 8483
rect 13829 8449 13863 8483
rect 13863 8449 13872 8483
rect 13820 8440 13872 8449
rect 11336 8415 11388 8424
rect 11336 8381 11345 8415
rect 11345 8381 11379 8415
rect 11379 8381 11388 8415
rect 11336 8372 11388 8381
rect 12072 8372 12124 8424
rect 11796 8304 11848 8356
rect 12256 8304 12308 8356
rect 13544 8372 13596 8424
rect 13912 8372 13964 8424
rect 14372 8440 14424 8492
rect 14648 8415 14700 8424
rect 14648 8381 14657 8415
rect 14657 8381 14691 8415
rect 14691 8381 14700 8415
rect 14648 8372 14700 8381
rect 19432 8440 19484 8492
rect 19984 8483 20036 8492
rect 19984 8449 19993 8483
rect 19993 8449 20027 8483
rect 20027 8449 20036 8483
rect 19984 8440 20036 8449
rect 20168 8440 20220 8492
rect 15568 8415 15620 8424
rect 15568 8381 15577 8415
rect 15577 8381 15611 8415
rect 15611 8381 15620 8415
rect 15568 8372 15620 8381
rect 16028 8415 16080 8424
rect 16028 8381 16037 8415
rect 16037 8381 16071 8415
rect 16071 8381 16080 8415
rect 16028 8372 16080 8381
rect 16764 8415 16816 8424
rect 16764 8381 16773 8415
rect 16773 8381 16807 8415
rect 16807 8381 16816 8415
rect 16764 8372 16816 8381
rect 18236 8415 18288 8424
rect 18236 8381 18245 8415
rect 18245 8381 18279 8415
rect 18279 8381 18288 8415
rect 18236 8372 18288 8381
rect 18604 8415 18656 8424
rect 18604 8381 18613 8415
rect 18613 8381 18647 8415
rect 18647 8381 18656 8415
rect 18604 8372 18656 8381
rect 19064 8415 19116 8424
rect 19064 8381 19073 8415
rect 19073 8381 19107 8415
rect 19107 8381 19116 8415
rect 19064 8372 19116 8381
rect 7380 8236 7432 8288
rect 10048 8236 10100 8288
rect 15568 8236 15620 8288
rect 19340 8304 19392 8356
rect 21916 8440 21968 8492
rect 24032 8508 24084 8560
rect 24676 8508 24728 8560
rect 28632 8551 28684 8560
rect 28632 8517 28641 8551
rect 28641 8517 28675 8551
rect 28675 8517 28684 8551
rect 28632 8508 28684 8517
rect 22376 8483 22428 8492
rect 22376 8449 22385 8483
rect 22385 8449 22419 8483
rect 22419 8449 22428 8483
rect 22376 8440 22428 8449
rect 23664 8440 23716 8492
rect 24952 8483 25004 8492
rect 22008 8415 22060 8424
rect 22008 8381 22017 8415
rect 22017 8381 22051 8415
rect 22051 8381 22060 8415
rect 22008 8372 22060 8381
rect 22284 8415 22336 8424
rect 22284 8381 22293 8415
rect 22293 8381 22327 8415
rect 22327 8381 22336 8415
rect 22284 8372 22336 8381
rect 22560 8415 22612 8424
rect 22560 8381 22569 8415
rect 22569 8381 22603 8415
rect 22603 8381 22612 8415
rect 22560 8372 22612 8381
rect 23940 8372 23992 8424
rect 24952 8449 24961 8483
rect 24961 8449 24995 8483
rect 24995 8449 25004 8483
rect 24952 8440 25004 8449
rect 25596 8440 25648 8492
rect 28908 8440 28960 8492
rect 31392 8440 31444 8492
rect 36820 8483 36872 8492
rect 36820 8449 36829 8483
rect 36829 8449 36863 8483
rect 36863 8449 36872 8483
rect 36820 8440 36872 8449
rect 23388 8304 23440 8356
rect 27620 8372 27672 8424
rect 28816 8372 28868 8424
rect 29184 8372 29236 8424
rect 29552 8415 29604 8424
rect 29552 8381 29561 8415
rect 29561 8381 29595 8415
rect 29595 8381 29604 8415
rect 29552 8372 29604 8381
rect 31576 8415 31628 8424
rect 31576 8381 31585 8415
rect 31585 8381 31619 8415
rect 31619 8381 31628 8415
rect 31576 8372 31628 8381
rect 32312 8304 32364 8356
rect 20996 8236 21048 8288
rect 21088 8236 21140 8288
rect 22192 8236 22244 8288
rect 22836 8236 22888 8288
rect 28540 8236 28592 8288
rect 28724 8236 28776 8288
rect 28908 8236 28960 8288
rect 32588 8372 32640 8424
rect 35900 8415 35952 8424
rect 34336 8304 34388 8356
rect 35900 8381 35909 8415
rect 35909 8381 35943 8415
rect 35943 8381 35952 8415
rect 35900 8372 35952 8381
rect 36544 8415 36596 8424
rect 36544 8381 36553 8415
rect 36553 8381 36587 8415
rect 36587 8381 36596 8415
rect 36544 8372 36596 8381
rect 36636 8372 36688 8424
rect 38108 8372 38160 8424
rect 35992 8304 36044 8356
rect 33876 8279 33928 8288
rect 33876 8245 33885 8279
rect 33885 8245 33919 8279
rect 33919 8245 33928 8279
rect 33876 8236 33928 8245
rect 19606 8134 19658 8186
rect 19670 8134 19722 8186
rect 19734 8134 19786 8186
rect 19798 8134 19850 8186
rect 3240 8075 3292 8084
rect 3240 8041 3249 8075
rect 3249 8041 3283 8075
rect 3283 8041 3292 8075
rect 3240 8032 3292 8041
rect 6460 8075 6512 8084
rect 6460 8041 6469 8075
rect 6469 8041 6503 8075
rect 6503 8041 6512 8075
rect 6460 8032 6512 8041
rect 11336 8032 11388 8084
rect 2872 7896 2924 7948
rect 4620 7896 4672 7948
rect 4712 7896 4764 7948
rect 5632 7896 5684 7948
rect 8024 7939 8076 7948
rect 3056 7828 3108 7880
rect 3792 7828 3844 7880
rect 4068 7692 4120 7744
rect 8024 7905 8033 7939
rect 8033 7905 8067 7939
rect 8067 7905 8076 7939
rect 8024 7896 8076 7905
rect 8392 7939 8444 7948
rect 8392 7905 8401 7939
rect 8401 7905 8435 7939
rect 8435 7905 8444 7939
rect 8392 7896 8444 7905
rect 9312 7896 9364 7948
rect 9864 7939 9916 7948
rect 9864 7905 9873 7939
rect 9873 7905 9907 7939
rect 9907 7905 9916 7939
rect 9864 7896 9916 7905
rect 10048 7939 10100 7948
rect 10048 7905 10057 7939
rect 10057 7905 10091 7939
rect 10091 7905 10100 7939
rect 10048 7896 10100 7905
rect 10508 7939 10560 7948
rect 10508 7905 10517 7939
rect 10517 7905 10551 7939
rect 10551 7905 10560 7939
rect 10508 7896 10560 7905
rect 10692 7896 10744 7948
rect 11796 7939 11848 7948
rect 11796 7905 11805 7939
rect 11805 7905 11839 7939
rect 11839 7905 11848 7939
rect 11796 7896 11848 7905
rect 14556 8032 14608 8084
rect 12532 7964 12584 8016
rect 7656 7871 7708 7880
rect 7656 7837 7665 7871
rect 7665 7837 7699 7871
rect 7699 7837 7708 7871
rect 7656 7828 7708 7837
rect 7840 7692 7892 7744
rect 12532 7828 12584 7880
rect 13820 7896 13872 7948
rect 15476 7896 15528 7948
rect 16212 7939 16264 7948
rect 16212 7905 16221 7939
rect 16221 7905 16255 7939
rect 16255 7905 16264 7939
rect 16212 7896 16264 7905
rect 17684 8032 17736 8084
rect 22100 8032 22152 8084
rect 22560 8032 22612 8084
rect 23756 8032 23808 8084
rect 24032 8075 24084 8084
rect 24032 8041 24041 8075
rect 24041 8041 24075 8075
rect 24075 8041 24084 8075
rect 24032 8032 24084 8041
rect 27620 8032 27672 8084
rect 31024 8032 31076 8084
rect 16856 7964 16908 8016
rect 23480 7964 23532 8016
rect 17960 7896 18012 7948
rect 18144 7896 18196 7948
rect 18604 7939 18656 7948
rect 18604 7905 18613 7939
rect 18613 7905 18647 7939
rect 18647 7905 18656 7939
rect 18604 7896 18656 7905
rect 19248 7939 19300 7948
rect 19248 7905 19257 7939
rect 19257 7905 19291 7939
rect 19291 7905 19300 7939
rect 19248 7896 19300 7905
rect 21088 7896 21140 7948
rect 23112 7896 23164 7948
rect 23940 7939 23992 7948
rect 23940 7905 23949 7939
rect 23949 7905 23983 7939
rect 23983 7905 23992 7939
rect 23940 7896 23992 7905
rect 25320 7939 25372 7948
rect 25320 7905 25329 7939
rect 25329 7905 25363 7939
rect 25363 7905 25372 7939
rect 25320 7896 25372 7905
rect 25504 7939 25556 7948
rect 25504 7905 25513 7939
rect 25513 7905 25547 7939
rect 25547 7905 25556 7939
rect 25504 7896 25556 7905
rect 29552 7964 29604 8016
rect 29828 7964 29880 8016
rect 34520 8032 34572 8084
rect 29276 7896 29328 7948
rect 29920 7896 29972 7948
rect 30380 7896 30432 7948
rect 37096 7964 37148 8016
rect 38292 7964 38344 8016
rect 31116 7939 31168 7948
rect 31116 7905 31125 7939
rect 31125 7905 31159 7939
rect 31159 7905 31168 7939
rect 31116 7896 31168 7905
rect 32496 7896 32548 7948
rect 33876 7896 33928 7948
rect 9680 7760 9732 7812
rect 12440 7760 12492 7812
rect 12624 7760 12676 7812
rect 13820 7692 13872 7744
rect 14648 7692 14700 7744
rect 16028 7735 16080 7744
rect 16028 7701 16037 7735
rect 16037 7701 16071 7735
rect 16071 7701 16080 7735
rect 16028 7692 16080 7701
rect 20996 7828 21048 7880
rect 21824 7871 21876 7880
rect 21824 7837 21833 7871
rect 21833 7837 21867 7871
rect 21867 7837 21876 7871
rect 21824 7828 21876 7837
rect 22284 7828 22336 7880
rect 24676 7871 24728 7880
rect 24676 7837 24685 7871
rect 24685 7837 24719 7871
rect 24719 7837 24728 7871
rect 24676 7828 24728 7837
rect 25780 7828 25832 7880
rect 28172 7828 28224 7880
rect 31392 7828 31444 7880
rect 32312 7828 32364 7880
rect 32956 7828 33008 7880
rect 34336 7896 34388 7948
rect 35900 7896 35952 7948
rect 36636 7939 36688 7948
rect 34796 7828 34848 7880
rect 36636 7905 36645 7939
rect 36645 7905 36679 7939
rect 36679 7905 36688 7939
rect 36636 7896 36688 7905
rect 37648 7896 37700 7948
rect 37740 7896 37792 7948
rect 37924 7939 37976 7948
rect 37924 7905 37933 7939
rect 37933 7905 37967 7939
rect 37967 7905 37976 7939
rect 37924 7896 37976 7905
rect 16580 7760 16632 7812
rect 17500 7803 17552 7812
rect 17500 7769 17509 7803
rect 17509 7769 17543 7803
rect 17543 7769 17552 7803
rect 17500 7760 17552 7769
rect 20628 7760 20680 7812
rect 18420 7692 18472 7744
rect 19984 7692 20036 7744
rect 22008 7692 22060 7744
rect 23848 7692 23900 7744
rect 24400 7692 24452 7744
rect 31760 7760 31812 7812
rect 28540 7692 28592 7744
rect 30932 7692 30984 7744
rect 35992 7760 36044 7812
rect 38476 7760 38528 7812
rect 34520 7692 34572 7744
rect 36728 7692 36780 7744
rect 4246 7590 4298 7642
rect 4310 7590 4362 7642
rect 4374 7590 4426 7642
rect 4438 7590 4490 7642
rect 34966 7590 35018 7642
rect 35030 7590 35082 7642
rect 35094 7590 35146 7642
rect 35158 7590 35210 7642
rect 2964 7488 3016 7540
rect 5172 7531 5224 7540
rect 5172 7497 5181 7531
rect 5181 7497 5215 7531
rect 5215 7497 5224 7531
rect 5172 7488 5224 7497
rect 1860 7352 1912 7404
rect 3240 7352 3292 7404
rect 4068 7395 4120 7404
rect 4068 7361 4077 7395
rect 4077 7361 4111 7395
rect 4111 7361 4120 7395
rect 4068 7352 4120 7361
rect 7196 7488 7248 7540
rect 12532 7488 12584 7540
rect 14372 7488 14424 7540
rect 19984 7488 20036 7540
rect 21088 7488 21140 7540
rect 23848 7488 23900 7540
rect 23940 7488 23992 7540
rect 26240 7531 26292 7540
rect 26240 7497 26249 7531
rect 26249 7497 26283 7531
rect 26283 7497 26292 7531
rect 26240 7488 26292 7497
rect 7288 7420 7340 7472
rect 9956 7420 10008 7472
rect 18144 7420 18196 7472
rect 22284 7463 22336 7472
rect 22284 7429 22293 7463
rect 22293 7429 22327 7463
rect 22327 7429 22336 7463
rect 22284 7420 22336 7429
rect 27436 7420 27488 7472
rect 31116 7488 31168 7540
rect 31392 7488 31444 7540
rect 35808 7488 35860 7540
rect 35900 7488 35952 7540
rect 32128 7420 32180 7472
rect 2780 7284 2832 7336
rect 3792 7327 3844 7336
rect 1584 7259 1636 7268
rect 1584 7225 1593 7259
rect 1593 7225 1627 7259
rect 1627 7225 1636 7259
rect 1584 7216 1636 7225
rect 1768 7216 1820 7268
rect 3792 7293 3801 7327
rect 3801 7293 3835 7327
rect 3835 7293 3844 7327
rect 3792 7284 3844 7293
rect 7380 7327 7432 7336
rect 7380 7293 7389 7327
rect 7389 7293 7423 7327
rect 7423 7293 7432 7327
rect 7380 7284 7432 7293
rect 7656 7327 7708 7336
rect 7656 7293 7665 7327
rect 7665 7293 7699 7327
rect 7699 7293 7708 7327
rect 7656 7284 7708 7293
rect 9772 7352 9824 7404
rect 10508 7352 10560 7404
rect 12992 7395 13044 7404
rect 12992 7361 13001 7395
rect 13001 7361 13035 7395
rect 13035 7361 13044 7395
rect 12992 7352 13044 7361
rect 14004 7395 14056 7404
rect 14004 7361 14013 7395
rect 14013 7361 14047 7395
rect 14047 7361 14056 7395
rect 14004 7352 14056 7361
rect 18972 7395 19024 7404
rect 8024 7216 8076 7268
rect 9312 7284 9364 7336
rect 10692 7284 10744 7336
rect 10876 7327 10928 7336
rect 10876 7293 10885 7327
rect 10885 7293 10919 7327
rect 10919 7293 10928 7327
rect 10876 7284 10928 7293
rect 11612 7284 11664 7336
rect 12440 7327 12492 7336
rect 12440 7293 12449 7327
rect 12449 7293 12483 7327
rect 12483 7293 12492 7327
rect 12440 7284 12492 7293
rect 12900 7327 12952 7336
rect 12900 7293 12909 7327
rect 12909 7293 12943 7327
rect 12943 7293 12952 7327
rect 12900 7284 12952 7293
rect 13176 7284 13228 7336
rect 13912 7327 13964 7336
rect 13912 7293 13921 7327
rect 13921 7293 13955 7327
rect 13955 7293 13964 7327
rect 14464 7327 14516 7336
rect 13912 7284 13964 7293
rect 14464 7293 14473 7327
rect 14473 7293 14507 7327
rect 14507 7293 14516 7327
rect 14464 7284 14516 7293
rect 14648 7327 14700 7336
rect 14648 7293 14657 7327
rect 14657 7293 14691 7327
rect 14691 7293 14700 7327
rect 14648 7284 14700 7293
rect 18972 7361 18981 7395
rect 18981 7361 19015 7395
rect 19015 7361 19024 7395
rect 18972 7352 19024 7361
rect 15568 7327 15620 7336
rect 15568 7293 15577 7327
rect 15577 7293 15611 7327
rect 15611 7293 15620 7327
rect 15568 7284 15620 7293
rect 16672 7327 16724 7336
rect 16672 7293 16681 7327
rect 16681 7293 16715 7327
rect 16715 7293 16724 7327
rect 16672 7284 16724 7293
rect 14372 7216 14424 7268
rect 16948 7284 17000 7336
rect 18420 7327 18472 7336
rect 17960 7216 18012 7268
rect 18420 7293 18429 7327
rect 18429 7293 18463 7327
rect 18463 7293 18472 7327
rect 18420 7284 18472 7293
rect 19340 7284 19392 7336
rect 21732 7352 21784 7404
rect 23664 7395 23716 7404
rect 23664 7361 23673 7395
rect 23673 7361 23707 7395
rect 23707 7361 23716 7395
rect 27620 7395 27672 7404
rect 23664 7352 23716 7361
rect 27620 7361 27629 7395
rect 27629 7361 27663 7395
rect 27663 7361 27672 7395
rect 27620 7352 27672 7361
rect 28172 7395 28224 7404
rect 28172 7361 28181 7395
rect 28181 7361 28215 7395
rect 28215 7361 28224 7395
rect 28172 7352 28224 7361
rect 32404 7352 32456 7404
rect 33140 7352 33192 7404
rect 37832 7395 37884 7404
rect 37832 7361 37841 7395
rect 37841 7361 37875 7395
rect 37875 7361 37884 7395
rect 37832 7352 37884 7361
rect 19984 7327 20036 7336
rect 19984 7293 19993 7327
rect 19993 7293 20027 7327
rect 20027 7293 20036 7327
rect 20444 7327 20496 7336
rect 19984 7284 20036 7293
rect 20444 7293 20453 7327
rect 20453 7293 20487 7327
rect 20487 7293 20496 7327
rect 20444 7284 20496 7293
rect 20628 7284 20680 7336
rect 22100 7284 22152 7336
rect 22376 7327 22428 7336
rect 22376 7293 22385 7327
rect 22385 7293 22419 7327
rect 22419 7293 22428 7327
rect 22376 7284 22428 7293
rect 23204 7327 23256 7336
rect 23204 7293 23213 7327
rect 23213 7293 23247 7327
rect 23247 7293 23256 7327
rect 23204 7284 23256 7293
rect 24216 7284 24268 7336
rect 26700 7284 26752 7336
rect 27252 7284 27304 7336
rect 28080 7284 28132 7336
rect 29276 7327 29328 7336
rect 29276 7293 29285 7327
rect 29285 7293 29319 7327
rect 29319 7293 29328 7327
rect 29276 7284 29328 7293
rect 30288 7284 30340 7336
rect 34336 7284 34388 7336
rect 37740 7327 37792 7336
rect 37740 7293 37749 7327
rect 37749 7293 37783 7327
rect 37783 7293 37792 7327
rect 37740 7284 37792 7293
rect 38292 7327 38344 7336
rect 38292 7293 38301 7327
rect 38301 7293 38335 7327
rect 38335 7293 38344 7327
rect 38292 7284 38344 7293
rect 38844 7327 38896 7336
rect 38844 7293 38853 7327
rect 38853 7293 38887 7327
rect 38887 7293 38896 7327
rect 38844 7284 38896 7293
rect 21456 7216 21508 7268
rect 34704 7216 34756 7268
rect 10324 7148 10376 7200
rect 10508 7148 10560 7200
rect 12440 7148 12492 7200
rect 12624 7148 12676 7200
rect 13084 7148 13136 7200
rect 15292 7148 15344 7200
rect 15476 7148 15528 7200
rect 16580 7148 16632 7200
rect 21088 7148 21140 7200
rect 22928 7148 22980 7200
rect 23204 7148 23256 7200
rect 27160 7148 27212 7200
rect 29092 7148 29144 7200
rect 19606 7046 19658 7098
rect 19670 7046 19722 7098
rect 19734 7046 19786 7098
rect 19798 7046 19850 7098
rect 7840 6987 7892 6996
rect 7840 6953 7849 6987
rect 7849 6953 7883 6987
rect 7883 6953 7892 6987
rect 7840 6944 7892 6953
rect 10232 6944 10284 6996
rect 18144 6944 18196 6996
rect 18236 6944 18288 6996
rect 29276 6987 29328 6996
rect 5172 6876 5224 6928
rect 2412 6851 2464 6860
rect 2412 6817 2421 6851
rect 2421 6817 2455 6851
rect 2455 6817 2464 6851
rect 2412 6808 2464 6817
rect 2504 6808 2556 6860
rect 3608 6808 3660 6860
rect 5080 6851 5132 6860
rect 5080 6817 5089 6851
rect 5089 6817 5123 6851
rect 5123 6817 5132 6851
rect 5080 6808 5132 6817
rect 5356 6808 5408 6860
rect 7288 6808 7340 6860
rect 9496 6808 9548 6860
rect 10140 6808 10192 6860
rect 4620 6783 4672 6792
rect 4620 6749 4629 6783
rect 4629 6749 4663 6783
rect 4663 6749 4672 6783
rect 4620 6740 4672 6749
rect 4712 6740 4764 6792
rect 6276 6783 6328 6792
rect 6276 6749 6285 6783
rect 6285 6749 6319 6783
rect 6319 6749 6328 6783
rect 6276 6740 6328 6749
rect 10508 6808 10560 6860
rect 12072 6808 12124 6860
rect 12900 6808 12952 6860
rect 14464 6876 14516 6928
rect 29276 6953 29285 6987
rect 29285 6953 29319 6987
rect 29319 6953 29328 6987
rect 29276 6944 29328 6953
rect 13084 6783 13136 6792
rect 13084 6749 13093 6783
rect 13093 6749 13127 6783
rect 13127 6749 13136 6783
rect 13084 6740 13136 6749
rect 14004 6808 14056 6860
rect 15476 6808 15528 6860
rect 17500 6808 17552 6860
rect 18328 6808 18380 6860
rect 2964 6715 3016 6724
rect 2964 6681 2973 6715
rect 2973 6681 3007 6715
rect 3007 6681 3016 6715
rect 2964 6672 3016 6681
rect 10324 6672 10376 6724
rect 12072 6672 12124 6724
rect 18236 6740 18288 6792
rect 19340 6783 19392 6792
rect 19340 6749 19349 6783
rect 19349 6749 19383 6783
rect 19383 6749 19392 6783
rect 19340 6740 19392 6749
rect 19984 6808 20036 6860
rect 20444 6808 20496 6860
rect 21088 6851 21140 6860
rect 21088 6817 21097 6851
rect 21097 6817 21131 6851
rect 21131 6817 21140 6851
rect 21088 6808 21140 6817
rect 20076 6740 20128 6792
rect 21272 6783 21324 6792
rect 21272 6749 21281 6783
rect 21281 6749 21315 6783
rect 21315 6749 21324 6783
rect 21272 6740 21324 6749
rect 11980 6604 12032 6656
rect 20904 6672 20956 6724
rect 22100 6808 22152 6860
rect 23204 6876 23256 6928
rect 23480 6808 23532 6860
rect 23756 6851 23808 6860
rect 23756 6817 23765 6851
rect 23765 6817 23799 6851
rect 23799 6817 23808 6851
rect 23756 6808 23808 6817
rect 24216 6876 24268 6928
rect 24492 6876 24544 6928
rect 26792 6876 26844 6928
rect 24584 6808 24636 6860
rect 24768 6808 24820 6860
rect 27252 6808 27304 6860
rect 31484 6851 31536 6860
rect 31484 6817 31493 6851
rect 31493 6817 31527 6851
rect 31527 6817 31536 6851
rect 31484 6808 31536 6817
rect 32588 6808 32640 6860
rect 33232 6808 33284 6860
rect 34612 6808 34664 6860
rect 25320 6740 25372 6792
rect 27436 6740 27488 6792
rect 27896 6740 27948 6792
rect 29920 6740 29972 6792
rect 30840 6783 30892 6792
rect 30840 6749 30849 6783
rect 30849 6749 30883 6783
rect 30883 6749 30892 6783
rect 30840 6740 30892 6749
rect 33968 6783 34020 6792
rect 24676 6672 24728 6724
rect 16764 6604 16816 6656
rect 22192 6604 22244 6656
rect 24768 6604 24820 6656
rect 25044 6604 25096 6656
rect 26240 6604 26292 6656
rect 33140 6672 33192 6724
rect 33968 6749 33977 6783
rect 33977 6749 34011 6783
rect 34011 6749 34020 6783
rect 33968 6740 34020 6749
rect 34428 6783 34480 6792
rect 34428 6749 34437 6783
rect 34437 6749 34471 6783
rect 34471 6749 34480 6783
rect 34428 6740 34480 6749
rect 36268 6808 36320 6860
rect 36728 6851 36780 6860
rect 35440 6783 35492 6792
rect 35440 6749 35449 6783
rect 35449 6749 35483 6783
rect 35483 6749 35492 6783
rect 35440 6740 35492 6749
rect 35900 6783 35952 6792
rect 35900 6749 35909 6783
rect 35909 6749 35943 6783
rect 35943 6749 35952 6783
rect 35900 6740 35952 6749
rect 36176 6740 36228 6792
rect 36728 6817 36737 6851
rect 36737 6817 36771 6851
rect 36771 6817 36780 6851
rect 36728 6808 36780 6817
rect 38016 6851 38068 6860
rect 38016 6817 38025 6851
rect 38025 6817 38059 6851
rect 38059 6817 38068 6851
rect 38016 6808 38068 6817
rect 38384 6851 38436 6860
rect 38384 6817 38393 6851
rect 38393 6817 38427 6851
rect 38427 6817 38436 6851
rect 38384 6808 38436 6817
rect 38476 6808 38528 6860
rect 37740 6672 37792 6724
rect 27344 6604 27396 6656
rect 28172 6604 28224 6656
rect 31208 6604 31260 6656
rect 31392 6604 31444 6656
rect 32312 6604 32364 6656
rect 4246 6502 4298 6554
rect 4310 6502 4362 6554
rect 4374 6502 4426 6554
rect 4438 6502 4490 6554
rect 34966 6502 35018 6554
rect 35030 6502 35082 6554
rect 35094 6502 35146 6554
rect 35158 6502 35210 6554
rect 3608 6332 3660 6384
rect 2412 6264 2464 6316
rect 3332 6239 3384 6248
rect 3332 6205 3341 6239
rect 3341 6205 3375 6239
rect 3375 6205 3384 6239
rect 3332 6196 3384 6205
rect 3608 6128 3660 6180
rect 5080 6400 5132 6452
rect 9496 6443 9548 6452
rect 9496 6409 9505 6443
rect 9505 6409 9539 6443
rect 9539 6409 9548 6443
rect 9496 6400 9548 6409
rect 13544 6443 13596 6452
rect 13544 6409 13553 6443
rect 13553 6409 13587 6443
rect 13587 6409 13596 6443
rect 13544 6400 13596 6409
rect 14096 6400 14148 6452
rect 14924 6400 14976 6452
rect 15844 6400 15896 6452
rect 20076 6443 20128 6452
rect 11612 6332 11664 6384
rect 16672 6375 16724 6384
rect 6276 6264 6328 6316
rect 8300 6264 8352 6316
rect 8576 6264 8628 6316
rect 14280 6307 14332 6316
rect 14280 6273 14289 6307
rect 14289 6273 14323 6307
rect 14323 6273 14332 6307
rect 14280 6264 14332 6273
rect 4160 6196 4212 6248
rect 4896 6239 4948 6248
rect 4528 6128 4580 6180
rect 3148 6060 3200 6112
rect 3792 6060 3844 6112
rect 4896 6205 4905 6239
rect 4905 6205 4939 6239
rect 4939 6205 4948 6239
rect 4896 6196 4948 6205
rect 8208 6239 8260 6248
rect 8208 6205 8217 6239
rect 8217 6205 8251 6239
rect 8251 6205 8260 6239
rect 8208 6196 8260 6205
rect 11428 6196 11480 6248
rect 13268 6196 13320 6248
rect 13820 6196 13872 6248
rect 13912 6196 13964 6248
rect 14556 6239 14608 6248
rect 14556 6205 14565 6239
rect 14565 6205 14599 6239
rect 14599 6205 14608 6239
rect 14556 6196 14608 6205
rect 14648 6196 14700 6248
rect 15568 6196 15620 6248
rect 16672 6341 16681 6375
rect 16681 6341 16715 6375
rect 16715 6341 16724 6375
rect 16672 6332 16724 6341
rect 18972 6307 19024 6316
rect 16856 6196 16908 6248
rect 18052 6239 18104 6248
rect 18052 6205 18061 6239
rect 18061 6205 18095 6239
rect 18095 6205 18104 6239
rect 18052 6196 18104 6205
rect 18512 6196 18564 6248
rect 18972 6273 18981 6307
rect 18981 6273 19015 6307
rect 19015 6273 19024 6307
rect 18972 6264 19024 6273
rect 20076 6409 20085 6443
rect 20085 6409 20119 6443
rect 20119 6409 20128 6443
rect 20076 6400 20128 6409
rect 20720 6400 20772 6452
rect 23388 6400 23440 6452
rect 23664 6400 23716 6452
rect 26700 6443 26752 6452
rect 24676 6332 24728 6384
rect 20352 6196 20404 6248
rect 20904 6196 20956 6248
rect 21272 6196 21324 6248
rect 22192 6196 22244 6248
rect 24584 6264 24636 6316
rect 24400 6239 24452 6248
rect 24400 6205 24409 6239
rect 24409 6205 24443 6239
rect 24443 6205 24452 6239
rect 24400 6196 24452 6205
rect 25044 6264 25096 6316
rect 26700 6409 26709 6443
rect 26709 6409 26743 6443
rect 26743 6409 26752 6443
rect 26700 6400 26752 6409
rect 27436 6375 27488 6384
rect 27436 6341 27445 6375
rect 27445 6341 27479 6375
rect 27479 6341 27488 6375
rect 27436 6332 27488 6341
rect 31484 6400 31536 6452
rect 25780 6264 25832 6316
rect 24768 6196 24820 6248
rect 25596 6239 25648 6248
rect 25596 6205 25605 6239
rect 25605 6205 25639 6239
rect 25639 6205 25648 6239
rect 25596 6196 25648 6205
rect 26240 6196 26292 6248
rect 31300 6332 31352 6384
rect 32312 6400 32364 6452
rect 33140 6400 33192 6452
rect 35992 6400 36044 6452
rect 38844 6443 38896 6452
rect 29920 6264 29972 6316
rect 28540 6239 28592 6248
rect 16764 6128 16816 6180
rect 5264 6060 5316 6112
rect 12532 6103 12584 6112
rect 12532 6069 12541 6103
rect 12541 6069 12575 6103
rect 12575 6069 12584 6103
rect 12532 6060 12584 6069
rect 25412 6128 25464 6180
rect 28540 6205 28549 6239
rect 28549 6205 28583 6239
rect 28583 6205 28592 6239
rect 28540 6196 28592 6205
rect 29092 6196 29144 6248
rect 29184 6196 29236 6248
rect 30196 6239 30248 6248
rect 30196 6205 30205 6239
rect 30205 6205 30239 6239
rect 30239 6205 30248 6239
rect 30196 6196 30248 6205
rect 30288 6239 30340 6248
rect 30288 6205 30297 6239
rect 30297 6205 30331 6239
rect 30331 6205 30340 6239
rect 31392 6264 31444 6316
rect 34428 6264 34480 6316
rect 30288 6196 30340 6205
rect 32128 6196 32180 6248
rect 32404 6239 32456 6248
rect 32404 6205 32413 6239
rect 32413 6205 32447 6239
rect 32447 6205 32456 6239
rect 32404 6196 32456 6205
rect 32956 6196 33008 6248
rect 33968 6196 34020 6248
rect 36084 6264 36136 6316
rect 38844 6409 38853 6443
rect 38853 6409 38887 6443
rect 38887 6409 38896 6443
rect 38844 6400 38896 6409
rect 37740 6307 37792 6316
rect 37740 6273 37749 6307
rect 37749 6273 37783 6307
rect 37783 6273 37792 6307
rect 37740 6264 37792 6273
rect 37372 6196 37424 6248
rect 30380 6128 30432 6180
rect 17776 6060 17828 6112
rect 20904 6060 20956 6112
rect 25044 6060 25096 6112
rect 29828 6060 29880 6112
rect 32312 6128 32364 6180
rect 33968 6060 34020 6112
rect 19606 5958 19658 6010
rect 19670 5958 19722 6010
rect 19734 5958 19786 6010
rect 19798 5958 19850 6010
rect 2504 5899 2556 5908
rect 2504 5865 2513 5899
rect 2513 5865 2547 5899
rect 2547 5865 2556 5899
rect 2504 5856 2556 5865
rect 3976 5788 4028 5840
rect 8208 5856 8260 5908
rect 12900 5856 12952 5908
rect 14556 5856 14608 5908
rect 16856 5856 16908 5908
rect 17960 5856 18012 5908
rect 24584 5899 24636 5908
rect 24584 5865 24593 5899
rect 24593 5865 24627 5899
rect 24627 5865 24636 5899
rect 24584 5856 24636 5865
rect 3332 5720 3384 5772
rect 4160 5720 4212 5772
rect 4988 5720 5040 5772
rect 5264 5720 5316 5772
rect 9680 5720 9732 5772
rect 4712 5652 4764 5704
rect 6276 5652 6328 5704
rect 4528 5584 4580 5636
rect 4804 5584 4856 5636
rect 9956 5763 10008 5772
rect 9956 5729 9965 5763
rect 9965 5729 9999 5763
rect 9999 5729 10008 5763
rect 10324 5763 10376 5772
rect 9956 5720 10008 5729
rect 10324 5729 10333 5763
rect 10333 5729 10367 5763
rect 10367 5729 10376 5763
rect 10324 5720 10376 5729
rect 10968 5720 11020 5772
rect 11980 5763 12032 5772
rect 11980 5729 11989 5763
rect 11989 5729 12023 5763
rect 12023 5729 12032 5763
rect 11980 5720 12032 5729
rect 11888 5652 11940 5704
rect 12624 5652 12676 5704
rect 12808 5652 12860 5704
rect 10416 5584 10468 5636
rect 13728 5584 13780 5636
rect 5356 5516 5408 5568
rect 10784 5516 10836 5568
rect 15292 5763 15344 5772
rect 15292 5729 15301 5763
rect 15301 5729 15335 5763
rect 15335 5729 15344 5763
rect 15292 5720 15344 5729
rect 15660 5584 15712 5636
rect 16304 5720 16356 5772
rect 17040 5720 17092 5772
rect 17684 5720 17736 5772
rect 18328 5788 18380 5840
rect 19340 5720 19392 5772
rect 20904 5763 20956 5772
rect 20904 5729 20913 5763
rect 20913 5729 20947 5763
rect 20947 5729 20956 5763
rect 20904 5720 20956 5729
rect 21272 5763 21324 5772
rect 21272 5729 21281 5763
rect 21281 5729 21315 5763
rect 21315 5729 21324 5763
rect 21272 5720 21324 5729
rect 22192 5720 22244 5772
rect 22744 5720 22796 5772
rect 28632 5856 28684 5908
rect 29736 5788 29788 5840
rect 36176 5831 36228 5840
rect 24860 5720 24912 5772
rect 27068 5763 27120 5772
rect 17224 5695 17276 5704
rect 17224 5661 17233 5695
rect 17233 5661 17267 5695
rect 17267 5661 17276 5695
rect 17224 5652 17276 5661
rect 17868 5695 17920 5704
rect 17868 5661 17877 5695
rect 17877 5661 17911 5695
rect 17911 5661 17920 5695
rect 17868 5652 17920 5661
rect 20352 5652 20404 5704
rect 22100 5652 22152 5704
rect 23020 5695 23072 5704
rect 23020 5661 23029 5695
rect 23029 5661 23063 5695
rect 23063 5661 23072 5695
rect 23020 5652 23072 5661
rect 25044 5652 25096 5704
rect 18880 5627 18932 5636
rect 18880 5593 18889 5627
rect 18889 5593 18923 5627
rect 18923 5593 18932 5627
rect 18880 5584 18932 5593
rect 21272 5584 21324 5636
rect 24400 5584 24452 5636
rect 27068 5729 27077 5763
rect 27077 5729 27111 5763
rect 27111 5729 27120 5763
rect 27068 5720 27120 5729
rect 27160 5720 27212 5772
rect 29276 5720 29328 5772
rect 30380 5720 30432 5772
rect 30840 5720 30892 5772
rect 31300 5720 31352 5772
rect 31852 5720 31904 5772
rect 26516 5695 26568 5704
rect 26516 5661 26525 5695
rect 26525 5661 26559 5695
rect 26559 5661 26568 5695
rect 26516 5652 26568 5661
rect 28264 5652 28316 5704
rect 27068 5584 27120 5636
rect 28816 5652 28868 5704
rect 30564 5652 30616 5704
rect 31484 5652 31536 5704
rect 31668 5652 31720 5704
rect 32956 5763 33008 5772
rect 32956 5729 32965 5763
rect 32965 5729 32999 5763
rect 32999 5729 33008 5763
rect 32956 5720 33008 5729
rect 32128 5695 32180 5704
rect 32128 5661 32137 5695
rect 32137 5661 32171 5695
rect 32171 5661 32180 5695
rect 32128 5652 32180 5661
rect 36176 5797 36185 5831
rect 36185 5797 36219 5831
rect 36219 5797 36228 5831
rect 36176 5788 36228 5797
rect 35900 5720 35952 5772
rect 37372 5856 37424 5908
rect 38384 5856 38436 5908
rect 37004 5763 37056 5772
rect 37004 5729 37013 5763
rect 37013 5729 37047 5763
rect 37047 5729 37056 5763
rect 37004 5720 37056 5729
rect 37832 5763 37884 5772
rect 37832 5729 37841 5763
rect 37841 5729 37875 5763
rect 37875 5729 37884 5763
rect 37832 5720 37884 5729
rect 38200 5763 38252 5772
rect 38200 5729 38209 5763
rect 38209 5729 38243 5763
rect 38243 5729 38252 5763
rect 38200 5720 38252 5729
rect 38844 5720 38896 5772
rect 32404 5584 32456 5636
rect 32956 5584 33008 5636
rect 35992 5652 36044 5704
rect 35440 5627 35492 5636
rect 35440 5593 35449 5627
rect 35449 5593 35483 5627
rect 35483 5593 35492 5627
rect 35440 5584 35492 5593
rect 19248 5516 19300 5568
rect 23296 5516 23348 5568
rect 28172 5516 28224 5568
rect 28356 5516 28408 5568
rect 4246 5414 4298 5466
rect 4310 5414 4362 5466
rect 4374 5414 4426 5466
rect 4438 5414 4490 5466
rect 34966 5414 35018 5466
rect 35030 5414 35082 5466
rect 35094 5414 35146 5466
rect 35158 5414 35210 5466
rect 3332 5312 3384 5364
rect 9680 5355 9732 5364
rect 9680 5321 9689 5355
rect 9689 5321 9723 5355
rect 9723 5321 9732 5355
rect 9680 5312 9732 5321
rect 10600 5312 10652 5364
rect 10784 5312 10836 5364
rect 2964 5176 3016 5228
rect 3148 5108 3200 5160
rect 5080 5244 5132 5296
rect 4712 5219 4764 5228
rect 4712 5185 4721 5219
rect 4721 5185 4755 5219
rect 4755 5185 4764 5219
rect 4712 5176 4764 5185
rect 5172 5176 5224 5228
rect 8300 5176 8352 5228
rect 11428 5244 11480 5296
rect 12532 5176 12584 5228
rect 4528 4972 4580 5024
rect 5356 5108 5408 5160
rect 10416 5151 10468 5160
rect 5172 5040 5224 5092
rect 10416 5117 10425 5151
rect 10425 5117 10459 5151
rect 10459 5117 10468 5151
rect 10416 5108 10468 5117
rect 10600 5108 10652 5160
rect 10784 5108 10836 5160
rect 10968 5151 11020 5160
rect 10968 5117 10977 5151
rect 10977 5117 11011 5151
rect 11011 5117 11020 5151
rect 10968 5108 11020 5117
rect 12072 5108 12124 5160
rect 12440 5108 12492 5160
rect 12624 5151 12676 5160
rect 12624 5117 12633 5151
rect 12633 5117 12667 5151
rect 12667 5117 12676 5151
rect 12624 5108 12676 5117
rect 11060 5040 11112 5092
rect 13912 5108 13964 5160
rect 15200 5176 15252 5228
rect 14648 5151 14700 5160
rect 14648 5117 14657 5151
rect 14657 5117 14691 5151
rect 14691 5117 14700 5151
rect 14648 5108 14700 5117
rect 15016 5151 15068 5160
rect 15016 5117 15025 5151
rect 15025 5117 15059 5151
rect 15059 5117 15068 5151
rect 15016 5108 15068 5117
rect 15568 5151 15620 5160
rect 15568 5117 15577 5151
rect 15577 5117 15611 5151
rect 15611 5117 15620 5151
rect 15568 5108 15620 5117
rect 15844 5108 15896 5160
rect 16212 5151 16264 5160
rect 16212 5117 16221 5151
rect 16221 5117 16255 5151
rect 16255 5117 16264 5151
rect 16212 5108 16264 5117
rect 16396 5108 16448 5160
rect 16764 5151 16816 5160
rect 16764 5117 16773 5151
rect 16773 5117 16807 5151
rect 16807 5117 16816 5151
rect 16764 5108 16816 5117
rect 5356 4972 5408 5024
rect 5816 4972 5868 5024
rect 12716 5015 12768 5024
rect 12716 4981 12725 5015
rect 12725 4981 12759 5015
rect 12759 4981 12768 5015
rect 12716 4972 12768 4981
rect 16580 4972 16632 5024
rect 18788 5312 18840 5364
rect 18880 5176 18932 5228
rect 17960 5108 18012 5160
rect 18512 5151 18564 5160
rect 18512 5117 18521 5151
rect 18521 5117 18555 5151
rect 18555 5117 18564 5151
rect 18512 5108 18564 5117
rect 19432 5108 19484 5160
rect 24492 5312 24544 5364
rect 27252 5355 27304 5364
rect 27252 5321 27261 5355
rect 27261 5321 27295 5355
rect 27295 5321 27304 5355
rect 27252 5312 27304 5321
rect 28264 5312 28316 5364
rect 28816 5312 28868 5364
rect 29368 5312 29420 5364
rect 31760 5355 31812 5364
rect 31760 5321 31769 5355
rect 31769 5321 31803 5355
rect 31803 5321 31812 5355
rect 31760 5312 31812 5321
rect 34796 5312 34848 5364
rect 22468 5244 22520 5296
rect 26516 5176 26568 5228
rect 30564 5176 30616 5228
rect 31392 5176 31444 5228
rect 31852 5244 31904 5296
rect 34612 5244 34664 5296
rect 37004 5312 37056 5364
rect 38016 5312 38068 5364
rect 22100 5151 22152 5160
rect 22100 5117 22109 5151
rect 22109 5117 22143 5151
rect 22143 5117 22152 5151
rect 22744 5151 22796 5160
rect 22100 5108 22152 5117
rect 22744 5117 22753 5151
rect 22753 5117 22787 5151
rect 22787 5117 22796 5151
rect 22744 5108 22796 5117
rect 22836 5108 22888 5160
rect 25228 5151 25280 5160
rect 25228 5117 25237 5151
rect 25237 5117 25271 5151
rect 25271 5117 25280 5151
rect 25228 5108 25280 5117
rect 25504 5108 25556 5160
rect 25780 5108 25832 5160
rect 26608 5108 26660 5160
rect 29092 5108 29144 5160
rect 29276 5151 29328 5160
rect 29276 5117 29285 5151
rect 29285 5117 29319 5151
rect 29319 5117 29328 5151
rect 29276 5108 29328 5117
rect 32128 5108 32180 5160
rect 33968 5176 34020 5228
rect 34704 5176 34756 5228
rect 23112 5040 23164 5092
rect 25596 5040 25648 5092
rect 31484 5040 31536 5092
rect 34520 5108 34572 5160
rect 35992 5176 36044 5228
rect 36360 5219 36412 5228
rect 36360 5185 36369 5219
rect 36369 5185 36403 5219
rect 36403 5185 36412 5219
rect 36360 5176 36412 5185
rect 37832 5176 37884 5228
rect 37648 5108 37700 5160
rect 32680 5040 32732 5092
rect 19432 4972 19484 5024
rect 19606 4870 19658 4922
rect 19670 4870 19722 4922
rect 19734 4870 19786 4922
rect 19798 4870 19850 4922
rect 4528 4675 4580 4684
rect 4528 4641 4537 4675
rect 4537 4641 4571 4675
rect 4571 4641 4580 4675
rect 4528 4632 4580 4641
rect 5172 4675 5224 4684
rect 5172 4641 5181 4675
rect 5181 4641 5215 4675
rect 5215 4641 5224 4675
rect 5172 4632 5224 4641
rect 10416 4768 10468 4820
rect 10416 4675 10468 4684
rect 10416 4641 10425 4675
rect 10425 4641 10459 4675
rect 10459 4641 10468 4675
rect 10968 4700 11020 4752
rect 10416 4632 10468 4641
rect 11060 4675 11112 4684
rect 11060 4641 11069 4675
rect 11069 4641 11103 4675
rect 11103 4641 11112 4675
rect 11060 4632 11112 4641
rect 14188 4675 14240 4684
rect 14188 4641 14197 4675
rect 14197 4641 14231 4675
rect 14231 4641 14240 4675
rect 14188 4632 14240 4641
rect 4988 4564 5040 4616
rect 6828 4607 6880 4616
rect 6828 4573 6837 4607
rect 6837 4573 6871 4607
rect 6871 4573 6880 4607
rect 6828 4564 6880 4573
rect 9588 4564 9640 4616
rect 11888 4564 11940 4616
rect 13912 4564 13964 4616
rect 14096 4607 14148 4616
rect 14096 4573 14105 4607
rect 14105 4573 14139 4607
rect 14139 4573 14148 4607
rect 14096 4564 14148 4573
rect 15016 4768 15068 4820
rect 22468 4768 22520 4820
rect 22836 4811 22888 4820
rect 22836 4777 22845 4811
rect 22845 4777 22879 4811
rect 22879 4777 22888 4811
rect 22836 4768 22888 4777
rect 15660 4632 15712 4684
rect 16304 4607 16356 4616
rect 16304 4573 16313 4607
rect 16313 4573 16347 4607
rect 16347 4573 16356 4607
rect 16304 4564 16356 4573
rect 20628 4700 20680 4752
rect 16580 4675 16632 4684
rect 16580 4641 16589 4675
rect 16589 4641 16623 4675
rect 16623 4641 16632 4675
rect 16580 4632 16632 4641
rect 18972 4675 19024 4684
rect 18972 4641 18981 4675
rect 18981 4641 19015 4675
rect 19015 4641 19024 4675
rect 18972 4632 19024 4641
rect 19156 4632 19208 4684
rect 23112 4700 23164 4752
rect 24400 4675 24452 4684
rect 24400 4641 24409 4675
rect 24409 4641 24443 4675
rect 24443 4641 24452 4675
rect 24400 4632 24452 4641
rect 24492 4632 24544 4684
rect 24768 4632 24820 4684
rect 19708 4607 19760 4616
rect 16212 4496 16264 4548
rect 19708 4573 19717 4607
rect 19717 4573 19751 4607
rect 19751 4573 19760 4607
rect 19708 4564 19760 4573
rect 21272 4607 21324 4616
rect 21272 4573 21281 4607
rect 21281 4573 21315 4607
rect 21315 4573 21324 4607
rect 21272 4564 21324 4573
rect 22836 4564 22888 4616
rect 23848 4607 23900 4616
rect 23848 4573 23857 4607
rect 23857 4573 23891 4607
rect 23891 4573 23900 4607
rect 23848 4564 23900 4573
rect 26516 4607 26568 4616
rect 26516 4573 26525 4607
rect 26525 4573 26559 4607
rect 26559 4573 26568 4607
rect 26516 4564 26568 4573
rect 27068 4607 27120 4616
rect 27068 4573 27077 4607
rect 27077 4573 27111 4607
rect 27111 4573 27120 4607
rect 27068 4564 27120 4573
rect 27344 4675 27396 4684
rect 27344 4641 27353 4675
rect 27353 4641 27387 4675
rect 27387 4641 27396 4675
rect 27344 4632 27396 4641
rect 27896 4632 27948 4684
rect 29276 4632 29328 4684
rect 38200 4768 38252 4820
rect 32128 4743 32180 4752
rect 32128 4709 32137 4743
rect 32137 4709 32171 4743
rect 32171 4709 32180 4743
rect 32128 4700 32180 4709
rect 33416 4700 33468 4752
rect 29736 4632 29788 4684
rect 32036 4632 32088 4684
rect 32680 4675 32732 4684
rect 32680 4641 32689 4675
rect 32689 4641 32723 4675
rect 32723 4641 32732 4675
rect 32680 4632 32732 4641
rect 34336 4632 34388 4684
rect 36084 4675 36136 4684
rect 28264 4564 28316 4616
rect 30380 4564 30432 4616
rect 31668 4564 31720 4616
rect 7564 4428 7616 4480
rect 12348 4428 12400 4480
rect 15568 4428 15620 4480
rect 16488 4428 16540 4480
rect 17776 4428 17828 4480
rect 18052 4428 18104 4480
rect 30012 4428 30064 4480
rect 30840 4428 30892 4480
rect 34520 4564 34572 4616
rect 34704 4564 34756 4616
rect 35624 4607 35676 4616
rect 35624 4573 35633 4607
rect 35633 4573 35667 4607
rect 35667 4573 35676 4607
rect 35624 4564 35676 4573
rect 36084 4641 36093 4675
rect 36093 4641 36127 4675
rect 36127 4641 36136 4675
rect 36084 4632 36136 4641
rect 37648 4632 37700 4684
rect 35992 4564 36044 4616
rect 36268 4564 36320 4616
rect 4246 4326 4298 4378
rect 4310 4326 4362 4378
rect 4374 4326 4426 4378
rect 4438 4326 4490 4378
rect 34966 4326 35018 4378
rect 35030 4326 35082 4378
rect 35094 4326 35146 4378
rect 35158 4326 35210 4378
rect 10416 4224 10468 4276
rect 20904 4224 20956 4276
rect 16396 4156 16448 4208
rect 19156 4156 19208 4208
rect 24860 4156 24912 4208
rect 25504 4156 25556 4208
rect 4804 4088 4856 4140
rect 4896 4088 4948 4140
rect 6276 4131 6328 4140
rect 6276 4097 6285 4131
rect 6285 4097 6319 4131
rect 6319 4097 6328 4131
rect 6276 4088 6328 4097
rect 9680 4088 9732 4140
rect 4620 4063 4672 4072
rect 4620 4029 4629 4063
rect 4629 4029 4663 4063
rect 4663 4029 4672 4063
rect 4620 4020 4672 4029
rect 5816 4063 5868 4072
rect 5816 4029 5825 4063
rect 5825 4029 5859 4063
rect 5859 4029 5868 4063
rect 5816 4020 5868 4029
rect 7564 4063 7616 4072
rect 7564 4029 7573 4063
rect 7573 4029 7607 4063
rect 7607 4029 7616 4063
rect 7564 4020 7616 4029
rect 8484 4063 8536 4072
rect 4712 3952 4764 4004
rect 4988 3952 5040 4004
rect 6828 3952 6880 4004
rect 8484 4029 8493 4063
rect 8493 4029 8527 4063
rect 8527 4029 8536 4063
rect 8484 4020 8536 4029
rect 8760 4063 8812 4072
rect 8760 4029 8769 4063
rect 8769 4029 8803 4063
rect 8803 4029 8812 4063
rect 8760 4020 8812 4029
rect 10968 4020 11020 4072
rect 13820 4088 13872 4140
rect 14280 4131 14332 4140
rect 11244 4063 11296 4072
rect 11244 4029 11253 4063
rect 11253 4029 11287 4063
rect 11287 4029 11296 4063
rect 11244 4020 11296 4029
rect 12808 4063 12860 4072
rect 12808 4029 12817 4063
rect 12817 4029 12851 4063
rect 12851 4029 12860 4063
rect 12808 4020 12860 4029
rect 14280 4097 14289 4131
rect 14289 4097 14323 4131
rect 14323 4097 14332 4131
rect 14280 4088 14332 4097
rect 15292 4088 15344 4140
rect 7748 3952 7800 4004
rect 10140 3995 10192 4004
rect 10140 3961 10149 3995
rect 10149 3961 10183 3995
rect 10183 3961 10192 3995
rect 10140 3952 10192 3961
rect 7472 3884 7524 3936
rect 16304 4020 16356 4072
rect 16672 4063 16724 4072
rect 16672 4029 16681 4063
rect 16681 4029 16715 4063
rect 16715 4029 16724 4063
rect 16672 4020 16724 4029
rect 17040 4063 17092 4072
rect 17040 4029 17049 4063
rect 17049 4029 17083 4063
rect 17083 4029 17092 4063
rect 17040 4020 17092 4029
rect 18052 4063 18104 4072
rect 18052 4029 18061 4063
rect 18061 4029 18095 4063
rect 18095 4029 18104 4063
rect 18052 4020 18104 4029
rect 18972 4088 19024 4140
rect 19708 4088 19760 4140
rect 20720 4088 20772 4140
rect 19340 4063 19392 4072
rect 19340 4029 19349 4063
rect 19349 4029 19383 4063
rect 19383 4029 19392 4063
rect 19340 4020 19392 4029
rect 20352 4020 20404 4072
rect 22100 4063 22152 4072
rect 22100 4029 22109 4063
rect 22109 4029 22143 4063
rect 22143 4029 22152 4063
rect 22100 4020 22152 4029
rect 13544 3995 13596 4004
rect 13544 3961 13553 3995
rect 13553 3961 13587 3995
rect 13587 3961 13596 3995
rect 13544 3952 13596 3961
rect 14556 3884 14608 3936
rect 16120 3884 16172 3936
rect 20628 3884 20680 3936
rect 22836 4088 22888 4140
rect 23848 4088 23900 4140
rect 23480 4020 23532 4072
rect 24492 4063 24544 4072
rect 24492 4029 24501 4063
rect 24501 4029 24535 4063
rect 24535 4029 24544 4063
rect 24492 4020 24544 4029
rect 24860 4020 24912 4072
rect 25044 4088 25096 4140
rect 25412 4088 25464 4140
rect 26516 4088 26568 4140
rect 28356 4156 28408 4208
rect 35992 4224 36044 4276
rect 30380 4088 30432 4140
rect 30564 4131 30616 4140
rect 30564 4097 30573 4131
rect 30573 4097 30607 4131
rect 30607 4097 30616 4131
rect 30564 4088 30616 4097
rect 30840 4131 30892 4140
rect 30840 4097 30849 4131
rect 30849 4097 30883 4131
rect 30883 4097 30892 4131
rect 30840 4088 30892 4097
rect 33600 4088 33652 4140
rect 26608 4063 26660 4072
rect 26608 4029 26617 4063
rect 26617 4029 26651 4063
rect 26651 4029 26660 4063
rect 26608 4020 26660 4029
rect 27436 4063 27488 4072
rect 27436 4029 27445 4063
rect 27445 4029 27479 4063
rect 27479 4029 27488 4063
rect 27436 4020 27488 4029
rect 29092 4020 29144 4072
rect 27160 3884 27212 3936
rect 27528 3952 27580 4004
rect 32588 4020 32640 4072
rect 33232 4063 33284 4072
rect 33232 4029 33241 4063
rect 33241 4029 33275 4063
rect 33275 4029 33284 4063
rect 33232 4020 33284 4029
rect 33416 4020 33468 4072
rect 33692 4063 33744 4072
rect 33692 4029 33701 4063
rect 33701 4029 33735 4063
rect 33735 4029 33744 4063
rect 33692 4020 33744 4029
rect 33876 4020 33928 4072
rect 34612 4088 34664 4140
rect 35624 4088 35676 4140
rect 34428 4020 34480 4072
rect 38936 4131 38988 4140
rect 38936 4097 38945 4131
rect 38945 4097 38979 4131
rect 38979 4097 38988 4131
rect 38936 4088 38988 4097
rect 32680 3995 32732 4004
rect 32680 3961 32689 3995
rect 32689 3961 32723 3995
rect 32723 3961 32732 3995
rect 32680 3952 32732 3961
rect 34336 3952 34388 4004
rect 31300 3884 31352 3936
rect 32036 3884 32088 3936
rect 33692 3884 33744 3936
rect 35440 3884 35492 3936
rect 37740 4063 37792 4072
rect 37740 4029 37749 4063
rect 37749 4029 37783 4063
rect 37783 4029 37792 4063
rect 37740 4020 37792 4029
rect 19606 3782 19658 3834
rect 19670 3782 19722 3834
rect 19734 3782 19786 3834
rect 19798 3782 19850 3834
rect 9680 3680 9732 3732
rect 14832 3680 14884 3732
rect 17040 3680 17092 3732
rect 23572 3680 23624 3732
rect 25136 3680 25188 3732
rect 27436 3680 27488 3732
rect 31208 3680 31260 3732
rect 31300 3680 31352 3732
rect 8760 3612 8812 3664
rect 24492 3612 24544 3664
rect 6828 3544 6880 3596
rect 7472 3587 7524 3596
rect 7472 3553 7481 3587
rect 7481 3553 7515 3587
rect 7515 3553 7524 3587
rect 7472 3544 7524 3553
rect 10968 3587 11020 3596
rect 10968 3553 10977 3587
rect 10977 3553 11011 3587
rect 11011 3553 11020 3587
rect 10968 3544 11020 3553
rect 12532 3544 12584 3596
rect 13544 3544 13596 3596
rect 17224 3544 17276 3596
rect 572 3476 624 3528
rect 1768 3476 1820 3528
rect 9680 3519 9732 3528
rect 9680 3485 9689 3519
rect 9689 3485 9723 3519
rect 9723 3485 9732 3519
rect 9680 3476 9732 3485
rect 12440 3519 12492 3528
rect 12440 3485 12449 3519
rect 12449 3485 12483 3519
rect 12483 3485 12492 3519
rect 12440 3476 12492 3485
rect 13176 3476 13228 3528
rect 15292 3519 15344 3528
rect 15292 3485 15301 3519
rect 15301 3485 15335 3519
rect 15335 3485 15344 3519
rect 15292 3476 15344 3485
rect 16304 3476 16356 3528
rect 17960 3476 18012 3528
rect 20352 3476 20404 3528
rect 22928 3544 22980 3596
rect 23020 3587 23072 3596
rect 23020 3553 23029 3587
rect 23029 3553 23063 3587
rect 23063 3553 23072 3587
rect 23020 3544 23072 3553
rect 25596 3544 25648 3596
rect 21088 3476 21140 3528
rect 23204 3476 23256 3528
rect 24584 3476 24636 3528
rect 27068 3519 27120 3528
rect 27068 3485 27077 3519
rect 27077 3485 27111 3519
rect 27111 3485 27120 3519
rect 27068 3476 27120 3485
rect 8668 3408 8720 3460
rect 9772 3408 9824 3460
rect 12624 3340 12676 3392
rect 14096 3340 14148 3392
rect 14924 3340 14976 3392
rect 22560 3340 22612 3392
rect 22652 3340 22704 3392
rect 24400 3340 24452 3392
rect 27620 3612 27672 3664
rect 27896 3612 27948 3664
rect 32680 3612 32732 3664
rect 31024 3587 31076 3596
rect 31024 3553 31033 3587
rect 31033 3553 31067 3587
rect 31067 3553 31076 3587
rect 31024 3544 31076 3553
rect 33600 3544 33652 3596
rect 34336 3680 34388 3732
rect 27896 3476 27948 3528
rect 28264 3476 28316 3528
rect 31208 3519 31260 3528
rect 29276 3408 29328 3460
rect 31208 3485 31217 3519
rect 31217 3485 31251 3519
rect 31251 3485 31260 3519
rect 31208 3476 31260 3485
rect 31668 3476 31720 3528
rect 32956 3519 33008 3528
rect 32956 3485 32965 3519
rect 32965 3485 32999 3519
rect 32999 3485 33008 3519
rect 32956 3476 33008 3485
rect 34704 3476 34756 3528
rect 31024 3340 31076 3392
rect 33416 3340 33468 3392
rect 33600 3340 33652 3392
rect 35440 3340 35492 3392
rect 37096 3383 37148 3392
rect 37096 3349 37105 3383
rect 37105 3349 37139 3383
rect 37139 3349 37148 3383
rect 37096 3340 37148 3349
rect 4246 3238 4298 3290
rect 4310 3238 4362 3290
rect 4374 3238 4426 3290
rect 4438 3238 4490 3290
rect 34966 3238 35018 3290
rect 35030 3238 35082 3290
rect 35094 3238 35146 3290
rect 35158 3238 35210 3290
rect 8024 3136 8076 3188
rect 8484 3068 8536 3120
rect 9404 3068 9456 3120
rect 11060 3068 11112 3120
rect 14188 3136 14240 3188
rect 20720 3136 20772 3188
rect 25228 3136 25280 3188
rect 25780 3136 25832 3188
rect 8024 3000 8076 3052
rect 12716 3043 12768 3052
rect 12716 3009 12725 3043
rect 12725 3009 12759 3043
rect 12759 3009 12768 3043
rect 12716 3000 12768 3009
rect 14832 3043 14884 3052
rect 14832 3009 14841 3043
rect 14841 3009 14875 3043
rect 14875 3009 14884 3043
rect 14832 3000 14884 3009
rect 16120 3043 16172 3052
rect 3148 2975 3200 2984
rect 3148 2941 3157 2975
rect 3157 2941 3191 2975
rect 3191 2941 3200 2975
rect 3148 2932 3200 2941
rect 7288 2975 7340 2984
rect 7288 2941 7297 2975
rect 7297 2941 7331 2975
rect 7331 2941 7340 2975
rect 7288 2932 7340 2941
rect 4620 2796 4672 2848
rect 8668 2932 8720 2984
rect 8852 2975 8904 2984
rect 8852 2941 8861 2975
rect 8861 2941 8895 2975
rect 8895 2941 8904 2975
rect 8852 2932 8904 2941
rect 9404 2932 9456 2984
rect 9220 2864 9272 2916
rect 9588 2864 9640 2916
rect 12348 2932 12400 2984
rect 12440 2975 12492 2984
rect 12440 2941 12449 2975
rect 12449 2941 12483 2975
rect 12483 2941 12492 2975
rect 12440 2932 12492 2941
rect 14188 2932 14240 2984
rect 14924 2975 14976 2984
rect 14924 2941 14933 2975
rect 14933 2941 14967 2975
rect 14967 2941 14976 2975
rect 14924 2932 14976 2941
rect 15292 2932 15344 2984
rect 16120 3009 16129 3043
rect 16129 3009 16163 3043
rect 16163 3009 16172 3043
rect 16120 3000 16172 3009
rect 22928 3068 22980 3120
rect 13912 2796 13964 2848
rect 15936 2796 15988 2848
rect 21088 3000 21140 3052
rect 24584 3043 24636 3052
rect 18972 2932 19024 2984
rect 19432 2932 19484 2984
rect 20352 2975 20404 2984
rect 20352 2941 20361 2975
rect 20361 2941 20395 2975
rect 20395 2941 20404 2975
rect 20352 2932 20404 2941
rect 20628 2975 20680 2984
rect 20628 2941 20637 2975
rect 20637 2941 20671 2975
rect 20671 2941 20680 2975
rect 20628 2932 20680 2941
rect 22100 2932 22152 2984
rect 22560 2975 22612 2984
rect 22560 2941 22569 2975
rect 22569 2941 22603 2975
rect 22603 2941 22612 2975
rect 22560 2932 22612 2941
rect 23112 2932 23164 2984
rect 24584 3009 24593 3043
rect 24593 3009 24627 3043
rect 24627 3009 24636 3043
rect 24584 3000 24636 3009
rect 27436 3136 27488 3188
rect 37740 3136 37792 3188
rect 29644 3068 29696 3120
rect 32588 3068 32640 3120
rect 28264 3000 28316 3052
rect 29276 3043 29328 3052
rect 29276 3009 29285 3043
rect 29285 3009 29319 3043
rect 29319 3009 29328 3043
rect 29276 3000 29328 3009
rect 29828 3043 29880 3052
rect 29828 3009 29837 3043
rect 29837 3009 29871 3043
rect 29871 3009 29880 3043
rect 29828 3000 29880 3009
rect 30196 3000 30248 3052
rect 27620 2932 27672 2984
rect 22744 2864 22796 2916
rect 23020 2907 23072 2916
rect 23020 2873 23029 2907
rect 23029 2873 23063 2907
rect 23063 2873 23072 2907
rect 23020 2864 23072 2873
rect 23388 2796 23440 2848
rect 23480 2796 23532 2848
rect 31852 2975 31904 2984
rect 29828 2864 29880 2916
rect 31852 2941 31861 2975
rect 31861 2941 31895 2975
rect 31895 2941 31904 2975
rect 31852 2932 31904 2941
rect 34520 3000 34572 3052
rect 35440 3068 35492 3120
rect 33600 2932 33652 2984
rect 33876 2932 33928 2984
rect 34428 2932 34480 2984
rect 35900 2975 35952 2984
rect 33324 2864 33376 2916
rect 35900 2941 35909 2975
rect 35909 2941 35943 2975
rect 35943 2941 35952 2975
rect 35900 2932 35952 2941
rect 33508 2796 33560 2848
rect 39028 2864 39080 2916
rect 19606 2694 19658 2746
rect 19670 2694 19722 2746
rect 19734 2694 19786 2746
rect 19798 2694 19850 2746
rect 3424 2592 3476 2644
rect 3148 2456 3200 2508
rect 7748 2456 7800 2508
rect 9220 2456 9272 2508
rect 12624 2499 12676 2508
rect 12624 2465 12633 2499
rect 12633 2465 12667 2499
rect 12667 2465 12676 2499
rect 12624 2456 12676 2465
rect 15568 2524 15620 2576
rect 19248 2524 19300 2576
rect 14096 2499 14148 2508
rect 14096 2465 14105 2499
rect 14105 2465 14139 2499
rect 14139 2465 14148 2499
rect 14096 2456 14148 2465
rect 16028 2456 16080 2508
rect 9680 2388 9732 2440
rect 12440 2388 12492 2440
rect 13176 2431 13228 2440
rect 13176 2397 13185 2431
rect 13185 2397 13219 2431
rect 13219 2397 13228 2431
rect 13176 2388 13228 2397
rect 13912 2388 13964 2440
rect 14188 2388 14240 2440
rect 23204 2524 23256 2576
rect 19708 2499 19760 2508
rect 19708 2465 19717 2499
rect 19717 2465 19751 2499
rect 19751 2465 19760 2499
rect 19708 2456 19760 2465
rect 22652 2456 22704 2508
rect 22744 2456 22796 2508
rect 24400 2592 24452 2644
rect 23388 2524 23440 2576
rect 27068 2592 27120 2644
rect 23480 2499 23532 2508
rect 23480 2465 23489 2499
rect 23489 2465 23523 2499
rect 23523 2465 23532 2499
rect 23480 2456 23532 2465
rect 26240 2524 26292 2576
rect 29828 2524 29880 2576
rect 24584 2431 24636 2440
rect 24584 2397 24593 2431
rect 24593 2397 24627 2431
rect 24627 2397 24636 2431
rect 24584 2388 24636 2397
rect 25780 2388 25832 2440
rect 27896 2499 27948 2508
rect 27896 2465 27905 2499
rect 27905 2465 27939 2499
rect 27939 2465 27948 2499
rect 27896 2456 27948 2465
rect 28908 2456 28960 2508
rect 29644 2456 29696 2508
rect 30012 2499 30064 2508
rect 30012 2465 30021 2499
rect 30021 2465 30055 2499
rect 30055 2465 30064 2499
rect 30012 2456 30064 2465
rect 30196 2388 30248 2440
rect 33232 2524 33284 2576
rect 33508 2456 33560 2508
rect 35440 2499 35492 2508
rect 35440 2465 35449 2499
rect 35449 2465 35483 2499
rect 35483 2465 35492 2499
rect 35440 2456 35492 2465
rect 33140 2431 33192 2440
rect 33140 2397 33149 2431
rect 33149 2397 33183 2431
rect 33183 2397 33192 2431
rect 33140 2388 33192 2397
rect 2412 2252 2464 2304
rect 11980 2295 12032 2304
rect 11980 2261 11989 2295
rect 11989 2261 12023 2295
rect 12023 2261 12032 2295
rect 11980 2252 12032 2261
rect 15844 2252 15896 2304
rect 23020 2252 23072 2304
rect 27436 2252 27488 2304
rect 31668 2320 31720 2372
rect 31300 2295 31352 2304
rect 31300 2261 31309 2295
rect 31309 2261 31343 2295
rect 31343 2261 31352 2295
rect 31300 2252 31352 2261
rect 33140 2252 33192 2304
rect 34428 2252 34480 2304
rect 37188 2252 37240 2304
rect 4246 2150 4298 2202
rect 4310 2150 4362 2202
rect 4374 2150 4426 2202
rect 4438 2150 4490 2202
rect 34966 2150 35018 2202
rect 35030 2150 35082 2202
rect 35094 2150 35146 2202
rect 35158 2150 35210 2202
rect 24584 2048 24636 2100
rect 31852 2048 31904 2100
rect 29736 1096 29788 1148
rect 35164 1096 35216 1148
<< metal2 >>
rect 754 40200 810 41000
rect 2778 40200 2834 41000
rect 4618 40200 4674 41000
rect 6642 40200 6698 41000
rect 8482 40200 8538 41000
rect 10506 40200 10562 41000
rect 12346 40200 12402 41000
rect 14370 40200 14426 41000
rect 16210 40200 16266 41000
rect 18234 40200 18290 41000
rect 20074 40200 20130 41000
rect 22098 40200 22154 41000
rect 23938 40200 23994 41000
rect 25962 40200 26018 41000
rect 27802 40200 27858 41000
rect 29826 40200 29882 41000
rect 31666 40200 31722 41000
rect 33690 40200 33746 41000
rect 35530 40200 35586 41000
rect 37554 40200 37610 41000
rect 39394 40200 39450 41000
rect 768 36038 796 40200
rect 2792 38026 2820 40200
rect 4220 38108 4516 38128
rect 4276 38106 4300 38108
rect 4356 38106 4380 38108
rect 4436 38106 4460 38108
rect 4298 38054 4300 38106
rect 4362 38054 4374 38106
rect 4436 38054 4438 38106
rect 4276 38052 4300 38054
rect 4356 38052 4380 38054
rect 4436 38052 4460 38054
rect 4220 38032 4516 38052
rect 2792 37998 3004 38026
rect 4632 38010 4660 40200
rect 6000 38480 6052 38486
rect 6000 38422 6052 38428
rect 2778 37904 2834 37913
rect 2778 37839 2834 37848
rect 2792 36922 2820 37839
rect 2976 36922 3004 37998
rect 4620 38004 4672 38010
rect 4620 37946 4672 37952
rect 3608 37868 3660 37874
rect 3608 37810 3660 37816
rect 5632 37868 5684 37874
rect 5632 37810 5684 37816
rect 2780 36916 2832 36922
rect 2780 36858 2832 36864
rect 2964 36916 3016 36922
rect 2964 36858 3016 36864
rect 3620 36786 3648 37810
rect 3976 37800 4028 37806
rect 3976 37742 4028 37748
rect 3608 36780 3660 36786
rect 3608 36722 3660 36728
rect 1952 36712 2004 36718
rect 1952 36654 2004 36660
rect 20 36032 72 36038
rect 20 35974 72 35980
rect 756 36032 808 36038
rect 756 35974 808 35980
rect 32 30841 60 35974
rect 1860 33992 1912 33998
rect 1860 33934 1912 33940
rect 1584 33584 1636 33590
rect 1584 33526 1636 33532
rect 1400 31884 1452 31890
rect 1400 31826 1452 31832
rect 18 30832 74 30841
rect 18 30767 74 30776
rect 1412 29714 1440 31826
rect 1596 31278 1624 33526
rect 1872 33046 1900 33934
rect 1860 33040 1912 33046
rect 1860 32982 1912 32988
rect 1860 32292 1912 32298
rect 1860 32234 1912 32240
rect 1676 31816 1728 31822
rect 1676 31758 1728 31764
rect 1688 31482 1716 31758
rect 1676 31476 1728 31482
rect 1676 31418 1728 31424
rect 1584 31272 1636 31278
rect 1584 31214 1636 31220
rect 1768 30252 1820 30258
rect 1768 30194 1820 30200
rect 1492 30116 1544 30122
rect 1492 30058 1544 30064
rect 1400 29708 1452 29714
rect 1400 29650 1452 29656
rect 1504 29306 1532 30058
rect 1676 29640 1728 29646
rect 1676 29582 1728 29588
rect 1688 29306 1716 29582
rect 1492 29300 1544 29306
rect 1492 29242 1544 29248
rect 1676 29300 1728 29306
rect 1676 29242 1728 29248
rect 1780 29102 1808 30194
rect 1872 29170 1900 32234
rect 1860 29164 1912 29170
rect 1860 29106 1912 29112
rect 1768 29096 1820 29102
rect 1768 29038 1820 29044
rect 1400 28552 1452 28558
rect 1400 28494 1452 28500
rect 1412 27402 1440 28494
rect 1400 27396 1452 27402
rect 1400 27338 1452 27344
rect 1412 26926 1440 27338
rect 1400 26920 1452 26926
rect 1400 26862 1452 26868
rect 1412 25378 1440 26862
rect 1964 26364 1992 36654
rect 3620 35154 3648 36722
rect 3608 35148 3660 35154
rect 3608 35090 3660 35096
rect 3332 34400 3384 34406
rect 3332 34342 3384 34348
rect 2688 34060 2740 34066
rect 2688 34002 2740 34008
rect 2136 33448 2188 33454
rect 2136 33390 2188 33396
rect 2044 33312 2096 33318
rect 2044 33254 2096 33260
rect 2056 29034 2084 33254
rect 2148 30870 2176 33390
rect 2700 32026 2728 34002
rect 3240 33856 3292 33862
rect 3240 33798 3292 33804
rect 3252 33522 3280 33798
rect 3240 33516 3292 33522
rect 3240 33458 3292 33464
rect 2780 33380 2832 33386
rect 2780 33322 2832 33328
rect 2872 33380 2924 33386
rect 2872 33322 2924 33328
rect 2792 32858 2820 33322
rect 2884 32978 2912 33322
rect 3252 32978 3280 33458
rect 3344 33454 3372 34342
rect 3620 34066 3648 35090
rect 3608 34060 3660 34066
rect 3608 34002 3660 34008
rect 3332 33448 3384 33454
rect 3332 33390 3384 33396
rect 2872 32972 2924 32978
rect 2872 32914 2924 32920
rect 3148 32972 3200 32978
rect 3148 32914 3200 32920
rect 3240 32972 3292 32978
rect 3240 32914 3292 32920
rect 2792 32830 2912 32858
rect 2780 32360 2832 32366
rect 2780 32302 2832 32308
rect 2688 32020 2740 32026
rect 2688 31962 2740 31968
rect 2792 31686 2820 32302
rect 2504 31680 2556 31686
rect 2504 31622 2556 31628
rect 2780 31680 2832 31686
rect 2780 31622 2832 31628
rect 2516 31278 2544 31622
rect 2884 31346 2912 32830
rect 3160 32434 3188 32914
rect 3148 32428 3200 32434
rect 3148 32370 3200 32376
rect 3056 32360 3108 32366
rect 3056 32302 3108 32308
rect 2962 32192 3018 32201
rect 2962 32127 3018 32136
rect 2872 31340 2924 31346
rect 2872 31282 2924 31288
rect 2504 31272 2556 31278
rect 2504 31214 2556 31220
rect 2780 31272 2832 31278
rect 2780 31214 2832 31220
rect 2136 30864 2188 30870
rect 2136 30806 2188 30812
rect 2792 30190 2820 31214
rect 2976 30274 3004 32127
rect 3068 31278 3096 32302
rect 3344 32230 3372 33390
rect 3608 33380 3660 33386
rect 3608 33322 3660 33328
rect 3620 32774 3648 33322
rect 3608 32768 3660 32774
rect 3608 32710 3660 32716
rect 3424 32496 3476 32502
rect 3424 32438 3476 32444
rect 3332 32224 3384 32230
rect 3332 32166 3384 32172
rect 3344 31278 3372 32166
rect 3056 31272 3108 31278
rect 3056 31214 3108 31220
rect 3332 31272 3384 31278
rect 3332 31214 3384 31220
rect 3332 30796 3384 30802
rect 3332 30738 3384 30744
rect 2976 30246 3096 30274
rect 2780 30184 2832 30190
rect 2780 30126 2832 30132
rect 2964 30184 3016 30190
rect 2964 30126 3016 30132
rect 2792 29850 2820 30126
rect 2780 29844 2832 29850
rect 2780 29786 2832 29792
rect 2792 29034 2820 29786
rect 2872 29708 2924 29714
rect 2872 29650 2924 29656
rect 2044 29028 2096 29034
rect 2044 28970 2096 28976
rect 2780 29028 2832 29034
rect 2780 28970 2832 28976
rect 2056 27538 2084 28970
rect 2884 28914 2912 29650
rect 2792 28886 2912 28914
rect 2792 28150 2820 28886
rect 2872 28756 2924 28762
rect 2872 28698 2924 28704
rect 2780 28144 2832 28150
rect 2780 28086 2832 28092
rect 2884 28082 2912 28698
rect 2976 28218 3004 30126
rect 2964 28212 3016 28218
rect 2964 28154 3016 28160
rect 2872 28076 2924 28082
rect 2872 28018 2924 28024
rect 2596 27872 2648 27878
rect 2596 27814 2648 27820
rect 2608 27538 2636 27814
rect 2044 27532 2096 27538
rect 2044 27474 2096 27480
rect 2504 27532 2556 27538
rect 2504 27474 2556 27480
rect 2596 27532 2648 27538
rect 2596 27474 2648 27480
rect 2044 27328 2096 27334
rect 2044 27270 2096 27276
rect 2056 26518 2084 27270
rect 2516 26790 2544 27474
rect 2780 27328 2832 27334
rect 2780 27270 2832 27276
rect 2792 26994 2820 27270
rect 2780 26988 2832 26994
rect 2780 26930 2832 26936
rect 2596 26920 2648 26926
rect 2596 26862 2648 26868
rect 2504 26784 2556 26790
rect 2504 26726 2556 26732
rect 2044 26512 2096 26518
rect 2044 26454 2096 26460
rect 1964 26336 2084 26364
rect 1768 25832 1820 25838
rect 1768 25774 1820 25780
rect 1676 25696 1728 25702
rect 1676 25638 1728 25644
rect 1412 25362 1532 25378
rect 1688 25362 1716 25638
rect 1412 25356 1544 25362
rect 1412 25350 1492 25356
rect 1492 25298 1544 25304
rect 1676 25356 1728 25362
rect 1676 25298 1728 25304
rect 1504 23526 1532 25298
rect 1780 24274 1808 25774
rect 1860 24404 1912 24410
rect 1860 24346 1912 24352
rect 1768 24268 1820 24274
rect 1768 24210 1820 24216
rect 1492 23520 1544 23526
rect 1492 23462 1544 23468
rect 1504 23186 1532 23462
rect 1492 23180 1544 23186
rect 1492 23122 1544 23128
rect 1504 21486 1532 23122
rect 1780 21554 1808 24210
rect 1872 23186 1900 24346
rect 1860 23180 1912 23186
rect 1860 23122 1912 23128
rect 1860 21956 1912 21962
rect 1860 21898 1912 21904
rect 1768 21548 1820 21554
rect 1768 21490 1820 21496
rect 1492 21480 1544 21486
rect 1492 21422 1544 21428
rect 1768 21072 1820 21078
rect 1768 21014 1820 21020
rect 1676 20936 1728 20942
rect 1676 20878 1728 20884
rect 1400 20392 1452 20398
rect 1400 20334 1452 20340
rect 1412 19174 1440 20334
rect 1688 19310 1716 20878
rect 1780 19310 1808 21014
rect 1872 21010 1900 21898
rect 1952 21480 2004 21486
rect 1952 21422 2004 21428
rect 1964 21146 1992 21422
rect 1952 21140 2004 21146
rect 1952 21082 2004 21088
rect 1860 21004 1912 21010
rect 1860 20946 1912 20952
rect 2056 20482 2084 26336
rect 2412 25900 2464 25906
rect 2412 25842 2464 25848
rect 2320 25832 2372 25838
rect 2318 25800 2320 25809
rect 2372 25800 2374 25809
rect 2318 25735 2374 25744
rect 2424 24886 2452 25842
rect 2412 24880 2464 24886
rect 2412 24822 2464 24828
rect 2320 22636 2372 22642
rect 2320 22578 2372 22584
rect 2332 22234 2360 22578
rect 2320 22228 2372 22234
rect 2320 22170 2372 22176
rect 2332 22098 2360 22170
rect 2320 22092 2372 22098
rect 2320 22034 2372 22040
rect 2516 21078 2544 26726
rect 2608 26450 2636 26862
rect 2870 26480 2926 26489
rect 2596 26444 2648 26450
rect 2596 26386 2648 26392
rect 2688 26444 2740 26450
rect 2870 26415 2926 26424
rect 2688 26386 2740 26392
rect 2700 26042 2728 26386
rect 2780 26308 2832 26314
rect 2780 26250 2832 26256
rect 2688 26036 2740 26042
rect 2688 25978 2740 25984
rect 2792 25158 2820 26250
rect 2780 25152 2832 25158
rect 2780 25094 2832 25100
rect 2792 24750 2820 25094
rect 2780 24744 2832 24750
rect 2780 24686 2832 24692
rect 2596 24268 2648 24274
rect 2596 24210 2648 24216
rect 2608 23798 2636 24210
rect 2596 23792 2648 23798
rect 2596 23734 2648 23740
rect 2778 23488 2834 23497
rect 2778 23423 2834 23432
rect 2688 22568 2740 22574
rect 2688 22510 2740 22516
rect 2700 22098 2728 22510
rect 2688 22092 2740 22098
rect 2688 22034 2740 22040
rect 2504 21072 2556 21078
rect 2504 21014 2556 21020
rect 1964 20454 2084 20482
rect 1676 19304 1728 19310
rect 1676 19246 1728 19252
rect 1768 19304 1820 19310
rect 1768 19246 1820 19252
rect 1400 19168 1452 19174
rect 1400 19110 1452 19116
rect 1412 18834 1440 19110
rect 1400 18828 1452 18834
rect 1400 18770 1452 18776
rect 1412 17746 1440 18770
rect 1964 18737 1992 20454
rect 2044 20392 2096 20398
rect 2044 20334 2096 20340
rect 2056 19514 2084 20334
rect 2044 19508 2096 19514
rect 2044 19450 2096 19456
rect 2792 18970 2820 23423
rect 2780 18964 2832 18970
rect 2780 18906 2832 18912
rect 1950 18728 2006 18737
rect 1950 18663 2006 18672
rect 1950 17776 2006 17785
rect 1400 17740 1452 17746
rect 1950 17711 2006 17720
rect 1400 17682 1452 17688
rect 1412 17202 1440 17682
rect 1400 17196 1452 17202
rect 1400 17138 1452 17144
rect 1412 15570 1440 17138
rect 1964 16794 1992 17711
rect 2884 17338 2912 26415
rect 2964 25832 3016 25838
rect 2964 25774 3016 25780
rect 2976 24750 3004 25774
rect 2964 24744 3016 24750
rect 2964 24686 3016 24692
rect 2976 23730 3004 24686
rect 3068 24154 3096 30246
rect 3240 30184 3292 30190
rect 3240 30126 3292 30132
rect 3148 29776 3200 29782
rect 3148 29718 3200 29724
rect 3160 29170 3188 29718
rect 3148 29164 3200 29170
rect 3148 29106 3200 29112
rect 3252 28762 3280 30126
rect 3344 29170 3372 30738
rect 3436 30190 3464 32438
rect 3516 31680 3568 31686
rect 3516 31622 3568 31628
rect 3528 30802 3556 31622
rect 3516 30796 3568 30802
rect 3516 30738 3568 30744
rect 3424 30184 3476 30190
rect 3424 30126 3476 30132
rect 3516 30184 3568 30190
rect 3516 30126 3568 30132
rect 3436 29782 3464 30126
rect 3528 29850 3556 30126
rect 3516 29844 3568 29850
rect 3516 29786 3568 29792
rect 3424 29776 3476 29782
rect 3424 29718 3476 29724
rect 3332 29164 3384 29170
rect 3332 29106 3384 29112
rect 3528 29102 3556 29786
rect 3516 29096 3568 29102
rect 3516 29038 3568 29044
rect 3514 28792 3570 28801
rect 3240 28756 3292 28762
rect 3514 28727 3570 28736
rect 3240 28698 3292 28704
rect 3424 28008 3476 28014
rect 3424 27950 3476 27956
rect 3436 27538 3464 27950
rect 3424 27532 3476 27538
rect 3424 27474 3476 27480
rect 3148 26444 3200 26450
rect 3148 26386 3200 26392
rect 3160 25702 3188 26386
rect 3148 25696 3200 25702
rect 3148 25638 3200 25644
rect 3240 24744 3292 24750
rect 3240 24686 3292 24692
rect 3068 24126 3188 24154
rect 2964 23724 3016 23730
rect 2964 23666 3016 23672
rect 2976 22642 3004 23666
rect 2964 22636 3016 22642
rect 2964 22578 3016 22584
rect 2964 22432 3016 22438
rect 2964 22374 3016 22380
rect 2976 22098 3004 22374
rect 2964 22092 3016 22098
rect 2964 22034 3016 22040
rect 2964 21412 3016 21418
rect 2964 21354 3016 21360
rect 2976 21010 3004 21354
rect 2964 21004 3016 21010
rect 2964 20946 3016 20952
rect 2976 20602 3004 20946
rect 2964 20596 3016 20602
rect 2964 20538 3016 20544
rect 2976 19990 3004 20538
rect 2964 19984 3016 19990
rect 2964 19926 3016 19932
rect 3056 19304 3108 19310
rect 3056 19246 3108 19252
rect 3068 18290 3096 19246
rect 3056 18284 3108 18290
rect 3056 18226 3108 18232
rect 3160 17814 3188 24126
rect 3252 23662 3280 24686
rect 3332 24268 3384 24274
rect 3332 24210 3384 24216
rect 3240 23656 3292 23662
rect 3240 23598 3292 23604
rect 3252 22574 3280 23598
rect 3240 22568 3292 22574
rect 3240 22510 3292 22516
rect 3252 22234 3280 22510
rect 3240 22228 3292 22234
rect 3240 22170 3292 22176
rect 3344 21894 3372 24210
rect 3424 24064 3476 24070
rect 3424 24006 3476 24012
rect 3436 23186 3464 24006
rect 3424 23180 3476 23186
rect 3424 23122 3476 23128
rect 3436 22574 3464 23122
rect 3424 22568 3476 22574
rect 3424 22510 3476 22516
rect 3332 21888 3384 21894
rect 3332 21830 3384 21836
rect 3344 21690 3372 21830
rect 3332 21684 3384 21690
rect 3332 21626 3384 21632
rect 3332 21004 3384 21010
rect 3332 20946 3384 20952
rect 3344 19922 3372 20946
rect 3422 20768 3478 20777
rect 3422 20703 3478 20712
rect 3332 19916 3384 19922
rect 3332 19858 3384 19864
rect 3148 17808 3200 17814
rect 3148 17750 3200 17756
rect 2872 17332 2924 17338
rect 2872 17274 2924 17280
rect 2504 17128 2556 17134
rect 2504 17070 2556 17076
rect 2516 16794 2544 17070
rect 1952 16788 2004 16794
rect 1952 16730 2004 16736
rect 2504 16788 2556 16794
rect 2504 16730 2556 16736
rect 1768 16652 1820 16658
rect 1768 16594 1820 16600
rect 1400 15564 1452 15570
rect 1400 15506 1452 15512
rect 1412 14958 1440 15506
rect 1400 14952 1452 14958
rect 1400 14894 1452 14900
rect 1674 14512 1730 14521
rect 1674 14447 1676 14456
rect 1728 14447 1730 14456
rect 1676 14418 1728 14424
rect 1400 14408 1452 14414
rect 1400 14350 1452 14356
rect 1412 13326 1440 14350
rect 1400 13320 1452 13326
rect 1400 13262 1452 13268
rect 1676 13320 1728 13326
rect 1676 13262 1728 13268
rect 1412 12850 1440 13262
rect 1688 12986 1716 13262
rect 1676 12980 1728 12986
rect 1676 12922 1728 12928
rect 1400 12844 1452 12850
rect 1400 12786 1452 12792
rect 1676 11212 1728 11218
rect 1676 11154 1728 11160
rect 1688 10606 1716 11154
rect 1400 10600 1452 10606
rect 1400 10542 1452 10548
rect 1676 10600 1728 10606
rect 1676 10542 1728 10548
rect 1412 10062 1440 10542
rect 1688 10266 1716 10542
rect 1676 10260 1728 10266
rect 1676 10202 1728 10208
rect 1400 10056 1452 10062
rect 1400 9998 1452 10004
rect 1780 8906 1808 16594
rect 2516 16114 2544 16730
rect 2504 16108 2556 16114
rect 2504 16050 2556 16056
rect 2516 15570 2544 16050
rect 2504 15564 2556 15570
rect 2504 15506 2556 15512
rect 2688 15564 2740 15570
rect 2688 15506 2740 15512
rect 2700 14958 2728 15506
rect 2872 15360 2924 15366
rect 2872 15302 2924 15308
rect 1952 14952 2004 14958
rect 1952 14894 2004 14900
rect 2688 14952 2740 14958
rect 2688 14894 2740 14900
rect 1964 14618 1992 14894
rect 1952 14612 2004 14618
rect 1952 14554 2004 14560
rect 2688 13864 2740 13870
rect 2688 13806 2740 13812
rect 1860 12844 1912 12850
rect 1860 12786 1912 12792
rect 1872 12306 1900 12786
rect 1860 12300 1912 12306
rect 1860 12242 1912 12248
rect 2136 12232 2188 12238
rect 2136 12174 2188 12180
rect 2700 12186 2728 13806
rect 2148 11898 2176 12174
rect 2700 12158 2820 12186
rect 2792 12102 2820 12158
rect 2780 12096 2832 12102
rect 2780 12038 2832 12044
rect 2136 11892 2188 11898
rect 2136 11834 2188 11840
rect 2688 11688 2740 11694
rect 2688 11630 2740 11636
rect 2596 11076 2648 11082
rect 2596 11018 2648 11024
rect 2608 9042 2636 11018
rect 2700 10810 2728 11630
rect 2780 11552 2832 11558
rect 2780 11494 2832 11500
rect 2792 11218 2820 11494
rect 2780 11212 2832 11218
rect 2780 11154 2832 11160
rect 2884 11200 2912 15302
rect 3240 12776 3292 12782
rect 3240 12718 3292 12724
rect 3252 12442 3280 12718
rect 3240 12436 3292 12442
rect 3240 12378 3292 12384
rect 3054 12064 3110 12073
rect 3054 11999 3110 12008
rect 2964 11212 3016 11218
rect 2884 11172 2964 11200
rect 2688 10804 2740 10810
rect 2688 10746 2740 10752
rect 2700 9586 2728 10746
rect 2884 10130 2912 11172
rect 2964 11154 3016 11160
rect 2872 10124 2924 10130
rect 2872 10066 2924 10072
rect 2964 9920 3016 9926
rect 2964 9862 3016 9868
rect 2688 9580 2740 9586
rect 2688 9522 2740 9528
rect 2976 9518 3004 9862
rect 2964 9512 3016 9518
rect 2964 9454 3016 9460
rect 2872 9172 2924 9178
rect 2872 9114 2924 9120
rect 2780 9104 2832 9110
rect 2780 9046 2832 9052
rect 2596 9036 2648 9042
rect 2424 8996 2596 9024
rect 1860 8968 1912 8974
rect 1860 8910 1912 8916
rect 1768 8900 1820 8906
rect 1768 8842 1820 8848
rect 1872 7410 1900 8910
rect 1860 7404 1912 7410
rect 1860 7346 1912 7352
rect 1582 7304 1638 7313
rect 1582 7239 1584 7248
rect 1636 7239 1638 7248
rect 1768 7268 1820 7274
rect 1584 7210 1636 7216
rect 1768 7210 1820 7216
rect 1780 3534 1808 7210
rect 2424 6866 2452 8996
rect 2596 8978 2648 8984
rect 2792 7342 2820 9046
rect 2884 7954 2912 9114
rect 2976 9058 3004 9454
rect 3068 9178 3096 11999
rect 3056 9172 3108 9178
rect 3056 9114 3108 9120
rect 2976 9030 3096 9058
rect 2964 8968 3016 8974
rect 2964 8910 3016 8916
rect 2872 7948 2924 7954
rect 2872 7890 2924 7896
rect 2976 7546 3004 8910
rect 3068 7886 3096 9030
rect 3332 9036 3384 9042
rect 3332 8978 3384 8984
rect 3344 8566 3372 8978
rect 3332 8560 3384 8566
rect 3332 8502 3384 8508
rect 3240 8424 3292 8430
rect 3240 8366 3292 8372
rect 3252 8090 3280 8366
rect 3436 8362 3464 20703
rect 3528 19938 3556 28727
rect 3620 25974 3648 32710
rect 3884 31884 3936 31890
rect 3884 31826 3936 31832
rect 3896 30054 3924 31826
rect 3884 30048 3936 30054
rect 3884 29990 3936 29996
rect 3896 27538 3924 29990
rect 3988 29073 4016 37742
rect 5644 37262 5672 37810
rect 5632 37256 5684 37262
rect 5632 37198 5684 37204
rect 6012 37126 6040 38422
rect 6656 37874 6684 40200
rect 8496 38570 8524 40200
rect 8496 38542 8708 38570
rect 10520 38554 10548 40200
rect 8680 38486 8708 38542
rect 10508 38548 10560 38554
rect 10508 38490 10560 38496
rect 8668 38480 8720 38486
rect 8668 38422 8720 38428
rect 9588 38480 9640 38486
rect 9588 38422 9640 38428
rect 8300 38412 8352 38418
rect 8300 38354 8352 38360
rect 6644 37868 6696 37874
rect 6644 37810 6696 37816
rect 8312 37466 8340 38354
rect 8668 38344 8720 38350
rect 8668 38286 8720 38292
rect 9312 38344 9364 38350
rect 9312 38286 9364 38292
rect 8392 37800 8444 37806
rect 8392 37742 8444 37748
rect 7656 37460 7708 37466
rect 7656 37402 7708 37408
rect 8300 37460 8352 37466
rect 8300 37402 8352 37408
rect 4804 37120 4856 37126
rect 4804 37062 4856 37068
rect 6000 37120 6052 37126
rect 6000 37062 6052 37068
rect 7196 37120 7248 37126
rect 7196 37062 7248 37068
rect 4220 37020 4516 37040
rect 4276 37018 4300 37020
rect 4356 37018 4380 37020
rect 4436 37018 4460 37020
rect 4298 36966 4300 37018
rect 4362 36966 4374 37018
rect 4436 36966 4438 37018
rect 4276 36964 4300 36966
rect 4356 36964 4380 36966
rect 4436 36964 4460 36966
rect 4220 36944 4516 36964
rect 4816 36786 4844 37062
rect 4804 36780 4856 36786
rect 4804 36722 4856 36728
rect 5356 36712 5408 36718
rect 5356 36654 5408 36660
rect 5368 36310 5396 36654
rect 5356 36304 5408 36310
rect 5356 36246 5408 36252
rect 4804 36236 4856 36242
rect 4804 36178 4856 36184
rect 4712 36168 4764 36174
rect 4712 36110 4764 36116
rect 4620 36100 4672 36106
rect 4620 36042 4672 36048
rect 4220 35932 4516 35952
rect 4276 35930 4300 35932
rect 4356 35930 4380 35932
rect 4436 35930 4460 35932
rect 4298 35878 4300 35930
rect 4362 35878 4374 35930
rect 4436 35878 4438 35930
rect 4276 35876 4300 35878
rect 4356 35876 4380 35878
rect 4436 35876 4460 35878
rect 4220 35856 4516 35876
rect 4068 35284 4120 35290
rect 4068 35226 4120 35232
rect 4080 34921 4108 35226
rect 4632 35154 4660 36042
rect 4724 35766 4752 36110
rect 4712 35760 4764 35766
rect 4712 35702 4764 35708
rect 4816 35698 4844 36178
rect 5080 36168 5132 36174
rect 5080 36110 5132 36116
rect 4804 35692 4856 35698
rect 4804 35634 4856 35640
rect 4620 35148 4672 35154
rect 4620 35090 4672 35096
rect 4816 35086 4844 35634
rect 5092 35562 5120 36110
rect 6012 36106 6040 37062
rect 6460 36780 6512 36786
rect 6460 36722 6512 36728
rect 6472 36174 6500 36722
rect 7208 36718 7236 37062
rect 7288 36780 7340 36786
rect 7288 36722 7340 36728
rect 6920 36712 6972 36718
rect 6920 36654 6972 36660
rect 7196 36712 7248 36718
rect 7196 36654 7248 36660
rect 6644 36236 6696 36242
rect 6644 36178 6696 36184
rect 6460 36168 6512 36174
rect 6460 36110 6512 36116
rect 6000 36100 6052 36106
rect 6000 36042 6052 36048
rect 6092 35624 6144 35630
rect 6092 35566 6144 35572
rect 5080 35556 5132 35562
rect 5080 35498 5132 35504
rect 4804 35080 4856 35086
rect 4804 35022 4856 35028
rect 4066 34912 4122 34921
rect 4066 34847 4122 34856
rect 4220 34844 4516 34864
rect 4276 34842 4300 34844
rect 4356 34842 4380 34844
rect 4436 34842 4460 34844
rect 4298 34790 4300 34842
rect 4362 34790 4374 34842
rect 4436 34790 4438 34842
rect 4276 34788 4300 34790
rect 4356 34788 4380 34790
rect 4436 34788 4460 34790
rect 4220 34768 4516 34788
rect 4816 34542 4844 35022
rect 5092 34678 5120 35498
rect 5080 34672 5132 34678
rect 5080 34614 5132 34620
rect 5264 34672 5316 34678
rect 5264 34614 5316 34620
rect 4712 34536 4764 34542
rect 4712 34478 4764 34484
rect 4804 34536 4856 34542
rect 4804 34478 4856 34484
rect 4220 33756 4516 33776
rect 4276 33754 4300 33756
rect 4356 33754 4380 33756
rect 4436 33754 4460 33756
rect 4298 33702 4300 33754
rect 4362 33702 4374 33754
rect 4436 33702 4438 33754
rect 4276 33700 4300 33702
rect 4356 33700 4380 33702
rect 4436 33700 4460 33702
rect 4220 33680 4516 33700
rect 4724 33538 4752 34478
rect 4724 33510 4844 33538
rect 4620 33448 4672 33454
rect 4620 33390 4672 33396
rect 4220 32668 4516 32688
rect 4276 32666 4300 32668
rect 4356 32666 4380 32668
rect 4436 32666 4460 32668
rect 4298 32614 4300 32666
rect 4362 32614 4374 32666
rect 4436 32614 4438 32666
rect 4276 32612 4300 32614
rect 4356 32612 4380 32614
rect 4436 32612 4460 32614
rect 4220 32592 4516 32612
rect 4632 31958 4660 33390
rect 4816 33114 4844 33510
rect 5080 33516 5132 33522
rect 5080 33458 5132 33464
rect 4896 33380 4948 33386
rect 4896 33322 4948 33328
rect 4804 33108 4856 33114
rect 4804 33050 4856 33056
rect 4908 32910 4936 33322
rect 5092 33046 5120 33458
rect 5276 33454 5304 34614
rect 5448 33992 5500 33998
rect 6104 33980 6132 35566
rect 6184 35556 6236 35562
rect 6184 35498 6236 35504
rect 6196 35154 6224 35498
rect 6184 35148 6236 35154
rect 6184 35090 6236 35096
rect 6276 35148 6328 35154
rect 6276 35090 6328 35096
rect 6288 34610 6316 35090
rect 6472 34950 6500 36110
rect 6656 35698 6684 36178
rect 6736 36100 6788 36106
rect 6736 36042 6788 36048
rect 6644 35692 6696 35698
rect 6644 35634 6696 35640
rect 6748 35630 6776 36042
rect 6932 36038 6960 36654
rect 7208 36378 7236 36654
rect 7196 36372 7248 36378
rect 7196 36314 7248 36320
rect 7300 36258 7328 36722
rect 7380 36576 7432 36582
rect 7380 36518 7432 36524
rect 7208 36230 7328 36258
rect 7392 36242 7420 36518
rect 7668 36310 7696 37402
rect 8116 37324 8168 37330
rect 8116 37266 8168 37272
rect 8128 36786 8156 37266
rect 8404 37262 8432 37742
rect 8680 37330 8708 38286
rect 9220 37800 9272 37806
rect 9324 37754 9352 38286
rect 9272 37748 9352 37754
rect 9220 37742 9352 37748
rect 9232 37726 9352 37742
rect 8668 37324 8720 37330
rect 8668 37266 8720 37272
rect 8392 37256 8444 37262
rect 8392 37198 8444 37204
rect 8116 36780 8168 36786
rect 8116 36722 8168 36728
rect 7840 36712 7892 36718
rect 7840 36654 7892 36660
rect 7656 36304 7708 36310
rect 7656 36246 7708 36252
rect 7380 36236 7432 36242
rect 7208 36038 7236 36230
rect 7380 36178 7432 36184
rect 6920 36032 6972 36038
rect 6920 35974 6972 35980
rect 7196 36032 7248 36038
rect 7196 35974 7248 35980
rect 6736 35624 6788 35630
rect 6736 35566 6788 35572
rect 6644 35488 6696 35494
rect 6644 35430 6696 35436
rect 6460 34944 6512 34950
rect 6460 34886 6512 34892
rect 6276 34604 6328 34610
rect 6276 34546 6328 34552
rect 6184 33992 6236 33998
rect 6104 33952 6184 33980
rect 5448 33934 5500 33940
rect 6184 33934 6236 33940
rect 5460 33658 5488 33934
rect 5632 33856 5684 33862
rect 5632 33798 5684 33804
rect 5448 33652 5500 33658
rect 5448 33594 5500 33600
rect 5264 33448 5316 33454
rect 5264 33390 5316 33396
rect 5172 33108 5224 33114
rect 5172 33050 5224 33056
rect 5080 33040 5132 33046
rect 5080 32982 5132 32988
rect 4896 32904 4948 32910
rect 4896 32846 4948 32852
rect 4712 32224 4764 32230
rect 4712 32166 4764 32172
rect 4620 31952 4672 31958
rect 4620 31894 4672 31900
rect 4724 31890 4752 32166
rect 4712 31884 4764 31890
rect 4712 31826 4764 31832
rect 4908 31872 4936 32846
rect 5092 32366 5120 32982
rect 5080 32360 5132 32366
rect 5080 32302 5132 32308
rect 5092 32026 5120 32302
rect 5080 32020 5132 32026
rect 5080 31962 5132 31968
rect 5184 31890 5212 33050
rect 5644 33046 5672 33798
rect 5632 33040 5684 33046
rect 5632 32982 5684 32988
rect 5264 32972 5316 32978
rect 5264 32914 5316 32920
rect 5276 32298 5304 32914
rect 5644 32434 5672 32982
rect 6196 32570 6224 33934
rect 6472 33046 6500 34886
rect 6460 33040 6512 33046
rect 6460 32982 6512 32988
rect 6276 32972 6328 32978
rect 6276 32914 6328 32920
rect 6184 32564 6236 32570
rect 6184 32506 6236 32512
rect 5632 32428 5684 32434
rect 5632 32370 5684 32376
rect 5540 32360 5592 32366
rect 5540 32302 5592 32308
rect 5264 32292 5316 32298
rect 5264 32234 5316 32240
rect 5276 31890 5304 32234
rect 4988 31884 5040 31890
rect 4908 31844 4988 31872
rect 4804 31748 4856 31754
rect 4804 31690 4856 31696
rect 4220 31580 4516 31600
rect 4276 31578 4300 31580
rect 4356 31578 4380 31580
rect 4436 31578 4460 31580
rect 4298 31526 4300 31578
rect 4362 31526 4374 31578
rect 4436 31526 4438 31578
rect 4276 31524 4300 31526
rect 4356 31524 4380 31526
rect 4436 31524 4460 31526
rect 4220 31504 4516 31524
rect 4816 31482 4844 31690
rect 4804 31476 4856 31482
rect 4804 31418 4856 31424
rect 4908 31328 4936 31844
rect 4988 31826 5040 31832
rect 5172 31884 5224 31890
rect 5172 31826 5224 31832
rect 5264 31884 5316 31890
rect 5264 31826 5316 31832
rect 5448 31816 5500 31822
rect 5448 31758 5500 31764
rect 4816 31300 4936 31328
rect 4068 31272 4120 31278
rect 4068 31214 4120 31220
rect 4080 30326 4108 31214
rect 4816 31210 4844 31300
rect 4988 31272 5040 31278
rect 4988 31214 5040 31220
rect 5356 31272 5408 31278
rect 5356 31214 5408 31220
rect 4804 31204 4856 31210
rect 4804 31146 4856 31152
rect 4712 30728 4764 30734
rect 4712 30670 4764 30676
rect 4220 30492 4516 30512
rect 4276 30490 4300 30492
rect 4356 30490 4380 30492
rect 4436 30490 4460 30492
rect 4298 30438 4300 30490
rect 4362 30438 4374 30490
rect 4436 30438 4438 30490
rect 4276 30436 4300 30438
rect 4356 30436 4380 30438
rect 4436 30436 4460 30438
rect 4220 30416 4516 30436
rect 4068 30320 4120 30326
rect 4068 30262 4120 30268
rect 4724 30122 4752 30670
rect 4712 30116 4764 30122
rect 4712 30058 4764 30064
rect 4816 29578 4844 31146
rect 4896 31136 4948 31142
rect 4896 31078 4948 31084
rect 4908 30802 4936 31078
rect 4896 30796 4948 30802
rect 4896 30738 4948 30744
rect 5000 30190 5028 31214
rect 5368 30190 5396 31214
rect 5460 31142 5488 31758
rect 5448 31136 5500 31142
rect 5448 31078 5500 31084
rect 4988 30184 5040 30190
rect 4988 30126 5040 30132
rect 5356 30184 5408 30190
rect 5356 30126 5408 30132
rect 4804 29572 4856 29578
rect 4804 29514 4856 29520
rect 4620 29504 4672 29510
rect 4620 29446 4672 29452
rect 4220 29404 4516 29424
rect 4276 29402 4300 29404
rect 4356 29402 4380 29404
rect 4436 29402 4460 29404
rect 4298 29350 4300 29402
rect 4362 29350 4374 29402
rect 4436 29350 4438 29402
rect 4276 29348 4300 29350
rect 4356 29348 4380 29350
rect 4436 29348 4460 29350
rect 4220 29328 4516 29348
rect 3974 29064 4030 29073
rect 4632 29034 4660 29446
rect 3974 28999 4030 29008
rect 4620 29028 4672 29034
rect 4620 28970 4672 28976
rect 4632 28626 4660 28970
rect 4816 28762 4844 29514
rect 5000 29170 5028 30126
rect 5368 29782 5396 30126
rect 5460 29850 5488 31078
rect 5552 30666 5580 32302
rect 6288 31958 6316 32914
rect 6656 32230 6684 35430
rect 6828 35012 6880 35018
rect 6828 34954 6880 34960
rect 6840 34542 6868 34954
rect 7104 34604 7156 34610
rect 7104 34546 7156 34552
rect 6828 34536 6880 34542
rect 6828 34478 6880 34484
rect 6840 34066 6868 34478
rect 6920 34400 6972 34406
rect 6920 34342 6972 34348
rect 6828 34060 6880 34066
rect 6828 34002 6880 34008
rect 6736 32360 6788 32366
rect 6736 32302 6788 32308
rect 6644 32224 6696 32230
rect 6644 32166 6696 32172
rect 6276 31952 6328 31958
rect 6276 31894 6328 31900
rect 5632 31476 5684 31482
rect 5632 31418 5684 31424
rect 5644 30734 5672 31418
rect 5632 30728 5684 30734
rect 5632 30670 5684 30676
rect 5540 30660 5592 30666
rect 5540 30602 5592 30608
rect 5552 29850 5580 30602
rect 5816 30320 5868 30326
rect 5816 30262 5868 30268
rect 5448 29844 5500 29850
rect 5448 29786 5500 29792
rect 5540 29844 5592 29850
rect 5540 29786 5592 29792
rect 5356 29776 5408 29782
rect 5356 29718 5408 29724
rect 5368 29306 5396 29718
rect 5448 29640 5500 29646
rect 5448 29582 5500 29588
rect 5356 29300 5408 29306
rect 5356 29242 5408 29248
rect 4988 29164 5040 29170
rect 4988 29106 5040 29112
rect 5264 29096 5316 29102
rect 5264 29038 5316 29044
rect 4804 28756 4856 28762
rect 4804 28698 4856 28704
rect 4620 28620 4672 28626
rect 4620 28562 4672 28568
rect 4068 28552 4120 28558
rect 4068 28494 4120 28500
rect 4080 28200 4108 28494
rect 4220 28316 4516 28336
rect 4276 28314 4300 28316
rect 4356 28314 4380 28316
rect 4436 28314 4460 28316
rect 4298 28262 4300 28314
rect 4362 28262 4374 28314
rect 4436 28262 4438 28314
rect 4276 28260 4300 28262
rect 4356 28260 4380 28262
rect 4436 28260 4460 28262
rect 4220 28240 4516 28260
rect 4080 28172 4200 28200
rect 4068 27940 4120 27946
rect 4068 27882 4120 27888
rect 4080 27538 4108 27882
rect 4172 27674 4200 28172
rect 4632 28150 4660 28562
rect 5276 28150 5304 29038
rect 5460 28558 5488 29582
rect 5724 29164 5776 29170
rect 5724 29106 5776 29112
rect 5632 29028 5684 29034
rect 5632 28970 5684 28976
rect 5644 28694 5672 28970
rect 5632 28688 5684 28694
rect 5632 28630 5684 28636
rect 5540 28620 5592 28626
rect 5540 28562 5592 28568
rect 5448 28552 5500 28558
rect 5448 28494 5500 28500
rect 4436 28144 4488 28150
rect 4436 28086 4488 28092
rect 4620 28144 4672 28150
rect 4620 28086 4672 28092
rect 5264 28144 5316 28150
rect 5264 28086 5316 28092
rect 4448 28014 4476 28086
rect 4436 28008 4488 28014
rect 4436 27950 4488 27956
rect 4160 27668 4212 27674
rect 4160 27610 4212 27616
rect 4632 27538 4660 28086
rect 5460 28014 5488 28494
rect 4988 28008 5040 28014
rect 4988 27950 5040 27956
rect 5448 28008 5500 28014
rect 5448 27950 5500 27956
rect 5000 27538 5028 27950
rect 5552 27606 5580 28562
rect 5644 28014 5672 28630
rect 5632 28008 5684 28014
rect 5632 27950 5684 27956
rect 5540 27600 5592 27606
rect 5540 27542 5592 27548
rect 3884 27532 3936 27538
rect 3884 27474 3936 27480
rect 4068 27532 4120 27538
rect 4068 27474 4120 27480
rect 4620 27532 4672 27538
rect 4620 27474 4672 27480
rect 4988 27532 5040 27538
rect 4988 27474 5040 27480
rect 3976 27396 4028 27402
rect 3976 27338 4028 27344
rect 3988 26450 4016 27338
rect 4220 27228 4516 27248
rect 4276 27226 4300 27228
rect 4356 27226 4380 27228
rect 4436 27226 4460 27228
rect 4298 27174 4300 27226
rect 4362 27174 4374 27226
rect 4436 27174 4438 27226
rect 4276 27172 4300 27174
rect 4356 27172 4380 27174
rect 4436 27172 4460 27174
rect 4220 27152 4516 27172
rect 5644 27130 5672 27950
rect 5736 27470 5764 29106
rect 5828 29102 5856 30262
rect 6000 29708 6052 29714
rect 6000 29650 6052 29656
rect 5816 29096 5868 29102
rect 5816 29038 5868 29044
rect 5724 27464 5776 27470
rect 5724 27406 5776 27412
rect 5828 27334 5856 29038
rect 6012 29034 6040 29650
rect 6000 29028 6052 29034
rect 6000 28970 6052 28976
rect 6552 28552 6604 28558
rect 6552 28494 6604 28500
rect 6000 27532 6052 27538
rect 6000 27474 6052 27480
rect 5724 27328 5776 27334
rect 5724 27270 5776 27276
rect 5816 27328 5868 27334
rect 5816 27270 5868 27276
rect 5632 27124 5684 27130
rect 5632 27066 5684 27072
rect 5736 26994 5764 27270
rect 5724 26988 5776 26994
rect 5724 26930 5776 26936
rect 6012 26926 6040 27474
rect 6564 27402 6592 28494
rect 6656 27946 6684 32166
rect 6748 31482 6776 32302
rect 6932 31890 6960 34342
rect 7116 34066 7144 34546
rect 7104 34060 7156 34066
rect 7104 34002 7156 34008
rect 7208 33454 7236 35974
rect 7392 35834 7420 36178
rect 7380 35828 7432 35834
rect 7380 35770 7432 35776
rect 7668 35154 7696 36246
rect 7748 35488 7800 35494
rect 7748 35430 7800 35436
rect 7656 35148 7708 35154
rect 7656 35090 7708 35096
rect 7668 35034 7696 35090
rect 7576 35006 7696 35034
rect 7196 33448 7248 33454
rect 7196 33390 7248 33396
rect 7208 32842 7236 33390
rect 7196 32836 7248 32842
rect 7196 32778 7248 32784
rect 7104 32360 7156 32366
rect 7104 32302 7156 32308
rect 7116 32026 7144 32302
rect 7104 32020 7156 32026
rect 7104 31962 7156 31968
rect 6920 31884 6972 31890
rect 6920 31826 6972 31832
rect 7012 31816 7064 31822
rect 7012 31758 7064 31764
rect 6736 31476 6788 31482
rect 6736 31418 6788 31424
rect 6828 31272 6880 31278
rect 6828 31214 6880 31220
rect 6840 30938 6868 31214
rect 6920 31136 6972 31142
rect 6920 31078 6972 31084
rect 6828 30932 6880 30938
rect 6828 30874 6880 30880
rect 6932 29782 6960 31078
rect 7024 30802 7052 31758
rect 7012 30796 7064 30802
rect 7012 30738 7064 30744
rect 7024 29866 7052 30738
rect 7576 30326 7604 35006
rect 7760 34678 7788 35430
rect 7852 35086 7880 36654
rect 8576 36644 8628 36650
rect 8576 36586 8628 36592
rect 8588 36378 8616 36586
rect 8576 36372 8628 36378
rect 8576 36314 8628 36320
rect 9324 36174 9352 37726
rect 9600 37194 9628 38422
rect 10876 38344 10928 38350
rect 10876 38286 10928 38292
rect 10888 38010 10916 38286
rect 10876 38004 10928 38010
rect 10876 37946 10928 37952
rect 12360 37942 12388 40200
rect 14384 38554 14412 40200
rect 14372 38548 14424 38554
rect 14372 38490 14424 38496
rect 12900 38412 12952 38418
rect 12900 38354 12952 38360
rect 14188 38412 14240 38418
rect 14188 38354 14240 38360
rect 14740 38412 14792 38418
rect 14740 38354 14792 38360
rect 12716 38208 12768 38214
rect 12716 38150 12768 38156
rect 9680 37936 9732 37942
rect 9680 37878 9732 37884
rect 12348 37936 12400 37942
rect 12348 37878 12400 37884
rect 9692 37330 9720 37878
rect 12728 37874 12756 38150
rect 12440 37868 12492 37874
rect 12440 37810 12492 37816
rect 12716 37868 12768 37874
rect 12716 37810 12768 37816
rect 10600 37800 10652 37806
rect 10600 37742 10652 37748
rect 11060 37800 11112 37806
rect 11060 37742 11112 37748
rect 10140 37392 10192 37398
rect 10140 37334 10192 37340
rect 9680 37324 9732 37330
rect 9680 37266 9732 37272
rect 9588 37188 9640 37194
rect 9588 37130 9640 37136
rect 9692 36854 9720 37266
rect 9680 36848 9732 36854
rect 9680 36790 9732 36796
rect 9956 36576 10008 36582
rect 9956 36518 10008 36524
rect 9680 36304 9732 36310
rect 9680 36246 9732 36252
rect 9312 36168 9364 36174
rect 9312 36110 9364 36116
rect 7932 36032 7984 36038
rect 7932 35974 7984 35980
rect 7944 35562 7972 35974
rect 8024 35828 8076 35834
rect 8024 35770 8076 35776
rect 7932 35556 7984 35562
rect 7932 35498 7984 35504
rect 7840 35080 7892 35086
rect 7840 35022 7892 35028
rect 7748 34672 7800 34678
rect 7748 34614 7800 34620
rect 7760 34542 7788 34614
rect 7656 34536 7708 34542
rect 7656 34478 7708 34484
rect 7748 34536 7800 34542
rect 7748 34478 7800 34484
rect 7668 33658 7696 34478
rect 7852 34202 7880 35022
rect 7840 34196 7892 34202
rect 7840 34138 7892 34144
rect 8036 34066 8064 35770
rect 9324 35698 9352 36110
rect 9692 36038 9720 36246
rect 9968 36242 9996 36518
rect 9956 36236 10008 36242
rect 9956 36178 10008 36184
rect 9680 36032 9732 36038
rect 9680 35974 9732 35980
rect 9312 35692 9364 35698
rect 9312 35634 9364 35640
rect 8024 34060 8076 34066
rect 8024 34002 8076 34008
rect 8944 34060 8996 34066
rect 8944 34002 8996 34008
rect 7656 33652 7708 33658
rect 7656 33594 7708 33600
rect 8036 32978 8064 34002
rect 8956 33590 8984 34002
rect 8944 33584 8996 33590
rect 8944 33526 8996 33532
rect 8208 33448 8260 33454
rect 8208 33390 8260 33396
rect 8024 32972 8076 32978
rect 8024 32914 8076 32920
rect 8220 32570 8248 33390
rect 8576 33312 8628 33318
rect 8576 33254 8628 33260
rect 8208 32564 8260 32570
rect 8208 32506 8260 32512
rect 8588 32434 8616 33254
rect 8668 32972 8720 32978
rect 8668 32914 8720 32920
rect 8576 32428 8628 32434
rect 8576 32370 8628 32376
rect 7748 31272 7800 31278
rect 7748 31214 7800 31220
rect 7760 30394 7788 31214
rect 8300 30796 8352 30802
rect 8300 30738 8352 30744
rect 7748 30388 7800 30394
rect 7748 30330 7800 30336
rect 7564 30320 7616 30326
rect 7564 30262 7616 30268
rect 7840 30116 7892 30122
rect 7840 30058 7892 30064
rect 7656 30048 7708 30054
rect 7656 29990 7708 29996
rect 7024 29838 7144 29866
rect 6920 29776 6972 29782
rect 6920 29718 6972 29724
rect 7012 29708 7064 29714
rect 7012 29650 7064 29656
rect 7024 29102 7052 29650
rect 7012 29096 7064 29102
rect 7012 29038 7064 29044
rect 7024 28762 7052 29038
rect 7012 28756 7064 28762
rect 7012 28698 7064 28704
rect 6920 28144 6972 28150
rect 6920 28086 6972 28092
rect 6644 27940 6696 27946
rect 6644 27882 6696 27888
rect 6656 27470 6684 27882
rect 6932 27606 6960 28086
rect 6920 27600 6972 27606
rect 6920 27542 6972 27548
rect 6644 27464 6696 27470
rect 6644 27406 6696 27412
rect 6552 27396 6604 27402
rect 6552 27338 6604 27344
rect 6564 26926 6592 27338
rect 6656 27130 6684 27406
rect 6644 27124 6696 27130
rect 6644 27066 6696 27072
rect 4252 26920 4304 26926
rect 4252 26862 4304 26868
rect 4804 26920 4856 26926
rect 4804 26862 4856 26868
rect 5632 26920 5684 26926
rect 5632 26862 5684 26868
rect 6000 26920 6052 26926
rect 6000 26862 6052 26868
rect 6552 26920 6604 26926
rect 6552 26862 6604 26868
rect 4068 26580 4120 26586
rect 4068 26522 4120 26528
rect 3976 26444 4028 26450
rect 3976 26386 4028 26392
rect 4080 25974 4108 26522
rect 4264 26382 4292 26862
rect 4252 26376 4304 26382
rect 4252 26318 4304 26324
rect 4712 26376 4764 26382
rect 4712 26318 4764 26324
rect 4220 26140 4516 26160
rect 4276 26138 4300 26140
rect 4356 26138 4380 26140
rect 4436 26138 4460 26140
rect 4298 26086 4300 26138
rect 4362 26086 4374 26138
rect 4436 26086 4438 26138
rect 4276 26084 4300 26086
rect 4356 26084 4380 26086
rect 4436 26084 4460 26086
rect 4220 26064 4516 26084
rect 3608 25968 3660 25974
rect 3608 25910 3660 25916
rect 4068 25968 4120 25974
rect 4068 25910 4120 25916
rect 4080 25838 4108 25910
rect 3608 25832 3660 25838
rect 4068 25832 4120 25838
rect 3608 25774 3660 25780
rect 3988 25792 4068 25820
rect 3620 24750 3648 25774
rect 3988 24818 4016 25792
rect 4068 25774 4120 25780
rect 4620 25764 4672 25770
rect 4620 25706 4672 25712
rect 4068 25696 4120 25702
rect 4068 25638 4120 25644
rect 3976 24812 4028 24818
rect 3976 24754 4028 24760
rect 4080 24750 4108 25638
rect 4632 25362 4660 25706
rect 4724 25430 4752 26318
rect 4712 25424 4764 25430
rect 4712 25366 4764 25372
rect 4816 25362 4844 26862
rect 5644 26586 5672 26862
rect 5724 26784 5776 26790
rect 5724 26726 5776 26732
rect 5736 26586 5764 26726
rect 5632 26580 5684 26586
rect 5632 26522 5684 26528
rect 5724 26580 5776 26586
rect 5724 26522 5776 26528
rect 5356 26240 5408 26246
rect 5356 26182 5408 26188
rect 5368 25702 5396 26182
rect 5448 26036 5500 26042
rect 5448 25978 5500 25984
rect 5460 25906 5488 25978
rect 5448 25900 5500 25906
rect 5448 25842 5500 25848
rect 5356 25696 5408 25702
rect 5356 25638 5408 25644
rect 4620 25356 4672 25362
rect 4620 25298 4672 25304
rect 4804 25356 4856 25362
rect 4804 25298 4856 25304
rect 4220 25052 4516 25072
rect 4276 25050 4300 25052
rect 4356 25050 4380 25052
rect 4436 25050 4460 25052
rect 4298 24998 4300 25050
rect 4362 24998 4374 25050
rect 4436 24998 4438 25050
rect 4276 24996 4300 24998
rect 4356 24996 4380 24998
rect 4436 24996 4460 24998
rect 4220 24976 4516 24996
rect 3608 24744 3660 24750
rect 3608 24686 3660 24692
rect 3700 24744 3752 24750
rect 3700 24686 3752 24692
rect 4068 24744 4120 24750
rect 4068 24686 4120 24692
rect 3712 23798 3740 24686
rect 3976 24268 4028 24274
rect 3976 24210 4028 24216
rect 3700 23792 3752 23798
rect 3700 23734 3752 23740
rect 3988 23662 4016 24210
rect 4816 24206 4844 25298
rect 4804 24200 4856 24206
rect 4804 24142 4856 24148
rect 4988 24200 5040 24206
rect 4988 24142 5040 24148
rect 4620 24064 4672 24070
rect 4620 24006 4672 24012
rect 4220 23964 4516 23984
rect 4276 23962 4300 23964
rect 4356 23962 4380 23964
rect 4436 23962 4460 23964
rect 4298 23910 4300 23962
rect 4362 23910 4374 23962
rect 4436 23910 4438 23962
rect 4276 23908 4300 23910
rect 4356 23908 4380 23910
rect 4436 23908 4460 23910
rect 4220 23888 4516 23908
rect 3976 23656 4028 23662
rect 3976 23598 4028 23604
rect 3988 23254 4016 23598
rect 3976 23248 4028 23254
rect 3976 23190 4028 23196
rect 4220 22876 4516 22896
rect 4276 22874 4300 22876
rect 4356 22874 4380 22876
rect 4436 22874 4460 22876
rect 4298 22822 4300 22874
rect 4362 22822 4374 22874
rect 4436 22822 4438 22874
rect 4276 22820 4300 22822
rect 4356 22820 4380 22822
rect 4436 22820 4460 22822
rect 4220 22800 4516 22820
rect 4632 22642 4660 24006
rect 4816 22710 4844 24142
rect 5000 23526 5028 24142
rect 4988 23520 5040 23526
rect 4988 23462 5040 23468
rect 4896 23180 4948 23186
rect 4896 23122 4948 23128
rect 4804 22704 4856 22710
rect 4804 22646 4856 22652
rect 4620 22636 4672 22642
rect 4620 22578 4672 22584
rect 4908 22574 4936 23122
rect 4528 22568 4580 22574
rect 4528 22510 4580 22516
rect 4896 22568 4948 22574
rect 4896 22510 4948 22516
rect 4540 22098 4568 22510
rect 4528 22092 4580 22098
rect 4528 22034 4580 22040
rect 4220 21788 4516 21808
rect 4276 21786 4300 21788
rect 4356 21786 4380 21788
rect 4436 21786 4460 21788
rect 4298 21734 4300 21786
rect 4362 21734 4374 21786
rect 4436 21734 4438 21786
rect 4276 21732 4300 21734
rect 4356 21732 4380 21734
rect 4436 21732 4460 21734
rect 4220 21712 4516 21732
rect 4908 21554 4936 22510
rect 5000 22098 5028 23462
rect 5460 23322 5488 25842
rect 5644 25362 5672 26522
rect 6012 26450 6040 26862
rect 6000 26444 6052 26450
rect 6000 26386 6052 26392
rect 5908 25968 5960 25974
rect 5908 25910 5960 25916
rect 5724 25832 5776 25838
rect 5724 25774 5776 25780
rect 5736 25498 5764 25774
rect 5920 25702 5948 25910
rect 6184 25832 6236 25838
rect 6182 25800 6184 25809
rect 6236 25800 6238 25809
rect 6182 25735 6238 25744
rect 5908 25696 5960 25702
rect 5908 25638 5960 25644
rect 5724 25492 5776 25498
rect 5724 25434 5776 25440
rect 6564 25362 6592 26862
rect 5632 25356 5684 25362
rect 5632 25298 5684 25304
rect 6552 25356 6604 25362
rect 6552 25298 6604 25304
rect 5724 24880 5776 24886
rect 5724 24822 5776 24828
rect 5632 24744 5684 24750
rect 5632 24686 5684 24692
rect 5644 24070 5672 24686
rect 5632 24064 5684 24070
rect 5632 24006 5684 24012
rect 5736 23662 5764 24822
rect 6184 24676 6236 24682
rect 6184 24618 6236 24624
rect 6196 23662 6224 24618
rect 5724 23656 5776 23662
rect 5724 23598 5776 23604
rect 6184 23656 6236 23662
rect 6184 23598 6236 23604
rect 5448 23316 5500 23322
rect 5448 23258 5500 23264
rect 5080 23180 5132 23186
rect 5080 23122 5132 23128
rect 6000 23180 6052 23186
rect 6000 23122 6052 23128
rect 5092 22778 5120 23122
rect 5908 22976 5960 22982
rect 5908 22918 5960 22924
rect 5080 22772 5132 22778
rect 5080 22714 5132 22720
rect 5920 22642 5948 22918
rect 5908 22636 5960 22642
rect 5908 22578 5960 22584
rect 6012 22574 6040 23122
rect 6196 22642 6224 23598
rect 6656 23186 6684 27066
rect 6920 25288 6972 25294
rect 6920 25230 6972 25236
rect 6932 24614 6960 25230
rect 7116 24750 7144 29838
rect 7472 29504 7524 29510
rect 7472 29446 7524 29452
rect 7484 29170 7512 29446
rect 7472 29164 7524 29170
rect 7472 29106 7524 29112
rect 7668 28422 7696 29990
rect 7656 28416 7708 28422
rect 7656 28358 7708 28364
rect 7196 28008 7248 28014
rect 7196 27950 7248 27956
rect 7380 28008 7432 28014
rect 7380 27950 7432 27956
rect 7208 26382 7236 27950
rect 7392 27606 7420 27950
rect 7380 27600 7432 27606
rect 7380 27542 7432 27548
rect 7668 27538 7696 28358
rect 7852 28218 7880 30058
rect 8312 29782 8340 30738
rect 8484 30728 8536 30734
rect 8484 30670 8536 30676
rect 8496 30394 8524 30670
rect 8484 30388 8536 30394
rect 8484 30330 8536 30336
rect 8300 29776 8352 29782
rect 8300 29718 8352 29724
rect 8484 29164 8536 29170
rect 8484 29106 8536 29112
rect 8300 29096 8352 29102
rect 8300 29038 8352 29044
rect 8312 28762 8340 29038
rect 8300 28756 8352 28762
rect 8300 28698 8352 28704
rect 8496 28626 8524 29106
rect 8484 28620 8536 28626
rect 8484 28562 8536 28568
rect 7840 28212 7892 28218
rect 7840 28154 7892 28160
rect 8300 28008 8352 28014
rect 8300 27950 8352 27956
rect 8312 27606 8340 27950
rect 8300 27600 8352 27606
rect 8300 27542 8352 27548
rect 7656 27532 7708 27538
rect 7576 27492 7656 27520
rect 7380 26444 7432 26450
rect 7380 26386 7432 26392
rect 7196 26376 7248 26382
rect 7196 26318 7248 26324
rect 7392 25906 7420 26386
rect 7380 25900 7432 25906
rect 7380 25842 7432 25848
rect 7576 24818 7604 27492
rect 7656 27474 7708 27480
rect 7932 27532 7984 27538
rect 7932 27474 7984 27480
rect 7748 26444 7800 26450
rect 7748 26386 7800 26392
rect 7760 25838 7788 26386
rect 7748 25832 7800 25838
rect 7748 25774 7800 25780
rect 7656 25696 7708 25702
rect 7656 25638 7708 25644
rect 7564 24812 7616 24818
rect 7564 24754 7616 24760
rect 7668 24750 7696 25638
rect 7760 25294 7788 25774
rect 7748 25288 7800 25294
rect 7748 25230 7800 25236
rect 7944 24818 7972 27474
rect 8312 27334 8340 27542
rect 8576 27464 8628 27470
rect 8576 27406 8628 27412
rect 8300 27328 8352 27334
rect 8300 27270 8352 27276
rect 8588 26858 8616 27406
rect 8576 26852 8628 26858
rect 8576 26794 8628 26800
rect 8588 26450 8616 26794
rect 8116 26444 8168 26450
rect 8116 26386 8168 26392
rect 8576 26444 8628 26450
rect 8576 26386 8628 26392
rect 8128 25838 8156 26386
rect 8116 25832 8168 25838
rect 8116 25774 8168 25780
rect 8128 25498 8156 25774
rect 8116 25492 8168 25498
rect 8116 25434 8168 25440
rect 7932 24812 7984 24818
rect 7932 24754 7984 24760
rect 7104 24744 7156 24750
rect 7104 24686 7156 24692
rect 7656 24744 7708 24750
rect 7656 24686 7708 24692
rect 6920 24608 6972 24614
rect 6920 24550 6972 24556
rect 7116 24410 7144 24686
rect 7104 24404 7156 24410
rect 7104 24346 7156 24352
rect 7748 24336 7800 24342
rect 7748 24278 7800 24284
rect 7104 24268 7156 24274
rect 7104 24210 7156 24216
rect 6828 24064 6880 24070
rect 6828 24006 6880 24012
rect 6840 23594 6868 24006
rect 7116 23798 7144 24210
rect 7760 23866 7788 24278
rect 7748 23860 7800 23866
rect 7748 23802 7800 23808
rect 8024 23860 8076 23866
rect 8024 23802 8076 23808
rect 7104 23792 7156 23798
rect 7104 23734 7156 23740
rect 7840 23656 7892 23662
rect 7840 23598 7892 23604
rect 6828 23588 6880 23594
rect 6828 23530 6880 23536
rect 6644 23180 6696 23186
rect 6644 23122 6696 23128
rect 6736 23112 6788 23118
rect 6736 23054 6788 23060
rect 6184 22636 6236 22642
rect 6184 22578 6236 22584
rect 5632 22568 5684 22574
rect 5552 22528 5632 22556
rect 4988 22092 5040 22098
rect 4988 22034 5040 22040
rect 5552 22030 5580 22528
rect 5632 22510 5684 22516
rect 6000 22568 6052 22574
rect 6000 22510 6052 22516
rect 5540 22024 5592 22030
rect 5540 21966 5592 21972
rect 5552 21622 5580 21966
rect 5540 21616 5592 21622
rect 5592 21564 5672 21570
rect 5540 21558 5672 21564
rect 3976 21548 4028 21554
rect 3976 21490 4028 21496
rect 4896 21548 4948 21554
rect 5552 21542 5672 21558
rect 4896 21490 4948 21496
rect 3988 20874 4016 21490
rect 4068 21480 4120 21486
rect 4068 21422 4120 21428
rect 4988 21480 5040 21486
rect 4988 21422 5040 21428
rect 3976 20868 4028 20874
rect 3976 20810 4028 20816
rect 3988 20244 4016 20810
rect 4080 20398 4108 21422
rect 5000 20942 5028 21422
rect 5540 21412 5592 21418
rect 5540 21354 5592 21360
rect 5552 21146 5580 21354
rect 5540 21140 5592 21146
rect 5540 21082 5592 21088
rect 5644 21010 5672 21542
rect 6748 21486 6776 23054
rect 6840 22574 6868 23530
rect 7852 23322 7880 23598
rect 7840 23316 7892 23322
rect 7840 23258 7892 23264
rect 7852 23186 7880 23258
rect 7380 23180 7432 23186
rect 7380 23122 7432 23128
rect 7840 23180 7892 23186
rect 7840 23122 7892 23128
rect 7196 23044 7248 23050
rect 7196 22986 7248 22992
rect 6828 22568 6880 22574
rect 6828 22510 6880 22516
rect 7208 22030 7236 22986
rect 7392 22574 7420 23122
rect 7472 22976 7524 22982
rect 7472 22918 7524 22924
rect 7380 22568 7432 22574
rect 7380 22510 7432 22516
rect 7392 22234 7420 22510
rect 7380 22228 7432 22234
rect 7380 22170 7432 22176
rect 6920 22024 6972 22030
rect 6920 21966 6972 21972
rect 7196 22024 7248 22030
rect 7196 21966 7248 21972
rect 6932 21622 6960 21966
rect 6920 21616 6972 21622
rect 6920 21558 6972 21564
rect 6736 21480 6788 21486
rect 6736 21422 6788 21428
rect 5908 21140 5960 21146
rect 5908 21082 5960 21088
rect 5632 21004 5684 21010
rect 5632 20946 5684 20952
rect 4988 20936 5040 20942
rect 4988 20878 5040 20884
rect 5816 20936 5868 20942
rect 5816 20878 5868 20884
rect 4620 20800 4672 20806
rect 4620 20742 4672 20748
rect 4220 20700 4516 20720
rect 4276 20698 4300 20700
rect 4356 20698 4380 20700
rect 4436 20698 4460 20700
rect 4298 20646 4300 20698
rect 4362 20646 4374 20698
rect 4436 20646 4438 20698
rect 4276 20644 4300 20646
rect 4356 20644 4380 20646
rect 4436 20644 4460 20646
rect 4220 20624 4516 20644
rect 4632 20602 4660 20742
rect 4620 20596 4672 20602
rect 4620 20538 4672 20544
rect 4068 20392 4120 20398
rect 4068 20334 4120 20340
rect 4160 20324 4212 20330
rect 4160 20266 4212 20272
rect 3988 20216 4108 20244
rect 3528 19910 3740 19938
rect 4080 19922 4108 20216
rect 3516 19848 3568 19854
rect 3516 19790 3568 19796
rect 3528 19378 3556 19790
rect 3516 19372 3568 19378
rect 3516 19314 3568 19320
rect 3528 18834 3556 19314
rect 3712 19258 3740 19910
rect 4068 19916 4120 19922
rect 4068 19858 4120 19864
rect 3976 19848 4028 19854
rect 4172 19802 4200 20266
rect 5000 19922 5028 20878
rect 5080 20800 5132 20806
rect 5080 20742 5132 20748
rect 5092 20466 5120 20742
rect 5080 20460 5132 20466
rect 5080 20402 5132 20408
rect 5828 20398 5856 20878
rect 5816 20392 5868 20398
rect 5816 20334 5868 20340
rect 5828 19922 5856 20334
rect 4804 19916 4856 19922
rect 4804 19858 4856 19864
rect 4988 19916 5040 19922
rect 4988 19858 5040 19864
rect 5816 19916 5868 19922
rect 5816 19858 5868 19864
rect 3976 19790 4028 19796
rect 3884 19304 3936 19310
rect 3712 19252 3884 19258
rect 3712 19246 3936 19252
rect 3712 19230 3924 19246
rect 3516 18828 3568 18834
rect 3516 18770 3568 18776
rect 3988 18222 4016 19790
rect 4080 19774 4200 19802
rect 4712 19780 4764 19786
rect 4080 19428 4108 19774
rect 4712 19722 4764 19728
rect 4220 19612 4516 19632
rect 4276 19610 4300 19612
rect 4356 19610 4380 19612
rect 4436 19610 4460 19612
rect 4298 19558 4300 19610
rect 4362 19558 4374 19610
rect 4436 19558 4438 19610
rect 4276 19556 4300 19558
rect 4356 19556 4380 19558
rect 4436 19556 4460 19558
rect 4220 19536 4516 19556
rect 4620 19508 4672 19514
rect 4620 19450 4672 19456
rect 4080 19400 4200 19428
rect 4172 18970 4200 19400
rect 4160 18964 4212 18970
rect 4160 18906 4212 18912
rect 4220 18524 4516 18544
rect 4276 18522 4300 18524
rect 4356 18522 4380 18524
rect 4436 18522 4460 18524
rect 4298 18470 4300 18522
rect 4362 18470 4374 18522
rect 4436 18470 4438 18522
rect 4276 18468 4300 18470
rect 4356 18468 4380 18470
rect 4436 18468 4460 18470
rect 4220 18448 4516 18468
rect 3976 18216 4028 18222
rect 3976 18158 4028 18164
rect 4632 18154 4660 19450
rect 4724 18290 4752 19722
rect 4816 19242 4844 19858
rect 5000 19514 5028 19858
rect 4988 19508 5040 19514
rect 4988 19450 5040 19456
rect 5920 19310 5948 21082
rect 6920 20936 6972 20942
rect 6920 20878 6972 20884
rect 6828 20460 6880 20466
rect 6828 20402 6880 20408
rect 6840 19922 6868 20402
rect 6828 19916 6880 19922
rect 6828 19858 6880 19864
rect 6000 19848 6052 19854
rect 6000 19790 6052 19796
rect 5908 19304 5960 19310
rect 5908 19246 5960 19252
rect 4804 19236 4856 19242
rect 4804 19178 4856 19184
rect 6012 18970 6040 19790
rect 6000 18964 6052 18970
rect 6000 18906 6052 18912
rect 6840 18834 6868 19858
rect 6932 19174 6960 20878
rect 7104 19712 7156 19718
rect 7104 19654 7156 19660
rect 6920 19168 6972 19174
rect 6920 19110 6972 19116
rect 7116 18834 7144 19654
rect 7208 19310 7236 21966
rect 7484 21486 7512 22918
rect 7852 22506 7880 23122
rect 7840 22500 7892 22506
rect 7840 22442 7892 22448
rect 8036 22098 8064 23802
rect 8680 23186 8708 32914
rect 9324 32366 9352 35634
rect 9496 34536 9548 34542
rect 9496 34478 9548 34484
rect 9508 34202 9536 34478
rect 9496 34196 9548 34202
rect 9496 34138 9548 34144
rect 9864 34060 9916 34066
rect 9864 34002 9916 34008
rect 9680 33856 9732 33862
rect 9680 33798 9732 33804
rect 9692 33454 9720 33798
rect 9876 33658 9904 34002
rect 9864 33652 9916 33658
rect 9864 33594 9916 33600
rect 9680 33448 9732 33454
rect 9680 33390 9732 33396
rect 10048 33448 10100 33454
rect 10048 33390 10100 33396
rect 9772 33380 9824 33386
rect 9772 33322 9824 33328
rect 9680 32428 9732 32434
rect 9680 32370 9732 32376
rect 9312 32360 9364 32366
rect 9312 32302 9364 32308
rect 8760 31884 8812 31890
rect 8760 31826 8812 31832
rect 8772 30938 8800 31826
rect 9220 31204 9272 31210
rect 9220 31146 9272 31152
rect 8760 30932 8812 30938
rect 8760 30874 8812 30880
rect 8944 30864 8996 30870
rect 8944 30806 8996 30812
rect 8760 30660 8812 30666
rect 8760 30602 8812 30608
rect 8772 29714 8800 30602
rect 8956 30394 8984 30806
rect 8944 30388 8996 30394
rect 8944 30330 8996 30336
rect 9232 30190 9260 31146
rect 9324 30598 9352 32302
rect 9496 32224 9548 32230
rect 9496 32166 9548 32172
rect 9508 31958 9536 32166
rect 9496 31952 9548 31958
rect 9692 31906 9720 32370
rect 9496 31894 9548 31900
rect 9600 31890 9720 31906
rect 9588 31884 9720 31890
rect 9640 31878 9720 31884
rect 9588 31826 9640 31832
rect 9692 30802 9720 31878
rect 9784 31754 9812 33322
rect 10060 33046 10088 33390
rect 10048 33040 10100 33046
rect 10048 32982 10100 32988
rect 9772 31748 9824 31754
rect 9772 31690 9824 31696
rect 9680 30796 9732 30802
rect 9680 30738 9732 30744
rect 9312 30592 9364 30598
rect 9312 30534 9364 30540
rect 9036 30184 9088 30190
rect 9036 30126 9088 30132
rect 9220 30184 9272 30190
rect 9220 30126 9272 30132
rect 8760 29708 8812 29714
rect 8760 29650 8812 29656
rect 8944 29708 8996 29714
rect 8944 29650 8996 29656
rect 8772 28218 8800 29650
rect 8956 28626 8984 29650
rect 9048 29034 9076 30126
rect 9232 29646 9260 30126
rect 9220 29640 9272 29646
rect 9220 29582 9272 29588
rect 9232 29238 9260 29582
rect 9220 29232 9272 29238
rect 9220 29174 9272 29180
rect 9324 29102 9352 30534
rect 9404 29708 9456 29714
rect 9404 29650 9456 29656
rect 9416 29209 9444 29650
rect 10046 29608 10102 29617
rect 10046 29543 10102 29552
rect 9402 29200 9458 29209
rect 9402 29135 9458 29144
rect 9312 29096 9364 29102
rect 9312 29038 9364 29044
rect 9956 29096 10008 29102
rect 9956 29038 10008 29044
rect 9036 29028 9088 29034
rect 9036 28970 9088 28976
rect 8944 28620 8996 28626
rect 8944 28562 8996 28568
rect 9128 28620 9180 28626
rect 9128 28562 9180 28568
rect 8760 28212 8812 28218
rect 8760 28154 8812 28160
rect 9140 28014 9168 28562
rect 9324 28558 9352 29038
rect 9864 28960 9916 28966
rect 9864 28902 9916 28908
rect 9312 28552 9364 28558
rect 9312 28494 9364 28500
rect 9128 28008 9180 28014
rect 9128 27950 9180 27956
rect 9140 27538 9168 27950
rect 9876 27878 9904 28902
rect 9968 28082 9996 29038
rect 9956 28076 10008 28082
rect 9956 28018 10008 28024
rect 10060 28014 10088 29543
rect 10152 29102 10180 37334
rect 10324 36712 10376 36718
rect 10612 36689 10640 37742
rect 10692 37324 10744 37330
rect 10744 37284 10824 37312
rect 10692 37266 10744 37272
rect 10324 36654 10376 36660
rect 10598 36680 10654 36689
rect 10232 29708 10284 29714
rect 10232 29650 10284 29656
rect 10140 29096 10192 29102
rect 10140 29038 10192 29044
rect 10152 28966 10180 29038
rect 10140 28960 10192 28966
rect 10140 28902 10192 28908
rect 10244 28014 10272 29650
rect 10048 28008 10100 28014
rect 10048 27950 10100 27956
rect 10232 28008 10284 28014
rect 10232 27950 10284 27956
rect 9864 27872 9916 27878
rect 9864 27814 9916 27820
rect 10244 27538 10272 27950
rect 9128 27532 9180 27538
rect 9128 27474 9180 27480
rect 10232 27532 10284 27538
rect 10232 27474 10284 27480
rect 9036 27328 9088 27334
rect 9036 27270 9088 27276
rect 9048 26926 9076 27270
rect 9036 26920 9088 26926
rect 9036 26862 9088 26868
rect 9036 25764 9088 25770
rect 9036 25706 9088 25712
rect 8852 25696 8904 25702
rect 8852 25638 8904 25644
rect 8864 25362 8892 25638
rect 9048 25498 9076 25706
rect 9036 25492 9088 25498
rect 9036 25434 9088 25440
rect 8852 25356 8904 25362
rect 8852 25298 8904 25304
rect 8760 24744 8812 24750
rect 8760 24686 8812 24692
rect 8772 24410 8800 24686
rect 8760 24404 8812 24410
rect 8760 24346 8812 24352
rect 9048 24274 9076 25434
rect 9036 24268 9088 24274
rect 9036 24210 9088 24216
rect 9036 23656 9088 23662
rect 9036 23598 9088 23604
rect 9048 23254 9076 23598
rect 9036 23248 9088 23254
rect 9036 23190 9088 23196
rect 8668 23180 8720 23186
rect 8588 23140 8668 23168
rect 8300 22568 8352 22574
rect 8300 22510 8352 22516
rect 8312 22234 8340 22510
rect 8300 22228 8352 22234
rect 8300 22170 8352 22176
rect 8024 22092 8076 22098
rect 8024 22034 8076 22040
rect 7472 21480 7524 21486
rect 7472 21422 7524 21428
rect 8208 20392 8260 20398
rect 8208 20334 8260 20340
rect 8220 19990 8248 20334
rect 8208 19984 8260 19990
rect 8208 19926 8260 19932
rect 8588 19310 8616 23140
rect 8668 23122 8720 23128
rect 9048 22098 9076 23190
rect 8852 22092 8904 22098
rect 8852 22034 8904 22040
rect 9036 22092 9088 22098
rect 9036 22034 9088 22040
rect 8864 21078 8892 22034
rect 9140 21978 9168 27474
rect 9680 26784 9732 26790
rect 9680 26726 9732 26732
rect 9692 26382 9720 26726
rect 9680 26376 9732 26382
rect 9680 26318 9732 26324
rect 9864 26376 9916 26382
rect 9864 26318 9916 26324
rect 9404 26036 9456 26042
rect 9404 25978 9456 25984
rect 9416 23186 9444 25978
rect 9496 25832 9548 25838
rect 9496 25774 9548 25780
rect 9508 25498 9536 25774
rect 9496 25492 9548 25498
rect 9496 25434 9548 25440
rect 9692 24614 9720 26318
rect 9876 25906 9904 26318
rect 9956 25968 10008 25974
rect 9956 25910 10008 25916
rect 9864 25900 9916 25906
rect 9864 25842 9916 25848
rect 9968 25838 9996 25910
rect 9956 25832 10008 25838
rect 9956 25774 10008 25780
rect 9968 25498 9996 25774
rect 9956 25492 10008 25498
rect 9956 25434 10008 25440
rect 9864 25356 9916 25362
rect 9864 25298 9916 25304
rect 9680 24608 9732 24614
rect 9680 24550 9732 24556
rect 9680 23724 9732 23730
rect 9680 23666 9732 23672
rect 9404 23180 9456 23186
rect 9404 23122 9456 23128
rect 9692 22098 9720 23666
rect 9772 23656 9824 23662
rect 9772 23598 9824 23604
rect 9784 23322 9812 23598
rect 9772 23316 9824 23322
rect 9772 23258 9824 23264
rect 9680 22092 9732 22098
rect 9680 22034 9732 22040
rect 9048 21950 9168 21978
rect 8852 21072 8904 21078
rect 8852 21014 8904 21020
rect 8668 20868 8720 20874
rect 8668 20810 8720 20816
rect 8680 19922 8708 20810
rect 8668 19916 8720 19922
rect 8668 19858 8720 19864
rect 9048 19310 9076 21950
rect 9876 21146 9904 25298
rect 9956 24608 10008 24614
rect 9956 24550 10008 24556
rect 9968 24070 9996 24550
rect 9956 24064 10008 24070
rect 9956 24006 10008 24012
rect 9968 22574 9996 24006
rect 9956 22568 10008 22574
rect 9956 22510 10008 22516
rect 9956 22092 10008 22098
rect 9956 22034 10008 22040
rect 9864 21140 9916 21146
rect 9864 21082 9916 21088
rect 9128 20936 9180 20942
rect 9128 20878 9180 20884
rect 9140 20262 9168 20878
rect 9128 20256 9180 20262
rect 9128 20198 9180 20204
rect 9140 19990 9168 20198
rect 9128 19984 9180 19990
rect 9128 19926 9180 19932
rect 7196 19304 7248 19310
rect 7196 19246 7248 19252
rect 8576 19304 8628 19310
rect 8576 19246 8628 19252
rect 9036 19304 9088 19310
rect 9036 19246 9088 19252
rect 5172 18828 5224 18834
rect 5172 18770 5224 18776
rect 6276 18828 6328 18834
rect 6276 18770 6328 18776
rect 6828 18828 6880 18834
rect 6828 18770 6880 18776
rect 7104 18828 7156 18834
rect 7104 18770 7156 18776
rect 5080 18760 5132 18766
rect 5080 18702 5132 18708
rect 4712 18284 4764 18290
rect 4712 18226 4764 18232
rect 4620 18148 4672 18154
rect 4620 18090 4672 18096
rect 4068 17672 4120 17678
rect 4068 17614 4120 17620
rect 4080 16454 4108 17614
rect 5092 17542 5120 18702
rect 5184 18426 5212 18770
rect 5172 18420 5224 18426
rect 5172 18362 5224 18368
rect 5448 18216 5500 18222
rect 5448 18158 5500 18164
rect 5264 17740 5316 17746
rect 5316 17700 5396 17728
rect 5264 17682 5316 17688
rect 5080 17536 5132 17542
rect 5080 17478 5132 17484
rect 4220 17436 4516 17456
rect 4276 17434 4300 17436
rect 4356 17434 4380 17436
rect 4436 17434 4460 17436
rect 4298 17382 4300 17434
rect 4362 17382 4374 17434
rect 4436 17382 4438 17434
rect 4276 17380 4300 17382
rect 4356 17380 4380 17382
rect 4436 17380 4460 17382
rect 4220 17360 4516 17380
rect 5092 17202 5120 17478
rect 4712 17196 4764 17202
rect 4712 17138 4764 17144
rect 5080 17196 5132 17202
rect 5080 17138 5132 17144
rect 4724 16658 4752 17138
rect 5264 16788 5316 16794
rect 5264 16730 5316 16736
rect 4620 16652 4672 16658
rect 4620 16594 4672 16600
rect 4712 16652 4764 16658
rect 4712 16594 4764 16600
rect 4068 16448 4120 16454
rect 4068 16390 4120 16396
rect 4220 16348 4516 16368
rect 4276 16346 4300 16348
rect 4356 16346 4380 16348
rect 4436 16346 4460 16348
rect 4298 16294 4300 16346
rect 4362 16294 4374 16346
rect 4436 16294 4438 16346
rect 4276 16292 4300 16294
rect 4356 16292 4380 16294
rect 4436 16292 4460 16294
rect 4220 16272 4516 16292
rect 4632 16250 4660 16594
rect 4620 16244 4672 16250
rect 4620 16186 4672 16192
rect 5276 16114 5304 16730
rect 5368 16522 5396 17700
rect 5460 17678 5488 18158
rect 6092 18148 6144 18154
rect 6092 18090 6144 18096
rect 6104 17678 6132 18090
rect 5448 17672 5500 17678
rect 5448 17614 5500 17620
rect 6092 17672 6144 17678
rect 6092 17614 6144 17620
rect 5540 17128 5592 17134
rect 5540 17070 5592 17076
rect 5356 16516 5408 16522
rect 5356 16458 5408 16464
rect 5264 16108 5316 16114
rect 5264 16050 5316 16056
rect 5368 16046 5396 16458
rect 5552 16114 5580 17070
rect 6288 16726 6316 18770
rect 6840 18086 6868 18770
rect 7932 18624 7984 18630
rect 7932 18566 7984 18572
rect 6828 18080 6880 18086
rect 6828 18022 6880 18028
rect 7380 18080 7432 18086
rect 7380 18022 7432 18028
rect 6840 17202 6868 18022
rect 7392 17746 7420 18022
rect 7944 17746 7972 18566
rect 8392 18284 8444 18290
rect 8392 18226 8444 18232
rect 8024 18216 8076 18222
rect 8024 18158 8076 18164
rect 8036 17814 8064 18158
rect 8024 17808 8076 17814
rect 8024 17750 8076 17756
rect 7380 17740 7432 17746
rect 7380 17682 7432 17688
rect 7932 17740 7984 17746
rect 7932 17682 7984 17688
rect 7196 17672 7248 17678
rect 7196 17614 7248 17620
rect 6828 17196 6880 17202
rect 6828 17138 6880 17144
rect 6276 16720 6328 16726
rect 6276 16662 6328 16668
rect 5724 16652 5776 16658
rect 5724 16594 5776 16600
rect 6552 16652 6604 16658
rect 6552 16594 6604 16600
rect 5540 16108 5592 16114
rect 5540 16050 5592 16056
rect 5356 16040 5408 16046
rect 5356 15982 5408 15988
rect 5172 15496 5224 15502
rect 5172 15438 5224 15444
rect 4220 15260 4516 15280
rect 4276 15258 4300 15260
rect 4356 15258 4380 15260
rect 4436 15258 4460 15260
rect 4298 15206 4300 15258
rect 4362 15206 4374 15258
rect 4436 15206 4438 15258
rect 4276 15204 4300 15206
rect 4356 15204 4380 15206
rect 4436 15204 4460 15206
rect 4220 15184 4516 15204
rect 5184 15162 5212 15438
rect 4068 15156 4120 15162
rect 4068 15098 4120 15104
rect 5172 15156 5224 15162
rect 5172 15098 5224 15104
rect 4080 15065 4108 15098
rect 4066 15056 4122 15065
rect 4066 14991 4122 15000
rect 3882 14648 3938 14657
rect 3882 14583 3938 14592
rect 3896 14482 3924 14583
rect 5078 14512 5134 14521
rect 3884 14476 3936 14482
rect 5078 14447 5134 14456
rect 3884 14418 3936 14424
rect 4068 14408 4120 14414
rect 4068 14350 4120 14356
rect 4080 13734 4108 14350
rect 5092 14346 5120 14447
rect 5632 14408 5684 14414
rect 5632 14350 5684 14356
rect 5080 14340 5132 14346
rect 5080 14282 5132 14288
rect 4712 14272 4764 14278
rect 4712 14214 4764 14220
rect 4220 14172 4516 14192
rect 4276 14170 4300 14172
rect 4356 14170 4380 14172
rect 4436 14170 4460 14172
rect 4298 14118 4300 14170
rect 4362 14118 4374 14170
rect 4436 14118 4438 14170
rect 4276 14116 4300 14118
rect 4356 14116 4380 14118
rect 4436 14116 4460 14118
rect 4220 14096 4516 14116
rect 4068 13728 4120 13734
rect 4068 13670 4120 13676
rect 4344 13728 4396 13734
rect 4344 13670 4396 13676
rect 4080 13394 4108 13670
rect 4356 13394 4384 13670
rect 4068 13388 4120 13394
rect 4068 13330 4120 13336
rect 4344 13388 4396 13394
rect 4344 13330 4396 13336
rect 3792 13184 3844 13190
rect 3792 13126 3844 13132
rect 3804 12850 3832 13126
rect 3792 12844 3844 12850
rect 3792 12786 3844 12792
rect 4080 12782 4108 13330
rect 4220 13084 4516 13104
rect 4276 13082 4300 13084
rect 4356 13082 4380 13084
rect 4436 13082 4460 13084
rect 4298 13030 4300 13082
rect 4362 13030 4374 13082
rect 4436 13030 4438 13082
rect 4276 13028 4300 13030
rect 4356 13028 4380 13030
rect 4436 13028 4460 13030
rect 4220 13008 4516 13028
rect 4068 12776 4120 12782
rect 4068 12718 4120 12724
rect 4724 12306 4752 14214
rect 5540 14000 5592 14006
rect 5540 13942 5592 13948
rect 4896 13864 4948 13870
rect 4896 13806 4948 13812
rect 4908 12986 4936 13806
rect 4896 12980 4948 12986
rect 4896 12922 4948 12928
rect 5552 12306 5580 13942
rect 5644 13530 5672 14350
rect 5632 13524 5684 13530
rect 5632 13466 5684 13472
rect 4712 12300 4764 12306
rect 4712 12242 4764 12248
rect 5540 12300 5592 12306
rect 5540 12242 5592 12248
rect 3700 12096 3752 12102
rect 3700 12038 3752 12044
rect 3516 11756 3568 11762
rect 3516 11698 3568 11704
rect 3528 10606 3556 11698
rect 3516 10600 3568 10606
rect 3516 10542 3568 10548
rect 3528 9926 3556 10542
rect 3712 10130 3740 12038
rect 4220 11996 4516 12016
rect 4276 11994 4300 11996
rect 4356 11994 4380 11996
rect 4436 11994 4460 11996
rect 4298 11942 4300 11994
rect 4362 11942 4374 11994
rect 4436 11942 4438 11994
rect 4276 11940 4300 11942
rect 4356 11940 4380 11942
rect 4436 11940 4460 11942
rect 4220 11920 4516 11940
rect 4896 11688 4948 11694
rect 4896 11630 4948 11636
rect 4220 10908 4516 10928
rect 4276 10906 4300 10908
rect 4356 10906 4380 10908
rect 4436 10906 4460 10908
rect 4298 10854 4300 10906
rect 4362 10854 4374 10906
rect 4436 10854 4438 10906
rect 4276 10852 4300 10854
rect 4356 10852 4380 10854
rect 4436 10852 4460 10854
rect 4220 10832 4516 10852
rect 4908 10810 4936 11630
rect 5552 11218 5580 12242
rect 5736 11218 5764 16594
rect 6184 16040 6236 16046
rect 6184 15982 6236 15988
rect 6000 15972 6052 15978
rect 6000 15914 6052 15920
rect 6012 13870 6040 15914
rect 6000 13864 6052 13870
rect 6000 13806 6052 13812
rect 6196 12986 6224 15982
rect 6460 14408 6512 14414
rect 6460 14350 6512 14356
rect 6472 14006 6500 14350
rect 6564 14278 6592 16594
rect 6840 15502 6868 17138
rect 7104 16176 7156 16182
rect 7104 16118 7156 16124
rect 6828 15496 6880 15502
rect 6828 15438 6880 15444
rect 7116 15026 7144 16118
rect 7208 15706 7236 17614
rect 7288 16652 7340 16658
rect 7288 16594 7340 16600
rect 7196 15700 7248 15706
rect 7196 15642 7248 15648
rect 7104 15020 7156 15026
rect 7104 14962 7156 14968
rect 6828 14952 6880 14958
rect 6880 14912 6960 14940
rect 6828 14894 6880 14900
rect 6932 14822 6960 14912
rect 6736 14816 6788 14822
rect 6736 14758 6788 14764
rect 6920 14816 6972 14822
rect 6920 14758 6972 14764
rect 6552 14272 6604 14278
rect 6552 14214 6604 14220
rect 6460 14000 6512 14006
rect 6460 13942 6512 13948
rect 6748 13938 6776 14758
rect 6932 14482 6960 14758
rect 6920 14476 6972 14482
rect 6920 14418 6972 14424
rect 6736 13932 6788 13938
rect 6736 13874 6788 13880
rect 6184 12980 6236 12986
rect 6184 12922 6236 12928
rect 6196 12374 6224 12922
rect 6748 12374 6776 13874
rect 6932 12850 6960 14418
rect 7300 13870 7328 16594
rect 7392 16046 7420 17682
rect 7564 17128 7616 17134
rect 7564 17070 7616 17076
rect 7576 16726 7604 17070
rect 7564 16720 7616 16726
rect 7564 16662 7616 16668
rect 7380 16040 7432 16046
rect 7380 15982 7432 15988
rect 7564 16040 7616 16046
rect 7564 15982 7616 15988
rect 7576 15502 7604 15982
rect 7944 15638 7972 17682
rect 8116 16584 8168 16590
rect 8116 16526 8168 16532
rect 7932 15632 7984 15638
rect 7932 15574 7984 15580
rect 7564 15496 7616 15502
rect 7564 15438 7616 15444
rect 7576 14958 7604 15438
rect 7564 14952 7616 14958
rect 7564 14894 7616 14900
rect 7748 14272 7800 14278
rect 7748 14214 7800 14220
rect 7760 13938 7788 14214
rect 7748 13932 7800 13938
rect 7748 13874 7800 13880
rect 7288 13864 7340 13870
rect 7288 13806 7340 13812
rect 7300 13530 7328 13806
rect 7288 13524 7340 13530
rect 7288 13466 7340 13472
rect 7760 13462 7788 13874
rect 8128 13530 8156 16526
rect 8208 16040 8260 16046
rect 8208 15982 8260 15988
rect 8220 15638 8248 15982
rect 8208 15632 8260 15638
rect 8208 15574 8260 15580
rect 8404 15570 8432 18226
rect 8588 17610 8616 19246
rect 9048 18970 9076 19246
rect 9876 19174 9904 21082
rect 9968 21010 9996 22034
rect 9956 21004 10008 21010
rect 9956 20946 10008 20952
rect 9956 20596 10008 20602
rect 9956 20538 10008 20544
rect 9968 19922 9996 20538
rect 10232 20460 10284 20466
rect 10232 20402 10284 20408
rect 10140 20256 10192 20262
rect 10140 20198 10192 20204
rect 10152 20058 10180 20198
rect 10140 20052 10192 20058
rect 10140 19994 10192 20000
rect 9956 19916 10008 19922
rect 9956 19858 10008 19864
rect 10244 19786 10272 20402
rect 10232 19780 10284 19786
rect 10232 19722 10284 19728
rect 9864 19168 9916 19174
rect 9864 19110 9916 19116
rect 9036 18964 9088 18970
rect 9036 18906 9088 18912
rect 10244 18766 10272 19722
rect 10232 18760 10284 18766
rect 9494 18728 9550 18737
rect 10232 18702 10284 18708
rect 9494 18663 9550 18672
rect 9404 18148 9456 18154
rect 9404 18090 9456 18096
rect 8852 17740 8904 17746
rect 8852 17682 8904 17688
rect 8576 17604 8628 17610
rect 8576 17546 8628 17552
rect 8588 17134 8616 17546
rect 8864 17338 8892 17682
rect 8852 17332 8904 17338
rect 8852 17274 8904 17280
rect 9036 17332 9088 17338
rect 9036 17274 9088 17280
rect 8576 17128 8628 17134
rect 8576 17070 8628 17076
rect 9048 16726 9076 17274
rect 9036 16720 9088 16726
rect 9036 16662 9088 16668
rect 9048 16046 9076 16662
rect 9128 16584 9180 16590
rect 9128 16526 9180 16532
rect 9140 16114 9168 16526
rect 9128 16108 9180 16114
rect 9128 16050 9180 16056
rect 9416 16046 9444 18090
rect 9508 17864 9536 18663
rect 10244 18426 10272 18702
rect 10232 18420 10284 18426
rect 10232 18362 10284 18368
rect 10232 18216 10284 18222
rect 10232 18158 10284 18164
rect 9588 17876 9640 17882
rect 9508 17836 9588 17864
rect 9588 17818 9640 17824
rect 10048 16652 10100 16658
rect 10048 16594 10100 16600
rect 10060 16454 10088 16594
rect 10048 16448 10100 16454
rect 10048 16390 10100 16396
rect 9036 16040 9088 16046
rect 9036 15982 9088 15988
rect 9404 16040 9456 16046
rect 9404 15982 9456 15988
rect 8392 15564 8444 15570
rect 8392 15506 8444 15512
rect 8208 15360 8260 15366
rect 8208 15302 8260 15308
rect 8220 13870 8248 15302
rect 8404 15162 8432 15506
rect 9416 15162 9444 15982
rect 8392 15156 8444 15162
rect 8392 15098 8444 15104
rect 9220 15156 9272 15162
rect 9220 15098 9272 15104
rect 9404 15156 9456 15162
rect 9404 15098 9456 15104
rect 8852 14952 8904 14958
rect 8852 14894 8904 14900
rect 8760 14272 8812 14278
rect 8760 14214 8812 14220
rect 8772 13870 8800 14214
rect 8208 13864 8260 13870
rect 8208 13806 8260 13812
rect 8760 13864 8812 13870
rect 8760 13806 8812 13812
rect 8116 13524 8168 13530
rect 8116 13466 8168 13472
rect 7748 13456 7800 13462
rect 7748 13398 7800 13404
rect 8128 13326 8156 13466
rect 7104 13320 7156 13326
rect 7104 13262 7156 13268
rect 7380 13320 7432 13326
rect 7380 13262 7432 13268
rect 8116 13320 8168 13326
rect 8116 13262 8168 13268
rect 6920 12844 6972 12850
rect 6920 12786 6972 12792
rect 6184 12368 6236 12374
rect 6184 12310 6236 12316
rect 6736 12368 6788 12374
rect 6736 12310 6788 12316
rect 6276 12300 6328 12306
rect 6276 12242 6328 12248
rect 5540 11212 5592 11218
rect 5724 11212 5776 11218
rect 5592 11172 5672 11200
rect 5540 11154 5592 11160
rect 5540 11076 5592 11082
rect 5540 11018 5592 11024
rect 4896 10804 4948 10810
rect 4896 10746 4948 10752
rect 4620 10668 4672 10674
rect 4620 10610 4672 10616
rect 3792 10600 3844 10606
rect 3792 10542 3844 10548
rect 3700 10124 3752 10130
rect 3700 10066 3752 10072
rect 3516 9920 3568 9926
rect 3516 9862 3568 9868
rect 3804 9722 3832 10542
rect 4632 10062 4660 10610
rect 5552 10130 5580 11018
rect 5644 10130 5672 11172
rect 6288 11200 6316 12242
rect 6932 11694 6960 12786
rect 7012 12368 7064 12374
rect 7012 12310 7064 12316
rect 7116 12322 7144 13262
rect 7288 13252 7340 13258
rect 7288 13194 7340 13200
rect 7300 12850 7328 13194
rect 7288 12844 7340 12850
rect 7288 12786 7340 12792
rect 6920 11688 6972 11694
rect 6920 11630 6972 11636
rect 7024 11286 7052 12310
rect 7116 12306 7236 12322
rect 7116 12300 7248 12306
rect 7116 12294 7196 12300
rect 7196 12242 7248 12248
rect 7104 12232 7156 12238
rect 7104 12174 7156 12180
rect 7116 11762 7144 12174
rect 7104 11756 7156 11762
rect 7104 11698 7156 11704
rect 7012 11280 7064 11286
rect 7012 11222 7064 11228
rect 6368 11212 6420 11218
rect 6288 11172 6368 11200
rect 5724 11154 5776 11160
rect 6368 11154 6420 11160
rect 6000 11144 6052 11150
rect 6000 11086 6052 11092
rect 6012 10810 6040 11086
rect 6000 10804 6052 10810
rect 6000 10746 6052 10752
rect 5908 10600 5960 10606
rect 5908 10542 5960 10548
rect 5920 10266 5948 10542
rect 5908 10260 5960 10266
rect 5908 10202 5960 10208
rect 6380 10198 6408 11154
rect 7024 10266 7052 11222
rect 7196 11212 7248 11218
rect 7196 11154 7248 11160
rect 7104 10600 7156 10606
rect 7104 10542 7156 10548
rect 7012 10260 7064 10266
rect 7012 10202 7064 10208
rect 6368 10192 6420 10198
rect 6368 10134 6420 10140
rect 5540 10124 5592 10130
rect 5540 10066 5592 10072
rect 5632 10124 5684 10130
rect 5632 10066 5684 10072
rect 4620 10056 4672 10062
rect 4620 9998 4672 10004
rect 5356 10056 5408 10062
rect 5356 9998 5408 10004
rect 4220 9820 4516 9840
rect 4276 9818 4300 9820
rect 4356 9818 4380 9820
rect 4436 9818 4460 9820
rect 4298 9766 4300 9818
rect 4362 9766 4374 9818
rect 4436 9766 4438 9818
rect 4276 9764 4300 9766
rect 4356 9764 4380 9766
rect 4436 9764 4460 9766
rect 4220 9744 4516 9764
rect 3792 9716 3844 9722
rect 3792 9658 3844 9664
rect 4068 9580 4120 9586
rect 4068 9522 4120 9528
rect 4080 9353 4108 9522
rect 4632 9518 4660 9998
rect 4620 9512 4672 9518
rect 4620 9454 4672 9460
rect 4896 9512 4948 9518
rect 4896 9454 4948 9460
rect 4066 9344 4122 9353
rect 4066 9279 4122 9288
rect 4632 9058 4660 9454
rect 4068 9036 4120 9042
rect 4632 9030 4752 9058
rect 4068 8978 4120 8984
rect 4080 8430 4108 8978
rect 4620 8968 4672 8974
rect 4620 8910 4672 8916
rect 4220 8732 4516 8752
rect 4276 8730 4300 8732
rect 4356 8730 4380 8732
rect 4436 8730 4460 8732
rect 4298 8678 4300 8730
rect 4362 8678 4374 8730
rect 4436 8678 4438 8730
rect 4276 8676 4300 8678
rect 4356 8676 4380 8678
rect 4436 8676 4460 8678
rect 4220 8656 4516 8676
rect 3608 8424 3660 8430
rect 3608 8366 3660 8372
rect 4068 8424 4120 8430
rect 4068 8366 4120 8372
rect 3424 8356 3476 8362
rect 3424 8298 3476 8304
rect 3240 8084 3292 8090
rect 3240 8026 3292 8032
rect 3056 7880 3108 7886
rect 3056 7822 3108 7828
rect 2964 7540 3016 7546
rect 2964 7482 3016 7488
rect 3252 7410 3280 8026
rect 3240 7404 3292 7410
rect 3240 7346 3292 7352
rect 2780 7336 2832 7342
rect 2780 7278 2832 7284
rect 3620 6866 3648 8366
rect 4632 7954 4660 8910
rect 4724 7954 4752 9030
rect 4908 8974 4936 9454
rect 5368 9042 5396 9998
rect 5632 9580 5684 9586
rect 5632 9522 5684 9528
rect 5172 9036 5224 9042
rect 5172 8978 5224 8984
rect 5356 9036 5408 9042
rect 5356 8978 5408 8984
rect 4896 8968 4948 8974
rect 4896 8910 4948 8916
rect 4620 7948 4672 7954
rect 4620 7890 4672 7896
rect 4712 7948 4764 7954
rect 4712 7890 4764 7896
rect 3792 7880 3844 7886
rect 3792 7822 3844 7828
rect 3804 7342 3832 7822
rect 4068 7744 4120 7750
rect 4068 7686 4120 7692
rect 4080 7410 4108 7686
rect 4220 7644 4516 7664
rect 4276 7642 4300 7644
rect 4356 7642 4380 7644
rect 4436 7642 4460 7644
rect 4298 7590 4300 7642
rect 4362 7590 4374 7642
rect 4436 7590 4438 7642
rect 4276 7588 4300 7590
rect 4356 7588 4380 7590
rect 4436 7588 4460 7590
rect 4220 7568 4516 7588
rect 4068 7404 4120 7410
rect 4068 7346 4120 7352
rect 3792 7336 3844 7342
rect 3792 7278 3844 7284
rect 2412 6860 2464 6866
rect 2412 6802 2464 6808
rect 2504 6860 2556 6866
rect 2504 6802 2556 6808
rect 3608 6860 3660 6866
rect 3608 6802 3660 6808
rect 2424 6322 2452 6802
rect 2412 6316 2464 6322
rect 2412 6258 2464 6264
rect 2516 5914 2544 6802
rect 2964 6724 3016 6730
rect 2964 6666 3016 6672
rect 2504 5908 2556 5914
rect 2504 5850 2556 5856
rect 2976 5234 3004 6666
rect 3620 6390 3648 6802
rect 3608 6384 3660 6390
rect 3608 6326 3660 6332
rect 3332 6248 3384 6254
rect 3332 6190 3384 6196
rect 3148 6112 3200 6118
rect 3148 6054 3200 6060
rect 2964 5228 3016 5234
rect 2964 5170 3016 5176
rect 3160 5166 3188 6054
rect 3344 5778 3372 6190
rect 3620 6186 3648 6326
rect 3608 6180 3660 6186
rect 3608 6122 3660 6128
rect 3804 6118 3832 7278
rect 4724 6798 4752 7890
rect 5184 7546 5212 8978
rect 5644 7954 5672 9522
rect 6380 9042 6408 10134
rect 6368 9036 6420 9042
rect 6368 8978 6420 8984
rect 6920 9036 6972 9042
rect 7024 9024 7052 10202
rect 7116 10062 7144 10542
rect 7104 10056 7156 10062
rect 7104 9998 7156 10004
rect 7208 9450 7236 11154
rect 7392 9518 7420 13262
rect 8024 12708 8076 12714
rect 8024 12650 8076 12656
rect 8036 12306 8064 12650
rect 8220 12374 8248 13806
rect 8300 13388 8352 13394
rect 8300 13330 8352 13336
rect 8208 12368 8260 12374
rect 8208 12310 8260 12316
rect 7840 12300 7892 12306
rect 7840 12242 7892 12248
rect 8024 12300 8076 12306
rect 8024 12242 8076 12248
rect 7852 11354 7880 12242
rect 7840 11348 7892 11354
rect 7840 11290 7892 11296
rect 8036 9654 8064 12242
rect 8312 12238 8340 13330
rect 8484 12640 8536 12646
rect 8484 12582 8536 12588
rect 8300 12232 8352 12238
rect 8300 12174 8352 12180
rect 8496 11898 8524 12582
rect 8760 12300 8812 12306
rect 8864 12288 8892 14894
rect 9232 14822 9260 15098
rect 9772 14952 9824 14958
rect 9772 14894 9824 14900
rect 9404 14884 9456 14890
rect 9324 14844 9404 14872
rect 9220 14816 9272 14822
rect 9220 14758 9272 14764
rect 9036 14408 9088 14414
rect 9088 14368 9168 14396
rect 9036 14350 9088 14356
rect 9140 12782 9168 14368
rect 9232 13870 9260 14758
rect 9324 13920 9352 14844
rect 9404 14826 9456 14832
rect 9494 14648 9550 14657
rect 9494 14583 9496 14592
rect 9548 14583 9550 14592
rect 9496 14554 9548 14560
rect 9784 14414 9812 14894
rect 10060 14482 10088 16390
rect 9956 14476 10008 14482
rect 9956 14418 10008 14424
rect 10048 14476 10100 14482
rect 10048 14418 10100 14424
rect 9772 14408 9824 14414
rect 9772 14350 9824 14356
rect 9968 14074 9996 14418
rect 9956 14068 10008 14074
rect 9956 14010 10008 14016
rect 9404 13932 9456 13938
rect 9324 13892 9404 13920
rect 9404 13874 9456 13880
rect 9220 13864 9272 13870
rect 9220 13806 9272 13812
rect 9680 13524 9732 13530
rect 9680 13466 9732 13472
rect 9128 12776 9180 12782
rect 9128 12718 9180 12724
rect 8812 12260 8892 12288
rect 8760 12242 8812 12248
rect 8484 11892 8536 11898
rect 8484 11834 8536 11840
rect 8392 11552 8444 11558
rect 8392 11494 8444 11500
rect 8404 11218 8432 11494
rect 8392 11212 8444 11218
rect 8392 11154 8444 11160
rect 8484 11212 8536 11218
rect 8484 11154 8536 11160
rect 8024 9648 8076 9654
rect 8024 9590 8076 9596
rect 7380 9512 7432 9518
rect 7380 9454 7432 9460
rect 7840 9512 7892 9518
rect 7840 9454 7892 9460
rect 7196 9444 7248 9450
rect 7196 9386 7248 9392
rect 6972 8996 7052 9024
rect 7196 9036 7248 9042
rect 6920 8978 6972 8984
rect 7196 8978 7248 8984
rect 6460 8356 6512 8362
rect 6460 8298 6512 8304
rect 6472 8090 6500 8298
rect 6460 8084 6512 8090
rect 6460 8026 6512 8032
rect 5632 7948 5684 7954
rect 5632 7890 5684 7896
rect 7208 7546 7236 8978
rect 7392 8294 7420 9454
rect 7748 9376 7800 9382
rect 7748 9318 7800 9324
rect 7760 9042 7788 9318
rect 7748 9036 7800 9042
rect 7748 8978 7800 8984
rect 7852 8498 7880 9454
rect 8496 9178 8524 11154
rect 8576 9512 8628 9518
rect 8576 9454 8628 9460
rect 8588 9178 8616 9454
rect 8484 9172 8536 9178
rect 8484 9114 8536 9120
rect 8576 9172 8628 9178
rect 8576 9114 8628 9120
rect 8576 8832 8628 8838
rect 8576 8774 8628 8780
rect 7840 8492 7892 8498
rect 7840 8434 7892 8440
rect 8392 8492 8444 8498
rect 8392 8434 8444 8440
rect 8024 8356 8076 8362
rect 8024 8298 8076 8304
rect 7380 8288 7432 8294
rect 7380 8230 7432 8236
rect 5172 7540 5224 7546
rect 5172 7482 5224 7488
rect 7196 7540 7248 7546
rect 7196 7482 7248 7488
rect 5184 6934 5212 7482
rect 7288 7472 7340 7478
rect 7288 7414 7340 7420
rect 5172 6928 5224 6934
rect 5172 6870 5224 6876
rect 5080 6860 5132 6866
rect 5080 6802 5132 6808
rect 4620 6792 4672 6798
rect 4620 6734 4672 6740
rect 4712 6792 4764 6798
rect 4712 6734 4764 6740
rect 4220 6556 4516 6576
rect 4276 6554 4300 6556
rect 4356 6554 4380 6556
rect 4436 6554 4460 6556
rect 4298 6502 4300 6554
rect 4362 6502 4374 6554
rect 4436 6502 4438 6554
rect 4276 6500 4300 6502
rect 4356 6500 4380 6502
rect 4436 6500 4460 6502
rect 4220 6480 4516 6500
rect 3974 6352 4030 6361
rect 3974 6287 4030 6296
rect 3792 6112 3844 6118
rect 3792 6054 3844 6060
rect 3988 5846 4016 6287
rect 4160 6248 4212 6254
rect 4160 6190 4212 6196
rect 3976 5840 4028 5846
rect 3976 5782 4028 5788
rect 4172 5778 4200 6190
rect 4528 6180 4580 6186
rect 4528 6122 4580 6128
rect 3332 5772 3384 5778
rect 3332 5714 3384 5720
rect 4160 5772 4212 5778
rect 4160 5714 4212 5720
rect 3344 5370 3372 5714
rect 4540 5642 4568 6122
rect 4528 5636 4580 5642
rect 4528 5578 4580 5584
rect 4220 5468 4516 5488
rect 4276 5466 4300 5468
rect 4356 5466 4380 5468
rect 4436 5466 4460 5468
rect 4298 5414 4300 5466
rect 4362 5414 4374 5466
rect 4436 5414 4438 5466
rect 4276 5412 4300 5414
rect 4356 5412 4380 5414
rect 4436 5412 4460 5414
rect 4220 5392 4516 5412
rect 3332 5364 3384 5370
rect 3332 5306 3384 5312
rect 3148 5160 3200 5166
rect 3148 5102 3200 5108
rect 572 3528 624 3534
rect 572 3470 624 3476
rect 1768 3528 1820 3534
rect 1768 3470 1820 3476
rect 584 800 612 3470
rect 3160 2990 3188 5102
rect 4528 5024 4580 5030
rect 4528 4966 4580 4972
rect 4540 4690 4568 4966
rect 4528 4684 4580 4690
rect 4528 4626 4580 4632
rect 4220 4380 4516 4400
rect 4276 4378 4300 4380
rect 4356 4378 4380 4380
rect 4436 4378 4460 4380
rect 4298 4326 4300 4378
rect 4362 4326 4374 4378
rect 4436 4326 4438 4378
rect 4276 4324 4300 4326
rect 4356 4324 4380 4326
rect 4436 4324 4460 4326
rect 4220 4304 4516 4324
rect 4632 4078 4660 6734
rect 5092 6458 5120 6802
rect 5080 6452 5132 6458
rect 5080 6394 5132 6400
rect 4896 6248 4948 6254
rect 4896 6190 4948 6196
rect 4712 5704 4764 5710
rect 4712 5646 4764 5652
rect 4724 5234 4752 5646
rect 4804 5636 4856 5642
rect 4804 5578 4856 5584
rect 4712 5228 4764 5234
rect 4712 5170 4764 5176
rect 4620 4072 4672 4078
rect 4620 4014 4672 4020
rect 4724 4010 4752 5170
rect 4816 4146 4844 5578
rect 4908 4146 4936 6190
rect 4988 5772 5040 5778
rect 4988 5714 5040 5720
rect 5000 4622 5028 5714
rect 5092 5302 5120 6394
rect 5080 5296 5132 5302
rect 5080 5238 5132 5244
rect 5184 5234 5212 6870
rect 7300 6866 7328 7414
rect 7392 7342 7420 8230
rect 8036 7954 8064 8298
rect 8404 7954 8432 8434
rect 8588 8430 8616 8774
rect 8772 8498 8800 12242
rect 9140 11558 9168 12718
rect 9692 11898 9720 13466
rect 9864 12844 9916 12850
rect 9864 12786 9916 12792
rect 9680 11892 9732 11898
rect 9680 11834 9732 11840
rect 9876 11694 9904 12786
rect 10060 12442 10088 14418
rect 10140 13388 10192 13394
rect 10140 13330 10192 13336
rect 10048 12436 10100 12442
rect 10048 12378 10100 12384
rect 10152 12238 10180 13330
rect 10140 12232 10192 12238
rect 10140 12174 10192 12180
rect 9864 11688 9916 11694
rect 9864 11630 9916 11636
rect 10140 11688 10192 11694
rect 10140 11630 10192 11636
rect 9128 11552 9180 11558
rect 9128 11494 9180 11500
rect 9680 11212 9732 11218
rect 9680 11154 9732 11160
rect 9312 10600 9364 10606
rect 9312 10542 9364 10548
rect 8944 10532 8996 10538
rect 8944 10474 8996 10480
rect 8852 10464 8904 10470
rect 8852 10406 8904 10412
rect 8864 9382 8892 10406
rect 8956 10130 8984 10474
rect 8944 10124 8996 10130
rect 8944 10066 8996 10072
rect 9324 9722 9352 10542
rect 9692 10130 9720 11154
rect 10152 11082 10180 11630
rect 10140 11076 10192 11082
rect 10140 11018 10192 11024
rect 9864 10600 9916 10606
rect 9864 10542 9916 10548
rect 9772 10260 9824 10266
rect 9772 10202 9824 10208
rect 9680 10124 9732 10130
rect 9680 10066 9732 10072
rect 9312 9716 9364 9722
rect 9312 9658 9364 9664
rect 9784 9518 9812 10202
rect 9772 9512 9824 9518
rect 9772 9454 9824 9460
rect 9496 9444 9548 9450
rect 9496 9386 9548 9392
rect 8852 9376 8904 9382
rect 8852 9318 8904 9324
rect 8760 8492 8812 8498
rect 8760 8434 8812 8440
rect 8576 8424 8628 8430
rect 8576 8366 8628 8372
rect 8024 7948 8076 7954
rect 8024 7890 8076 7896
rect 8392 7948 8444 7954
rect 8392 7890 8444 7896
rect 7656 7880 7708 7886
rect 7656 7822 7708 7828
rect 7668 7342 7696 7822
rect 7840 7744 7892 7750
rect 7840 7686 7892 7692
rect 7380 7336 7432 7342
rect 7380 7278 7432 7284
rect 7656 7336 7708 7342
rect 7656 7278 7708 7284
rect 7852 7002 7880 7686
rect 8036 7274 8064 7890
rect 8024 7268 8076 7274
rect 8024 7210 8076 7216
rect 7840 6996 7892 7002
rect 7840 6938 7892 6944
rect 5356 6860 5408 6866
rect 5356 6802 5408 6808
rect 7288 6860 7340 6866
rect 7288 6802 7340 6808
rect 5264 6112 5316 6118
rect 5264 6054 5316 6060
rect 5276 5778 5304 6054
rect 5264 5772 5316 5778
rect 5264 5714 5316 5720
rect 5368 5574 5396 6802
rect 6276 6792 6328 6798
rect 6276 6734 6328 6740
rect 6288 6322 6316 6734
rect 8588 6322 8616 8366
rect 6276 6316 6328 6322
rect 6276 6258 6328 6264
rect 8300 6316 8352 6322
rect 8300 6258 8352 6264
rect 8576 6316 8628 6322
rect 8576 6258 8628 6264
rect 8208 6248 8260 6254
rect 8208 6190 8260 6196
rect 8220 5914 8248 6190
rect 8208 5908 8260 5914
rect 8208 5850 8260 5856
rect 6276 5704 6328 5710
rect 6276 5646 6328 5652
rect 5356 5568 5408 5574
rect 5356 5510 5408 5516
rect 5172 5228 5224 5234
rect 5172 5170 5224 5176
rect 5184 5098 5212 5170
rect 5368 5166 5396 5510
rect 5356 5160 5408 5166
rect 5356 5102 5408 5108
rect 5172 5092 5224 5098
rect 5172 5034 5224 5040
rect 5184 4690 5212 5034
rect 5368 5030 5396 5102
rect 5356 5024 5408 5030
rect 5356 4966 5408 4972
rect 5816 5024 5868 5030
rect 5816 4966 5868 4972
rect 5172 4684 5224 4690
rect 5172 4626 5224 4632
rect 4988 4616 5040 4622
rect 4988 4558 5040 4564
rect 4804 4140 4856 4146
rect 4804 4082 4856 4088
rect 4896 4140 4948 4146
rect 4896 4082 4948 4088
rect 5000 4010 5028 4558
rect 5828 4078 5856 4966
rect 6288 4146 6316 5646
rect 8312 5234 8340 6258
rect 8300 5228 8352 5234
rect 8300 5170 8352 5176
rect 6828 4616 6880 4622
rect 6828 4558 6880 4564
rect 6276 4140 6328 4146
rect 6276 4082 6328 4088
rect 5816 4072 5868 4078
rect 5816 4014 5868 4020
rect 6840 4010 6868 4558
rect 7564 4480 7616 4486
rect 7564 4422 7616 4428
rect 7576 4078 7604 4422
rect 7564 4072 7616 4078
rect 7564 4014 7616 4020
rect 8484 4072 8536 4078
rect 8484 4014 8536 4020
rect 8760 4072 8812 4078
rect 8760 4014 8812 4020
rect 4712 4004 4764 4010
rect 4712 3946 4764 3952
rect 4988 4004 5040 4010
rect 4988 3946 5040 3952
rect 6828 4004 6880 4010
rect 6828 3946 6880 3952
rect 7748 4004 7800 4010
rect 7748 3946 7800 3952
rect 3422 3632 3478 3641
rect 6840 3602 6868 3946
rect 7472 3936 7524 3942
rect 7472 3878 7524 3884
rect 7484 3602 7512 3878
rect 3422 3567 3478 3576
rect 6828 3596 6880 3602
rect 3148 2984 3200 2990
rect 3148 2926 3200 2932
rect 3160 2514 3188 2926
rect 3436 2650 3464 3567
rect 6828 3538 6880 3544
rect 7472 3596 7524 3602
rect 7472 3538 7524 3544
rect 6274 3360 6330 3369
rect 4220 3292 4516 3312
rect 6274 3295 6330 3304
rect 4276 3290 4300 3292
rect 4356 3290 4380 3292
rect 4436 3290 4460 3292
rect 4298 3238 4300 3290
rect 4362 3238 4374 3290
rect 4436 3238 4438 3290
rect 4276 3236 4300 3238
rect 4356 3236 4380 3238
rect 4436 3236 4460 3238
rect 4220 3216 4516 3236
rect 4620 2848 4672 2854
rect 4620 2790 4672 2796
rect 3424 2644 3476 2650
rect 3424 2586 3476 2592
rect 3148 2508 3200 2514
rect 3148 2450 3200 2456
rect 2412 2304 2464 2310
rect 2412 2246 2464 2252
rect 2424 800 2452 2246
rect 4220 2204 4516 2224
rect 4276 2202 4300 2204
rect 4356 2202 4380 2204
rect 4436 2202 4460 2204
rect 4298 2150 4300 2202
rect 4362 2150 4374 2202
rect 4436 2150 4438 2202
rect 4276 2148 4300 2150
rect 4356 2148 4380 2150
rect 4436 2148 4460 2150
rect 4220 2128 4516 2148
rect 4632 1442 4660 2790
rect 4264 1414 4660 1442
rect 4264 800 4292 1414
rect 6288 800 6316 3295
rect 7288 2984 7340 2990
rect 7286 2952 7288 2961
rect 7340 2952 7342 2961
rect 7286 2887 7342 2896
rect 7760 2514 7788 3946
rect 8114 3496 8170 3505
rect 8114 3431 8170 3440
rect 8024 3188 8076 3194
rect 8024 3130 8076 3136
rect 8036 3058 8064 3130
rect 8024 3052 8076 3058
rect 8024 2994 8076 3000
rect 7748 2508 7800 2514
rect 7748 2450 7800 2456
rect 8128 800 8156 3431
rect 8496 3126 8524 4014
rect 8772 3670 8800 4014
rect 8760 3664 8812 3670
rect 8760 3606 8812 3612
rect 8668 3460 8720 3466
rect 8668 3402 8720 3408
rect 8484 3120 8536 3126
rect 8484 3062 8536 3068
rect 8680 2990 8708 3402
rect 8864 2990 8892 9318
rect 9312 7948 9364 7954
rect 9312 7890 9364 7896
rect 9324 7342 9352 7890
rect 9312 7336 9364 7342
rect 9312 7278 9364 7284
rect 9508 6866 9536 9386
rect 9876 9110 9904 10542
rect 9956 10192 10008 10198
rect 9956 10134 10008 10140
rect 9864 9104 9916 9110
rect 9864 9046 9916 9052
rect 9864 8968 9916 8974
rect 9864 8910 9916 8916
rect 9876 8498 9904 8910
rect 9864 8492 9916 8498
rect 9864 8434 9916 8440
rect 9680 8424 9732 8430
rect 9876 8378 9904 8434
rect 9680 8366 9732 8372
rect 9692 7818 9720 8366
rect 9784 8350 9904 8378
rect 9680 7812 9732 7818
rect 9680 7754 9732 7760
rect 9784 7410 9812 8350
rect 9864 7948 9916 7954
rect 9968 7936 9996 10134
rect 10048 10124 10100 10130
rect 10048 10066 10100 10072
rect 10060 9625 10088 10066
rect 10046 9616 10102 9625
rect 10046 9551 10102 9560
rect 10152 9518 10180 11018
rect 10140 9512 10192 9518
rect 10140 9454 10192 9460
rect 10152 9382 10180 9454
rect 10140 9376 10192 9382
rect 10140 9318 10192 9324
rect 10048 8288 10100 8294
rect 10048 8230 10100 8236
rect 10060 7954 10088 8230
rect 9916 7908 9996 7936
rect 10048 7948 10100 7954
rect 9864 7890 9916 7896
rect 10048 7890 10100 7896
rect 9876 7857 9904 7890
rect 9862 7848 9918 7857
rect 9862 7783 9918 7792
rect 9956 7472 10008 7478
rect 9956 7414 10008 7420
rect 9772 7404 9824 7410
rect 9772 7346 9824 7352
rect 9496 6860 9548 6866
rect 9496 6802 9548 6808
rect 9508 6458 9536 6802
rect 9496 6452 9548 6458
rect 9496 6394 9548 6400
rect 9968 5778 9996 7414
rect 10244 7002 10272 18158
rect 10336 17542 10364 36654
rect 10598 36615 10654 36624
rect 10416 35624 10468 35630
rect 10416 35566 10468 35572
rect 10428 35290 10456 35566
rect 10416 35284 10468 35290
rect 10416 35226 10468 35232
rect 10416 33516 10468 33522
rect 10416 33458 10468 33464
rect 10428 33318 10456 33458
rect 10416 33312 10468 33318
rect 10416 33254 10468 33260
rect 10428 32978 10456 33254
rect 10416 32972 10468 32978
rect 10416 32914 10468 32920
rect 10416 32768 10468 32774
rect 10416 32710 10468 32716
rect 10428 32298 10456 32710
rect 10416 32292 10468 32298
rect 10416 32234 10468 32240
rect 10428 31822 10456 32234
rect 10508 31884 10560 31890
rect 10508 31826 10560 31832
rect 10416 31816 10468 31822
rect 10416 31758 10468 31764
rect 10520 30258 10548 31826
rect 10692 31272 10744 31278
rect 10692 31214 10744 31220
rect 10704 30802 10732 31214
rect 10692 30796 10744 30802
rect 10692 30738 10744 30744
rect 10508 30252 10560 30258
rect 10508 30194 10560 30200
rect 10506 29744 10562 29753
rect 10704 29714 10732 30738
rect 10506 29679 10508 29688
rect 10560 29679 10562 29688
rect 10692 29708 10744 29714
rect 10508 29650 10560 29656
rect 10692 29650 10744 29656
rect 10704 29617 10732 29650
rect 10690 29608 10746 29617
rect 10690 29543 10746 29552
rect 10416 29096 10468 29102
rect 10416 29038 10468 29044
rect 10428 28762 10456 29038
rect 10416 28756 10468 28762
rect 10416 28698 10468 28704
rect 10508 28212 10560 28218
rect 10508 28154 10560 28160
rect 10520 26994 10548 28154
rect 10796 27996 10824 37284
rect 11072 36378 11100 37742
rect 12452 37262 12480 37810
rect 12808 37392 12860 37398
rect 12808 37334 12860 37340
rect 12440 37256 12492 37262
rect 12440 37198 12492 37204
rect 11152 36916 11204 36922
rect 11152 36858 11204 36864
rect 11164 36378 11192 36858
rect 12820 36718 12848 37334
rect 12912 36786 12940 38354
rect 14096 38276 14148 38282
rect 14096 38218 14148 38224
rect 13820 37800 13872 37806
rect 13820 37742 13872 37748
rect 12992 37392 13044 37398
rect 12992 37334 13044 37340
rect 12900 36780 12952 36786
rect 12900 36722 12952 36728
rect 11428 36712 11480 36718
rect 11428 36654 11480 36660
rect 12808 36712 12860 36718
rect 12808 36654 12860 36660
rect 11060 36372 11112 36378
rect 11060 36314 11112 36320
rect 11152 36372 11204 36378
rect 11152 36314 11204 36320
rect 11440 36242 11468 36654
rect 13004 36650 13032 37334
rect 13832 37330 13860 37742
rect 13084 37324 13136 37330
rect 13084 37266 13136 37272
rect 13820 37324 13872 37330
rect 13820 37266 13872 37272
rect 12992 36644 13044 36650
rect 12992 36586 13044 36592
rect 12164 36576 12216 36582
rect 12164 36518 12216 36524
rect 12808 36576 12860 36582
rect 12808 36518 12860 36524
rect 11428 36236 11480 36242
rect 11428 36178 11480 36184
rect 12176 35766 12204 36518
rect 12820 36242 12848 36518
rect 13004 36242 13032 36586
rect 12808 36236 12860 36242
rect 12808 36178 12860 36184
rect 12992 36236 13044 36242
rect 12992 36178 13044 36184
rect 12164 35760 12216 35766
rect 12164 35702 12216 35708
rect 11152 35624 11204 35630
rect 11152 35566 11204 35572
rect 10968 35080 11020 35086
rect 10968 35022 11020 35028
rect 10980 34610 11008 35022
rect 10968 34604 11020 34610
rect 10968 34546 11020 34552
rect 11164 33998 11192 35566
rect 11244 35488 11296 35494
rect 11244 35430 11296 35436
rect 11256 35154 11284 35430
rect 11244 35148 11296 35154
rect 11244 35090 11296 35096
rect 11336 35148 11388 35154
rect 11336 35090 11388 35096
rect 11348 34542 11376 35090
rect 11336 34536 11388 34542
rect 11336 34478 11388 34484
rect 11704 34400 11756 34406
rect 11704 34342 11756 34348
rect 11716 33998 11744 34342
rect 11888 34060 11940 34066
rect 11888 34002 11940 34008
rect 11152 33992 11204 33998
rect 11152 33934 11204 33940
rect 11704 33992 11756 33998
rect 11704 33934 11756 33940
rect 11060 33924 11112 33930
rect 11060 33866 11112 33872
rect 11072 33386 11100 33866
rect 11520 33584 11572 33590
rect 11520 33526 11572 33532
rect 11152 33448 11204 33454
rect 11152 33390 11204 33396
rect 11060 33380 11112 33386
rect 11060 33322 11112 33328
rect 11060 32972 11112 32978
rect 11164 32960 11192 33390
rect 11112 32932 11192 32960
rect 11060 32914 11112 32920
rect 11072 32502 11100 32914
rect 11060 32496 11112 32502
rect 11060 32438 11112 32444
rect 10876 31884 10928 31890
rect 10876 31826 10928 31832
rect 10888 30190 10916 31826
rect 10968 30728 11020 30734
rect 10968 30670 11020 30676
rect 10876 30184 10928 30190
rect 10876 30126 10928 30132
rect 10876 29300 10928 29306
rect 10876 29242 10928 29248
rect 10612 27968 10824 27996
rect 10612 26994 10640 27968
rect 10784 27872 10836 27878
rect 10784 27814 10836 27820
rect 10508 26988 10560 26994
rect 10508 26930 10560 26936
rect 10600 26988 10652 26994
rect 10600 26930 10652 26936
rect 10600 26784 10652 26790
rect 10600 26726 10652 26732
rect 10612 25906 10640 26726
rect 10692 26036 10744 26042
rect 10692 25978 10744 25984
rect 10600 25900 10652 25906
rect 10600 25842 10652 25848
rect 10612 25498 10640 25842
rect 10600 25492 10652 25498
rect 10600 25434 10652 25440
rect 10612 25362 10640 25434
rect 10600 25356 10652 25362
rect 10600 25298 10652 25304
rect 10704 25294 10732 25978
rect 10692 25288 10744 25294
rect 10692 25230 10744 25236
rect 10704 24614 10732 25230
rect 10692 24608 10744 24614
rect 10692 24550 10744 24556
rect 10508 23588 10560 23594
rect 10508 23530 10560 23536
rect 10520 23186 10548 23530
rect 10600 23316 10652 23322
rect 10600 23258 10652 23264
rect 10508 23180 10560 23186
rect 10508 23122 10560 23128
rect 10612 22642 10640 23258
rect 10600 22636 10652 22642
rect 10600 22578 10652 22584
rect 10416 22568 10468 22574
rect 10416 22510 10468 22516
rect 10428 22234 10456 22510
rect 10416 22228 10468 22234
rect 10416 22170 10468 22176
rect 10612 22098 10640 22578
rect 10600 22092 10652 22098
rect 10600 22034 10652 22040
rect 10796 21554 10824 27814
rect 10888 27606 10916 29242
rect 10980 28218 11008 30670
rect 11072 30190 11100 32438
rect 11532 32366 11560 33526
rect 11612 33380 11664 33386
rect 11612 33322 11664 33328
rect 11624 32978 11652 33322
rect 11716 33318 11744 33934
rect 11704 33312 11756 33318
rect 11704 33254 11756 33260
rect 11612 32972 11664 32978
rect 11612 32914 11664 32920
rect 11796 32904 11848 32910
rect 11796 32846 11848 32852
rect 11520 32360 11572 32366
rect 11520 32302 11572 32308
rect 11532 31346 11560 32302
rect 11808 32230 11836 32846
rect 11796 32224 11848 32230
rect 11796 32166 11848 32172
rect 11808 32026 11836 32166
rect 11796 32020 11848 32026
rect 11796 31962 11848 31968
rect 11520 31340 11572 31346
rect 11520 31282 11572 31288
rect 11152 31272 11204 31278
rect 11152 31214 11204 31220
rect 11704 31272 11756 31278
rect 11704 31214 11756 31220
rect 11164 30802 11192 31214
rect 11520 31204 11572 31210
rect 11520 31146 11572 31152
rect 11532 30802 11560 31146
rect 11716 30938 11744 31214
rect 11704 30932 11756 30938
rect 11704 30874 11756 30880
rect 11152 30796 11204 30802
rect 11152 30738 11204 30744
rect 11520 30796 11572 30802
rect 11520 30738 11572 30744
rect 11164 30326 11192 30738
rect 11152 30320 11204 30326
rect 11152 30262 11204 30268
rect 11808 30190 11836 31962
rect 11900 31142 11928 34002
rect 11980 32836 12032 32842
rect 11980 32778 12032 32784
rect 11992 31822 12020 32778
rect 11980 31816 12032 31822
rect 11980 31758 12032 31764
rect 11888 31136 11940 31142
rect 11888 31078 11940 31084
rect 11060 30184 11112 30190
rect 11060 30126 11112 30132
rect 11796 30184 11848 30190
rect 11796 30126 11848 30132
rect 11428 29776 11480 29782
rect 11428 29718 11480 29724
rect 11244 29708 11296 29714
rect 11244 29650 11296 29656
rect 11256 29306 11284 29650
rect 11336 29572 11388 29578
rect 11336 29514 11388 29520
rect 11244 29300 11296 29306
rect 11244 29242 11296 29248
rect 11348 28626 11376 29514
rect 11440 29306 11468 29718
rect 11796 29708 11848 29714
rect 11796 29650 11848 29656
rect 11808 29306 11836 29650
rect 11428 29300 11480 29306
rect 11428 29242 11480 29248
rect 11796 29300 11848 29306
rect 11796 29242 11848 29248
rect 11440 28642 11468 29242
rect 11440 28626 11560 28642
rect 11336 28620 11388 28626
rect 11336 28562 11388 28568
rect 11440 28620 11572 28626
rect 11440 28614 11520 28620
rect 10968 28212 11020 28218
rect 10968 28154 11020 28160
rect 10968 28076 11020 28082
rect 10968 28018 11020 28024
rect 10876 27600 10928 27606
rect 10876 27542 10928 27548
rect 10876 26988 10928 26994
rect 10876 26930 10928 26936
rect 10784 21548 10836 21554
rect 10784 21490 10836 21496
rect 10692 21480 10744 21486
rect 10888 21434 10916 26930
rect 10980 25770 11008 28018
rect 11440 28014 11468 28614
rect 11520 28562 11572 28568
rect 11428 28008 11480 28014
rect 11428 27950 11480 27956
rect 11336 27532 11388 27538
rect 11336 27474 11388 27480
rect 11060 27328 11112 27334
rect 11060 27270 11112 27276
rect 11072 26926 11100 27270
rect 11060 26920 11112 26926
rect 11060 26862 11112 26868
rect 11072 26246 11100 26862
rect 11348 26382 11376 27474
rect 11808 27470 11836 29242
rect 12072 27872 12124 27878
rect 12072 27814 12124 27820
rect 12084 27538 12112 27814
rect 12072 27532 12124 27538
rect 12072 27474 12124 27480
rect 11796 27464 11848 27470
rect 11796 27406 11848 27412
rect 11980 27396 12032 27402
rect 11980 27338 12032 27344
rect 11428 26920 11480 26926
rect 11428 26862 11480 26868
rect 11888 26920 11940 26926
rect 11888 26862 11940 26868
rect 11336 26376 11388 26382
rect 11336 26318 11388 26324
rect 11060 26240 11112 26246
rect 11060 26182 11112 26188
rect 10968 25764 11020 25770
rect 10968 25706 11020 25712
rect 11072 25498 11100 26182
rect 11440 26042 11468 26862
rect 11900 26586 11928 26862
rect 11992 26858 12020 27338
rect 11980 26852 12032 26858
rect 11980 26794 12032 26800
rect 11888 26580 11940 26586
rect 11888 26522 11940 26528
rect 12084 26450 12112 27474
rect 12072 26444 12124 26450
rect 12072 26386 12124 26392
rect 11428 26036 11480 26042
rect 11428 25978 11480 25984
rect 11336 25832 11388 25838
rect 11336 25774 11388 25780
rect 11060 25492 11112 25498
rect 11060 25434 11112 25440
rect 11244 25492 11296 25498
rect 11244 25434 11296 25440
rect 11152 25424 11204 25430
rect 11152 25366 11204 25372
rect 11060 25288 11112 25294
rect 11060 25230 11112 25236
rect 11072 24750 11100 25230
rect 11060 24744 11112 24750
rect 11060 24686 11112 24692
rect 11072 24274 11100 24686
rect 11164 24682 11192 25366
rect 11256 24750 11284 25434
rect 11244 24744 11296 24750
rect 11244 24686 11296 24692
rect 11152 24676 11204 24682
rect 11152 24618 11204 24624
rect 11164 24410 11192 24618
rect 11256 24614 11284 24686
rect 11348 24614 11376 25774
rect 11980 25696 12032 25702
rect 11980 25638 12032 25644
rect 11992 24682 12020 25638
rect 11980 24676 12032 24682
rect 11980 24618 12032 24624
rect 11244 24608 11296 24614
rect 11244 24550 11296 24556
rect 11336 24608 11388 24614
rect 11336 24550 11388 24556
rect 11152 24404 11204 24410
rect 11152 24346 11204 24352
rect 11992 24342 12020 24618
rect 11980 24336 12032 24342
rect 11980 24278 12032 24284
rect 11060 24268 11112 24274
rect 11244 24268 11296 24274
rect 11060 24210 11112 24216
rect 11164 24228 11244 24256
rect 11072 23526 11100 24210
rect 11164 23662 11192 24228
rect 11244 24210 11296 24216
rect 11888 24268 11940 24274
rect 11888 24210 11940 24216
rect 11900 23798 11928 24210
rect 11888 23792 11940 23798
rect 11888 23734 11940 23740
rect 11152 23656 11204 23662
rect 11152 23598 11204 23604
rect 12072 23656 12124 23662
rect 12072 23598 12124 23604
rect 11060 23520 11112 23526
rect 11060 23462 11112 23468
rect 11060 22568 11112 22574
rect 11164 22556 11192 23598
rect 12084 23186 12112 23598
rect 11428 23180 11480 23186
rect 11428 23122 11480 23128
rect 12072 23180 12124 23186
rect 12072 23122 12124 23128
rect 11440 22982 11468 23122
rect 11428 22976 11480 22982
rect 11428 22918 11480 22924
rect 11112 22528 11192 22556
rect 11060 22510 11112 22516
rect 11072 22098 11100 22510
rect 11440 22234 11468 22918
rect 11428 22228 11480 22234
rect 11428 22170 11480 22176
rect 11060 22092 11112 22098
rect 11060 22034 11112 22040
rect 12176 21962 12204 35702
rect 12532 34944 12584 34950
rect 12532 34886 12584 34892
rect 12624 34944 12676 34950
rect 12624 34886 12676 34892
rect 12544 33998 12572 34886
rect 12636 34542 12664 34886
rect 12624 34536 12676 34542
rect 12624 34478 12676 34484
rect 12716 34468 12768 34474
rect 12716 34410 12768 34416
rect 12728 34066 12756 34410
rect 12716 34060 12768 34066
rect 12716 34002 12768 34008
rect 12900 34060 12952 34066
rect 12900 34002 12952 34008
rect 12532 33992 12584 33998
rect 12532 33934 12584 33940
rect 12348 33924 12400 33930
rect 12348 33866 12400 33872
rect 12360 33522 12388 33866
rect 12348 33516 12400 33522
rect 12348 33458 12400 33464
rect 12912 33454 12940 34002
rect 13004 33862 13032 36178
rect 13096 36174 13124 37266
rect 13176 37120 13228 37126
rect 13176 37062 13228 37068
rect 13188 36718 13216 37062
rect 13176 36712 13228 36718
rect 13176 36654 13228 36660
rect 13084 36168 13136 36174
rect 13084 36110 13136 36116
rect 13268 35624 13320 35630
rect 13268 35566 13320 35572
rect 13636 35624 13688 35630
rect 13636 35566 13688 35572
rect 12992 33856 13044 33862
rect 12992 33798 13044 33804
rect 13280 33522 13308 35566
rect 13648 35154 13676 35566
rect 13636 35148 13688 35154
rect 13636 35090 13688 35096
rect 13648 33998 13676 35090
rect 13820 34536 13872 34542
rect 13820 34478 13872 34484
rect 13636 33992 13688 33998
rect 13636 33934 13688 33940
rect 13268 33516 13320 33522
rect 13268 33458 13320 33464
rect 12900 33448 12952 33454
rect 12900 33390 12952 33396
rect 12440 33040 12492 33046
rect 12440 32982 12492 32988
rect 12624 33040 12676 33046
rect 12624 32982 12676 32988
rect 12256 32972 12308 32978
rect 12256 32914 12308 32920
rect 12268 31890 12296 32914
rect 12452 32502 12480 32982
rect 12440 32496 12492 32502
rect 12440 32438 12492 32444
rect 12636 32434 12664 32982
rect 12716 32496 12768 32502
rect 12716 32438 12768 32444
rect 12624 32428 12676 32434
rect 12624 32370 12676 32376
rect 12532 32360 12584 32366
rect 12532 32302 12584 32308
rect 12256 31884 12308 31890
rect 12256 31826 12308 31832
rect 12268 31414 12296 31826
rect 12440 31816 12492 31822
rect 12440 31758 12492 31764
rect 12256 31408 12308 31414
rect 12256 31350 12308 31356
rect 12452 31346 12480 31758
rect 12440 31340 12492 31346
rect 12440 31282 12492 31288
rect 12544 30938 12572 32302
rect 12728 31958 12756 32438
rect 12912 32366 12940 33390
rect 12900 32360 12952 32366
rect 12900 32302 12952 32308
rect 12716 31952 12768 31958
rect 12716 31894 12768 31900
rect 13084 31476 13136 31482
rect 13084 31418 13136 31424
rect 12716 31204 12768 31210
rect 12716 31146 12768 31152
rect 12532 30932 12584 30938
rect 12532 30874 12584 30880
rect 12728 30258 12756 31146
rect 12808 30728 12860 30734
rect 12808 30670 12860 30676
rect 12716 30252 12768 30258
rect 12716 30194 12768 30200
rect 12624 29776 12676 29782
rect 12622 29744 12624 29753
rect 12676 29744 12678 29753
rect 12440 29708 12492 29714
rect 12622 29679 12678 29688
rect 12440 29650 12492 29656
rect 12452 29170 12480 29650
rect 12440 29164 12492 29170
rect 12440 29106 12492 29112
rect 12452 28694 12480 29106
rect 12440 28688 12492 28694
rect 12440 28630 12492 28636
rect 12452 27538 12480 28630
rect 12636 28218 12664 29679
rect 12624 28212 12676 28218
rect 12624 28154 12676 28160
rect 12820 28014 12848 30670
rect 13096 30190 13124 31418
rect 13084 30184 13136 30190
rect 13084 30126 13136 30132
rect 12898 29608 12954 29617
rect 12898 29543 12900 29552
rect 12952 29543 12954 29552
rect 12900 29514 12952 29520
rect 13096 28558 13124 30126
rect 13544 29640 13596 29646
rect 13544 29582 13596 29588
rect 13556 29102 13584 29582
rect 13648 29578 13676 33934
rect 13832 33658 13860 34478
rect 13912 34128 13964 34134
rect 13912 34070 13964 34076
rect 13820 33652 13872 33658
rect 13820 33594 13872 33600
rect 13832 33386 13860 33594
rect 13924 33454 13952 34070
rect 13912 33448 13964 33454
rect 13912 33390 13964 33396
rect 13820 33380 13872 33386
rect 13820 33322 13872 33328
rect 13924 33114 13952 33390
rect 13912 33108 13964 33114
rect 13912 33050 13964 33056
rect 13820 32904 13872 32910
rect 13820 32846 13872 32852
rect 13832 32434 13860 32846
rect 13820 32428 13872 32434
rect 13820 32370 13872 32376
rect 13820 31340 13872 31346
rect 13820 31282 13872 31288
rect 13728 30796 13780 30802
rect 13832 30784 13860 31282
rect 14004 31204 14056 31210
rect 14004 31146 14056 31152
rect 14016 30802 14044 31146
rect 13780 30756 13860 30784
rect 14004 30796 14056 30802
rect 13728 30738 13780 30744
rect 14004 30738 14056 30744
rect 13728 29708 13780 29714
rect 13728 29650 13780 29656
rect 13636 29572 13688 29578
rect 13636 29514 13688 29520
rect 13740 29102 13768 29650
rect 13360 29096 13412 29102
rect 13360 29038 13412 29044
rect 13544 29096 13596 29102
rect 13544 29038 13596 29044
rect 13728 29096 13780 29102
rect 13728 29038 13780 29044
rect 13084 28552 13136 28558
rect 13084 28494 13136 28500
rect 12808 28008 12860 28014
rect 12808 27950 12860 27956
rect 12440 27532 12492 27538
rect 12440 27474 12492 27480
rect 12440 26784 12492 26790
rect 12440 26726 12492 26732
rect 12452 26518 12480 26726
rect 12440 26512 12492 26518
rect 12440 26454 12492 26460
rect 12624 26512 12676 26518
rect 12624 26454 12676 26460
rect 12348 26444 12400 26450
rect 12268 26404 12348 26432
rect 12268 25702 12296 26404
rect 12348 26386 12400 26392
rect 12452 25838 12480 26454
rect 12636 26314 12664 26454
rect 12820 26382 12848 27950
rect 12808 26376 12860 26382
rect 12808 26318 12860 26324
rect 12624 26308 12676 26314
rect 12624 26250 12676 26256
rect 12440 25832 12492 25838
rect 12440 25774 12492 25780
rect 12256 25696 12308 25702
rect 12256 25638 12308 25644
rect 12452 25362 12480 25774
rect 12440 25356 12492 25362
rect 12440 25298 12492 25304
rect 12808 25356 12860 25362
rect 12808 25298 12860 25304
rect 12820 24682 12848 25298
rect 12808 24676 12860 24682
rect 12808 24618 12860 24624
rect 12256 24268 12308 24274
rect 12256 24210 12308 24216
rect 12268 23594 12296 24210
rect 12624 23656 12676 23662
rect 12624 23598 12676 23604
rect 12256 23588 12308 23594
rect 12256 23530 12308 23536
rect 12348 23180 12400 23186
rect 12348 23122 12400 23128
rect 12360 22438 12388 23122
rect 12440 23112 12492 23118
rect 12440 23054 12492 23060
rect 12348 22432 12400 22438
rect 12348 22374 12400 22380
rect 12452 22098 12480 23054
rect 12636 22778 12664 23598
rect 12992 23520 13044 23526
rect 12992 23462 13044 23468
rect 12624 22772 12676 22778
rect 12624 22714 12676 22720
rect 12636 22166 12664 22714
rect 13004 22574 13032 23462
rect 12992 22568 13044 22574
rect 12992 22510 13044 22516
rect 12624 22160 12676 22166
rect 12624 22102 12676 22108
rect 12440 22092 12492 22098
rect 12440 22034 12492 22040
rect 12532 22092 12584 22098
rect 12532 22034 12584 22040
rect 12164 21956 12216 21962
rect 12164 21898 12216 21904
rect 10692 21422 10744 21428
rect 10416 21004 10468 21010
rect 10416 20946 10468 20952
rect 10428 20874 10456 20946
rect 10416 20868 10468 20874
rect 10416 20810 10468 20816
rect 10428 20534 10456 20810
rect 10416 20528 10468 20534
rect 10416 20470 10468 20476
rect 10704 20466 10732 21422
rect 10796 21406 10916 21434
rect 11704 21412 11756 21418
rect 10692 20460 10744 20466
rect 10692 20402 10744 20408
rect 10692 19916 10744 19922
rect 10692 19858 10744 19864
rect 10704 19514 10732 19858
rect 10692 19508 10744 19514
rect 10692 19450 10744 19456
rect 10600 18760 10652 18766
rect 10600 18702 10652 18708
rect 10324 17536 10376 17542
rect 10324 17478 10376 17484
rect 10612 16998 10640 18702
rect 10796 17814 10824 21406
rect 11704 21354 11756 21360
rect 11152 21004 11204 21010
rect 11152 20946 11204 20952
rect 11612 21004 11664 21010
rect 11612 20946 11664 20952
rect 10876 20392 10928 20398
rect 10876 20334 10928 20340
rect 10888 19854 10916 20334
rect 11164 20330 11192 20946
rect 11624 20330 11652 20946
rect 11716 20398 11744 21354
rect 12176 20874 12204 21898
rect 12544 21554 12572 22034
rect 12532 21548 12584 21554
rect 12532 21490 12584 21496
rect 12440 21480 12492 21486
rect 12440 21422 12492 21428
rect 12716 21480 12768 21486
rect 12716 21422 12768 21428
rect 12164 20868 12216 20874
rect 12164 20810 12216 20816
rect 12452 20466 12480 21422
rect 12728 21010 12756 21422
rect 12716 21004 12768 21010
rect 12716 20946 12768 20952
rect 12728 20602 12756 20946
rect 13004 20806 13032 22510
rect 13096 21350 13124 28494
rect 13372 28422 13400 29038
rect 13452 28756 13504 28762
rect 13452 28698 13504 28704
rect 13360 28416 13412 28422
rect 13360 28358 13412 28364
rect 13176 27940 13228 27946
rect 13176 27882 13228 27888
rect 13188 26382 13216 27882
rect 13268 26444 13320 26450
rect 13268 26386 13320 26392
rect 13176 26376 13228 26382
rect 13176 26318 13228 26324
rect 13280 25362 13308 26386
rect 13372 25838 13400 28358
rect 13464 27130 13492 28698
rect 13740 28422 13768 29038
rect 13728 28416 13780 28422
rect 13728 28358 13780 28364
rect 13740 27402 13768 28358
rect 13820 28144 13872 28150
rect 13820 28086 13872 28092
rect 13728 27396 13780 27402
rect 13728 27338 13780 27344
rect 13740 27130 13768 27338
rect 13452 27124 13504 27130
rect 13452 27066 13504 27072
rect 13728 27124 13780 27130
rect 13728 27066 13780 27072
rect 13832 26926 13860 28086
rect 13544 26920 13596 26926
rect 13544 26862 13596 26868
rect 13820 26920 13872 26926
rect 13820 26862 13872 26868
rect 13360 25832 13412 25838
rect 13360 25774 13412 25780
rect 13268 25356 13320 25362
rect 13268 25298 13320 25304
rect 13280 24614 13308 25298
rect 13452 25288 13504 25294
rect 13452 25230 13504 25236
rect 13268 24608 13320 24614
rect 13268 24550 13320 24556
rect 13464 24274 13492 25230
rect 13556 24750 13584 26862
rect 13636 26852 13688 26858
rect 13636 26794 13688 26800
rect 13648 26314 13676 26794
rect 13820 26784 13872 26790
rect 13740 26744 13820 26772
rect 13740 26450 13768 26744
rect 13820 26726 13872 26732
rect 13728 26444 13780 26450
rect 13728 26386 13780 26392
rect 13820 26444 13872 26450
rect 13820 26386 13872 26392
rect 13636 26308 13688 26314
rect 13636 26250 13688 26256
rect 13832 25838 13860 26386
rect 13636 25832 13688 25838
rect 13636 25774 13688 25780
rect 13820 25832 13872 25838
rect 13820 25774 13872 25780
rect 13648 24818 13676 25774
rect 13832 25294 13860 25774
rect 13912 25764 13964 25770
rect 13912 25706 13964 25712
rect 13820 25288 13872 25294
rect 13820 25230 13872 25236
rect 13636 24812 13688 24818
rect 13636 24754 13688 24760
rect 13544 24744 13596 24750
rect 13544 24686 13596 24692
rect 13924 24274 13952 25706
rect 14004 24744 14056 24750
rect 14004 24686 14056 24692
rect 13452 24268 13504 24274
rect 13452 24210 13504 24216
rect 13912 24268 13964 24274
rect 13912 24210 13964 24216
rect 14016 24070 14044 24686
rect 14004 24064 14056 24070
rect 14004 24006 14056 24012
rect 14016 23730 14044 24006
rect 14004 23724 14056 23730
rect 14004 23666 14056 23672
rect 13728 23656 13780 23662
rect 13728 23598 13780 23604
rect 13740 23186 13768 23598
rect 13728 23180 13780 23186
rect 13728 23122 13780 23128
rect 13176 23112 13228 23118
rect 13176 23054 13228 23060
rect 13188 22098 13216 23054
rect 13740 22438 13768 23122
rect 14016 22642 14044 23666
rect 13820 22636 13872 22642
rect 13820 22578 13872 22584
rect 14004 22636 14056 22642
rect 14004 22578 14056 22584
rect 13728 22432 13780 22438
rect 13728 22374 13780 22380
rect 13176 22092 13228 22098
rect 13176 22034 13228 22040
rect 13728 22024 13780 22030
rect 13728 21966 13780 21972
rect 13740 21554 13768 21966
rect 13832 21554 13860 22578
rect 13728 21548 13780 21554
rect 13728 21490 13780 21496
rect 13820 21548 13872 21554
rect 13820 21490 13872 21496
rect 13176 21480 13228 21486
rect 13176 21422 13228 21428
rect 13084 21344 13136 21350
rect 13084 21286 13136 21292
rect 13188 21078 13216 21422
rect 13728 21412 13780 21418
rect 13728 21354 13780 21360
rect 13176 21072 13228 21078
rect 13176 21014 13228 21020
rect 13084 20936 13136 20942
rect 13084 20878 13136 20884
rect 12992 20800 13044 20806
rect 12992 20742 13044 20748
rect 12716 20596 12768 20602
rect 12716 20538 12768 20544
rect 12440 20460 12492 20466
rect 12440 20402 12492 20408
rect 11704 20392 11756 20398
rect 11704 20334 11756 20340
rect 11152 20324 11204 20330
rect 11152 20266 11204 20272
rect 11612 20324 11664 20330
rect 11612 20266 11664 20272
rect 11796 20256 11848 20262
rect 11796 20198 11848 20204
rect 11428 20052 11480 20058
rect 11428 19994 11480 20000
rect 10876 19848 10928 19854
rect 10876 19790 10928 19796
rect 10784 17808 10836 17814
rect 10784 17750 10836 17756
rect 10600 16992 10652 16998
rect 10600 16934 10652 16940
rect 10692 16992 10744 16998
rect 10692 16934 10744 16940
rect 10704 16794 10732 16934
rect 10692 16788 10744 16794
rect 10692 16730 10744 16736
rect 10888 16726 10916 19790
rect 11244 19304 11296 19310
rect 11244 19246 11296 19252
rect 11256 18426 11284 19246
rect 11244 18420 11296 18426
rect 11244 18362 11296 18368
rect 11440 17746 11468 19994
rect 11808 19922 11836 20198
rect 13096 19990 13124 20878
rect 13188 20806 13216 21014
rect 13740 21010 13768 21354
rect 13728 21004 13780 21010
rect 13728 20946 13780 20952
rect 13176 20800 13228 20806
rect 13176 20742 13228 20748
rect 13188 20466 13216 20742
rect 13176 20460 13228 20466
rect 13176 20402 13228 20408
rect 13452 20460 13504 20466
rect 13452 20402 13504 20408
rect 13268 20392 13320 20398
rect 13268 20334 13320 20340
rect 13084 19984 13136 19990
rect 13084 19926 13136 19932
rect 11796 19916 11848 19922
rect 11796 19858 11848 19864
rect 12440 19848 12492 19854
rect 12440 19790 12492 19796
rect 12452 19446 12480 19790
rect 12440 19440 12492 19446
rect 12440 19382 12492 19388
rect 12992 19304 13044 19310
rect 12992 19246 13044 19252
rect 11704 19168 11756 19174
rect 11704 19110 11756 19116
rect 11716 18222 11744 19110
rect 12440 18760 12492 18766
rect 12440 18702 12492 18708
rect 11980 18692 12032 18698
rect 11980 18634 12032 18640
rect 11888 18624 11940 18630
rect 11888 18566 11940 18572
rect 11900 18290 11928 18566
rect 11888 18284 11940 18290
rect 11888 18226 11940 18232
rect 11704 18216 11756 18222
rect 11704 18158 11756 18164
rect 11428 17740 11480 17746
rect 11428 17682 11480 17688
rect 11336 17604 11388 17610
rect 11336 17546 11388 17552
rect 10876 16720 10928 16726
rect 10876 16662 10928 16668
rect 11348 16658 11376 17546
rect 10416 16652 10468 16658
rect 10416 16594 10468 16600
rect 11336 16652 11388 16658
rect 11336 16594 11388 16600
rect 10428 14482 10456 16594
rect 11348 16250 11376 16594
rect 11336 16244 11388 16250
rect 11336 16186 11388 16192
rect 10876 15564 10928 15570
rect 10876 15506 10928 15512
rect 10692 14952 10744 14958
rect 10692 14894 10744 14900
rect 10704 14550 10732 14894
rect 10692 14544 10744 14550
rect 10692 14486 10744 14492
rect 10416 14476 10468 14482
rect 10416 14418 10468 14424
rect 10428 13870 10456 14418
rect 10416 13864 10468 13870
rect 10416 13806 10468 13812
rect 10428 13530 10456 13806
rect 10416 13524 10468 13530
rect 10416 13466 10468 13472
rect 10784 13388 10836 13394
rect 10784 13330 10836 13336
rect 10692 12776 10744 12782
rect 10692 12718 10744 12724
rect 10704 12306 10732 12718
rect 10416 12300 10468 12306
rect 10416 12242 10468 12248
rect 10692 12300 10744 12306
rect 10692 12242 10744 12248
rect 10428 9042 10456 12242
rect 10796 11762 10824 13330
rect 10888 12782 10916 15506
rect 11348 14958 11376 16186
rect 11440 15910 11468 17682
rect 11716 17678 11744 18158
rect 11992 17746 12020 18634
rect 11796 17740 11848 17746
rect 11796 17682 11848 17688
rect 11980 17740 12032 17746
rect 11980 17682 12032 17688
rect 11704 17672 11756 17678
rect 11704 17614 11756 17620
rect 11808 17134 11836 17682
rect 11520 17128 11572 17134
rect 11520 17070 11572 17076
rect 11796 17128 11848 17134
rect 11796 17070 11848 17076
rect 11532 16046 11560 17070
rect 11808 16794 11836 17070
rect 11796 16788 11848 16794
rect 11796 16730 11848 16736
rect 11520 16040 11572 16046
rect 11520 15982 11572 15988
rect 11428 15904 11480 15910
rect 11428 15846 11480 15852
rect 11440 15570 11468 15846
rect 11428 15564 11480 15570
rect 11428 15506 11480 15512
rect 11428 15156 11480 15162
rect 11428 15098 11480 15104
rect 11060 14952 11112 14958
rect 11060 14894 11112 14900
rect 11336 14952 11388 14958
rect 11336 14894 11388 14900
rect 11072 13394 11100 14894
rect 11244 14816 11296 14822
rect 11244 14758 11296 14764
rect 11336 14816 11388 14822
rect 11336 14758 11388 14764
rect 11152 14340 11204 14346
rect 11152 14282 11204 14288
rect 11060 13388 11112 13394
rect 11060 13330 11112 13336
rect 11060 12912 11112 12918
rect 11060 12854 11112 12860
rect 10876 12776 10928 12782
rect 10876 12718 10928 12724
rect 10784 11756 10836 11762
rect 10784 11698 10836 11704
rect 11072 11694 11100 12854
rect 11164 12374 11192 14282
rect 11256 14074 11284 14758
rect 11244 14068 11296 14074
rect 11244 14010 11296 14016
rect 11152 12368 11204 12374
rect 11152 12310 11204 12316
rect 11060 11688 11112 11694
rect 11060 11630 11112 11636
rect 11242 11248 11298 11257
rect 11242 11183 11244 11192
rect 11296 11183 11298 11192
rect 11244 11154 11296 11160
rect 10876 11144 10928 11150
rect 10876 11086 10928 11092
rect 10508 11008 10560 11014
rect 10508 10950 10560 10956
rect 10324 9036 10376 9042
rect 10324 8978 10376 8984
rect 10416 9036 10468 9042
rect 10416 8978 10468 8984
rect 10336 7206 10364 8978
rect 10520 8566 10548 10950
rect 10600 10532 10652 10538
rect 10600 10474 10652 10480
rect 10508 8560 10560 8566
rect 10508 8502 10560 8508
rect 10508 7948 10560 7954
rect 10508 7890 10560 7896
rect 10520 7410 10548 7890
rect 10508 7404 10560 7410
rect 10508 7346 10560 7352
rect 10324 7200 10376 7206
rect 10508 7200 10560 7206
rect 10324 7142 10376 7148
rect 10428 7160 10508 7188
rect 10232 6996 10284 7002
rect 10232 6938 10284 6944
rect 10140 6860 10192 6866
rect 10428 6848 10456 7160
rect 10508 7142 10560 7148
rect 10192 6820 10456 6848
rect 10508 6860 10560 6866
rect 10140 6802 10192 6808
rect 10508 6802 10560 6808
rect 10324 6724 10376 6730
rect 10324 6666 10376 6672
rect 10336 5778 10364 6666
rect 9680 5772 9732 5778
rect 9680 5714 9732 5720
rect 9956 5772 10008 5778
rect 9956 5714 10008 5720
rect 10324 5772 10376 5778
rect 10324 5714 10376 5720
rect 9692 5370 9720 5714
rect 10520 5658 10548 6802
rect 10428 5642 10548 5658
rect 10416 5636 10548 5642
rect 10468 5630 10548 5636
rect 10416 5578 10468 5584
rect 9680 5364 9732 5370
rect 9680 5306 9732 5312
rect 10428 5166 10456 5578
rect 10612 5370 10640 10474
rect 10888 10130 10916 11086
rect 11244 10600 11296 10606
rect 11244 10542 11296 10548
rect 10876 10124 10928 10130
rect 10876 10066 10928 10072
rect 11256 9897 11284 10542
rect 11242 9888 11298 9897
rect 11242 9823 11298 9832
rect 11152 9580 11204 9586
rect 11152 9522 11204 9528
rect 11060 9512 11112 9518
rect 11060 9454 11112 9460
rect 10968 9104 11020 9110
rect 10968 9046 11020 9052
rect 10980 8498 11008 9046
rect 11072 8974 11100 9454
rect 11060 8968 11112 8974
rect 11060 8910 11112 8916
rect 11164 8634 11192 9522
rect 11256 9518 11284 9823
rect 11244 9512 11296 9518
rect 11244 9454 11296 9460
rect 11152 8628 11204 8634
rect 11152 8570 11204 8576
rect 11348 8514 11376 14758
rect 11440 14482 11468 15098
rect 11428 14476 11480 14482
rect 11428 14418 11480 14424
rect 11532 14362 11560 15982
rect 11992 15570 12020 17682
rect 12452 17202 12480 18702
rect 12624 18624 12676 18630
rect 12624 18566 12676 18572
rect 12636 17746 12664 18566
rect 12624 17740 12676 17746
rect 12624 17682 12676 17688
rect 12440 17196 12492 17202
rect 12440 17138 12492 17144
rect 12452 16658 12480 17138
rect 12440 16652 12492 16658
rect 12440 16594 12492 16600
rect 11796 15564 11848 15570
rect 11796 15506 11848 15512
rect 11980 15564 12032 15570
rect 11980 15506 12032 15512
rect 11612 15428 11664 15434
rect 11612 15370 11664 15376
rect 11624 14482 11652 15370
rect 11808 14822 11836 15506
rect 11888 15496 11940 15502
rect 11888 15438 11940 15444
rect 11796 14816 11848 14822
rect 11796 14758 11848 14764
rect 11612 14476 11664 14482
rect 11612 14418 11664 14424
rect 11532 14334 11652 14362
rect 11518 12336 11574 12345
rect 11518 12271 11520 12280
rect 11572 12271 11574 12280
rect 11520 12242 11572 12248
rect 11520 12164 11572 12170
rect 11520 12106 11572 12112
rect 11428 11076 11480 11082
rect 11428 11018 11480 11024
rect 11440 9518 11468 11018
rect 11532 10742 11560 12106
rect 11520 10736 11572 10742
rect 11520 10678 11572 10684
rect 11520 10600 11572 10606
rect 11520 10542 11572 10548
rect 11532 10198 11560 10542
rect 11520 10192 11572 10198
rect 11520 10134 11572 10140
rect 11428 9512 11480 9518
rect 11428 9454 11480 9460
rect 10784 8492 10836 8498
rect 10784 8434 10836 8440
rect 10968 8492 11020 8498
rect 10968 8434 11020 8440
rect 11256 8486 11376 8514
rect 10692 7948 10744 7954
rect 10692 7890 10744 7896
rect 10704 7342 10732 7890
rect 10692 7336 10744 7342
rect 10692 7278 10744 7284
rect 10796 5658 10824 8434
rect 10874 7440 10930 7449
rect 10874 7375 10930 7384
rect 10888 7342 10916 7375
rect 10876 7336 10928 7342
rect 10876 7278 10928 7284
rect 10968 5772 11020 5778
rect 10968 5714 11020 5720
rect 10704 5630 10824 5658
rect 10600 5364 10652 5370
rect 10600 5306 10652 5312
rect 10704 5250 10732 5630
rect 10784 5568 10836 5574
rect 10784 5510 10836 5516
rect 10796 5370 10824 5510
rect 10784 5364 10836 5370
rect 10784 5306 10836 5312
rect 10612 5222 10732 5250
rect 10612 5166 10640 5222
rect 10796 5166 10824 5306
rect 10980 5166 11008 5714
rect 10416 5160 10468 5166
rect 10416 5102 10468 5108
rect 10600 5160 10652 5166
rect 10600 5102 10652 5108
rect 10784 5160 10836 5166
rect 10784 5102 10836 5108
rect 10968 5160 11020 5166
rect 10968 5102 11020 5108
rect 10428 4826 10456 5102
rect 10416 4820 10468 4826
rect 10416 4762 10468 4768
rect 10980 4758 11008 5102
rect 11060 5092 11112 5098
rect 11060 5034 11112 5040
rect 10968 4752 11020 4758
rect 10968 4694 11020 4700
rect 11072 4690 11100 5034
rect 10416 4684 10468 4690
rect 10416 4626 10468 4632
rect 11060 4684 11112 4690
rect 11060 4626 11112 4632
rect 9588 4616 9640 4622
rect 9588 4558 9640 4564
rect 9600 3346 9628 4558
rect 10428 4282 10456 4626
rect 10416 4276 10468 4282
rect 10416 4218 10468 4224
rect 9680 4140 9732 4146
rect 9680 4082 9732 4088
rect 9692 3738 9720 4082
rect 10968 4072 11020 4078
rect 10968 4014 11020 4020
rect 10140 4004 10192 4010
rect 10140 3946 10192 3952
rect 9680 3732 9732 3738
rect 9680 3674 9732 3680
rect 9692 3534 9720 3674
rect 9680 3528 9732 3534
rect 9680 3470 9732 3476
rect 9772 3460 9824 3466
rect 9772 3402 9824 3408
rect 9784 3346 9812 3402
rect 9600 3318 9812 3346
rect 9404 3120 9456 3126
rect 9456 3068 9720 3074
rect 9404 3062 9720 3068
rect 9416 3046 9720 3062
rect 9416 2990 9444 3046
rect 8668 2984 8720 2990
rect 8668 2926 8720 2932
rect 8852 2984 8904 2990
rect 8852 2926 8904 2932
rect 9404 2984 9456 2990
rect 9404 2926 9456 2932
rect 9586 2952 9642 2961
rect 9220 2916 9272 2922
rect 9586 2887 9588 2896
rect 9220 2858 9272 2864
rect 9640 2887 9642 2896
rect 9588 2858 9640 2864
rect 9232 2514 9260 2858
rect 9220 2508 9272 2514
rect 9220 2450 9272 2456
rect 9692 2446 9720 3046
rect 9680 2440 9732 2446
rect 9680 2382 9732 2388
rect 10152 800 10180 3946
rect 10980 3602 11008 4014
rect 10968 3596 11020 3602
rect 10968 3538 11020 3544
rect 11072 3126 11100 4626
rect 11256 4078 11284 8486
rect 11336 8424 11388 8430
rect 11336 8366 11388 8372
rect 11348 8090 11376 8366
rect 11336 8084 11388 8090
rect 11336 8026 11388 8032
rect 11624 7342 11652 14334
rect 11796 12776 11848 12782
rect 11796 12718 11848 12724
rect 11704 10600 11756 10606
rect 11704 10542 11756 10548
rect 11716 9110 11744 10542
rect 11808 10062 11836 12718
rect 11900 12306 11928 15438
rect 12452 15162 12480 16594
rect 12636 15638 12664 17682
rect 12716 17672 12768 17678
rect 12716 17614 12768 17620
rect 12728 17202 12756 17614
rect 12716 17196 12768 17202
rect 12716 17138 12768 17144
rect 12808 16040 12860 16046
rect 12808 15982 12860 15988
rect 12820 15638 12848 15982
rect 12624 15632 12676 15638
rect 12624 15574 12676 15580
rect 12808 15632 12860 15638
rect 12808 15574 12860 15580
rect 12440 15156 12492 15162
rect 12440 15098 12492 15104
rect 12164 15088 12216 15094
rect 12164 15030 12216 15036
rect 12072 14952 12124 14958
rect 12072 14894 12124 14900
rect 12084 14074 12112 14894
rect 12176 14074 12204 15030
rect 12440 14952 12492 14958
rect 12440 14894 12492 14900
rect 12452 14414 12480 14894
rect 12440 14408 12492 14414
rect 12440 14350 12492 14356
rect 12072 14068 12124 14074
rect 12072 14010 12124 14016
rect 12164 14068 12216 14074
rect 12164 14010 12216 14016
rect 12440 13864 12492 13870
rect 12492 13812 12756 13818
rect 12440 13806 12756 13812
rect 12452 13790 12756 13806
rect 11980 13388 12032 13394
rect 11980 13330 12032 13336
rect 11992 12442 12020 13330
rect 12440 12640 12492 12646
rect 12440 12582 12492 12588
rect 11980 12436 12032 12442
rect 11980 12378 12032 12384
rect 11888 12300 11940 12306
rect 11888 12242 11940 12248
rect 11888 11552 11940 11558
rect 11888 11494 11940 11500
rect 11900 10606 11928 11494
rect 11992 11082 12020 12378
rect 12348 12232 12400 12238
rect 12348 12174 12400 12180
rect 12360 11898 12388 12174
rect 12348 11892 12400 11898
rect 12348 11834 12400 11840
rect 12452 11694 12480 12582
rect 12532 12232 12584 12238
rect 12532 12174 12584 12180
rect 12440 11688 12492 11694
rect 12440 11630 12492 11636
rect 12072 11280 12124 11286
rect 12072 11222 12124 11228
rect 11980 11076 12032 11082
rect 11980 11018 12032 11024
rect 11888 10600 11940 10606
rect 11888 10542 11940 10548
rect 11796 10056 11848 10062
rect 11796 9998 11848 10004
rect 11808 9586 11836 9998
rect 11796 9580 11848 9586
rect 11796 9522 11848 9528
rect 11704 9104 11756 9110
rect 11704 9046 11756 9052
rect 12084 8974 12112 11222
rect 12544 11218 12572 12174
rect 12728 11354 12756 13790
rect 12716 11348 12768 11354
rect 12716 11290 12768 11296
rect 12348 11212 12400 11218
rect 12348 11154 12400 11160
rect 12532 11212 12584 11218
rect 12532 11154 12584 11160
rect 12254 9616 12310 9625
rect 12254 9551 12310 9560
rect 12164 9036 12216 9042
rect 12164 8978 12216 8984
rect 12072 8968 12124 8974
rect 12072 8910 12124 8916
rect 12084 8430 12112 8910
rect 12176 8498 12204 8978
rect 12164 8492 12216 8498
rect 12164 8434 12216 8440
rect 12072 8424 12124 8430
rect 12072 8366 12124 8372
rect 12268 8362 12296 9551
rect 11796 8356 11848 8362
rect 11796 8298 11848 8304
rect 12256 8356 12308 8362
rect 12256 8298 12308 8304
rect 11808 7954 11836 8298
rect 11796 7948 11848 7954
rect 11796 7890 11848 7896
rect 11612 7336 11664 7342
rect 11612 7278 11664 7284
rect 11624 6390 11652 7278
rect 12072 6860 12124 6866
rect 12072 6802 12124 6808
rect 12084 6730 12112 6802
rect 12072 6724 12124 6730
rect 12072 6666 12124 6672
rect 11980 6656 12032 6662
rect 11980 6598 12032 6604
rect 11612 6384 11664 6390
rect 11612 6326 11664 6332
rect 11428 6248 11480 6254
rect 11428 6190 11480 6196
rect 11440 5302 11468 6190
rect 11992 5778 12020 6598
rect 11980 5772 12032 5778
rect 11980 5714 12032 5720
rect 11888 5704 11940 5710
rect 11888 5646 11940 5652
rect 11428 5296 11480 5302
rect 11428 5238 11480 5244
rect 11900 4622 11928 5646
rect 12084 5166 12112 6666
rect 12072 5160 12124 5166
rect 12072 5102 12124 5108
rect 11888 4616 11940 4622
rect 11888 4558 11940 4564
rect 12360 4486 12388 11154
rect 12820 10282 12848 15574
rect 12900 15156 12952 15162
rect 12900 15098 12952 15104
rect 12912 13802 12940 15098
rect 12900 13796 12952 13802
rect 12900 13738 12952 13744
rect 12912 11626 12940 13738
rect 12900 11620 12952 11626
rect 12900 11562 12952 11568
rect 12728 10254 12848 10282
rect 12624 10056 12676 10062
rect 12624 9998 12676 10004
rect 12440 9988 12492 9994
rect 12440 9930 12492 9936
rect 12452 7818 12480 9930
rect 12532 9648 12584 9654
rect 12530 9616 12532 9625
rect 12584 9616 12586 9625
rect 12530 9551 12586 9560
rect 12532 9512 12584 9518
rect 12530 9480 12532 9489
rect 12584 9480 12586 9489
rect 12530 9415 12586 9424
rect 12636 9042 12664 9998
rect 12532 9036 12584 9042
rect 12532 8978 12584 8984
rect 12624 9036 12676 9042
rect 12624 8978 12676 8984
rect 12544 8022 12572 8978
rect 12532 8016 12584 8022
rect 12532 7958 12584 7964
rect 12532 7880 12584 7886
rect 12532 7822 12584 7828
rect 12440 7812 12492 7818
rect 12440 7754 12492 7760
rect 12544 7546 12572 7822
rect 12624 7812 12676 7818
rect 12624 7754 12676 7760
rect 12532 7540 12584 7546
rect 12532 7482 12584 7488
rect 12440 7336 12492 7342
rect 12440 7278 12492 7284
rect 12452 7206 12480 7278
rect 12636 7206 12664 7754
rect 12440 7200 12492 7206
rect 12440 7142 12492 7148
rect 12624 7200 12676 7206
rect 12624 7142 12676 7148
rect 12452 5166 12480 7142
rect 12532 6112 12584 6118
rect 12532 6054 12584 6060
rect 12544 5234 12572 6054
rect 12636 5710 12664 7142
rect 12624 5704 12676 5710
rect 12624 5646 12676 5652
rect 12532 5228 12584 5234
rect 12532 5170 12584 5176
rect 12440 5160 12492 5166
rect 12440 5102 12492 5108
rect 12348 4480 12400 4486
rect 12348 4422 12400 4428
rect 11244 4072 11296 4078
rect 11244 4014 11296 4020
rect 11060 3120 11112 3126
rect 11060 3062 11112 3068
rect 12360 2990 12388 4422
rect 12544 3602 12572 5170
rect 12624 5160 12676 5166
rect 12728 5148 12756 10254
rect 12808 10124 12860 10130
rect 12808 10066 12860 10072
rect 12820 5710 12848 10066
rect 12912 9489 12940 11562
rect 12898 9480 12954 9489
rect 12898 9415 12954 9424
rect 13004 7410 13032 19246
rect 13176 17740 13228 17746
rect 13176 17682 13228 17688
rect 13188 15910 13216 17682
rect 13280 17610 13308 20334
rect 13268 17604 13320 17610
rect 13268 17546 13320 17552
rect 13464 16046 13492 20402
rect 13740 20398 13768 20946
rect 13728 20392 13780 20398
rect 13728 20334 13780 20340
rect 13820 20392 13872 20398
rect 13820 20334 13872 20340
rect 13832 19310 13860 20334
rect 14108 19718 14136 38218
rect 14200 37262 14228 38354
rect 14188 37256 14240 37262
rect 14188 37198 14240 37204
rect 14752 36310 14780 38354
rect 15568 38208 15620 38214
rect 15568 38150 15620 38156
rect 15016 37800 15068 37806
rect 15016 37742 15068 37748
rect 14924 37664 14976 37670
rect 14924 37606 14976 37612
rect 14936 36582 14964 37606
rect 15028 36718 15056 37742
rect 15108 37188 15160 37194
rect 15108 37130 15160 37136
rect 15016 36712 15068 36718
rect 15016 36654 15068 36660
rect 14924 36576 14976 36582
rect 14924 36518 14976 36524
rect 15016 36576 15068 36582
rect 15120 36530 15148 37130
rect 15580 36786 15608 38150
rect 16224 38010 16252 40200
rect 17316 38548 17368 38554
rect 17316 38490 17368 38496
rect 16580 38480 16632 38486
rect 16580 38422 16632 38428
rect 16212 38004 16264 38010
rect 16212 37946 16264 37952
rect 16212 37868 16264 37874
rect 16212 37810 16264 37816
rect 15752 37800 15804 37806
rect 15752 37742 15804 37748
rect 15568 36780 15620 36786
rect 15568 36722 15620 36728
rect 15068 36524 15148 36530
rect 15016 36518 15148 36524
rect 14936 36310 14964 36518
rect 15028 36502 15148 36518
rect 14740 36304 14792 36310
rect 14740 36246 14792 36252
rect 14924 36304 14976 36310
rect 14924 36246 14976 36252
rect 15028 36174 15056 36502
rect 15108 36236 15160 36242
rect 15108 36178 15160 36184
rect 15016 36168 15068 36174
rect 15016 36110 15068 36116
rect 14924 36032 14976 36038
rect 14924 35974 14976 35980
rect 14936 35630 14964 35974
rect 15120 35698 15148 36178
rect 15108 35692 15160 35698
rect 15108 35634 15160 35640
rect 14924 35624 14976 35630
rect 14924 35566 14976 35572
rect 14936 34610 14964 35566
rect 14924 34604 14976 34610
rect 14924 34546 14976 34552
rect 14372 34536 14424 34542
rect 14372 34478 14424 34484
rect 14280 32904 14332 32910
rect 14280 32846 14332 32852
rect 14292 32434 14320 32846
rect 14280 32428 14332 32434
rect 14280 32370 14332 32376
rect 14384 32366 14412 34478
rect 15120 34066 15148 35634
rect 15568 35624 15620 35630
rect 15568 35566 15620 35572
rect 15580 34610 15608 35566
rect 15292 34604 15344 34610
rect 15292 34546 15344 34552
rect 15568 34604 15620 34610
rect 15568 34546 15620 34552
rect 15108 34060 15160 34066
rect 15108 34002 15160 34008
rect 14832 32428 14884 32434
rect 14832 32370 14884 32376
rect 14372 32360 14424 32366
rect 14372 32302 14424 32308
rect 14556 32360 14608 32366
rect 14556 32302 14608 32308
rect 14188 31272 14240 31278
rect 14188 31214 14240 31220
rect 14200 30054 14228 31214
rect 14384 31142 14412 32302
rect 14464 32292 14516 32298
rect 14464 32234 14516 32240
rect 14476 31822 14504 32234
rect 14464 31816 14516 31822
rect 14464 31758 14516 31764
rect 14372 31136 14424 31142
rect 14372 31078 14424 31084
rect 14384 30258 14412 31078
rect 14372 30252 14424 30258
rect 14372 30194 14424 30200
rect 14476 30190 14504 31758
rect 14568 31482 14596 32302
rect 14844 31686 14872 32370
rect 14832 31680 14884 31686
rect 14832 31622 14884 31628
rect 14556 31476 14608 31482
rect 14556 31418 14608 31424
rect 14844 30870 14872 31622
rect 14832 30864 14884 30870
rect 14832 30806 14884 30812
rect 14464 30184 14516 30190
rect 14464 30126 14516 30132
rect 14844 30122 14872 30806
rect 15120 30666 15148 34002
rect 15200 33992 15252 33998
rect 15200 33934 15252 33940
rect 15212 33454 15240 33934
rect 15304 33522 15332 34546
rect 15292 33516 15344 33522
rect 15292 33458 15344 33464
rect 15200 33448 15252 33454
rect 15200 33390 15252 33396
rect 15660 33448 15712 33454
rect 15660 33390 15712 33396
rect 15476 32972 15528 32978
rect 15476 32914 15528 32920
rect 15568 32972 15620 32978
rect 15568 32914 15620 32920
rect 15292 32904 15344 32910
rect 15292 32846 15344 32852
rect 15200 31816 15252 31822
rect 15200 31758 15252 31764
rect 15212 31346 15240 31758
rect 15200 31340 15252 31346
rect 15200 31282 15252 31288
rect 15304 30870 15332 32846
rect 15488 32570 15516 32914
rect 15476 32564 15528 32570
rect 15476 32506 15528 32512
rect 15384 32428 15436 32434
rect 15384 32370 15436 32376
rect 15396 31482 15424 32370
rect 15488 31890 15516 32506
rect 15476 31884 15528 31890
rect 15476 31826 15528 31832
rect 15384 31476 15436 31482
rect 15384 31418 15436 31424
rect 15396 31278 15424 31418
rect 15384 31272 15436 31278
rect 15384 31214 15436 31220
rect 15292 30864 15344 30870
rect 15292 30806 15344 30812
rect 15384 30728 15436 30734
rect 15384 30670 15436 30676
rect 15108 30660 15160 30666
rect 15108 30602 15160 30608
rect 15292 30592 15344 30598
rect 15292 30534 15344 30540
rect 14832 30116 14884 30122
rect 14832 30058 14884 30064
rect 14188 30048 14240 30054
rect 14188 29990 14240 29996
rect 15200 30048 15252 30054
rect 15200 29990 15252 29996
rect 14280 29708 14332 29714
rect 14280 29650 14332 29656
rect 14292 29306 14320 29650
rect 15212 29510 15240 29990
rect 15304 29714 15332 30534
rect 15396 29714 15424 30670
rect 15580 30054 15608 32914
rect 15672 32434 15700 33390
rect 15660 32428 15712 32434
rect 15660 32370 15712 32376
rect 15660 31952 15712 31958
rect 15660 31894 15712 31900
rect 15568 30048 15620 30054
rect 15568 29990 15620 29996
rect 15292 29708 15344 29714
rect 15292 29650 15344 29656
rect 15384 29708 15436 29714
rect 15384 29650 15436 29656
rect 15672 29646 15700 31894
rect 15660 29640 15712 29646
rect 15660 29582 15712 29588
rect 15200 29504 15252 29510
rect 15200 29446 15252 29452
rect 14280 29300 14332 29306
rect 14280 29242 14332 29248
rect 14292 29102 14320 29242
rect 14280 29096 14332 29102
rect 14280 29038 14332 29044
rect 14648 29096 14700 29102
rect 14648 29038 14700 29044
rect 15660 29096 15712 29102
rect 15660 29038 15712 29044
rect 14556 29028 14608 29034
rect 14556 28970 14608 28976
rect 14464 28008 14516 28014
rect 14464 27950 14516 27956
rect 14280 27600 14332 27606
rect 14280 27542 14332 27548
rect 14292 26042 14320 27542
rect 14476 27538 14504 27950
rect 14568 27538 14596 28970
rect 14660 28422 14688 29038
rect 15672 28626 15700 29038
rect 15660 28620 15712 28626
rect 15660 28562 15712 28568
rect 15200 28552 15252 28558
rect 15200 28494 15252 28500
rect 14648 28416 14700 28422
rect 14648 28358 14700 28364
rect 15212 28218 15240 28494
rect 15200 28212 15252 28218
rect 15200 28154 15252 28160
rect 14924 28144 14976 28150
rect 14924 28086 14976 28092
rect 14464 27532 14516 27538
rect 14464 27474 14516 27480
rect 14556 27532 14608 27538
rect 14556 27474 14608 27480
rect 14936 26246 14964 28086
rect 15384 27940 15436 27946
rect 15384 27882 15436 27888
rect 15396 27606 15424 27882
rect 15384 27600 15436 27606
rect 15384 27542 15436 27548
rect 15476 26852 15528 26858
rect 15476 26794 15528 26800
rect 15108 26444 15160 26450
rect 15108 26386 15160 26392
rect 14924 26240 14976 26246
rect 14924 26182 14976 26188
rect 14280 26036 14332 26042
rect 14280 25978 14332 25984
rect 14292 25922 14320 25978
rect 14200 25894 14320 25922
rect 14200 25362 14228 25894
rect 14280 25832 14332 25838
rect 14280 25774 14332 25780
rect 14292 25430 14320 25774
rect 14280 25424 14332 25430
rect 14280 25366 14332 25372
rect 14188 25356 14240 25362
rect 14188 25298 14240 25304
rect 14556 23656 14608 23662
rect 14556 23598 14608 23604
rect 14188 23180 14240 23186
rect 14188 23122 14240 23128
rect 14200 22982 14228 23122
rect 14188 22976 14240 22982
rect 14188 22918 14240 22924
rect 14200 22642 14228 22918
rect 14188 22636 14240 22642
rect 14188 22578 14240 22584
rect 14188 22228 14240 22234
rect 14188 22170 14240 22176
rect 14200 22098 14228 22170
rect 14568 22098 14596 23598
rect 14188 22092 14240 22098
rect 14188 22034 14240 22040
rect 14556 22092 14608 22098
rect 14556 22034 14608 22040
rect 14200 21078 14228 22034
rect 14464 21480 14516 21486
rect 14464 21422 14516 21428
rect 14188 21072 14240 21078
rect 14188 21014 14240 21020
rect 14280 21072 14332 21078
rect 14280 21014 14332 21020
rect 14188 19916 14240 19922
rect 14188 19858 14240 19864
rect 14096 19712 14148 19718
rect 14096 19654 14148 19660
rect 14200 19514 14228 19858
rect 14188 19508 14240 19514
rect 14188 19450 14240 19456
rect 13820 19304 13872 19310
rect 13820 19246 13872 19252
rect 13544 19236 13596 19242
rect 13544 19178 13596 19184
rect 13556 18766 13584 19178
rect 13544 18760 13596 18766
rect 13544 18702 13596 18708
rect 13728 18624 13780 18630
rect 13728 18566 13780 18572
rect 13452 16040 13504 16046
rect 13452 15982 13504 15988
rect 13176 15904 13228 15910
rect 13176 15846 13228 15852
rect 13188 15026 13216 15846
rect 13636 15360 13688 15366
rect 13636 15302 13688 15308
rect 13176 15020 13228 15026
rect 13176 14962 13228 14968
rect 13544 14816 13596 14822
rect 13544 14758 13596 14764
rect 13556 14618 13584 14758
rect 13544 14612 13596 14618
rect 13544 14554 13596 14560
rect 13544 14476 13596 14482
rect 13648 14464 13676 15302
rect 13740 14482 13768 18566
rect 13832 18222 13860 19246
rect 13820 18216 13872 18222
rect 13820 18158 13872 18164
rect 13832 17202 13860 18158
rect 13820 17196 13872 17202
rect 13820 17138 13872 17144
rect 13820 16992 13872 16998
rect 13820 16934 13872 16940
rect 13832 16726 13860 16934
rect 13820 16720 13872 16726
rect 13820 16662 13872 16668
rect 13832 15094 13860 16662
rect 14004 16652 14056 16658
rect 14004 16594 14056 16600
rect 13912 16448 13964 16454
rect 13912 16390 13964 16396
rect 13924 15706 13952 16390
rect 14016 16182 14044 16594
rect 14004 16176 14056 16182
rect 14004 16118 14056 16124
rect 14292 16046 14320 21014
rect 14372 18964 14424 18970
rect 14372 18906 14424 18912
rect 14384 18630 14412 18906
rect 14372 18624 14424 18630
rect 14372 18566 14424 18572
rect 14280 16040 14332 16046
rect 14280 15982 14332 15988
rect 13912 15700 13964 15706
rect 13912 15642 13964 15648
rect 13820 15088 13872 15094
rect 13820 15030 13872 15036
rect 13924 14940 13952 15642
rect 14096 15020 14148 15026
rect 14096 14962 14148 14968
rect 13832 14912 13952 14940
rect 14004 14952 14056 14958
rect 13596 14436 13676 14464
rect 13544 14418 13596 14424
rect 13268 13864 13320 13870
rect 13268 13806 13320 13812
rect 13360 13864 13412 13870
rect 13360 13806 13412 13812
rect 13280 13258 13308 13806
rect 13268 13252 13320 13258
rect 13268 13194 13320 13200
rect 13268 12708 13320 12714
rect 13268 12650 13320 12656
rect 13176 10668 13228 10674
rect 13176 10610 13228 10616
rect 13188 10130 13216 10610
rect 13176 10124 13228 10130
rect 13176 10066 13228 10072
rect 13176 9036 13228 9042
rect 13176 8978 13228 8984
rect 13188 8838 13216 8978
rect 13176 8832 13228 8838
rect 13176 8774 13228 8780
rect 12992 7404 13044 7410
rect 12992 7346 13044 7352
rect 13188 7342 13216 8774
rect 12900 7336 12952 7342
rect 12900 7278 12952 7284
rect 13176 7336 13228 7342
rect 13176 7278 13228 7284
rect 12912 6866 12940 7278
rect 13084 7200 13136 7206
rect 13084 7142 13136 7148
rect 12900 6860 12952 6866
rect 12900 6802 12952 6808
rect 12912 5914 12940 6802
rect 13096 6798 13124 7142
rect 13084 6792 13136 6798
rect 13084 6734 13136 6740
rect 13280 6254 13308 12650
rect 13372 12646 13400 13806
rect 13544 13184 13596 13190
rect 13544 13126 13596 13132
rect 13360 12640 13412 12646
rect 13360 12582 13412 12588
rect 13360 11348 13412 11354
rect 13360 11290 13412 11296
rect 13372 9042 13400 11290
rect 13556 11218 13584 13126
rect 13648 12442 13676 14436
rect 13728 14476 13780 14482
rect 13728 14418 13780 14424
rect 13740 13870 13768 14418
rect 13728 13864 13780 13870
rect 13728 13806 13780 13812
rect 13728 13388 13780 13394
rect 13728 13330 13780 13336
rect 13740 12918 13768 13330
rect 13832 13326 13860 14912
rect 14004 14894 14056 14900
rect 13912 14476 13964 14482
rect 13912 14418 13964 14424
rect 13924 13870 13952 14418
rect 13912 13864 13964 13870
rect 13912 13806 13964 13812
rect 13820 13320 13872 13326
rect 13820 13262 13872 13268
rect 13728 12912 13780 12918
rect 13728 12854 13780 12860
rect 13740 12782 13768 12854
rect 13820 12844 13872 12850
rect 13924 12832 13952 13806
rect 14016 13258 14044 14894
rect 14004 13252 14056 13258
rect 14004 13194 14056 13200
rect 13872 12804 13952 12832
rect 13820 12786 13872 12792
rect 13728 12776 13780 12782
rect 13728 12718 13780 12724
rect 13636 12436 13688 12442
rect 13636 12378 13688 12384
rect 13924 12374 13952 12804
rect 14016 12782 14044 13194
rect 14004 12776 14056 12782
rect 14004 12718 14056 12724
rect 14004 12640 14056 12646
rect 14004 12582 14056 12588
rect 13912 12368 13964 12374
rect 13912 12310 13964 12316
rect 13636 12096 13688 12102
rect 13636 12038 13688 12044
rect 13544 11212 13596 11218
rect 13544 11154 13596 11160
rect 13648 11150 13676 12038
rect 13820 11756 13872 11762
rect 13820 11698 13872 11704
rect 13636 11144 13688 11150
rect 13636 11086 13688 11092
rect 13832 9042 13860 11698
rect 13912 11688 13964 11694
rect 13912 11630 13964 11636
rect 13924 11558 13952 11630
rect 13912 11552 13964 11558
rect 13912 11494 13964 11500
rect 14016 10606 14044 12582
rect 14108 11762 14136 14962
rect 14188 12776 14240 12782
rect 14188 12718 14240 12724
rect 14096 11756 14148 11762
rect 14096 11698 14148 11704
rect 14200 11218 14228 12718
rect 14292 12646 14320 15982
rect 14476 15706 14504 21422
rect 15120 20534 15148 26386
rect 15200 26308 15252 26314
rect 15200 26250 15252 26256
rect 15212 23594 15240 26250
rect 15384 24744 15436 24750
rect 15384 24686 15436 24692
rect 15396 24410 15424 24686
rect 15384 24404 15436 24410
rect 15384 24346 15436 24352
rect 15488 23866 15516 26794
rect 15672 25770 15700 28562
rect 15660 25764 15712 25770
rect 15660 25706 15712 25712
rect 15660 25288 15712 25294
rect 15660 25230 15712 25236
rect 15672 24818 15700 25230
rect 15660 24812 15712 24818
rect 15660 24754 15712 24760
rect 15476 23860 15528 23866
rect 15476 23802 15528 23808
rect 15292 23792 15344 23798
rect 15292 23734 15344 23740
rect 15200 23588 15252 23594
rect 15200 23530 15252 23536
rect 15304 23186 15332 23734
rect 15292 23180 15344 23186
rect 15292 23122 15344 23128
rect 15200 23112 15252 23118
rect 15200 23054 15252 23060
rect 15212 22166 15240 23054
rect 15304 22234 15332 23122
rect 15384 22568 15436 22574
rect 15384 22510 15436 22516
rect 15292 22228 15344 22234
rect 15292 22170 15344 22176
rect 15200 22160 15252 22166
rect 15200 22102 15252 22108
rect 15292 21956 15344 21962
rect 15292 21898 15344 21904
rect 15304 21010 15332 21898
rect 15396 21146 15424 22510
rect 15384 21140 15436 21146
rect 15384 21082 15436 21088
rect 15292 21004 15344 21010
rect 15292 20946 15344 20952
rect 15108 20528 15160 20534
rect 15108 20470 15160 20476
rect 15016 20392 15068 20398
rect 15016 20334 15068 20340
rect 14740 19848 14792 19854
rect 15028 19802 15056 20334
rect 14740 19790 14792 19796
rect 14752 19378 14780 19790
rect 14844 19786 15056 19802
rect 14832 19780 15056 19786
rect 14884 19774 15056 19780
rect 14832 19722 14884 19728
rect 14740 19372 14792 19378
rect 14740 19314 14792 19320
rect 14924 19372 14976 19378
rect 14924 19314 14976 19320
rect 14556 19168 14608 19174
rect 14556 19110 14608 19116
rect 14568 18834 14596 19110
rect 14556 18828 14608 18834
rect 14556 18770 14608 18776
rect 14556 16040 14608 16046
rect 14556 15982 14608 15988
rect 14568 15706 14596 15982
rect 14464 15700 14516 15706
rect 14464 15642 14516 15648
rect 14556 15700 14608 15706
rect 14556 15642 14608 15648
rect 14648 15564 14700 15570
rect 14648 15506 14700 15512
rect 14556 14952 14608 14958
rect 14556 14894 14608 14900
rect 14568 14618 14596 14894
rect 14556 14612 14608 14618
rect 14556 14554 14608 14560
rect 14280 12640 14332 12646
rect 14280 12582 14332 12588
rect 14372 12368 14424 12374
rect 14372 12310 14424 12316
rect 14280 12300 14332 12306
rect 14280 12242 14332 12248
rect 14188 11212 14240 11218
rect 14188 11154 14240 11160
rect 14004 10600 14056 10606
rect 14004 10542 14056 10548
rect 14016 10130 14044 10542
rect 14004 10124 14056 10130
rect 14004 10066 14056 10072
rect 14292 9042 14320 12242
rect 14384 11354 14412 12310
rect 14556 12300 14608 12306
rect 14556 12242 14608 12248
rect 14372 11348 14424 11354
rect 14372 11290 14424 11296
rect 14568 10198 14596 12242
rect 14556 10192 14608 10198
rect 14556 10134 14608 10140
rect 14372 9512 14424 9518
rect 14372 9454 14424 9460
rect 13360 9036 13412 9042
rect 13360 8978 13412 8984
rect 13820 9036 13872 9042
rect 13820 8978 13872 8984
rect 14280 9036 14332 9042
rect 14280 8978 14332 8984
rect 14096 8900 14148 8906
rect 14096 8842 14148 8848
rect 13820 8492 13872 8498
rect 13820 8434 13872 8440
rect 13544 8424 13596 8430
rect 13544 8366 13596 8372
rect 13556 6458 13584 8366
rect 13832 7954 13860 8434
rect 13912 8424 13964 8430
rect 13912 8366 13964 8372
rect 13820 7948 13872 7954
rect 13820 7890 13872 7896
rect 13820 7744 13872 7750
rect 13820 7686 13872 7692
rect 13544 6452 13596 6458
rect 13544 6394 13596 6400
rect 13832 6254 13860 7686
rect 13924 7342 13952 8366
rect 14004 7404 14056 7410
rect 14004 7346 14056 7352
rect 13912 7336 13964 7342
rect 13912 7278 13964 7284
rect 13924 6254 13952 7278
rect 14016 6866 14044 7346
rect 14004 6860 14056 6866
rect 14004 6802 14056 6808
rect 14108 6712 14136 8842
rect 14384 8498 14412 9454
rect 14568 9178 14596 10134
rect 14660 9518 14688 15506
rect 14648 9512 14700 9518
rect 14648 9454 14700 9460
rect 14740 9512 14792 9518
rect 14740 9454 14792 9460
rect 14556 9172 14608 9178
rect 14556 9114 14608 9120
rect 14372 8492 14424 8498
rect 14372 8434 14424 8440
rect 14648 8424 14700 8430
rect 14752 8412 14780 9454
rect 14700 8384 14780 8412
rect 14648 8366 14700 8372
rect 14556 8084 14608 8090
rect 14556 8026 14608 8032
rect 14372 7540 14424 7546
rect 14372 7482 14424 7488
rect 14384 7274 14412 7482
rect 14462 7440 14518 7449
rect 14462 7375 14518 7384
rect 14476 7342 14504 7375
rect 14464 7336 14516 7342
rect 14464 7278 14516 7284
rect 14372 7268 14424 7274
rect 14372 7210 14424 7216
rect 14476 6934 14504 7278
rect 14464 6928 14516 6934
rect 14464 6870 14516 6876
rect 14016 6684 14136 6712
rect 13268 6248 13320 6254
rect 13268 6190 13320 6196
rect 13820 6248 13872 6254
rect 13820 6190 13872 6196
rect 13912 6248 13964 6254
rect 13912 6190 13964 6196
rect 12900 5908 12952 5914
rect 12900 5850 12952 5856
rect 12808 5704 12860 5710
rect 12808 5646 12860 5652
rect 13728 5636 13780 5642
rect 13728 5578 13780 5584
rect 12728 5120 12848 5148
rect 12624 5102 12676 5108
rect 12532 3596 12584 3602
rect 12532 3538 12584 3544
rect 12440 3528 12492 3534
rect 12440 3470 12492 3476
rect 12452 2990 12480 3470
rect 12636 3398 12664 5102
rect 12716 5024 12768 5030
rect 12716 4966 12768 4972
rect 12624 3392 12676 3398
rect 12624 3334 12676 3340
rect 12348 2984 12400 2990
rect 12348 2926 12400 2932
rect 12440 2984 12492 2990
rect 12440 2926 12492 2932
rect 12452 2446 12480 2926
rect 12636 2514 12664 3334
rect 12728 3058 12756 4966
rect 12820 4078 12848 5120
rect 13740 4162 13768 5578
rect 13924 5166 13952 6190
rect 13912 5160 13964 5166
rect 13912 5102 13964 5108
rect 13912 4616 13964 4622
rect 13912 4558 13964 4564
rect 13740 4146 13860 4162
rect 13740 4140 13872 4146
rect 13740 4134 13820 4140
rect 13820 4082 13872 4088
rect 12808 4072 12860 4078
rect 12808 4014 12860 4020
rect 13544 4004 13596 4010
rect 13544 3946 13596 3952
rect 13556 3602 13584 3946
rect 13544 3596 13596 3602
rect 13544 3538 13596 3544
rect 13176 3528 13228 3534
rect 13176 3470 13228 3476
rect 12716 3052 12768 3058
rect 12716 2994 12768 3000
rect 12624 2508 12676 2514
rect 12624 2450 12676 2456
rect 13188 2446 13216 3470
rect 13924 2854 13952 4558
rect 13912 2848 13964 2854
rect 13912 2790 13964 2796
rect 13924 2446 13952 2790
rect 12440 2440 12492 2446
rect 12440 2382 12492 2388
rect 13176 2440 13228 2446
rect 13176 2382 13228 2388
rect 13912 2440 13964 2446
rect 13912 2382 13964 2388
rect 11980 2304 12032 2310
rect 11980 2246 12032 2252
rect 11992 800 12020 2246
rect 14016 800 14044 6684
rect 14096 6452 14148 6458
rect 14096 6394 14148 6400
rect 14108 4622 14136 6394
rect 14280 6316 14332 6322
rect 14280 6258 14332 6264
rect 14188 4684 14240 4690
rect 14188 4626 14240 4632
rect 14096 4616 14148 4622
rect 14096 4558 14148 4564
rect 14096 3392 14148 3398
rect 14096 3334 14148 3340
rect 14108 2514 14136 3334
rect 14200 3194 14228 4626
rect 14292 4146 14320 6258
rect 14568 6254 14596 8026
rect 14660 7750 14688 8366
rect 14648 7744 14700 7750
rect 14648 7686 14700 7692
rect 14660 7342 14688 7686
rect 14648 7336 14700 7342
rect 14648 7278 14700 7284
rect 14660 6254 14688 7278
rect 14936 6458 14964 19314
rect 15028 19310 15056 19774
rect 15016 19304 15068 19310
rect 15016 19246 15068 19252
rect 14924 6452 14976 6458
rect 14924 6394 14976 6400
rect 15028 6338 15056 19246
rect 15120 15434 15148 20470
rect 15292 20256 15344 20262
rect 15292 20198 15344 20204
rect 15200 19916 15252 19922
rect 15200 19858 15252 19864
rect 15212 19446 15240 19858
rect 15200 19440 15252 19446
rect 15200 19382 15252 19388
rect 15212 18170 15240 19382
rect 15304 19310 15332 20198
rect 15292 19304 15344 19310
rect 15292 19246 15344 19252
rect 15384 18896 15436 18902
rect 15384 18838 15436 18844
rect 15396 18426 15424 18838
rect 15384 18420 15436 18426
rect 15384 18362 15436 18368
rect 15212 18142 15332 18170
rect 15200 18080 15252 18086
rect 15200 18022 15252 18028
rect 15212 17746 15240 18022
rect 15200 17740 15252 17746
rect 15200 17682 15252 17688
rect 15304 16658 15332 18142
rect 15660 17672 15712 17678
rect 15660 17614 15712 17620
rect 15476 17196 15528 17202
rect 15476 17138 15528 17144
rect 15488 17082 15516 17138
rect 15488 17054 15608 17082
rect 15292 16652 15344 16658
rect 15292 16594 15344 16600
rect 15108 15428 15160 15434
rect 15108 15370 15160 15376
rect 15476 15428 15528 15434
rect 15476 15370 15528 15376
rect 15292 14952 15344 14958
rect 15292 14894 15344 14900
rect 15200 13864 15252 13870
rect 15200 13806 15252 13812
rect 15108 13184 15160 13190
rect 15108 13126 15160 13132
rect 15120 12782 15148 13126
rect 15108 12776 15160 12782
rect 15108 12718 15160 12724
rect 15108 11212 15160 11218
rect 15108 11154 15160 11160
rect 15120 9586 15148 11154
rect 15108 9580 15160 9586
rect 15108 9522 15160 9528
rect 15108 8900 15160 8906
rect 15108 8842 15160 8848
rect 15120 8537 15148 8842
rect 15106 8528 15162 8537
rect 15106 8463 15162 8472
rect 14844 6310 15056 6338
rect 14556 6248 14608 6254
rect 14556 6190 14608 6196
rect 14648 6248 14700 6254
rect 14648 6190 14700 6196
rect 14568 5914 14596 6190
rect 14556 5908 14608 5914
rect 14556 5850 14608 5856
rect 14280 4140 14332 4146
rect 14280 4082 14332 4088
rect 14568 3942 14596 5850
rect 14660 5166 14688 6190
rect 14648 5160 14700 5166
rect 14648 5102 14700 5108
rect 14556 3936 14608 3942
rect 14556 3878 14608 3884
rect 14844 3738 14872 6310
rect 15212 5234 15240 13806
rect 15304 13734 15332 14894
rect 15384 14476 15436 14482
rect 15488 14464 15516 15370
rect 15436 14436 15516 14464
rect 15384 14418 15436 14424
rect 15292 13728 15344 13734
rect 15292 13670 15344 13676
rect 15396 11898 15424 14418
rect 15580 14362 15608 17054
rect 15672 16794 15700 17614
rect 15764 17542 15792 37742
rect 15844 37324 15896 37330
rect 15844 37266 15896 37272
rect 15856 35630 15884 37266
rect 16224 37262 16252 37810
rect 16488 37324 16540 37330
rect 16488 37266 16540 37272
rect 16212 37256 16264 37262
rect 16212 37198 16264 37204
rect 16224 36922 16252 37198
rect 16212 36916 16264 36922
rect 16212 36858 16264 36864
rect 16224 36786 16252 36858
rect 16304 36848 16356 36854
rect 16304 36790 16356 36796
rect 16212 36780 16264 36786
rect 16212 36722 16264 36728
rect 15844 35624 15896 35630
rect 15844 35566 15896 35572
rect 15856 34542 15884 35566
rect 16120 35148 16172 35154
rect 16120 35090 16172 35096
rect 16132 34746 16160 35090
rect 16224 34950 16252 36722
rect 16316 36242 16344 36790
rect 16304 36236 16356 36242
rect 16304 36178 16356 36184
rect 16304 35080 16356 35086
rect 16304 35022 16356 35028
rect 16396 35080 16448 35086
rect 16396 35022 16448 35028
rect 16212 34944 16264 34950
rect 16212 34886 16264 34892
rect 16120 34740 16172 34746
rect 16120 34682 16172 34688
rect 16028 34672 16080 34678
rect 16028 34614 16080 34620
rect 15844 34536 15896 34542
rect 15844 34478 15896 34484
rect 15936 33856 15988 33862
rect 15936 33798 15988 33804
rect 15948 33522 15976 33798
rect 15936 33516 15988 33522
rect 15936 33458 15988 33464
rect 15936 32836 15988 32842
rect 15936 32778 15988 32784
rect 15948 32434 15976 32778
rect 15936 32428 15988 32434
rect 15936 32370 15988 32376
rect 15936 29708 15988 29714
rect 15936 29650 15988 29656
rect 15948 29102 15976 29650
rect 15936 29096 15988 29102
rect 15936 29038 15988 29044
rect 15844 28008 15896 28014
rect 15844 27950 15896 27956
rect 15856 24342 15884 27950
rect 15936 27872 15988 27878
rect 15936 27814 15988 27820
rect 15948 27674 15976 27814
rect 15936 27668 15988 27674
rect 15936 27610 15988 27616
rect 15844 24336 15896 24342
rect 15844 24278 15896 24284
rect 16040 22148 16068 34614
rect 16316 34066 16344 35022
rect 16304 34060 16356 34066
rect 16304 34002 16356 34008
rect 16408 33454 16436 35022
rect 16500 34678 16528 37266
rect 16592 36689 16620 38422
rect 17224 38004 17276 38010
rect 17224 37946 17276 37952
rect 17236 37466 17264 37946
rect 17224 37460 17276 37466
rect 17224 37402 17276 37408
rect 17328 37194 17356 38490
rect 18248 37398 18276 40200
rect 19580 38652 19876 38672
rect 19636 38650 19660 38652
rect 19716 38650 19740 38652
rect 19796 38650 19820 38652
rect 19658 38598 19660 38650
rect 19722 38598 19734 38650
rect 19796 38598 19798 38650
rect 19636 38596 19660 38598
rect 19716 38596 19740 38598
rect 19796 38596 19820 38598
rect 19580 38576 19876 38596
rect 18512 37800 18564 37806
rect 18512 37742 18564 37748
rect 18696 37800 18748 37806
rect 18696 37742 18748 37748
rect 19156 37800 19208 37806
rect 19156 37742 19208 37748
rect 19432 37800 19484 37806
rect 19432 37742 19484 37748
rect 18236 37392 18288 37398
rect 18236 37334 18288 37340
rect 18524 37330 18552 37742
rect 18512 37324 18564 37330
rect 18512 37266 18564 37272
rect 17316 37188 17368 37194
rect 17316 37130 17368 37136
rect 18236 36780 18288 36786
rect 18236 36722 18288 36728
rect 18420 36780 18472 36786
rect 18420 36722 18472 36728
rect 16578 36680 16634 36689
rect 16578 36615 16634 36624
rect 16592 36242 16620 36615
rect 18144 36576 18196 36582
rect 18144 36518 18196 36524
rect 17040 36304 17092 36310
rect 17040 36246 17092 36252
rect 16580 36236 16632 36242
rect 16580 36178 16632 36184
rect 16856 36236 16908 36242
rect 16856 36178 16908 36184
rect 16592 35306 16620 36178
rect 16672 36168 16724 36174
rect 16672 36110 16724 36116
rect 16684 35834 16712 36110
rect 16672 35828 16724 35834
rect 16672 35770 16724 35776
rect 16868 35698 16896 36178
rect 16856 35692 16908 35698
rect 16856 35634 16908 35640
rect 16764 35624 16816 35630
rect 16764 35566 16816 35572
rect 16948 35624 17000 35630
rect 16948 35566 17000 35572
rect 16592 35278 16712 35306
rect 16580 35012 16632 35018
rect 16580 34954 16632 34960
rect 16488 34672 16540 34678
rect 16488 34614 16540 34620
rect 16488 34536 16540 34542
rect 16488 34478 16540 34484
rect 16500 33998 16528 34478
rect 16488 33992 16540 33998
rect 16488 33934 16540 33940
rect 16396 33448 16448 33454
rect 16396 33390 16448 33396
rect 16592 33114 16620 34954
rect 16580 33108 16632 33114
rect 16580 33050 16632 33056
rect 16396 32428 16448 32434
rect 16396 32370 16448 32376
rect 16408 31142 16436 32370
rect 16396 31136 16448 31142
rect 16396 31078 16448 31084
rect 16120 30796 16172 30802
rect 16120 30738 16172 30744
rect 16132 30258 16160 30738
rect 16408 30734 16436 31078
rect 16396 30728 16448 30734
rect 16396 30670 16448 30676
rect 16120 30252 16172 30258
rect 16120 30194 16172 30200
rect 16396 29096 16448 29102
rect 16396 29038 16448 29044
rect 16408 28626 16436 29038
rect 16684 28762 16712 35278
rect 16776 35222 16804 35566
rect 16764 35216 16816 35222
rect 16764 35158 16816 35164
rect 16776 34746 16804 35158
rect 16960 35154 16988 35566
rect 16948 35148 17000 35154
rect 16948 35090 17000 35096
rect 16764 34740 16816 34746
rect 16764 34682 16816 34688
rect 16948 34060 17000 34066
rect 16948 34002 17000 34008
rect 16960 33658 16988 34002
rect 16948 33652 17000 33658
rect 16948 33594 17000 33600
rect 16948 32972 17000 32978
rect 16948 32914 17000 32920
rect 16856 32836 16908 32842
rect 16856 32778 16908 32784
rect 16672 28756 16724 28762
rect 16672 28698 16724 28704
rect 16396 28620 16448 28626
rect 16396 28562 16448 28568
rect 16408 26450 16436 28562
rect 16672 28484 16724 28490
rect 16672 28426 16724 28432
rect 16684 28082 16712 28426
rect 16672 28076 16724 28082
rect 16672 28018 16724 28024
rect 16868 26926 16896 32778
rect 16960 31822 16988 32914
rect 16948 31816 17000 31822
rect 16948 31758 17000 31764
rect 16948 29096 17000 29102
rect 16948 29038 17000 29044
rect 16960 28626 16988 29038
rect 16948 28620 17000 28626
rect 16948 28562 17000 28568
rect 16580 26920 16632 26926
rect 16580 26862 16632 26868
rect 16856 26920 16908 26926
rect 16856 26862 16908 26868
rect 16120 26444 16172 26450
rect 16120 26386 16172 26392
rect 16396 26444 16448 26450
rect 16396 26386 16448 26392
rect 16132 25838 16160 26386
rect 16408 25838 16436 26386
rect 16592 26042 16620 26862
rect 16580 26036 16632 26042
rect 16580 25978 16632 25984
rect 16120 25832 16172 25838
rect 16120 25774 16172 25780
rect 16396 25832 16448 25838
rect 16396 25774 16448 25780
rect 16132 25362 16160 25774
rect 16120 25356 16172 25362
rect 16120 25298 16172 25304
rect 16132 24614 16160 25298
rect 16960 25158 16988 28562
rect 17052 27538 17080 36246
rect 18156 36242 18184 36518
rect 18144 36236 18196 36242
rect 18144 36178 18196 36184
rect 17316 36168 17368 36174
rect 17316 36110 17368 36116
rect 17132 35080 17184 35086
rect 17132 35022 17184 35028
rect 17144 34202 17172 35022
rect 17132 34196 17184 34202
rect 17132 34138 17184 34144
rect 17328 34066 17356 36110
rect 18248 34066 18276 36722
rect 18328 35624 18380 35630
rect 18328 35566 18380 35572
rect 18340 34542 18368 35566
rect 18432 35494 18460 36722
rect 18524 36310 18552 37266
rect 18708 37262 18736 37742
rect 18880 37664 18932 37670
rect 18880 37606 18932 37612
rect 18788 37460 18840 37466
rect 18788 37402 18840 37408
rect 18696 37256 18748 37262
rect 18696 37198 18748 37204
rect 18512 36304 18564 36310
rect 18512 36246 18564 36252
rect 18708 36174 18736 37198
rect 18800 36922 18828 37402
rect 18788 36916 18840 36922
rect 18788 36858 18840 36864
rect 18696 36168 18748 36174
rect 18696 36110 18748 36116
rect 18800 35698 18828 36858
rect 18788 35692 18840 35698
rect 18788 35634 18840 35640
rect 18892 35630 18920 37606
rect 19168 36242 19196 37742
rect 19340 37732 19392 37738
rect 19340 37674 19392 37680
rect 19352 37398 19380 37674
rect 19340 37392 19392 37398
rect 19340 37334 19392 37340
rect 19352 36242 19380 37334
rect 19444 37262 19472 37742
rect 19580 37564 19876 37584
rect 19636 37562 19660 37564
rect 19716 37562 19740 37564
rect 19796 37562 19820 37564
rect 19658 37510 19660 37562
rect 19722 37510 19734 37562
rect 19796 37510 19798 37562
rect 19636 37508 19660 37510
rect 19716 37508 19740 37510
rect 19796 37508 19820 37510
rect 19580 37488 19876 37508
rect 19892 37324 19944 37330
rect 19892 37266 19944 37272
rect 19432 37256 19484 37262
rect 19432 37198 19484 37204
rect 19444 36310 19472 37198
rect 19904 36854 19932 37266
rect 19892 36848 19944 36854
rect 19892 36790 19944 36796
rect 19800 36712 19852 36718
rect 19798 36680 19800 36689
rect 19852 36680 19854 36689
rect 19798 36615 19854 36624
rect 19580 36476 19876 36496
rect 19636 36474 19660 36476
rect 19716 36474 19740 36476
rect 19796 36474 19820 36476
rect 19658 36422 19660 36474
rect 19722 36422 19734 36474
rect 19796 36422 19798 36474
rect 19636 36420 19660 36422
rect 19716 36420 19740 36422
rect 19796 36420 19820 36422
rect 19580 36400 19876 36420
rect 19432 36304 19484 36310
rect 19432 36246 19484 36252
rect 19156 36236 19208 36242
rect 19156 36178 19208 36184
rect 19340 36236 19392 36242
rect 19340 36178 19392 36184
rect 19168 36106 19196 36178
rect 19156 36100 19208 36106
rect 19156 36042 19208 36048
rect 19352 35630 19380 36178
rect 18880 35624 18932 35630
rect 18880 35566 18932 35572
rect 19340 35624 19392 35630
rect 19340 35566 19392 35572
rect 18420 35488 18472 35494
rect 18420 35430 18472 35436
rect 19352 35154 19380 35566
rect 19904 35562 19932 36790
rect 20088 36650 20116 40200
rect 20996 38412 21048 38418
rect 20996 38354 21048 38360
rect 21548 38412 21600 38418
rect 21548 38354 21600 38360
rect 20720 38344 20772 38350
rect 20720 38286 20772 38292
rect 20536 38208 20588 38214
rect 20536 38150 20588 38156
rect 20548 37806 20576 38150
rect 20536 37800 20588 37806
rect 20536 37742 20588 37748
rect 20076 36644 20128 36650
rect 20076 36586 20128 36592
rect 20260 36576 20312 36582
rect 20260 36518 20312 36524
rect 20444 36576 20496 36582
rect 20444 36518 20496 36524
rect 20272 35766 20300 36518
rect 20456 36310 20484 36518
rect 20444 36304 20496 36310
rect 20444 36246 20496 36252
rect 20536 36236 20588 36242
rect 20536 36178 20588 36184
rect 20260 35760 20312 35766
rect 20260 35702 20312 35708
rect 19892 35556 19944 35562
rect 19892 35498 19944 35504
rect 19580 35388 19876 35408
rect 19636 35386 19660 35388
rect 19716 35386 19740 35388
rect 19796 35386 19820 35388
rect 19658 35334 19660 35386
rect 19722 35334 19734 35386
rect 19796 35334 19798 35386
rect 19636 35332 19660 35334
rect 19716 35332 19740 35334
rect 19796 35332 19820 35334
rect 19580 35312 19876 35332
rect 19432 35284 19484 35290
rect 19432 35226 19484 35232
rect 18972 35148 19024 35154
rect 18972 35090 19024 35096
rect 19340 35148 19392 35154
rect 19340 35090 19392 35096
rect 18984 34610 19012 35090
rect 19444 34746 19472 35226
rect 20260 35148 20312 35154
rect 20260 35090 20312 35096
rect 19432 34740 19484 34746
rect 19432 34682 19484 34688
rect 18972 34604 19024 34610
rect 18972 34546 19024 34552
rect 18328 34536 18380 34542
rect 18328 34478 18380 34484
rect 18696 34400 18748 34406
rect 18696 34342 18748 34348
rect 18708 34066 18736 34342
rect 17316 34060 17368 34066
rect 17316 34002 17368 34008
rect 18236 34060 18288 34066
rect 18236 34002 18288 34008
rect 18696 34060 18748 34066
rect 18696 34002 18748 34008
rect 17224 33992 17276 33998
rect 17224 33934 17276 33940
rect 17236 33658 17264 33934
rect 17224 33652 17276 33658
rect 17224 33594 17276 33600
rect 18984 33454 19012 34546
rect 20168 34468 20220 34474
rect 20168 34410 20220 34416
rect 19580 34300 19876 34320
rect 19636 34298 19660 34300
rect 19716 34298 19740 34300
rect 19796 34298 19820 34300
rect 19658 34246 19660 34298
rect 19722 34246 19734 34298
rect 19796 34246 19798 34298
rect 19636 34244 19660 34246
rect 19716 34244 19740 34246
rect 19796 34244 19820 34246
rect 19580 34224 19876 34244
rect 19984 33856 20036 33862
rect 19984 33798 20036 33804
rect 19064 33584 19116 33590
rect 19064 33526 19116 33532
rect 18328 33448 18380 33454
rect 18328 33390 18380 33396
rect 18972 33448 19024 33454
rect 18972 33390 19024 33396
rect 17684 33312 17736 33318
rect 17684 33254 17736 33260
rect 18144 33312 18196 33318
rect 18144 33254 18196 33260
rect 17316 33108 17368 33114
rect 17316 33050 17368 33056
rect 17224 33040 17276 33046
rect 17224 32982 17276 32988
rect 17132 31952 17184 31958
rect 17132 31894 17184 31900
rect 17144 31770 17172 31894
rect 17236 31890 17264 32982
rect 17224 31884 17276 31890
rect 17224 31826 17276 31832
rect 17144 31754 17264 31770
rect 17144 31748 17276 31754
rect 17144 31742 17224 31748
rect 17224 31690 17276 31696
rect 17236 30802 17264 31690
rect 17328 31278 17356 33050
rect 17500 32972 17552 32978
rect 17500 32914 17552 32920
rect 17512 32502 17540 32914
rect 17500 32496 17552 32502
rect 17500 32438 17552 32444
rect 17592 31816 17644 31822
rect 17592 31758 17644 31764
rect 17316 31272 17368 31278
rect 17316 31214 17368 31220
rect 17604 30802 17632 31758
rect 17696 30802 17724 33254
rect 18156 32978 18184 33254
rect 18340 32978 18368 33390
rect 19076 33386 19104 33526
rect 19892 33448 19944 33454
rect 19892 33390 19944 33396
rect 19064 33380 19116 33386
rect 19064 33322 19116 33328
rect 19076 32978 19104 33322
rect 19248 33312 19300 33318
rect 19248 33254 19300 33260
rect 18144 32972 18196 32978
rect 18144 32914 18196 32920
rect 18328 32972 18380 32978
rect 18328 32914 18380 32920
rect 19064 32972 19116 32978
rect 19064 32914 19116 32920
rect 17868 32768 17920 32774
rect 17868 32710 17920 32716
rect 17880 32026 17908 32710
rect 17868 32020 17920 32026
rect 17868 31962 17920 31968
rect 17880 30870 17908 31962
rect 17868 30864 17920 30870
rect 17868 30806 17920 30812
rect 17132 30796 17184 30802
rect 17132 30738 17184 30744
rect 17224 30796 17276 30802
rect 17224 30738 17276 30744
rect 17592 30796 17644 30802
rect 17592 30738 17644 30744
rect 17684 30796 17736 30802
rect 17684 30738 17736 30744
rect 17144 28762 17172 30738
rect 17236 29102 17264 30738
rect 18236 30660 18288 30666
rect 18236 30602 18288 30608
rect 18248 29714 18276 30602
rect 17592 29708 17644 29714
rect 17592 29650 17644 29656
rect 18236 29708 18288 29714
rect 18236 29650 18288 29656
rect 17604 29306 17632 29650
rect 18340 29306 18368 32914
rect 19260 32910 19288 33254
rect 19580 33212 19876 33232
rect 19636 33210 19660 33212
rect 19716 33210 19740 33212
rect 19796 33210 19820 33212
rect 19658 33158 19660 33210
rect 19722 33158 19734 33210
rect 19796 33158 19798 33210
rect 19636 33156 19660 33158
rect 19716 33156 19740 33158
rect 19796 33156 19820 33158
rect 19580 33136 19876 33156
rect 19248 32904 19300 32910
rect 19248 32846 19300 32852
rect 19064 32836 19116 32842
rect 19064 32778 19116 32784
rect 19156 32836 19208 32842
rect 19156 32778 19208 32784
rect 18604 32360 18656 32366
rect 18604 32302 18656 32308
rect 18418 32192 18474 32201
rect 18418 32127 18474 32136
rect 18432 31958 18460 32127
rect 18616 31958 18644 32302
rect 18788 32020 18840 32026
rect 18788 31962 18840 31968
rect 18420 31952 18472 31958
rect 18420 31894 18472 31900
rect 18604 31952 18656 31958
rect 18604 31894 18656 31900
rect 18512 30252 18564 30258
rect 18512 30194 18564 30200
rect 18420 29572 18472 29578
rect 18420 29514 18472 29520
rect 17592 29300 17644 29306
rect 17592 29242 17644 29248
rect 18328 29300 18380 29306
rect 18328 29242 18380 29248
rect 17316 29232 17368 29238
rect 17316 29174 17368 29180
rect 17224 29096 17276 29102
rect 17224 29038 17276 29044
rect 17132 28756 17184 28762
rect 17132 28698 17184 28704
rect 17040 27532 17092 27538
rect 17040 27474 17092 27480
rect 17224 27464 17276 27470
rect 17224 27406 17276 27412
rect 17040 27396 17092 27402
rect 17040 27338 17092 27344
rect 17052 25158 17080 27338
rect 17132 26444 17184 26450
rect 17132 26386 17184 26392
rect 17144 25838 17172 26386
rect 17132 25832 17184 25838
rect 17132 25774 17184 25780
rect 16672 25152 16724 25158
rect 16672 25094 16724 25100
rect 16948 25152 17000 25158
rect 16948 25094 17000 25100
rect 17040 25152 17092 25158
rect 17040 25094 17092 25100
rect 16580 24676 16632 24682
rect 16580 24618 16632 24624
rect 16120 24608 16172 24614
rect 16120 24550 16172 24556
rect 16132 23118 16160 24550
rect 16592 23186 16620 24618
rect 16684 24206 16712 25094
rect 16672 24200 16724 24206
rect 16672 24142 16724 24148
rect 17236 23186 17264 27406
rect 17328 27402 17356 29174
rect 18432 29102 18460 29514
rect 17960 29096 18012 29102
rect 17960 29038 18012 29044
rect 18420 29096 18472 29102
rect 18420 29038 18472 29044
rect 17500 29028 17552 29034
rect 17500 28970 17552 28976
rect 17408 28688 17460 28694
rect 17408 28630 17460 28636
rect 17420 27470 17448 28630
rect 17408 27464 17460 27470
rect 17408 27406 17460 27412
rect 17316 27396 17368 27402
rect 17316 27338 17368 27344
rect 17408 26920 17460 26926
rect 17408 26862 17460 26868
rect 17316 25696 17368 25702
rect 17316 25638 17368 25644
rect 17328 25362 17356 25638
rect 17316 25356 17368 25362
rect 17316 25298 17368 25304
rect 17316 25152 17368 25158
rect 17316 25094 17368 25100
rect 16488 23180 16540 23186
rect 16488 23122 16540 23128
rect 16580 23180 16632 23186
rect 16580 23122 16632 23128
rect 16672 23180 16724 23186
rect 16672 23122 16724 23128
rect 17224 23180 17276 23186
rect 17224 23122 17276 23128
rect 16120 23112 16172 23118
rect 16120 23054 16172 23060
rect 16132 22574 16160 23054
rect 16500 22574 16528 23122
rect 16684 22982 16712 23122
rect 16672 22976 16724 22982
rect 16672 22918 16724 22924
rect 16684 22574 16712 22918
rect 17236 22778 17264 23122
rect 17224 22772 17276 22778
rect 17224 22714 17276 22720
rect 17236 22574 17264 22714
rect 16120 22568 16172 22574
rect 16120 22510 16172 22516
rect 16488 22568 16540 22574
rect 16488 22510 16540 22516
rect 16672 22568 16724 22574
rect 17224 22568 17276 22574
rect 16724 22528 16804 22556
rect 16672 22510 16724 22516
rect 15948 22120 16068 22148
rect 15948 19310 15976 22120
rect 16500 21962 16528 22510
rect 16776 22098 16804 22528
rect 17224 22510 17276 22516
rect 17132 22500 17184 22506
rect 17132 22442 17184 22448
rect 16764 22092 16816 22098
rect 16948 22092 17000 22098
rect 16816 22052 16896 22080
rect 16764 22034 16816 22040
rect 16580 22024 16632 22030
rect 16580 21966 16632 21972
rect 16488 21956 16540 21962
rect 16488 21898 16540 21904
rect 16500 21418 16528 21898
rect 16592 21486 16620 21966
rect 16580 21480 16632 21486
rect 16580 21422 16632 21428
rect 16120 21412 16172 21418
rect 16120 21354 16172 21360
rect 16488 21412 16540 21418
rect 16488 21354 16540 21360
rect 16132 20398 16160 21354
rect 16868 21010 16896 22052
rect 16948 22034 17000 22040
rect 16960 21690 16988 22034
rect 16948 21684 17000 21690
rect 16948 21626 17000 21632
rect 17144 21486 17172 22442
rect 17236 22098 17264 22510
rect 17224 22092 17276 22098
rect 17224 22034 17276 22040
rect 17132 21480 17184 21486
rect 17132 21422 17184 21428
rect 17328 21010 17356 25094
rect 17420 22030 17448 26862
rect 17512 22642 17540 28970
rect 17972 28694 18000 29038
rect 17960 28688 18012 28694
rect 17960 28630 18012 28636
rect 18236 28620 18288 28626
rect 18236 28562 18288 28568
rect 18248 28082 18276 28562
rect 18328 28552 18380 28558
rect 18328 28494 18380 28500
rect 18236 28076 18288 28082
rect 18236 28018 18288 28024
rect 18340 28014 18368 28494
rect 17868 28008 17920 28014
rect 17868 27950 17920 27956
rect 18328 28008 18380 28014
rect 18328 27950 18380 27956
rect 17592 27940 17644 27946
rect 17592 27882 17644 27888
rect 17604 23866 17632 27882
rect 17880 27402 17908 27950
rect 17960 27600 18012 27606
rect 17960 27542 18012 27548
rect 17868 27396 17920 27402
rect 17868 27338 17920 27344
rect 17972 26994 18000 27542
rect 17960 26988 18012 26994
rect 17960 26930 18012 26936
rect 17868 26784 17920 26790
rect 17868 26726 17920 26732
rect 17880 26450 17908 26726
rect 17868 26444 17920 26450
rect 17868 26386 17920 26392
rect 17880 25362 17908 26386
rect 17972 25838 18000 26930
rect 18144 26444 18196 26450
rect 18144 26386 18196 26392
rect 18156 25838 18184 26386
rect 18340 26042 18368 27950
rect 18524 26586 18552 30194
rect 18800 29578 18828 31962
rect 18880 31884 18932 31890
rect 18880 31826 18932 31832
rect 18972 31884 19024 31890
rect 18972 31826 19024 31832
rect 18892 31278 18920 31826
rect 18984 31754 19012 31826
rect 18972 31748 19024 31754
rect 18972 31690 19024 31696
rect 18880 31272 18932 31278
rect 18880 31214 18932 31220
rect 18880 30796 18932 30802
rect 18880 30738 18932 30744
rect 18788 29572 18840 29578
rect 18708 29532 18788 29560
rect 18604 27328 18656 27334
rect 18604 27270 18656 27276
rect 18616 26926 18644 27270
rect 18604 26920 18656 26926
rect 18604 26862 18656 26868
rect 18512 26580 18564 26586
rect 18512 26522 18564 26528
rect 18708 26466 18736 29532
rect 18788 29514 18840 29520
rect 18788 29232 18840 29238
rect 18786 29200 18788 29209
rect 18840 29200 18842 29209
rect 18786 29135 18842 29144
rect 18788 26920 18840 26926
rect 18788 26862 18840 26868
rect 18432 26438 18736 26466
rect 18800 26450 18828 26862
rect 18788 26444 18840 26450
rect 18328 26036 18380 26042
rect 18328 25978 18380 25984
rect 17960 25832 18012 25838
rect 17960 25774 18012 25780
rect 18144 25832 18196 25838
rect 18144 25774 18196 25780
rect 18328 25832 18380 25838
rect 18328 25774 18380 25780
rect 18052 25492 18104 25498
rect 18052 25434 18104 25440
rect 17868 25356 17920 25362
rect 17868 25298 17920 25304
rect 17776 24268 17828 24274
rect 17776 24210 17828 24216
rect 17592 23860 17644 23866
rect 17592 23802 17644 23808
rect 17500 22636 17552 22642
rect 17500 22578 17552 22584
rect 17592 22092 17644 22098
rect 17592 22034 17644 22040
rect 17408 22024 17460 22030
rect 17408 21966 17460 21972
rect 17604 21146 17632 22034
rect 17592 21140 17644 21146
rect 17592 21082 17644 21088
rect 17604 21010 17632 21082
rect 16672 21004 16724 21010
rect 16672 20946 16724 20952
rect 16856 21004 16908 21010
rect 16856 20946 16908 20952
rect 17132 21004 17184 21010
rect 17132 20946 17184 20952
rect 17316 21004 17368 21010
rect 17316 20946 17368 20952
rect 17592 21004 17644 21010
rect 17592 20946 17644 20952
rect 16304 20596 16356 20602
rect 16304 20538 16356 20544
rect 16120 20392 16172 20398
rect 16316 20369 16344 20538
rect 16120 20334 16172 20340
rect 16302 20360 16358 20369
rect 16302 20295 16358 20304
rect 16212 19916 16264 19922
rect 16212 19858 16264 19864
rect 16224 19310 16252 19858
rect 16684 19854 16712 20946
rect 16868 19922 16896 20946
rect 17144 19922 17172 20946
rect 17224 20052 17276 20058
rect 17224 19994 17276 20000
rect 16856 19916 16908 19922
rect 16856 19858 16908 19864
rect 16948 19916 17000 19922
rect 16948 19858 17000 19864
rect 17132 19916 17184 19922
rect 17132 19858 17184 19864
rect 16672 19848 16724 19854
rect 16672 19790 16724 19796
rect 16960 19446 16988 19858
rect 17040 19508 17092 19514
rect 17040 19450 17092 19456
rect 16948 19440 17000 19446
rect 16948 19382 17000 19388
rect 15936 19304 15988 19310
rect 15936 19246 15988 19252
rect 16212 19304 16264 19310
rect 16212 19246 16264 19252
rect 15844 19168 15896 19174
rect 15844 19110 15896 19116
rect 15856 18834 15884 19110
rect 15844 18828 15896 18834
rect 15844 18770 15896 18776
rect 16224 18358 16252 19246
rect 16856 19168 16908 19174
rect 16856 19110 16908 19116
rect 16948 19168 17000 19174
rect 16948 19110 17000 19116
rect 16764 18760 16816 18766
rect 16764 18702 16816 18708
rect 16212 18352 16264 18358
rect 16212 18294 16264 18300
rect 16120 18284 16172 18290
rect 16120 18226 16172 18232
rect 15936 18080 15988 18086
rect 15936 18022 15988 18028
rect 15844 17740 15896 17746
rect 15844 17682 15896 17688
rect 15752 17536 15804 17542
rect 15752 17478 15804 17484
rect 15856 17338 15884 17682
rect 15844 17332 15896 17338
rect 15844 17274 15896 17280
rect 15660 16788 15712 16794
rect 15660 16730 15712 16736
rect 15844 16788 15896 16794
rect 15844 16730 15896 16736
rect 15660 14476 15712 14482
rect 15660 14418 15712 14424
rect 15488 14334 15608 14362
rect 15384 11892 15436 11898
rect 15384 11834 15436 11840
rect 15292 10600 15344 10606
rect 15292 10542 15344 10548
rect 15304 9722 15332 10542
rect 15488 10470 15516 14334
rect 15568 14000 15620 14006
rect 15568 13942 15620 13948
rect 15580 10674 15608 13942
rect 15568 10668 15620 10674
rect 15568 10610 15620 10616
rect 15476 10464 15528 10470
rect 15476 10406 15528 10412
rect 15488 9738 15516 10406
rect 15580 10198 15608 10610
rect 15568 10192 15620 10198
rect 15568 10134 15620 10140
rect 15292 9716 15344 9722
rect 15292 9658 15344 9664
rect 15396 9710 15516 9738
rect 15292 8968 15344 8974
rect 15292 8910 15344 8916
rect 15304 7206 15332 8910
rect 15292 7200 15344 7206
rect 15292 7142 15344 7148
rect 15292 5772 15344 5778
rect 15292 5714 15344 5720
rect 15200 5228 15252 5234
rect 15200 5170 15252 5176
rect 15016 5160 15068 5166
rect 15016 5102 15068 5108
rect 15028 4826 15056 5102
rect 15016 4820 15068 4826
rect 15016 4762 15068 4768
rect 15304 4146 15332 5714
rect 15292 4140 15344 4146
rect 15292 4082 15344 4088
rect 15396 4026 15424 9710
rect 15580 9602 15608 10134
rect 15488 9574 15608 9602
rect 15488 7954 15516 9574
rect 15568 9512 15620 9518
rect 15568 9454 15620 9460
rect 15580 8430 15608 9454
rect 15568 8424 15620 8430
rect 15568 8366 15620 8372
rect 15580 8294 15608 8366
rect 15568 8288 15620 8294
rect 15568 8230 15620 8236
rect 15476 7948 15528 7954
rect 15476 7890 15528 7896
rect 15580 7342 15608 8230
rect 15672 7834 15700 14418
rect 15752 13388 15804 13394
rect 15752 13330 15804 13336
rect 15764 13190 15792 13330
rect 15752 13184 15804 13190
rect 15752 13126 15804 13132
rect 15856 13138 15884 16730
rect 15948 16046 15976 18022
rect 16132 17202 16160 18226
rect 16212 17604 16264 17610
rect 16212 17546 16264 17552
rect 16224 17338 16252 17546
rect 16212 17332 16264 17338
rect 16212 17274 16264 17280
rect 16120 17196 16172 17202
rect 16120 17138 16172 17144
rect 16224 16794 16252 17274
rect 16212 16788 16264 16794
rect 16212 16730 16264 16736
rect 16776 16590 16804 18702
rect 16764 16584 16816 16590
rect 16764 16526 16816 16532
rect 16120 16176 16172 16182
rect 16120 16118 16172 16124
rect 15936 16040 15988 16046
rect 15988 16000 16068 16028
rect 15936 15982 15988 15988
rect 15936 14476 15988 14482
rect 15936 14418 15988 14424
rect 15948 13326 15976 14418
rect 15936 13320 15988 13326
rect 15936 13262 15988 13268
rect 15856 13110 15976 13138
rect 15844 12776 15896 12782
rect 15844 12718 15896 12724
rect 15856 11694 15884 12718
rect 15844 11688 15896 11694
rect 15844 11630 15896 11636
rect 15844 9376 15896 9382
rect 15844 9318 15896 9324
rect 15856 9110 15884 9318
rect 15844 9104 15896 9110
rect 15844 9046 15896 9052
rect 15672 7806 15884 7834
rect 15568 7336 15620 7342
rect 15568 7278 15620 7284
rect 15476 7200 15528 7206
rect 15476 7142 15528 7148
rect 15488 6866 15516 7142
rect 15476 6860 15528 6866
rect 15476 6802 15528 6808
rect 15580 6254 15608 7278
rect 15856 6458 15884 7806
rect 15844 6452 15896 6458
rect 15844 6394 15896 6400
rect 15568 6248 15620 6254
rect 15568 6190 15620 6196
rect 15580 5166 15608 6190
rect 15660 5636 15712 5642
rect 15660 5578 15712 5584
rect 15568 5160 15620 5166
rect 15568 5102 15620 5108
rect 15672 4690 15700 5578
rect 15856 5166 15884 6394
rect 15844 5160 15896 5166
rect 15844 5102 15896 5108
rect 15660 4684 15712 4690
rect 15660 4626 15712 4632
rect 15568 4480 15620 4486
rect 15568 4422 15620 4428
rect 15304 3998 15424 4026
rect 14832 3732 14884 3738
rect 14832 3674 14884 3680
rect 14188 3188 14240 3194
rect 14188 3130 14240 3136
rect 14844 3058 14872 3674
rect 15304 3534 15332 3998
rect 15292 3528 15344 3534
rect 15292 3470 15344 3476
rect 14924 3392 14976 3398
rect 14924 3334 14976 3340
rect 14832 3052 14884 3058
rect 14832 2994 14884 3000
rect 14936 2990 14964 3334
rect 15304 2990 15332 3470
rect 14188 2984 14240 2990
rect 14188 2926 14240 2932
rect 14924 2984 14976 2990
rect 14924 2926 14976 2932
rect 15292 2984 15344 2990
rect 15292 2926 15344 2932
rect 14096 2508 14148 2514
rect 14096 2450 14148 2456
rect 14200 2446 14228 2926
rect 15580 2582 15608 4422
rect 15948 2854 15976 13110
rect 16040 10674 16068 16000
rect 16132 15706 16160 16118
rect 16120 15700 16172 15706
rect 16120 15642 16172 15648
rect 16132 14006 16160 15642
rect 16776 15570 16804 16526
rect 16764 15564 16816 15570
rect 16764 15506 16816 15512
rect 16304 15496 16356 15502
rect 16304 15438 16356 15444
rect 16212 14340 16264 14346
rect 16212 14282 16264 14288
rect 16120 14000 16172 14006
rect 16120 13942 16172 13948
rect 16120 13388 16172 13394
rect 16120 13330 16172 13336
rect 16132 11830 16160 13330
rect 16120 11824 16172 11830
rect 16120 11766 16172 11772
rect 16224 11150 16252 14282
rect 16316 11694 16344 15438
rect 16776 14958 16804 15506
rect 16764 14952 16816 14958
rect 16764 14894 16816 14900
rect 16776 14346 16804 14894
rect 16764 14340 16816 14346
rect 16764 14282 16816 14288
rect 16580 14000 16632 14006
rect 16580 13942 16632 13948
rect 16592 12850 16620 13942
rect 16764 13864 16816 13870
rect 16764 13806 16816 13812
rect 16672 13728 16724 13734
rect 16672 13670 16724 13676
rect 16684 13002 16712 13670
rect 16776 13394 16804 13806
rect 16764 13388 16816 13394
rect 16764 13330 16816 13336
rect 16684 12986 16804 13002
rect 16684 12980 16816 12986
rect 16684 12974 16764 12980
rect 16580 12844 16632 12850
rect 16580 12786 16632 12792
rect 16684 12730 16712 12974
rect 16764 12922 16816 12928
rect 16592 12702 16712 12730
rect 16592 11830 16620 12702
rect 16762 12336 16818 12345
rect 16762 12271 16818 12280
rect 16580 11824 16632 11830
rect 16580 11766 16632 11772
rect 16304 11688 16356 11694
rect 16304 11630 16356 11636
rect 16316 11354 16344 11630
rect 16304 11348 16356 11354
rect 16304 11290 16356 11296
rect 16212 11144 16264 11150
rect 16212 11086 16264 11092
rect 16776 10810 16804 12271
rect 16764 10804 16816 10810
rect 16764 10746 16816 10752
rect 16028 10668 16080 10674
rect 16028 10610 16080 10616
rect 16040 10062 16068 10610
rect 16212 10600 16264 10606
rect 16212 10542 16264 10548
rect 16028 10056 16080 10062
rect 16028 9998 16080 10004
rect 16040 8430 16068 9998
rect 16120 9988 16172 9994
rect 16120 9930 16172 9936
rect 16132 9042 16160 9930
rect 16120 9036 16172 9042
rect 16120 8978 16172 8984
rect 16224 8634 16252 10542
rect 16488 10124 16540 10130
rect 16488 10066 16540 10072
rect 16304 8968 16356 8974
rect 16304 8910 16356 8916
rect 16212 8628 16264 8634
rect 16212 8570 16264 8576
rect 16028 8424 16080 8430
rect 16028 8366 16080 8372
rect 16224 7954 16252 8570
rect 16212 7948 16264 7954
rect 16212 7890 16264 7896
rect 16028 7744 16080 7750
rect 16028 7686 16080 7692
rect 15936 2848 15988 2854
rect 15936 2790 15988 2796
rect 15568 2576 15620 2582
rect 15568 2518 15620 2524
rect 16040 2514 16068 7686
rect 16316 5778 16344 8910
rect 16304 5772 16356 5778
rect 16304 5714 16356 5720
rect 16212 5160 16264 5166
rect 16212 5102 16264 5108
rect 16396 5160 16448 5166
rect 16396 5102 16448 5108
rect 16224 4554 16252 5102
rect 16304 4616 16356 4622
rect 16304 4558 16356 4564
rect 16212 4548 16264 4554
rect 16212 4490 16264 4496
rect 16316 4078 16344 4558
rect 16408 4214 16436 5102
rect 16500 4486 16528 10066
rect 16764 9920 16816 9926
rect 16764 9862 16816 9868
rect 16670 9616 16726 9625
rect 16670 9551 16726 9560
rect 16684 9518 16712 9551
rect 16580 9512 16632 9518
rect 16580 9454 16632 9460
rect 16672 9512 16724 9518
rect 16672 9454 16724 9460
rect 16592 7818 16620 9454
rect 16776 8430 16804 9862
rect 16764 8424 16816 8430
rect 16764 8366 16816 8372
rect 16868 8022 16896 19110
rect 16960 18834 16988 19110
rect 16948 18828 17000 18834
rect 16948 18770 17000 18776
rect 16960 18222 16988 18770
rect 17052 18222 17080 19450
rect 17236 19310 17264 19994
rect 17328 19990 17356 20946
rect 17500 20392 17552 20398
rect 17500 20334 17552 20340
rect 17316 19984 17368 19990
rect 17316 19926 17368 19932
rect 17512 19922 17540 20334
rect 17788 20058 17816 24210
rect 17880 23186 17908 25298
rect 17868 23180 17920 23186
rect 17868 23122 17920 23128
rect 17880 22166 17908 23122
rect 18064 22574 18092 25434
rect 18156 25362 18184 25774
rect 18340 25430 18368 25774
rect 18328 25424 18380 25430
rect 18328 25366 18380 25372
rect 18144 25356 18196 25362
rect 18144 25298 18196 25304
rect 18328 24744 18380 24750
rect 18328 24686 18380 24692
rect 18340 24274 18368 24686
rect 18328 24268 18380 24274
rect 18328 24210 18380 24216
rect 18340 24138 18368 24210
rect 18328 24132 18380 24138
rect 18328 24074 18380 24080
rect 18340 23730 18368 24074
rect 18328 23724 18380 23730
rect 18328 23666 18380 23672
rect 18144 23112 18196 23118
rect 18144 23054 18196 23060
rect 18052 22568 18104 22574
rect 18052 22510 18104 22516
rect 17868 22160 17920 22166
rect 17868 22102 17920 22108
rect 18156 21690 18184 23054
rect 18144 21684 18196 21690
rect 18144 21626 18196 21632
rect 17776 20052 17828 20058
rect 17776 19994 17828 20000
rect 17500 19916 17552 19922
rect 17500 19858 17552 19864
rect 17684 19916 17736 19922
rect 17684 19858 17736 19864
rect 17512 19786 17540 19858
rect 17500 19780 17552 19786
rect 17500 19722 17552 19728
rect 17512 19310 17540 19722
rect 17696 19310 17724 19858
rect 18144 19848 18196 19854
rect 18144 19790 18196 19796
rect 17224 19304 17276 19310
rect 17224 19246 17276 19252
rect 17500 19304 17552 19310
rect 17500 19246 17552 19252
rect 17684 19304 17736 19310
rect 17684 19246 17736 19252
rect 17316 18828 17368 18834
rect 17316 18770 17368 18776
rect 17328 18290 17356 18770
rect 17500 18692 17552 18698
rect 17500 18634 17552 18640
rect 17316 18284 17368 18290
rect 17316 18226 17368 18232
rect 16948 18216 17000 18222
rect 16948 18158 17000 18164
rect 17040 18216 17092 18222
rect 17040 18158 17092 18164
rect 17040 17604 17092 17610
rect 17040 17546 17092 17552
rect 17052 16658 17080 17546
rect 17328 17134 17356 18226
rect 17316 17128 17368 17134
rect 17316 17070 17368 17076
rect 17224 16992 17276 16998
rect 17224 16934 17276 16940
rect 17040 16652 17092 16658
rect 17040 16594 17092 16600
rect 17040 15020 17092 15026
rect 17040 14962 17092 14968
rect 16948 14952 17000 14958
rect 16948 14894 17000 14900
rect 16960 13802 16988 14894
rect 16948 13796 17000 13802
rect 16948 13738 17000 13744
rect 16948 13524 17000 13530
rect 16948 13466 17000 13472
rect 16856 8016 16908 8022
rect 16856 7958 16908 7964
rect 16580 7812 16632 7818
rect 16580 7754 16632 7760
rect 16592 7206 16620 7754
rect 16672 7336 16724 7342
rect 16672 7278 16724 7284
rect 16580 7200 16632 7206
rect 16580 7142 16632 7148
rect 16684 6390 16712 7278
rect 16764 6656 16816 6662
rect 16764 6598 16816 6604
rect 16672 6384 16724 6390
rect 16672 6326 16724 6332
rect 16580 5024 16632 5030
rect 16580 4966 16632 4972
rect 16592 4690 16620 4966
rect 16580 4684 16632 4690
rect 16580 4626 16632 4632
rect 16488 4480 16540 4486
rect 16488 4422 16540 4428
rect 16396 4208 16448 4214
rect 16396 4150 16448 4156
rect 16684 4078 16712 6326
rect 16776 6186 16804 6598
rect 16868 6254 16896 7958
rect 16960 7342 16988 13466
rect 16948 7336 17000 7342
rect 16948 7278 17000 7284
rect 16856 6248 16908 6254
rect 16856 6190 16908 6196
rect 16764 6180 16816 6186
rect 16764 6122 16816 6128
rect 16776 5166 16804 6122
rect 16868 5914 16896 6190
rect 16856 5908 16908 5914
rect 16856 5850 16908 5856
rect 17052 5778 17080 14962
rect 17132 14816 17184 14822
rect 17132 14758 17184 14764
rect 17144 14482 17172 14758
rect 17132 14476 17184 14482
rect 17132 14418 17184 14424
rect 17236 13530 17264 16934
rect 17512 15162 17540 18634
rect 17684 18148 17736 18154
rect 17684 18090 17736 18096
rect 17776 18148 17828 18154
rect 17776 18090 17828 18096
rect 17500 15156 17552 15162
rect 17500 15098 17552 15104
rect 17408 14816 17460 14822
rect 17408 14758 17460 14764
rect 17224 13524 17276 13530
rect 17224 13466 17276 13472
rect 17132 13184 17184 13190
rect 17132 13126 17184 13132
rect 17144 12714 17172 13126
rect 17132 12708 17184 12714
rect 17132 12650 17184 12656
rect 17132 12436 17184 12442
rect 17132 12378 17184 12384
rect 17144 10810 17172 12378
rect 17420 12306 17448 14758
rect 17408 12300 17460 12306
rect 17408 12242 17460 12248
rect 17224 12232 17276 12238
rect 17224 12174 17276 12180
rect 17236 11694 17264 12174
rect 17224 11688 17276 11694
rect 17224 11630 17276 11636
rect 17132 10804 17184 10810
rect 17132 10746 17184 10752
rect 17224 10736 17276 10742
rect 17276 10684 17448 10690
rect 17224 10678 17448 10684
rect 17236 10674 17448 10678
rect 17236 10668 17460 10674
rect 17236 10662 17408 10668
rect 17408 10610 17460 10616
rect 17512 10606 17540 15098
rect 17316 10600 17368 10606
rect 17316 10542 17368 10548
rect 17500 10600 17552 10606
rect 17500 10542 17552 10548
rect 17132 10532 17184 10538
rect 17132 10474 17184 10480
rect 17144 9518 17172 10474
rect 17224 10464 17276 10470
rect 17224 10406 17276 10412
rect 17236 10266 17264 10406
rect 17224 10260 17276 10266
rect 17224 10202 17276 10208
rect 17328 9926 17356 10542
rect 17408 9988 17460 9994
rect 17408 9930 17460 9936
rect 17316 9920 17368 9926
rect 17420 9897 17448 9930
rect 17316 9862 17368 9868
rect 17406 9888 17462 9897
rect 17406 9823 17462 9832
rect 17132 9512 17184 9518
rect 17132 9454 17184 9460
rect 17224 9104 17276 9110
rect 17224 9046 17276 9052
rect 17236 8566 17264 9046
rect 17224 8560 17276 8566
rect 17224 8502 17276 8508
rect 17696 8090 17724 18090
rect 17788 16590 17816 18090
rect 18052 17740 18104 17746
rect 18052 17682 18104 17688
rect 17776 16584 17828 16590
rect 17776 16526 17828 16532
rect 17960 16448 18012 16454
rect 17960 16390 18012 16396
rect 17972 16046 18000 16390
rect 18064 16182 18092 17682
rect 18052 16176 18104 16182
rect 18052 16118 18104 16124
rect 17960 16040 18012 16046
rect 17960 15982 18012 15988
rect 17972 12306 18000 15982
rect 18052 14884 18104 14890
rect 18052 14826 18104 14832
rect 18064 13870 18092 14826
rect 18156 14482 18184 19790
rect 18432 18834 18460 26438
rect 18788 26386 18840 26392
rect 18892 25226 18920 30738
rect 19076 29714 19104 32778
rect 19168 32502 19196 32778
rect 19156 32496 19208 32502
rect 19156 32438 19208 32444
rect 19340 32360 19392 32366
rect 19340 32302 19392 32308
rect 19154 32192 19210 32201
rect 19154 32127 19210 32136
rect 19168 32042 19196 32127
rect 19352 32042 19380 32302
rect 19580 32124 19876 32144
rect 19636 32122 19660 32124
rect 19716 32122 19740 32124
rect 19796 32122 19820 32124
rect 19658 32070 19660 32122
rect 19722 32070 19734 32122
rect 19796 32070 19798 32122
rect 19636 32068 19660 32070
rect 19716 32068 19740 32070
rect 19796 32068 19820 32070
rect 19580 32048 19876 32068
rect 19168 32014 19380 32042
rect 19432 32020 19484 32026
rect 19432 31962 19484 31968
rect 19248 31952 19300 31958
rect 19248 31894 19300 31900
rect 19338 31920 19394 31929
rect 19156 30184 19208 30190
rect 19156 30126 19208 30132
rect 19064 29708 19116 29714
rect 19064 29650 19116 29656
rect 19168 28762 19196 30126
rect 19156 28756 19208 28762
rect 19156 28698 19208 28704
rect 18972 28620 19024 28626
rect 19024 28580 19196 28608
rect 18972 28562 19024 28568
rect 19168 28014 19196 28580
rect 19156 28008 19208 28014
rect 19156 27950 19208 27956
rect 19168 26994 19196 27950
rect 19156 26988 19208 26994
rect 19156 26930 19208 26936
rect 19168 26790 19196 26930
rect 19156 26784 19208 26790
rect 19156 26726 19208 26732
rect 19168 26450 19196 26726
rect 19156 26444 19208 26450
rect 19156 26386 19208 26392
rect 19156 25356 19208 25362
rect 19156 25298 19208 25304
rect 18880 25220 18932 25226
rect 18880 25162 18932 25168
rect 18788 24608 18840 24614
rect 18788 24550 18840 24556
rect 18800 24274 18828 24550
rect 18788 24268 18840 24274
rect 18788 24210 18840 24216
rect 18696 24200 18748 24206
rect 18696 24142 18748 24148
rect 18708 23662 18736 24142
rect 18800 23662 18828 24210
rect 18892 23866 18920 25162
rect 19168 24818 19196 25298
rect 19156 24812 19208 24818
rect 19156 24754 19208 24760
rect 19156 24676 19208 24682
rect 19156 24618 19208 24624
rect 19168 24342 19196 24618
rect 18972 24336 19024 24342
rect 18972 24278 19024 24284
rect 19156 24336 19208 24342
rect 19156 24278 19208 24284
rect 18880 23860 18932 23866
rect 18880 23802 18932 23808
rect 18696 23656 18748 23662
rect 18696 23598 18748 23604
rect 18788 23656 18840 23662
rect 18788 23598 18840 23604
rect 18604 23180 18656 23186
rect 18708 23168 18736 23598
rect 18800 23186 18828 23598
rect 18656 23140 18736 23168
rect 18604 23122 18656 23128
rect 18708 22166 18736 23140
rect 18788 23180 18840 23186
rect 18788 23122 18840 23128
rect 18800 22574 18828 23122
rect 18984 22778 19012 24278
rect 19064 24268 19116 24274
rect 19064 24210 19116 24216
rect 18972 22772 19024 22778
rect 18972 22714 19024 22720
rect 18788 22568 18840 22574
rect 18788 22510 18840 22516
rect 18984 22386 19012 22714
rect 18800 22358 19012 22386
rect 18696 22160 18748 22166
rect 18696 22102 18748 22108
rect 18604 20596 18656 20602
rect 18604 20538 18656 20544
rect 18512 20324 18564 20330
rect 18512 20266 18564 20272
rect 18524 19854 18552 20266
rect 18616 19922 18644 20538
rect 18800 20330 18828 22358
rect 18972 22228 19024 22234
rect 18972 22170 19024 22176
rect 18984 22030 19012 22170
rect 18972 22024 19024 22030
rect 18972 21966 19024 21972
rect 18880 20936 18932 20942
rect 18880 20878 18932 20884
rect 18788 20324 18840 20330
rect 18788 20266 18840 20272
rect 18696 20256 18748 20262
rect 18696 20198 18748 20204
rect 18604 19916 18656 19922
rect 18604 19858 18656 19864
rect 18512 19848 18564 19854
rect 18708 19802 18736 20198
rect 18788 19848 18840 19854
rect 18512 19790 18564 19796
rect 18616 19796 18788 19802
rect 18616 19790 18840 19796
rect 18524 19514 18552 19790
rect 18616 19774 18828 19790
rect 18512 19508 18564 19514
rect 18512 19450 18564 19456
rect 18420 18828 18472 18834
rect 18420 18770 18472 18776
rect 18432 18222 18460 18770
rect 18420 18216 18472 18222
rect 18420 18158 18472 18164
rect 18328 17128 18380 17134
rect 18328 17070 18380 17076
rect 18340 16250 18368 17070
rect 18328 16244 18380 16250
rect 18328 16186 18380 16192
rect 18420 16040 18472 16046
rect 18420 15982 18472 15988
rect 18432 15638 18460 15982
rect 18420 15632 18472 15638
rect 18420 15574 18472 15580
rect 18328 15020 18380 15026
rect 18328 14962 18380 14968
rect 18236 14952 18288 14958
rect 18236 14894 18288 14900
rect 18144 14476 18196 14482
rect 18144 14418 18196 14424
rect 18052 13864 18104 13870
rect 18052 13806 18104 13812
rect 18248 13682 18276 14894
rect 18340 14482 18368 14962
rect 18328 14476 18380 14482
rect 18328 14418 18380 14424
rect 18512 13932 18564 13938
rect 18512 13874 18564 13880
rect 18420 13864 18472 13870
rect 18420 13806 18472 13812
rect 18248 13654 18368 13682
rect 18236 13320 18288 13326
rect 18236 13262 18288 13268
rect 18144 12844 18196 12850
rect 18144 12786 18196 12792
rect 18052 12776 18104 12782
rect 18052 12718 18104 12724
rect 18064 12374 18092 12718
rect 18052 12368 18104 12374
rect 18052 12310 18104 12316
rect 17960 12300 18012 12306
rect 17960 12242 18012 12248
rect 17960 11688 18012 11694
rect 17960 11630 18012 11636
rect 17776 11620 17828 11626
rect 17776 11562 17828 11568
rect 17788 11082 17816 11562
rect 17972 11218 18000 11630
rect 17960 11212 18012 11218
rect 17960 11154 18012 11160
rect 17776 11076 17828 11082
rect 17776 11018 17828 11024
rect 17972 10538 18000 11154
rect 18052 11008 18104 11014
rect 18052 10950 18104 10956
rect 17960 10532 18012 10538
rect 17960 10474 18012 10480
rect 18064 9586 18092 10950
rect 18052 9580 18104 9586
rect 18052 9522 18104 9528
rect 17868 9512 17920 9518
rect 17868 9454 17920 9460
rect 17684 8084 17736 8090
rect 17684 8026 17736 8032
rect 17500 7812 17552 7818
rect 17500 7754 17552 7760
rect 17512 6866 17540 7754
rect 17500 6860 17552 6866
rect 17500 6802 17552 6808
rect 17696 5778 17724 8026
rect 17776 6112 17828 6118
rect 17776 6054 17828 6060
rect 17040 5772 17092 5778
rect 17040 5714 17092 5720
rect 17684 5772 17736 5778
rect 17684 5714 17736 5720
rect 16764 5160 16816 5166
rect 16764 5102 16816 5108
rect 17052 4078 17080 5714
rect 17224 5704 17276 5710
rect 17224 5646 17276 5652
rect 16304 4072 16356 4078
rect 16304 4014 16356 4020
rect 16672 4072 16724 4078
rect 16672 4014 16724 4020
rect 17040 4072 17092 4078
rect 17040 4014 17092 4020
rect 16120 3936 16172 3942
rect 16120 3878 16172 3884
rect 16132 3058 16160 3878
rect 16316 3534 16344 4014
rect 17052 3738 17080 4014
rect 17040 3732 17092 3738
rect 17040 3674 17092 3680
rect 17236 3602 17264 5646
rect 17788 4486 17816 6054
rect 17880 5710 17908 9454
rect 18156 9178 18184 12786
rect 18248 12374 18276 13262
rect 18236 12368 18288 12374
rect 18236 12310 18288 12316
rect 18236 12232 18288 12238
rect 18236 12174 18288 12180
rect 18248 11898 18276 12174
rect 18236 11892 18288 11898
rect 18236 11834 18288 11840
rect 18248 11354 18276 11834
rect 18236 11348 18288 11354
rect 18236 11290 18288 11296
rect 18340 11286 18368 13654
rect 18432 12782 18460 13806
rect 18524 13394 18552 13874
rect 18512 13388 18564 13394
rect 18512 13330 18564 13336
rect 18420 12776 18472 12782
rect 18420 12718 18472 12724
rect 18328 11280 18380 11286
rect 18328 11222 18380 11228
rect 18236 10464 18288 10470
rect 18236 10406 18288 10412
rect 18248 10130 18276 10406
rect 18236 10124 18288 10130
rect 18236 10066 18288 10072
rect 18328 9920 18380 9926
rect 18328 9862 18380 9868
rect 18144 9172 18196 9178
rect 18144 9114 18196 9120
rect 18156 9058 18184 9114
rect 18064 9030 18184 9058
rect 17960 7948 18012 7954
rect 17960 7890 18012 7896
rect 17972 7274 18000 7890
rect 17960 7268 18012 7274
rect 17960 7210 18012 7216
rect 17972 5914 18000 7210
rect 18064 6254 18092 9030
rect 18236 8424 18288 8430
rect 18236 8366 18288 8372
rect 18144 7948 18196 7954
rect 18144 7890 18196 7896
rect 18156 7478 18184 7890
rect 18144 7472 18196 7478
rect 18144 7414 18196 7420
rect 18156 7002 18184 7414
rect 18248 7002 18276 8366
rect 18144 6996 18196 7002
rect 18144 6938 18196 6944
rect 18236 6996 18288 7002
rect 18236 6938 18288 6944
rect 18248 6798 18276 6938
rect 18340 6866 18368 9862
rect 18616 9518 18644 19774
rect 18788 19304 18840 19310
rect 18788 19246 18840 19252
rect 18800 18834 18828 19246
rect 18788 18828 18840 18834
rect 18788 18770 18840 18776
rect 18800 17746 18828 18770
rect 18788 17740 18840 17746
rect 18788 17682 18840 17688
rect 18696 17672 18748 17678
rect 18892 17626 18920 20878
rect 19076 20806 19104 24210
rect 19156 23656 19208 23662
rect 19156 23598 19208 23604
rect 19168 23186 19196 23598
rect 19156 23180 19208 23186
rect 19156 23122 19208 23128
rect 19168 22234 19196 23122
rect 19156 22228 19208 22234
rect 19156 22170 19208 22176
rect 19156 21480 19208 21486
rect 19156 21422 19208 21428
rect 19168 21078 19196 21422
rect 19156 21072 19208 21078
rect 19156 21014 19208 21020
rect 19064 20800 19116 20806
rect 19064 20742 19116 20748
rect 19064 20460 19116 20466
rect 19064 20402 19116 20408
rect 19076 18970 19104 20402
rect 19156 19508 19208 19514
rect 19156 19450 19208 19456
rect 19064 18964 19116 18970
rect 19064 18906 19116 18912
rect 18972 18692 19024 18698
rect 18972 18634 19024 18640
rect 18696 17614 18748 17620
rect 18708 10198 18736 17614
rect 18800 17598 18920 17626
rect 18800 15910 18828 17598
rect 18788 15904 18840 15910
rect 18788 15846 18840 15852
rect 18800 15638 18828 15846
rect 18788 15632 18840 15638
rect 18788 15574 18840 15580
rect 18800 12646 18828 15574
rect 18984 15570 19012 18634
rect 19076 17542 19104 18906
rect 19168 18358 19196 19450
rect 19156 18352 19208 18358
rect 19156 18294 19208 18300
rect 19156 18216 19208 18222
rect 19154 18184 19156 18193
rect 19208 18184 19210 18193
rect 19154 18119 19210 18128
rect 19156 17604 19208 17610
rect 19156 17546 19208 17552
rect 19064 17536 19116 17542
rect 19064 17478 19116 17484
rect 19076 17270 19104 17478
rect 19064 17264 19116 17270
rect 19064 17206 19116 17212
rect 19168 16658 19196 17546
rect 19156 16652 19208 16658
rect 19156 16594 19208 16600
rect 18972 15564 19024 15570
rect 18972 15506 19024 15512
rect 19156 15564 19208 15570
rect 19156 15506 19208 15512
rect 18880 15496 18932 15502
rect 18880 15438 18932 15444
rect 18788 12640 18840 12646
rect 18788 12582 18840 12588
rect 18892 12442 18920 15438
rect 19168 14414 19196 15506
rect 19156 14408 19208 14414
rect 19156 14350 19208 14356
rect 19156 14272 19208 14278
rect 19156 14214 19208 14220
rect 19168 13938 19196 14214
rect 19156 13932 19208 13938
rect 19156 13874 19208 13880
rect 19156 13252 19208 13258
rect 19156 13194 19208 13200
rect 19168 12850 19196 13194
rect 19260 12918 19288 31894
rect 19444 31890 19472 31962
rect 19338 31855 19340 31864
rect 19392 31855 19394 31864
rect 19432 31884 19484 31890
rect 19340 31826 19392 31832
rect 19432 31826 19484 31832
rect 19800 31748 19852 31754
rect 19800 31690 19852 31696
rect 19812 31278 19840 31690
rect 19904 31482 19932 33390
rect 19996 32978 20024 33798
rect 20076 33312 20128 33318
rect 20076 33254 20128 33260
rect 19984 32972 20036 32978
rect 19984 32914 20036 32920
rect 19984 32564 20036 32570
rect 19984 32506 20036 32512
rect 19996 31890 20024 32506
rect 20088 32434 20116 33254
rect 20180 33114 20208 34410
rect 20272 33658 20300 35090
rect 20548 34542 20576 36178
rect 20628 36168 20680 36174
rect 20628 36110 20680 36116
rect 20640 35698 20668 36110
rect 20732 36106 20760 38286
rect 21008 37466 21036 38354
rect 21180 37664 21232 37670
rect 21180 37606 21232 37612
rect 20996 37460 21048 37466
rect 20996 37402 21048 37408
rect 20902 37360 20958 37369
rect 20902 37295 20904 37304
rect 20956 37295 20958 37304
rect 20904 37266 20956 37272
rect 20916 36242 20944 37266
rect 21192 36718 21220 37606
rect 21560 36922 21588 38354
rect 21824 38276 21876 38282
rect 21824 38218 21876 38224
rect 21640 38208 21692 38214
rect 21640 38150 21692 38156
rect 21652 37330 21680 38150
rect 21732 37732 21784 37738
rect 21732 37674 21784 37680
rect 21744 37466 21772 37674
rect 21836 37466 21864 38218
rect 22112 38010 22140 40200
rect 22284 38412 22336 38418
rect 22284 38354 22336 38360
rect 22100 38004 22152 38010
rect 22100 37946 22152 37952
rect 21732 37460 21784 37466
rect 21732 37402 21784 37408
rect 21824 37460 21876 37466
rect 21824 37402 21876 37408
rect 22296 37398 22324 38354
rect 22468 37868 22520 37874
rect 22468 37810 22520 37816
rect 22480 37670 22508 37810
rect 22652 37800 22704 37806
rect 22652 37742 22704 37748
rect 23388 37800 23440 37806
rect 23388 37742 23440 37748
rect 22468 37664 22520 37670
rect 22468 37606 22520 37612
rect 22284 37392 22336 37398
rect 22284 37334 22336 37340
rect 21640 37324 21692 37330
rect 21640 37266 21692 37272
rect 21916 37256 21968 37262
rect 21916 37198 21968 37204
rect 21548 36916 21600 36922
rect 21548 36858 21600 36864
rect 21272 36848 21324 36854
rect 21272 36790 21324 36796
rect 21180 36712 21232 36718
rect 21180 36654 21232 36660
rect 20904 36236 20956 36242
rect 20904 36178 20956 36184
rect 20720 36100 20772 36106
rect 20720 36042 20772 36048
rect 20628 35692 20680 35698
rect 20628 35634 20680 35640
rect 20904 35556 20956 35562
rect 20904 35498 20956 35504
rect 20916 35222 20944 35498
rect 20904 35216 20956 35222
rect 20904 35158 20956 35164
rect 21192 35204 21220 36654
rect 21284 36242 21312 36790
rect 21928 36718 21956 37198
rect 21916 36712 21968 36718
rect 21730 36680 21786 36689
rect 21916 36654 21968 36660
rect 21730 36615 21786 36624
rect 21272 36236 21324 36242
rect 21272 36178 21324 36184
rect 21364 35760 21416 35766
rect 21364 35702 21416 35708
rect 21272 35216 21324 35222
rect 21192 35176 21272 35204
rect 20720 35148 20772 35154
rect 20640 35108 20720 35136
rect 20536 34536 20588 34542
rect 20536 34478 20588 34484
rect 20640 34474 20668 35108
rect 20720 35090 20772 35096
rect 20996 35080 21048 35086
rect 20996 35022 21048 35028
rect 21008 34610 21036 35022
rect 20996 34604 21048 34610
rect 20996 34546 21048 34552
rect 20628 34468 20680 34474
rect 20628 34410 20680 34416
rect 21192 34066 21220 35176
rect 21272 35158 21324 35164
rect 21376 34066 21404 35702
rect 21640 35624 21692 35630
rect 21640 35566 21692 35572
rect 21652 35290 21680 35566
rect 21640 35284 21692 35290
rect 21640 35226 21692 35232
rect 21456 35148 21508 35154
rect 21456 35090 21508 35096
rect 21468 34542 21496 35090
rect 21456 34536 21508 34542
rect 21456 34478 21508 34484
rect 21548 34400 21600 34406
rect 21548 34342 21600 34348
rect 21180 34060 21232 34066
rect 21180 34002 21232 34008
rect 21364 34060 21416 34066
rect 21364 34002 21416 34008
rect 20260 33652 20312 33658
rect 20260 33594 20312 33600
rect 20168 33108 20220 33114
rect 20168 33050 20220 33056
rect 20272 32910 20300 33594
rect 20260 32904 20312 32910
rect 20260 32846 20312 32852
rect 21192 32434 21220 34002
rect 21376 33454 21404 34002
rect 21560 33522 21588 34342
rect 21652 34066 21680 35226
rect 21640 34060 21692 34066
rect 21640 34002 21692 34008
rect 21744 33946 21772 36615
rect 21824 35760 21876 35766
rect 21824 35702 21876 35708
rect 21836 35630 21864 35702
rect 21928 35698 21956 36654
rect 21916 35692 21968 35698
rect 21916 35634 21968 35640
rect 21824 35624 21876 35630
rect 21824 35566 21876 35572
rect 22008 35624 22060 35630
rect 22008 35566 22060 35572
rect 22020 35222 22048 35566
rect 22480 35290 22508 37606
rect 22664 37194 22692 37742
rect 23400 37670 23428 37742
rect 23756 37732 23808 37738
rect 23756 37674 23808 37680
rect 23388 37664 23440 37670
rect 23388 37606 23440 37612
rect 23480 37664 23532 37670
rect 23480 37606 23532 37612
rect 22926 37360 22982 37369
rect 23204 37324 23256 37330
rect 22982 37304 23152 37312
rect 22926 37295 22928 37304
rect 22980 37284 23152 37304
rect 22928 37266 22980 37272
rect 22652 37188 22704 37194
rect 22652 37130 22704 37136
rect 22836 36236 22888 36242
rect 22836 36178 22888 36184
rect 22560 36032 22612 36038
rect 22560 35974 22612 35980
rect 22572 35562 22600 35974
rect 22652 35624 22704 35630
rect 22652 35566 22704 35572
rect 22560 35556 22612 35562
rect 22560 35498 22612 35504
rect 22468 35284 22520 35290
rect 22468 35226 22520 35232
rect 22008 35216 22060 35222
rect 22008 35158 22060 35164
rect 22664 35154 22692 35566
rect 22560 35148 22612 35154
rect 22560 35090 22612 35096
rect 22652 35148 22704 35154
rect 22652 35090 22704 35096
rect 22100 34468 22152 34474
rect 22100 34410 22152 34416
rect 22112 34066 22140 34410
rect 22572 34116 22600 35090
rect 22848 35086 22876 36178
rect 23124 35154 23152 37284
rect 23204 37266 23256 37272
rect 23388 37324 23440 37330
rect 23388 37266 23440 37272
rect 23216 37194 23244 37266
rect 23204 37188 23256 37194
rect 23204 37130 23256 37136
rect 23216 35154 23244 37130
rect 23400 35834 23428 37266
rect 23492 37262 23520 37606
rect 23768 37330 23796 37674
rect 23572 37324 23624 37330
rect 23572 37266 23624 37272
rect 23756 37324 23808 37330
rect 23756 37266 23808 37272
rect 23480 37256 23532 37262
rect 23480 37198 23532 37204
rect 23492 36718 23520 37198
rect 23480 36712 23532 36718
rect 23480 36654 23532 36660
rect 23584 36650 23612 37266
rect 23952 36786 23980 40200
rect 25976 38842 26004 40200
rect 25976 38814 26188 38842
rect 26160 38570 26188 38814
rect 26160 38542 26280 38570
rect 26252 38486 26280 38542
rect 26240 38480 26292 38486
rect 26240 38422 26292 38428
rect 24952 38344 25004 38350
rect 24952 38286 25004 38292
rect 27436 38344 27488 38350
rect 27436 38286 27488 38292
rect 24860 38208 24912 38214
rect 24860 38150 24912 38156
rect 24308 38004 24360 38010
rect 24308 37946 24360 37952
rect 23940 36780 23992 36786
rect 23940 36722 23992 36728
rect 24320 36718 24348 37946
rect 24872 37806 24900 38150
rect 24860 37800 24912 37806
rect 24860 37742 24912 37748
rect 24872 37330 24900 37742
rect 24860 37324 24912 37330
rect 24860 37266 24912 37272
rect 24124 36712 24176 36718
rect 24124 36654 24176 36660
rect 24308 36712 24360 36718
rect 24308 36654 24360 36660
rect 23572 36644 23624 36650
rect 23572 36586 23624 36592
rect 23388 35828 23440 35834
rect 23388 35770 23440 35776
rect 23112 35148 23164 35154
rect 23032 35108 23112 35136
rect 22836 35080 22888 35086
rect 22836 35022 22888 35028
rect 22836 34536 22888 34542
rect 22836 34478 22888 34484
rect 22652 34128 22704 34134
rect 22572 34088 22652 34116
rect 22652 34070 22704 34076
rect 22100 34060 22152 34066
rect 22100 34002 22152 34008
rect 21744 33918 21956 33946
rect 21548 33516 21600 33522
rect 21548 33458 21600 33464
rect 21364 33448 21416 33454
rect 21364 33390 21416 33396
rect 20076 32428 20128 32434
rect 20076 32370 20128 32376
rect 21180 32428 21232 32434
rect 21180 32370 21232 32376
rect 20260 32292 20312 32298
rect 20260 32234 20312 32240
rect 20076 32224 20128 32230
rect 20076 32166 20128 32172
rect 19984 31884 20036 31890
rect 19984 31826 20036 31832
rect 19892 31476 19944 31482
rect 19892 31418 19944 31424
rect 19340 31272 19392 31278
rect 19340 31214 19392 31220
rect 19800 31272 19852 31278
rect 19800 31214 19852 31220
rect 19892 31272 19944 31278
rect 19892 31214 19944 31220
rect 19352 30376 19380 31214
rect 19580 31036 19876 31056
rect 19636 31034 19660 31036
rect 19716 31034 19740 31036
rect 19796 31034 19820 31036
rect 19658 30982 19660 31034
rect 19722 30982 19734 31034
rect 19796 30982 19798 31034
rect 19636 30980 19660 30982
rect 19716 30980 19740 30982
rect 19796 30980 19820 30982
rect 19580 30960 19876 30980
rect 19524 30388 19576 30394
rect 19352 30348 19524 30376
rect 19524 30330 19576 30336
rect 19536 30190 19564 30330
rect 19904 30190 19932 31214
rect 19984 30660 20036 30666
rect 19984 30602 20036 30608
rect 19524 30184 19576 30190
rect 19800 30184 19852 30190
rect 19524 30126 19576 30132
rect 19798 30152 19800 30161
rect 19892 30184 19944 30190
rect 19852 30152 19854 30161
rect 19340 30116 19392 30122
rect 19892 30126 19944 30132
rect 19798 30087 19854 30096
rect 19340 30058 19392 30064
rect 19352 28744 19380 30058
rect 19580 29948 19876 29968
rect 19636 29946 19660 29948
rect 19716 29946 19740 29948
rect 19796 29946 19820 29948
rect 19658 29894 19660 29946
rect 19722 29894 19734 29946
rect 19796 29894 19798 29946
rect 19636 29892 19660 29894
rect 19716 29892 19740 29894
rect 19796 29892 19820 29894
rect 19580 29872 19876 29892
rect 19800 29708 19852 29714
rect 19904 29696 19932 30126
rect 19996 29782 20024 30602
rect 19984 29776 20036 29782
rect 19984 29718 20036 29724
rect 19852 29668 19932 29696
rect 19800 29650 19852 29656
rect 19616 29640 19668 29646
rect 19614 29608 19616 29617
rect 19668 29608 19670 29617
rect 19614 29543 19670 29552
rect 19812 29345 19840 29650
rect 19982 29608 20038 29617
rect 19982 29543 20038 29552
rect 19798 29336 19854 29345
rect 19798 29271 19854 29280
rect 19432 29096 19484 29102
rect 19432 29038 19484 29044
rect 19444 28937 19472 29038
rect 19430 28928 19486 28937
rect 19430 28863 19486 28872
rect 19580 28860 19876 28880
rect 19636 28858 19660 28860
rect 19716 28858 19740 28860
rect 19796 28858 19820 28860
rect 19658 28806 19660 28858
rect 19722 28806 19734 28858
rect 19796 28806 19798 28858
rect 19636 28804 19660 28806
rect 19716 28804 19740 28806
rect 19796 28804 19820 28806
rect 19580 28784 19876 28804
rect 19352 28716 19748 28744
rect 19340 28620 19392 28626
rect 19340 28562 19392 28568
rect 19432 28620 19484 28626
rect 19432 28562 19484 28568
rect 19352 28529 19380 28562
rect 19338 28520 19394 28529
rect 19338 28455 19394 28464
rect 19444 28404 19472 28562
rect 19616 28416 19668 28422
rect 19444 28376 19616 28404
rect 19616 28358 19668 28364
rect 19432 28076 19484 28082
rect 19432 28018 19484 28024
rect 19340 28008 19392 28014
rect 19340 27950 19392 27956
rect 19352 22098 19380 27950
rect 19444 27538 19472 28018
rect 19628 28014 19656 28358
rect 19720 28150 19748 28716
rect 19708 28144 19760 28150
rect 19708 28086 19760 28092
rect 19616 28008 19668 28014
rect 19616 27950 19668 27956
rect 19580 27772 19876 27792
rect 19636 27770 19660 27772
rect 19716 27770 19740 27772
rect 19796 27770 19820 27772
rect 19658 27718 19660 27770
rect 19722 27718 19734 27770
rect 19796 27718 19798 27770
rect 19636 27716 19660 27718
rect 19716 27716 19740 27718
rect 19796 27716 19820 27718
rect 19580 27696 19876 27716
rect 19996 27538 20024 29543
rect 19432 27532 19484 27538
rect 19432 27474 19484 27480
rect 19892 27532 19944 27538
rect 19892 27474 19944 27480
rect 19984 27532 20036 27538
rect 19984 27474 20036 27480
rect 19580 26684 19876 26704
rect 19636 26682 19660 26684
rect 19716 26682 19740 26684
rect 19796 26682 19820 26684
rect 19658 26630 19660 26682
rect 19722 26630 19734 26682
rect 19796 26630 19798 26682
rect 19636 26628 19660 26630
rect 19716 26628 19740 26630
rect 19796 26628 19820 26630
rect 19580 26608 19876 26628
rect 19580 25596 19876 25616
rect 19636 25594 19660 25596
rect 19716 25594 19740 25596
rect 19796 25594 19820 25596
rect 19658 25542 19660 25594
rect 19722 25542 19734 25594
rect 19796 25542 19798 25594
rect 19636 25540 19660 25542
rect 19716 25540 19740 25542
rect 19796 25540 19820 25542
rect 19580 25520 19876 25540
rect 19580 24508 19876 24528
rect 19636 24506 19660 24508
rect 19716 24506 19740 24508
rect 19796 24506 19820 24508
rect 19658 24454 19660 24506
rect 19722 24454 19734 24506
rect 19796 24454 19798 24506
rect 19636 24452 19660 24454
rect 19716 24452 19740 24454
rect 19796 24452 19820 24454
rect 19580 24432 19876 24452
rect 19524 24268 19576 24274
rect 19524 24210 19576 24216
rect 19536 23866 19564 24210
rect 19524 23860 19576 23866
rect 19524 23802 19576 23808
rect 19580 23420 19876 23440
rect 19636 23418 19660 23420
rect 19716 23418 19740 23420
rect 19796 23418 19820 23420
rect 19658 23366 19660 23418
rect 19722 23366 19734 23418
rect 19796 23366 19798 23418
rect 19636 23364 19660 23366
rect 19716 23364 19740 23366
rect 19796 23364 19820 23366
rect 19430 23352 19486 23361
rect 19580 23344 19876 23364
rect 19430 23287 19432 23296
rect 19484 23287 19486 23296
rect 19432 23258 19484 23264
rect 19904 22710 19932 27474
rect 20088 25906 20116 32166
rect 20168 31204 20220 31210
rect 20168 31146 20220 31152
rect 20180 29578 20208 31146
rect 20272 30938 20300 32234
rect 20350 31920 20406 31929
rect 20350 31855 20352 31864
rect 20404 31855 20406 31864
rect 20996 31884 21048 31890
rect 20352 31826 20404 31832
rect 21272 31884 21324 31890
rect 21048 31844 21128 31872
rect 20996 31826 21048 31832
rect 20352 31680 20404 31686
rect 20352 31622 20404 31628
rect 20364 31278 20392 31622
rect 20628 31476 20680 31482
rect 20628 31418 20680 31424
rect 20352 31272 20404 31278
rect 20352 31214 20404 31220
rect 20260 30932 20312 30938
rect 20260 30874 20312 30880
rect 20352 30728 20404 30734
rect 20352 30670 20404 30676
rect 20260 30388 20312 30394
rect 20260 30330 20312 30336
rect 20168 29572 20220 29578
rect 20168 29514 20220 29520
rect 20166 29336 20222 29345
rect 20166 29271 20222 29280
rect 20180 28558 20208 29271
rect 20272 28966 20300 30330
rect 20260 28960 20312 28966
rect 20260 28902 20312 28908
rect 20260 28756 20312 28762
rect 20260 28698 20312 28704
rect 20168 28552 20220 28558
rect 20168 28494 20220 28500
rect 20076 25900 20128 25906
rect 20076 25842 20128 25848
rect 19984 25832 20036 25838
rect 19984 25774 20036 25780
rect 19996 23254 20024 25774
rect 20168 24744 20220 24750
rect 20168 24686 20220 24692
rect 20180 24206 20208 24686
rect 20272 24274 20300 28698
rect 20364 27554 20392 30670
rect 20536 30184 20588 30190
rect 20536 30126 20588 30132
rect 20548 29782 20576 30126
rect 20536 29776 20588 29782
rect 20536 29718 20588 29724
rect 20536 29096 20588 29102
rect 20536 29038 20588 29044
rect 20364 27526 20484 27554
rect 20352 27464 20404 27470
rect 20352 27406 20404 27412
rect 20364 26926 20392 27406
rect 20352 26920 20404 26926
rect 20352 26862 20404 26868
rect 20352 24880 20404 24886
rect 20352 24822 20404 24828
rect 20364 24410 20392 24822
rect 20352 24404 20404 24410
rect 20352 24346 20404 24352
rect 20260 24268 20312 24274
rect 20260 24210 20312 24216
rect 20168 24200 20220 24206
rect 20168 24142 20220 24148
rect 20168 23792 20220 23798
rect 20168 23734 20220 23740
rect 19984 23248 20036 23254
rect 19984 23190 20036 23196
rect 19892 22704 19944 22710
rect 19892 22646 19944 22652
rect 20076 22500 20128 22506
rect 20076 22442 20128 22448
rect 19580 22332 19876 22352
rect 19636 22330 19660 22332
rect 19716 22330 19740 22332
rect 19796 22330 19820 22332
rect 19658 22278 19660 22330
rect 19722 22278 19734 22330
rect 19796 22278 19798 22330
rect 19636 22276 19660 22278
rect 19716 22276 19740 22278
rect 19796 22276 19820 22278
rect 19580 22256 19876 22276
rect 19340 22092 19392 22098
rect 19340 22034 19392 22040
rect 19892 22092 19944 22098
rect 19892 22034 19944 22040
rect 19340 21888 19392 21894
rect 19340 21830 19392 21836
rect 19352 19802 19380 21830
rect 19580 21244 19876 21264
rect 19636 21242 19660 21244
rect 19716 21242 19740 21244
rect 19796 21242 19820 21244
rect 19658 21190 19660 21242
rect 19722 21190 19734 21242
rect 19796 21190 19798 21242
rect 19636 21188 19660 21190
rect 19716 21188 19740 21190
rect 19796 21188 19820 21190
rect 19580 21168 19876 21188
rect 19432 21072 19484 21078
rect 19432 21014 19484 21020
rect 19444 20466 19472 21014
rect 19904 21010 19932 22034
rect 19984 21072 20036 21078
rect 19984 21014 20036 21020
rect 19892 21004 19944 21010
rect 19892 20946 19944 20952
rect 19432 20460 19484 20466
rect 19432 20402 19484 20408
rect 19432 20324 19484 20330
rect 19432 20266 19484 20272
rect 19444 19961 19472 20266
rect 19580 20156 19876 20176
rect 19636 20154 19660 20156
rect 19716 20154 19740 20156
rect 19796 20154 19820 20156
rect 19658 20102 19660 20154
rect 19722 20102 19734 20154
rect 19796 20102 19798 20154
rect 19636 20100 19660 20102
rect 19716 20100 19740 20102
rect 19796 20100 19820 20102
rect 19580 20080 19876 20100
rect 19708 19984 19760 19990
rect 19430 19952 19486 19961
rect 19430 19887 19486 19896
rect 19706 19952 19708 19961
rect 19760 19952 19762 19961
rect 19706 19887 19762 19896
rect 19800 19848 19852 19854
rect 19352 19774 19564 19802
rect 19800 19790 19852 19796
rect 19340 19712 19392 19718
rect 19340 19654 19392 19660
rect 19352 19378 19380 19654
rect 19340 19372 19392 19378
rect 19340 19314 19392 19320
rect 19536 19156 19564 19774
rect 19708 19712 19760 19718
rect 19708 19654 19760 19660
rect 19616 19440 19668 19446
rect 19616 19382 19668 19388
rect 19628 19310 19656 19382
rect 19720 19310 19748 19654
rect 19616 19304 19668 19310
rect 19616 19246 19668 19252
rect 19708 19304 19760 19310
rect 19708 19246 19760 19252
rect 19352 19128 19564 19156
rect 19812 19156 19840 19790
rect 19904 19292 19932 20946
rect 19996 20058 20024 21014
rect 19984 20052 20036 20058
rect 19984 19994 20036 20000
rect 19996 19553 20024 19994
rect 19982 19544 20038 19553
rect 19982 19479 20038 19488
rect 19984 19304 20036 19310
rect 19904 19264 19984 19292
rect 19984 19246 20036 19252
rect 19812 19128 19932 19156
rect 19352 17814 19380 19128
rect 19580 19068 19876 19088
rect 19636 19066 19660 19068
rect 19716 19066 19740 19068
rect 19796 19066 19820 19068
rect 19658 19014 19660 19066
rect 19722 19014 19734 19066
rect 19796 19014 19798 19066
rect 19636 19012 19660 19014
rect 19716 19012 19740 19014
rect 19796 19012 19820 19014
rect 19580 18992 19876 19012
rect 19524 18896 19576 18902
rect 19522 18864 19524 18873
rect 19616 18896 19668 18902
rect 19576 18864 19578 18873
rect 19616 18838 19668 18844
rect 19522 18799 19578 18808
rect 19628 18737 19656 18838
rect 19614 18728 19670 18737
rect 19614 18663 19670 18672
rect 19616 18284 19668 18290
rect 19616 18226 19668 18232
rect 19708 18284 19760 18290
rect 19708 18226 19760 18232
rect 19628 18170 19656 18226
rect 19720 18193 19748 18226
rect 19444 18142 19656 18170
rect 19706 18184 19762 18193
rect 19340 17808 19392 17814
rect 19340 17750 19392 17756
rect 19444 17270 19472 18142
rect 19706 18119 19762 18128
rect 19580 17980 19876 18000
rect 19636 17978 19660 17980
rect 19716 17978 19740 17980
rect 19796 17978 19820 17980
rect 19658 17926 19660 17978
rect 19722 17926 19734 17978
rect 19796 17926 19798 17978
rect 19636 17924 19660 17926
rect 19716 17924 19740 17926
rect 19796 17924 19820 17926
rect 19580 17904 19876 17924
rect 19708 17740 19760 17746
rect 19708 17682 19760 17688
rect 19720 17270 19748 17682
rect 19432 17264 19484 17270
rect 19432 17206 19484 17212
rect 19708 17264 19760 17270
rect 19708 17206 19760 17212
rect 19340 17128 19392 17134
rect 19340 17070 19392 17076
rect 19352 16454 19380 17070
rect 19580 16892 19876 16912
rect 19636 16890 19660 16892
rect 19716 16890 19740 16892
rect 19796 16890 19820 16892
rect 19658 16838 19660 16890
rect 19722 16838 19734 16890
rect 19796 16838 19798 16890
rect 19636 16836 19660 16838
rect 19716 16836 19740 16838
rect 19796 16836 19820 16838
rect 19580 16816 19876 16836
rect 19340 16448 19392 16454
rect 19340 16390 19392 16396
rect 19432 16448 19484 16454
rect 19432 16390 19484 16396
rect 19352 16046 19380 16390
rect 19340 16040 19392 16046
rect 19340 15982 19392 15988
rect 19352 14958 19380 15982
rect 19444 15978 19472 16390
rect 19432 15972 19484 15978
rect 19432 15914 19484 15920
rect 19580 15804 19876 15824
rect 19636 15802 19660 15804
rect 19716 15802 19740 15804
rect 19796 15802 19820 15804
rect 19658 15750 19660 15802
rect 19722 15750 19734 15802
rect 19796 15750 19798 15802
rect 19636 15748 19660 15750
rect 19716 15748 19740 15750
rect 19796 15748 19820 15750
rect 19580 15728 19876 15748
rect 19904 15162 19932 19128
rect 20088 18970 20116 22442
rect 20180 21894 20208 23734
rect 20260 22568 20312 22574
rect 20260 22510 20312 22516
rect 20168 21888 20220 21894
rect 20168 21830 20220 21836
rect 20168 21004 20220 21010
rect 20168 20946 20220 20952
rect 20180 19718 20208 20946
rect 20168 19712 20220 19718
rect 20168 19654 20220 19660
rect 20166 19544 20222 19553
rect 20166 19479 20222 19488
rect 20076 18964 20128 18970
rect 20076 18906 20128 18912
rect 20180 18902 20208 19479
rect 20168 18896 20220 18902
rect 20168 18838 20220 18844
rect 20272 18170 20300 22510
rect 20364 21622 20392 24346
rect 20456 23236 20484 27526
rect 20548 26994 20576 29038
rect 20640 28218 20668 31418
rect 21100 31278 21128 31844
rect 21272 31826 21324 31832
rect 21088 31272 21140 31278
rect 21088 31214 21140 31220
rect 21100 30190 21128 31214
rect 21088 30184 21140 30190
rect 20718 30152 20774 30161
rect 21088 30126 21140 30132
rect 20718 30087 20774 30096
rect 20732 29714 20760 30087
rect 21180 29776 21232 29782
rect 21180 29718 21232 29724
rect 20720 29708 20772 29714
rect 20720 29650 20772 29656
rect 20904 29708 20956 29714
rect 20904 29650 20956 29656
rect 21088 29708 21140 29714
rect 21088 29650 21140 29656
rect 20720 28484 20772 28490
rect 20720 28426 20772 28432
rect 20628 28212 20680 28218
rect 20628 28154 20680 28160
rect 20732 27538 20760 28426
rect 20812 28008 20864 28014
rect 20812 27950 20864 27956
rect 20720 27532 20772 27538
rect 20720 27474 20772 27480
rect 20824 27402 20852 27950
rect 20812 27396 20864 27402
rect 20812 27338 20864 27344
rect 20536 26988 20588 26994
rect 20536 26930 20588 26936
rect 20812 26444 20864 26450
rect 20812 26386 20864 26392
rect 20720 25832 20772 25838
rect 20720 25774 20772 25780
rect 20732 25430 20760 25774
rect 20720 25424 20772 25430
rect 20720 25366 20772 25372
rect 20824 25294 20852 26386
rect 20916 25362 20944 29650
rect 20996 29640 21048 29646
rect 20996 29582 21048 29588
rect 21008 29306 21036 29582
rect 20996 29300 21048 29306
rect 20996 29242 21048 29248
rect 20996 28552 21048 28558
rect 20996 28494 21048 28500
rect 21008 27418 21036 28494
rect 21100 27538 21128 29650
rect 21088 27532 21140 27538
rect 21088 27474 21140 27480
rect 21008 27390 21128 27418
rect 21100 26246 21128 27390
rect 21088 26240 21140 26246
rect 21088 26182 21140 26188
rect 21100 25362 21128 26182
rect 20904 25356 20956 25362
rect 20904 25298 20956 25304
rect 21088 25356 21140 25362
rect 21088 25298 21140 25304
rect 20812 25288 20864 25294
rect 20812 25230 20864 25236
rect 20536 24812 20588 24818
rect 20536 24754 20588 24760
rect 20548 23662 20576 24754
rect 20916 24426 20944 25298
rect 20824 24410 20944 24426
rect 20824 24404 20956 24410
rect 20824 24398 20904 24404
rect 20824 23662 20852 24398
rect 20904 24346 20956 24352
rect 20904 24268 20956 24274
rect 20904 24210 20956 24216
rect 20916 23662 20944 24210
rect 21192 23866 21220 29718
rect 21180 23860 21232 23866
rect 21180 23802 21232 23808
rect 21284 23746 21312 31826
rect 21560 29714 21588 33458
rect 21824 33448 21876 33454
rect 21824 33390 21876 33396
rect 21836 32842 21864 33390
rect 21824 32836 21876 32842
rect 21824 32778 21876 32784
rect 21732 32768 21784 32774
rect 21732 32710 21784 32716
rect 21744 32570 21772 32710
rect 21732 32564 21784 32570
rect 21732 32506 21784 32512
rect 21824 32360 21876 32366
rect 21824 32302 21876 32308
rect 21836 31754 21864 32302
rect 21824 31748 21876 31754
rect 21824 31690 21876 31696
rect 21640 31340 21692 31346
rect 21640 31282 21692 31288
rect 21732 31340 21784 31346
rect 21732 31282 21784 31288
rect 21652 30802 21680 31282
rect 21744 30938 21772 31282
rect 21732 30932 21784 30938
rect 21732 30874 21784 30880
rect 21640 30796 21692 30802
rect 21640 30738 21692 30744
rect 21640 30184 21692 30190
rect 21640 30126 21692 30132
rect 21548 29708 21600 29714
rect 21548 29650 21600 29656
rect 21364 29096 21416 29102
rect 21364 29038 21416 29044
rect 21376 28626 21404 29038
rect 21456 28756 21508 28762
rect 21456 28698 21508 28704
rect 21364 28620 21416 28626
rect 21364 28562 21416 28568
rect 21376 28014 21404 28562
rect 21364 28008 21416 28014
rect 21364 27950 21416 27956
rect 21376 27334 21404 27950
rect 21364 27328 21416 27334
rect 21364 27270 21416 27276
rect 21008 23718 21312 23746
rect 20536 23656 20588 23662
rect 20536 23598 20588 23604
rect 20812 23656 20864 23662
rect 20812 23598 20864 23604
rect 20904 23656 20956 23662
rect 20904 23598 20956 23604
rect 20456 23208 20852 23236
rect 20720 23112 20772 23118
rect 20720 23054 20772 23060
rect 20628 22568 20680 22574
rect 20628 22510 20680 22516
rect 20536 21888 20588 21894
rect 20536 21830 20588 21836
rect 20352 21616 20404 21622
rect 20352 21558 20404 21564
rect 20364 21162 20392 21558
rect 20364 21134 20484 21162
rect 20352 19916 20404 19922
rect 20352 19858 20404 19864
rect 20364 19786 20392 19858
rect 20352 19780 20404 19786
rect 20352 19722 20404 19728
rect 20364 19310 20392 19722
rect 20456 19446 20484 21134
rect 20444 19440 20496 19446
rect 20444 19382 20496 19388
rect 20352 19304 20404 19310
rect 20352 19246 20404 19252
rect 20364 18630 20392 19246
rect 20548 18873 20576 21830
rect 20534 18864 20590 18873
rect 20534 18799 20590 18808
rect 20548 18630 20576 18799
rect 20352 18624 20404 18630
rect 20352 18566 20404 18572
rect 20536 18624 20588 18630
rect 20536 18566 20588 18572
rect 20536 18216 20588 18222
rect 20272 18142 20484 18170
rect 20536 18158 20588 18164
rect 20352 18080 20404 18086
rect 20352 18022 20404 18028
rect 20168 17808 20220 17814
rect 20168 17750 20220 17756
rect 19984 17128 20036 17134
rect 19984 17070 20036 17076
rect 20076 17128 20128 17134
rect 20076 17070 20128 17076
rect 19996 16794 20024 17070
rect 19984 16788 20036 16794
rect 19984 16730 20036 16736
rect 19984 16108 20036 16114
rect 19984 16050 20036 16056
rect 19432 15156 19484 15162
rect 19432 15098 19484 15104
rect 19892 15156 19944 15162
rect 19892 15098 19944 15104
rect 19340 14952 19392 14958
rect 19340 14894 19392 14900
rect 19444 14600 19472 15098
rect 19580 14716 19876 14736
rect 19636 14714 19660 14716
rect 19716 14714 19740 14716
rect 19796 14714 19820 14716
rect 19658 14662 19660 14714
rect 19722 14662 19734 14714
rect 19796 14662 19798 14714
rect 19636 14660 19660 14662
rect 19716 14660 19740 14662
rect 19796 14660 19820 14662
rect 19580 14640 19876 14660
rect 19352 14572 19472 14600
rect 19352 13394 19380 14572
rect 19432 14476 19484 14482
rect 19432 14418 19484 14424
rect 19444 14278 19472 14418
rect 19432 14272 19484 14278
rect 19432 14214 19484 14220
rect 19340 13388 19392 13394
rect 19340 13330 19392 13336
rect 19248 12912 19300 12918
rect 19248 12854 19300 12860
rect 19156 12844 19208 12850
rect 19156 12786 19208 12792
rect 18880 12436 18932 12442
rect 18880 12378 18932 12384
rect 18788 11212 18840 11218
rect 18788 11154 18840 11160
rect 18696 10192 18748 10198
rect 18696 10134 18748 10140
rect 18604 9512 18656 9518
rect 18604 9454 18656 9460
rect 18616 9042 18644 9454
rect 18604 9036 18656 9042
rect 18604 8978 18656 8984
rect 18616 8430 18644 8978
rect 18708 8906 18736 10134
rect 18696 8900 18748 8906
rect 18696 8842 18748 8848
rect 18604 8424 18656 8430
rect 18604 8366 18656 8372
rect 18616 7954 18644 8366
rect 18604 7948 18656 7954
rect 18604 7890 18656 7896
rect 18420 7744 18472 7750
rect 18420 7686 18472 7692
rect 18432 7342 18460 7686
rect 18420 7336 18472 7342
rect 18420 7278 18472 7284
rect 18328 6860 18380 6866
rect 18328 6802 18380 6808
rect 18236 6792 18288 6798
rect 18236 6734 18288 6740
rect 18052 6248 18104 6254
rect 18052 6190 18104 6196
rect 17960 5908 18012 5914
rect 17960 5850 18012 5856
rect 18340 5846 18368 6802
rect 18512 6248 18564 6254
rect 18512 6190 18564 6196
rect 18328 5840 18380 5846
rect 18328 5782 18380 5788
rect 17868 5704 17920 5710
rect 17868 5646 17920 5652
rect 18524 5166 18552 6190
rect 18800 5370 18828 11154
rect 18892 8974 18920 12378
rect 19064 12300 19116 12306
rect 19064 12242 19116 12248
rect 19076 11354 19104 12242
rect 19168 11558 19196 12786
rect 19340 12640 19392 12646
rect 19340 12582 19392 12588
rect 19248 12232 19300 12238
rect 19248 12174 19300 12180
rect 19260 12102 19288 12174
rect 19248 12096 19300 12102
rect 19248 12038 19300 12044
rect 19352 11830 19380 12582
rect 19444 12306 19472 14214
rect 19996 13870 20024 16050
rect 19984 13864 20036 13870
rect 19984 13806 20036 13812
rect 19580 13628 19876 13648
rect 19636 13626 19660 13628
rect 19716 13626 19740 13628
rect 19796 13626 19820 13628
rect 19658 13574 19660 13626
rect 19722 13574 19734 13626
rect 19796 13574 19798 13626
rect 19636 13572 19660 13574
rect 19716 13572 19740 13574
rect 19796 13572 19820 13574
rect 19580 13552 19876 13572
rect 19892 13388 19944 13394
rect 19892 13330 19944 13336
rect 19580 12540 19876 12560
rect 19636 12538 19660 12540
rect 19716 12538 19740 12540
rect 19796 12538 19820 12540
rect 19658 12486 19660 12538
rect 19722 12486 19734 12538
rect 19796 12486 19798 12538
rect 19636 12484 19660 12486
rect 19716 12484 19740 12486
rect 19796 12484 19820 12486
rect 19580 12464 19876 12484
rect 19524 12368 19576 12374
rect 19524 12310 19576 12316
rect 19432 12300 19484 12306
rect 19432 12242 19484 12248
rect 19340 11824 19392 11830
rect 19340 11766 19392 11772
rect 19156 11552 19208 11558
rect 19536 11540 19564 12310
rect 19904 12238 19932 13330
rect 20088 12782 20116 17070
rect 20180 15162 20208 17750
rect 20364 16658 20392 18022
rect 20352 16652 20404 16658
rect 20352 16594 20404 16600
rect 20260 16040 20312 16046
rect 20260 15982 20312 15988
rect 20168 15156 20220 15162
rect 20168 15098 20220 15104
rect 20168 15020 20220 15026
rect 20168 14962 20220 14968
rect 20180 14278 20208 14962
rect 20168 14272 20220 14278
rect 20168 14214 20220 14220
rect 19984 12776 20036 12782
rect 19984 12718 20036 12724
rect 20076 12776 20128 12782
rect 20076 12718 20128 12724
rect 19892 12232 19944 12238
rect 19892 12174 19944 12180
rect 19616 11892 19668 11898
rect 19616 11834 19668 11840
rect 19628 11694 19656 11834
rect 19996 11762 20024 12718
rect 20272 12374 20300 15982
rect 20364 13394 20392 16594
rect 20456 13394 20484 18142
rect 20548 17678 20576 18158
rect 20536 17672 20588 17678
rect 20536 17614 20588 17620
rect 20536 16652 20588 16658
rect 20536 16594 20588 16600
rect 20548 15910 20576 16594
rect 20536 15904 20588 15910
rect 20536 15846 20588 15852
rect 20548 15570 20576 15846
rect 20536 15564 20588 15570
rect 20536 15506 20588 15512
rect 20536 15156 20588 15162
rect 20536 15098 20588 15104
rect 20352 13388 20404 13394
rect 20352 13330 20404 13336
rect 20444 13388 20496 13394
rect 20444 13330 20496 13336
rect 20548 12866 20576 15098
rect 20640 13530 20668 22510
rect 20732 19514 20760 23054
rect 20824 19854 20852 23208
rect 20916 23186 20944 23598
rect 20904 23180 20956 23186
rect 20904 23122 20956 23128
rect 20904 21412 20956 21418
rect 20904 21354 20956 21360
rect 20916 21010 20944 21354
rect 20904 21004 20956 21010
rect 20904 20946 20956 20952
rect 20812 19848 20864 19854
rect 20812 19790 20864 19796
rect 20812 19712 20864 19718
rect 20812 19654 20864 19660
rect 20720 19508 20772 19514
rect 20720 19450 20772 19456
rect 20720 17128 20772 17134
rect 20720 17070 20772 17076
rect 20732 16046 20760 17070
rect 20720 16040 20772 16046
rect 20720 15982 20772 15988
rect 20732 14958 20760 15982
rect 20720 14952 20772 14958
rect 20720 14894 20772 14900
rect 20628 13524 20680 13530
rect 20628 13466 20680 13472
rect 20628 13388 20680 13394
rect 20628 13330 20680 13336
rect 20456 12838 20576 12866
rect 20352 12776 20404 12782
rect 20352 12718 20404 12724
rect 20260 12368 20312 12374
rect 20260 12310 20312 12316
rect 20076 12300 20128 12306
rect 20076 12242 20128 12248
rect 19984 11756 20036 11762
rect 19984 11698 20036 11704
rect 19616 11688 19668 11694
rect 19616 11630 19668 11636
rect 19156 11494 19208 11500
rect 19444 11512 19564 11540
rect 19064 11348 19116 11354
rect 19064 11290 19116 11296
rect 19064 11212 19116 11218
rect 19064 11154 19116 11160
rect 18972 10600 19024 10606
rect 18972 10542 19024 10548
rect 18984 10198 19012 10542
rect 18972 10192 19024 10198
rect 18972 10134 19024 10140
rect 19076 10146 19104 11154
rect 19168 10538 19196 11494
rect 19156 10532 19208 10538
rect 19156 10474 19208 10480
rect 19340 10464 19392 10470
rect 19340 10406 19392 10412
rect 19076 10118 19196 10146
rect 18972 9512 19024 9518
rect 18972 9454 19024 9460
rect 18984 9024 19012 9454
rect 19064 9376 19116 9382
rect 19168 9364 19196 10118
rect 19116 9336 19196 9364
rect 19064 9318 19116 9324
rect 19064 9036 19116 9042
rect 18984 8996 19064 9024
rect 19064 8978 19116 8984
rect 18880 8968 18932 8974
rect 18880 8910 18932 8916
rect 19076 8430 19104 8978
rect 19168 8906 19196 9336
rect 19156 8900 19208 8906
rect 19156 8842 19208 8848
rect 19064 8424 19116 8430
rect 19062 8392 19064 8401
rect 19116 8392 19118 8401
rect 19062 8327 19118 8336
rect 19246 8392 19302 8401
rect 19352 8362 19380 10406
rect 19444 10248 19472 11512
rect 19580 11452 19876 11472
rect 19636 11450 19660 11452
rect 19716 11450 19740 11452
rect 19796 11450 19820 11452
rect 19658 11398 19660 11450
rect 19722 11398 19734 11450
rect 19796 11398 19798 11450
rect 19636 11396 19660 11398
rect 19716 11396 19740 11398
rect 19796 11396 19820 11398
rect 19580 11376 19876 11396
rect 19800 11212 19852 11218
rect 19800 11154 19852 11160
rect 19812 10849 19840 11154
rect 19996 11082 20024 11698
rect 20088 11354 20116 12242
rect 20168 12232 20220 12238
rect 20168 12174 20220 12180
rect 20076 11348 20128 11354
rect 20076 11290 20128 11296
rect 20088 11218 20116 11290
rect 20076 11212 20128 11218
rect 20076 11154 20128 11160
rect 20180 11098 20208 12174
rect 20260 12096 20312 12102
rect 20260 12038 20312 12044
rect 20272 11762 20300 12038
rect 20260 11756 20312 11762
rect 20260 11698 20312 11704
rect 20258 11656 20314 11665
rect 20258 11591 20314 11600
rect 19984 11076 20036 11082
rect 19984 11018 20036 11024
rect 20088 11070 20208 11098
rect 19798 10840 19854 10849
rect 19996 10826 20024 11018
rect 19798 10775 19854 10784
rect 19904 10798 20024 10826
rect 19580 10364 19876 10384
rect 19636 10362 19660 10364
rect 19716 10362 19740 10364
rect 19796 10362 19820 10364
rect 19658 10310 19660 10362
rect 19722 10310 19734 10362
rect 19796 10310 19798 10362
rect 19636 10308 19660 10310
rect 19716 10308 19740 10310
rect 19796 10308 19820 10310
rect 19580 10288 19876 10308
rect 19444 10220 19564 10248
rect 19432 10124 19484 10130
rect 19432 10066 19484 10072
rect 19444 9178 19472 10066
rect 19536 9722 19564 10220
rect 19904 10062 19932 10798
rect 19984 10124 20036 10130
rect 19984 10066 20036 10072
rect 19892 10056 19944 10062
rect 19892 9998 19944 10004
rect 19524 9716 19576 9722
rect 19524 9658 19576 9664
rect 19890 9480 19946 9489
rect 19890 9415 19946 9424
rect 19580 9276 19876 9296
rect 19636 9274 19660 9276
rect 19716 9274 19740 9276
rect 19796 9274 19820 9276
rect 19658 9222 19660 9274
rect 19722 9222 19734 9274
rect 19796 9222 19798 9274
rect 19636 9220 19660 9222
rect 19716 9220 19740 9222
rect 19796 9220 19820 9222
rect 19580 9200 19876 9220
rect 19432 9172 19484 9178
rect 19432 9114 19484 9120
rect 19904 9110 19932 9415
rect 19892 9104 19944 9110
rect 19892 9046 19944 9052
rect 19996 9024 20024 10066
rect 20088 10062 20116 11070
rect 20076 10056 20128 10062
rect 20076 9998 20128 10004
rect 20088 9926 20116 9998
rect 20076 9920 20128 9926
rect 20076 9862 20128 9868
rect 20168 9648 20220 9654
rect 20168 9590 20220 9596
rect 19996 8996 20116 9024
rect 19708 8968 19760 8974
rect 19536 8916 19708 8922
rect 19536 8910 19760 8916
rect 19536 8894 19748 8910
rect 19432 8492 19484 8498
rect 19536 8480 19564 8894
rect 19982 8664 20038 8673
rect 19982 8599 20038 8608
rect 19996 8498 20024 8599
rect 19484 8452 19564 8480
rect 19984 8492 20036 8498
rect 19432 8434 19484 8440
rect 19984 8434 20036 8440
rect 19246 8327 19302 8336
rect 19340 8356 19392 8362
rect 19260 7954 19288 8327
rect 19340 8298 19392 8304
rect 19580 8188 19876 8208
rect 19636 8186 19660 8188
rect 19716 8186 19740 8188
rect 19796 8186 19820 8188
rect 19658 8134 19660 8186
rect 19722 8134 19734 8186
rect 19796 8134 19798 8186
rect 19636 8132 19660 8134
rect 19716 8132 19740 8134
rect 19796 8132 19820 8134
rect 19580 8112 19876 8132
rect 19248 7948 19300 7954
rect 19248 7890 19300 7896
rect 19984 7744 20036 7750
rect 19984 7686 20036 7692
rect 19996 7546 20024 7686
rect 19984 7540 20036 7546
rect 19984 7482 20036 7488
rect 18972 7404 19024 7410
rect 18972 7346 19024 7352
rect 18984 6322 19012 7346
rect 19996 7342 20024 7482
rect 19340 7336 19392 7342
rect 19340 7278 19392 7284
rect 19984 7336 20036 7342
rect 19984 7278 20036 7284
rect 19246 6896 19302 6905
rect 19246 6831 19302 6840
rect 18972 6316 19024 6322
rect 18972 6258 19024 6264
rect 18880 5636 18932 5642
rect 18880 5578 18932 5584
rect 18788 5364 18840 5370
rect 18788 5306 18840 5312
rect 18892 5234 18920 5578
rect 19260 5574 19288 6831
rect 19352 6798 19380 7278
rect 19580 7100 19876 7120
rect 19636 7098 19660 7100
rect 19716 7098 19740 7100
rect 19796 7098 19820 7100
rect 19658 7046 19660 7098
rect 19722 7046 19734 7098
rect 19796 7046 19798 7098
rect 19636 7044 19660 7046
rect 19716 7044 19740 7046
rect 19796 7044 19820 7046
rect 19580 7024 19876 7044
rect 19996 6866 20024 7278
rect 19984 6860 20036 6866
rect 19984 6802 20036 6808
rect 20088 6798 20116 8996
rect 20180 8498 20208 9590
rect 20272 9382 20300 11591
rect 20260 9376 20312 9382
rect 20260 9318 20312 9324
rect 20260 9036 20312 9042
rect 20260 8978 20312 8984
rect 20272 8838 20300 8978
rect 20260 8832 20312 8838
rect 20260 8774 20312 8780
rect 20168 8492 20220 8498
rect 20168 8434 20220 8440
rect 19340 6792 19392 6798
rect 19340 6734 19392 6740
rect 20076 6792 20128 6798
rect 20076 6734 20128 6740
rect 20088 6458 20116 6734
rect 20076 6452 20128 6458
rect 20076 6394 20128 6400
rect 20364 6254 20392 12718
rect 20456 8906 20484 12838
rect 20536 12776 20588 12782
rect 20536 12718 20588 12724
rect 20640 12730 20668 13330
rect 20548 9042 20576 12718
rect 20640 12702 20760 12730
rect 20628 12640 20680 12646
rect 20628 12582 20680 12588
rect 20640 11898 20668 12582
rect 20628 11892 20680 11898
rect 20628 11834 20680 11840
rect 20628 11688 20680 11694
rect 20732 11665 20760 12702
rect 20824 11914 20852 19654
rect 20916 19310 20944 20946
rect 20904 19304 20956 19310
rect 20904 19246 20956 19252
rect 21008 16130 21036 23718
rect 21468 23322 21496 28698
rect 21546 28112 21602 28121
rect 21546 28047 21548 28056
rect 21600 28047 21602 28056
rect 21548 28018 21600 28024
rect 21652 27878 21680 30126
rect 21824 30116 21876 30122
rect 21824 30058 21876 30064
rect 21836 29782 21864 30058
rect 21824 29776 21876 29782
rect 21824 29718 21876 29724
rect 21822 29200 21878 29209
rect 21822 29135 21878 29144
rect 21836 29102 21864 29135
rect 21824 29096 21876 29102
rect 21744 29056 21824 29084
rect 21744 28218 21772 29056
rect 21928 29084 21956 33918
rect 22376 33856 22428 33862
rect 22376 33798 22428 33804
rect 22388 33454 22416 33798
rect 22664 33658 22692 34070
rect 22652 33652 22704 33658
rect 22652 33594 22704 33600
rect 22376 33448 22428 33454
rect 22376 33390 22428 33396
rect 22192 33040 22244 33046
rect 22192 32982 22244 32988
rect 22100 32972 22152 32978
rect 22100 32914 22152 32920
rect 22112 32366 22140 32914
rect 22100 32360 22152 32366
rect 22100 32302 22152 32308
rect 22204 32298 22232 32982
rect 22848 32978 22876 34478
rect 23032 34474 23060 35108
rect 23112 35090 23164 35096
rect 23204 35148 23256 35154
rect 23204 35090 23256 35096
rect 23400 35086 23428 35770
rect 23388 35080 23440 35086
rect 23388 35022 23440 35028
rect 23400 34678 23428 35022
rect 23584 35018 23612 36586
rect 23756 36168 23808 36174
rect 23808 36128 23888 36156
rect 23756 36110 23808 36116
rect 23756 35148 23808 35154
rect 23756 35090 23808 35096
rect 23572 35012 23624 35018
rect 23572 34954 23624 34960
rect 23388 34672 23440 34678
rect 23388 34614 23440 34620
rect 23480 34536 23532 34542
rect 23480 34478 23532 34484
rect 23664 34536 23716 34542
rect 23664 34478 23716 34484
rect 23020 34468 23072 34474
rect 23020 34410 23072 34416
rect 23492 34066 23520 34478
rect 23480 34060 23532 34066
rect 23532 34020 23612 34048
rect 23480 34002 23532 34008
rect 23584 33590 23612 34020
rect 23480 33584 23532 33590
rect 23480 33526 23532 33532
rect 23572 33584 23624 33590
rect 23572 33526 23624 33532
rect 23492 32978 23520 33526
rect 23572 33448 23624 33454
rect 23572 33390 23624 33396
rect 22836 32972 22888 32978
rect 22836 32914 22888 32920
rect 23480 32972 23532 32978
rect 23480 32914 23532 32920
rect 22468 32768 22520 32774
rect 22468 32710 22520 32716
rect 23480 32768 23532 32774
rect 23480 32710 23532 32716
rect 22192 32292 22244 32298
rect 22192 32234 22244 32240
rect 22008 31816 22060 31822
rect 22008 31758 22060 31764
rect 22020 31142 22048 31758
rect 22008 31136 22060 31142
rect 22008 31078 22060 31084
rect 22100 30660 22152 30666
rect 22100 30602 22152 30608
rect 22112 30190 22140 30602
rect 22100 30184 22152 30190
rect 22100 30126 22152 30132
rect 22008 29096 22060 29102
rect 21928 29056 22008 29084
rect 21824 29038 21876 29044
rect 22008 29038 22060 29044
rect 22100 28620 22152 28626
rect 22100 28562 22152 28568
rect 21824 28552 21876 28558
rect 21824 28494 21876 28500
rect 21732 28212 21784 28218
rect 21732 28154 21784 28160
rect 21732 27940 21784 27946
rect 21732 27882 21784 27888
rect 21640 27872 21692 27878
rect 21640 27814 21692 27820
rect 21548 27532 21600 27538
rect 21548 27474 21600 27480
rect 21456 23316 21508 23322
rect 21456 23258 21508 23264
rect 21364 22976 21416 22982
rect 21364 22918 21416 22924
rect 21376 22574 21404 22918
rect 21364 22568 21416 22574
rect 21364 22510 21416 22516
rect 21376 22030 21404 22510
rect 21180 22024 21232 22030
rect 21180 21966 21232 21972
rect 21364 22024 21416 22030
rect 21364 21966 21416 21972
rect 21088 19440 21140 19446
rect 21088 19382 21140 19388
rect 20916 16102 21036 16130
rect 20916 12918 20944 16102
rect 20996 16040 21048 16046
rect 20996 15982 21048 15988
rect 21008 15910 21036 15982
rect 20996 15904 21048 15910
rect 20996 15846 21048 15852
rect 21008 14958 21036 15846
rect 21100 15042 21128 19382
rect 21192 18970 21220 21966
rect 21456 21616 21508 21622
rect 21456 21558 21508 21564
rect 21468 21486 21496 21558
rect 21456 21480 21508 21486
rect 21456 21422 21508 21428
rect 21272 21004 21324 21010
rect 21272 20946 21324 20952
rect 21284 19310 21312 20946
rect 21272 19304 21324 19310
rect 21272 19246 21324 19252
rect 21180 18964 21232 18970
rect 21180 18906 21232 18912
rect 21284 18834 21312 19246
rect 21456 18964 21508 18970
rect 21456 18906 21508 18912
rect 21364 18896 21416 18902
rect 21364 18838 21416 18844
rect 21272 18828 21324 18834
rect 21272 18770 21324 18776
rect 21180 18624 21232 18630
rect 21180 18566 21232 18572
rect 21192 18086 21220 18566
rect 21376 18222 21404 18838
rect 21468 18358 21496 18906
rect 21456 18352 21508 18358
rect 21456 18294 21508 18300
rect 21364 18216 21416 18222
rect 21364 18158 21416 18164
rect 21180 18080 21232 18086
rect 21560 18068 21588 27474
rect 21744 27402 21772 27882
rect 21836 27606 21864 28494
rect 21916 28008 21968 28014
rect 21916 27950 21968 27956
rect 21824 27600 21876 27606
rect 21824 27542 21876 27548
rect 21732 27396 21784 27402
rect 21732 27338 21784 27344
rect 21640 26444 21692 26450
rect 21640 26386 21692 26392
rect 21652 23118 21680 26386
rect 21824 25356 21876 25362
rect 21824 25298 21876 25304
rect 21836 24818 21864 25298
rect 21928 24886 21956 27950
rect 22112 26994 22140 28562
rect 22204 27062 22232 32234
rect 22284 32224 22336 32230
rect 22284 32166 22336 32172
rect 22296 30734 22324 32166
rect 22480 31890 22508 32710
rect 23492 32570 23520 32710
rect 23584 32570 23612 33390
rect 23480 32564 23532 32570
rect 23480 32506 23532 32512
rect 23572 32564 23624 32570
rect 23572 32506 23624 32512
rect 23572 32360 23624 32366
rect 23676 32314 23704 34478
rect 23768 33998 23796 35090
rect 23860 34202 23888 36128
rect 23848 34196 23900 34202
rect 23848 34138 23900 34144
rect 23756 33992 23808 33998
rect 23756 33934 23808 33940
rect 23756 33448 23808 33454
rect 23860 33436 23888 34138
rect 23808 33408 23888 33436
rect 23940 33448 23992 33454
rect 23756 33390 23808 33396
rect 23940 33390 23992 33396
rect 23848 32360 23900 32366
rect 23624 32308 23796 32314
rect 23572 32302 23796 32308
rect 23848 32302 23900 32308
rect 23584 32298 23796 32302
rect 23584 32292 23808 32298
rect 23584 32286 23756 32292
rect 23756 32234 23808 32240
rect 22560 32224 22612 32230
rect 23860 32178 23888 32302
rect 22560 32166 22612 32172
rect 22468 31884 22520 31890
rect 22468 31826 22520 31832
rect 22376 31408 22428 31414
rect 22376 31350 22428 31356
rect 22388 30802 22416 31350
rect 22468 31136 22520 31142
rect 22468 31078 22520 31084
rect 22376 30796 22428 30802
rect 22376 30738 22428 30744
rect 22284 30728 22336 30734
rect 22284 30670 22336 30676
rect 22480 28762 22508 31078
rect 22572 29714 22600 32166
rect 23492 32150 23888 32178
rect 23296 31816 23348 31822
rect 23294 31784 23296 31793
rect 23348 31784 23350 31793
rect 23294 31719 23350 31728
rect 23308 31346 23336 31719
rect 23296 31340 23348 31346
rect 23296 31282 23348 31288
rect 23112 31204 23164 31210
rect 23112 31146 23164 31152
rect 22560 29708 22612 29714
rect 22560 29650 22612 29656
rect 22928 29708 22980 29714
rect 22928 29650 22980 29656
rect 22940 29617 22968 29650
rect 22926 29608 22982 29617
rect 22926 29543 22982 29552
rect 22836 29096 22888 29102
rect 22888 29056 23060 29084
rect 22836 29038 22888 29044
rect 22836 28960 22888 28966
rect 22836 28902 22888 28908
rect 22468 28756 22520 28762
rect 22468 28698 22520 28704
rect 22848 28626 22876 28902
rect 22836 28620 22888 28626
rect 22836 28562 22888 28568
rect 22848 28422 22876 28562
rect 22928 28552 22980 28558
rect 22928 28494 22980 28500
rect 22376 28416 22428 28422
rect 22376 28358 22428 28364
rect 22836 28416 22888 28422
rect 22836 28358 22888 28364
rect 22284 28212 22336 28218
rect 22284 28154 22336 28160
rect 22296 28014 22324 28154
rect 22284 28008 22336 28014
rect 22284 27950 22336 27956
rect 22284 27532 22336 27538
rect 22284 27474 22336 27480
rect 22192 27056 22244 27062
rect 22192 26998 22244 27004
rect 22100 26988 22152 26994
rect 22100 26930 22152 26936
rect 22112 26586 22140 26930
rect 22192 26920 22244 26926
rect 22296 26874 22324 27474
rect 22244 26868 22324 26874
rect 22192 26862 22324 26868
rect 22204 26846 22324 26862
rect 22100 26580 22152 26586
rect 22100 26522 22152 26528
rect 22204 26518 22232 26846
rect 22192 26512 22244 26518
rect 22192 26454 22244 26460
rect 22388 26450 22416 28358
rect 22744 27872 22796 27878
rect 22744 27814 22796 27820
rect 22468 27328 22520 27334
rect 22468 27270 22520 27276
rect 22376 26444 22428 26450
rect 22376 26386 22428 26392
rect 22008 25832 22060 25838
rect 22008 25774 22060 25780
rect 22284 25832 22336 25838
rect 22388 25820 22416 26386
rect 22336 25792 22416 25820
rect 22284 25774 22336 25780
rect 22020 25430 22048 25774
rect 22008 25424 22060 25430
rect 22008 25366 22060 25372
rect 22008 25288 22060 25294
rect 22008 25230 22060 25236
rect 21916 24880 21968 24886
rect 21916 24822 21968 24828
rect 21824 24812 21876 24818
rect 21824 24754 21876 24760
rect 21732 24744 21784 24750
rect 21732 24686 21784 24692
rect 21744 24274 21772 24686
rect 21732 24268 21784 24274
rect 21732 24210 21784 24216
rect 21744 23662 21772 24210
rect 21732 23656 21784 23662
rect 21732 23598 21784 23604
rect 21732 23316 21784 23322
rect 21732 23258 21784 23264
rect 21640 23112 21692 23118
rect 21640 23054 21692 23060
rect 21640 22568 21692 22574
rect 21640 22510 21692 22516
rect 21652 21146 21680 22510
rect 21640 21140 21692 21146
rect 21640 21082 21692 21088
rect 21640 20324 21692 20330
rect 21640 20266 21692 20272
rect 21652 19417 21680 20266
rect 21744 19446 21772 23258
rect 21836 23186 21864 24754
rect 22020 24596 22048 25230
rect 22192 25152 22244 25158
rect 22192 25094 22244 25100
rect 22020 24568 22140 24596
rect 22112 24410 22140 24568
rect 22100 24404 22152 24410
rect 22100 24346 22152 24352
rect 22204 24342 22232 25094
rect 22192 24336 22244 24342
rect 22192 24278 22244 24284
rect 22296 24138 22324 25774
rect 22480 25752 22508 27270
rect 22756 26926 22784 27814
rect 22744 26920 22796 26926
rect 22744 26862 22796 26868
rect 22560 26784 22612 26790
rect 22560 26726 22612 26732
rect 22572 26042 22600 26726
rect 22560 26036 22612 26042
rect 22560 25978 22612 25984
rect 22652 25832 22704 25838
rect 22652 25774 22704 25780
rect 22388 25724 22508 25752
rect 22560 25764 22612 25770
rect 22284 24132 22336 24138
rect 22284 24074 22336 24080
rect 22100 23724 22152 23730
rect 22100 23666 22152 23672
rect 21824 23180 21876 23186
rect 21824 23122 21876 23128
rect 21916 21412 21968 21418
rect 21916 21354 21968 21360
rect 21824 20936 21876 20942
rect 21824 20878 21876 20884
rect 21732 19440 21784 19446
rect 21638 19408 21694 19417
rect 21732 19382 21784 19388
rect 21638 19343 21694 19352
rect 21836 19310 21864 20878
rect 21928 19938 21956 21354
rect 22112 20806 22140 23666
rect 22284 23588 22336 23594
rect 22284 23530 22336 23536
rect 22296 23186 22324 23530
rect 22284 23180 22336 23186
rect 22284 23122 22336 23128
rect 22296 22778 22324 23122
rect 22284 22772 22336 22778
rect 22284 22714 22336 22720
rect 22388 20942 22416 25724
rect 22560 25706 22612 25712
rect 22572 25226 22600 25706
rect 22560 25220 22612 25226
rect 22560 25162 22612 25168
rect 22664 24834 22692 25774
rect 22756 24954 22784 26862
rect 22940 26450 22968 28494
rect 23032 26790 23060 29056
rect 23020 26784 23072 26790
rect 23020 26726 23072 26732
rect 23124 26738 23152 31146
rect 23204 29708 23256 29714
rect 23204 29650 23256 29656
rect 23216 29306 23244 29650
rect 23296 29572 23348 29578
rect 23296 29514 23348 29520
rect 23308 29345 23336 29514
rect 23294 29336 23350 29345
rect 23204 29300 23256 29306
rect 23294 29271 23350 29280
rect 23204 29242 23256 29248
rect 23492 28626 23520 32150
rect 23952 32026 23980 33390
rect 23940 32020 23992 32026
rect 23940 31962 23992 31968
rect 23664 31884 23716 31890
rect 23664 31826 23716 31832
rect 23572 31816 23624 31822
rect 23572 31758 23624 31764
rect 23584 31278 23612 31758
rect 23572 31272 23624 31278
rect 23572 31214 23624 31220
rect 23572 31136 23624 31142
rect 23572 31078 23624 31084
rect 23584 30802 23612 31078
rect 23572 30796 23624 30802
rect 23572 30738 23624 30744
rect 23480 28620 23532 28626
rect 23480 28562 23532 28568
rect 23572 27600 23624 27606
rect 23572 27542 23624 27548
rect 23584 27130 23612 27542
rect 23572 27124 23624 27130
rect 23572 27066 23624 27072
rect 23572 26920 23624 26926
rect 23572 26862 23624 26868
rect 22928 26444 22980 26450
rect 22928 26386 22980 26392
rect 22744 24948 22796 24954
rect 22744 24890 22796 24896
rect 22836 24880 22888 24886
rect 22664 24806 22784 24834
rect 22836 24822 22888 24828
rect 22652 24744 22704 24750
rect 22652 24686 22704 24692
rect 22664 24274 22692 24686
rect 22652 24268 22704 24274
rect 22572 24228 22652 24256
rect 22468 24064 22520 24070
rect 22468 24006 22520 24012
rect 22376 20936 22428 20942
rect 22376 20878 22428 20884
rect 22100 20800 22152 20806
rect 22100 20742 22152 20748
rect 21928 19910 22048 19938
rect 21916 19848 21968 19854
rect 21916 19790 21968 19796
rect 21824 19304 21876 19310
rect 21824 19246 21876 19252
rect 21928 18834 21956 19790
rect 22020 18902 22048 19910
rect 22112 19310 22140 20742
rect 22284 19848 22336 19854
rect 22284 19790 22336 19796
rect 22192 19712 22244 19718
rect 22192 19654 22244 19660
rect 22204 19446 22232 19654
rect 22192 19440 22244 19446
rect 22192 19382 22244 19388
rect 22100 19304 22152 19310
rect 22100 19246 22152 19252
rect 22008 18896 22060 18902
rect 22008 18838 22060 18844
rect 21916 18828 21968 18834
rect 21916 18770 21968 18776
rect 21824 18760 21876 18766
rect 21824 18702 21876 18708
rect 21836 18222 21864 18702
rect 21928 18290 21956 18770
rect 22112 18737 22140 19246
rect 22098 18728 22154 18737
rect 22098 18663 22154 18672
rect 21916 18284 21968 18290
rect 21916 18226 21968 18232
rect 21824 18216 21876 18222
rect 21824 18158 21876 18164
rect 21560 18040 21772 18068
rect 21180 18022 21232 18028
rect 21272 17128 21324 17134
rect 21272 17070 21324 17076
rect 21284 16998 21312 17070
rect 21272 16992 21324 16998
rect 21272 16934 21324 16940
rect 21180 16040 21232 16046
rect 21180 15982 21232 15988
rect 21192 15706 21220 15982
rect 21284 15910 21312 16934
rect 21640 16448 21692 16454
rect 21640 16390 21692 16396
rect 21364 16176 21416 16182
rect 21364 16118 21416 16124
rect 21272 15904 21324 15910
rect 21272 15846 21324 15852
rect 21180 15700 21232 15706
rect 21180 15642 21232 15648
rect 21100 15014 21220 15042
rect 20996 14952 21048 14958
rect 20996 14894 21048 14900
rect 21088 14952 21140 14958
rect 21088 14894 21140 14900
rect 21100 13938 21128 14894
rect 21088 13932 21140 13938
rect 21088 13874 21140 13880
rect 20996 12980 21048 12986
rect 20996 12922 21048 12928
rect 20904 12912 20956 12918
rect 20904 12854 20956 12860
rect 20904 12776 20956 12782
rect 20904 12718 20956 12724
rect 20916 12170 20944 12718
rect 20904 12164 20956 12170
rect 20904 12106 20956 12112
rect 20824 11886 20944 11914
rect 20628 11630 20680 11636
rect 20718 11656 20774 11665
rect 20640 11558 20668 11630
rect 20718 11591 20774 11600
rect 20628 11552 20680 11558
rect 20628 11494 20680 11500
rect 20720 11008 20772 11014
rect 20720 10950 20772 10956
rect 20628 10464 20680 10470
rect 20628 10406 20680 10412
rect 20640 9382 20668 10406
rect 20628 9376 20680 9382
rect 20628 9318 20680 9324
rect 20536 9036 20588 9042
rect 20536 8978 20588 8984
rect 20444 8900 20496 8906
rect 20444 8842 20496 8848
rect 20456 7342 20484 8842
rect 20628 7812 20680 7818
rect 20628 7754 20680 7760
rect 20640 7342 20668 7754
rect 20444 7336 20496 7342
rect 20444 7278 20496 7284
rect 20628 7336 20680 7342
rect 20628 7278 20680 7284
rect 20456 6866 20484 7278
rect 20444 6860 20496 6866
rect 20444 6802 20496 6808
rect 20352 6248 20404 6254
rect 20352 6190 20404 6196
rect 19580 6012 19876 6032
rect 19636 6010 19660 6012
rect 19716 6010 19740 6012
rect 19796 6010 19820 6012
rect 19658 5958 19660 6010
rect 19722 5958 19734 6010
rect 19796 5958 19798 6010
rect 19636 5956 19660 5958
rect 19716 5956 19740 5958
rect 19796 5956 19820 5958
rect 19580 5936 19876 5956
rect 19340 5772 19392 5778
rect 19340 5714 19392 5720
rect 19248 5568 19300 5574
rect 19248 5510 19300 5516
rect 18880 5228 18932 5234
rect 18880 5170 18932 5176
rect 17960 5160 18012 5166
rect 17960 5102 18012 5108
rect 18512 5160 18564 5166
rect 18512 5102 18564 5108
rect 17776 4480 17828 4486
rect 17776 4422 17828 4428
rect 17866 3632 17922 3641
rect 17224 3596 17276 3602
rect 17866 3567 17922 3576
rect 17224 3538 17276 3544
rect 16304 3528 16356 3534
rect 16304 3470 16356 3476
rect 16120 3052 16172 3058
rect 16120 2994 16172 3000
rect 16028 2508 16080 2514
rect 16028 2450 16080 2456
rect 14188 2440 14240 2446
rect 14188 2382 14240 2388
rect 15844 2304 15896 2310
rect 15844 2246 15896 2252
rect 15856 800 15884 2246
rect 17880 800 17908 3567
rect 17972 3534 18000 5102
rect 18972 4684 19024 4690
rect 18972 4626 19024 4632
rect 19156 4684 19208 4690
rect 19156 4626 19208 4632
rect 18052 4480 18104 4486
rect 18052 4422 18104 4428
rect 18064 4078 18092 4422
rect 18984 4146 19012 4626
rect 19168 4214 19196 4626
rect 19156 4208 19208 4214
rect 19156 4150 19208 4156
rect 18972 4140 19024 4146
rect 18972 4082 19024 4088
rect 18052 4072 18104 4078
rect 18052 4014 18104 4020
rect 17960 3528 18012 3534
rect 17960 3470 18012 3476
rect 18984 2990 19012 4082
rect 18972 2984 19024 2990
rect 18972 2926 19024 2932
rect 19260 2582 19288 5510
rect 19352 5148 19380 5714
rect 20364 5710 20392 6190
rect 20352 5704 20404 5710
rect 20352 5646 20404 5652
rect 19432 5160 19484 5166
rect 19352 5120 19432 5148
rect 19352 4078 19380 5120
rect 19432 5102 19484 5108
rect 19432 5024 19484 5030
rect 19432 4966 19484 4972
rect 19340 4072 19392 4078
rect 19340 4014 19392 4020
rect 19444 2990 19472 4966
rect 19580 4924 19876 4944
rect 19636 4922 19660 4924
rect 19716 4922 19740 4924
rect 19796 4922 19820 4924
rect 19658 4870 19660 4922
rect 19722 4870 19734 4922
rect 19796 4870 19798 4922
rect 19636 4868 19660 4870
rect 19716 4868 19740 4870
rect 19796 4868 19820 4870
rect 19580 4848 19876 4868
rect 20640 4758 20668 7278
rect 20732 6458 20760 10950
rect 20812 10804 20864 10810
rect 20812 10746 20864 10752
rect 20824 10606 20852 10746
rect 20812 10600 20864 10606
rect 20812 10542 20864 10548
rect 20916 6730 20944 11886
rect 21008 11694 21036 12922
rect 21100 12306 21128 13874
rect 21192 13394 21220 15014
rect 21272 15020 21324 15026
rect 21272 14962 21324 14968
rect 21180 13388 21232 13394
rect 21180 13330 21232 13336
rect 21088 12300 21140 12306
rect 21088 12242 21140 12248
rect 20996 11688 21048 11694
rect 20996 11630 21048 11636
rect 20996 11212 21048 11218
rect 20996 11154 21048 11160
rect 21008 10606 21036 11154
rect 20996 10600 21048 10606
rect 20996 10542 21048 10548
rect 21088 10464 21140 10470
rect 21088 10406 21140 10412
rect 21100 9518 21128 10406
rect 21192 9586 21220 13330
rect 21284 11014 21312 14962
rect 21272 11008 21324 11014
rect 21272 10950 21324 10956
rect 21272 10056 21324 10062
rect 21272 9998 21324 10004
rect 21284 9586 21312 9998
rect 21180 9580 21232 9586
rect 21180 9522 21232 9528
rect 21272 9580 21324 9586
rect 21272 9522 21324 9528
rect 21088 9512 21140 9518
rect 21376 9466 21404 16118
rect 21652 15910 21680 16390
rect 21640 15904 21692 15910
rect 21640 15846 21692 15852
rect 21456 13388 21508 13394
rect 21456 13330 21508 13336
rect 21468 11354 21496 13330
rect 21548 11620 21600 11626
rect 21548 11562 21600 11568
rect 21560 11354 21588 11562
rect 21456 11348 21508 11354
rect 21456 11290 21508 11296
rect 21548 11348 21600 11354
rect 21548 11290 21600 11296
rect 21456 10124 21508 10130
rect 21456 10066 21508 10072
rect 21088 9454 21140 9460
rect 21284 9438 21404 9466
rect 21180 8900 21232 8906
rect 21180 8842 21232 8848
rect 21192 8673 21220 8842
rect 21178 8664 21234 8673
rect 21178 8599 21234 8608
rect 20996 8288 21048 8294
rect 20996 8230 21048 8236
rect 21088 8288 21140 8294
rect 21088 8230 21140 8236
rect 21008 7886 21036 8230
rect 21100 7954 21128 8230
rect 21088 7948 21140 7954
rect 21088 7890 21140 7896
rect 20996 7880 21048 7886
rect 20996 7822 21048 7828
rect 21088 7540 21140 7546
rect 21088 7482 21140 7488
rect 21100 7206 21128 7482
rect 21088 7200 21140 7206
rect 21088 7142 21140 7148
rect 21100 6866 21128 7142
rect 21088 6860 21140 6866
rect 21088 6802 21140 6808
rect 21284 6798 21312 9438
rect 21468 8634 21496 10066
rect 21652 9654 21680 15846
rect 21744 15042 21772 18040
rect 21824 17672 21876 17678
rect 21824 17614 21876 17620
rect 21836 16590 21864 17614
rect 22192 16992 22244 16998
rect 22192 16934 22244 16940
rect 22204 16726 22232 16934
rect 22192 16720 22244 16726
rect 22192 16662 22244 16668
rect 21916 16652 21968 16658
rect 21916 16594 21968 16600
rect 21824 16584 21876 16590
rect 21824 16526 21876 16532
rect 21928 16182 21956 16594
rect 21916 16176 21968 16182
rect 21916 16118 21968 16124
rect 21824 15972 21876 15978
rect 21824 15914 21876 15920
rect 21836 15162 21864 15914
rect 22100 15564 22152 15570
rect 22100 15506 22152 15512
rect 21824 15156 21876 15162
rect 21824 15098 21876 15104
rect 21744 15014 21864 15042
rect 21640 9648 21692 9654
rect 21640 9590 21692 9596
rect 21652 9450 21680 9590
rect 21836 9450 21864 15014
rect 22112 14822 22140 15506
rect 22192 15496 22244 15502
rect 22192 15438 22244 15444
rect 22100 14816 22152 14822
rect 22100 14758 22152 14764
rect 21916 13184 21968 13190
rect 21916 13126 21968 13132
rect 21928 12782 21956 13126
rect 22112 12850 22140 14758
rect 22204 14482 22232 15438
rect 22296 15366 22324 19790
rect 22480 18834 22508 24006
rect 22572 23322 22600 24228
rect 22652 24210 22704 24216
rect 22756 23730 22784 24806
rect 22744 23724 22796 23730
rect 22744 23666 22796 23672
rect 22652 23656 22704 23662
rect 22652 23598 22704 23604
rect 22560 23316 22612 23322
rect 22560 23258 22612 23264
rect 22664 23254 22692 23598
rect 22652 23248 22704 23254
rect 22652 23190 22704 23196
rect 22664 22098 22692 23190
rect 22652 22092 22704 22098
rect 22652 22034 22704 22040
rect 22560 21616 22612 21622
rect 22560 21558 22612 21564
rect 22572 21486 22600 21558
rect 22848 21486 22876 24822
rect 22560 21480 22612 21486
rect 22836 21480 22888 21486
rect 22612 21440 22692 21468
rect 22560 21422 22612 21428
rect 22560 21344 22612 21350
rect 22560 21286 22612 21292
rect 22572 21010 22600 21286
rect 22560 21004 22612 21010
rect 22560 20946 22612 20952
rect 22664 20942 22692 21440
rect 22836 21422 22888 21428
rect 22848 21078 22876 21422
rect 22836 21072 22888 21078
rect 22836 21014 22888 21020
rect 22652 20936 22704 20942
rect 22652 20878 22704 20884
rect 22744 20800 22796 20806
rect 22744 20742 22796 20748
rect 22468 18828 22520 18834
rect 22468 18770 22520 18776
rect 22376 18624 22428 18630
rect 22376 18566 22428 18572
rect 22388 16658 22416 18566
rect 22480 17882 22508 18770
rect 22468 17876 22520 17882
rect 22468 17818 22520 17824
rect 22560 17740 22612 17746
rect 22560 17682 22612 17688
rect 22572 16998 22600 17682
rect 22560 16992 22612 16998
rect 22560 16934 22612 16940
rect 22376 16652 22428 16658
rect 22376 16594 22428 16600
rect 22388 16114 22416 16594
rect 22468 16584 22520 16590
rect 22468 16526 22520 16532
rect 22376 16108 22428 16114
rect 22376 16050 22428 16056
rect 22388 15722 22416 16050
rect 22480 16046 22508 16526
rect 22468 16040 22520 16046
rect 22468 15982 22520 15988
rect 22388 15694 22508 15722
rect 22480 15570 22508 15694
rect 22376 15564 22428 15570
rect 22376 15506 22428 15512
rect 22468 15564 22520 15570
rect 22468 15506 22520 15512
rect 22284 15360 22336 15366
rect 22284 15302 22336 15308
rect 22192 14476 22244 14482
rect 22192 14418 22244 14424
rect 22192 13932 22244 13938
rect 22192 13874 22244 13880
rect 22284 13932 22336 13938
rect 22284 13874 22336 13880
rect 22204 13530 22232 13874
rect 22192 13524 22244 13530
rect 22192 13466 22244 13472
rect 22296 13258 22324 13874
rect 22284 13252 22336 13258
rect 22284 13194 22336 13200
rect 22284 12980 22336 12986
rect 22284 12922 22336 12928
rect 22100 12844 22152 12850
rect 22100 12786 22152 12792
rect 21916 12776 21968 12782
rect 21916 12718 21968 12724
rect 21928 11150 21956 12718
rect 22008 11688 22060 11694
rect 22060 11636 22232 11642
rect 22008 11630 22232 11636
rect 22020 11626 22232 11630
rect 22020 11620 22244 11626
rect 22020 11614 22192 11620
rect 22192 11562 22244 11568
rect 22008 11552 22060 11558
rect 22008 11494 22060 11500
rect 21916 11144 21968 11150
rect 21916 11086 21968 11092
rect 21928 10606 21956 11086
rect 22020 10674 22048 11494
rect 22192 11212 22244 11218
rect 22192 11154 22244 11160
rect 22008 10668 22060 10674
rect 22008 10610 22060 10616
rect 21916 10600 21968 10606
rect 21916 10542 21968 10548
rect 21640 9444 21692 9450
rect 21640 9386 21692 9392
rect 21824 9444 21876 9450
rect 21824 9386 21876 9392
rect 21916 9104 21968 9110
rect 21916 9046 21968 9052
rect 21732 9036 21784 9042
rect 21732 8978 21784 8984
rect 21456 8628 21508 8634
rect 21456 8570 21508 8576
rect 21468 7274 21496 8570
rect 21744 7410 21772 8978
rect 21928 8498 21956 9046
rect 21916 8492 21968 8498
rect 21916 8434 21968 8440
rect 22020 8430 22048 10610
rect 22204 9994 22232 11154
rect 22192 9988 22244 9994
rect 22192 9930 22244 9936
rect 22296 9330 22324 12922
rect 22204 9302 22324 9330
rect 22204 9042 22232 9302
rect 22284 9172 22336 9178
rect 22284 9114 22336 9120
rect 22192 9036 22244 9042
rect 22192 8978 22244 8984
rect 22008 8424 22060 8430
rect 22008 8366 22060 8372
rect 21822 7984 21878 7993
rect 21822 7919 21878 7928
rect 21836 7886 21864 7919
rect 21824 7880 21876 7886
rect 21824 7822 21876 7828
rect 22020 7750 22048 8366
rect 22204 8294 22232 8978
rect 22296 8430 22324 9114
rect 22388 8650 22416 15506
rect 22572 15450 22600 16934
rect 22652 16652 22704 16658
rect 22652 16594 22704 16600
rect 22664 15570 22692 16594
rect 22652 15564 22704 15570
rect 22652 15506 22704 15512
rect 22480 15422 22600 15450
rect 22480 12986 22508 15422
rect 22560 13864 22612 13870
rect 22560 13806 22612 13812
rect 22468 12980 22520 12986
rect 22468 12922 22520 12928
rect 22572 12102 22600 13806
rect 22652 13320 22704 13326
rect 22652 13262 22704 13268
rect 22664 12918 22692 13262
rect 22652 12912 22704 12918
rect 22652 12854 22704 12860
rect 22652 12776 22704 12782
rect 22652 12718 22704 12724
rect 22560 12096 22612 12102
rect 22560 12038 22612 12044
rect 22664 11830 22692 12718
rect 22652 11824 22704 11830
rect 22652 11766 22704 11772
rect 22652 11688 22704 11694
rect 22652 11630 22704 11636
rect 22560 11076 22612 11082
rect 22664 11064 22692 11630
rect 22612 11036 22692 11064
rect 22560 11018 22612 11024
rect 22560 10260 22612 10266
rect 22560 10202 22612 10208
rect 22572 9518 22600 10202
rect 22560 9512 22612 9518
rect 22560 9454 22612 9460
rect 22756 8906 22784 20742
rect 22928 20392 22980 20398
rect 22928 20334 22980 20340
rect 22836 20256 22888 20262
rect 22836 20198 22888 20204
rect 22848 19990 22876 20198
rect 22836 19984 22888 19990
rect 22836 19926 22888 19932
rect 22836 19848 22888 19854
rect 22940 19836 22968 20334
rect 23032 19961 23060 26726
rect 23124 26710 23244 26738
rect 23112 26376 23164 26382
rect 23112 26318 23164 26324
rect 23124 24070 23152 26318
rect 23112 24064 23164 24070
rect 23112 24006 23164 24012
rect 23112 20868 23164 20874
rect 23112 20810 23164 20816
rect 23018 19952 23074 19961
rect 23018 19887 23020 19896
rect 23072 19887 23074 19896
rect 23020 19858 23072 19864
rect 22888 19808 22968 19836
rect 22836 19790 22888 19796
rect 22848 19310 22876 19790
rect 22836 19304 22888 19310
rect 22836 19246 22888 19252
rect 22928 19304 22980 19310
rect 22928 19246 22980 19252
rect 22848 18902 22876 19246
rect 22836 18896 22888 18902
rect 22836 18838 22888 18844
rect 22836 18352 22888 18358
rect 22836 18294 22888 18300
rect 22848 17542 22876 18294
rect 22836 17536 22888 17542
rect 22836 17478 22888 17484
rect 22848 17134 22876 17478
rect 22836 17128 22888 17134
rect 22836 17070 22888 17076
rect 22940 15910 22968 19246
rect 22928 15904 22980 15910
rect 22928 15846 22980 15852
rect 23020 15496 23072 15502
rect 23020 15438 23072 15444
rect 22928 14952 22980 14958
rect 22928 14894 22980 14900
rect 22836 14884 22888 14890
rect 22836 14826 22888 14832
rect 22848 12986 22876 14826
rect 22940 14618 22968 14894
rect 23032 14822 23060 15438
rect 23020 14816 23072 14822
rect 23020 14758 23072 14764
rect 22928 14612 22980 14618
rect 22928 14554 22980 14560
rect 23124 13138 23152 20810
rect 23216 14006 23244 26710
rect 23584 26382 23612 26862
rect 23572 26376 23624 26382
rect 23572 26318 23624 26324
rect 23296 26240 23348 26246
rect 23296 26182 23348 26188
rect 23308 25362 23336 26182
rect 23572 26036 23624 26042
rect 23572 25978 23624 25984
rect 23584 25838 23612 25978
rect 23572 25832 23624 25838
rect 23572 25774 23624 25780
rect 23296 25356 23348 25362
rect 23296 25298 23348 25304
rect 23480 24812 23532 24818
rect 23480 24754 23532 24760
rect 23492 23186 23520 24754
rect 23676 24154 23704 31826
rect 23848 31680 23900 31686
rect 23848 31622 23900 31628
rect 23756 31272 23808 31278
rect 23756 31214 23808 31220
rect 23768 30394 23796 31214
rect 23756 30388 23808 30394
rect 23756 30330 23808 30336
rect 23860 30190 23888 31622
rect 23848 30184 23900 30190
rect 23848 30126 23900 30132
rect 23940 29232 23992 29238
rect 23940 29174 23992 29180
rect 23848 29096 23900 29102
rect 23952 29073 23980 29174
rect 24032 29096 24084 29102
rect 23848 29038 23900 29044
rect 23938 29064 23994 29073
rect 23756 28620 23808 28626
rect 23756 28562 23808 28568
rect 23768 25362 23796 28562
rect 23860 28064 23888 29038
rect 24136 29084 24164 36654
rect 24320 34610 24348 36654
rect 24872 35630 24900 37266
rect 24964 36922 24992 38286
rect 26424 38208 26476 38214
rect 26424 38150 26476 38156
rect 26436 37874 26464 38150
rect 26424 37868 26476 37874
rect 26424 37810 26476 37816
rect 25780 37800 25832 37806
rect 25780 37742 25832 37748
rect 25792 37262 25820 37742
rect 26608 37324 26660 37330
rect 26608 37266 26660 37272
rect 25780 37256 25832 37262
rect 25780 37198 25832 37204
rect 24952 36916 25004 36922
rect 24952 36858 25004 36864
rect 25792 36786 25820 37198
rect 25780 36780 25832 36786
rect 25780 36722 25832 36728
rect 25136 36576 25188 36582
rect 25136 36518 25188 36524
rect 24860 35624 24912 35630
rect 24860 35566 24912 35572
rect 25044 35624 25096 35630
rect 25044 35566 25096 35572
rect 25056 34610 25084 35566
rect 24308 34604 24360 34610
rect 24308 34546 24360 34552
rect 25044 34604 25096 34610
rect 25044 34546 25096 34552
rect 24584 33992 24636 33998
rect 24584 33934 24636 33940
rect 24596 33658 24624 33934
rect 24584 33652 24636 33658
rect 24584 33594 24636 33600
rect 24400 33516 24452 33522
rect 24400 33458 24452 33464
rect 24412 32366 24440 33458
rect 25044 33448 25096 33454
rect 25044 33390 25096 33396
rect 24492 33108 24544 33114
rect 24492 33050 24544 33056
rect 24400 32360 24452 32366
rect 24400 32302 24452 32308
rect 24308 31952 24360 31958
rect 24308 31894 24360 31900
rect 24216 30796 24268 30802
rect 24216 30738 24268 30744
rect 24228 30326 24256 30738
rect 24216 30320 24268 30326
rect 24216 30262 24268 30268
rect 24320 30190 24348 31894
rect 24504 30258 24532 33050
rect 24860 32904 24912 32910
rect 24860 32846 24912 32852
rect 24584 32768 24636 32774
rect 24584 32710 24636 32716
rect 24492 30252 24544 30258
rect 24492 30194 24544 30200
rect 24308 30184 24360 30190
rect 24308 30126 24360 30132
rect 24492 29776 24544 29782
rect 24492 29718 24544 29724
rect 24400 29708 24452 29714
rect 24400 29650 24452 29656
rect 24214 29608 24270 29617
rect 24214 29543 24216 29552
rect 24268 29543 24270 29552
rect 24216 29514 24268 29520
rect 24412 29238 24440 29650
rect 24400 29232 24452 29238
rect 24400 29174 24452 29180
rect 24504 29102 24532 29718
rect 24596 29102 24624 32710
rect 24768 31952 24820 31958
rect 24768 31894 24820 31900
rect 24674 29336 24730 29345
rect 24674 29271 24730 29280
rect 24084 29056 24164 29084
rect 24492 29096 24544 29102
rect 24032 29038 24084 29044
rect 24492 29038 24544 29044
rect 24584 29096 24636 29102
rect 24584 29038 24636 29044
rect 23938 28999 23994 29008
rect 24400 28552 24452 28558
rect 24504 28540 24532 29038
rect 24688 28948 24716 29271
rect 24596 28920 24716 28948
rect 24596 28626 24624 28920
rect 24584 28620 24636 28626
rect 24584 28562 24636 28568
rect 24452 28512 24532 28540
rect 24400 28494 24452 28500
rect 24124 28416 24176 28422
rect 24124 28358 24176 28364
rect 24136 28150 24164 28358
rect 24124 28144 24176 28150
rect 24124 28086 24176 28092
rect 24032 28076 24084 28082
rect 23860 28036 24032 28064
rect 24032 28018 24084 28024
rect 24308 28076 24360 28082
rect 24308 28018 24360 28024
rect 24032 27872 24084 27878
rect 24032 27814 24084 27820
rect 24044 27674 24072 27814
rect 24032 27668 24084 27674
rect 24032 27610 24084 27616
rect 23940 27464 23992 27470
rect 23940 27406 23992 27412
rect 23848 26444 23900 26450
rect 23848 26386 23900 26392
rect 23860 25702 23888 26386
rect 23952 26314 23980 27406
rect 24032 27396 24084 27402
rect 24032 27338 24084 27344
rect 24044 26994 24072 27338
rect 24032 26988 24084 26994
rect 24032 26930 24084 26936
rect 23940 26308 23992 26314
rect 23940 26250 23992 26256
rect 23848 25696 23900 25702
rect 23848 25638 23900 25644
rect 23952 25430 23980 26250
rect 23940 25424 23992 25430
rect 23940 25366 23992 25372
rect 23756 25356 23808 25362
rect 23756 25298 23808 25304
rect 23848 25356 23900 25362
rect 23848 25298 23900 25304
rect 23860 24954 23888 25298
rect 23848 24948 23900 24954
rect 23848 24890 23900 24896
rect 23940 24948 23992 24954
rect 23940 24890 23992 24896
rect 23860 24410 23888 24890
rect 23848 24404 23900 24410
rect 23848 24346 23900 24352
rect 23848 24268 23900 24274
rect 23848 24210 23900 24216
rect 23676 24126 23796 24154
rect 23664 23724 23716 23730
rect 23664 23666 23716 23672
rect 23480 23180 23532 23186
rect 23480 23122 23532 23128
rect 23492 21554 23520 23122
rect 23676 23118 23704 23666
rect 23572 23112 23624 23118
rect 23572 23054 23624 23060
rect 23664 23112 23716 23118
rect 23664 23054 23716 23060
rect 23480 21548 23532 21554
rect 23480 21490 23532 21496
rect 23296 21344 23348 21350
rect 23296 21286 23348 21292
rect 23388 21344 23440 21350
rect 23388 21286 23440 21292
rect 23308 16590 23336 21286
rect 23400 21010 23428 21286
rect 23388 21004 23440 21010
rect 23388 20946 23440 20952
rect 23400 19378 23428 20946
rect 23388 19372 23440 19378
rect 23388 19314 23440 19320
rect 23584 19174 23612 23054
rect 23676 22574 23704 23054
rect 23664 22568 23716 22574
rect 23664 22510 23716 22516
rect 23768 22522 23796 24126
rect 23860 23662 23888 24210
rect 23848 23656 23900 23662
rect 23848 23598 23900 23604
rect 23952 22642 23980 24890
rect 24320 24410 24348 28018
rect 24504 27538 24532 28512
rect 24780 28422 24808 31894
rect 24768 28416 24820 28422
rect 24768 28358 24820 28364
rect 24768 27940 24820 27946
rect 24768 27882 24820 27888
rect 24780 27606 24808 27882
rect 24768 27600 24820 27606
rect 24768 27542 24820 27548
rect 24492 27532 24544 27538
rect 24492 27474 24544 27480
rect 24780 26994 24808 27542
rect 24872 27334 24900 32846
rect 24952 29028 25004 29034
rect 24952 28970 25004 28976
rect 24964 28626 24992 28970
rect 24952 28620 25004 28626
rect 24952 28562 25004 28568
rect 24860 27328 24912 27334
rect 24860 27270 24912 27276
rect 24768 26988 24820 26994
rect 24768 26930 24820 26936
rect 24492 26444 24544 26450
rect 24492 26386 24544 26392
rect 24504 25158 24532 26386
rect 24584 26240 24636 26246
rect 24584 26182 24636 26188
rect 24596 25838 24624 26182
rect 25056 25888 25084 33390
rect 25148 31278 25176 36518
rect 25412 36168 25464 36174
rect 25412 36110 25464 36116
rect 25424 35086 25452 36110
rect 25792 35834 25820 36722
rect 26056 36712 26108 36718
rect 26056 36654 26108 36660
rect 26068 36310 26096 36654
rect 26424 36576 26476 36582
rect 26424 36518 26476 36524
rect 26056 36304 26108 36310
rect 26056 36246 26108 36252
rect 25872 36032 25924 36038
rect 25872 35974 25924 35980
rect 25780 35828 25832 35834
rect 25780 35770 25832 35776
rect 25504 35488 25556 35494
rect 25504 35430 25556 35436
rect 25516 35154 25544 35430
rect 25884 35222 25912 35974
rect 26332 35828 26384 35834
rect 26332 35770 26384 35776
rect 26240 35760 26292 35766
rect 26240 35702 26292 35708
rect 25872 35216 25924 35222
rect 25872 35158 25924 35164
rect 25504 35148 25556 35154
rect 25504 35090 25556 35096
rect 25412 35080 25464 35086
rect 25412 35022 25464 35028
rect 25688 34740 25740 34746
rect 25688 34682 25740 34688
rect 25504 32972 25556 32978
rect 25504 32914 25556 32920
rect 25320 32360 25372 32366
rect 25320 32302 25372 32308
rect 25228 32224 25280 32230
rect 25228 32166 25280 32172
rect 25240 31890 25268 32166
rect 25228 31884 25280 31890
rect 25228 31826 25280 31832
rect 25136 31272 25188 31278
rect 25136 31214 25188 31220
rect 25226 30832 25282 30841
rect 25226 30767 25228 30776
rect 25280 30767 25282 30776
rect 25228 30738 25280 30744
rect 25332 30258 25360 32302
rect 25516 31793 25544 32914
rect 25700 31890 25728 34682
rect 25688 31884 25740 31890
rect 25688 31826 25740 31832
rect 25502 31784 25558 31793
rect 25502 31719 25558 31728
rect 25688 31748 25740 31754
rect 25412 30796 25464 30802
rect 25412 30738 25464 30744
rect 25320 30252 25372 30258
rect 25320 30194 25372 30200
rect 25320 29776 25372 29782
rect 25320 29718 25372 29724
rect 25332 29306 25360 29718
rect 25320 29300 25372 29306
rect 25320 29242 25372 29248
rect 25424 28098 25452 30738
rect 25516 30394 25544 31719
rect 25688 31690 25740 31696
rect 25700 31210 25728 31690
rect 25780 31272 25832 31278
rect 25780 31214 25832 31220
rect 25688 31204 25740 31210
rect 25688 31146 25740 31152
rect 25504 30388 25556 30394
rect 25504 30330 25556 30336
rect 25504 30252 25556 30258
rect 25504 30194 25556 30200
rect 25516 29714 25544 30194
rect 25504 29708 25556 29714
rect 25504 29650 25556 29656
rect 25516 28218 25544 29650
rect 25700 29578 25728 31146
rect 25792 30802 25820 31214
rect 25780 30796 25832 30802
rect 25780 30738 25832 30744
rect 25688 29572 25740 29578
rect 25688 29514 25740 29520
rect 25504 28212 25556 28218
rect 25504 28154 25556 28160
rect 25424 28070 25544 28098
rect 25412 28008 25464 28014
rect 25412 27950 25464 27956
rect 25424 27674 25452 27950
rect 25412 27668 25464 27674
rect 25412 27610 25464 27616
rect 25412 27532 25464 27538
rect 25412 27474 25464 27480
rect 25320 27056 25372 27062
rect 25320 26998 25372 27004
rect 25332 26450 25360 26998
rect 25424 26858 25452 27474
rect 25412 26852 25464 26858
rect 25412 26794 25464 26800
rect 25320 26444 25372 26450
rect 25320 26386 25372 26392
rect 25228 25968 25280 25974
rect 25228 25910 25280 25916
rect 25056 25860 25176 25888
rect 24584 25832 24636 25838
rect 24584 25774 24636 25780
rect 24492 25152 24544 25158
rect 24492 25094 24544 25100
rect 24596 24750 24624 25774
rect 25044 25764 25096 25770
rect 25044 25706 25096 25712
rect 25056 25362 25084 25706
rect 25044 25356 25096 25362
rect 25044 25298 25096 25304
rect 24952 25220 25004 25226
rect 24952 25162 25004 25168
rect 24964 24818 24992 25162
rect 25148 24834 25176 25860
rect 25240 25362 25268 25910
rect 25228 25356 25280 25362
rect 25228 25298 25280 25304
rect 24952 24812 25004 24818
rect 25148 24806 25268 24834
rect 24952 24754 25004 24760
rect 24400 24744 24452 24750
rect 24400 24686 24452 24692
rect 24584 24744 24636 24750
rect 24584 24686 24636 24692
rect 24308 24404 24360 24410
rect 24308 24346 24360 24352
rect 24412 23662 24440 24686
rect 24400 23656 24452 23662
rect 24400 23598 24452 23604
rect 24412 23322 24440 23598
rect 24400 23316 24452 23322
rect 24400 23258 24452 23264
rect 24216 23180 24268 23186
rect 24216 23122 24268 23128
rect 23940 22636 23992 22642
rect 23940 22578 23992 22584
rect 23768 22494 23980 22522
rect 23664 22092 23716 22098
rect 23664 22034 23716 22040
rect 23676 21894 23704 22034
rect 23848 21956 23900 21962
rect 23848 21898 23900 21904
rect 23664 21888 23716 21894
rect 23664 21830 23716 21836
rect 23676 19310 23704 21830
rect 23860 21554 23888 21898
rect 23848 21548 23900 21554
rect 23848 21490 23900 21496
rect 23756 21004 23808 21010
rect 23756 20946 23808 20952
rect 23768 20534 23796 20946
rect 23756 20528 23808 20534
rect 23756 20470 23808 20476
rect 23664 19304 23716 19310
rect 23664 19246 23716 19252
rect 23480 19168 23532 19174
rect 23480 19110 23532 19116
rect 23572 19168 23624 19174
rect 23572 19110 23624 19116
rect 23492 18986 23520 19110
rect 23492 18958 23796 18986
rect 23388 17536 23440 17542
rect 23388 17478 23440 17484
rect 23400 16658 23428 17478
rect 23572 16788 23624 16794
rect 23572 16730 23624 16736
rect 23388 16652 23440 16658
rect 23388 16594 23440 16600
rect 23480 16652 23532 16658
rect 23480 16594 23532 16600
rect 23296 16584 23348 16590
rect 23296 16526 23348 16532
rect 23388 16516 23440 16522
rect 23388 16458 23440 16464
rect 23400 15910 23428 16458
rect 23492 16114 23520 16594
rect 23584 16454 23612 16730
rect 23572 16448 23624 16454
rect 23572 16390 23624 16396
rect 23480 16108 23532 16114
rect 23480 16050 23532 16056
rect 23664 16040 23716 16046
rect 23664 15982 23716 15988
rect 23388 15904 23440 15910
rect 23388 15846 23440 15852
rect 23204 14000 23256 14006
rect 23204 13942 23256 13948
rect 23032 13110 23152 13138
rect 22836 12980 22888 12986
rect 22836 12922 22888 12928
rect 22848 12306 22876 12922
rect 23032 12442 23060 13110
rect 23020 12436 23072 12442
rect 23020 12378 23072 12384
rect 22836 12300 22888 12306
rect 22836 12242 22888 12248
rect 22836 12164 22888 12170
rect 22836 12106 22888 12112
rect 22744 8900 22796 8906
rect 22744 8842 22796 8848
rect 22388 8622 22508 8650
rect 22376 8492 22428 8498
rect 22376 8434 22428 8440
rect 22284 8424 22336 8430
rect 22284 8366 22336 8372
rect 22192 8288 22244 8294
rect 22192 8230 22244 8236
rect 22100 8084 22152 8090
rect 22100 8026 22152 8032
rect 22008 7744 22060 7750
rect 22008 7686 22060 7692
rect 21732 7404 21784 7410
rect 21732 7346 21784 7352
rect 22112 7342 22140 8026
rect 22100 7336 22152 7342
rect 22100 7278 22152 7284
rect 21456 7268 21508 7274
rect 21456 7210 21508 7216
rect 22100 6860 22152 6866
rect 22100 6802 22152 6808
rect 21272 6792 21324 6798
rect 21272 6734 21324 6740
rect 20904 6724 20956 6730
rect 20904 6666 20956 6672
rect 20720 6452 20772 6458
rect 20720 6394 20772 6400
rect 20916 6254 20944 6666
rect 22112 6474 22140 6802
rect 22204 6662 22232 8230
rect 22284 7880 22336 7886
rect 22284 7822 22336 7828
rect 22296 7478 22324 7822
rect 22284 7472 22336 7478
rect 22284 7414 22336 7420
rect 22388 7342 22416 8434
rect 22376 7336 22428 7342
rect 22376 7278 22428 7284
rect 22192 6656 22244 6662
rect 22192 6598 22244 6604
rect 22112 6446 22232 6474
rect 22204 6254 22232 6446
rect 20904 6248 20956 6254
rect 20904 6190 20956 6196
rect 21272 6248 21324 6254
rect 21272 6190 21324 6196
rect 22192 6248 22244 6254
rect 22192 6190 22244 6196
rect 20904 6112 20956 6118
rect 20904 6054 20956 6060
rect 20916 5778 20944 6054
rect 21284 5778 21312 6190
rect 22204 5778 22232 6190
rect 20904 5772 20956 5778
rect 20904 5714 20956 5720
rect 21272 5772 21324 5778
rect 21272 5714 21324 5720
rect 22192 5772 22244 5778
rect 22192 5714 22244 5720
rect 20628 4752 20680 4758
rect 20628 4694 20680 4700
rect 19708 4616 19760 4622
rect 19708 4558 19760 4564
rect 19720 4146 19748 4558
rect 20916 4282 20944 5714
rect 22100 5704 22152 5710
rect 22100 5646 22152 5652
rect 21272 5636 21324 5642
rect 21272 5578 21324 5584
rect 21284 4622 21312 5578
rect 22112 5166 22140 5646
rect 22480 5302 22508 8622
rect 22652 8628 22704 8634
rect 22652 8570 22704 8576
rect 22560 8424 22612 8430
rect 22664 8401 22692 8570
rect 22560 8366 22612 8372
rect 22650 8392 22706 8401
rect 22572 8090 22600 8366
rect 22650 8327 22706 8336
rect 22848 8294 22876 12106
rect 22928 11688 22980 11694
rect 22928 11630 22980 11636
rect 22940 10606 22968 11630
rect 23032 11218 23060 12378
rect 23400 11778 23428 15846
rect 23676 15570 23704 15982
rect 23664 15564 23716 15570
rect 23664 15506 23716 15512
rect 23480 14408 23532 14414
rect 23480 14350 23532 14356
rect 23124 11750 23428 11778
rect 23020 11212 23072 11218
rect 23020 11154 23072 11160
rect 22928 10600 22980 10606
rect 22928 10542 22980 10548
rect 22940 10266 22968 10542
rect 22928 10260 22980 10266
rect 22928 10202 22980 10208
rect 23032 9024 23060 11154
rect 23124 9178 23152 11750
rect 23204 11688 23256 11694
rect 23204 11630 23256 11636
rect 23216 11286 23244 11630
rect 23204 11280 23256 11286
rect 23204 11222 23256 11228
rect 23296 11144 23348 11150
rect 23296 11086 23348 11092
rect 23204 10532 23256 10538
rect 23204 10474 23256 10480
rect 23216 9382 23244 10474
rect 23308 9586 23336 11086
rect 23492 10470 23520 14350
rect 23676 13870 23704 15506
rect 23664 13864 23716 13870
rect 23664 13806 23716 13812
rect 23572 13388 23624 13394
rect 23572 13330 23624 13336
rect 23584 12646 23612 13330
rect 23664 13252 23716 13258
rect 23664 13194 23716 13200
rect 23572 12640 23624 12646
rect 23572 12582 23624 12588
rect 23676 11898 23704 13194
rect 23768 12374 23796 18958
rect 23848 18692 23900 18698
rect 23848 18634 23900 18640
rect 23860 17746 23888 18634
rect 23848 17740 23900 17746
rect 23848 17682 23900 17688
rect 23848 17536 23900 17542
rect 23848 17478 23900 17484
rect 23756 12368 23808 12374
rect 23756 12310 23808 12316
rect 23664 11892 23716 11898
rect 23664 11834 23716 11840
rect 23768 11234 23796 12310
rect 23860 11694 23888 17478
rect 23952 13462 23980 22494
rect 24228 22438 24256 23122
rect 24860 22568 24912 22574
rect 24860 22510 24912 22516
rect 24308 22500 24360 22506
rect 24308 22442 24360 22448
rect 24584 22500 24636 22506
rect 24584 22442 24636 22448
rect 24216 22432 24268 22438
rect 24216 22374 24268 22380
rect 24124 22024 24176 22030
rect 24124 21966 24176 21972
rect 24136 21010 24164 21966
rect 24124 21004 24176 21010
rect 24124 20946 24176 20952
rect 24228 20398 24256 22374
rect 24320 22098 24348 22442
rect 24308 22092 24360 22098
rect 24308 22034 24360 22040
rect 24596 21010 24624 22442
rect 24872 21146 24900 22510
rect 24860 21140 24912 21146
rect 24860 21082 24912 21088
rect 24584 21004 24636 21010
rect 24584 20946 24636 20952
rect 24216 20392 24268 20398
rect 24216 20334 24268 20340
rect 24492 20324 24544 20330
rect 24492 20266 24544 20272
rect 24400 20256 24452 20262
rect 24400 20198 24452 20204
rect 24032 19780 24084 19786
rect 24032 19722 24084 19728
rect 24124 19780 24176 19786
rect 24124 19722 24176 19728
rect 24044 19310 24072 19722
rect 24032 19304 24084 19310
rect 24032 19246 24084 19252
rect 24044 18834 24072 19246
rect 24136 19242 24164 19722
rect 24124 19236 24176 19242
rect 24124 19178 24176 19184
rect 24032 18828 24084 18834
rect 24032 18770 24084 18776
rect 24032 17128 24084 17134
rect 24032 17070 24084 17076
rect 24308 17128 24360 17134
rect 24308 17070 24360 17076
rect 24044 16590 24072 17070
rect 24032 16584 24084 16590
rect 24084 16544 24164 16572
rect 24032 16526 24084 16532
rect 24136 14958 24164 16544
rect 24216 16448 24268 16454
rect 24216 16390 24268 16396
rect 24228 16046 24256 16390
rect 24320 16114 24348 17070
rect 24308 16108 24360 16114
rect 24308 16050 24360 16056
rect 24216 16040 24268 16046
rect 24216 15982 24268 15988
rect 24124 14952 24176 14958
rect 24124 14894 24176 14900
rect 24136 14414 24164 14894
rect 24124 14408 24176 14414
rect 24124 14350 24176 14356
rect 24124 14272 24176 14278
rect 24124 14214 24176 14220
rect 24136 13870 24164 14214
rect 24124 13864 24176 13870
rect 24124 13806 24176 13812
rect 23940 13456 23992 13462
rect 23940 13398 23992 13404
rect 24228 13326 24256 15982
rect 24412 15722 24440 20198
rect 24504 17626 24532 20266
rect 24596 19922 24624 20946
rect 24768 20800 24820 20806
rect 24768 20742 24820 20748
rect 24780 20058 24808 20742
rect 24860 20392 24912 20398
rect 24860 20334 24912 20340
rect 24768 20052 24820 20058
rect 24768 19994 24820 20000
rect 24584 19916 24636 19922
rect 24584 19858 24636 19864
rect 24596 17746 24624 19858
rect 24676 19304 24728 19310
rect 24676 19246 24728 19252
rect 24688 18766 24716 19246
rect 24676 18760 24728 18766
rect 24676 18702 24728 18708
rect 24768 18216 24820 18222
rect 24872 18204 24900 20334
rect 25136 18896 25188 18902
rect 25136 18838 25188 18844
rect 25148 18222 25176 18838
rect 24820 18176 24900 18204
rect 24952 18216 25004 18222
rect 24768 18158 24820 18164
rect 24952 18158 25004 18164
rect 25136 18216 25188 18222
rect 25136 18158 25188 18164
rect 24584 17740 24636 17746
rect 24584 17682 24636 17688
rect 24768 17672 24820 17678
rect 24504 17598 24716 17626
rect 24768 17614 24820 17620
rect 24412 15694 24624 15722
rect 24400 15496 24452 15502
rect 24400 15438 24452 15444
rect 24308 15020 24360 15026
rect 24308 14962 24360 14968
rect 24320 13938 24348 14962
rect 24412 14482 24440 15438
rect 24492 15020 24544 15026
rect 24492 14962 24544 14968
rect 24400 14476 24452 14482
rect 24400 14418 24452 14424
rect 24308 13932 24360 13938
rect 24308 13874 24360 13880
rect 24216 13320 24268 13326
rect 24216 13262 24268 13268
rect 24504 12238 24532 14962
rect 24124 12232 24176 12238
rect 24124 12174 24176 12180
rect 24492 12232 24544 12238
rect 24492 12174 24544 12180
rect 23848 11688 23900 11694
rect 23848 11630 23900 11636
rect 23940 11620 23992 11626
rect 23940 11562 23992 11568
rect 23768 11218 23888 11234
rect 23768 11212 23900 11218
rect 23768 11206 23848 11212
rect 23768 10606 23796 11206
rect 23848 11154 23900 11160
rect 23756 10600 23808 10606
rect 23756 10542 23808 10548
rect 23848 10532 23900 10538
rect 23848 10474 23900 10480
rect 23480 10464 23532 10470
rect 23480 10406 23532 10412
rect 23492 10130 23520 10406
rect 23480 10124 23532 10130
rect 23480 10066 23532 10072
rect 23296 9580 23348 9586
rect 23296 9522 23348 9528
rect 23204 9376 23256 9382
rect 23204 9318 23256 9324
rect 23112 9172 23164 9178
rect 23112 9114 23164 9120
rect 23112 9036 23164 9042
rect 23032 8996 23112 9024
rect 23112 8978 23164 8984
rect 22836 8288 22888 8294
rect 22836 8230 22888 8236
rect 22560 8084 22612 8090
rect 22560 8026 22612 8032
rect 23018 7984 23074 7993
rect 23124 7954 23152 8978
rect 23018 7919 23074 7928
rect 23112 7948 23164 7954
rect 22928 7200 22980 7206
rect 22928 7142 22980 7148
rect 22744 5772 22796 5778
rect 22744 5714 22796 5720
rect 22468 5296 22520 5302
rect 22468 5238 22520 5244
rect 22100 5160 22152 5166
rect 22100 5102 22152 5108
rect 22480 4826 22508 5238
rect 22756 5166 22784 5714
rect 22744 5160 22796 5166
rect 22744 5102 22796 5108
rect 22836 5160 22888 5166
rect 22836 5102 22888 5108
rect 22848 4826 22876 5102
rect 22468 4820 22520 4826
rect 22468 4762 22520 4768
rect 22836 4820 22888 4826
rect 22836 4762 22888 4768
rect 21272 4616 21324 4622
rect 21272 4558 21324 4564
rect 22836 4616 22888 4622
rect 22836 4558 22888 4564
rect 20904 4276 20956 4282
rect 20904 4218 20956 4224
rect 22848 4146 22876 4558
rect 19708 4140 19760 4146
rect 19708 4082 19760 4088
rect 20720 4140 20772 4146
rect 20720 4082 20772 4088
rect 22836 4140 22888 4146
rect 22836 4082 22888 4088
rect 20352 4072 20404 4078
rect 20352 4014 20404 4020
rect 19580 3836 19876 3856
rect 19636 3834 19660 3836
rect 19716 3834 19740 3836
rect 19796 3834 19820 3836
rect 19658 3782 19660 3834
rect 19722 3782 19734 3834
rect 19796 3782 19798 3834
rect 19636 3780 19660 3782
rect 19716 3780 19740 3782
rect 19796 3780 19820 3782
rect 19580 3760 19876 3780
rect 20364 3534 20392 4014
rect 20628 3936 20680 3942
rect 20628 3878 20680 3884
rect 20352 3528 20404 3534
rect 20352 3470 20404 3476
rect 20364 2990 20392 3470
rect 20640 2990 20668 3878
rect 20732 3194 20760 4082
rect 22100 4072 22152 4078
rect 21730 4040 21786 4049
rect 22100 4014 22152 4020
rect 21730 3975 21786 3984
rect 21088 3528 21140 3534
rect 21088 3470 21140 3476
rect 20720 3188 20772 3194
rect 20720 3130 20772 3136
rect 21100 3058 21128 3470
rect 21088 3052 21140 3058
rect 21088 2994 21140 3000
rect 19432 2984 19484 2990
rect 19432 2926 19484 2932
rect 20352 2984 20404 2990
rect 20352 2926 20404 2932
rect 20628 2984 20680 2990
rect 20628 2926 20680 2932
rect 19580 2748 19876 2768
rect 19636 2746 19660 2748
rect 19716 2746 19740 2748
rect 19796 2746 19820 2748
rect 19658 2694 19660 2746
rect 19722 2694 19734 2746
rect 19796 2694 19798 2746
rect 19636 2692 19660 2694
rect 19716 2692 19740 2694
rect 19796 2692 19820 2694
rect 19580 2672 19876 2692
rect 19248 2576 19300 2582
rect 19248 2518 19300 2524
rect 19708 2508 19760 2514
rect 19708 2450 19760 2456
rect 19720 800 19748 2450
rect 21744 800 21772 3975
rect 22112 2990 22140 4014
rect 22940 3602 22968 7142
rect 23032 5710 23060 7919
rect 23112 7890 23164 7896
rect 23216 7342 23244 9318
rect 23204 7336 23256 7342
rect 23204 7278 23256 7284
rect 23204 7200 23256 7206
rect 23204 7142 23256 7148
rect 23216 6934 23244 7142
rect 23204 6928 23256 6934
rect 23204 6870 23256 6876
rect 23020 5704 23072 5710
rect 23020 5646 23072 5652
rect 23032 3602 23060 5646
rect 23308 5574 23336 9522
rect 23860 9518 23888 10474
rect 23664 9512 23716 9518
rect 23662 9480 23664 9489
rect 23848 9512 23900 9518
rect 23716 9480 23718 9489
rect 23848 9454 23900 9460
rect 23662 9415 23718 9424
rect 23388 9376 23440 9382
rect 23388 9318 23440 9324
rect 23400 8362 23428 9318
rect 23860 9178 23888 9454
rect 23480 9172 23532 9178
rect 23480 9114 23532 9120
rect 23848 9172 23900 9178
rect 23848 9114 23900 9120
rect 23388 8356 23440 8362
rect 23388 8298 23440 8304
rect 23400 6458 23428 8298
rect 23492 8022 23520 9114
rect 23860 9042 23888 9114
rect 23848 9036 23900 9042
rect 23848 8978 23900 8984
rect 23664 8492 23716 8498
rect 23664 8434 23716 8440
rect 23480 8016 23532 8022
rect 23676 7993 23704 8434
rect 23952 8430 23980 11562
rect 24136 10198 24164 12174
rect 24308 11824 24360 11830
rect 24308 11766 24360 11772
rect 24320 10674 24348 11766
rect 24398 11248 24454 11257
rect 24398 11183 24454 11192
rect 24308 10668 24360 10674
rect 24308 10610 24360 10616
rect 24124 10192 24176 10198
rect 24124 10134 24176 10140
rect 24136 9994 24164 10134
rect 24216 10056 24268 10062
rect 24216 9998 24268 10004
rect 24124 9988 24176 9994
rect 24124 9930 24176 9936
rect 24228 9654 24256 9998
rect 24216 9648 24268 9654
rect 24216 9590 24268 9596
rect 24320 9518 24348 10610
rect 24412 10470 24440 11183
rect 24492 11008 24544 11014
rect 24492 10950 24544 10956
rect 24400 10464 24452 10470
rect 24400 10406 24452 10412
rect 24504 10062 24532 10950
rect 24596 10606 24624 15694
rect 24688 14618 24716 17598
rect 24780 15026 24808 17614
rect 24964 16998 24992 18158
rect 24952 16992 25004 16998
rect 24952 16934 25004 16940
rect 24768 15020 24820 15026
rect 24768 14962 24820 14968
rect 24860 14952 24912 14958
rect 24860 14894 24912 14900
rect 24676 14612 24728 14618
rect 24676 14554 24728 14560
rect 24872 14074 24900 14894
rect 24860 14068 24912 14074
rect 24860 14010 24912 14016
rect 24860 10736 24912 10742
rect 24860 10678 24912 10684
rect 24584 10600 24636 10606
rect 24584 10542 24636 10548
rect 24584 10464 24636 10470
rect 24584 10406 24636 10412
rect 24492 10056 24544 10062
rect 24492 9998 24544 10004
rect 24596 9722 24624 10406
rect 24584 9716 24636 9722
rect 24584 9658 24636 9664
rect 24872 9518 24900 10678
rect 24964 9625 24992 16934
rect 25044 14272 25096 14278
rect 25044 14214 25096 14220
rect 25056 13870 25084 14214
rect 25044 13864 25096 13870
rect 25044 13806 25096 13812
rect 25136 11348 25188 11354
rect 25136 11290 25188 11296
rect 25148 11218 25176 11290
rect 25136 11212 25188 11218
rect 25136 11154 25188 11160
rect 25044 10736 25096 10742
rect 25044 10678 25096 10684
rect 25056 10606 25084 10678
rect 25044 10600 25096 10606
rect 25044 10542 25096 10548
rect 24950 9616 25006 9625
rect 24950 9551 25006 9560
rect 24308 9512 24360 9518
rect 24308 9454 24360 9460
rect 24860 9512 24912 9518
rect 24860 9454 24912 9460
rect 24400 9036 24452 9042
rect 24400 8978 24452 8984
rect 24676 9036 24728 9042
rect 24676 8978 24728 8984
rect 24032 8560 24084 8566
rect 24032 8502 24084 8508
rect 23940 8424 23992 8430
rect 23940 8366 23992 8372
rect 24044 8090 24072 8502
rect 23756 8084 23808 8090
rect 23756 8026 23808 8032
rect 24032 8084 24084 8090
rect 24032 8026 24084 8032
rect 23480 7958 23532 7964
rect 23662 7984 23718 7993
rect 23492 6866 23520 7958
rect 23662 7919 23718 7928
rect 23676 7410 23704 7919
rect 23664 7404 23716 7410
rect 23664 7346 23716 7352
rect 23480 6860 23532 6866
rect 23480 6802 23532 6808
rect 23676 6458 23704 7346
rect 23768 6866 23796 8026
rect 23940 7948 23992 7954
rect 23940 7890 23992 7896
rect 23848 7744 23900 7750
rect 23848 7686 23900 7692
rect 23860 7546 23888 7686
rect 23952 7546 23980 7890
rect 24412 7750 24440 8978
rect 24688 8566 24716 8978
rect 24952 8900 25004 8906
rect 24952 8842 25004 8848
rect 24676 8560 24728 8566
rect 24676 8502 24728 8508
rect 24964 8498 24992 8842
rect 24952 8492 25004 8498
rect 24952 8434 25004 8440
rect 24676 7880 24728 7886
rect 24676 7822 24728 7828
rect 24400 7744 24452 7750
rect 24400 7686 24452 7692
rect 23848 7540 23900 7546
rect 23848 7482 23900 7488
rect 23940 7540 23992 7546
rect 23940 7482 23992 7488
rect 24216 7336 24268 7342
rect 24216 7278 24268 7284
rect 24228 6934 24256 7278
rect 24216 6928 24268 6934
rect 24216 6870 24268 6876
rect 24492 6928 24544 6934
rect 24492 6870 24544 6876
rect 23756 6860 23808 6866
rect 23756 6802 23808 6808
rect 23388 6452 23440 6458
rect 23388 6394 23440 6400
rect 23664 6452 23716 6458
rect 23664 6394 23716 6400
rect 24400 6248 24452 6254
rect 24400 6190 24452 6196
rect 24412 5642 24440 6190
rect 24400 5636 24452 5642
rect 24400 5578 24452 5584
rect 23296 5568 23348 5574
rect 23296 5510 23348 5516
rect 23112 5092 23164 5098
rect 23112 5034 23164 5040
rect 23124 4758 23152 5034
rect 23112 4752 23164 4758
rect 23112 4694 23164 4700
rect 24412 4690 24440 5578
rect 24504 5370 24532 6870
rect 24584 6860 24636 6866
rect 24584 6802 24636 6808
rect 24596 6322 24624 6802
rect 24688 6730 24716 7822
rect 24768 6860 24820 6866
rect 24768 6802 24820 6808
rect 24676 6724 24728 6730
rect 24676 6666 24728 6672
rect 24688 6390 24716 6666
rect 24780 6662 24808 6802
rect 25056 6662 25084 10542
rect 24768 6656 24820 6662
rect 24768 6598 24820 6604
rect 25044 6656 25096 6662
rect 25044 6598 25096 6604
rect 24676 6384 24728 6390
rect 24676 6326 24728 6332
rect 24780 6338 24808 6598
rect 24584 6316 24636 6322
rect 24780 6310 24900 6338
rect 25056 6322 25084 6598
rect 24584 6258 24636 6264
rect 24596 5914 24624 6258
rect 24768 6248 24820 6254
rect 24768 6190 24820 6196
rect 24584 5908 24636 5914
rect 24584 5850 24636 5856
rect 24492 5364 24544 5370
rect 24492 5306 24544 5312
rect 24504 4690 24532 5306
rect 24780 4690 24808 6190
rect 24872 5778 24900 6310
rect 25044 6316 25096 6322
rect 25044 6258 25096 6264
rect 25056 6118 25084 6258
rect 25044 6112 25096 6118
rect 25044 6054 25096 6060
rect 24860 5772 24912 5778
rect 24860 5714 24912 5720
rect 25044 5704 25096 5710
rect 25044 5646 25096 5652
rect 24400 4684 24452 4690
rect 24400 4626 24452 4632
rect 24492 4684 24544 4690
rect 24492 4626 24544 4632
rect 24768 4684 24820 4690
rect 24768 4626 24820 4632
rect 23848 4616 23900 4622
rect 23848 4558 23900 4564
rect 23860 4146 23888 4558
rect 24860 4208 24912 4214
rect 24860 4150 24912 4156
rect 23848 4140 23900 4146
rect 23848 4082 23900 4088
rect 24872 4078 24900 4150
rect 25056 4146 25084 5646
rect 25240 5250 25268 24806
rect 25332 22234 25360 26386
rect 25412 25832 25464 25838
rect 25412 25774 25464 25780
rect 25424 23186 25452 25774
rect 25516 25158 25544 28070
rect 25780 28008 25832 28014
rect 25780 27950 25832 27956
rect 25688 27872 25740 27878
rect 25688 27814 25740 27820
rect 25700 27674 25728 27814
rect 25688 27668 25740 27674
rect 25688 27610 25740 27616
rect 25596 27532 25648 27538
rect 25596 27474 25648 27480
rect 25608 26586 25636 27474
rect 25596 26580 25648 26586
rect 25596 26522 25648 26528
rect 25608 26042 25636 26522
rect 25792 26450 25820 27950
rect 25884 27878 25912 35158
rect 25964 35080 26016 35086
rect 25964 35022 26016 35028
rect 25976 34610 26004 35022
rect 25964 34604 26016 34610
rect 25964 34546 26016 34552
rect 26252 34474 26280 35702
rect 26344 34542 26372 35770
rect 26332 34536 26384 34542
rect 26332 34478 26384 34484
rect 26240 34468 26292 34474
rect 26240 34410 26292 34416
rect 26252 33522 26280 34410
rect 26344 34066 26372 34478
rect 26332 34060 26384 34066
rect 26332 34002 26384 34008
rect 26240 33516 26292 33522
rect 26240 33458 26292 33464
rect 26344 32910 26372 34002
rect 26332 32904 26384 32910
rect 26332 32846 26384 32852
rect 26056 32292 26108 32298
rect 26056 32234 26108 32240
rect 26068 30190 26096 32234
rect 26332 31884 26384 31890
rect 26332 31826 26384 31832
rect 26148 31816 26200 31822
rect 26148 31758 26200 31764
rect 26160 30870 26188 31758
rect 26344 31414 26372 31826
rect 26332 31408 26384 31414
rect 26332 31350 26384 31356
rect 26148 30864 26200 30870
rect 26148 30806 26200 30812
rect 26344 30258 26372 31350
rect 26332 30252 26384 30258
rect 26332 30194 26384 30200
rect 26056 30184 26108 30190
rect 25976 30144 26056 30172
rect 25976 29102 26004 30144
rect 26056 30126 26108 30132
rect 26344 29306 26372 30194
rect 26436 30190 26464 36518
rect 26620 36242 26648 37266
rect 27448 36650 27476 38286
rect 27620 38208 27672 38214
rect 27620 38150 27672 38156
rect 27528 37664 27580 37670
rect 27528 37606 27580 37612
rect 27436 36644 27488 36650
rect 27436 36586 27488 36592
rect 26608 36236 26660 36242
rect 26608 36178 26660 36184
rect 27252 36100 27304 36106
rect 27252 36042 27304 36048
rect 27264 35834 27292 36042
rect 27252 35828 27304 35834
rect 27252 35770 27304 35776
rect 27448 35290 27476 36586
rect 27436 35284 27488 35290
rect 27436 35226 27488 35232
rect 26608 35148 26660 35154
rect 26608 35090 26660 35096
rect 26620 34134 26648 35090
rect 27448 35086 27476 35226
rect 27436 35080 27488 35086
rect 27436 35022 27488 35028
rect 26792 34944 26844 34950
rect 26792 34886 26844 34892
rect 26608 34128 26660 34134
rect 26608 34070 26660 34076
rect 26804 34066 26832 34886
rect 26792 34060 26844 34066
rect 26792 34002 26844 34008
rect 26700 33856 26752 33862
rect 26700 33798 26752 33804
rect 26712 31278 26740 33798
rect 27160 33448 27212 33454
rect 27160 33390 27212 33396
rect 27344 33448 27396 33454
rect 27344 33390 27396 33396
rect 26792 33380 26844 33386
rect 26792 33322 26844 33328
rect 26804 32502 26832 33322
rect 27172 32978 27200 33390
rect 27160 32972 27212 32978
rect 27160 32914 27212 32920
rect 26792 32496 26844 32502
rect 26792 32438 26844 32444
rect 27172 32366 27200 32914
rect 27356 32366 27384 33390
rect 27160 32360 27212 32366
rect 27160 32302 27212 32308
rect 27344 32360 27396 32366
rect 27344 32302 27396 32308
rect 27172 31278 27200 32302
rect 27356 32230 27384 32302
rect 27344 32224 27396 32230
rect 27344 32166 27396 32172
rect 27252 31680 27304 31686
rect 27356 31668 27384 32166
rect 27540 31890 27568 37606
rect 27632 37330 27660 38150
rect 27816 38010 27844 40200
rect 29840 38434 29868 40200
rect 29840 38418 29960 38434
rect 29840 38412 29972 38418
rect 29840 38406 29920 38412
rect 29920 38354 29972 38360
rect 28632 38344 28684 38350
rect 28632 38286 28684 38292
rect 27804 38004 27856 38010
rect 27804 37946 27856 37952
rect 28080 37800 28132 37806
rect 28080 37742 28132 37748
rect 27620 37324 27672 37330
rect 27620 37266 27672 37272
rect 27988 37120 28040 37126
rect 28092 37074 28120 37742
rect 28040 37068 28120 37074
rect 27988 37062 28120 37068
rect 28000 37046 28120 37062
rect 27804 36916 27856 36922
rect 27804 36858 27856 36864
rect 27816 36242 27844 36858
rect 27804 36236 27856 36242
rect 27804 36178 27856 36184
rect 27804 36032 27856 36038
rect 27804 35974 27856 35980
rect 27620 35624 27672 35630
rect 27620 35566 27672 35572
rect 27632 35154 27660 35566
rect 27620 35148 27672 35154
rect 27620 35090 27672 35096
rect 27816 33454 27844 35974
rect 27804 33448 27856 33454
rect 27804 33390 27856 33396
rect 27896 33448 27948 33454
rect 27896 33390 27948 33396
rect 27712 32904 27764 32910
rect 27712 32846 27764 32852
rect 27528 31884 27580 31890
rect 27528 31826 27580 31832
rect 27724 31686 27752 32846
rect 27908 32366 27936 33390
rect 27896 32360 27948 32366
rect 27896 32302 27948 32308
rect 27908 31822 27936 32302
rect 27896 31816 27948 31822
rect 27896 31758 27948 31764
rect 27304 31640 27384 31668
rect 27712 31680 27764 31686
rect 27252 31622 27304 31628
rect 27712 31622 27764 31628
rect 27264 31278 27292 31622
rect 26516 31272 26568 31278
rect 26516 31214 26568 31220
rect 26700 31272 26752 31278
rect 26700 31214 26752 31220
rect 27160 31272 27212 31278
rect 27160 31214 27212 31220
rect 27252 31272 27304 31278
rect 27252 31214 27304 31220
rect 26424 30184 26476 30190
rect 26424 30126 26476 30132
rect 26528 29510 26556 31214
rect 27988 31136 28040 31142
rect 27988 31078 28040 31084
rect 27068 30796 27120 30802
rect 27068 30738 27120 30744
rect 27080 30705 27108 30738
rect 27620 30728 27672 30734
rect 27066 30696 27122 30705
rect 27620 30670 27672 30676
rect 27066 30631 27122 30640
rect 27252 30660 27304 30666
rect 27252 30602 27304 30608
rect 27160 30048 27212 30054
rect 27264 30002 27292 30602
rect 27212 29996 27292 30002
rect 27160 29990 27292 29996
rect 27172 29974 27292 29990
rect 26608 29708 26660 29714
rect 26608 29650 26660 29656
rect 26516 29504 26568 29510
rect 26516 29446 26568 29452
rect 26332 29300 26384 29306
rect 26332 29242 26384 29248
rect 25964 29096 26016 29102
rect 25964 29038 26016 29044
rect 26056 29096 26108 29102
rect 26108 29056 26280 29084
rect 26056 29038 26108 29044
rect 26252 29050 26280 29056
rect 26252 29022 26464 29050
rect 25964 28960 26016 28966
rect 25964 28902 26016 28908
rect 26240 28960 26292 28966
rect 26240 28902 26292 28908
rect 25976 28014 26004 28902
rect 26252 28558 26280 28902
rect 26332 28620 26384 28626
rect 26332 28562 26384 28568
rect 26240 28552 26292 28558
rect 26240 28494 26292 28500
rect 25964 28008 26016 28014
rect 25964 27950 26016 27956
rect 25872 27872 25924 27878
rect 25872 27814 25924 27820
rect 25976 26994 26004 27950
rect 25964 26988 26016 26994
rect 25964 26930 26016 26936
rect 25780 26444 25832 26450
rect 25780 26386 25832 26392
rect 25596 26036 25648 26042
rect 25596 25978 25648 25984
rect 25504 25152 25556 25158
rect 25504 25094 25556 25100
rect 25792 24818 25820 26386
rect 25964 25832 26016 25838
rect 25964 25774 26016 25780
rect 25872 25288 25924 25294
rect 25872 25230 25924 25236
rect 25780 24812 25832 24818
rect 25780 24754 25832 24760
rect 25596 24336 25648 24342
rect 25596 24278 25648 24284
rect 25412 23180 25464 23186
rect 25412 23122 25464 23128
rect 25424 22642 25452 23122
rect 25412 22636 25464 22642
rect 25412 22578 25464 22584
rect 25320 22228 25372 22234
rect 25320 22170 25372 22176
rect 25504 22092 25556 22098
rect 25504 22034 25556 22040
rect 25516 19922 25544 22034
rect 25608 21010 25636 24278
rect 25792 23662 25820 24754
rect 25780 23656 25832 23662
rect 25780 23598 25832 23604
rect 25688 22092 25740 22098
rect 25688 22034 25740 22040
rect 25700 21690 25728 22034
rect 25688 21684 25740 21690
rect 25688 21626 25740 21632
rect 25780 21684 25832 21690
rect 25780 21626 25832 21632
rect 25700 21078 25728 21626
rect 25792 21350 25820 21626
rect 25780 21344 25832 21350
rect 25780 21286 25832 21292
rect 25688 21072 25740 21078
rect 25688 21014 25740 21020
rect 25596 21004 25648 21010
rect 25596 20946 25648 20952
rect 25700 20398 25728 21014
rect 25688 20392 25740 20398
rect 25688 20334 25740 20340
rect 25504 19916 25556 19922
rect 25504 19858 25556 19864
rect 25884 19378 25912 25230
rect 25976 24342 26004 25774
rect 25964 24336 26016 24342
rect 25964 24278 26016 24284
rect 26240 23656 26292 23662
rect 26240 23598 26292 23604
rect 26252 23322 26280 23598
rect 26240 23316 26292 23322
rect 26240 23258 26292 23264
rect 26148 21480 26200 21486
rect 26148 21422 26200 21428
rect 25964 20936 26016 20942
rect 25964 20878 26016 20884
rect 25976 20058 26004 20878
rect 26160 20874 26188 21422
rect 26240 21344 26292 21350
rect 26240 21286 26292 21292
rect 26148 20868 26200 20874
rect 26148 20810 26200 20816
rect 26252 20466 26280 21286
rect 26240 20460 26292 20466
rect 26240 20402 26292 20408
rect 25964 20052 26016 20058
rect 25964 19994 26016 20000
rect 25872 19372 25924 19378
rect 25872 19314 25924 19320
rect 25502 19000 25558 19009
rect 25502 18935 25558 18944
rect 25516 18834 25544 18935
rect 25504 18828 25556 18834
rect 25504 18770 25556 18776
rect 25688 18828 25740 18834
rect 25688 18770 25740 18776
rect 25318 18592 25374 18601
rect 25318 18527 25374 18536
rect 25332 10742 25360 18527
rect 25700 18358 25728 18770
rect 26240 18760 26292 18766
rect 26240 18702 26292 18708
rect 25688 18352 25740 18358
rect 25688 18294 25740 18300
rect 25872 18284 25924 18290
rect 25872 18226 25924 18232
rect 25884 17882 25912 18226
rect 25872 17876 25924 17882
rect 25872 17818 25924 17824
rect 26252 17814 26280 18702
rect 26240 17808 26292 17814
rect 26240 17750 26292 17756
rect 25412 17536 25464 17542
rect 25412 17478 25464 17484
rect 25320 10736 25372 10742
rect 25320 10678 25372 10684
rect 25320 9512 25372 9518
rect 25424 9489 25452 17478
rect 26148 17332 26200 17338
rect 26148 17274 26200 17280
rect 26160 17202 26188 17274
rect 26148 17196 26200 17202
rect 26148 17138 26200 17144
rect 26160 15502 26188 17138
rect 26344 16946 26372 28562
rect 26436 28014 26464 29022
rect 26528 28762 26556 29446
rect 26620 29102 26648 29650
rect 27264 29646 27292 29974
rect 27632 29714 27660 30670
rect 27712 30048 27764 30054
rect 27712 29990 27764 29996
rect 27620 29708 27672 29714
rect 27620 29650 27672 29656
rect 26700 29640 26752 29646
rect 26700 29582 26752 29588
rect 27252 29640 27304 29646
rect 27252 29582 27304 29588
rect 26608 29096 26660 29102
rect 26608 29038 26660 29044
rect 26516 28756 26568 28762
rect 26516 28698 26568 28704
rect 26620 28642 26648 29038
rect 26528 28614 26648 28642
rect 26424 28008 26476 28014
rect 26424 27950 26476 27956
rect 26528 27946 26556 28614
rect 26712 28558 26740 29582
rect 26976 29164 27028 29170
rect 26976 29106 27028 29112
rect 26608 28552 26660 28558
rect 26608 28494 26660 28500
rect 26700 28552 26752 28558
rect 26700 28494 26752 28500
rect 26620 28422 26648 28494
rect 26608 28416 26660 28422
rect 26608 28358 26660 28364
rect 26884 28008 26936 28014
rect 26884 27950 26936 27956
rect 26516 27940 26568 27946
rect 26516 27882 26568 27888
rect 26896 26926 26924 27950
rect 26988 27334 27016 29106
rect 27068 27940 27120 27946
rect 27068 27882 27120 27888
rect 27080 27606 27108 27882
rect 27068 27600 27120 27606
rect 27068 27542 27120 27548
rect 26976 27328 27028 27334
rect 26976 27270 27028 27276
rect 26884 26920 26936 26926
rect 26884 26862 26936 26868
rect 26896 26518 26924 26862
rect 26884 26512 26936 26518
rect 26884 26454 26936 26460
rect 26608 26308 26660 26314
rect 26608 26250 26660 26256
rect 26620 25362 26648 26250
rect 26896 25702 26924 26454
rect 26988 25906 27016 27270
rect 27264 26382 27292 29582
rect 27618 29064 27674 29073
rect 27618 28999 27674 29008
rect 27632 28694 27660 28999
rect 27620 28688 27672 28694
rect 27620 28630 27672 28636
rect 27724 28626 27752 29990
rect 27804 29504 27856 29510
rect 27804 29446 27856 29452
rect 27816 29102 27844 29446
rect 27804 29096 27856 29102
rect 27804 29038 27856 29044
rect 27712 28620 27764 28626
rect 27712 28562 27764 28568
rect 27526 28520 27582 28529
rect 27816 28506 27844 29038
rect 27526 28455 27582 28464
rect 27724 28478 27844 28506
rect 27540 28422 27568 28455
rect 27436 28416 27488 28422
rect 27436 28358 27488 28364
rect 27528 28416 27580 28422
rect 27528 28358 27580 28364
rect 27252 26376 27304 26382
rect 27252 26318 27304 26324
rect 26976 25900 27028 25906
rect 26976 25842 27028 25848
rect 27252 25832 27304 25838
rect 27252 25774 27304 25780
rect 26884 25696 26936 25702
rect 26884 25638 26936 25644
rect 27264 25362 27292 25774
rect 26608 25356 26660 25362
rect 26608 25298 26660 25304
rect 27252 25356 27304 25362
rect 27252 25298 27304 25304
rect 27264 24818 27292 25298
rect 26516 24812 26568 24818
rect 26516 24754 26568 24760
rect 27252 24812 27304 24818
rect 27252 24754 27304 24760
rect 26528 24274 26556 24754
rect 26884 24676 26936 24682
rect 26884 24618 26936 24624
rect 26516 24268 26568 24274
rect 26516 24210 26568 24216
rect 26424 23180 26476 23186
rect 26424 23122 26476 23128
rect 26436 22574 26464 23122
rect 26424 22568 26476 22574
rect 26422 22536 26424 22545
rect 26476 22536 26478 22545
rect 26422 22471 26478 22480
rect 26424 21412 26476 21418
rect 26424 21354 26476 21360
rect 26436 20398 26464 21354
rect 26528 21146 26556 24210
rect 26896 23746 26924 24618
rect 27448 24614 27476 28358
rect 27528 27940 27580 27946
rect 27528 27882 27580 27888
rect 27540 27674 27568 27882
rect 27528 27668 27580 27674
rect 27528 27610 27580 27616
rect 27620 26376 27672 26382
rect 27620 26318 27672 26324
rect 27436 24608 27488 24614
rect 27436 24550 27488 24556
rect 27160 24200 27212 24206
rect 27160 24142 27212 24148
rect 26712 23718 26924 23746
rect 26712 23662 26740 23718
rect 26700 23656 26752 23662
rect 26700 23598 26752 23604
rect 26884 23656 26936 23662
rect 26884 23598 26936 23604
rect 26712 22778 26740 23598
rect 26700 22772 26752 22778
rect 26700 22714 26752 22720
rect 26792 22568 26844 22574
rect 26896 22545 26924 23598
rect 27068 23180 27120 23186
rect 27068 23122 27120 23128
rect 27080 22574 27108 23122
rect 27172 22574 27200 24142
rect 27344 23724 27396 23730
rect 27344 23666 27396 23672
rect 27252 23112 27304 23118
rect 27252 23054 27304 23060
rect 27264 22642 27292 23054
rect 27252 22636 27304 22642
rect 27252 22578 27304 22584
rect 27068 22568 27120 22574
rect 26792 22510 26844 22516
rect 26882 22536 26938 22545
rect 26804 22166 26832 22510
rect 27068 22510 27120 22516
rect 27160 22568 27212 22574
rect 27356 22522 27384 23666
rect 27448 23066 27476 24550
rect 27632 24410 27660 26318
rect 27724 26246 27752 28478
rect 27802 28112 27858 28121
rect 27802 28047 27804 28056
rect 27856 28047 27858 28056
rect 27804 28018 27856 28024
rect 27712 26240 27764 26246
rect 27712 26182 27764 26188
rect 27620 24404 27672 24410
rect 27620 24346 27672 24352
rect 27528 24132 27580 24138
rect 27528 24074 27580 24080
rect 27540 23186 27568 24074
rect 27724 23526 27752 26182
rect 28000 24954 28028 31078
rect 27988 24948 28040 24954
rect 27988 24890 28040 24896
rect 27896 24200 27948 24206
rect 27896 24142 27948 24148
rect 27908 23798 27936 24142
rect 27896 23792 27948 23798
rect 27896 23734 27948 23740
rect 27908 23662 27936 23734
rect 27896 23656 27948 23662
rect 27896 23598 27948 23604
rect 27712 23520 27764 23526
rect 27712 23462 27764 23468
rect 27620 23248 27672 23254
rect 27620 23190 27672 23196
rect 27528 23180 27580 23186
rect 27528 23122 27580 23128
rect 27448 23038 27568 23066
rect 27160 22510 27212 22516
rect 26882 22471 26938 22480
rect 26976 22500 27028 22506
rect 26976 22442 27028 22448
rect 26792 22160 26844 22166
rect 26792 22102 26844 22108
rect 26988 22098 27016 22442
rect 27080 22098 27108 22510
rect 27264 22494 27384 22522
rect 26976 22092 27028 22098
rect 26976 22034 27028 22040
rect 27068 22092 27120 22098
rect 27068 22034 27120 22040
rect 26792 21616 26844 21622
rect 26792 21558 26844 21564
rect 26516 21140 26568 21146
rect 26516 21082 26568 21088
rect 26804 21010 26832 21558
rect 26976 21480 27028 21486
rect 26976 21422 27028 21428
rect 26792 21004 26844 21010
rect 26792 20946 26844 20952
rect 26804 20466 26832 20946
rect 26792 20460 26844 20466
rect 26792 20402 26844 20408
rect 26424 20392 26476 20398
rect 26424 20334 26476 20340
rect 26608 19304 26660 19310
rect 26608 19246 26660 19252
rect 26424 18216 26476 18222
rect 26424 18158 26476 18164
rect 26436 16998 26464 18158
rect 26620 17542 26648 19246
rect 26792 19168 26844 19174
rect 26792 19110 26844 19116
rect 26804 18834 26832 19110
rect 26988 18834 27016 21422
rect 27080 20942 27108 22034
rect 27068 20936 27120 20942
rect 27068 20878 27120 20884
rect 27160 19236 27212 19242
rect 27160 19178 27212 19184
rect 27068 19168 27120 19174
rect 27068 19110 27120 19116
rect 26792 18828 26844 18834
rect 26792 18770 26844 18776
rect 26976 18828 27028 18834
rect 26976 18770 27028 18776
rect 26804 18426 26832 18770
rect 27080 18698 27108 19110
rect 27172 18834 27200 19178
rect 27160 18828 27212 18834
rect 27160 18770 27212 18776
rect 27172 18737 27200 18770
rect 27158 18728 27214 18737
rect 27068 18692 27120 18698
rect 27158 18663 27214 18672
rect 27068 18634 27120 18640
rect 26792 18420 26844 18426
rect 26792 18362 26844 18368
rect 26804 18222 26832 18362
rect 27172 18222 27200 18663
rect 26792 18216 26844 18222
rect 26792 18158 26844 18164
rect 27160 18216 27212 18222
rect 27160 18158 27212 18164
rect 26884 18148 26936 18154
rect 26884 18090 26936 18096
rect 27068 18148 27120 18154
rect 27068 18090 27120 18096
rect 26896 17746 26924 18090
rect 27080 17814 27108 18090
rect 27068 17808 27120 17814
rect 27068 17750 27120 17756
rect 26884 17740 26936 17746
rect 26884 17682 26936 17688
rect 26608 17536 26660 17542
rect 26608 17478 26660 17484
rect 26252 16918 26372 16946
rect 26424 16992 26476 16998
rect 26424 16934 26476 16940
rect 26792 16992 26844 16998
rect 26792 16934 26844 16940
rect 26148 15496 26200 15502
rect 26148 15438 26200 15444
rect 26160 14414 26188 15438
rect 26148 14408 26200 14414
rect 26148 14350 26200 14356
rect 26160 14074 26188 14350
rect 26148 14068 26200 14074
rect 26148 14010 26200 14016
rect 25780 12776 25832 12782
rect 25780 12718 25832 12724
rect 25792 12374 25820 12718
rect 25780 12368 25832 12374
rect 25780 12310 25832 12316
rect 25504 11552 25556 11558
rect 25504 11494 25556 11500
rect 25516 10849 25544 11494
rect 25688 11212 25740 11218
rect 25688 11154 25740 11160
rect 25502 10840 25558 10849
rect 25502 10775 25558 10784
rect 25320 9454 25372 9460
rect 25410 9480 25466 9489
rect 25332 9110 25360 9454
rect 25410 9415 25466 9424
rect 25320 9104 25372 9110
rect 25320 9046 25372 9052
rect 25332 7954 25360 9046
rect 25424 8974 25452 9415
rect 25412 8968 25464 8974
rect 25412 8910 25464 8916
rect 25516 8514 25544 10775
rect 25700 10520 25728 11154
rect 26252 10810 26280 16918
rect 26804 16794 26832 16934
rect 26792 16788 26844 16794
rect 26792 16730 26844 16736
rect 26804 16658 26832 16730
rect 26608 16652 26660 16658
rect 26608 16594 26660 16600
rect 26792 16652 26844 16658
rect 26792 16594 26844 16600
rect 26516 15972 26568 15978
rect 26516 15914 26568 15920
rect 26528 15026 26556 15914
rect 26620 15570 26648 16594
rect 26608 15564 26660 15570
rect 26608 15506 26660 15512
rect 26516 15020 26568 15026
rect 26516 14962 26568 14968
rect 26608 14816 26660 14822
rect 26608 14758 26660 14764
rect 26620 14482 26648 14758
rect 26608 14476 26660 14482
rect 26608 14418 26660 14424
rect 26804 14362 26832 16594
rect 26884 16584 26936 16590
rect 26884 16526 26936 16532
rect 26896 16114 26924 16526
rect 26884 16108 26936 16114
rect 26884 16050 26936 16056
rect 26804 14334 27016 14362
rect 26792 14272 26844 14278
rect 26792 14214 26844 14220
rect 26884 14272 26936 14278
rect 26884 14214 26936 14220
rect 26424 13524 26476 13530
rect 26424 13466 26476 13472
rect 26436 11218 26464 13466
rect 26804 12442 26832 14214
rect 26896 13870 26924 14214
rect 26884 13864 26936 13870
rect 26884 13806 26936 13812
rect 26988 13462 27016 14334
rect 26976 13456 27028 13462
rect 26976 13398 27028 13404
rect 26792 12436 26844 12442
rect 26792 12378 26844 12384
rect 27080 12322 27108 17750
rect 27172 17746 27200 18158
rect 27160 17740 27212 17746
rect 27160 17682 27212 17688
rect 27264 17202 27292 22494
rect 27540 22386 27568 23038
rect 27632 22438 27660 23190
rect 27908 22438 27936 23598
rect 27356 22358 27568 22386
rect 27620 22432 27672 22438
rect 27620 22374 27672 22380
rect 27896 22432 27948 22438
rect 27896 22374 27948 22380
rect 27252 17196 27304 17202
rect 27252 17138 27304 17144
rect 27264 16658 27292 17138
rect 27356 16726 27384 22358
rect 27528 22228 27580 22234
rect 27528 22170 27580 22176
rect 27436 18828 27488 18834
rect 27436 18770 27488 18776
rect 27448 18601 27476 18770
rect 27434 18592 27490 18601
rect 27434 18527 27490 18536
rect 27436 18420 27488 18426
rect 27436 18362 27488 18368
rect 27448 17746 27476 18362
rect 27436 17740 27488 17746
rect 27436 17682 27488 17688
rect 27344 16720 27396 16726
rect 27344 16662 27396 16668
rect 27252 16652 27304 16658
rect 27252 16594 27304 16600
rect 27160 15360 27212 15366
rect 27160 15302 27212 15308
rect 27172 13870 27200 15302
rect 27252 14000 27304 14006
rect 27252 13942 27304 13948
rect 27160 13864 27212 13870
rect 27160 13806 27212 13812
rect 27264 13802 27292 13942
rect 27252 13796 27304 13802
rect 27252 13738 27304 13744
rect 27356 13462 27384 16662
rect 27436 13864 27488 13870
rect 27436 13806 27488 13812
rect 27344 13456 27396 13462
rect 27344 13398 27396 13404
rect 27356 12850 27384 13398
rect 27344 12844 27396 12850
rect 27344 12786 27396 12792
rect 27344 12708 27396 12714
rect 27344 12650 27396 12656
rect 26804 12294 27108 12322
rect 26424 11212 26476 11218
rect 26424 11154 26476 11160
rect 26608 11212 26660 11218
rect 26608 11154 26660 11160
rect 26436 10810 26464 11154
rect 26240 10804 26292 10810
rect 26240 10746 26292 10752
rect 26424 10804 26476 10810
rect 26424 10746 26476 10752
rect 26148 10736 26200 10742
rect 26148 10678 26200 10684
rect 25780 10532 25832 10538
rect 25700 10492 25780 10520
rect 25700 10266 25728 10492
rect 25780 10474 25832 10480
rect 25964 10464 26016 10470
rect 25964 10406 26016 10412
rect 25688 10260 25740 10266
rect 25688 10202 25740 10208
rect 25688 9920 25740 9926
rect 25688 9862 25740 9868
rect 25700 9586 25728 9862
rect 25976 9586 26004 10406
rect 25688 9580 25740 9586
rect 25688 9522 25740 9528
rect 25964 9580 26016 9586
rect 25964 9522 26016 9528
rect 26160 9178 26188 10678
rect 26620 10606 26648 11154
rect 26608 10600 26660 10606
rect 26608 10542 26660 10548
rect 26620 9178 26648 10542
rect 26148 9172 26200 9178
rect 26148 9114 26200 9120
rect 26608 9172 26660 9178
rect 26608 9114 26660 9120
rect 25516 8498 25636 8514
rect 25516 8492 25648 8498
rect 25516 8486 25596 8492
rect 25516 7954 25544 8486
rect 25596 8434 25648 8440
rect 25320 7948 25372 7954
rect 25320 7890 25372 7896
rect 25504 7948 25556 7954
rect 25504 7890 25556 7896
rect 25332 6798 25360 7890
rect 25780 7880 25832 7886
rect 25780 7822 25832 7828
rect 26238 7848 26294 7857
rect 25320 6792 25372 6798
rect 25320 6734 25372 6740
rect 25792 6322 25820 7822
rect 26238 7783 26294 7792
rect 26252 7546 26280 7783
rect 26240 7540 26292 7546
rect 26240 7482 26292 7488
rect 26700 7336 26752 7342
rect 26700 7278 26752 7284
rect 26240 6656 26292 6662
rect 26240 6598 26292 6604
rect 25780 6316 25832 6322
rect 25780 6258 25832 6264
rect 25596 6248 25648 6254
rect 25596 6190 25648 6196
rect 25412 6180 25464 6186
rect 25412 6122 25464 6128
rect 25148 5222 25268 5250
rect 25044 4140 25096 4146
rect 25044 4082 25096 4088
rect 23480 4072 23532 4078
rect 23480 4014 23532 4020
rect 24492 4072 24544 4078
rect 24492 4014 24544 4020
rect 24860 4072 24912 4078
rect 24860 4014 24912 4020
rect 22928 3596 22980 3602
rect 22928 3538 22980 3544
rect 23020 3596 23072 3602
rect 23072 3556 23152 3584
rect 23020 3538 23072 3544
rect 22560 3392 22612 3398
rect 22560 3334 22612 3340
rect 22652 3392 22704 3398
rect 22652 3334 22704 3340
rect 22572 2990 22600 3334
rect 22100 2984 22152 2990
rect 22100 2926 22152 2932
rect 22560 2984 22612 2990
rect 22560 2926 22612 2932
rect 22664 2514 22692 3334
rect 22940 3126 22968 3538
rect 22928 3120 22980 3126
rect 22928 3062 22980 3068
rect 23124 2990 23152 3556
rect 23204 3528 23256 3534
rect 23204 3470 23256 3476
rect 23112 2984 23164 2990
rect 23112 2926 23164 2932
rect 22744 2916 22796 2922
rect 22744 2858 22796 2864
rect 23020 2916 23072 2922
rect 23020 2858 23072 2864
rect 22756 2514 22784 2858
rect 22652 2508 22704 2514
rect 22652 2450 22704 2456
rect 22744 2508 22796 2514
rect 22744 2450 22796 2456
rect 23032 2310 23060 2858
rect 23216 2582 23244 3470
rect 23492 2854 23520 4014
rect 23572 3732 23624 3738
rect 23572 3674 23624 3680
rect 23388 2848 23440 2854
rect 23388 2790 23440 2796
rect 23480 2848 23532 2854
rect 23480 2790 23532 2796
rect 23400 2582 23428 2790
rect 23204 2576 23256 2582
rect 23204 2518 23256 2524
rect 23388 2576 23440 2582
rect 23388 2518 23440 2524
rect 23492 2514 23520 2790
rect 23480 2508 23532 2514
rect 23480 2450 23532 2456
rect 23020 2304 23072 2310
rect 23020 2246 23072 2252
rect 23584 800 23612 3674
rect 24504 3670 24532 4014
rect 25148 3738 25176 5222
rect 25228 5160 25280 5166
rect 25228 5102 25280 5108
rect 25136 3732 25188 3738
rect 25136 3674 25188 3680
rect 24492 3664 24544 3670
rect 24492 3606 24544 3612
rect 24584 3528 24636 3534
rect 24584 3470 24636 3476
rect 24400 3392 24452 3398
rect 24400 3334 24452 3340
rect 24412 2650 24440 3334
rect 24596 3058 24624 3470
rect 25240 3194 25268 5102
rect 25424 4146 25452 6122
rect 25504 5160 25556 5166
rect 25504 5102 25556 5108
rect 25516 4214 25544 5102
rect 25608 5098 25636 6190
rect 25792 5166 25820 6258
rect 26252 6254 26280 6598
rect 26712 6458 26740 7278
rect 26804 6934 26832 12294
rect 26884 11892 26936 11898
rect 26884 11834 26936 11840
rect 26896 11234 26924 11834
rect 27356 11694 27384 12650
rect 27344 11688 27396 11694
rect 27344 11630 27396 11636
rect 26896 11218 27384 11234
rect 26896 11212 27396 11218
rect 26896 11206 27344 11212
rect 26896 9654 26924 11206
rect 27344 11154 27396 11160
rect 26976 11076 27028 11082
rect 26976 11018 27028 11024
rect 26988 10606 27016 11018
rect 27160 10804 27212 10810
rect 27160 10746 27212 10752
rect 27172 10674 27200 10746
rect 27160 10668 27212 10674
rect 27160 10610 27212 10616
rect 26976 10600 27028 10606
rect 26976 10542 27028 10548
rect 26988 10266 27016 10542
rect 26976 10260 27028 10266
rect 26976 10202 27028 10208
rect 27160 10056 27212 10062
rect 27160 9998 27212 10004
rect 26884 9648 26936 9654
rect 26884 9590 26936 9596
rect 26896 9042 26924 9590
rect 27172 9110 27200 9998
rect 27344 9512 27396 9518
rect 27344 9454 27396 9460
rect 27356 9110 27384 9454
rect 27160 9104 27212 9110
rect 27160 9046 27212 9052
rect 27344 9104 27396 9110
rect 27344 9046 27396 9052
rect 26884 9036 26936 9042
rect 26884 8978 26936 8984
rect 27448 7478 27476 13806
rect 27540 13394 27568 22170
rect 27632 22166 27660 22374
rect 27620 22160 27672 22166
rect 27620 22102 27672 22108
rect 27712 22092 27764 22098
rect 27712 22034 27764 22040
rect 27724 21486 27752 22034
rect 27712 21480 27764 21486
rect 27712 21422 27764 21428
rect 27620 21344 27672 21350
rect 27620 21286 27672 21292
rect 27632 21010 27660 21286
rect 27908 21026 27936 22374
rect 27988 21412 28040 21418
rect 27988 21354 28040 21360
rect 27620 21004 27672 21010
rect 27620 20946 27672 20952
rect 27816 20998 27936 21026
rect 27632 19922 27660 20946
rect 27712 20936 27764 20942
rect 27712 20878 27764 20884
rect 27724 20262 27752 20878
rect 27712 20256 27764 20262
rect 27712 20198 27764 20204
rect 27724 19990 27752 20198
rect 27712 19984 27764 19990
rect 27712 19926 27764 19932
rect 27620 19916 27672 19922
rect 27620 19858 27672 19864
rect 27712 19304 27764 19310
rect 27712 19246 27764 19252
rect 27618 19136 27674 19145
rect 27618 19071 27674 19080
rect 27632 17134 27660 19071
rect 27724 18834 27752 19246
rect 27712 18828 27764 18834
rect 27712 18770 27764 18776
rect 27724 18630 27752 18770
rect 27712 18624 27764 18630
rect 27712 18566 27764 18572
rect 27724 18222 27752 18566
rect 27712 18216 27764 18222
rect 27712 18158 27764 18164
rect 27816 17202 27844 20998
rect 27896 20868 27948 20874
rect 27896 20810 27948 20816
rect 27908 19922 27936 20810
rect 27896 19916 27948 19922
rect 27896 19858 27948 19864
rect 28000 19854 28028 21354
rect 27988 19848 28040 19854
rect 27988 19790 28040 19796
rect 28092 18612 28120 37046
rect 28172 36712 28224 36718
rect 28172 36654 28224 36660
rect 28184 36174 28212 36654
rect 28172 36168 28224 36174
rect 28172 36110 28224 36116
rect 28184 35494 28212 36110
rect 28448 35624 28500 35630
rect 28448 35566 28500 35572
rect 28172 35488 28224 35494
rect 28172 35430 28224 35436
rect 28184 33522 28212 35430
rect 28460 34678 28488 35566
rect 28448 34672 28500 34678
rect 28448 34614 28500 34620
rect 28172 33516 28224 33522
rect 28172 33458 28224 33464
rect 28184 31890 28212 33458
rect 28460 33454 28488 34614
rect 28644 33658 28672 38286
rect 30012 38208 30064 38214
rect 30012 38150 30064 38156
rect 31024 38208 31076 38214
rect 31024 38150 31076 38156
rect 29000 37868 29052 37874
rect 29000 37810 29052 37816
rect 28724 37120 28776 37126
rect 28724 37062 28776 37068
rect 28736 35154 28764 37062
rect 29012 36718 29040 37810
rect 29828 37664 29880 37670
rect 29828 37606 29880 37612
rect 29840 37466 29868 37606
rect 29828 37460 29880 37466
rect 29828 37402 29880 37408
rect 29276 37324 29328 37330
rect 29276 37266 29328 37272
rect 29288 36786 29316 37266
rect 30024 36786 30052 38150
rect 30104 37800 30156 37806
rect 30104 37742 30156 37748
rect 30116 37466 30144 37742
rect 30104 37460 30156 37466
rect 30104 37402 30156 37408
rect 31036 37330 31064 38150
rect 31680 38010 31708 40200
rect 31668 38004 31720 38010
rect 31668 37946 31720 37952
rect 32036 37800 32088 37806
rect 32036 37742 32088 37748
rect 32772 37800 32824 37806
rect 32772 37742 32824 37748
rect 31024 37324 31076 37330
rect 31024 37266 31076 37272
rect 31944 37324 31996 37330
rect 31944 37266 31996 37272
rect 31852 37256 31904 37262
rect 31852 37198 31904 37204
rect 29276 36780 29328 36786
rect 30012 36780 30064 36786
rect 29328 36740 29408 36768
rect 29276 36722 29328 36728
rect 29000 36712 29052 36718
rect 29000 36654 29052 36660
rect 29380 35698 29408 36740
rect 30012 36722 30064 36728
rect 30656 36576 30708 36582
rect 30656 36518 30708 36524
rect 29368 35692 29420 35698
rect 29368 35634 29420 35640
rect 28724 35148 28776 35154
rect 28724 35090 28776 35096
rect 29380 35086 29408 35634
rect 30196 35624 30248 35630
rect 30196 35566 30248 35572
rect 29736 35488 29788 35494
rect 29736 35430 29788 35436
rect 29748 35154 29776 35430
rect 29736 35148 29788 35154
rect 29736 35090 29788 35096
rect 29276 35080 29328 35086
rect 29276 35022 29328 35028
rect 29368 35080 29420 35086
rect 29368 35022 29420 35028
rect 29288 34610 29316 35022
rect 30208 34746 30236 35566
rect 30288 35284 30340 35290
rect 30288 35226 30340 35232
rect 30196 34740 30248 34746
rect 30196 34682 30248 34688
rect 29276 34604 29328 34610
rect 29276 34546 29328 34552
rect 29828 34604 29880 34610
rect 29828 34546 29880 34552
rect 28724 34536 28776 34542
rect 28724 34478 28776 34484
rect 28632 33652 28684 33658
rect 28632 33594 28684 33600
rect 28448 33448 28500 33454
rect 28448 33390 28500 33396
rect 28172 31884 28224 31890
rect 28172 31826 28224 31832
rect 28644 31822 28672 33594
rect 28448 31816 28500 31822
rect 28448 31758 28500 31764
rect 28632 31816 28684 31822
rect 28632 31758 28684 31764
rect 28460 31142 28488 31758
rect 28448 31136 28500 31142
rect 28448 31078 28500 31084
rect 28460 30054 28488 31078
rect 28644 30802 28672 31758
rect 28632 30796 28684 30802
rect 28632 30738 28684 30744
rect 28540 30184 28592 30190
rect 28540 30126 28592 30132
rect 28448 30048 28500 30054
rect 28448 29990 28500 29996
rect 28172 29232 28224 29238
rect 28172 29174 28224 29180
rect 28184 29102 28212 29174
rect 28172 29096 28224 29102
rect 28172 29038 28224 29044
rect 28264 28620 28316 28626
rect 28264 28562 28316 28568
rect 28276 27606 28304 28562
rect 28264 27600 28316 27606
rect 28264 27542 28316 27548
rect 28356 26852 28408 26858
rect 28356 26794 28408 26800
rect 28368 26518 28396 26794
rect 28356 26512 28408 26518
rect 28356 26454 28408 26460
rect 28172 26444 28224 26450
rect 28172 26386 28224 26392
rect 28184 26246 28212 26386
rect 28172 26240 28224 26246
rect 28172 26182 28224 26188
rect 28184 25838 28212 26182
rect 28172 25832 28224 25838
rect 28172 25774 28224 25780
rect 28264 25832 28316 25838
rect 28264 25774 28316 25780
rect 28276 25430 28304 25774
rect 28264 25424 28316 25430
rect 28264 25366 28316 25372
rect 28172 25288 28224 25294
rect 28172 25230 28224 25236
rect 28184 23322 28212 25230
rect 28172 23316 28224 23322
rect 28172 23258 28224 23264
rect 28276 22574 28304 25366
rect 28356 25288 28408 25294
rect 28356 25230 28408 25236
rect 28368 24274 28396 25230
rect 28356 24268 28408 24274
rect 28356 24210 28408 24216
rect 28460 23662 28488 29990
rect 28552 29510 28580 30126
rect 28540 29504 28592 29510
rect 28540 29446 28592 29452
rect 28632 26920 28684 26926
rect 28632 26862 28684 26868
rect 28644 26586 28672 26862
rect 28632 26580 28684 26586
rect 28632 26522 28684 26528
rect 28540 24676 28592 24682
rect 28540 24618 28592 24624
rect 28552 24274 28580 24618
rect 28540 24268 28592 24274
rect 28540 24210 28592 24216
rect 28448 23656 28500 23662
rect 28448 23598 28500 23604
rect 28356 23588 28408 23594
rect 28356 23530 28408 23536
rect 28368 23186 28396 23530
rect 28448 23520 28500 23526
rect 28448 23462 28500 23468
rect 28356 23180 28408 23186
rect 28356 23122 28408 23128
rect 28356 23044 28408 23050
rect 28356 22986 28408 22992
rect 28264 22568 28316 22574
rect 28264 22510 28316 22516
rect 28172 22092 28224 22098
rect 28172 22034 28224 22040
rect 28184 21486 28212 22034
rect 28172 21480 28224 21486
rect 28172 21422 28224 21428
rect 28276 21146 28304 22510
rect 28264 21140 28316 21146
rect 28264 21082 28316 21088
rect 28262 18864 28318 18873
rect 28262 18799 28318 18808
rect 28276 18698 28304 18799
rect 28264 18692 28316 18698
rect 28264 18634 28316 18640
rect 28092 18584 28212 18612
rect 27804 17196 27856 17202
rect 27804 17138 27856 17144
rect 27620 17128 27672 17134
rect 27620 17070 27672 17076
rect 27816 16658 27844 17138
rect 27896 17060 27948 17066
rect 27896 17002 27948 17008
rect 27804 16652 27856 16658
rect 27804 16594 27856 16600
rect 27620 16040 27672 16046
rect 27620 15982 27672 15988
rect 27632 14414 27660 15982
rect 27908 14890 27936 17002
rect 28080 16040 28132 16046
rect 28080 15982 28132 15988
rect 27896 14884 27948 14890
rect 27896 14826 27948 14832
rect 27804 14612 27856 14618
rect 27804 14554 27856 14560
rect 27712 14476 27764 14482
rect 27712 14418 27764 14424
rect 27620 14408 27672 14414
rect 27620 14350 27672 14356
rect 27620 13932 27672 13938
rect 27620 13874 27672 13880
rect 27528 13388 27580 13394
rect 27528 13330 27580 13336
rect 27540 12850 27568 13330
rect 27528 12844 27580 12850
rect 27528 12786 27580 12792
rect 27528 12436 27580 12442
rect 27528 12378 27580 12384
rect 27436 7472 27488 7478
rect 27436 7414 27488 7420
rect 27252 7336 27304 7342
rect 27252 7278 27304 7284
rect 27160 7200 27212 7206
rect 27160 7142 27212 7148
rect 26792 6928 26844 6934
rect 26792 6870 26844 6876
rect 26700 6452 26752 6458
rect 26700 6394 26752 6400
rect 26240 6248 26292 6254
rect 26240 6190 26292 6196
rect 25780 5160 25832 5166
rect 25780 5102 25832 5108
rect 25596 5092 25648 5098
rect 25596 5034 25648 5040
rect 25504 4208 25556 4214
rect 25504 4150 25556 4156
rect 25412 4140 25464 4146
rect 25412 4082 25464 4088
rect 25596 3596 25648 3602
rect 25596 3538 25648 3544
rect 25228 3188 25280 3194
rect 25228 3130 25280 3136
rect 24584 3052 24636 3058
rect 24584 2994 24636 3000
rect 24400 2644 24452 2650
rect 24400 2586 24452 2592
rect 24584 2440 24636 2446
rect 24584 2382 24636 2388
rect 24596 2106 24624 2382
rect 24584 2100 24636 2106
rect 24584 2042 24636 2048
rect 25608 800 25636 3538
rect 25780 3188 25832 3194
rect 25780 3130 25832 3136
rect 25792 2446 25820 3130
rect 26252 2582 26280 6190
rect 27172 5778 27200 7142
rect 27264 6866 27292 7278
rect 27252 6860 27304 6866
rect 27252 6802 27304 6808
rect 27068 5772 27120 5778
rect 27068 5714 27120 5720
rect 27160 5772 27212 5778
rect 27160 5714 27212 5720
rect 26516 5704 26568 5710
rect 26516 5646 26568 5652
rect 26528 5234 26556 5646
rect 27080 5642 27108 5714
rect 27068 5636 27120 5642
rect 27068 5578 27120 5584
rect 26516 5228 26568 5234
rect 26516 5170 26568 5176
rect 26608 5160 26660 5166
rect 26608 5102 26660 5108
rect 26516 4616 26568 4622
rect 26516 4558 26568 4564
rect 26528 4146 26556 4558
rect 26516 4140 26568 4146
rect 26516 4082 26568 4088
rect 26620 4078 26648 5102
rect 27080 4622 27108 5578
rect 27264 5370 27292 6802
rect 27436 6792 27488 6798
rect 27436 6734 27488 6740
rect 27344 6656 27396 6662
rect 27344 6598 27396 6604
rect 27252 5364 27304 5370
rect 27252 5306 27304 5312
rect 27356 4690 27384 6598
rect 27448 6390 27476 6734
rect 27436 6384 27488 6390
rect 27436 6326 27488 6332
rect 27344 4684 27396 4690
rect 27344 4626 27396 4632
rect 27068 4616 27120 4622
rect 27068 4558 27120 4564
rect 26608 4072 26660 4078
rect 26608 4014 26660 4020
rect 27436 4072 27488 4078
rect 27436 4014 27488 4020
rect 27160 3936 27212 3942
rect 27212 3896 27384 3924
rect 27160 3878 27212 3884
rect 27068 3528 27120 3534
rect 27068 3470 27120 3476
rect 27080 2650 27108 3470
rect 27356 3210 27384 3896
rect 27448 3738 27476 4014
rect 27540 4010 27568 12378
rect 27632 12306 27660 13874
rect 27724 13326 27752 14418
rect 27712 13320 27764 13326
rect 27712 13262 27764 13268
rect 27724 12714 27752 13262
rect 27712 12708 27764 12714
rect 27712 12650 27764 12656
rect 27712 12436 27764 12442
rect 27712 12378 27764 12384
rect 27620 12300 27672 12306
rect 27620 12242 27672 12248
rect 27620 11892 27672 11898
rect 27620 11834 27672 11840
rect 27632 11064 27660 11834
rect 27724 11778 27752 12378
rect 27816 12102 27844 14554
rect 28092 14550 28120 15982
rect 28080 14544 28132 14550
rect 28080 14486 28132 14492
rect 28080 14408 28132 14414
rect 28080 14350 28132 14356
rect 28092 13938 28120 14350
rect 28080 13932 28132 13938
rect 28080 13874 28132 13880
rect 27896 13864 27948 13870
rect 27896 13806 27948 13812
rect 27804 12096 27856 12102
rect 27804 12038 27856 12044
rect 27816 11898 27844 12038
rect 27804 11892 27856 11898
rect 27804 11834 27856 11840
rect 27724 11750 27844 11778
rect 27816 11694 27844 11750
rect 27712 11688 27764 11694
rect 27712 11630 27764 11636
rect 27804 11688 27856 11694
rect 27804 11630 27856 11636
rect 27724 11286 27752 11630
rect 27712 11280 27764 11286
rect 27712 11222 27764 11228
rect 27632 11036 27752 11064
rect 27620 8424 27672 8430
rect 27620 8366 27672 8372
rect 27632 8090 27660 8366
rect 27620 8084 27672 8090
rect 27620 8026 27672 8032
rect 27724 7970 27752 11036
rect 27804 10532 27856 10538
rect 27804 10474 27856 10480
rect 27816 9042 27844 10474
rect 27908 9518 27936 13806
rect 28080 13388 28132 13394
rect 28080 13330 28132 13336
rect 28092 12442 28120 13330
rect 28080 12436 28132 12442
rect 28080 12378 28132 12384
rect 28080 12164 28132 12170
rect 28080 12106 28132 12112
rect 27988 11688 28040 11694
rect 27988 11630 28040 11636
rect 28000 11354 28028 11630
rect 27988 11348 28040 11354
rect 27988 11290 28040 11296
rect 27896 9512 27948 9518
rect 27896 9454 27948 9460
rect 28092 9042 28120 12106
rect 28184 9926 28212 18584
rect 28276 16998 28304 18634
rect 28368 18290 28396 22986
rect 28460 21078 28488 23462
rect 28538 22536 28594 22545
rect 28538 22471 28594 22480
rect 28552 22438 28580 22471
rect 28540 22432 28592 22438
rect 28540 22374 28592 22380
rect 28448 21072 28500 21078
rect 28448 21014 28500 21020
rect 28448 19304 28500 19310
rect 28448 19246 28500 19252
rect 28356 18284 28408 18290
rect 28356 18226 28408 18232
rect 28264 16992 28316 16998
rect 28264 16934 28316 16940
rect 28264 16652 28316 16658
rect 28264 16594 28316 16600
rect 28276 16046 28304 16594
rect 28264 16040 28316 16046
rect 28264 15982 28316 15988
rect 28276 14482 28304 15982
rect 28356 14884 28408 14890
rect 28356 14826 28408 14832
rect 28264 14476 28316 14482
rect 28264 14418 28316 14424
rect 28368 12918 28396 14826
rect 28356 12912 28408 12918
rect 28356 12854 28408 12860
rect 28356 12708 28408 12714
rect 28356 12650 28408 12656
rect 28368 12374 28396 12650
rect 28356 12368 28408 12374
rect 28356 12310 28408 12316
rect 28264 12300 28316 12306
rect 28264 12242 28316 12248
rect 28276 11150 28304 12242
rect 28264 11144 28316 11150
rect 28264 11086 28316 11092
rect 28172 9920 28224 9926
rect 28172 9862 28224 9868
rect 28460 9738 28488 19246
rect 28736 18873 28764 34478
rect 28908 34196 28960 34202
rect 28908 34138 28960 34144
rect 28920 33658 28948 34138
rect 28908 33652 28960 33658
rect 28908 33594 28960 33600
rect 29184 33652 29236 33658
rect 29184 33594 29236 33600
rect 29092 32768 29144 32774
rect 29092 32710 29144 32716
rect 29104 32502 29132 32710
rect 29092 32496 29144 32502
rect 29196 32473 29224 33594
rect 29288 32586 29316 34546
rect 29644 34060 29696 34066
rect 29644 34002 29696 34008
rect 29552 33992 29604 33998
rect 29552 33934 29604 33940
rect 29564 33658 29592 33934
rect 29552 33652 29604 33658
rect 29552 33594 29604 33600
rect 29552 32904 29604 32910
rect 29552 32846 29604 32852
rect 29288 32570 29408 32586
rect 29288 32564 29420 32570
rect 29288 32558 29368 32564
rect 29092 32438 29144 32444
rect 29182 32464 29238 32473
rect 29182 32399 29238 32408
rect 29000 32292 29052 32298
rect 29000 32234 29052 32240
rect 28816 31884 28868 31890
rect 28816 31826 28868 31832
rect 28828 19281 28856 31826
rect 28908 31816 28960 31822
rect 28908 31758 28960 31764
rect 28920 29714 28948 31758
rect 29012 30598 29040 32234
rect 29000 30592 29052 30598
rect 29000 30534 29052 30540
rect 29184 30592 29236 30598
rect 29184 30534 29236 30540
rect 28908 29708 28960 29714
rect 28908 29650 28960 29656
rect 29000 29232 29052 29238
rect 29000 29174 29052 29180
rect 29012 28762 29040 29174
rect 29196 29102 29224 30534
rect 29092 29096 29144 29102
rect 29092 29038 29144 29044
rect 29184 29096 29236 29102
rect 29184 29038 29236 29044
rect 29000 28756 29052 28762
rect 29000 28698 29052 28704
rect 29104 28694 29132 29038
rect 29092 28688 29144 28694
rect 29092 28630 29144 28636
rect 29092 28416 29144 28422
rect 29092 28358 29144 28364
rect 29104 27538 29132 28358
rect 29196 28150 29224 29038
rect 29184 28144 29236 28150
rect 29184 28086 29236 28092
rect 29288 28082 29316 32558
rect 29368 32506 29420 32512
rect 29564 32366 29592 32846
rect 29552 32360 29604 32366
rect 29552 32302 29604 32308
rect 29460 31136 29512 31142
rect 29460 31078 29512 31084
rect 29368 29504 29420 29510
rect 29368 29446 29420 29452
rect 29276 28076 29328 28082
rect 29276 28018 29328 28024
rect 29380 28014 29408 29446
rect 29368 28008 29420 28014
rect 29368 27950 29420 27956
rect 29472 27878 29500 31078
rect 29656 30870 29684 34002
rect 29840 33998 29868 34546
rect 30196 34468 30248 34474
rect 30196 34410 30248 34416
rect 29828 33992 29880 33998
rect 29828 33934 29880 33940
rect 29736 33924 29788 33930
rect 29736 33866 29788 33872
rect 29748 31346 29776 33866
rect 29920 33312 29972 33318
rect 29920 33254 29972 33260
rect 29736 31340 29788 31346
rect 29736 31282 29788 31288
rect 29644 30864 29696 30870
rect 29644 30806 29696 30812
rect 29736 30728 29788 30734
rect 29736 30670 29788 30676
rect 29644 30116 29696 30122
rect 29644 30058 29696 30064
rect 29656 29782 29684 30058
rect 29644 29776 29696 29782
rect 29644 29718 29696 29724
rect 29552 29096 29604 29102
rect 29552 29038 29604 29044
rect 29564 28218 29592 29038
rect 29552 28212 29604 28218
rect 29552 28154 29604 28160
rect 29460 27872 29512 27878
rect 29460 27814 29512 27820
rect 29092 27532 29144 27538
rect 29092 27474 29144 27480
rect 29184 27532 29236 27538
rect 29472 27520 29500 27814
rect 29656 27674 29684 29718
rect 29748 29510 29776 30670
rect 29828 30184 29880 30190
rect 29828 30126 29880 30132
rect 29840 29646 29868 30126
rect 29828 29640 29880 29646
rect 29828 29582 29880 29588
rect 29736 29504 29788 29510
rect 29736 29446 29788 29452
rect 29644 27668 29696 27674
rect 29644 27610 29696 27616
rect 29472 27492 29592 27520
rect 29184 27474 29236 27480
rect 29000 27396 29052 27402
rect 29196 27384 29224 27474
rect 29052 27356 29224 27384
rect 29460 27396 29512 27402
rect 29000 27338 29052 27344
rect 29460 27338 29512 27344
rect 29472 26994 29500 27338
rect 29460 26988 29512 26994
rect 29460 26930 29512 26936
rect 29564 26450 29592 27492
rect 29736 27328 29788 27334
rect 29736 27270 29788 27276
rect 29748 27062 29776 27270
rect 29736 27056 29788 27062
rect 29736 26998 29788 27004
rect 29552 26444 29604 26450
rect 29552 26386 29604 26392
rect 29368 26376 29420 26382
rect 29368 26318 29420 26324
rect 29276 24744 29328 24750
rect 29276 24686 29328 24692
rect 29000 22772 29052 22778
rect 29000 22714 29052 22720
rect 29012 21554 29040 22714
rect 29092 22092 29144 22098
rect 29092 22034 29144 22040
rect 29000 21548 29052 21554
rect 29000 21490 29052 21496
rect 28908 21072 28960 21078
rect 28908 21014 28960 21020
rect 28814 19272 28870 19281
rect 28814 19207 28870 19216
rect 28920 19145 28948 21014
rect 29000 19712 29052 19718
rect 29000 19654 29052 19660
rect 28906 19136 28962 19145
rect 28906 19071 28962 19080
rect 28722 18864 28778 18873
rect 28722 18799 28778 18808
rect 28906 18728 28962 18737
rect 28906 18663 28962 18672
rect 28920 18630 28948 18663
rect 28908 18624 28960 18630
rect 28908 18566 28960 18572
rect 28538 18456 28594 18465
rect 28538 18391 28540 18400
rect 28592 18391 28594 18400
rect 28540 18362 28592 18368
rect 28632 18216 28684 18222
rect 28632 18158 28684 18164
rect 28644 17814 28672 18158
rect 29012 18086 29040 19654
rect 29104 19553 29132 22034
rect 29184 21888 29236 21894
rect 29184 21830 29236 21836
rect 29196 21486 29224 21830
rect 29184 21480 29236 21486
rect 29184 21422 29236 21428
rect 29288 20482 29316 24686
rect 29380 22420 29408 26318
rect 29564 25838 29592 26386
rect 29552 25832 29604 25838
rect 29472 25792 29552 25820
rect 29472 24886 29500 25792
rect 29552 25774 29604 25780
rect 29552 25356 29604 25362
rect 29552 25298 29604 25304
rect 29460 24880 29512 24886
rect 29460 24822 29512 24828
rect 29460 24200 29512 24206
rect 29460 24142 29512 24148
rect 29472 22778 29500 24142
rect 29564 23866 29592 25298
rect 29644 25288 29696 25294
rect 29644 25230 29696 25236
rect 29552 23860 29604 23866
rect 29552 23802 29604 23808
rect 29460 22772 29512 22778
rect 29460 22714 29512 22720
rect 29472 22574 29500 22714
rect 29460 22568 29512 22574
rect 29460 22510 29512 22516
rect 29380 22392 29500 22420
rect 29368 21344 29420 21350
rect 29368 21286 29420 21292
rect 29196 20454 29316 20482
rect 29196 20398 29224 20454
rect 29184 20392 29236 20398
rect 29184 20334 29236 20340
rect 29276 20324 29328 20330
rect 29276 20266 29328 20272
rect 29184 20256 29236 20262
rect 29184 20198 29236 20204
rect 29090 19544 29146 19553
rect 29090 19479 29146 19488
rect 29104 19310 29132 19479
rect 29092 19304 29144 19310
rect 29092 19246 29144 19252
rect 29092 18760 29144 18766
rect 29092 18702 29144 18708
rect 29000 18080 29052 18086
rect 29000 18022 29052 18028
rect 29000 17876 29052 17882
rect 29000 17818 29052 17824
rect 28632 17808 28684 17814
rect 28632 17750 28684 17756
rect 28540 17740 28592 17746
rect 28540 17682 28592 17688
rect 28552 15434 28580 17682
rect 28632 17672 28684 17678
rect 28632 17614 28684 17620
rect 28644 16658 28672 17614
rect 29012 17270 29040 17818
rect 29000 17264 29052 17270
rect 29000 17206 29052 17212
rect 28816 16992 28868 16998
rect 28816 16934 28868 16940
rect 28632 16652 28684 16658
rect 28632 16594 28684 16600
rect 28724 15700 28776 15706
rect 28724 15642 28776 15648
rect 28736 15570 28764 15642
rect 28724 15564 28776 15570
rect 28724 15506 28776 15512
rect 28540 15428 28592 15434
rect 28540 15370 28592 15376
rect 28630 14512 28686 14521
rect 28540 14476 28592 14482
rect 28630 14447 28686 14456
rect 28540 14418 28592 14424
rect 28552 13938 28580 14418
rect 28540 13932 28592 13938
rect 28540 13874 28592 13880
rect 28540 13796 28592 13802
rect 28540 13738 28592 13744
rect 28552 10606 28580 13738
rect 28540 10600 28592 10606
rect 28540 10542 28592 10548
rect 28368 9710 28488 9738
rect 27804 9036 27856 9042
rect 27804 8978 27856 8984
rect 28080 9036 28132 9042
rect 28080 8978 28132 8984
rect 27632 7942 27752 7970
rect 27632 7410 27660 7942
rect 28172 7880 28224 7886
rect 28172 7822 28224 7828
rect 28184 7410 28212 7822
rect 27620 7404 27672 7410
rect 27620 7346 27672 7352
rect 28172 7404 28224 7410
rect 28172 7346 28224 7352
rect 28080 7336 28132 7342
rect 28080 7278 28132 7284
rect 27896 6792 27948 6798
rect 27896 6734 27948 6740
rect 27908 4690 27936 6734
rect 27896 4684 27948 4690
rect 27896 4626 27948 4632
rect 27528 4004 27580 4010
rect 27528 3946 27580 3952
rect 27436 3732 27488 3738
rect 27436 3674 27488 3680
rect 27908 3670 27936 4626
rect 27620 3664 27672 3670
rect 27620 3606 27672 3612
rect 27896 3664 27948 3670
rect 27896 3606 27948 3612
rect 27356 3194 27476 3210
rect 27356 3188 27488 3194
rect 27356 3182 27436 3188
rect 27436 3130 27488 3136
rect 27632 2990 27660 3606
rect 27896 3528 27948 3534
rect 28092 3505 28120 7278
rect 28172 6656 28224 6662
rect 28172 6598 28224 6604
rect 28184 5574 28212 6598
rect 28264 5704 28316 5710
rect 28264 5646 28316 5652
rect 28172 5568 28224 5574
rect 28172 5510 28224 5516
rect 28276 5370 28304 5646
rect 28368 5574 28396 9710
rect 28448 9648 28500 9654
rect 28448 9590 28500 9596
rect 28460 9042 28488 9590
rect 28552 9382 28580 10542
rect 28540 9376 28592 9382
rect 28540 9318 28592 9324
rect 28448 9036 28500 9042
rect 28448 8978 28500 8984
rect 28644 8650 28672 14447
rect 28736 13870 28764 15506
rect 28724 13864 28776 13870
rect 28724 13806 28776 13812
rect 28724 13728 28776 13734
rect 28724 13670 28776 13676
rect 28460 8622 28672 8650
rect 28356 5568 28408 5574
rect 28356 5510 28408 5516
rect 28264 5364 28316 5370
rect 28264 5306 28316 5312
rect 28276 4622 28304 5306
rect 28264 4616 28316 4622
rect 28264 4558 28316 4564
rect 28368 4214 28396 5510
rect 28356 4208 28408 4214
rect 28356 4150 28408 4156
rect 28460 4049 28488 8622
rect 28632 8560 28684 8566
rect 28632 8502 28684 8508
rect 28540 8288 28592 8294
rect 28540 8230 28592 8236
rect 28552 7750 28580 8230
rect 28540 7744 28592 7750
rect 28540 7686 28592 7692
rect 28552 6254 28580 7686
rect 28540 6248 28592 6254
rect 28540 6190 28592 6196
rect 28644 5914 28672 8502
rect 28736 8294 28764 13670
rect 28828 9042 28856 16934
rect 29104 16590 29132 18702
rect 29196 17814 29224 20198
rect 29288 18170 29316 20266
rect 29380 20058 29408 21286
rect 29368 20052 29420 20058
rect 29368 19994 29420 20000
rect 29368 19236 29420 19242
rect 29368 19178 29420 19184
rect 29380 18834 29408 19178
rect 29368 18828 29420 18834
rect 29368 18770 29420 18776
rect 29288 18142 29408 18170
rect 29380 17882 29408 18142
rect 29368 17876 29420 17882
rect 29368 17818 29420 17824
rect 29184 17808 29236 17814
rect 29184 17750 29236 17756
rect 29368 17740 29420 17746
rect 29368 17682 29420 17688
rect 29276 17604 29328 17610
rect 29276 17546 29328 17552
rect 29092 16584 29144 16590
rect 29092 16526 29144 16532
rect 28908 16176 28960 16182
rect 28908 16118 28960 16124
rect 28920 15026 28948 16118
rect 29184 15564 29236 15570
rect 29184 15506 29236 15512
rect 29000 15496 29052 15502
rect 29000 15438 29052 15444
rect 29012 15162 29040 15438
rect 29000 15156 29052 15162
rect 29000 15098 29052 15104
rect 28908 15020 28960 15026
rect 28908 14962 28960 14968
rect 29196 14958 29224 15506
rect 29184 14952 29236 14958
rect 29184 14894 29236 14900
rect 28908 14816 28960 14822
rect 28908 14758 28960 14764
rect 28920 13870 28948 14758
rect 29092 14476 29144 14482
rect 29092 14418 29144 14424
rect 29104 13870 29132 14418
rect 28908 13864 28960 13870
rect 28908 13806 28960 13812
rect 29092 13864 29144 13870
rect 29092 13806 29144 13812
rect 28908 13728 28960 13734
rect 28908 13670 28960 13676
rect 28920 13326 28948 13670
rect 29000 13388 29052 13394
rect 29000 13330 29052 13336
rect 28908 13320 28960 13326
rect 28908 13262 28960 13268
rect 28920 12170 28948 13262
rect 28908 12164 28960 12170
rect 28908 12106 28960 12112
rect 29012 11762 29040 13330
rect 29092 12708 29144 12714
rect 29092 12650 29144 12656
rect 29104 12442 29132 12650
rect 29092 12436 29144 12442
rect 29092 12378 29144 12384
rect 29000 11756 29052 11762
rect 29000 11698 29052 11704
rect 29000 11076 29052 11082
rect 29000 11018 29052 11024
rect 28908 11008 28960 11014
rect 28908 10950 28960 10956
rect 28920 9994 28948 10950
rect 29012 10198 29040 11018
rect 29092 11008 29144 11014
rect 29092 10950 29144 10956
rect 29104 10266 29132 10950
rect 29196 10538 29224 14894
rect 29288 11778 29316 17546
rect 29380 14346 29408 17682
rect 29368 14340 29420 14346
rect 29368 14282 29420 14288
rect 29368 13864 29420 13870
rect 29368 13806 29420 13812
rect 29380 13530 29408 13806
rect 29368 13524 29420 13530
rect 29368 13466 29420 13472
rect 29472 11880 29500 22392
rect 29552 22092 29604 22098
rect 29552 22034 29604 22040
rect 29564 20874 29592 22034
rect 29552 20868 29604 20874
rect 29552 20810 29604 20816
rect 29552 20392 29604 20398
rect 29552 20334 29604 20340
rect 29564 19514 29592 20334
rect 29552 19508 29604 19514
rect 29552 19450 29604 19456
rect 29656 19394 29684 25230
rect 29828 22568 29880 22574
rect 29828 22510 29880 22516
rect 29840 22234 29868 22510
rect 29828 22228 29880 22234
rect 29828 22170 29880 22176
rect 29828 20936 29880 20942
rect 29828 20878 29880 20884
rect 29736 19916 29788 19922
rect 29736 19858 29788 19864
rect 29748 19718 29776 19858
rect 29736 19712 29788 19718
rect 29736 19654 29788 19660
rect 29656 19378 29776 19394
rect 29656 19372 29788 19378
rect 29656 19366 29736 19372
rect 29736 19314 29788 19320
rect 29644 19304 29696 19310
rect 29644 19246 29696 19252
rect 29656 19145 29684 19246
rect 29642 19136 29698 19145
rect 29564 19094 29642 19122
rect 29564 18290 29592 19094
rect 29642 19071 29698 19080
rect 29734 19000 29790 19009
rect 29734 18935 29790 18944
rect 29552 18284 29604 18290
rect 29552 18226 29604 18232
rect 29644 18216 29696 18222
rect 29644 18158 29696 18164
rect 29656 17746 29684 18158
rect 29552 17740 29604 17746
rect 29552 17682 29604 17688
rect 29644 17740 29696 17746
rect 29644 17682 29696 17688
rect 29564 17202 29592 17682
rect 29552 17196 29604 17202
rect 29552 17138 29604 17144
rect 29748 16776 29776 18935
rect 29656 16748 29776 16776
rect 29552 13728 29604 13734
rect 29552 13670 29604 13676
rect 29564 13462 29592 13670
rect 29552 13456 29604 13462
rect 29552 13398 29604 13404
rect 29564 12646 29592 13398
rect 29552 12640 29604 12646
rect 29552 12582 29604 12588
rect 29564 12306 29592 12582
rect 29552 12300 29604 12306
rect 29552 12242 29604 12248
rect 29472 11852 29592 11880
rect 29288 11750 29408 11778
rect 29276 11688 29328 11694
rect 29276 11630 29328 11636
rect 29288 11218 29316 11630
rect 29276 11212 29328 11218
rect 29276 11154 29328 11160
rect 29380 11098 29408 11750
rect 29460 11756 29512 11762
rect 29460 11698 29512 11704
rect 29288 11070 29408 11098
rect 29184 10532 29236 10538
rect 29184 10474 29236 10480
rect 29092 10260 29144 10266
rect 29092 10202 29144 10208
rect 29000 10192 29052 10198
rect 29000 10134 29052 10140
rect 28908 9988 28960 9994
rect 28908 9930 28960 9936
rect 28920 9654 28948 9930
rect 29000 9716 29052 9722
rect 29000 9658 29052 9664
rect 28908 9648 28960 9654
rect 28908 9590 28960 9596
rect 28816 9036 28868 9042
rect 28816 8978 28868 8984
rect 28828 8430 28856 8978
rect 28920 8498 28948 9590
rect 29012 9042 29040 9658
rect 29092 9580 29144 9586
rect 29092 9522 29144 9528
rect 29104 9110 29132 9522
rect 29196 9178 29224 10474
rect 29184 9172 29236 9178
rect 29184 9114 29236 9120
rect 29092 9104 29144 9110
rect 29092 9046 29144 9052
rect 29000 9036 29052 9042
rect 29000 8978 29052 8984
rect 29288 8514 29316 11070
rect 29368 10668 29420 10674
rect 29368 10610 29420 10616
rect 29380 10198 29408 10610
rect 29472 10266 29500 11698
rect 29460 10260 29512 10266
rect 29460 10202 29512 10208
rect 29368 10192 29420 10198
rect 29368 10134 29420 10140
rect 29368 8968 29420 8974
rect 29368 8910 29420 8916
rect 28908 8492 28960 8498
rect 28908 8434 28960 8440
rect 29104 8486 29316 8514
rect 28816 8424 28868 8430
rect 28816 8366 28868 8372
rect 28724 8288 28776 8294
rect 28724 8230 28776 8236
rect 28908 8288 28960 8294
rect 28908 8230 28960 8236
rect 28632 5908 28684 5914
rect 28632 5850 28684 5856
rect 28816 5704 28868 5710
rect 28816 5646 28868 5652
rect 28828 5370 28856 5646
rect 28816 5364 28868 5370
rect 28816 5306 28868 5312
rect 28446 4040 28502 4049
rect 28446 3975 28502 3984
rect 28264 3528 28316 3534
rect 27896 3470 27948 3476
rect 28078 3496 28134 3505
rect 27620 2984 27672 2990
rect 27620 2926 27672 2932
rect 27068 2644 27120 2650
rect 27068 2586 27120 2592
rect 26240 2576 26292 2582
rect 26240 2518 26292 2524
rect 27908 2514 27936 3470
rect 28264 3470 28316 3476
rect 28078 3431 28134 3440
rect 28276 3058 28304 3470
rect 28264 3052 28316 3058
rect 28264 2994 28316 3000
rect 28920 2514 28948 8230
rect 29104 7206 29132 8486
rect 29184 8424 29236 8430
rect 29184 8366 29236 8372
rect 29092 7200 29144 7206
rect 29092 7142 29144 7148
rect 29196 6254 29224 8366
rect 29276 7948 29328 7954
rect 29276 7890 29328 7896
rect 29288 7342 29316 7890
rect 29276 7336 29328 7342
rect 29276 7278 29328 7284
rect 29288 7002 29316 7278
rect 29276 6996 29328 7002
rect 29276 6938 29328 6944
rect 29092 6248 29144 6254
rect 29090 6216 29092 6225
rect 29184 6248 29236 6254
rect 29144 6216 29146 6225
rect 29184 6190 29236 6196
rect 29090 6151 29146 6160
rect 29104 5166 29132 6151
rect 29276 5772 29328 5778
rect 29276 5714 29328 5720
rect 29288 5166 29316 5714
rect 29380 5370 29408 8910
rect 29460 8900 29512 8906
rect 29460 8842 29512 8848
rect 29368 5364 29420 5370
rect 29368 5306 29420 5312
rect 29092 5160 29144 5166
rect 29092 5102 29144 5108
rect 29276 5160 29328 5166
rect 29276 5102 29328 5108
rect 29104 4078 29132 5102
rect 29288 4690 29316 5102
rect 29276 4684 29328 4690
rect 29276 4626 29328 4632
rect 29092 4072 29144 4078
rect 29092 4014 29144 4020
rect 29276 3460 29328 3466
rect 29276 3402 29328 3408
rect 29288 3058 29316 3402
rect 29276 3052 29328 3058
rect 29276 2994 29328 3000
rect 27896 2508 27948 2514
rect 27896 2450 27948 2456
rect 28908 2508 28960 2514
rect 28908 2450 28960 2456
rect 25780 2440 25832 2446
rect 25780 2382 25832 2388
rect 27436 2304 27488 2310
rect 27436 2246 27488 2252
rect 27448 800 27476 2246
rect 29472 800 29500 8842
rect 29564 8514 29592 11852
rect 29656 8906 29684 16748
rect 29840 14618 29868 20878
rect 29828 14612 29880 14618
rect 29828 14554 29880 14560
rect 29736 13252 29788 13258
rect 29736 13194 29788 13200
rect 29748 10062 29776 13194
rect 29840 12850 29868 14554
rect 29828 12844 29880 12850
rect 29828 12786 29880 12792
rect 29828 12436 29880 12442
rect 29828 12378 29880 12384
rect 29840 11218 29868 12378
rect 29828 11212 29880 11218
rect 29828 11154 29880 11160
rect 29828 10736 29880 10742
rect 29828 10678 29880 10684
rect 29840 10198 29868 10678
rect 29828 10192 29880 10198
rect 29828 10134 29880 10140
rect 29736 10056 29788 10062
rect 29736 9998 29788 10004
rect 29748 9081 29776 9998
rect 29828 9580 29880 9586
rect 29828 9522 29880 9528
rect 29734 9072 29790 9081
rect 29734 9007 29790 9016
rect 29644 8900 29696 8906
rect 29644 8842 29696 8848
rect 29564 8486 29684 8514
rect 29552 8424 29604 8430
rect 29552 8366 29604 8372
rect 29564 8022 29592 8366
rect 29552 8016 29604 8022
rect 29552 7958 29604 7964
rect 29656 3210 29684 8486
rect 29840 8022 29868 9522
rect 29932 9217 29960 33254
rect 30012 32224 30064 32230
rect 30012 32166 30064 32172
rect 30024 31890 30052 32166
rect 30012 31884 30064 31890
rect 30012 31826 30064 31832
rect 30104 31884 30156 31890
rect 30104 31826 30156 31832
rect 30116 30190 30144 31826
rect 30208 31822 30236 34410
rect 30196 31816 30248 31822
rect 30196 31758 30248 31764
rect 30300 30258 30328 35226
rect 30668 34542 30696 36518
rect 31208 36372 31260 36378
rect 31208 36314 31260 36320
rect 31220 36106 31248 36314
rect 31208 36100 31260 36106
rect 31208 36042 31260 36048
rect 30840 35488 30892 35494
rect 30840 35430 30892 35436
rect 30656 34536 30708 34542
rect 30656 34478 30708 34484
rect 30380 33856 30432 33862
rect 30380 33798 30432 33804
rect 30392 33454 30420 33798
rect 30564 33652 30616 33658
rect 30564 33594 30616 33600
rect 30380 33448 30432 33454
rect 30380 33390 30432 33396
rect 30576 32978 30604 33594
rect 30852 33114 30880 35430
rect 30932 34944 30984 34950
rect 30932 34886 30984 34892
rect 30840 33108 30892 33114
rect 30840 33050 30892 33056
rect 30564 32972 30616 32978
rect 30564 32914 30616 32920
rect 30380 32428 30432 32434
rect 30380 32370 30432 32376
rect 30392 31226 30420 32370
rect 30840 31952 30892 31958
rect 30840 31894 30892 31900
rect 30392 31198 30696 31226
rect 30380 31136 30432 31142
rect 30380 31078 30432 31084
rect 30288 30252 30340 30258
rect 30288 30194 30340 30200
rect 30104 30184 30156 30190
rect 30104 30126 30156 30132
rect 30012 30048 30064 30054
rect 30012 29990 30064 29996
rect 30104 30048 30156 30054
rect 30392 30002 30420 31078
rect 30564 30728 30616 30734
rect 30564 30670 30616 30676
rect 30576 30258 30604 30670
rect 30564 30252 30616 30258
rect 30564 30194 30616 30200
rect 30472 30116 30524 30122
rect 30472 30058 30524 30064
rect 30156 29996 30420 30002
rect 30104 29990 30420 29996
rect 30024 29714 30052 29990
rect 30116 29974 30420 29990
rect 30104 29844 30156 29850
rect 30104 29786 30156 29792
rect 30012 29708 30064 29714
rect 30012 29650 30064 29656
rect 30024 29306 30052 29650
rect 30012 29300 30064 29306
rect 30012 29242 30064 29248
rect 30012 28484 30064 28490
rect 30012 28426 30064 28432
rect 30024 28218 30052 28426
rect 30012 28212 30064 28218
rect 30012 28154 30064 28160
rect 30012 28076 30064 28082
rect 30012 28018 30064 28024
rect 30024 26926 30052 28018
rect 30012 26920 30064 26926
rect 30012 26862 30064 26868
rect 30116 25974 30144 29786
rect 30288 29232 30340 29238
rect 30288 29174 30340 29180
rect 30300 28626 30328 29174
rect 30288 28620 30340 28626
rect 30288 28562 30340 28568
rect 30300 27062 30328 28562
rect 30392 27470 30420 29974
rect 30484 29850 30512 30058
rect 30668 30002 30696 31198
rect 30748 30592 30800 30598
rect 30748 30534 30800 30540
rect 30760 30258 30788 30534
rect 30748 30252 30800 30258
rect 30748 30194 30800 30200
rect 30576 29974 30696 30002
rect 30472 29844 30524 29850
rect 30472 29786 30524 29792
rect 30472 28620 30524 28626
rect 30472 28562 30524 28568
rect 30484 27538 30512 28562
rect 30472 27532 30524 27538
rect 30472 27474 30524 27480
rect 30380 27464 30432 27470
rect 30380 27406 30432 27412
rect 30576 27334 30604 29974
rect 30656 29844 30708 29850
rect 30656 29786 30708 29792
rect 30668 27538 30696 29786
rect 30852 29782 30880 31894
rect 30944 31890 30972 34886
rect 31220 34678 31248 36042
rect 31300 35488 31352 35494
rect 31300 35430 31352 35436
rect 31208 34672 31260 34678
rect 31208 34614 31260 34620
rect 31116 33108 31168 33114
rect 31116 33050 31168 33056
rect 30932 31884 30984 31890
rect 30932 31826 30984 31832
rect 30840 29776 30892 29782
rect 30840 29718 30892 29724
rect 30656 27532 30708 27538
rect 30656 27474 30708 27480
rect 30944 27402 30972 31826
rect 31024 31816 31076 31822
rect 31024 31758 31076 31764
rect 31036 29714 31064 31758
rect 31128 30734 31156 33050
rect 31116 30728 31168 30734
rect 31116 30670 31168 30676
rect 31220 30274 31248 34614
rect 31128 30246 31248 30274
rect 31024 29708 31076 29714
rect 31024 29650 31076 29656
rect 30932 27396 30984 27402
rect 30932 27338 30984 27344
rect 30564 27328 30616 27334
rect 30564 27270 30616 27276
rect 31024 27328 31076 27334
rect 31024 27270 31076 27276
rect 30288 27056 30340 27062
rect 30288 26998 30340 27004
rect 30932 26920 30984 26926
rect 30932 26862 30984 26868
rect 30564 26852 30616 26858
rect 30616 26812 30696 26840
rect 30564 26794 30616 26800
rect 30104 25968 30156 25974
rect 30104 25910 30156 25916
rect 30564 25832 30616 25838
rect 30564 25774 30616 25780
rect 30576 25362 30604 25774
rect 30564 25356 30616 25362
rect 30564 25298 30616 25304
rect 30564 24812 30616 24818
rect 30564 24754 30616 24760
rect 30012 24744 30064 24750
rect 30012 24686 30064 24692
rect 30024 21350 30052 24686
rect 30104 24676 30156 24682
rect 30104 24618 30156 24624
rect 30116 24274 30144 24618
rect 30104 24268 30156 24274
rect 30104 24210 30156 24216
rect 30288 24200 30340 24206
rect 30340 24160 30420 24188
rect 30288 24142 30340 24148
rect 30288 23520 30340 23526
rect 30288 23462 30340 23468
rect 30300 23186 30328 23462
rect 30288 23180 30340 23186
rect 30288 23122 30340 23128
rect 30300 22574 30328 23122
rect 30288 22568 30340 22574
rect 30288 22510 30340 22516
rect 30300 22098 30328 22510
rect 30288 22092 30340 22098
rect 30288 22034 30340 22040
rect 30012 21344 30064 21350
rect 30012 21286 30064 21292
rect 30288 21072 30340 21078
rect 30288 21014 30340 21020
rect 30300 20602 30328 21014
rect 30288 20596 30340 20602
rect 30288 20538 30340 20544
rect 30104 20460 30156 20466
rect 30104 20402 30156 20408
rect 30012 20256 30064 20262
rect 30012 20198 30064 20204
rect 30024 18465 30052 20198
rect 30116 19990 30144 20402
rect 30104 19984 30156 19990
rect 30104 19926 30156 19932
rect 30286 19544 30342 19553
rect 30286 19479 30342 19488
rect 30104 19304 30156 19310
rect 30104 19246 30156 19252
rect 30010 18456 30066 18465
rect 30010 18391 30066 18400
rect 30024 18290 30052 18391
rect 30012 18284 30064 18290
rect 30012 18226 30064 18232
rect 30116 17610 30144 19246
rect 30300 18426 30328 19479
rect 30392 19174 30420 24160
rect 30472 23112 30524 23118
rect 30472 23054 30524 23060
rect 30484 22778 30512 23054
rect 30472 22772 30524 22778
rect 30472 22714 30524 22720
rect 30484 20398 30512 22714
rect 30576 20398 30604 24754
rect 30472 20392 30524 20398
rect 30472 20334 30524 20340
rect 30564 20392 30616 20398
rect 30564 20334 30616 20340
rect 30484 19854 30512 20334
rect 30668 20040 30696 26812
rect 30748 26376 30800 26382
rect 30748 26318 30800 26324
rect 30760 25362 30788 26318
rect 30748 25356 30800 25362
rect 30748 25298 30800 25304
rect 30760 25158 30788 25298
rect 30748 25152 30800 25158
rect 30748 25094 30800 25100
rect 30840 24744 30892 24750
rect 30840 24686 30892 24692
rect 30852 23322 30880 24686
rect 30840 23316 30892 23322
rect 30840 23258 30892 23264
rect 30852 22098 30880 23258
rect 30840 22092 30892 22098
rect 30840 22034 30892 22040
rect 30576 20012 30696 20040
rect 30472 19848 30524 19854
rect 30472 19790 30524 19796
rect 30380 19168 30432 19174
rect 30380 19110 30432 19116
rect 30392 18737 30420 19110
rect 30378 18728 30434 18737
rect 30378 18663 30434 18672
rect 30288 18420 30340 18426
rect 30288 18362 30340 18368
rect 30576 18170 30604 20012
rect 30656 19916 30708 19922
rect 30656 19858 30708 19864
rect 30748 19916 30800 19922
rect 30748 19858 30800 19864
rect 30668 19242 30696 19858
rect 30760 19378 30788 19858
rect 30748 19372 30800 19378
rect 30748 19314 30800 19320
rect 30656 19236 30708 19242
rect 30656 19178 30708 19184
rect 30668 18970 30696 19178
rect 30656 18964 30708 18970
rect 30656 18906 30708 18912
rect 30760 18902 30788 19314
rect 30838 19136 30894 19145
rect 30838 19071 30894 19080
rect 30748 18896 30800 18902
rect 30748 18838 30800 18844
rect 30300 18142 30604 18170
rect 30104 17604 30156 17610
rect 30104 17546 30156 17552
rect 30300 17184 30328 18142
rect 30564 18080 30616 18086
rect 30564 18022 30616 18028
rect 30208 17156 30328 17184
rect 30104 16584 30156 16590
rect 30104 16526 30156 16532
rect 30116 16046 30144 16526
rect 30104 16040 30156 16046
rect 30104 15982 30156 15988
rect 30104 15904 30156 15910
rect 30104 15846 30156 15852
rect 30116 15706 30144 15846
rect 30104 15700 30156 15706
rect 30104 15642 30156 15648
rect 30104 15564 30156 15570
rect 30104 15506 30156 15512
rect 30012 15088 30064 15094
rect 30012 15030 30064 15036
rect 30024 14770 30052 15030
rect 30116 14958 30144 15506
rect 30104 14952 30156 14958
rect 30104 14894 30156 14900
rect 30024 14742 30144 14770
rect 30012 14476 30064 14482
rect 30012 14418 30064 14424
rect 30024 13938 30052 14418
rect 30116 14278 30144 14742
rect 30104 14272 30156 14278
rect 30104 14214 30156 14220
rect 30012 13932 30064 13938
rect 30012 13874 30064 13880
rect 30116 12714 30144 14214
rect 30104 12708 30156 12714
rect 30104 12650 30156 12656
rect 30208 12594 30236 17156
rect 30380 17128 30432 17134
rect 30380 17070 30432 17076
rect 30288 17060 30340 17066
rect 30288 17002 30340 17008
rect 30300 16658 30328 17002
rect 30288 16652 30340 16658
rect 30288 16594 30340 16600
rect 30288 16448 30340 16454
rect 30288 16390 30340 16396
rect 30300 15162 30328 16390
rect 30392 15434 30420 17070
rect 30472 17060 30524 17066
rect 30472 17002 30524 17008
rect 30484 16114 30512 17002
rect 30472 16108 30524 16114
rect 30472 16050 30524 16056
rect 30380 15428 30432 15434
rect 30380 15370 30432 15376
rect 30288 15156 30340 15162
rect 30288 15098 30340 15104
rect 30300 14414 30328 15098
rect 30576 14958 30604 18022
rect 30656 17808 30708 17814
rect 30656 17750 30708 17756
rect 30668 17134 30696 17750
rect 30852 17746 30880 19071
rect 30840 17740 30892 17746
rect 30840 17682 30892 17688
rect 30656 17128 30708 17134
rect 30656 17070 30708 17076
rect 30840 16788 30892 16794
rect 30840 16730 30892 16736
rect 30564 14952 30616 14958
rect 30564 14894 30616 14900
rect 30748 14952 30800 14958
rect 30748 14894 30800 14900
rect 30288 14408 30340 14414
rect 30288 14350 30340 14356
rect 30300 13394 30328 14350
rect 30288 13388 30340 13394
rect 30288 13330 30340 13336
rect 30656 13320 30708 13326
rect 30656 13262 30708 13268
rect 30116 12566 30236 12594
rect 30116 9602 30144 12566
rect 30288 12300 30340 12306
rect 30288 12242 30340 12248
rect 30300 11150 30328 12242
rect 30564 12232 30616 12238
rect 30564 12174 30616 12180
rect 30472 11824 30524 11830
rect 30472 11766 30524 11772
rect 30288 11144 30340 11150
rect 30288 11086 30340 11092
rect 30484 10606 30512 11766
rect 30576 11694 30604 12174
rect 30668 11762 30696 13262
rect 30760 12442 30788 14894
rect 30852 13938 30880 16730
rect 30840 13932 30892 13938
rect 30840 13874 30892 13880
rect 30840 13388 30892 13394
rect 30840 13330 30892 13336
rect 30852 12850 30880 13330
rect 30840 12844 30892 12850
rect 30840 12786 30892 12792
rect 30748 12436 30800 12442
rect 30748 12378 30800 12384
rect 30656 11756 30708 11762
rect 30656 11698 30708 11704
rect 30564 11688 30616 11694
rect 30564 11630 30616 11636
rect 30576 11354 30604 11630
rect 30840 11552 30892 11558
rect 30840 11494 30892 11500
rect 30564 11348 30616 11354
rect 30564 11290 30616 11296
rect 30852 11218 30880 11494
rect 30564 11212 30616 11218
rect 30564 11154 30616 11160
rect 30840 11212 30892 11218
rect 30840 11154 30892 11160
rect 30576 10674 30604 11154
rect 30840 11076 30892 11082
rect 30840 11018 30892 11024
rect 30564 10668 30616 10674
rect 30564 10610 30616 10616
rect 30472 10600 30524 10606
rect 30472 10542 30524 10548
rect 30380 9988 30432 9994
rect 30380 9930 30432 9936
rect 30024 9574 30144 9602
rect 29918 9208 29974 9217
rect 29918 9143 29974 9152
rect 29920 8968 29972 8974
rect 29920 8910 29972 8916
rect 29828 8016 29880 8022
rect 29828 7958 29880 7964
rect 29932 7954 29960 8910
rect 29920 7948 29972 7954
rect 29920 7890 29972 7896
rect 29920 6792 29972 6798
rect 29920 6734 29972 6740
rect 29932 6322 29960 6734
rect 29920 6316 29972 6322
rect 29920 6258 29972 6264
rect 29828 6112 29880 6118
rect 29828 6054 29880 6060
rect 29736 5840 29788 5846
rect 29736 5782 29788 5788
rect 29748 4690 29776 5782
rect 29736 4684 29788 4690
rect 29736 4626 29788 4632
rect 29656 3182 29776 3210
rect 29644 3120 29696 3126
rect 29644 3062 29696 3068
rect 29656 2514 29684 3062
rect 29644 2508 29696 2514
rect 29644 2450 29696 2456
rect 29748 1154 29776 3182
rect 29840 3058 29868 6054
rect 30024 4842 30052 9574
rect 30288 9512 30340 9518
rect 30288 9454 30340 9460
rect 30300 9178 30328 9454
rect 30288 9172 30340 9178
rect 30288 9114 30340 9120
rect 30300 7834 30328 9114
rect 30392 7954 30420 9930
rect 30484 9636 30512 10542
rect 30852 9994 30880 11018
rect 30840 9988 30892 9994
rect 30840 9930 30892 9936
rect 30852 9654 30880 9930
rect 30840 9648 30892 9654
rect 30484 9608 30696 9636
rect 30668 9110 30696 9608
rect 30840 9590 30892 9596
rect 30656 9104 30708 9110
rect 30656 9046 30708 9052
rect 30380 7948 30432 7954
rect 30380 7890 30432 7896
rect 30208 7806 30328 7834
rect 30208 6254 30236 7806
rect 30944 7750 30972 26862
rect 31036 26790 31064 27270
rect 31024 26784 31076 26790
rect 31024 26726 31076 26732
rect 31128 24834 31156 30246
rect 31208 30184 31260 30190
rect 31208 30126 31260 30132
rect 31220 29782 31248 30126
rect 31312 29850 31340 35430
rect 31668 32904 31720 32910
rect 31668 32846 31720 32852
rect 31680 32366 31708 32846
rect 31668 32360 31720 32366
rect 31668 32302 31720 32308
rect 31760 31816 31812 31822
rect 31760 31758 31812 31764
rect 31772 31346 31800 31758
rect 31760 31340 31812 31346
rect 31760 31282 31812 31288
rect 31300 29844 31352 29850
rect 31300 29786 31352 29792
rect 31208 29776 31260 29782
rect 31208 29718 31260 29724
rect 31392 28620 31444 28626
rect 31392 28562 31444 28568
rect 31404 27878 31432 28562
rect 31864 27962 31892 37198
rect 31956 35578 31984 37266
rect 32048 35698 32076 37742
rect 32128 37664 32180 37670
rect 32128 37606 32180 37612
rect 32140 37330 32168 37606
rect 32128 37324 32180 37330
rect 32128 37266 32180 37272
rect 32784 36922 32812 37742
rect 33704 37466 33732 40200
rect 34940 38108 35236 38128
rect 34996 38106 35020 38108
rect 35076 38106 35100 38108
rect 35156 38106 35180 38108
rect 35018 38054 35020 38106
rect 35082 38054 35094 38106
rect 35156 38054 35158 38106
rect 34996 38052 35020 38054
rect 35076 38052 35100 38054
rect 35156 38052 35180 38054
rect 34940 38032 35236 38052
rect 35544 37466 35572 40200
rect 35898 38720 35954 38729
rect 35898 38655 35954 38664
rect 35912 38554 35940 38655
rect 35900 38548 35952 38554
rect 35900 38490 35952 38496
rect 33692 37460 33744 37466
rect 33692 37402 33744 37408
rect 35532 37460 35584 37466
rect 35532 37402 35584 37408
rect 35532 37324 35584 37330
rect 35532 37266 35584 37272
rect 34940 37020 35236 37040
rect 34996 37018 35020 37020
rect 35076 37018 35100 37020
rect 35156 37018 35180 37020
rect 35018 36966 35020 37018
rect 35082 36966 35094 37018
rect 35156 36966 35158 37018
rect 34996 36964 35020 36966
rect 35076 36964 35100 36966
rect 35156 36964 35180 36966
rect 34940 36944 35236 36964
rect 32772 36916 32824 36922
rect 32772 36858 32824 36864
rect 32496 36712 32548 36718
rect 32496 36654 32548 36660
rect 32508 36242 32536 36654
rect 34520 36304 34572 36310
rect 34520 36246 34572 36252
rect 32496 36236 32548 36242
rect 32496 36178 32548 36184
rect 33140 36236 33192 36242
rect 33140 36178 33192 36184
rect 33968 36236 34020 36242
rect 33968 36178 34020 36184
rect 32312 36168 32364 36174
rect 32312 36110 32364 36116
rect 32324 35698 32352 36110
rect 33152 35766 33180 36178
rect 33980 35834 34008 36178
rect 34152 36032 34204 36038
rect 34152 35974 34204 35980
rect 33968 35828 34020 35834
rect 33968 35770 34020 35776
rect 33140 35760 33192 35766
rect 33140 35702 33192 35708
rect 32036 35692 32088 35698
rect 32036 35634 32088 35640
rect 32312 35692 32364 35698
rect 32312 35634 32364 35640
rect 31956 35550 32168 35578
rect 32036 35488 32088 35494
rect 32036 35430 32088 35436
rect 32048 35086 32076 35430
rect 32036 35080 32088 35086
rect 32036 35022 32088 35028
rect 31944 33448 31996 33454
rect 31944 33390 31996 33396
rect 31956 30326 31984 33390
rect 32036 31272 32088 31278
rect 32036 31214 32088 31220
rect 32048 30598 32076 31214
rect 32036 30592 32088 30598
rect 32036 30534 32088 30540
rect 32048 30326 32076 30534
rect 31944 30320 31996 30326
rect 31944 30262 31996 30268
rect 32036 30320 32088 30326
rect 32036 30262 32088 30268
rect 32036 29096 32088 29102
rect 32036 29038 32088 29044
rect 31864 27934 31984 27962
rect 31392 27872 31444 27878
rect 31392 27814 31444 27820
rect 31852 27872 31904 27878
rect 31852 27814 31904 27820
rect 31864 27470 31892 27814
rect 31852 27464 31904 27470
rect 31852 27406 31904 27412
rect 31484 27396 31536 27402
rect 31484 27338 31536 27344
rect 31208 26784 31260 26790
rect 31208 26726 31260 26732
rect 31220 26518 31248 26726
rect 31496 26586 31524 27338
rect 31484 26580 31536 26586
rect 31484 26522 31536 26528
rect 31208 26512 31260 26518
rect 31208 26454 31260 26460
rect 31852 25356 31904 25362
rect 31852 25298 31904 25304
rect 31036 24818 31156 24834
rect 31024 24812 31156 24818
rect 31076 24806 31156 24812
rect 31024 24754 31076 24760
rect 31036 24410 31064 24754
rect 31864 24750 31892 25298
rect 31116 24744 31168 24750
rect 31116 24686 31168 24692
rect 31852 24744 31904 24750
rect 31852 24686 31904 24692
rect 31024 24404 31076 24410
rect 31024 24346 31076 24352
rect 31128 23730 31156 24686
rect 31576 24676 31628 24682
rect 31576 24618 31628 24624
rect 31484 24064 31536 24070
rect 31484 24006 31536 24012
rect 31116 23724 31168 23730
rect 31116 23666 31168 23672
rect 31496 23594 31524 24006
rect 31588 23730 31616 24618
rect 31864 24274 31892 24686
rect 31852 24268 31904 24274
rect 31852 24210 31904 24216
rect 31576 23724 31628 23730
rect 31576 23666 31628 23672
rect 31484 23588 31536 23594
rect 31484 23530 31536 23536
rect 31588 22710 31616 23666
rect 31668 23656 31720 23662
rect 31668 23598 31720 23604
rect 31680 23186 31708 23598
rect 31760 23248 31812 23254
rect 31760 23190 31812 23196
rect 31668 23180 31720 23186
rect 31668 23122 31720 23128
rect 31576 22704 31628 22710
rect 31576 22646 31628 22652
rect 31680 22438 31708 23122
rect 31772 22982 31800 23190
rect 31852 23180 31904 23186
rect 31852 23122 31904 23128
rect 31760 22976 31812 22982
rect 31760 22918 31812 22924
rect 31772 22642 31800 22918
rect 31760 22636 31812 22642
rect 31760 22578 31812 22584
rect 31024 22432 31076 22438
rect 31024 22374 31076 22380
rect 31668 22432 31720 22438
rect 31668 22374 31720 22380
rect 31036 20398 31064 22374
rect 31392 22092 31444 22098
rect 31392 22034 31444 22040
rect 31208 20800 31260 20806
rect 31208 20742 31260 20748
rect 31024 20392 31076 20398
rect 31024 20334 31076 20340
rect 31220 18630 31248 20742
rect 31404 20534 31432 22034
rect 31484 21956 31536 21962
rect 31484 21898 31536 21904
rect 31496 21486 31524 21898
rect 31484 21480 31536 21486
rect 31484 21422 31536 21428
rect 31392 20528 31444 20534
rect 31392 20470 31444 20476
rect 31484 20392 31536 20398
rect 31484 20334 31536 20340
rect 31392 19304 31444 19310
rect 31390 19272 31392 19281
rect 31444 19272 31446 19281
rect 31300 19236 31352 19242
rect 31390 19207 31446 19216
rect 31300 19178 31352 19184
rect 31312 18834 31340 19178
rect 31300 18828 31352 18834
rect 31300 18770 31352 18776
rect 31208 18624 31260 18630
rect 31208 18566 31260 18572
rect 31220 18222 31248 18566
rect 31208 18216 31260 18222
rect 31208 18158 31260 18164
rect 31300 17128 31352 17134
rect 31300 17070 31352 17076
rect 31208 14544 31260 14550
rect 31208 14486 31260 14492
rect 31220 14346 31248 14486
rect 31208 14340 31260 14346
rect 31208 14282 31260 14288
rect 31208 13796 31260 13802
rect 31208 13738 31260 13744
rect 31220 13394 31248 13738
rect 31208 13388 31260 13394
rect 31208 13330 31260 13336
rect 31220 12918 31248 13330
rect 31312 13258 31340 17070
rect 31496 15366 31524 20334
rect 31680 20058 31708 22374
rect 31760 21888 31812 21894
rect 31760 21830 31812 21836
rect 31668 20052 31720 20058
rect 31668 19994 31720 20000
rect 31574 19408 31630 19417
rect 31574 19343 31630 19352
rect 31588 18902 31616 19343
rect 31668 19304 31720 19310
rect 31668 19246 31720 19252
rect 31576 18896 31628 18902
rect 31680 18873 31708 19246
rect 31576 18838 31628 18844
rect 31666 18864 31722 18873
rect 31666 18799 31722 18808
rect 31772 18714 31800 21830
rect 31864 21350 31892 23122
rect 31852 21344 31904 21350
rect 31852 21286 31904 21292
rect 31772 18686 31892 18714
rect 31760 17672 31812 17678
rect 31760 17614 31812 17620
rect 31772 17134 31800 17614
rect 31760 17128 31812 17134
rect 31760 17070 31812 17076
rect 31760 16788 31812 16794
rect 31760 16730 31812 16736
rect 31668 15904 31720 15910
rect 31668 15846 31720 15852
rect 31392 15360 31444 15366
rect 31392 15302 31444 15308
rect 31484 15360 31536 15366
rect 31484 15302 31536 15308
rect 31404 15162 31432 15302
rect 31392 15156 31444 15162
rect 31392 15098 31444 15104
rect 31404 13870 31432 15098
rect 31496 14074 31524 15302
rect 31576 15020 31628 15026
rect 31576 14962 31628 14968
rect 31588 14550 31616 14962
rect 31680 14958 31708 15846
rect 31668 14952 31720 14958
rect 31668 14894 31720 14900
rect 31576 14544 31628 14550
rect 31576 14486 31628 14492
rect 31484 14068 31536 14074
rect 31484 14010 31536 14016
rect 31392 13864 31444 13870
rect 31392 13806 31444 13812
rect 31404 13326 31432 13806
rect 31392 13320 31444 13326
rect 31392 13262 31444 13268
rect 31300 13252 31352 13258
rect 31300 13194 31352 13200
rect 31208 12912 31260 12918
rect 31208 12854 31260 12860
rect 31404 12850 31432 13262
rect 31392 12844 31444 12850
rect 31392 12786 31444 12792
rect 31392 12300 31444 12306
rect 31392 12242 31444 12248
rect 31300 12096 31352 12102
rect 31300 12038 31352 12044
rect 31312 10674 31340 12038
rect 31300 10668 31352 10674
rect 31300 10610 31352 10616
rect 31312 10130 31340 10610
rect 31024 10124 31076 10130
rect 31024 10066 31076 10072
rect 31300 10124 31352 10130
rect 31300 10066 31352 10072
rect 31036 8090 31064 10066
rect 31116 9512 31168 9518
rect 31116 9454 31168 9460
rect 31128 9042 31156 9454
rect 31404 9382 31432 12242
rect 31484 11688 31536 11694
rect 31484 11630 31536 11636
rect 31496 11150 31524 11630
rect 31484 11144 31536 11150
rect 31484 11086 31536 11092
rect 31496 10810 31524 11086
rect 31484 10804 31536 10810
rect 31484 10746 31536 10752
rect 31588 10538 31616 14486
rect 31772 13870 31800 16730
rect 31864 15570 31892 18686
rect 31852 15564 31904 15570
rect 31852 15506 31904 15512
rect 31956 15502 31984 27934
rect 32048 27538 32076 29038
rect 32140 28694 32168 35550
rect 34164 35154 34192 35974
rect 34532 35154 34560 36246
rect 35256 36032 35308 36038
rect 35256 35974 35308 35980
rect 34940 35932 35236 35952
rect 34996 35930 35020 35932
rect 35076 35930 35100 35932
rect 35156 35930 35180 35932
rect 35018 35878 35020 35930
rect 35082 35878 35094 35930
rect 35156 35878 35158 35930
rect 34996 35876 35020 35878
rect 35076 35876 35100 35878
rect 35156 35876 35180 35878
rect 34940 35856 35236 35876
rect 35268 35698 35296 35974
rect 35256 35692 35308 35698
rect 35256 35634 35308 35640
rect 35440 35624 35492 35630
rect 35440 35566 35492 35572
rect 34152 35148 34204 35154
rect 34152 35090 34204 35096
rect 34520 35148 34572 35154
rect 34520 35090 34572 35096
rect 35452 35086 35480 35566
rect 32864 35080 32916 35086
rect 32864 35022 32916 35028
rect 35440 35080 35492 35086
rect 35440 35022 35492 35028
rect 32496 34604 32548 34610
rect 32496 34546 32548 34552
rect 32220 34536 32272 34542
rect 32220 34478 32272 34484
rect 32232 31414 32260 34478
rect 32404 33992 32456 33998
rect 32404 33934 32456 33940
rect 32416 33522 32444 33934
rect 32404 33516 32456 33522
rect 32404 33458 32456 33464
rect 32312 33380 32364 33386
rect 32312 33322 32364 33328
rect 32324 32842 32352 33322
rect 32312 32836 32364 32842
rect 32312 32778 32364 32784
rect 32508 31822 32536 34546
rect 32876 34066 32904 35022
rect 33232 34944 33284 34950
rect 33232 34886 33284 34892
rect 33140 34536 33192 34542
rect 33140 34478 33192 34484
rect 33152 34066 33180 34478
rect 32864 34060 32916 34066
rect 32864 34002 32916 34008
rect 33140 34060 33192 34066
rect 33140 34002 33192 34008
rect 32876 33522 32904 34002
rect 32864 33516 32916 33522
rect 32864 33458 32916 33464
rect 33244 33114 33272 34886
rect 34940 34844 35236 34864
rect 34996 34842 35020 34844
rect 35076 34842 35100 34844
rect 35156 34842 35180 34844
rect 35018 34790 35020 34842
rect 35082 34790 35094 34842
rect 35156 34790 35158 34842
rect 34996 34788 35020 34790
rect 35076 34788 35100 34790
rect 35156 34788 35180 34790
rect 34940 34768 35236 34788
rect 35452 34610 35480 35022
rect 34060 34604 34112 34610
rect 34060 34546 34112 34552
rect 35440 34604 35492 34610
rect 35440 34546 35492 34552
rect 33324 34536 33376 34542
rect 33324 34478 33376 34484
rect 33232 33108 33284 33114
rect 33232 33050 33284 33056
rect 33336 32978 33364 34478
rect 33508 33856 33560 33862
rect 33508 33798 33560 33804
rect 33520 33402 33548 33798
rect 34072 33658 34100 34546
rect 35348 34400 35400 34406
rect 35348 34342 35400 34348
rect 34796 34060 34848 34066
rect 34796 34002 34848 34008
rect 34336 33856 34388 33862
rect 34336 33798 34388 33804
rect 34060 33652 34112 33658
rect 34060 33594 34112 33600
rect 33600 33448 33652 33454
rect 33520 33396 33600 33402
rect 33520 33390 33652 33396
rect 33520 33374 33640 33390
rect 33520 33046 33548 33374
rect 33508 33040 33560 33046
rect 33508 32982 33560 32988
rect 34072 32978 34100 33594
rect 34348 33522 34376 33798
rect 34336 33516 34388 33522
rect 34336 33458 34388 33464
rect 34520 33312 34572 33318
rect 34520 33254 34572 33260
rect 34532 32978 34560 33254
rect 33324 32972 33376 32978
rect 33324 32914 33376 32920
rect 34060 32972 34112 32978
rect 34060 32914 34112 32920
rect 34520 32972 34572 32978
rect 34520 32914 34572 32920
rect 33336 32858 33364 32914
rect 32772 32836 32824 32842
rect 33336 32830 33548 32858
rect 32772 32778 32824 32784
rect 32496 31816 32548 31822
rect 32496 31758 32548 31764
rect 32680 31680 32732 31686
rect 32680 31622 32732 31628
rect 32220 31408 32272 31414
rect 32220 31350 32272 31356
rect 32692 31210 32720 31622
rect 32680 31204 32732 31210
rect 32680 31146 32732 31152
rect 32692 30734 32720 31146
rect 32680 30728 32732 30734
rect 32680 30670 32732 30676
rect 32692 30054 32720 30670
rect 32680 30048 32732 30054
rect 32680 29990 32732 29996
rect 32128 28688 32180 28694
rect 32128 28630 32180 28636
rect 32404 28416 32456 28422
rect 32404 28358 32456 28364
rect 32416 28082 32444 28358
rect 32404 28076 32456 28082
rect 32404 28018 32456 28024
rect 32036 27532 32088 27538
rect 32036 27474 32088 27480
rect 32048 26450 32076 27474
rect 32496 27396 32548 27402
rect 32496 27338 32548 27344
rect 32036 26444 32088 26450
rect 32036 26386 32088 26392
rect 32508 26314 32536 27338
rect 32496 26308 32548 26314
rect 32496 26250 32548 26256
rect 32404 25424 32456 25430
rect 32404 25366 32456 25372
rect 32128 24268 32180 24274
rect 32128 24210 32180 24216
rect 32036 23520 32088 23526
rect 32036 23462 32088 23468
rect 32048 23118 32076 23462
rect 32140 23186 32168 24210
rect 32220 23316 32272 23322
rect 32220 23258 32272 23264
rect 32128 23180 32180 23186
rect 32128 23122 32180 23128
rect 32036 23112 32088 23118
rect 32036 23054 32088 23060
rect 32048 22574 32076 23054
rect 32140 22778 32168 23122
rect 32128 22772 32180 22778
rect 32128 22714 32180 22720
rect 32036 22568 32088 22574
rect 32036 22510 32088 22516
rect 32232 22166 32260 23258
rect 32416 22778 32444 25366
rect 32508 25294 32536 26250
rect 32680 25356 32732 25362
rect 32680 25298 32732 25304
rect 32496 25288 32548 25294
rect 32496 25230 32548 25236
rect 32588 24268 32640 24274
rect 32588 24210 32640 24216
rect 32496 24200 32548 24206
rect 32496 24142 32548 24148
rect 32508 23798 32536 24142
rect 32600 23798 32628 24210
rect 32692 23866 32720 25298
rect 32784 24614 32812 32778
rect 32956 32360 33008 32366
rect 32956 32302 33008 32308
rect 33324 32360 33376 32366
rect 33324 32302 33376 32308
rect 32968 30802 32996 32302
rect 33232 32292 33284 32298
rect 33232 32234 33284 32240
rect 32956 30796 33008 30802
rect 32956 30738 33008 30744
rect 33244 30546 33272 32234
rect 33060 30518 33272 30546
rect 33060 30394 33088 30518
rect 33336 30410 33364 32302
rect 33520 32230 33548 32830
rect 33784 32360 33836 32366
rect 33784 32302 33836 32308
rect 33508 32224 33560 32230
rect 33508 32166 33560 32172
rect 33416 31272 33468 31278
rect 33416 31214 33468 31220
rect 33428 30938 33456 31214
rect 33416 30932 33468 30938
rect 33416 30874 33468 30880
rect 33048 30388 33100 30394
rect 33048 30330 33100 30336
rect 33152 30382 33364 30410
rect 33048 30048 33100 30054
rect 33048 29990 33100 29996
rect 33060 29714 33088 29990
rect 33048 29708 33100 29714
rect 33048 29650 33100 29656
rect 33060 28626 33088 29650
rect 33152 28966 33180 30382
rect 33428 30274 33456 30874
rect 33336 30246 33456 30274
rect 33336 30190 33364 30246
rect 33520 30190 33548 32166
rect 33796 32026 33824 32302
rect 34532 32298 34560 32914
rect 34520 32292 34572 32298
rect 34520 32234 34572 32240
rect 33784 32020 33836 32026
rect 33784 31962 33836 31968
rect 34532 31346 34560 32234
rect 34704 31816 34756 31822
rect 34704 31758 34756 31764
rect 34520 31340 34572 31346
rect 34520 31282 34572 31288
rect 34532 30394 34560 31282
rect 34520 30388 34572 30394
rect 34520 30330 34572 30336
rect 34152 30320 34204 30326
rect 34152 30262 34204 30268
rect 33324 30184 33376 30190
rect 33324 30126 33376 30132
rect 33508 30184 33560 30190
rect 33508 30126 33560 30132
rect 33232 29640 33284 29646
rect 33232 29582 33284 29588
rect 33244 29238 33272 29582
rect 33232 29232 33284 29238
rect 33232 29174 33284 29180
rect 33140 28960 33192 28966
rect 33140 28902 33192 28908
rect 33048 28620 33100 28626
rect 33048 28562 33100 28568
rect 33416 28552 33468 28558
rect 33416 28494 33468 28500
rect 33428 28082 33456 28494
rect 33520 28218 33548 30126
rect 34164 29102 34192 30262
rect 34428 30184 34480 30190
rect 34428 30126 34480 30132
rect 34520 30184 34572 30190
rect 34520 30126 34572 30132
rect 34440 29578 34468 30126
rect 34428 29572 34480 29578
rect 34428 29514 34480 29520
rect 34152 29096 34204 29102
rect 34152 29038 34204 29044
rect 33508 28212 33560 28218
rect 33508 28154 33560 28160
rect 33416 28076 33468 28082
rect 33416 28018 33468 28024
rect 33324 28008 33376 28014
rect 33324 27950 33376 27956
rect 33336 27538 33364 27950
rect 33520 27946 33548 28154
rect 33968 28008 34020 28014
rect 33968 27950 34020 27956
rect 33508 27940 33560 27946
rect 33508 27882 33560 27888
rect 33980 27538 34008 27950
rect 34060 27872 34112 27878
rect 34060 27814 34112 27820
rect 33324 27532 33376 27538
rect 33324 27474 33376 27480
rect 33968 27532 34020 27538
rect 33968 27474 34020 27480
rect 33048 27464 33100 27470
rect 33048 27406 33100 27412
rect 33060 26790 33088 27406
rect 33980 27402 34008 27474
rect 33968 27396 34020 27402
rect 33968 27338 34020 27344
rect 34072 26926 34100 27814
rect 34164 27334 34192 29038
rect 34440 28694 34468 29514
rect 34532 29510 34560 30126
rect 34520 29504 34572 29510
rect 34520 29446 34572 29452
rect 34532 29034 34560 29446
rect 34520 29028 34572 29034
rect 34520 28970 34572 28976
rect 34428 28688 34480 28694
rect 34428 28630 34480 28636
rect 34244 27532 34296 27538
rect 34244 27474 34296 27480
rect 34152 27328 34204 27334
rect 34152 27270 34204 27276
rect 34164 26994 34192 27270
rect 34152 26988 34204 26994
rect 34152 26930 34204 26936
rect 33140 26920 33192 26926
rect 33140 26862 33192 26868
rect 34060 26920 34112 26926
rect 34060 26862 34112 26868
rect 33048 26784 33100 26790
rect 33048 26726 33100 26732
rect 33152 26518 33180 26862
rect 33784 26784 33836 26790
rect 33784 26726 33836 26732
rect 33140 26512 33192 26518
rect 33140 26454 33192 26460
rect 33796 26450 33824 26726
rect 33784 26444 33836 26450
rect 33784 26386 33836 26392
rect 33324 26376 33376 26382
rect 33324 26318 33376 26324
rect 33508 26376 33560 26382
rect 33508 26318 33560 26324
rect 33336 26042 33364 26318
rect 33324 26036 33376 26042
rect 33324 25978 33376 25984
rect 33520 25906 33548 26318
rect 33508 25900 33560 25906
rect 33508 25842 33560 25848
rect 34072 25838 34100 26862
rect 34256 26042 34284 27474
rect 34244 26036 34296 26042
rect 34244 25978 34296 25984
rect 33876 25832 33928 25838
rect 33876 25774 33928 25780
rect 34060 25832 34112 25838
rect 34060 25774 34112 25780
rect 33140 25356 33192 25362
rect 33140 25298 33192 25304
rect 33152 24818 33180 25298
rect 33140 24812 33192 24818
rect 33140 24754 33192 24760
rect 33324 24744 33376 24750
rect 33324 24686 33376 24692
rect 32772 24608 32824 24614
rect 32772 24550 32824 24556
rect 33048 24608 33100 24614
rect 33048 24550 33100 24556
rect 32680 23860 32732 23866
rect 32680 23802 32732 23808
rect 32496 23792 32548 23798
rect 32496 23734 32548 23740
rect 32588 23792 32640 23798
rect 32588 23734 32640 23740
rect 32600 23594 32628 23734
rect 32588 23588 32640 23594
rect 32588 23530 32640 23536
rect 32772 23588 32824 23594
rect 32772 23530 32824 23536
rect 32600 23186 32628 23530
rect 32588 23180 32640 23186
rect 32588 23122 32640 23128
rect 32404 22772 32456 22778
rect 32404 22714 32456 22720
rect 32312 22636 32364 22642
rect 32312 22578 32364 22584
rect 32220 22160 32272 22166
rect 32220 22102 32272 22108
rect 32128 22092 32180 22098
rect 32128 22034 32180 22040
rect 32140 21842 32168 22034
rect 32140 21814 32260 21842
rect 32232 21146 32260 21814
rect 32324 21554 32352 22578
rect 32416 22574 32444 22714
rect 32404 22568 32456 22574
rect 32404 22510 32456 22516
rect 32496 22568 32548 22574
rect 32496 22510 32548 22516
rect 32312 21548 32364 21554
rect 32312 21490 32364 21496
rect 32220 21140 32272 21146
rect 32220 21082 32272 21088
rect 32128 20936 32180 20942
rect 32128 20878 32180 20884
rect 32140 20466 32168 20878
rect 32128 20460 32180 20466
rect 32128 20402 32180 20408
rect 32140 19854 32168 20402
rect 32232 20210 32260 21082
rect 32312 21004 32364 21010
rect 32312 20946 32364 20952
rect 32324 20330 32352 20946
rect 32312 20324 32364 20330
rect 32312 20266 32364 20272
rect 32232 20182 32352 20210
rect 32220 19916 32272 19922
rect 32220 19858 32272 19864
rect 32128 19848 32180 19854
rect 32128 19790 32180 19796
rect 32036 19780 32088 19786
rect 32036 19722 32088 19728
rect 32048 17202 32076 19722
rect 32232 19514 32260 19858
rect 32220 19508 32272 19514
rect 32220 19450 32272 19456
rect 32126 19408 32182 19417
rect 32126 19343 32182 19352
rect 32140 19174 32168 19343
rect 32220 19304 32272 19310
rect 32324 19292 32352 20182
rect 32508 19446 32536 22510
rect 32784 22098 32812 23530
rect 33060 23474 33088 24550
rect 33336 24274 33364 24686
rect 33324 24268 33376 24274
rect 33324 24210 33376 24216
rect 33140 24132 33192 24138
rect 33140 24074 33192 24080
rect 33152 23730 33180 24074
rect 33140 23724 33192 23730
rect 33140 23666 33192 23672
rect 33232 23656 33284 23662
rect 33232 23598 33284 23604
rect 33060 23446 33180 23474
rect 33152 22114 33180 23446
rect 33244 23118 33272 23598
rect 33692 23316 33744 23322
rect 33692 23258 33744 23264
rect 33508 23180 33560 23186
rect 33508 23122 33560 23128
rect 33232 23112 33284 23118
rect 33232 23054 33284 23060
rect 33244 22234 33272 23054
rect 33324 23044 33376 23050
rect 33324 22986 33376 22992
rect 33232 22228 33284 22234
rect 33232 22170 33284 22176
rect 32772 22092 32824 22098
rect 33152 22086 33272 22114
rect 32772 22034 32824 22040
rect 32956 21548 33008 21554
rect 32956 21490 33008 21496
rect 32968 21078 32996 21490
rect 33244 21486 33272 22086
rect 33232 21480 33284 21486
rect 33232 21422 33284 21428
rect 33048 21344 33100 21350
rect 33048 21286 33100 21292
rect 32956 21072 33008 21078
rect 32956 21014 33008 21020
rect 32864 20392 32916 20398
rect 32864 20334 32916 20340
rect 32496 19440 32548 19446
rect 32496 19382 32548 19388
rect 32876 19378 32904 20334
rect 32864 19372 32916 19378
rect 32864 19314 32916 19320
rect 32272 19264 32352 19292
rect 32220 19246 32272 19252
rect 32128 19168 32180 19174
rect 32128 19110 32180 19116
rect 32036 17196 32088 17202
rect 32036 17138 32088 17144
rect 32128 16992 32180 16998
rect 32128 16934 32180 16940
rect 32036 15564 32088 15570
rect 32036 15506 32088 15512
rect 31944 15496 31996 15502
rect 31944 15438 31996 15444
rect 31760 13864 31812 13870
rect 31760 13806 31812 13812
rect 31668 13796 31720 13802
rect 31668 13738 31720 13744
rect 31680 12646 31708 13738
rect 31772 12782 31800 13806
rect 32048 13326 32076 15506
rect 32140 14482 32168 16934
rect 32232 16658 32260 19246
rect 32876 18902 32904 19314
rect 32864 18896 32916 18902
rect 32864 18838 32916 18844
rect 32956 18896 33008 18902
rect 32956 18838 33008 18844
rect 32588 18828 32640 18834
rect 32588 18770 32640 18776
rect 32496 18692 32548 18698
rect 32496 18634 32548 18640
rect 32312 18352 32364 18358
rect 32310 18320 32312 18329
rect 32364 18320 32366 18329
rect 32310 18255 32366 18264
rect 32324 17746 32352 18255
rect 32508 18222 32536 18634
rect 32496 18216 32548 18222
rect 32496 18158 32548 18164
rect 32600 17882 32628 18770
rect 32680 18352 32732 18358
rect 32680 18294 32732 18300
rect 32588 17876 32640 17882
rect 32588 17818 32640 17824
rect 32312 17740 32364 17746
rect 32312 17682 32364 17688
rect 32220 16652 32272 16658
rect 32220 16594 32272 16600
rect 32324 16114 32352 17682
rect 32600 17270 32628 17818
rect 32692 17746 32720 18294
rect 32968 18154 32996 18838
rect 33060 18834 33088 21286
rect 33140 20868 33192 20874
rect 33140 20810 33192 20816
rect 33152 20466 33180 20810
rect 33140 20460 33192 20466
rect 33140 20402 33192 20408
rect 33336 19394 33364 22986
rect 33520 22098 33548 23122
rect 33600 22568 33652 22574
rect 33600 22510 33652 22516
rect 33508 22092 33560 22098
rect 33508 22034 33560 22040
rect 33612 21962 33640 22510
rect 33704 22166 33732 23258
rect 33784 22432 33836 22438
rect 33784 22374 33836 22380
rect 33692 22160 33744 22166
rect 33692 22102 33744 22108
rect 33600 21956 33652 21962
rect 33600 21898 33652 21904
rect 33612 21570 33640 21898
rect 33520 21542 33640 21570
rect 33416 20936 33468 20942
rect 33416 20878 33468 20884
rect 33428 19854 33456 20878
rect 33520 20398 33548 21542
rect 33704 21010 33732 22102
rect 33796 22030 33824 22374
rect 33784 22024 33836 22030
rect 33784 21966 33836 21972
rect 33692 21004 33744 21010
rect 33692 20946 33744 20952
rect 33508 20392 33560 20398
rect 33508 20334 33560 20340
rect 33416 19848 33468 19854
rect 33416 19790 33468 19796
rect 33336 19366 33456 19394
rect 33140 19304 33192 19310
rect 33140 19246 33192 19252
rect 33324 19304 33376 19310
rect 33324 19246 33376 19252
rect 33152 19145 33180 19246
rect 33138 19136 33194 19145
rect 33138 19071 33194 19080
rect 33048 18828 33100 18834
rect 33048 18770 33100 18776
rect 33336 18290 33364 19246
rect 33324 18284 33376 18290
rect 33324 18226 33376 18232
rect 33048 18216 33100 18222
rect 33048 18158 33100 18164
rect 33232 18216 33284 18222
rect 33232 18158 33284 18164
rect 32956 18148 33008 18154
rect 32956 18090 33008 18096
rect 32680 17740 32732 17746
rect 32680 17682 32732 17688
rect 32772 17536 32824 17542
rect 32772 17478 32824 17484
rect 32784 17338 32812 17478
rect 32968 17338 32996 18090
rect 32772 17332 32824 17338
rect 32772 17274 32824 17280
rect 32956 17332 33008 17338
rect 32956 17274 33008 17280
rect 32588 17264 32640 17270
rect 32588 17206 32640 17212
rect 33060 17202 33088 18158
rect 33048 17196 33100 17202
rect 33048 17138 33100 17144
rect 32404 16652 32456 16658
rect 32404 16594 32456 16600
rect 32312 16108 32364 16114
rect 32312 16050 32364 16056
rect 32416 16046 32444 16594
rect 32404 16040 32456 16046
rect 32404 15982 32456 15988
rect 32220 15904 32272 15910
rect 32220 15846 32272 15852
rect 32232 15434 32260 15846
rect 32772 15564 32824 15570
rect 32772 15506 32824 15512
rect 32312 15496 32364 15502
rect 32312 15438 32364 15444
rect 32220 15428 32272 15434
rect 32220 15370 32272 15376
rect 32232 14890 32260 15370
rect 32324 14958 32352 15438
rect 32784 14958 32812 15506
rect 33244 15162 33272 18158
rect 33428 16794 33456 19366
rect 33784 18896 33836 18902
rect 33784 18838 33836 18844
rect 33508 18760 33560 18766
rect 33508 18702 33560 18708
rect 33520 18222 33548 18702
rect 33690 18320 33746 18329
rect 33690 18255 33746 18264
rect 33508 18216 33560 18222
rect 33508 18158 33560 18164
rect 33520 17882 33548 18158
rect 33508 17876 33560 17882
rect 33508 17818 33560 17824
rect 33416 16788 33468 16794
rect 33416 16730 33468 16736
rect 33324 15428 33376 15434
rect 33324 15370 33376 15376
rect 33232 15156 33284 15162
rect 33232 15098 33284 15104
rect 33048 15020 33100 15026
rect 33048 14962 33100 14968
rect 32312 14952 32364 14958
rect 32312 14894 32364 14900
rect 32772 14952 32824 14958
rect 32772 14894 32824 14900
rect 32220 14884 32272 14890
rect 32220 14826 32272 14832
rect 32128 14476 32180 14482
rect 32128 14418 32180 14424
rect 32036 13320 32088 13326
rect 32036 13262 32088 13268
rect 32036 12980 32088 12986
rect 32036 12922 32088 12928
rect 31760 12776 31812 12782
rect 31760 12718 31812 12724
rect 31852 12708 31904 12714
rect 31852 12650 31904 12656
rect 31668 12640 31720 12646
rect 31668 12582 31720 12588
rect 31680 11830 31708 12582
rect 31864 11898 31892 12650
rect 31852 11892 31904 11898
rect 31852 11834 31904 11840
rect 31668 11824 31720 11830
rect 31668 11766 31720 11772
rect 31576 10532 31628 10538
rect 31576 10474 31628 10480
rect 31588 9518 31616 10474
rect 32048 9654 32076 12922
rect 32140 12306 32168 14418
rect 32128 12300 32180 12306
rect 32128 12242 32180 12248
rect 32128 11212 32180 11218
rect 32128 11154 32180 11160
rect 32036 9648 32088 9654
rect 31850 9616 31906 9625
rect 32036 9590 32088 9596
rect 31850 9551 31906 9560
rect 31864 9518 31892 9551
rect 31576 9512 31628 9518
rect 31576 9454 31628 9460
rect 31852 9512 31904 9518
rect 31852 9454 31904 9460
rect 31300 9376 31352 9382
rect 31300 9318 31352 9324
rect 31392 9376 31444 9382
rect 31392 9318 31444 9324
rect 31116 9036 31168 9042
rect 31116 8978 31168 8984
rect 31312 8838 31340 9318
rect 31300 8832 31352 8838
rect 31300 8774 31352 8780
rect 31404 8498 31432 9318
rect 32048 8974 32076 9590
rect 32036 8968 32088 8974
rect 32036 8910 32088 8916
rect 31574 8528 31630 8537
rect 31392 8492 31444 8498
rect 31574 8463 31630 8472
rect 31392 8434 31444 8440
rect 31588 8430 31616 8463
rect 31576 8424 31628 8430
rect 31576 8366 31628 8372
rect 31024 8084 31076 8090
rect 31024 8026 31076 8032
rect 31116 7948 31168 7954
rect 31116 7890 31168 7896
rect 30932 7744 30984 7750
rect 30932 7686 30984 7692
rect 31128 7546 31156 7890
rect 31392 7880 31444 7886
rect 31392 7822 31444 7828
rect 31404 7546 31432 7822
rect 31760 7812 31812 7818
rect 31760 7754 31812 7760
rect 31116 7540 31168 7546
rect 31116 7482 31168 7488
rect 31392 7540 31444 7546
rect 31392 7482 31444 7488
rect 30288 7336 30340 7342
rect 30288 7278 30340 7284
rect 30300 6254 30328 7278
rect 31484 6860 31536 6866
rect 31484 6802 31536 6808
rect 30840 6792 30892 6798
rect 30840 6734 30892 6740
rect 30392 6446 30604 6474
rect 30196 6248 30248 6254
rect 30196 6190 30248 6196
rect 30288 6248 30340 6254
rect 30288 6190 30340 6196
rect 30392 6186 30420 6446
rect 30380 6180 30432 6186
rect 30380 6122 30432 6128
rect 30380 5772 30432 5778
rect 30380 5714 30432 5720
rect 29932 4814 30052 4842
rect 29932 3369 29960 4814
rect 30392 4622 30420 5714
rect 30576 5710 30604 6446
rect 30852 5778 30880 6734
rect 31208 6656 31260 6662
rect 31208 6598 31260 6604
rect 31392 6656 31444 6662
rect 31392 6598 31444 6604
rect 31220 6474 31248 6598
rect 31220 6446 31340 6474
rect 31312 6390 31340 6446
rect 31300 6384 31352 6390
rect 31300 6326 31352 6332
rect 31312 5778 31340 6326
rect 31404 6322 31432 6598
rect 31496 6458 31524 6802
rect 31484 6452 31536 6458
rect 31484 6394 31536 6400
rect 31392 6316 31444 6322
rect 31392 6258 31444 6264
rect 30840 5772 30892 5778
rect 30840 5714 30892 5720
rect 31300 5772 31352 5778
rect 31300 5714 31352 5720
rect 30564 5704 30616 5710
rect 30564 5646 30616 5652
rect 31404 5234 31432 6258
rect 31484 5704 31536 5710
rect 31484 5646 31536 5652
rect 31668 5704 31720 5710
rect 31668 5646 31720 5652
rect 30564 5228 30616 5234
rect 30564 5170 30616 5176
rect 31392 5228 31444 5234
rect 31392 5170 31444 5176
rect 30380 4616 30432 4622
rect 30380 4558 30432 4564
rect 30012 4480 30064 4486
rect 30012 4422 30064 4428
rect 29918 3360 29974 3369
rect 29918 3295 29974 3304
rect 29828 3052 29880 3058
rect 29828 2994 29880 3000
rect 29828 2916 29880 2922
rect 29828 2858 29880 2864
rect 29840 2582 29868 2858
rect 29828 2576 29880 2582
rect 29828 2518 29880 2524
rect 30024 2514 30052 4422
rect 30392 4146 30420 4558
rect 30576 4146 30604 5170
rect 31496 5098 31524 5646
rect 31484 5092 31536 5098
rect 31484 5034 31536 5040
rect 31680 4622 31708 5646
rect 31772 5370 31800 7754
rect 32140 7478 32168 11154
rect 32232 10606 32260 14826
rect 32324 13530 32352 14894
rect 32784 14346 32812 14894
rect 32772 14340 32824 14346
rect 32772 14282 32824 14288
rect 32588 14272 32640 14278
rect 32588 14214 32640 14220
rect 32496 13864 32548 13870
rect 32496 13806 32548 13812
rect 32312 13524 32364 13530
rect 32312 13466 32364 13472
rect 32324 13410 32352 13466
rect 32324 13382 32444 13410
rect 32312 13320 32364 13326
rect 32312 13262 32364 13268
rect 32324 12442 32352 13262
rect 32312 12436 32364 12442
rect 32312 12378 32364 12384
rect 32312 11688 32364 11694
rect 32312 11630 32364 11636
rect 32324 11354 32352 11630
rect 32416 11626 32444 13382
rect 32508 12986 32536 13806
rect 32496 12980 32548 12986
rect 32496 12922 32548 12928
rect 32496 12776 32548 12782
rect 32496 12718 32548 12724
rect 32404 11620 32456 11626
rect 32404 11562 32456 11568
rect 32312 11348 32364 11354
rect 32312 11290 32364 11296
rect 32312 11212 32364 11218
rect 32312 11154 32364 11160
rect 32220 10600 32272 10606
rect 32220 10542 32272 10548
rect 32220 10124 32272 10130
rect 32220 10066 32272 10072
rect 32232 9926 32260 10066
rect 32220 9920 32272 9926
rect 32220 9862 32272 9868
rect 32324 9586 32352 11154
rect 32508 10606 32536 12718
rect 32600 11218 32628 14214
rect 32680 12844 32732 12850
rect 32680 12786 32732 12792
rect 32692 12306 32720 12786
rect 32680 12300 32732 12306
rect 32680 12242 32732 12248
rect 32772 11688 32824 11694
rect 32772 11630 32824 11636
rect 32588 11212 32640 11218
rect 32588 11154 32640 11160
rect 32784 11150 32812 11630
rect 32956 11280 33008 11286
rect 32956 11222 33008 11228
rect 32772 11144 32824 11150
rect 32772 11086 32824 11092
rect 32588 11076 32640 11082
rect 32588 11018 32640 11024
rect 32496 10600 32548 10606
rect 32496 10542 32548 10548
rect 32404 9920 32456 9926
rect 32404 9862 32456 9868
rect 32312 9580 32364 9586
rect 32312 9522 32364 9528
rect 32312 8356 32364 8362
rect 32312 8298 32364 8304
rect 32324 7886 32352 8298
rect 32312 7880 32364 7886
rect 32312 7822 32364 7828
rect 32128 7472 32180 7478
rect 32128 7414 32180 7420
rect 32416 7410 32444 9862
rect 32508 7954 32536 10542
rect 32600 8906 32628 11018
rect 32772 10668 32824 10674
rect 32772 10610 32824 10616
rect 32680 10600 32732 10606
rect 32680 10542 32732 10548
rect 32692 9654 32720 10542
rect 32680 9648 32732 9654
rect 32680 9590 32732 9596
rect 32784 9518 32812 10610
rect 32864 10600 32916 10606
rect 32864 10542 32916 10548
rect 32772 9512 32824 9518
rect 32772 9454 32824 9460
rect 32876 9042 32904 10542
rect 32968 10062 32996 11222
rect 33060 11218 33088 14962
rect 33336 14414 33364 15370
rect 33324 14408 33376 14414
rect 33324 14350 33376 14356
rect 33232 14272 33284 14278
rect 33232 14214 33284 14220
rect 33244 13870 33272 14214
rect 33336 13870 33364 14350
rect 33428 14074 33456 16730
rect 33704 16658 33732 18255
rect 33796 17134 33824 18838
rect 33888 18086 33916 25774
rect 33968 25696 34020 25702
rect 33968 25638 34020 25644
rect 33980 25226 34008 25638
rect 34060 25492 34112 25498
rect 34060 25434 34112 25440
rect 33968 25220 34020 25226
rect 33968 25162 34020 25168
rect 34072 24750 34100 25434
rect 34060 24744 34112 24750
rect 34060 24686 34112 24692
rect 33968 24200 34020 24206
rect 33968 24142 34020 24148
rect 33980 23798 34008 24142
rect 33968 23792 34020 23798
rect 33968 23734 34020 23740
rect 33980 23322 34008 23734
rect 34072 23526 34100 24686
rect 34244 24200 34296 24206
rect 34244 24142 34296 24148
rect 34152 23656 34204 23662
rect 34152 23598 34204 23604
rect 34060 23520 34112 23526
rect 34060 23462 34112 23468
rect 33968 23316 34020 23322
rect 33968 23258 34020 23264
rect 34072 23202 34100 23462
rect 33980 23174 34100 23202
rect 33980 22506 34008 23174
rect 34060 22636 34112 22642
rect 34060 22578 34112 22584
rect 33968 22500 34020 22506
rect 33968 22442 34020 22448
rect 33980 21554 34008 22442
rect 33968 21548 34020 21554
rect 33968 21490 34020 21496
rect 34072 21468 34100 22578
rect 34164 21690 34192 23598
rect 34256 23254 34284 24142
rect 34244 23248 34296 23254
rect 34244 23190 34296 23196
rect 34440 22642 34468 28630
rect 34520 28416 34572 28422
rect 34520 28358 34572 28364
rect 34532 27606 34560 28358
rect 34520 27600 34572 27606
rect 34520 27542 34572 27548
rect 34716 23866 34744 31758
rect 34808 30734 34836 34002
rect 34940 33756 35236 33776
rect 34996 33754 35020 33756
rect 35076 33754 35100 33756
rect 35156 33754 35180 33756
rect 35018 33702 35020 33754
rect 35082 33702 35094 33754
rect 35156 33702 35158 33754
rect 34996 33700 35020 33702
rect 35076 33700 35100 33702
rect 35156 33700 35180 33702
rect 34940 33680 35236 33700
rect 35360 33046 35388 34342
rect 35452 34066 35480 34546
rect 35440 34060 35492 34066
rect 35440 34002 35492 34008
rect 35348 33040 35400 33046
rect 35348 32982 35400 32988
rect 34940 32668 35236 32688
rect 34996 32666 35020 32668
rect 35076 32666 35100 32668
rect 35156 32666 35180 32668
rect 35018 32614 35020 32666
rect 35082 32614 35094 32666
rect 35156 32614 35158 32666
rect 34996 32612 35020 32614
rect 35076 32612 35100 32614
rect 35156 32612 35180 32614
rect 34940 32592 35236 32612
rect 35348 32496 35400 32502
rect 35348 32438 35400 32444
rect 35256 31816 35308 31822
rect 35256 31758 35308 31764
rect 34940 31580 35236 31600
rect 34996 31578 35020 31580
rect 35076 31578 35100 31580
rect 35156 31578 35180 31580
rect 35018 31526 35020 31578
rect 35082 31526 35094 31578
rect 35156 31526 35158 31578
rect 34996 31524 35020 31526
rect 35076 31524 35100 31526
rect 35156 31524 35180 31526
rect 34940 31504 35236 31524
rect 35164 31272 35216 31278
rect 35164 31214 35216 31220
rect 34796 30728 34848 30734
rect 34796 30670 34848 30676
rect 35176 30682 35204 31214
rect 35268 30938 35296 31758
rect 35256 30932 35308 30938
rect 35256 30874 35308 30880
rect 35360 30802 35388 32438
rect 35544 31890 35572 37266
rect 37568 36718 37596 40200
rect 39408 38010 39436 40200
rect 39396 38004 39448 38010
rect 39396 37946 39448 37952
rect 38292 37664 38344 37670
rect 38292 37606 38344 37612
rect 37556 36712 37608 36718
rect 37556 36654 37608 36660
rect 35900 36236 35952 36242
rect 35900 36178 35952 36184
rect 35912 36009 35940 36178
rect 35898 36000 35954 36009
rect 35898 35935 35954 35944
rect 37924 35148 37976 35154
rect 37924 35090 37976 35096
rect 38200 35148 38252 35154
rect 38200 35090 38252 35096
rect 36084 34536 36136 34542
rect 36084 34478 36136 34484
rect 36360 34536 36412 34542
rect 36360 34478 36412 34484
rect 37372 34536 37424 34542
rect 37372 34478 37424 34484
rect 35716 34400 35768 34406
rect 35716 34342 35768 34348
rect 35728 34066 35756 34342
rect 35716 34060 35768 34066
rect 35716 34002 35768 34008
rect 35808 34060 35860 34066
rect 35808 34002 35860 34008
rect 35820 33590 35848 34002
rect 35808 33584 35860 33590
rect 35808 33526 35860 33532
rect 35808 33448 35860 33454
rect 35808 33390 35860 33396
rect 35820 32978 35848 33390
rect 35808 32972 35860 32978
rect 35808 32914 35860 32920
rect 35820 32366 35848 32914
rect 36096 32842 36124 34478
rect 36372 33318 36400 34478
rect 37384 34202 37412 34478
rect 37372 34196 37424 34202
rect 37372 34138 37424 34144
rect 37648 33992 37700 33998
rect 37648 33934 37700 33940
rect 36636 33856 36688 33862
rect 36636 33798 36688 33804
rect 36648 33454 36676 33798
rect 36636 33448 36688 33454
rect 36636 33390 36688 33396
rect 36360 33312 36412 33318
rect 36360 33254 36412 33260
rect 36452 32972 36504 32978
rect 36452 32914 36504 32920
rect 36268 32904 36320 32910
rect 36268 32846 36320 32852
rect 36084 32836 36136 32842
rect 36084 32778 36136 32784
rect 35808 32360 35860 32366
rect 35808 32302 35860 32308
rect 35532 31884 35584 31890
rect 35532 31826 35584 31832
rect 35440 31680 35492 31686
rect 35440 31622 35492 31628
rect 35452 31362 35480 31622
rect 35820 31482 35848 32302
rect 36280 32026 36308 32846
rect 36268 32020 36320 32026
rect 36268 31962 36320 31968
rect 35808 31476 35860 31482
rect 35808 31418 35860 31424
rect 35452 31334 35572 31362
rect 35544 31210 35572 31334
rect 35716 31340 35768 31346
rect 35716 31282 35768 31288
rect 35440 31204 35492 31210
rect 35440 31146 35492 31152
rect 35532 31204 35584 31210
rect 35532 31146 35584 31152
rect 35348 30796 35400 30802
rect 35348 30738 35400 30744
rect 35176 30654 35296 30682
rect 34940 30492 35236 30512
rect 34996 30490 35020 30492
rect 35076 30490 35100 30492
rect 35156 30490 35180 30492
rect 35018 30438 35020 30490
rect 35082 30438 35094 30490
rect 35156 30438 35158 30490
rect 34996 30436 35020 30438
rect 35076 30436 35100 30438
rect 35156 30436 35180 30438
rect 34940 30416 35236 30436
rect 34940 29404 35236 29424
rect 34996 29402 35020 29404
rect 35076 29402 35100 29404
rect 35156 29402 35180 29404
rect 35018 29350 35020 29402
rect 35082 29350 35094 29402
rect 35156 29350 35158 29402
rect 34996 29348 35020 29350
rect 35076 29348 35100 29350
rect 35156 29348 35180 29350
rect 34940 29328 35236 29348
rect 34796 28620 34848 28626
rect 34796 28562 34848 28568
rect 34808 27130 34836 28562
rect 34940 28316 35236 28336
rect 34996 28314 35020 28316
rect 35076 28314 35100 28316
rect 35156 28314 35180 28316
rect 35018 28262 35020 28314
rect 35082 28262 35094 28314
rect 35156 28262 35158 28314
rect 34996 28260 35020 28262
rect 35076 28260 35100 28262
rect 35156 28260 35180 28262
rect 34940 28240 35236 28260
rect 34940 27228 35236 27248
rect 34996 27226 35020 27228
rect 35076 27226 35100 27228
rect 35156 27226 35180 27228
rect 35018 27174 35020 27226
rect 35082 27174 35094 27226
rect 35156 27174 35158 27226
rect 34996 27172 35020 27174
rect 35076 27172 35100 27174
rect 35156 27172 35180 27174
rect 34940 27152 35236 27172
rect 34796 27124 34848 27130
rect 34796 27066 34848 27072
rect 35268 26926 35296 30654
rect 35452 29102 35480 31146
rect 35544 29714 35572 31146
rect 35728 30802 35756 31282
rect 35716 30796 35768 30802
rect 35716 30738 35768 30744
rect 35820 30190 35848 31418
rect 35992 31272 36044 31278
rect 35992 31214 36044 31220
rect 35624 30184 35676 30190
rect 35624 30126 35676 30132
rect 35808 30184 35860 30190
rect 35808 30126 35860 30132
rect 35532 29708 35584 29714
rect 35532 29650 35584 29656
rect 35440 29096 35492 29102
rect 35440 29038 35492 29044
rect 35636 29050 35664 30126
rect 35716 29640 35768 29646
rect 35716 29582 35768 29588
rect 35728 29238 35756 29582
rect 35716 29232 35768 29238
rect 35716 29174 35768 29180
rect 35636 29022 35756 29050
rect 35728 28626 35756 29022
rect 35716 28620 35768 28626
rect 35716 28562 35768 28568
rect 35808 28620 35860 28626
rect 35808 28562 35860 28568
rect 35728 28422 35756 28562
rect 35716 28416 35768 28422
rect 35716 28358 35768 28364
rect 35728 27538 35756 28358
rect 35820 27538 35848 28562
rect 35716 27532 35768 27538
rect 35716 27474 35768 27480
rect 35808 27532 35860 27538
rect 35808 27474 35860 27480
rect 35624 27124 35676 27130
rect 35624 27066 35676 27072
rect 35256 26920 35308 26926
rect 35256 26862 35308 26868
rect 35348 26376 35400 26382
rect 35348 26318 35400 26324
rect 34940 26140 35236 26160
rect 34996 26138 35020 26140
rect 35076 26138 35100 26140
rect 35156 26138 35180 26140
rect 35018 26086 35020 26138
rect 35082 26086 35094 26138
rect 35156 26086 35158 26138
rect 34996 26084 35020 26086
rect 35076 26084 35100 26086
rect 35156 26084 35180 26086
rect 34940 26064 35236 26084
rect 34940 25052 35236 25072
rect 34996 25050 35020 25052
rect 35076 25050 35100 25052
rect 35156 25050 35180 25052
rect 35018 24998 35020 25050
rect 35082 24998 35094 25050
rect 35156 24998 35158 25050
rect 34996 24996 35020 24998
rect 35076 24996 35100 24998
rect 35156 24996 35180 24998
rect 34940 24976 35236 24996
rect 35360 24750 35388 26318
rect 35440 25832 35492 25838
rect 35440 25774 35492 25780
rect 35452 25498 35480 25774
rect 35440 25492 35492 25498
rect 35440 25434 35492 25440
rect 35532 25356 35584 25362
rect 35532 25298 35584 25304
rect 35348 24744 35400 24750
rect 35348 24686 35400 24692
rect 35256 24676 35308 24682
rect 35256 24618 35308 24624
rect 34940 23964 35236 23984
rect 34996 23962 35020 23964
rect 35076 23962 35100 23964
rect 35156 23962 35180 23964
rect 35018 23910 35020 23962
rect 35082 23910 35094 23962
rect 35156 23910 35158 23962
rect 34996 23908 35020 23910
rect 35076 23908 35100 23910
rect 35156 23908 35180 23910
rect 34940 23888 35236 23908
rect 34520 23860 34572 23866
rect 34520 23802 34572 23808
rect 34704 23860 34756 23866
rect 34704 23802 34756 23808
rect 34428 22636 34480 22642
rect 34428 22578 34480 22584
rect 34428 22160 34480 22166
rect 34428 22102 34480 22108
rect 34440 22030 34468 22102
rect 34428 22024 34480 22030
rect 34428 21966 34480 21972
rect 34152 21684 34204 21690
rect 34152 21626 34204 21632
rect 34164 21570 34192 21626
rect 34336 21616 34388 21622
rect 34164 21542 34284 21570
rect 34336 21558 34388 21564
rect 34152 21480 34204 21486
rect 34072 21440 34152 21468
rect 34152 21422 34204 21428
rect 34060 21344 34112 21350
rect 34060 21286 34112 21292
rect 33968 19304 34020 19310
rect 33968 19246 34020 19252
rect 33980 18834 34008 19246
rect 33968 18828 34020 18834
rect 33968 18770 34020 18776
rect 33876 18080 33928 18086
rect 33876 18022 33928 18028
rect 33784 17128 33836 17134
rect 33784 17070 33836 17076
rect 33692 16652 33744 16658
rect 33692 16594 33744 16600
rect 33508 16040 33560 16046
rect 33508 15982 33560 15988
rect 33520 15706 33548 15982
rect 33508 15700 33560 15706
rect 33508 15642 33560 15648
rect 33600 15700 33652 15706
rect 33600 15642 33652 15648
rect 33612 14958 33640 15642
rect 33796 14958 33824 17070
rect 33888 16980 33916 18022
rect 34072 16998 34100 21286
rect 34164 21146 34192 21422
rect 34152 21140 34204 21146
rect 34152 21082 34204 21088
rect 34256 20806 34284 21542
rect 34244 20800 34296 20806
rect 34244 20742 34296 20748
rect 34244 20460 34296 20466
rect 34244 20402 34296 20408
rect 34256 19514 34284 20402
rect 34348 20058 34376 21558
rect 34336 20052 34388 20058
rect 34336 19994 34388 20000
rect 34428 19916 34480 19922
rect 34428 19858 34480 19864
rect 34244 19508 34296 19514
rect 34244 19450 34296 19456
rect 34152 19304 34204 19310
rect 34152 19246 34204 19252
rect 34164 18873 34192 19246
rect 34150 18864 34206 18873
rect 34150 18799 34206 18808
rect 34152 17672 34204 17678
rect 34152 17614 34204 17620
rect 34164 17134 34192 17614
rect 34152 17128 34204 17134
rect 34152 17070 34204 17076
rect 34060 16992 34112 16998
rect 33888 16952 34008 16980
rect 33600 14952 33652 14958
rect 33600 14894 33652 14900
rect 33784 14952 33836 14958
rect 33784 14894 33836 14900
rect 33876 14408 33928 14414
rect 33876 14350 33928 14356
rect 33416 14068 33468 14074
rect 33416 14010 33468 14016
rect 33232 13864 33284 13870
rect 33232 13806 33284 13812
rect 33324 13864 33376 13870
rect 33324 13806 33376 13812
rect 33244 12782 33272 13806
rect 33232 12776 33284 12782
rect 33232 12718 33284 12724
rect 33232 12232 33284 12238
rect 33232 12174 33284 12180
rect 33048 11212 33100 11218
rect 33048 11154 33100 11160
rect 33140 11008 33192 11014
rect 33140 10950 33192 10956
rect 33152 10266 33180 10950
rect 33244 10674 33272 12174
rect 33428 11694 33456 14010
rect 33888 13530 33916 14350
rect 33980 13530 34008 16952
rect 34060 16934 34112 16940
rect 34072 14414 34100 16934
rect 34336 15904 34388 15910
rect 34336 15846 34388 15852
rect 34348 15570 34376 15846
rect 34440 15706 34468 19858
rect 34532 19174 34560 23802
rect 35268 23186 35296 24618
rect 35440 24608 35492 24614
rect 35440 24550 35492 24556
rect 35256 23180 35308 23186
rect 35256 23122 35308 23128
rect 35268 23066 35296 23122
rect 35452 23118 35480 24550
rect 35440 23112 35492 23118
rect 35268 23038 35388 23066
rect 35440 23054 35492 23060
rect 34940 22876 35236 22896
rect 34996 22874 35020 22876
rect 35076 22874 35100 22876
rect 35156 22874 35180 22876
rect 35018 22822 35020 22874
rect 35082 22822 35094 22874
rect 35156 22822 35158 22874
rect 34996 22820 35020 22822
rect 35076 22820 35100 22822
rect 35156 22820 35180 22822
rect 34940 22800 35236 22820
rect 35256 22568 35308 22574
rect 35256 22510 35308 22516
rect 34940 21788 35236 21808
rect 34996 21786 35020 21788
rect 35076 21786 35100 21788
rect 35156 21786 35180 21788
rect 35018 21734 35020 21786
rect 35082 21734 35094 21786
rect 35156 21734 35158 21786
rect 34996 21732 35020 21734
rect 35076 21732 35100 21734
rect 35156 21732 35180 21734
rect 34940 21712 35236 21732
rect 35268 21078 35296 22510
rect 34796 21072 34848 21078
rect 34796 21014 34848 21020
rect 35256 21072 35308 21078
rect 35256 21014 35308 21020
rect 34808 20398 34836 21014
rect 34940 20700 35236 20720
rect 34996 20698 35020 20700
rect 35076 20698 35100 20700
rect 35156 20698 35180 20700
rect 35018 20646 35020 20698
rect 35082 20646 35094 20698
rect 35156 20646 35158 20698
rect 34996 20644 35020 20646
rect 35076 20644 35100 20646
rect 35156 20644 35180 20646
rect 34940 20624 35236 20644
rect 34796 20392 34848 20398
rect 34796 20334 34848 20340
rect 35256 20392 35308 20398
rect 35360 20380 35388 23038
rect 35452 22982 35480 23054
rect 35440 22976 35492 22982
rect 35440 22918 35492 22924
rect 35544 22710 35572 25298
rect 35636 24750 35664 27066
rect 35728 26382 35756 27474
rect 35716 26376 35768 26382
rect 35716 26318 35768 26324
rect 35624 24744 35676 24750
rect 35624 24686 35676 24692
rect 35532 22704 35584 22710
rect 35532 22646 35584 22652
rect 35532 22432 35584 22438
rect 35532 22374 35584 22380
rect 35440 22024 35492 22030
rect 35440 21966 35492 21972
rect 35452 21554 35480 21966
rect 35440 21548 35492 21554
rect 35440 21490 35492 21496
rect 35440 21140 35492 21146
rect 35440 21082 35492 21088
rect 35308 20352 35388 20380
rect 35256 20334 35308 20340
rect 34704 20256 34756 20262
rect 34704 20198 34756 20204
rect 34520 19168 34572 19174
rect 34520 19110 34572 19116
rect 34520 18828 34572 18834
rect 34520 18770 34572 18776
rect 34532 18154 34560 18770
rect 34520 18148 34572 18154
rect 34520 18090 34572 18096
rect 34716 17678 34744 20198
rect 34808 19378 34836 20334
rect 34940 19612 35236 19632
rect 34996 19610 35020 19612
rect 35076 19610 35100 19612
rect 35156 19610 35180 19612
rect 35018 19558 35020 19610
rect 35082 19558 35094 19610
rect 35156 19558 35158 19610
rect 34996 19556 35020 19558
rect 35076 19556 35100 19558
rect 35156 19556 35180 19558
rect 34940 19536 35236 19556
rect 35268 19514 35296 20334
rect 35256 19508 35308 19514
rect 35256 19450 35308 19456
rect 34796 19372 34848 19378
rect 34796 19314 34848 19320
rect 35452 18834 35480 21082
rect 35256 18828 35308 18834
rect 35256 18770 35308 18776
rect 35440 18828 35492 18834
rect 35440 18770 35492 18776
rect 34940 18524 35236 18544
rect 34996 18522 35020 18524
rect 35076 18522 35100 18524
rect 35156 18522 35180 18524
rect 35018 18470 35020 18522
rect 35082 18470 35094 18522
rect 35156 18470 35158 18522
rect 34996 18468 35020 18470
rect 35076 18468 35100 18470
rect 35156 18468 35180 18470
rect 34940 18448 35236 18468
rect 35268 18222 35296 18770
rect 35452 18222 35480 18770
rect 35256 18216 35308 18222
rect 35256 18158 35308 18164
rect 35440 18216 35492 18222
rect 35440 18158 35492 18164
rect 34796 17740 34848 17746
rect 34796 17682 34848 17688
rect 34704 17672 34756 17678
rect 34704 17614 34756 17620
rect 34612 16652 34664 16658
rect 34612 16594 34664 16600
rect 34624 16250 34652 16594
rect 34612 16244 34664 16250
rect 34612 16186 34664 16192
rect 34716 15978 34744 17614
rect 34808 17134 34836 17682
rect 34940 17436 35236 17456
rect 34996 17434 35020 17436
rect 35076 17434 35100 17436
rect 35156 17434 35180 17436
rect 35018 17382 35020 17434
rect 35082 17382 35094 17434
rect 35156 17382 35158 17434
rect 34996 17380 35020 17382
rect 35076 17380 35100 17382
rect 35156 17380 35180 17382
rect 34940 17360 35236 17380
rect 35452 17338 35480 18158
rect 35544 17746 35572 22374
rect 35624 21616 35676 21622
rect 35624 21558 35676 21564
rect 35532 17740 35584 17746
rect 35532 17682 35584 17688
rect 35440 17332 35492 17338
rect 35440 17274 35492 17280
rect 34796 17128 34848 17134
rect 34796 17070 34848 17076
rect 34808 16454 34836 17070
rect 34796 16448 34848 16454
rect 34796 16390 34848 16396
rect 34808 16114 34836 16390
rect 34940 16348 35236 16368
rect 34996 16346 35020 16348
rect 35076 16346 35100 16348
rect 35156 16346 35180 16348
rect 35018 16294 35020 16346
rect 35082 16294 35094 16346
rect 35156 16294 35158 16346
rect 34996 16292 35020 16294
rect 35076 16292 35100 16294
rect 35156 16292 35180 16294
rect 34940 16272 35236 16292
rect 34796 16108 34848 16114
rect 34796 16050 34848 16056
rect 34704 15972 34756 15978
rect 34704 15914 34756 15920
rect 34428 15700 34480 15706
rect 34428 15642 34480 15648
rect 34336 15564 34388 15570
rect 34336 15506 34388 15512
rect 34520 15564 34572 15570
rect 34520 15506 34572 15512
rect 34348 14618 34376 15506
rect 34532 14822 34560 15506
rect 34940 15260 35236 15280
rect 34996 15258 35020 15260
rect 35076 15258 35100 15260
rect 35156 15258 35180 15260
rect 35018 15206 35020 15258
rect 35082 15206 35094 15258
rect 35156 15206 35158 15258
rect 34996 15204 35020 15206
rect 35076 15204 35100 15206
rect 35156 15204 35180 15206
rect 34940 15184 35236 15204
rect 34520 14816 34572 14822
rect 34520 14758 34572 14764
rect 34336 14612 34388 14618
rect 34336 14554 34388 14560
rect 34060 14408 34112 14414
rect 34060 14350 34112 14356
rect 33876 13524 33928 13530
rect 33876 13466 33928 13472
rect 33968 13524 34020 13530
rect 33968 13466 34020 13472
rect 34072 13462 34100 14350
rect 34152 13932 34204 13938
rect 34152 13874 34204 13880
rect 34060 13456 34112 13462
rect 34060 13398 34112 13404
rect 34164 13394 34192 13874
rect 34348 13870 34376 14554
rect 34612 14476 34664 14482
rect 34612 14418 34664 14424
rect 35532 14476 35584 14482
rect 35532 14418 35584 14424
rect 34336 13864 34388 13870
rect 34336 13806 34388 13812
rect 33692 13388 33744 13394
rect 33692 13330 33744 13336
rect 34152 13388 34204 13394
rect 34152 13330 34204 13336
rect 33704 11898 33732 13330
rect 34060 12776 34112 12782
rect 34060 12718 34112 12724
rect 34072 12306 34100 12718
rect 34244 12708 34296 12714
rect 34244 12650 34296 12656
rect 34060 12300 34112 12306
rect 34060 12242 34112 12248
rect 33692 11892 33744 11898
rect 33692 11834 33744 11840
rect 34072 11762 34100 12242
rect 34256 11762 34284 12650
rect 34520 12232 34572 12238
rect 34624 12186 34652 14418
rect 34940 14172 35236 14192
rect 34996 14170 35020 14172
rect 35076 14170 35100 14172
rect 35156 14170 35180 14172
rect 35018 14118 35020 14170
rect 35082 14118 35094 14170
rect 35156 14118 35158 14170
rect 34996 14116 35020 14118
rect 35076 14116 35100 14118
rect 35156 14116 35180 14118
rect 34940 14096 35236 14116
rect 34704 14000 34756 14006
rect 34704 13942 34756 13948
rect 34572 12180 34652 12186
rect 34520 12174 34652 12180
rect 34532 12158 34652 12174
rect 34060 11756 34112 11762
rect 34060 11698 34112 11704
rect 34244 11756 34296 11762
rect 34244 11698 34296 11704
rect 33416 11688 33468 11694
rect 33416 11630 33468 11636
rect 33692 11688 33744 11694
rect 33692 11630 33744 11636
rect 33600 11348 33652 11354
rect 33600 11290 33652 11296
rect 33324 10804 33376 10810
rect 33324 10746 33376 10752
rect 33232 10668 33284 10674
rect 33232 10610 33284 10616
rect 33336 10266 33364 10746
rect 33612 10470 33640 11290
rect 33704 11218 33732 11630
rect 33692 11212 33744 11218
rect 33692 11154 33744 11160
rect 33784 11212 33836 11218
rect 33784 11154 33836 11160
rect 33600 10464 33652 10470
rect 33600 10406 33652 10412
rect 33140 10260 33192 10266
rect 33140 10202 33192 10208
rect 33324 10260 33376 10266
rect 33324 10202 33376 10208
rect 32956 10056 33008 10062
rect 32956 9998 33008 10004
rect 33416 10056 33468 10062
rect 33416 9998 33468 10004
rect 32864 9036 32916 9042
rect 32864 8978 32916 8984
rect 32588 8900 32640 8906
rect 32588 8842 32640 8848
rect 32588 8424 32640 8430
rect 32588 8366 32640 8372
rect 32496 7948 32548 7954
rect 32496 7890 32548 7896
rect 32404 7404 32456 7410
rect 32404 7346 32456 7352
rect 32600 6866 32628 8366
rect 32968 7886 32996 9998
rect 33428 9722 33456 9998
rect 33416 9716 33468 9722
rect 33416 9658 33468 9664
rect 33612 9518 33640 10406
rect 33796 9518 33824 11154
rect 34624 11150 34652 12158
rect 34612 11144 34664 11150
rect 34612 11086 34664 11092
rect 33968 11076 34020 11082
rect 33968 11018 34020 11024
rect 33980 10130 34008 11018
rect 34336 11008 34388 11014
rect 34336 10950 34388 10956
rect 33968 10124 34020 10130
rect 33968 10066 34020 10072
rect 33600 9512 33652 9518
rect 33600 9454 33652 9460
rect 33784 9512 33836 9518
rect 33784 9454 33836 9460
rect 33138 9072 33194 9081
rect 34348 9042 34376 10950
rect 34716 10130 34744 13942
rect 35544 13938 35572 14418
rect 35532 13932 35584 13938
rect 35532 13874 35584 13880
rect 34940 13084 35236 13104
rect 34996 13082 35020 13084
rect 35076 13082 35100 13084
rect 35156 13082 35180 13084
rect 35018 13030 35020 13082
rect 35082 13030 35094 13082
rect 35156 13030 35158 13082
rect 34996 13028 35020 13030
rect 35076 13028 35100 13030
rect 35156 13028 35180 13030
rect 34940 13008 35236 13028
rect 35256 12776 35308 12782
rect 35256 12718 35308 12724
rect 34796 12232 34848 12238
rect 34796 12174 34848 12180
rect 34808 11830 34836 12174
rect 34940 11996 35236 12016
rect 34996 11994 35020 11996
rect 35076 11994 35100 11996
rect 35156 11994 35180 11996
rect 35018 11942 35020 11994
rect 35082 11942 35094 11994
rect 35156 11942 35158 11994
rect 34996 11940 35020 11942
rect 35076 11940 35100 11942
rect 35156 11940 35180 11942
rect 34940 11920 35236 11940
rect 34796 11824 34848 11830
rect 34796 11766 34848 11772
rect 35268 11762 35296 12718
rect 35256 11756 35308 11762
rect 35256 11698 35308 11704
rect 34796 11688 34848 11694
rect 34796 11630 34848 11636
rect 34808 10810 34836 11630
rect 34940 10908 35236 10928
rect 34996 10906 35020 10908
rect 35076 10906 35100 10908
rect 35156 10906 35180 10908
rect 35018 10854 35020 10906
rect 35082 10854 35094 10906
rect 35156 10854 35158 10906
rect 34996 10852 35020 10854
rect 35076 10852 35100 10854
rect 35156 10852 35180 10854
rect 34940 10832 35236 10852
rect 34796 10804 34848 10810
rect 34796 10746 34848 10752
rect 34704 10124 34756 10130
rect 34704 10066 34756 10072
rect 34940 9820 35236 9840
rect 34996 9818 35020 9820
rect 35076 9818 35100 9820
rect 35156 9818 35180 9820
rect 35018 9766 35020 9818
rect 35082 9766 35094 9818
rect 35156 9766 35158 9818
rect 34996 9764 35020 9766
rect 35076 9764 35100 9766
rect 35156 9764 35180 9766
rect 34940 9744 35236 9764
rect 35636 9636 35664 21558
rect 35728 21026 35756 26318
rect 35820 25702 35848 27474
rect 35900 27396 35952 27402
rect 35900 27338 35952 27344
rect 35912 26926 35940 27338
rect 35900 26920 35952 26926
rect 35900 26862 35952 26868
rect 36004 26450 36032 31214
rect 36280 30870 36308 31962
rect 36464 31278 36492 32914
rect 36648 32366 36676 33390
rect 36728 33380 36780 33386
rect 36728 33322 36780 33328
rect 36740 32978 36768 33322
rect 37660 33318 37688 33934
rect 37648 33312 37700 33318
rect 37648 33254 37700 33260
rect 36728 32972 36780 32978
rect 36728 32914 36780 32920
rect 36912 32972 36964 32978
rect 36912 32914 36964 32920
rect 36924 32434 36952 32914
rect 37462 32464 37518 32473
rect 36912 32428 36964 32434
rect 37462 32399 37518 32408
rect 36912 32370 36964 32376
rect 37476 32366 37504 32399
rect 36636 32360 36688 32366
rect 36636 32302 36688 32308
rect 37464 32360 37516 32366
rect 37464 32302 37516 32308
rect 36544 32292 36596 32298
rect 36544 32234 36596 32240
rect 36452 31272 36504 31278
rect 36452 31214 36504 31220
rect 36268 30864 36320 30870
rect 36556 30818 36584 32234
rect 36636 31272 36688 31278
rect 36636 31214 36688 31220
rect 36820 31272 36872 31278
rect 36820 31214 36872 31220
rect 36268 30806 36320 30812
rect 36464 30802 36584 30818
rect 36452 30796 36584 30802
rect 36504 30790 36584 30796
rect 36452 30738 36504 30744
rect 36360 30728 36412 30734
rect 36360 30670 36412 30676
rect 36268 29844 36320 29850
rect 36372 29832 36400 30670
rect 36464 30122 36492 30738
rect 36452 30116 36504 30122
rect 36452 30058 36504 30064
rect 36320 29804 36400 29832
rect 36268 29786 36320 29792
rect 36176 29504 36228 29510
rect 36176 29446 36228 29452
rect 36188 29102 36216 29446
rect 36372 29186 36400 29804
rect 36464 29306 36492 30058
rect 36648 29782 36676 31214
rect 36832 30938 36860 31214
rect 36820 30932 36872 30938
rect 36820 30874 36872 30880
rect 36912 30796 36964 30802
rect 36912 30738 36964 30744
rect 36924 30326 36952 30738
rect 36912 30320 36964 30326
rect 36912 30262 36964 30268
rect 37476 30258 37504 32302
rect 37660 30734 37688 33254
rect 37936 33046 37964 35090
rect 38108 34944 38160 34950
rect 38108 34886 38160 34892
rect 38016 34604 38068 34610
rect 38016 34546 38068 34552
rect 37924 33040 37976 33046
rect 37924 32982 37976 32988
rect 37936 32434 37964 32982
rect 37924 32428 37976 32434
rect 37924 32370 37976 32376
rect 37740 32360 37792 32366
rect 37740 32302 37792 32308
rect 37752 32065 37780 32302
rect 37738 32056 37794 32065
rect 37738 31991 37794 32000
rect 38028 31890 38056 34546
rect 38120 33454 38148 34886
rect 38212 34610 38240 35090
rect 38200 34604 38252 34610
rect 38200 34546 38252 34552
rect 38304 34490 38332 37606
rect 38212 34462 38332 34490
rect 38108 33448 38160 33454
rect 38108 33390 38160 33396
rect 38016 31884 38068 31890
rect 38016 31826 38068 31832
rect 37740 31272 37792 31278
rect 37740 31214 37792 31220
rect 37752 30938 37780 31214
rect 38108 31136 38160 31142
rect 38108 31078 38160 31084
rect 37740 30932 37792 30938
rect 37740 30874 37792 30880
rect 37648 30728 37700 30734
rect 37648 30670 37700 30676
rect 37832 30728 37884 30734
rect 37832 30670 37884 30676
rect 37464 30252 37516 30258
rect 37464 30194 37516 30200
rect 36912 30184 36964 30190
rect 36912 30126 36964 30132
rect 37372 30184 37424 30190
rect 37372 30126 37424 30132
rect 36636 29776 36688 29782
rect 36636 29718 36688 29724
rect 36924 29510 36952 30126
rect 36912 29504 36964 29510
rect 36912 29446 36964 29452
rect 36452 29300 36504 29306
rect 36452 29242 36504 29248
rect 36372 29170 36492 29186
rect 36372 29164 36504 29170
rect 36372 29158 36452 29164
rect 36452 29106 36504 29112
rect 36176 29096 36228 29102
rect 36176 29038 36228 29044
rect 36360 29096 36412 29102
rect 36360 29038 36412 29044
rect 36372 28694 36400 29038
rect 36360 28688 36412 28694
rect 36360 28630 36412 28636
rect 36084 28008 36136 28014
rect 36084 27950 36136 27956
rect 36096 27062 36124 27950
rect 36084 27056 36136 27062
rect 36084 26998 36136 27004
rect 35992 26444 36044 26450
rect 35992 26386 36044 26392
rect 36268 26444 36320 26450
rect 36268 26386 36320 26392
rect 36084 26240 36136 26246
rect 36084 26182 36136 26188
rect 35808 25696 35860 25702
rect 35808 25638 35860 25644
rect 36096 25362 36124 26182
rect 36280 26042 36308 26386
rect 36268 26036 36320 26042
rect 36268 25978 36320 25984
rect 36084 25356 36136 25362
rect 36084 25298 36136 25304
rect 35900 25288 35952 25294
rect 35900 25230 35952 25236
rect 35912 24818 35940 25230
rect 36084 25152 36136 25158
rect 36084 25094 36136 25100
rect 35900 24812 35952 24818
rect 35900 24754 35952 24760
rect 35808 24744 35860 24750
rect 35808 24686 35860 24692
rect 35820 21622 35848 24686
rect 35992 23656 36044 23662
rect 35992 23598 36044 23604
rect 36004 23322 36032 23598
rect 35992 23316 36044 23322
rect 35992 23258 36044 23264
rect 35808 21616 35860 21622
rect 35808 21558 35860 21564
rect 35808 21480 35860 21486
rect 35808 21422 35860 21428
rect 35992 21480 36044 21486
rect 35992 21422 36044 21428
rect 35820 21146 35848 21422
rect 35808 21140 35860 21146
rect 35808 21082 35860 21088
rect 35728 20998 35848 21026
rect 35820 19922 35848 20998
rect 35808 19916 35860 19922
rect 35808 19858 35860 19864
rect 35900 19848 35952 19854
rect 35900 19790 35952 19796
rect 35912 19145 35940 19790
rect 35898 19136 35954 19145
rect 35898 19071 35954 19080
rect 35716 18964 35768 18970
rect 35716 18906 35768 18912
rect 35728 17202 35756 18906
rect 35808 18216 35860 18222
rect 35808 18158 35860 18164
rect 35716 17196 35768 17202
rect 35716 17138 35768 17144
rect 35820 16046 35848 18158
rect 35912 17882 35940 19071
rect 35900 17876 35952 17882
rect 35900 17818 35952 17824
rect 35900 17740 35952 17746
rect 35900 17682 35952 17688
rect 35912 16658 35940 17682
rect 35900 16652 35952 16658
rect 35900 16594 35952 16600
rect 35912 16114 35940 16594
rect 35900 16108 35952 16114
rect 35900 16050 35952 16056
rect 35808 16040 35860 16046
rect 35808 15982 35860 15988
rect 35912 15706 35940 16050
rect 36004 16046 36032 21422
rect 36096 18873 36124 25094
rect 36464 24342 36492 29106
rect 36636 27396 36688 27402
rect 36636 27338 36688 27344
rect 36648 26926 36676 27338
rect 36636 26920 36688 26926
rect 36636 26862 36688 26868
rect 36924 24750 36952 29446
rect 37280 28008 37332 28014
rect 37280 27950 37332 27956
rect 37096 27600 37148 27606
rect 37096 27542 37148 27548
rect 37108 26858 37136 27542
rect 37096 26852 37148 26858
rect 37096 26794 37148 26800
rect 37108 25158 37136 26794
rect 37292 25906 37320 27950
rect 37280 25900 37332 25906
rect 37280 25842 37332 25848
rect 37096 25152 37148 25158
rect 37096 25094 37148 25100
rect 36912 24744 36964 24750
rect 36912 24686 36964 24692
rect 36268 24336 36320 24342
rect 36268 24278 36320 24284
rect 36452 24336 36504 24342
rect 36452 24278 36504 24284
rect 36176 22568 36228 22574
rect 36176 22510 36228 22516
rect 36188 21690 36216 22510
rect 36176 21684 36228 21690
rect 36176 21626 36228 21632
rect 36188 20398 36216 21626
rect 36280 21486 36308 24278
rect 36360 24268 36412 24274
rect 36360 24210 36412 24216
rect 36372 23526 36400 24210
rect 36452 24200 36504 24206
rect 36452 24142 36504 24148
rect 36360 23520 36412 23526
rect 36360 23462 36412 23468
rect 36372 23254 36400 23462
rect 36360 23248 36412 23254
rect 36360 23190 36412 23196
rect 36464 23186 36492 24142
rect 36452 23180 36504 23186
rect 36452 23122 36504 23128
rect 36636 23112 36688 23118
rect 36636 23054 36688 23060
rect 36820 23112 36872 23118
rect 36820 23054 36872 23060
rect 36544 22976 36596 22982
rect 36544 22918 36596 22924
rect 36360 22704 36412 22710
rect 36360 22646 36412 22652
rect 36268 21480 36320 21486
rect 36268 21422 36320 21428
rect 36176 20392 36228 20398
rect 36176 20334 36228 20340
rect 36268 19780 36320 19786
rect 36268 19722 36320 19728
rect 36280 19281 36308 19722
rect 36372 19310 36400 22646
rect 36452 21548 36504 21554
rect 36452 21490 36504 21496
rect 36464 20942 36492 21490
rect 36556 21486 36584 22918
rect 36648 22778 36676 23054
rect 36636 22772 36688 22778
rect 36636 22714 36688 22720
rect 36832 22098 36860 23054
rect 37004 22772 37056 22778
rect 37004 22714 37056 22720
rect 36820 22092 36872 22098
rect 36820 22034 36872 22040
rect 36544 21480 36596 21486
rect 36544 21422 36596 21428
rect 36912 21480 36964 21486
rect 36912 21422 36964 21428
rect 36452 20936 36504 20942
rect 36452 20878 36504 20884
rect 36464 20466 36492 20878
rect 36544 20868 36596 20874
rect 36544 20810 36596 20816
rect 36452 20460 36504 20466
rect 36452 20402 36504 20408
rect 36464 19378 36492 20402
rect 36556 19990 36584 20810
rect 36636 20800 36688 20806
rect 36636 20742 36688 20748
rect 36820 20800 36872 20806
rect 36820 20742 36872 20748
rect 36544 19984 36596 19990
rect 36544 19926 36596 19932
rect 36452 19372 36504 19378
rect 36452 19314 36504 19320
rect 36360 19304 36412 19310
rect 36266 19272 36322 19281
rect 36360 19246 36412 19252
rect 36266 19207 36322 19216
rect 36082 18864 36138 18873
rect 36082 18799 36138 18808
rect 36372 18737 36400 19246
rect 36556 19174 36584 19926
rect 36544 19168 36596 19174
rect 36544 19110 36596 19116
rect 36556 18834 36584 19110
rect 36648 18834 36676 20742
rect 36832 19990 36860 20742
rect 36924 20058 36952 21422
rect 37016 21010 37044 22714
rect 37004 21004 37056 21010
rect 37004 20946 37056 20952
rect 37004 20256 37056 20262
rect 37004 20198 37056 20204
rect 36912 20052 36964 20058
rect 36912 19994 36964 20000
rect 36820 19984 36872 19990
rect 36820 19926 36872 19932
rect 36728 19848 36780 19854
rect 36924 19802 36952 19994
rect 37016 19922 37044 20198
rect 37004 19916 37056 19922
rect 37004 19858 37056 19864
rect 36728 19790 36780 19796
rect 36740 19310 36768 19790
rect 36832 19774 36952 19802
rect 36728 19304 36780 19310
rect 36728 19246 36780 19252
rect 36728 19168 36780 19174
rect 36728 19110 36780 19116
rect 36544 18828 36596 18834
rect 36464 18788 36544 18816
rect 36358 18728 36414 18737
rect 36358 18663 36414 18672
rect 36174 18320 36230 18329
rect 36084 18284 36136 18290
rect 36174 18255 36176 18264
rect 36084 18226 36136 18232
rect 36228 18255 36230 18264
rect 36176 18226 36228 18232
rect 35992 16040 36044 16046
rect 35992 15982 36044 15988
rect 35900 15700 35952 15706
rect 35900 15642 35952 15648
rect 36096 14958 36124 18226
rect 36372 17610 36400 18663
rect 36464 18222 36492 18788
rect 36544 18770 36596 18776
rect 36636 18828 36688 18834
rect 36636 18770 36688 18776
rect 36544 18624 36596 18630
rect 36544 18566 36596 18572
rect 36636 18624 36688 18630
rect 36636 18566 36688 18572
rect 36452 18216 36504 18222
rect 36452 18158 36504 18164
rect 36360 17604 36412 17610
rect 36360 17546 36412 17552
rect 36268 17060 36320 17066
rect 36268 17002 36320 17008
rect 36176 16992 36228 16998
rect 36176 16934 36228 16940
rect 36188 16794 36216 16934
rect 36176 16788 36228 16794
rect 36176 16730 36228 16736
rect 36280 14958 36308 17002
rect 36360 16992 36412 16998
rect 36360 16934 36412 16940
rect 36084 14952 36136 14958
rect 36084 14894 36136 14900
rect 36268 14952 36320 14958
rect 36268 14894 36320 14900
rect 35808 14884 35860 14890
rect 35808 14826 35860 14832
rect 35820 14482 35848 14826
rect 35808 14476 35860 14482
rect 35808 14418 35860 14424
rect 35808 14340 35860 14346
rect 35808 14282 35860 14288
rect 35820 13938 35848 14282
rect 35808 13932 35860 13938
rect 35808 13874 35860 13880
rect 36084 13388 36136 13394
rect 36084 13330 36136 13336
rect 35808 13184 35860 13190
rect 35808 13126 35860 13132
rect 35716 11756 35768 11762
rect 35716 11698 35768 11704
rect 35728 10742 35756 11698
rect 35820 11354 35848 13126
rect 36096 12782 36124 13330
rect 36084 12776 36136 12782
rect 36084 12718 36136 12724
rect 36096 11354 36124 12718
rect 36176 12708 36228 12714
rect 36176 12650 36228 12656
rect 36188 11694 36216 12650
rect 36176 11688 36228 11694
rect 36176 11630 36228 11636
rect 35808 11348 35860 11354
rect 35808 11290 35860 11296
rect 36084 11348 36136 11354
rect 36084 11290 36136 11296
rect 35820 11014 35848 11290
rect 36176 11144 36228 11150
rect 36176 11086 36228 11092
rect 35808 11008 35860 11014
rect 35808 10950 35860 10956
rect 35716 10736 35768 10742
rect 35716 10678 35768 10684
rect 36188 10674 36216 11086
rect 36176 10668 36228 10674
rect 36176 10610 36228 10616
rect 35636 9608 35848 9636
rect 35346 9208 35402 9217
rect 35346 9143 35402 9152
rect 33138 9007 33140 9016
rect 33192 9007 33194 9016
rect 34336 9036 34388 9042
rect 33140 8978 33192 8984
rect 34336 8978 34388 8984
rect 34348 8362 34376 8978
rect 34520 8968 34572 8974
rect 34520 8910 34572 8916
rect 34336 8356 34388 8362
rect 34336 8298 34388 8304
rect 33876 8288 33928 8294
rect 33876 8230 33928 8236
rect 33888 7954 33916 8230
rect 34348 7954 34376 8298
rect 34532 8090 34560 8910
rect 34940 8732 35236 8752
rect 34996 8730 35020 8732
rect 35076 8730 35100 8732
rect 35156 8730 35180 8732
rect 35018 8678 35020 8730
rect 35082 8678 35094 8730
rect 35156 8678 35158 8730
rect 34996 8676 35020 8678
rect 35076 8676 35100 8678
rect 35156 8676 35180 8678
rect 34940 8656 35236 8676
rect 34520 8084 34572 8090
rect 34520 8026 34572 8032
rect 33876 7948 33928 7954
rect 33876 7890 33928 7896
rect 34336 7948 34388 7954
rect 34336 7890 34388 7896
rect 32956 7880 33008 7886
rect 32956 7822 33008 7828
rect 33140 7404 33192 7410
rect 33140 7346 33192 7352
rect 32588 6860 32640 6866
rect 32588 6802 32640 6808
rect 33152 6730 33180 7346
rect 34348 7342 34376 7890
rect 34796 7880 34848 7886
rect 34796 7822 34848 7828
rect 34520 7744 34572 7750
rect 34520 7686 34572 7692
rect 34336 7336 34388 7342
rect 34336 7278 34388 7284
rect 33232 6860 33284 6866
rect 33232 6802 33284 6808
rect 33140 6724 33192 6730
rect 33140 6666 33192 6672
rect 32312 6656 32364 6662
rect 32364 6616 32444 6644
rect 32312 6598 32364 6604
rect 32312 6452 32364 6458
rect 32312 6394 32364 6400
rect 32128 6248 32180 6254
rect 31850 6216 31906 6225
rect 32128 6190 32180 6196
rect 31850 6151 31906 6160
rect 31864 5778 31892 6151
rect 31852 5772 31904 5778
rect 31852 5714 31904 5720
rect 31760 5364 31812 5370
rect 31760 5306 31812 5312
rect 31864 5302 31892 5714
rect 32140 5710 32168 6190
rect 32324 6186 32352 6394
rect 32416 6254 32444 6616
rect 33244 6610 33272 6802
rect 33968 6792 34020 6798
rect 33968 6734 34020 6740
rect 34428 6792 34480 6798
rect 34428 6734 34480 6740
rect 33152 6582 33272 6610
rect 33152 6458 33180 6582
rect 33140 6452 33192 6458
rect 33140 6394 33192 6400
rect 32404 6248 32456 6254
rect 32404 6190 32456 6196
rect 32956 6248 33008 6254
rect 32956 6190 33008 6196
rect 32312 6180 32364 6186
rect 32312 6122 32364 6128
rect 32128 5704 32180 5710
rect 32128 5646 32180 5652
rect 32416 5642 32444 6190
rect 32968 5778 32996 6190
rect 32956 5772 33008 5778
rect 32956 5714 33008 5720
rect 32404 5636 32456 5642
rect 32404 5578 32456 5584
rect 32956 5636 33008 5642
rect 32956 5578 33008 5584
rect 31852 5296 31904 5302
rect 31852 5238 31904 5244
rect 32128 5160 32180 5166
rect 32128 5102 32180 5108
rect 32140 4758 32168 5102
rect 32680 5092 32732 5098
rect 32680 5034 32732 5040
rect 32128 4752 32180 4758
rect 32128 4694 32180 4700
rect 32692 4690 32720 5034
rect 32036 4684 32088 4690
rect 32036 4626 32088 4632
rect 32680 4684 32732 4690
rect 32680 4626 32732 4632
rect 31668 4616 31720 4622
rect 31668 4558 31720 4564
rect 30840 4480 30892 4486
rect 30840 4422 30892 4428
rect 30852 4146 30880 4422
rect 30380 4140 30432 4146
rect 30380 4082 30432 4088
rect 30564 4140 30616 4146
rect 30564 4082 30616 4088
rect 30840 4140 30892 4146
rect 30840 4082 30892 4088
rect 32048 3942 32076 4626
rect 32588 4072 32640 4078
rect 32588 4014 32640 4020
rect 31300 3936 31352 3942
rect 31300 3878 31352 3884
rect 32036 3936 32088 3942
rect 32036 3878 32088 3884
rect 31312 3738 31340 3878
rect 31208 3732 31260 3738
rect 31208 3674 31260 3680
rect 31300 3732 31352 3738
rect 31300 3674 31352 3680
rect 31024 3596 31076 3602
rect 31024 3538 31076 3544
rect 31036 3398 31064 3538
rect 31220 3534 31248 3674
rect 31208 3528 31260 3534
rect 31208 3470 31260 3476
rect 31668 3528 31720 3534
rect 31668 3470 31720 3476
rect 31024 3392 31076 3398
rect 31024 3334 31076 3340
rect 30196 3052 30248 3058
rect 30196 2994 30248 3000
rect 30012 2508 30064 2514
rect 30012 2450 30064 2456
rect 30208 2446 30236 2994
rect 30196 2440 30248 2446
rect 30196 2382 30248 2388
rect 31680 2378 31708 3470
rect 32600 3126 32628 4014
rect 32680 4004 32732 4010
rect 32680 3946 32732 3952
rect 32692 3670 32720 3946
rect 32680 3664 32732 3670
rect 32680 3606 32732 3612
rect 32968 3534 32996 5578
rect 32956 3528 33008 3534
rect 32956 3470 33008 3476
rect 32588 3120 32640 3126
rect 32588 3062 32640 3068
rect 31852 2984 31904 2990
rect 31852 2926 31904 2932
rect 31668 2372 31720 2378
rect 31668 2314 31720 2320
rect 31300 2304 31352 2310
rect 31300 2246 31352 2252
rect 29736 1148 29788 1154
rect 29736 1090 29788 1096
rect 31312 800 31340 2246
rect 31864 2106 31892 2926
rect 33152 2446 33180 6394
rect 33980 6254 34008 6734
rect 34440 6322 34468 6734
rect 34428 6316 34480 6322
rect 34428 6258 34480 6264
rect 33968 6248 34020 6254
rect 33968 6190 34020 6196
rect 33968 6112 34020 6118
rect 33968 6054 34020 6060
rect 33980 5234 34008 6054
rect 33968 5228 34020 5234
rect 33968 5170 34020 5176
rect 34532 5166 34560 7686
rect 34704 7268 34756 7274
rect 34704 7210 34756 7216
rect 34612 6860 34664 6866
rect 34612 6802 34664 6808
rect 34624 5302 34652 6802
rect 34612 5296 34664 5302
rect 34612 5238 34664 5244
rect 34520 5160 34572 5166
rect 34520 5102 34572 5108
rect 33416 4752 33468 4758
rect 33416 4694 33468 4700
rect 33428 4078 33456 4694
rect 34336 4684 34388 4690
rect 34336 4626 34388 4632
rect 33600 4140 33652 4146
rect 33600 4082 33652 4088
rect 33232 4072 33284 4078
rect 33232 4014 33284 4020
rect 33416 4072 33468 4078
rect 33416 4014 33468 4020
rect 33244 2582 33272 4014
rect 33428 3398 33456 4014
rect 33612 3602 33640 4082
rect 33692 4072 33744 4078
rect 33692 4014 33744 4020
rect 33876 4072 33928 4078
rect 33876 4014 33928 4020
rect 33704 3942 33732 4014
rect 33692 3936 33744 3942
rect 33690 3904 33692 3913
rect 33744 3904 33746 3913
rect 33690 3839 33746 3848
rect 33704 3813 33732 3839
rect 33600 3596 33652 3602
rect 33600 3538 33652 3544
rect 33416 3392 33468 3398
rect 33416 3334 33468 3340
rect 33600 3392 33652 3398
rect 33600 3334 33652 3340
rect 33612 2990 33640 3334
rect 33888 2990 33916 4014
rect 34348 4010 34376 4626
rect 34520 4616 34572 4622
rect 34520 4558 34572 4564
rect 34428 4072 34480 4078
rect 34428 4014 34480 4020
rect 34336 4004 34388 4010
rect 34336 3946 34388 3952
rect 34348 3738 34376 3946
rect 34336 3732 34388 3738
rect 34336 3674 34388 3680
rect 34440 2990 34468 4014
rect 34532 3058 34560 4558
rect 34624 4146 34652 5238
rect 34716 5234 34744 7210
rect 34808 5370 34836 7822
rect 34940 7644 35236 7664
rect 34996 7642 35020 7644
rect 35076 7642 35100 7644
rect 35156 7642 35180 7644
rect 35018 7590 35020 7642
rect 35082 7590 35094 7642
rect 35156 7590 35158 7642
rect 34996 7588 35020 7590
rect 35076 7588 35100 7590
rect 35156 7588 35180 7590
rect 34940 7568 35236 7588
rect 34940 6556 35236 6576
rect 34996 6554 35020 6556
rect 35076 6554 35100 6556
rect 35156 6554 35180 6556
rect 35018 6502 35020 6554
rect 35082 6502 35094 6554
rect 35156 6502 35158 6554
rect 34996 6500 35020 6502
rect 35076 6500 35100 6502
rect 35156 6500 35180 6502
rect 34940 6480 35236 6500
rect 34940 5468 35236 5488
rect 34996 5466 35020 5468
rect 35076 5466 35100 5468
rect 35156 5466 35180 5468
rect 35018 5414 35020 5466
rect 35082 5414 35094 5466
rect 35156 5414 35158 5466
rect 34996 5412 35020 5414
rect 35076 5412 35100 5414
rect 35156 5412 35180 5414
rect 34940 5392 35236 5412
rect 34796 5364 34848 5370
rect 34796 5306 34848 5312
rect 34704 5228 34756 5234
rect 34704 5170 34756 5176
rect 34704 4616 34756 4622
rect 34704 4558 34756 4564
rect 34612 4140 34664 4146
rect 34612 4082 34664 4088
rect 34716 3534 34744 4558
rect 35360 4457 35388 9143
rect 35820 8974 35848 9608
rect 36176 9512 36228 9518
rect 36176 9454 36228 9460
rect 35808 8968 35860 8974
rect 35808 8910 35860 8916
rect 35820 7546 35848 8910
rect 36188 8634 36216 9454
rect 36176 8628 36228 8634
rect 36176 8570 36228 8576
rect 35900 8424 35952 8430
rect 35900 8366 35952 8372
rect 35912 7954 35940 8366
rect 35992 8356 36044 8362
rect 35992 8298 36044 8304
rect 35900 7948 35952 7954
rect 35900 7890 35952 7896
rect 35912 7546 35940 7890
rect 36004 7818 36032 8298
rect 35992 7812 36044 7818
rect 35992 7754 36044 7760
rect 35808 7540 35860 7546
rect 35808 7482 35860 7488
rect 35900 7540 35952 7546
rect 35900 7482 35952 7488
rect 36268 6860 36320 6866
rect 36268 6802 36320 6808
rect 35440 6792 35492 6798
rect 35440 6734 35492 6740
rect 35900 6792 35952 6798
rect 35900 6734 35952 6740
rect 36176 6792 36228 6798
rect 36176 6734 36228 6740
rect 35452 5642 35480 6734
rect 35912 5778 35940 6734
rect 35992 6452 36044 6458
rect 35992 6394 36044 6400
rect 35900 5772 35952 5778
rect 35900 5714 35952 5720
rect 36004 5710 36032 6394
rect 36084 6316 36136 6322
rect 36084 6258 36136 6264
rect 35992 5704 36044 5710
rect 35992 5646 36044 5652
rect 35440 5636 35492 5642
rect 35440 5578 35492 5584
rect 36004 5234 36032 5646
rect 35992 5228 36044 5234
rect 35992 5170 36044 5176
rect 36096 4690 36124 6258
rect 36188 5846 36216 6734
rect 36176 5840 36228 5846
rect 36176 5782 36228 5788
rect 36084 4684 36136 4690
rect 36084 4626 36136 4632
rect 36280 4622 36308 6802
rect 36372 5234 36400 16934
rect 36556 14482 36584 18566
rect 36648 17746 36676 18566
rect 36740 17746 36768 19110
rect 36636 17740 36688 17746
rect 36636 17682 36688 17688
rect 36728 17740 36780 17746
rect 36728 17682 36780 17688
rect 36832 16658 36860 19774
rect 36912 19304 36964 19310
rect 36912 19246 36964 19252
rect 36924 18426 36952 19246
rect 36912 18420 36964 18426
rect 36912 18362 36964 18368
rect 36636 16652 36688 16658
rect 36636 16594 36688 16600
rect 36820 16652 36872 16658
rect 36820 16594 36872 16600
rect 36648 15706 36676 16594
rect 36636 15700 36688 15706
rect 36636 15642 36688 15648
rect 36544 14476 36596 14482
rect 36544 14418 36596 14424
rect 36544 13728 36596 13734
rect 36544 13670 36596 13676
rect 36556 13394 36584 13670
rect 36544 13388 36596 13394
rect 36544 13330 36596 13336
rect 36728 13388 36780 13394
rect 36728 13330 36780 13336
rect 36556 12782 36584 13330
rect 36544 12776 36596 12782
rect 36544 12718 36596 12724
rect 36556 12306 36584 12718
rect 36544 12300 36596 12306
rect 36544 12242 36596 12248
rect 36740 11830 36768 13330
rect 36728 11824 36780 11830
rect 36728 11766 36780 11772
rect 36544 10668 36596 10674
rect 36544 10610 36596 10616
rect 36452 10600 36504 10606
rect 36452 10542 36504 10548
rect 36464 8838 36492 10542
rect 36452 8832 36504 8838
rect 36452 8774 36504 8780
rect 36556 8430 36584 10610
rect 37004 10056 37056 10062
rect 37004 9998 37056 10004
rect 37016 9586 37044 9998
rect 37004 9580 37056 9586
rect 37004 9522 37056 9528
rect 37108 9042 37136 25094
rect 37292 24750 37320 25842
rect 37280 24744 37332 24750
rect 37280 24686 37332 24692
rect 37292 23730 37320 24686
rect 37384 24018 37412 30126
rect 37740 29708 37792 29714
rect 37740 29650 37792 29656
rect 37556 29232 37608 29238
rect 37556 29174 37608 29180
rect 37568 28082 37596 29174
rect 37752 28218 37780 29650
rect 37844 29102 37872 30670
rect 37924 29708 37976 29714
rect 37924 29650 37976 29656
rect 37832 29096 37884 29102
rect 37832 29038 37884 29044
rect 37740 28212 37792 28218
rect 37740 28154 37792 28160
rect 37556 28076 37608 28082
rect 37556 28018 37608 28024
rect 37752 26926 37780 28154
rect 37844 26994 37872 29038
rect 37832 26988 37884 26994
rect 37832 26930 37884 26936
rect 37740 26920 37792 26926
rect 37740 26862 37792 26868
rect 37936 26586 37964 29650
rect 38120 28626 38148 31078
rect 38108 28620 38160 28626
rect 38108 28562 38160 28568
rect 38016 27872 38068 27878
rect 38016 27814 38068 27820
rect 38028 27538 38056 27814
rect 38016 27532 38068 27538
rect 38016 27474 38068 27480
rect 37924 26580 37976 26586
rect 37924 26522 37976 26528
rect 37740 26444 37792 26450
rect 37740 26386 37792 26392
rect 37556 25832 37608 25838
rect 37556 25774 37608 25780
rect 37568 24818 37596 25774
rect 37752 25294 37780 26386
rect 37924 25696 37976 25702
rect 37924 25638 37976 25644
rect 37740 25288 37792 25294
rect 37740 25230 37792 25236
rect 37556 24812 37608 24818
rect 37556 24754 37608 24760
rect 37464 24744 37516 24750
rect 37464 24686 37516 24692
rect 37476 24138 37504 24686
rect 37464 24132 37516 24138
rect 37464 24074 37516 24080
rect 37384 23990 37504 24018
rect 37280 23724 37332 23730
rect 37280 23666 37332 23672
rect 37280 22636 37332 22642
rect 37280 22578 37332 22584
rect 37188 22500 37240 22506
rect 37188 22442 37240 22448
rect 37200 19922 37228 22442
rect 37292 20942 37320 22578
rect 37372 22432 37424 22438
rect 37372 22374 37424 22380
rect 37384 22098 37412 22374
rect 37372 22092 37424 22098
rect 37372 22034 37424 22040
rect 37280 20936 37332 20942
rect 37280 20878 37332 20884
rect 37188 19916 37240 19922
rect 37188 19858 37240 19864
rect 37384 18970 37412 22034
rect 37372 18964 37424 18970
rect 37372 18906 37424 18912
rect 37188 18692 37240 18698
rect 37188 18634 37240 18640
rect 37200 18222 37228 18634
rect 37372 18420 37424 18426
rect 37372 18362 37424 18368
rect 37188 18216 37240 18222
rect 37188 18158 37240 18164
rect 37384 17116 37412 18362
rect 37476 17542 37504 23990
rect 37740 23656 37792 23662
rect 37740 23598 37792 23604
rect 37752 23050 37780 23598
rect 37740 23044 37792 23050
rect 37740 22986 37792 22992
rect 37936 22642 37964 25638
rect 38108 24200 38160 24206
rect 38108 24142 38160 24148
rect 38016 23180 38068 23186
rect 38016 23122 38068 23128
rect 37924 22636 37976 22642
rect 37924 22578 37976 22584
rect 37832 22228 37884 22234
rect 37832 22170 37884 22176
rect 37844 21554 37872 22170
rect 37922 21584 37978 21593
rect 37832 21548 37884 21554
rect 37922 21519 37978 21528
rect 37832 21490 37884 21496
rect 37740 20392 37792 20398
rect 37740 20334 37792 20340
rect 37752 19990 37780 20334
rect 37740 19984 37792 19990
rect 37740 19926 37792 19932
rect 37740 18964 37792 18970
rect 37740 18906 37792 18912
rect 37648 18216 37700 18222
rect 37648 18158 37700 18164
rect 37660 17882 37688 18158
rect 37648 17876 37700 17882
rect 37648 17818 37700 17824
rect 37464 17536 37516 17542
rect 37464 17478 37516 17484
rect 37464 17128 37516 17134
rect 37384 17088 37464 17116
rect 37384 16046 37412 17088
rect 37464 17070 37516 17076
rect 37556 16584 37608 16590
rect 37556 16526 37608 16532
rect 37568 16114 37596 16526
rect 37556 16108 37608 16114
rect 37556 16050 37608 16056
rect 37372 16040 37424 16046
rect 37372 15982 37424 15988
rect 37384 15502 37412 15982
rect 37752 15586 37780 18906
rect 37660 15558 37780 15586
rect 37936 15570 37964 21519
rect 38028 17882 38056 23122
rect 38120 22574 38148 24142
rect 38108 22568 38160 22574
rect 38108 22510 38160 22516
rect 38120 22098 38148 22510
rect 38108 22092 38160 22098
rect 38108 22034 38160 22040
rect 38108 20596 38160 20602
rect 38108 20538 38160 20544
rect 38016 17876 38068 17882
rect 38016 17818 38068 17824
rect 38028 16794 38056 17818
rect 38016 16788 38068 16794
rect 38016 16730 38068 16736
rect 37924 15564 37976 15570
rect 37372 15496 37424 15502
rect 37372 15438 37424 15444
rect 37384 15026 37412 15438
rect 37372 15020 37424 15026
rect 37372 14962 37424 14968
rect 37188 12776 37240 12782
rect 37188 12718 37240 12724
rect 37200 11762 37228 12718
rect 37188 11756 37240 11762
rect 37188 11698 37240 11704
rect 37200 10674 37228 11698
rect 37188 10668 37240 10674
rect 37188 10610 37240 10616
rect 37186 10160 37242 10169
rect 37186 10095 37188 10104
rect 37240 10095 37242 10104
rect 37188 10066 37240 10072
rect 37464 9988 37516 9994
rect 37464 9930 37516 9936
rect 37476 9518 37504 9930
rect 37464 9512 37516 9518
rect 37464 9454 37516 9460
rect 37280 9376 37332 9382
rect 37280 9318 37332 9324
rect 37292 9178 37320 9318
rect 37280 9172 37332 9178
rect 37280 9114 37332 9120
rect 37096 9036 37148 9042
rect 37096 8978 37148 8984
rect 36820 8968 36872 8974
rect 36820 8910 36872 8916
rect 36832 8498 36860 8910
rect 36820 8492 36872 8498
rect 36820 8434 36872 8440
rect 36544 8424 36596 8430
rect 36544 8366 36596 8372
rect 36636 8424 36688 8430
rect 36636 8366 36688 8372
rect 36648 7954 36676 8366
rect 37108 8022 37136 8978
rect 37096 8016 37148 8022
rect 37096 7958 37148 7964
rect 37660 7954 37688 15558
rect 37924 15506 37976 15512
rect 37924 15360 37976 15366
rect 37924 15302 37976 15308
rect 37740 14952 37792 14958
rect 37740 14894 37792 14900
rect 37752 14618 37780 14894
rect 37740 14612 37792 14618
rect 37740 14554 37792 14560
rect 37740 14476 37792 14482
rect 37740 14418 37792 14424
rect 37832 14476 37884 14482
rect 37832 14418 37884 14424
rect 37752 14074 37780 14418
rect 37740 14068 37792 14074
rect 37740 14010 37792 14016
rect 37752 13394 37780 14010
rect 37844 13462 37872 14418
rect 37832 13456 37884 13462
rect 37832 13398 37884 13404
rect 37740 13388 37792 13394
rect 37740 13330 37792 13336
rect 37740 13252 37792 13258
rect 37740 13194 37792 13200
rect 37752 12850 37780 13194
rect 37740 12844 37792 12850
rect 37740 12786 37792 12792
rect 37936 11762 37964 15302
rect 38120 15162 38148 20538
rect 38212 19009 38240 34462
rect 38292 34060 38344 34066
rect 38292 34002 38344 34008
rect 38304 33522 38332 34002
rect 38476 33584 38528 33590
rect 38476 33526 38528 33532
rect 38292 33516 38344 33522
rect 38292 33458 38344 33464
rect 38488 31958 38516 33526
rect 39026 33008 39082 33017
rect 38568 32972 38620 32978
rect 39026 32943 39082 32952
rect 38568 32914 38620 32920
rect 38476 31952 38528 31958
rect 38476 31894 38528 31900
rect 38292 31884 38344 31890
rect 38292 31826 38344 31832
rect 38304 28626 38332 31826
rect 38476 31816 38528 31822
rect 38476 31758 38528 31764
rect 38488 30802 38516 31758
rect 38580 31142 38608 32914
rect 38752 32904 38804 32910
rect 38752 32846 38804 32852
rect 38764 31890 38792 32846
rect 39040 32570 39068 32943
rect 39028 32564 39080 32570
rect 39028 32506 39080 32512
rect 38752 31884 38804 31890
rect 38752 31826 38804 31832
rect 38568 31136 38620 31142
rect 38568 31078 38620 31084
rect 38476 30796 38528 30802
rect 38476 30738 38528 30744
rect 39118 30288 39174 30297
rect 39118 30223 39120 30232
rect 39172 30223 39174 30232
rect 39120 30194 39172 30200
rect 38568 30048 38620 30054
rect 38568 29990 38620 29996
rect 38580 29714 38608 29990
rect 38568 29708 38620 29714
rect 38568 29650 38620 29656
rect 38476 29096 38528 29102
rect 38476 29038 38528 29044
rect 38292 28620 38344 28626
rect 38292 28562 38344 28568
rect 38384 28620 38436 28626
rect 38384 28562 38436 28568
rect 38304 27538 38332 28562
rect 38396 27606 38424 28562
rect 38384 27600 38436 27606
rect 38384 27542 38436 27548
rect 38292 27532 38344 27538
rect 38292 27474 38344 27480
rect 38304 26382 38332 27474
rect 38488 27418 38516 29038
rect 38660 29028 38712 29034
rect 38660 28970 38712 28976
rect 38672 28490 38700 28970
rect 38660 28484 38712 28490
rect 38660 28426 38712 28432
rect 38568 27532 38620 27538
rect 38568 27474 38620 27480
rect 38396 27390 38516 27418
rect 38396 26450 38424 27390
rect 38580 26994 38608 27474
rect 38844 27328 38896 27334
rect 38844 27270 38896 27276
rect 39946 27296 40002 27305
rect 38568 26988 38620 26994
rect 38568 26930 38620 26936
rect 38476 26580 38528 26586
rect 38476 26522 38528 26528
rect 38384 26444 38436 26450
rect 38384 26386 38436 26392
rect 38292 26376 38344 26382
rect 38292 26318 38344 26324
rect 38488 25362 38516 26522
rect 38660 26512 38712 26518
rect 38660 26454 38712 26460
rect 38672 26042 38700 26454
rect 38752 26444 38804 26450
rect 38752 26386 38804 26392
rect 38660 26036 38712 26042
rect 38660 25978 38712 25984
rect 38764 25362 38792 26386
rect 38476 25356 38528 25362
rect 38476 25298 38528 25304
rect 38752 25356 38804 25362
rect 38752 25298 38804 25304
rect 38856 25294 38884 27270
rect 39946 27231 39948 27240
rect 40000 27231 40002 27240
rect 39948 27202 40000 27208
rect 39120 25356 39172 25362
rect 39120 25298 39172 25304
rect 38384 25288 38436 25294
rect 38384 25230 38436 25236
rect 38844 25288 38896 25294
rect 38844 25230 38896 25236
rect 38292 25220 38344 25226
rect 38292 25162 38344 25168
rect 38304 24585 38332 25162
rect 38290 24576 38346 24585
rect 38290 24511 38346 24520
rect 38292 24268 38344 24274
rect 38292 24210 38344 24216
rect 38304 23186 38332 24210
rect 38292 23180 38344 23186
rect 38292 23122 38344 23128
rect 38292 22636 38344 22642
rect 38292 22578 38344 22584
rect 38304 20482 38332 22578
rect 38396 20618 38424 25230
rect 38568 24608 38620 24614
rect 38568 24550 38620 24556
rect 38580 22574 38608 24550
rect 38936 24268 38988 24274
rect 38936 24210 38988 24216
rect 38948 23866 38976 24210
rect 38936 23860 38988 23866
rect 38936 23802 38988 23808
rect 39028 22976 39080 22982
rect 39028 22918 39080 22924
rect 38568 22568 38620 22574
rect 38488 22528 38568 22556
rect 38488 22030 38516 22528
rect 38568 22510 38620 22516
rect 38476 22024 38528 22030
rect 38476 21966 38528 21972
rect 39040 21418 39068 22918
rect 39028 21412 39080 21418
rect 39028 21354 39080 21360
rect 38660 21344 38712 21350
rect 38660 21286 38712 21292
rect 38672 21010 38700 21286
rect 38660 21004 38712 21010
rect 38660 20946 38712 20952
rect 38396 20590 38516 20618
rect 38304 20454 38424 20482
rect 38292 20392 38344 20398
rect 38292 20334 38344 20340
rect 38304 19854 38332 20334
rect 38292 19848 38344 19854
rect 38292 19790 38344 19796
rect 38198 19000 38254 19009
rect 38198 18935 38254 18944
rect 38304 18834 38332 19790
rect 38292 18828 38344 18834
rect 38292 18770 38344 18776
rect 38292 18080 38344 18086
rect 38292 18022 38344 18028
rect 38304 17218 38332 18022
rect 38212 17202 38332 17218
rect 38200 17196 38332 17202
rect 38252 17190 38332 17196
rect 38200 17138 38252 17144
rect 38304 16726 38332 17190
rect 38292 16720 38344 16726
rect 38292 16662 38344 16668
rect 38396 16590 38424 20454
rect 38488 17270 38516 20590
rect 38752 20256 38804 20262
rect 38752 20198 38804 20204
rect 38764 19922 38792 20198
rect 38752 19916 38804 19922
rect 38752 19858 38804 19864
rect 38660 17740 38712 17746
rect 38660 17682 38712 17688
rect 38476 17264 38528 17270
rect 38476 17206 38528 17212
rect 38384 16584 38436 16590
rect 38384 16526 38436 16532
rect 38396 15502 38424 16526
rect 38488 15994 38516 17206
rect 38568 17128 38620 17134
rect 38568 17070 38620 17076
rect 38580 16726 38608 17070
rect 38672 16998 38700 17682
rect 38660 16992 38712 16998
rect 38660 16934 38712 16940
rect 38568 16720 38620 16726
rect 38568 16662 38620 16668
rect 38672 16658 38700 16934
rect 38660 16652 38712 16658
rect 38660 16594 38712 16600
rect 38488 15966 38608 15994
rect 38474 15872 38530 15881
rect 38474 15807 38530 15816
rect 38488 15570 38516 15807
rect 38476 15564 38528 15570
rect 38476 15506 38528 15512
rect 38384 15496 38436 15502
rect 38384 15438 38436 15444
rect 38580 15348 38608 15966
rect 38396 15320 38608 15348
rect 38108 15156 38160 15162
rect 38108 15098 38160 15104
rect 38120 13870 38148 15098
rect 38108 13864 38160 13870
rect 38108 13806 38160 13812
rect 38200 13388 38252 13394
rect 38200 13330 38252 13336
rect 38212 12986 38240 13330
rect 38200 12980 38252 12986
rect 38200 12922 38252 12928
rect 37924 11756 37976 11762
rect 37924 11698 37976 11704
rect 37832 11552 37884 11558
rect 37832 11494 37884 11500
rect 37844 11218 37872 11494
rect 37832 11212 37884 11218
rect 37832 11154 37884 11160
rect 37924 11212 37976 11218
rect 37924 11154 37976 11160
rect 37936 10810 37964 11154
rect 37924 10804 37976 10810
rect 37924 10746 37976 10752
rect 38396 10130 38424 15320
rect 38476 14816 38528 14822
rect 38476 14758 38528 14764
rect 38488 13870 38516 14758
rect 38568 14408 38620 14414
rect 38568 14350 38620 14356
rect 38580 13938 38608 14350
rect 38568 13932 38620 13938
rect 38568 13874 38620 13880
rect 38476 13864 38528 13870
rect 38476 13806 38528 13812
rect 38488 12238 38516 13806
rect 38568 13320 38620 13326
rect 38568 13262 38620 13268
rect 38580 12306 38608 13262
rect 38568 12300 38620 12306
rect 38568 12242 38620 12248
rect 38476 12232 38528 12238
rect 38476 12174 38528 12180
rect 38672 11354 38700 16594
rect 38660 11348 38712 11354
rect 38660 11290 38712 11296
rect 37924 10124 37976 10130
rect 37924 10066 37976 10072
rect 38108 10124 38160 10130
rect 38108 10066 38160 10072
rect 38384 10124 38436 10130
rect 38384 10066 38436 10072
rect 37740 9512 37792 9518
rect 37740 9454 37792 9460
rect 37752 9382 37780 9454
rect 37740 9376 37792 9382
rect 37740 9318 37792 9324
rect 37936 9110 37964 10066
rect 38120 9586 38148 10066
rect 38292 9920 38344 9926
rect 38292 9862 38344 9868
rect 38108 9580 38160 9586
rect 38108 9522 38160 9528
rect 37924 9104 37976 9110
rect 37924 9046 37976 9052
rect 37936 8634 37964 9046
rect 37924 8628 37976 8634
rect 37924 8570 37976 8576
rect 37936 7954 37964 8570
rect 38120 8430 38148 9522
rect 38304 9042 38332 9862
rect 38764 9654 38792 19858
rect 38936 19780 38988 19786
rect 38936 19722 38988 19728
rect 38948 18834 38976 19722
rect 38936 18828 38988 18834
rect 38936 18770 38988 18776
rect 38936 17740 38988 17746
rect 38936 17682 38988 17688
rect 38948 17338 38976 17682
rect 38936 17332 38988 17338
rect 38936 17274 38988 17280
rect 38948 16250 38976 17274
rect 38936 16244 38988 16250
rect 38936 16186 38988 16192
rect 38934 13152 38990 13161
rect 38934 13087 38990 13096
rect 38752 9648 38804 9654
rect 38752 9590 38804 9596
rect 38568 9376 38620 9382
rect 38568 9318 38620 9324
rect 38292 9036 38344 9042
rect 38292 8978 38344 8984
rect 38108 8424 38160 8430
rect 38108 8366 38160 8372
rect 38292 8016 38344 8022
rect 38292 7958 38344 7964
rect 36636 7948 36688 7954
rect 36636 7890 36688 7896
rect 37648 7948 37700 7954
rect 37648 7890 37700 7896
rect 37740 7948 37792 7954
rect 37740 7890 37792 7896
rect 37924 7948 37976 7954
rect 37924 7890 37976 7896
rect 36728 7744 36780 7750
rect 36728 7686 36780 7692
rect 36740 6866 36768 7686
rect 36728 6860 36780 6866
rect 36728 6802 36780 6808
rect 37372 6248 37424 6254
rect 37372 6190 37424 6196
rect 37384 5914 37412 6190
rect 37372 5908 37424 5914
rect 37372 5850 37424 5856
rect 37004 5772 37056 5778
rect 37004 5714 37056 5720
rect 37016 5370 37044 5714
rect 37004 5364 37056 5370
rect 37004 5306 37056 5312
rect 36360 5228 36412 5234
rect 36360 5170 36412 5176
rect 37660 5166 37688 7890
rect 37752 7342 37780 7890
rect 37832 7404 37884 7410
rect 37832 7346 37884 7352
rect 37740 7336 37792 7342
rect 37740 7278 37792 7284
rect 37740 6724 37792 6730
rect 37740 6666 37792 6672
rect 37752 6322 37780 6666
rect 37740 6316 37792 6322
rect 37740 6258 37792 6264
rect 37844 5778 37872 7346
rect 38304 7342 38332 7958
rect 38476 7812 38528 7818
rect 38476 7754 38528 7760
rect 38292 7336 38344 7342
rect 38292 7278 38344 7284
rect 38488 6866 38516 7754
rect 38580 7449 38608 9318
rect 38566 7440 38622 7449
rect 38566 7375 38622 7384
rect 38844 7336 38896 7342
rect 38844 7278 38896 7284
rect 38016 6860 38068 6866
rect 38016 6802 38068 6808
rect 38384 6860 38436 6866
rect 38384 6802 38436 6808
rect 38476 6860 38528 6866
rect 38476 6802 38528 6808
rect 37832 5772 37884 5778
rect 37832 5714 37884 5720
rect 37844 5234 37872 5714
rect 38028 5370 38056 6802
rect 38396 5914 38424 6802
rect 38856 6458 38884 7278
rect 38844 6452 38896 6458
rect 38844 6394 38896 6400
rect 38384 5908 38436 5914
rect 38384 5850 38436 5856
rect 38856 5778 38884 6394
rect 38200 5772 38252 5778
rect 38200 5714 38252 5720
rect 38844 5772 38896 5778
rect 38844 5714 38896 5720
rect 38016 5364 38068 5370
rect 38016 5306 38068 5312
rect 37832 5228 37884 5234
rect 37832 5170 37884 5176
rect 37648 5160 37700 5166
rect 37648 5102 37700 5108
rect 37660 4690 37688 5102
rect 38212 4826 38240 5714
rect 38200 4820 38252 4826
rect 38200 4762 38252 4768
rect 37648 4684 37700 4690
rect 37648 4626 37700 4632
rect 35624 4616 35676 4622
rect 35624 4558 35676 4564
rect 35992 4616 36044 4622
rect 35992 4558 36044 4564
rect 36268 4616 36320 4622
rect 36268 4558 36320 4564
rect 35346 4448 35402 4457
rect 34940 4380 35236 4400
rect 35346 4383 35402 4392
rect 34996 4378 35020 4380
rect 35076 4378 35100 4380
rect 35156 4378 35180 4380
rect 35018 4326 35020 4378
rect 35082 4326 35094 4378
rect 35156 4326 35158 4378
rect 34996 4324 35020 4326
rect 35076 4324 35100 4326
rect 35156 4324 35180 4326
rect 34940 4304 35236 4324
rect 35636 4146 35664 4558
rect 36004 4282 36032 4558
rect 35992 4276 36044 4282
rect 35992 4218 36044 4224
rect 38948 4146 38976 13087
rect 39132 12850 39160 25298
rect 39120 12844 39172 12850
rect 39120 12786 39172 12792
rect 39132 12374 39160 12786
rect 39120 12368 39172 12374
rect 39120 12310 39172 12316
rect 35624 4140 35676 4146
rect 35624 4082 35676 4088
rect 38936 4140 38988 4146
rect 38936 4082 38988 4088
rect 37740 4072 37792 4078
rect 37740 4014 37792 4020
rect 35440 3936 35492 3942
rect 35440 3878 35492 3884
rect 35898 3904 35954 3913
rect 34704 3528 34756 3534
rect 34704 3470 34756 3476
rect 35452 3398 35480 3878
rect 35898 3839 35954 3848
rect 35440 3392 35492 3398
rect 35440 3334 35492 3340
rect 34940 3292 35236 3312
rect 34996 3290 35020 3292
rect 35076 3290 35100 3292
rect 35156 3290 35180 3292
rect 35018 3238 35020 3290
rect 35082 3238 35094 3290
rect 35156 3238 35158 3290
rect 34996 3236 35020 3238
rect 35076 3236 35100 3238
rect 35156 3236 35180 3238
rect 34940 3216 35236 3236
rect 35452 3126 35480 3334
rect 35440 3120 35492 3126
rect 35440 3062 35492 3068
rect 34520 3052 34572 3058
rect 34520 2994 34572 3000
rect 33600 2984 33652 2990
rect 33600 2926 33652 2932
rect 33876 2984 33928 2990
rect 33876 2926 33928 2932
rect 34428 2984 34480 2990
rect 34428 2926 34480 2932
rect 33324 2916 33376 2922
rect 33324 2858 33376 2864
rect 33232 2576 33284 2582
rect 33232 2518 33284 2524
rect 33140 2440 33192 2446
rect 33140 2382 33192 2388
rect 33152 2310 33180 2382
rect 33140 2304 33192 2310
rect 33140 2246 33192 2252
rect 31852 2100 31904 2106
rect 31852 2042 31904 2048
rect 33336 800 33364 2858
rect 33508 2848 33560 2854
rect 33508 2790 33560 2796
rect 33520 2514 33548 2790
rect 33508 2508 33560 2514
rect 33508 2450 33560 2456
rect 34440 2310 34468 2926
rect 35452 2514 35480 3062
rect 35912 2990 35940 3839
rect 37096 3392 37148 3398
rect 37096 3334 37148 3340
rect 35900 2984 35952 2990
rect 35900 2926 35952 2932
rect 35440 2508 35492 2514
rect 35440 2450 35492 2456
rect 34428 2304 34480 2310
rect 34428 2246 34480 2252
rect 34940 2204 35236 2224
rect 34996 2202 35020 2204
rect 35076 2202 35100 2204
rect 35156 2202 35180 2204
rect 35018 2150 35020 2202
rect 35082 2150 35094 2202
rect 35156 2150 35158 2202
rect 34996 2148 35020 2150
rect 35076 2148 35100 2150
rect 35156 2148 35180 2150
rect 34940 2128 35236 2148
rect 37108 1737 37136 3334
rect 37752 3194 37780 4014
rect 37740 3188 37792 3194
rect 37740 3130 37792 3136
rect 39028 2916 39080 2922
rect 39028 2858 39080 2864
rect 37188 2304 37240 2310
rect 37188 2246 37240 2252
rect 37094 1728 37150 1737
rect 37094 1663 37150 1672
rect 35164 1148 35216 1154
rect 35164 1090 35216 1096
rect 35176 800 35204 1090
rect 37200 800 37228 2246
rect 39040 800 39068 2858
rect 570 0 626 800
rect 2410 0 2466 800
rect 4250 0 4306 800
rect 6274 0 6330 800
rect 8114 0 8170 800
rect 10138 0 10194 800
rect 11978 0 12034 800
rect 14002 0 14058 800
rect 15842 0 15898 800
rect 17866 0 17922 800
rect 19706 0 19762 800
rect 21730 0 21786 800
rect 23570 0 23626 800
rect 25594 0 25650 800
rect 27434 0 27490 800
rect 29458 0 29514 800
rect 31298 0 31354 800
rect 33322 0 33378 800
rect 35162 0 35218 800
rect 37186 0 37242 800
rect 39026 0 39082 800
<< via2 >>
rect 4220 38106 4276 38108
rect 4300 38106 4356 38108
rect 4380 38106 4436 38108
rect 4460 38106 4516 38108
rect 4220 38054 4246 38106
rect 4246 38054 4276 38106
rect 4300 38054 4310 38106
rect 4310 38054 4356 38106
rect 4380 38054 4426 38106
rect 4426 38054 4436 38106
rect 4460 38054 4490 38106
rect 4490 38054 4516 38106
rect 4220 38052 4276 38054
rect 4300 38052 4356 38054
rect 4380 38052 4436 38054
rect 4460 38052 4516 38054
rect 2778 37848 2834 37904
rect 18 30776 74 30832
rect 2962 32136 3018 32192
rect 2318 25780 2320 25800
rect 2320 25780 2372 25800
rect 2372 25780 2374 25800
rect 2318 25744 2374 25780
rect 2870 26424 2926 26480
rect 2778 23432 2834 23488
rect 1950 18672 2006 18728
rect 1950 17720 2006 17776
rect 3514 28736 3570 28792
rect 3422 20712 3478 20768
rect 1674 14476 1730 14512
rect 1674 14456 1676 14476
rect 1676 14456 1728 14476
rect 1728 14456 1730 14476
rect 3054 12008 3110 12064
rect 1582 7268 1638 7304
rect 1582 7248 1584 7268
rect 1584 7248 1636 7268
rect 1636 7248 1638 7268
rect 4220 37018 4276 37020
rect 4300 37018 4356 37020
rect 4380 37018 4436 37020
rect 4460 37018 4516 37020
rect 4220 36966 4246 37018
rect 4246 36966 4276 37018
rect 4300 36966 4310 37018
rect 4310 36966 4356 37018
rect 4380 36966 4426 37018
rect 4426 36966 4436 37018
rect 4460 36966 4490 37018
rect 4490 36966 4516 37018
rect 4220 36964 4276 36966
rect 4300 36964 4356 36966
rect 4380 36964 4436 36966
rect 4460 36964 4516 36966
rect 4220 35930 4276 35932
rect 4300 35930 4356 35932
rect 4380 35930 4436 35932
rect 4460 35930 4516 35932
rect 4220 35878 4246 35930
rect 4246 35878 4276 35930
rect 4300 35878 4310 35930
rect 4310 35878 4356 35930
rect 4380 35878 4426 35930
rect 4426 35878 4436 35930
rect 4460 35878 4490 35930
rect 4490 35878 4516 35930
rect 4220 35876 4276 35878
rect 4300 35876 4356 35878
rect 4380 35876 4436 35878
rect 4460 35876 4516 35878
rect 4066 34856 4122 34912
rect 4220 34842 4276 34844
rect 4300 34842 4356 34844
rect 4380 34842 4436 34844
rect 4460 34842 4516 34844
rect 4220 34790 4246 34842
rect 4246 34790 4276 34842
rect 4300 34790 4310 34842
rect 4310 34790 4356 34842
rect 4380 34790 4426 34842
rect 4426 34790 4436 34842
rect 4460 34790 4490 34842
rect 4490 34790 4516 34842
rect 4220 34788 4276 34790
rect 4300 34788 4356 34790
rect 4380 34788 4436 34790
rect 4460 34788 4516 34790
rect 4220 33754 4276 33756
rect 4300 33754 4356 33756
rect 4380 33754 4436 33756
rect 4460 33754 4516 33756
rect 4220 33702 4246 33754
rect 4246 33702 4276 33754
rect 4300 33702 4310 33754
rect 4310 33702 4356 33754
rect 4380 33702 4426 33754
rect 4426 33702 4436 33754
rect 4460 33702 4490 33754
rect 4490 33702 4516 33754
rect 4220 33700 4276 33702
rect 4300 33700 4356 33702
rect 4380 33700 4436 33702
rect 4460 33700 4516 33702
rect 4220 32666 4276 32668
rect 4300 32666 4356 32668
rect 4380 32666 4436 32668
rect 4460 32666 4516 32668
rect 4220 32614 4246 32666
rect 4246 32614 4276 32666
rect 4300 32614 4310 32666
rect 4310 32614 4356 32666
rect 4380 32614 4426 32666
rect 4426 32614 4436 32666
rect 4460 32614 4490 32666
rect 4490 32614 4516 32666
rect 4220 32612 4276 32614
rect 4300 32612 4356 32614
rect 4380 32612 4436 32614
rect 4460 32612 4516 32614
rect 4220 31578 4276 31580
rect 4300 31578 4356 31580
rect 4380 31578 4436 31580
rect 4460 31578 4516 31580
rect 4220 31526 4246 31578
rect 4246 31526 4276 31578
rect 4300 31526 4310 31578
rect 4310 31526 4356 31578
rect 4380 31526 4426 31578
rect 4426 31526 4436 31578
rect 4460 31526 4490 31578
rect 4490 31526 4516 31578
rect 4220 31524 4276 31526
rect 4300 31524 4356 31526
rect 4380 31524 4436 31526
rect 4460 31524 4516 31526
rect 4220 30490 4276 30492
rect 4300 30490 4356 30492
rect 4380 30490 4436 30492
rect 4460 30490 4516 30492
rect 4220 30438 4246 30490
rect 4246 30438 4276 30490
rect 4300 30438 4310 30490
rect 4310 30438 4356 30490
rect 4380 30438 4426 30490
rect 4426 30438 4436 30490
rect 4460 30438 4490 30490
rect 4490 30438 4516 30490
rect 4220 30436 4276 30438
rect 4300 30436 4356 30438
rect 4380 30436 4436 30438
rect 4460 30436 4516 30438
rect 4220 29402 4276 29404
rect 4300 29402 4356 29404
rect 4380 29402 4436 29404
rect 4460 29402 4516 29404
rect 4220 29350 4246 29402
rect 4246 29350 4276 29402
rect 4300 29350 4310 29402
rect 4310 29350 4356 29402
rect 4380 29350 4426 29402
rect 4426 29350 4436 29402
rect 4460 29350 4490 29402
rect 4490 29350 4516 29402
rect 4220 29348 4276 29350
rect 4300 29348 4356 29350
rect 4380 29348 4436 29350
rect 4460 29348 4516 29350
rect 3974 29008 4030 29064
rect 4220 28314 4276 28316
rect 4300 28314 4356 28316
rect 4380 28314 4436 28316
rect 4460 28314 4516 28316
rect 4220 28262 4246 28314
rect 4246 28262 4276 28314
rect 4300 28262 4310 28314
rect 4310 28262 4356 28314
rect 4380 28262 4426 28314
rect 4426 28262 4436 28314
rect 4460 28262 4490 28314
rect 4490 28262 4516 28314
rect 4220 28260 4276 28262
rect 4300 28260 4356 28262
rect 4380 28260 4436 28262
rect 4460 28260 4516 28262
rect 4220 27226 4276 27228
rect 4300 27226 4356 27228
rect 4380 27226 4436 27228
rect 4460 27226 4516 27228
rect 4220 27174 4246 27226
rect 4246 27174 4276 27226
rect 4300 27174 4310 27226
rect 4310 27174 4356 27226
rect 4380 27174 4426 27226
rect 4426 27174 4436 27226
rect 4460 27174 4490 27226
rect 4490 27174 4516 27226
rect 4220 27172 4276 27174
rect 4300 27172 4356 27174
rect 4380 27172 4436 27174
rect 4460 27172 4516 27174
rect 4220 26138 4276 26140
rect 4300 26138 4356 26140
rect 4380 26138 4436 26140
rect 4460 26138 4516 26140
rect 4220 26086 4246 26138
rect 4246 26086 4276 26138
rect 4300 26086 4310 26138
rect 4310 26086 4356 26138
rect 4380 26086 4426 26138
rect 4426 26086 4436 26138
rect 4460 26086 4490 26138
rect 4490 26086 4516 26138
rect 4220 26084 4276 26086
rect 4300 26084 4356 26086
rect 4380 26084 4436 26086
rect 4460 26084 4516 26086
rect 4220 25050 4276 25052
rect 4300 25050 4356 25052
rect 4380 25050 4436 25052
rect 4460 25050 4516 25052
rect 4220 24998 4246 25050
rect 4246 24998 4276 25050
rect 4300 24998 4310 25050
rect 4310 24998 4356 25050
rect 4380 24998 4426 25050
rect 4426 24998 4436 25050
rect 4460 24998 4490 25050
rect 4490 24998 4516 25050
rect 4220 24996 4276 24998
rect 4300 24996 4356 24998
rect 4380 24996 4436 24998
rect 4460 24996 4516 24998
rect 4220 23962 4276 23964
rect 4300 23962 4356 23964
rect 4380 23962 4436 23964
rect 4460 23962 4516 23964
rect 4220 23910 4246 23962
rect 4246 23910 4276 23962
rect 4300 23910 4310 23962
rect 4310 23910 4356 23962
rect 4380 23910 4426 23962
rect 4426 23910 4436 23962
rect 4460 23910 4490 23962
rect 4490 23910 4516 23962
rect 4220 23908 4276 23910
rect 4300 23908 4356 23910
rect 4380 23908 4436 23910
rect 4460 23908 4516 23910
rect 4220 22874 4276 22876
rect 4300 22874 4356 22876
rect 4380 22874 4436 22876
rect 4460 22874 4516 22876
rect 4220 22822 4246 22874
rect 4246 22822 4276 22874
rect 4300 22822 4310 22874
rect 4310 22822 4356 22874
rect 4380 22822 4426 22874
rect 4426 22822 4436 22874
rect 4460 22822 4490 22874
rect 4490 22822 4516 22874
rect 4220 22820 4276 22822
rect 4300 22820 4356 22822
rect 4380 22820 4436 22822
rect 4460 22820 4516 22822
rect 4220 21786 4276 21788
rect 4300 21786 4356 21788
rect 4380 21786 4436 21788
rect 4460 21786 4516 21788
rect 4220 21734 4246 21786
rect 4246 21734 4276 21786
rect 4300 21734 4310 21786
rect 4310 21734 4356 21786
rect 4380 21734 4426 21786
rect 4426 21734 4436 21786
rect 4460 21734 4490 21786
rect 4490 21734 4516 21786
rect 4220 21732 4276 21734
rect 4300 21732 4356 21734
rect 4380 21732 4436 21734
rect 4460 21732 4516 21734
rect 6182 25780 6184 25800
rect 6184 25780 6236 25800
rect 6236 25780 6238 25800
rect 6182 25744 6238 25780
rect 4220 20698 4276 20700
rect 4300 20698 4356 20700
rect 4380 20698 4436 20700
rect 4460 20698 4516 20700
rect 4220 20646 4246 20698
rect 4246 20646 4276 20698
rect 4300 20646 4310 20698
rect 4310 20646 4356 20698
rect 4380 20646 4426 20698
rect 4426 20646 4436 20698
rect 4460 20646 4490 20698
rect 4490 20646 4516 20698
rect 4220 20644 4276 20646
rect 4300 20644 4356 20646
rect 4380 20644 4436 20646
rect 4460 20644 4516 20646
rect 4220 19610 4276 19612
rect 4300 19610 4356 19612
rect 4380 19610 4436 19612
rect 4460 19610 4516 19612
rect 4220 19558 4246 19610
rect 4246 19558 4276 19610
rect 4300 19558 4310 19610
rect 4310 19558 4356 19610
rect 4380 19558 4426 19610
rect 4426 19558 4436 19610
rect 4460 19558 4490 19610
rect 4490 19558 4516 19610
rect 4220 19556 4276 19558
rect 4300 19556 4356 19558
rect 4380 19556 4436 19558
rect 4460 19556 4516 19558
rect 4220 18522 4276 18524
rect 4300 18522 4356 18524
rect 4380 18522 4436 18524
rect 4460 18522 4516 18524
rect 4220 18470 4246 18522
rect 4246 18470 4276 18522
rect 4300 18470 4310 18522
rect 4310 18470 4356 18522
rect 4380 18470 4426 18522
rect 4426 18470 4436 18522
rect 4460 18470 4490 18522
rect 4490 18470 4516 18522
rect 4220 18468 4276 18470
rect 4300 18468 4356 18470
rect 4380 18468 4436 18470
rect 4460 18468 4516 18470
rect 10046 29552 10102 29608
rect 9402 29144 9458 29200
rect 4220 17434 4276 17436
rect 4300 17434 4356 17436
rect 4380 17434 4436 17436
rect 4460 17434 4516 17436
rect 4220 17382 4246 17434
rect 4246 17382 4276 17434
rect 4300 17382 4310 17434
rect 4310 17382 4356 17434
rect 4380 17382 4426 17434
rect 4426 17382 4436 17434
rect 4460 17382 4490 17434
rect 4490 17382 4516 17434
rect 4220 17380 4276 17382
rect 4300 17380 4356 17382
rect 4380 17380 4436 17382
rect 4460 17380 4516 17382
rect 4220 16346 4276 16348
rect 4300 16346 4356 16348
rect 4380 16346 4436 16348
rect 4460 16346 4516 16348
rect 4220 16294 4246 16346
rect 4246 16294 4276 16346
rect 4300 16294 4310 16346
rect 4310 16294 4356 16346
rect 4380 16294 4426 16346
rect 4426 16294 4436 16346
rect 4460 16294 4490 16346
rect 4490 16294 4516 16346
rect 4220 16292 4276 16294
rect 4300 16292 4356 16294
rect 4380 16292 4436 16294
rect 4460 16292 4516 16294
rect 4220 15258 4276 15260
rect 4300 15258 4356 15260
rect 4380 15258 4436 15260
rect 4460 15258 4516 15260
rect 4220 15206 4246 15258
rect 4246 15206 4276 15258
rect 4300 15206 4310 15258
rect 4310 15206 4356 15258
rect 4380 15206 4426 15258
rect 4426 15206 4436 15258
rect 4460 15206 4490 15258
rect 4490 15206 4516 15258
rect 4220 15204 4276 15206
rect 4300 15204 4356 15206
rect 4380 15204 4436 15206
rect 4460 15204 4516 15206
rect 4066 15000 4122 15056
rect 3882 14592 3938 14648
rect 5078 14456 5134 14512
rect 4220 14170 4276 14172
rect 4300 14170 4356 14172
rect 4380 14170 4436 14172
rect 4460 14170 4516 14172
rect 4220 14118 4246 14170
rect 4246 14118 4276 14170
rect 4300 14118 4310 14170
rect 4310 14118 4356 14170
rect 4380 14118 4426 14170
rect 4426 14118 4436 14170
rect 4460 14118 4490 14170
rect 4490 14118 4516 14170
rect 4220 14116 4276 14118
rect 4300 14116 4356 14118
rect 4380 14116 4436 14118
rect 4460 14116 4516 14118
rect 4220 13082 4276 13084
rect 4300 13082 4356 13084
rect 4380 13082 4436 13084
rect 4460 13082 4516 13084
rect 4220 13030 4246 13082
rect 4246 13030 4276 13082
rect 4300 13030 4310 13082
rect 4310 13030 4356 13082
rect 4380 13030 4426 13082
rect 4426 13030 4436 13082
rect 4460 13030 4490 13082
rect 4490 13030 4516 13082
rect 4220 13028 4276 13030
rect 4300 13028 4356 13030
rect 4380 13028 4436 13030
rect 4460 13028 4516 13030
rect 4220 11994 4276 11996
rect 4300 11994 4356 11996
rect 4380 11994 4436 11996
rect 4460 11994 4516 11996
rect 4220 11942 4246 11994
rect 4246 11942 4276 11994
rect 4300 11942 4310 11994
rect 4310 11942 4356 11994
rect 4380 11942 4426 11994
rect 4426 11942 4436 11994
rect 4460 11942 4490 11994
rect 4490 11942 4516 11994
rect 4220 11940 4276 11942
rect 4300 11940 4356 11942
rect 4380 11940 4436 11942
rect 4460 11940 4516 11942
rect 4220 10906 4276 10908
rect 4300 10906 4356 10908
rect 4380 10906 4436 10908
rect 4460 10906 4516 10908
rect 4220 10854 4246 10906
rect 4246 10854 4276 10906
rect 4300 10854 4310 10906
rect 4310 10854 4356 10906
rect 4380 10854 4426 10906
rect 4426 10854 4436 10906
rect 4460 10854 4490 10906
rect 4490 10854 4516 10906
rect 4220 10852 4276 10854
rect 4300 10852 4356 10854
rect 4380 10852 4436 10854
rect 4460 10852 4516 10854
rect 9494 18672 9550 18728
rect 4220 9818 4276 9820
rect 4300 9818 4356 9820
rect 4380 9818 4436 9820
rect 4460 9818 4516 9820
rect 4220 9766 4246 9818
rect 4246 9766 4276 9818
rect 4300 9766 4310 9818
rect 4310 9766 4356 9818
rect 4380 9766 4426 9818
rect 4426 9766 4436 9818
rect 4460 9766 4490 9818
rect 4490 9766 4516 9818
rect 4220 9764 4276 9766
rect 4300 9764 4356 9766
rect 4380 9764 4436 9766
rect 4460 9764 4516 9766
rect 4066 9288 4122 9344
rect 4220 8730 4276 8732
rect 4300 8730 4356 8732
rect 4380 8730 4436 8732
rect 4460 8730 4516 8732
rect 4220 8678 4246 8730
rect 4246 8678 4276 8730
rect 4300 8678 4310 8730
rect 4310 8678 4356 8730
rect 4380 8678 4426 8730
rect 4426 8678 4436 8730
rect 4460 8678 4490 8730
rect 4490 8678 4516 8730
rect 4220 8676 4276 8678
rect 4300 8676 4356 8678
rect 4380 8676 4436 8678
rect 4460 8676 4516 8678
rect 4220 7642 4276 7644
rect 4300 7642 4356 7644
rect 4380 7642 4436 7644
rect 4460 7642 4516 7644
rect 4220 7590 4246 7642
rect 4246 7590 4276 7642
rect 4300 7590 4310 7642
rect 4310 7590 4356 7642
rect 4380 7590 4426 7642
rect 4426 7590 4436 7642
rect 4460 7590 4490 7642
rect 4490 7590 4516 7642
rect 4220 7588 4276 7590
rect 4300 7588 4356 7590
rect 4380 7588 4436 7590
rect 4460 7588 4516 7590
rect 9494 14612 9550 14648
rect 9494 14592 9496 14612
rect 9496 14592 9548 14612
rect 9548 14592 9550 14612
rect 4220 6554 4276 6556
rect 4300 6554 4356 6556
rect 4380 6554 4436 6556
rect 4460 6554 4516 6556
rect 4220 6502 4246 6554
rect 4246 6502 4276 6554
rect 4300 6502 4310 6554
rect 4310 6502 4356 6554
rect 4380 6502 4426 6554
rect 4426 6502 4436 6554
rect 4460 6502 4490 6554
rect 4490 6502 4516 6554
rect 4220 6500 4276 6502
rect 4300 6500 4356 6502
rect 4380 6500 4436 6502
rect 4460 6500 4516 6502
rect 3974 6296 4030 6352
rect 4220 5466 4276 5468
rect 4300 5466 4356 5468
rect 4380 5466 4436 5468
rect 4460 5466 4516 5468
rect 4220 5414 4246 5466
rect 4246 5414 4276 5466
rect 4300 5414 4310 5466
rect 4310 5414 4356 5466
rect 4380 5414 4426 5466
rect 4426 5414 4436 5466
rect 4460 5414 4490 5466
rect 4490 5414 4516 5466
rect 4220 5412 4276 5414
rect 4300 5412 4356 5414
rect 4380 5412 4436 5414
rect 4460 5412 4516 5414
rect 4220 4378 4276 4380
rect 4300 4378 4356 4380
rect 4380 4378 4436 4380
rect 4460 4378 4516 4380
rect 4220 4326 4246 4378
rect 4246 4326 4276 4378
rect 4300 4326 4310 4378
rect 4310 4326 4356 4378
rect 4380 4326 4426 4378
rect 4426 4326 4436 4378
rect 4460 4326 4490 4378
rect 4490 4326 4516 4378
rect 4220 4324 4276 4326
rect 4300 4324 4356 4326
rect 4380 4324 4436 4326
rect 4460 4324 4516 4326
rect 3422 3576 3478 3632
rect 6274 3304 6330 3360
rect 4220 3290 4276 3292
rect 4300 3290 4356 3292
rect 4380 3290 4436 3292
rect 4460 3290 4516 3292
rect 4220 3238 4246 3290
rect 4246 3238 4276 3290
rect 4300 3238 4310 3290
rect 4310 3238 4356 3290
rect 4380 3238 4426 3290
rect 4426 3238 4436 3290
rect 4460 3238 4490 3290
rect 4490 3238 4516 3290
rect 4220 3236 4276 3238
rect 4300 3236 4356 3238
rect 4380 3236 4436 3238
rect 4460 3236 4516 3238
rect 4220 2202 4276 2204
rect 4300 2202 4356 2204
rect 4380 2202 4436 2204
rect 4460 2202 4516 2204
rect 4220 2150 4246 2202
rect 4246 2150 4276 2202
rect 4300 2150 4310 2202
rect 4310 2150 4356 2202
rect 4380 2150 4426 2202
rect 4426 2150 4436 2202
rect 4460 2150 4490 2202
rect 4490 2150 4516 2202
rect 4220 2148 4276 2150
rect 4300 2148 4356 2150
rect 4380 2148 4436 2150
rect 4460 2148 4516 2150
rect 7286 2932 7288 2952
rect 7288 2932 7340 2952
rect 7340 2932 7342 2952
rect 7286 2896 7342 2932
rect 8114 3440 8170 3496
rect 10046 9560 10102 9616
rect 9862 7792 9918 7848
rect 10598 36624 10654 36680
rect 10506 29708 10562 29744
rect 10506 29688 10508 29708
rect 10508 29688 10560 29708
rect 10560 29688 10562 29708
rect 10690 29552 10746 29608
rect 12622 29724 12624 29744
rect 12624 29724 12676 29744
rect 12676 29724 12678 29744
rect 12622 29688 12678 29724
rect 12898 29572 12954 29608
rect 12898 29552 12900 29572
rect 12900 29552 12952 29572
rect 12952 29552 12954 29572
rect 11242 11212 11298 11248
rect 11242 11192 11244 11212
rect 11244 11192 11296 11212
rect 11296 11192 11298 11212
rect 11242 9832 11298 9888
rect 11518 12300 11574 12336
rect 11518 12280 11520 12300
rect 11520 12280 11572 12300
rect 11572 12280 11574 12300
rect 10874 7384 10930 7440
rect 9586 2916 9642 2952
rect 9586 2896 9588 2916
rect 9588 2896 9640 2916
rect 9640 2896 9642 2916
rect 12254 9560 12310 9616
rect 12530 9596 12532 9616
rect 12532 9596 12584 9616
rect 12584 9596 12586 9616
rect 12530 9560 12586 9596
rect 12530 9460 12532 9480
rect 12532 9460 12584 9480
rect 12584 9460 12586 9480
rect 12530 9424 12586 9460
rect 12898 9424 12954 9480
rect 14462 7384 14518 7440
rect 15106 8472 15162 8528
rect 19580 38650 19636 38652
rect 19660 38650 19716 38652
rect 19740 38650 19796 38652
rect 19820 38650 19876 38652
rect 19580 38598 19606 38650
rect 19606 38598 19636 38650
rect 19660 38598 19670 38650
rect 19670 38598 19716 38650
rect 19740 38598 19786 38650
rect 19786 38598 19796 38650
rect 19820 38598 19850 38650
rect 19850 38598 19876 38650
rect 19580 38596 19636 38598
rect 19660 38596 19716 38598
rect 19740 38596 19796 38598
rect 19820 38596 19876 38598
rect 16578 36624 16634 36680
rect 19580 37562 19636 37564
rect 19660 37562 19716 37564
rect 19740 37562 19796 37564
rect 19820 37562 19876 37564
rect 19580 37510 19606 37562
rect 19606 37510 19636 37562
rect 19660 37510 19670 37562
rect 19670 37510 19716 37562
rect 19740 37510 19786 37562
rect 19786 37510 19796 37562
rect 19820 37510 19850 37562
rect 19850 37510 19876 37562
rect 19580 37508 19636 37510
rect 19660 37508 19716 37510
rect 19740 37508 19796 37510
rect 19820 37508 19876 37510
rect 19798 36660 19800 36680
rect 19800 36660 19852 36680
rect 19852 36660 19854 36680
rect 19798 36624 19854 36660
rect 19580 36474 19636 36476
rect 19660 36474 19716 36476
rect 19740 36474 19796 36476
rect 19820 36474 19876 36476
rect 19580 36422 19606 36474
rect 19606 36422 19636 36474
rect 19660 36422 19670 36474
rect 19670 36422 19716 36474
rect 19740 36422 19786 36474
rect 19786 36422 19796 36474
rect 19820 36422 19850 36474
rect 19850 36422 19876 36474
rect 19580 36420 19636 36422
rect 19660 36420 19716 36422
rect 19740 36420 19796 36422
rect 19820 36420 19876 36422
rect 19580 35386 19636 35388
rect 19660 35386 19716 35388
rect 19740 35386 19796 35388
rect 19820 35386 19876 35388
rect 19580 35334 19606 35386
rect 19606 35334 19636 35386
rect 19660 35334 19670 35386
rect 19670 35334 19716 35386
rect 19740 35334 19786 35386
rect 19786 35334 19796 35386
rect 19820 35334 19850 35386
rect 19850 35334 19876 35386
rect 19580 35332 19636 35334
rect 19660 35332 19716 35334
rect 19740 35332 19796 35334
rect 19820 35332 19876 35334
rect 19580 34298 19636 34300
rect 19660 34298 19716 34300
rect 19740 34298 19796 34300
rect 19820 34298 19876 34300
rect 19580 34246 19606 34298
rect 19606 34246 19636 34298
rect 19660 34246 19670 34298
rect 19670 34246 19716 34298
rect 19740 34246 19786 34298
rect 19786 34246 19796 34298
rect 19820 34246 19850 34298
rect 19850 34246 19876 34298
rect 19580 34244 19636 34246
rect 19660 34244 19716 34246
rect 19740 34244 19796 34246
rect 19820 34244 19876 34246
rect 19580 33210 19636 33212
rect 19660 33210 19716 33212
rect 19740 33210 19796 33212
rect 19820 33210 19876 33212
rect 19580 33158 19606 33210
rect 19606 33158 19636 33210
rect 19660 33158 19670 33210
rect 19670 33158 19716 33210
rect 19740 33158 19786 33210
rect 19786 33158 19796 33210
rect 19820 33158 19850 33210
rect 19850 33158 19876 33210
rect 19580 33156 19636 33158
rect 19660 33156 19716 33158
rect 19740 33156 19796 33158
rect 19820 33156 19876 33158
rect 18418 32136 18474 32192
rect 18786 29180 18788 29200
rect 18788 29180 18840 29200
rect 18840 29180 18842 29200
rect 18786 29144 18842 29180
rect 16302 20304 16358 20360
rect 16762 12280 16818 12336
rect 16670 9560 16726 9616
rect 17406 9832 17462 9888
rect 19154 32136 19210 32192
rect 19580 32122 19636 32124
rect 19660 32122 19716 32124
rect 19740 32122 19796 32124
rect 19820 32122 19876 32124
rect 19580 32070 19606 32122
rect 19606 32070 19636 32122
rect 19660 32070 19670 32122
rect 19670 32070 19716 32122
rect 19740 32070 19786 32122
rect 19786 32070 19796 32122
rect 19820 32070 19850 32122
rect 19850 32070 19876 32122
rect 19580 32068 19636 32070
rect 19660 32068 19716 32070
rect 19740 32068 19796 32070
rect 19820 32068 19876 32070
rect 19154 18164 19156 18184
rect 19156 18164 19208 18184
rect 19208 18164 19210 18184
rect 19154 18128 19210 18164
rect 19338 31884 19394 31920
rect 19338 31864 19340 31884
rect 19340 31864 19392 31884
rect 19392 31864 19394 31884
rect 20902 37324 20958 37360
rect 20902 37304 20904 37324
rect 20904 37304 20956 37324
rect 20956 37304 20958 37324
rect 21730 36624 21786 36680
rect 22926 37324 22982 37360
rect 22926 37304 22928 37324
rect 22928 37304 22980 37324
rect 22980 37304 22982 37324
rect 19580 31034 19636 31036
rect 19660 31034 19716 31036
rect 19740 31034 19796 31036
rect 19820 31034 19876 31036
rect 19580 30982 19606 31034
rect 19606 30982 19636 31034
rect 19660 30982 19670 31034
rect 19670 30982 19716 31034
rect 19740 30982 19786 31034
rect 19786 30982 19796 31034
rect 19820 30982 19850 31034
rect 19850 30982 19876 31034
rect 19580 30980 19636 30982
rect 19660 30980 19716 30982
rect 19740 30980 19796 30982
rect 19820 30980 19876 30982
rect 19798 30132 19800 30152
rect 19800 30132 19852 30152
rect 19852 30132 19854 30152
rect 19798 30096 19854 30132
rect 19580 29946 19636 29948
rect 19660 29946 19716 29948
rect 19740 29946 19796 29948
rect 19820 29946 19876 29948
rect 19580 29894 19606 29946
rect 19606 29894 19636 29946
rect 19660 29894 19670 29946
rect 19670 29894 19716 29946
rect 19740 29894 19786 29946
rect 19786 29894 19796 29946
rect 19820 29894 19850 29946
rect 19850 29894 19876 29946
rect 19580 29892 19636 29894
rect 19660 29892 19716 29894
rect 19740 29892 19796 29894
rect 19820 29892 19876 29894
rect 19614 29588 19616 29608
rect 19616 29588 19668 29608
rect 19668 29588 19670 29608
rect 19614 29552 19670 29588
rect 19982 29552 20038 29608
rect 19798 29280 19854 29336
rect 19430 28872 19486 28928
rect 19580 28858 19636 28860
rect 19660 28858 19716 28860
rect 19740 28858 19796 28860
rect 19820 28858 19876 28860
rect 19580 28806 19606 28858
rect 19606 28806 19636 28858
rect 19660 28806 19670 28858
rect 19670 28806 19716 28858
rect 19740 28806 19786 28858
rect 19786 28806 19796 28858
rect 19820 28806 19850 28858
rect 19850 28806 19876 28858
rect 19580 28804 19636 28806
rect 19660 28804 19716 28806
rect 19740 28804 19796 28806
rect 19820 28804 19876 28806
rect 19338 28464 19394 28520
rect 19580 27770 19636 27772
rect 19660 27770 19716 27772
rect 19740 27770 19796 27772
rect 19820 27770 19876 27772
rect 19580 27718 19606 27770
rect 19606 27718 19636 27770
rect 19660 27718 19670 27770
rect 19670 27718 19716 27770
rect 19740 27718 19786 27770
rect 19786 27718 19796 27770
rect 19820 27718 19850 27770
rect 19850 27718 19876 27770
rect 19580 27716 19636 27718
rect 19660 27716 19716 27718
rect 19740 27716 19796 27718
rect 19820 27716 19876 27718
rect 19580 26682 19636 26684
rect 19660 26682 19716 26684
rect 19740 26682 19796 26684
rect 19820 26682 19876 26684
rect 19580 26630 19606 26682
rect 19606 26630 19636 26682
rect 19660 26630 19670 26682
rect 19670 26630 19716 26682
rect 19740 26630 19786 26682
rect 19786 26630 19796 26682
rect 19820 26630 19850 26682
rect 19850 26630 19876 26682
rect 19580 26628 19636 26630
rect 19660 26628 19716 26630
rect 19740 26628 19796 26630
rect 19820 26628 19876 26630
rect 19580 25594 19636 25596
rect 19660 25594 19716 25596
rect 19740 25594 19796 25596
rect 19820 25594 19876 25596
rect 19580 25542 19606 25594
rect 19606 25542 19636 25594
rect 19660 25542 19670 25594
rect 19670 25542 19716 25594
rect 19740 25542 19786 25594
rect 19786 25542 19796 25594
rect 19820 25542 19850 25594
rect 19850 25542 19876 25594
rect 19580 25540 19636 25542
rect 19660 25540 19716 25542
rect 19740 25540 19796 25542
rect 19820 25540 19876 25542
rect 19580 24506 19636 24508
rect 19660 24506 19716 24508
rect 19740 24506 19796 24508
rect 19820 24506 19876 24508
rect 19580 24454 19606 24506
rect 19606 24454 19636 24506
rect 19660 24454 19670 24506
rect 19670 24454 19716 24506
rect 19740 24454 19786 24506
rect 19786 24454 19796 24506
rect 19820 24454 19850 24506
rect 19850 24454 19876 24506
rect 19580 24452 19636 24454
rect 19660 24452 19716 24454
rect 19740 24452 19796 24454
rect 19820 24452 19876 24454
rect 19580 23418 19636 23420
rect 19660 23418 19716 23420
rect 19740 23418 19796 23420
rect 19820 23418 19876 23420
rect 19580 23366 19606 23418
rect 19606 23366 19636 23418
rect 19660 23366 19670 23418
rect 19670 23366 19716 23418
rect 19740 23366 19786 23418
rect 19786 23366 19796 23418
rect 19820 23366 19850 23418
rect 19850 23366 19876 23418
rect 19580 23364 19636 23366
rect 19660 23364 19716 23366
rect 19740 23364 19796 23366
rect 19820 23364 19876 23366
rect 19430 23316 19486 23352
rect 19430 23296 19432 23316
rect 19432 23296 19484 23316
rect 19484 23296 19486 23316
rect 20350 31884 20406 31920
rect 20350 31864 20352 31884
rect 20352 31864 20404 31884
rect 20404 31864 20406 31884
rect 20166 29280 20222 29336
rect 19580 22330 19636 22332
rect 19660 22330 19716 22332
rect 19740 22330 19796 22332
rect 19820 22330 19876 22332
rect 19580 22278 19606 22330
rect 19606 22278 19636 22330
rect 19660 22278 19670 22330
rect 19670 22278 19716 22330
rect 19740 22278 19786 22330
rect 19786 22278 19796 22330
rect 19820 22278 19850 22330
rect 19850 22278 19876 22330
rect 19580 22276 19636 22278
rect 19660 22276 19716 22278
rect 19740 22276 19796 22278
rect 19820 22276 19876 22278
rect 19580 21242 19636 21244
rect 19660 21242 19716 21244
rect 19740 21242 19796 21244
rect 19820 21242 19876 21244
rect 19580 21190 19606 21242
rect 19606 21190 19636 21242
rect 19660 21190 19670 21242
rect 19670 21190 19716 21242
rect 19740 21190 19786 21242
rect 19786 21190 19796 21242
rect 19820 21190 19850 21242
rect 19850 21190 19876 21242
rect 19580 21188 19636 21190
rect 19660 21188 19716 21190
rect 19740 21188 19796 21190
rect 19820 21188 19876 21190
rect 19580 20154 19636 20156
rect 19660 20154 19716 20156
rect 19740 20154 19796 20156
rect 19820 20154 19876 20156
rect 19580 20102 19606 20154
rect 19606 20102 19636 20154
rect 19660 20102 19670 20154
rect 19670 20102 19716 20154
rect 19740 20102 19786 20154
rect 19786 20102 19796 20154
rect 19820 20102 19850 20154
rect 19850 20102 19876 20154
rect 19580 20100 19636 20102
rect 19660 20100 19716 20102
rect 19740 20100 19796 20102
rect 19820 20100 19876 20102
rect 19430 19896 19486 19952
rect 19706 19932 19708 19952
rect 19708 19932 19760 19952
rect 19760 19932 19762 19952
rect 19706 19896 19762 19932
rect 19982 19488 20038 19544
rect 19580 19066 19636 19068
rect 19660 19066 19716 19068
rect 19740 19066 19796 19068
rect 19820 19066 19876 19068
rect 19580 19014 19606 19066
rect 19606 19014 19636 19066
rect 19660 19014 19670 19066
rect 19670 19014 19716 19066
rect 19740 19014 19786 19066
rect 19786 19014 19796 19066
rect 19820 19014 19850 19066
rect 19850 19014 19876 19066
rect 19580 19012 19636 19014
rect 19660 19012 19716 19014
rect 19740 19012 19796 19014
rect 19820 19012 19876 19014
rect 19522 18844 19524 18864
rect 19524 18844 19576 18864
rect 19576 18844 19578 18864
rect 19522 18808 19578 18844
rect 19614 18672 19670 18728
rect 19706 18128 19762 18184
rect 19580 17978 19636 17980
rect 19660 17978 19716 17980
rect 19740 17978 19796 17980
rect 19820 17978 19876 17980
rect 19580 17926 19606 17978
rect 19606 17926 19636 17978
rect 19660 17926 19670 17978
rect 19670 17926 19716 17978
rect 19740 17926 19786 17978
rect 19786 17926 19796 17978
rect 19820 17926 19850 17978
rect 19850 17926 19876 17978
rect 19580 17924 19636 17926
rect 19660 17924 19716 17926
rect 19740 17924 19796 17926
rect 19820 17924 19876 17926
rect 19580 16890 19636 16892
rect 19660 16890 19716 16892
rect 19740 16890 19796 16892
rect 19820 16890 19876 16892
rect 19580 16838 19606 16890
rect 19606 16838 19636 16890
rect 19660 16838 19670 16890
rect 19670 16838 19716 16890
rect 19740 16838 19786 16890
rect 19786 16838 19796 16890
rect 19820 16838 19850 16890
rect 19850 16838 19876 16890
rect 19580 16836 19636 16838
rect 19660 16836 19716 16838
rect 19740 16836 19796 16838
rect 19820 16836 19876 16838
rect 19580 15802 19636 15804
rect 19660 15802 19716 15804
rect 19740 15802 19796 15804
rect 19820 15802 19876 15804
rect 19580 15750 19606 15802
rect 19606 15750 19636 15802
rect 19660 15750 19670 15802
rect 19670 15750 19716 15802
rect 19740 15750 19786 15802
rect 19786 15750 19796 15802
rect 19820 15750 19850 15802
rect 19850 15750 19876 15802
rect 19580 15748 19636 15750
rect 19660 15748 19716 15750
rect 19740 15748 19796 15750
rect 19820 15748 19876 15750
rect 20166 19488 20222 19544
rect 20718 30096 20774 30152
rect 20534 18808 20590 18864
rect 19580 14714 19636 14716
rect 19660 14714 19716 14716
rect 19740 14714 19796 14716
rect 19820 14714 19876 14716
rect 19580 14662 19606 14714
rect 19606 14662 19636 14714
rect 19660 14662 19670 14714
rect 19670 14662 19716 14714
rect 19740 14662 19786 14714
rect 19786 14662 19796 14714
rect 19820 14662 19850 14714
rect 19850 14662 19876 14714
rect 19580 14660 19636 14662
rect 19660 14660 19716 14662
rect 19740 14660 19796 14662
rect 19820 14660 19876 14662
rect 19580 13626 19636 13628
rect 19660 13626 19716 13628
rect 19740 13626 19796 13628
rect 19820 13626 19876 13628
rect 19580 13574 19606 13626
rect 19606 13574 19636 13626
rect 19660 13574 19670 13626
rect 19670 13574 19716 13626
rect 19740 13574 19786 13626
rect 19786 13574 19796 13626
rect 19820 13574 19850 13626
rect 19850 13574 19876 13626
rect 19580 13572 19636 13574
rect 19660 13572 19716 13574
rect 19740 13572 19796 13574
rect 19820 13572 19876 13574
rect 19580 12538 19636 12540
rect 19660 12538 19716 12540
rect 19740 12538 19796 12540
rect 19820 12538 19876 12540
rect 19580 12486 19606 12538
rect 19606 12486 19636 12538
rect 19660 12486 19670 12538
rect 19670 12486 19716 12538
rect 19740 12486 19786 12538
rect 19786 12486 19796 12538
rect 19820 12486 19850 12538
rect 19850 12486 19876 12538
rect 19580 12484 19636 12486
rect 19660 12484 19716 12486
rect 19740 12484 19796 12486
rect 19820 12484 19876 12486
rect 19062 8372 19064 8392
rect 19064 8372 19116 8392
rect 19116 8372 19118 8392
rect 19062 8336 19118 8372
rect 19246 8336 19302 8392
rect 19580 11450 19636 11452
rect 19660 11450 19716 11452
rect 19740 11450 19796 11452
rect 19820 11450 19876 11452
rect 19580 11398 19606 11450
rect 19606 11398 19636 11450
rect 19660 11398 19670 11450
rect 19670 11398 19716 11450
rect 19740 11398 19786 11450
rect 19786 11398 19796 11450
rect 19820 11398 19850 11450
rect 19850 11398 19876 11450
rect 19580 11396 19636 11398
rect 19660 11396 19716 11398
rect 19740 11396 19796 11398
rect 19820 11396 19876 11398
rect 20258 11600 20314 11656
rect 19798 10784 19854 10840
rect 19580 10362 19636 10364
rect 19660 10362 19716 10364
rect 19740 10362 19796 10364
rect 19820 10362 19876 10364
rect 19580 10310 19606 10362
rect 19606 10310 19636 10362
rect 19660 10310 19670 10362
rect 19670 10310 19716 10362
rect 19740 10310 19786 10362
rect 19786 10310 19796 10362
rect 19820 10310 19850 10362
rect 19850 10310 19876 10362
rect 19580 10308 19636 10310
rect 19660 10308 19716 10310
rect 19740 10308 19796 10310
rect 19820 10308 19876 10310
rect 19890 9424 19946 9480
rect 19580 9274 19636 9276
rect 19660 9274 19716 9276
rect 19740 9274 19796 9276
rect 19820 9274 19876 9276
rect 19580 9222 19606 9274
rect 19606 9222 19636 9274
rect 19660 9222 19670 9274
rect 19670 9222 19716 9274
rect 19740 9222 19786 9274
rect 19786 9222 19796 9274
rect 19820 9222 19850 9274
rect 19850 9222 19876 9274
rect 19580 9220 19636 9222
rect 19660 9220 19716 9222
rect 19740 9220 19796 9222
rect 19820 9220 19876 9222
rect 19982 8608 20038 8664
rect 19580 8186 19636 8188
rect 19660 8186 19716 8188
rect 19740 8186 19796 8188
rect 19820 8186 19876 8188
rect 19580 8134 19606 8186
rect 19606 8134 19636 8186
rect 19660 8134 19670 8186
rect 19670 8134 19716 8186
rect 19740 8134 19786 8186
rect 19786 8134 19796 8186
rect 19820 8134 19850 8186
rect 19850 8134 19876 8186
rect 19580 8132 19636 8134
rect 19660 8132 19716 8134
rect 19740 8132 19796 8134
rect 19820 8132 19876 8134
rect 19246 6840 19302 6896
rect 19580 7098 19636 7100
rect 19660 7098 19716 7100
rect 19740 7098 19796 7100
rect 19820 7098 19876 7100
rect 19580 7046 19606 7098
rect 19606 7046 19636 7098
rect 19660 7046 19670 7098
rect 19670 7046 19716 7098
rect 19740 7046 19786 7098
rect 19786 7046 19796 7098
rect 19820 7046 19850 7098
rect 19850 7046 19876 7098
rect 19580 7044 19636 7046
rect 19660 7044 19716 7046
rect 19740 7044 19796 7046
rect 19820 7044 19876 7046
rect 21546 28076 21602 28112
rect 21546 28056 21548 28076
rect 21548 28056 21600 28076
rect 21600 28056 21602 28076
rect 21822 29144 21878 29200
rect 23294 31764 23296 31784
rect 23296 31764 23348 31784
rect 23348 31764 23350 31784
rect 23294 31728 23350 31764
rect 22926 29552 22982 29608
rect 21638 19352 21694 19408
rect 23294 29280 23350 29336
rect 22098 18672 22154 18728
rect 20718 11600 20774 11656
rect 19580 6010 19636 6012
rect 19660 6010 19716 6012
rect 19740 6010 19796 6012
rect 19820 6010 19876 6012
rect 19580 5958 19606 6010
rect 19606 5958 19636 6010
rect 19660 5958 19670 6010
rect 19670 5958 19716 6010
rect 19740 5958 19786 6010
rect 19786 5958 19796 6010
rect 19820 5958 19850 6010
rect 19850 5958 19876 6010
rect 19580 5956 19636 5958
rect 19660 5956 19716 5958
rect 19740 5956 19796 5958
rect 19820 5956 19876 5958
rect 17866 3576 17922 3632
rect 19580 4922 19636 4924
rect 19660 4922 19716 4924
rect 19740 4922 19796 4924
rect 19820 4922 19876 4924
rect 19580 4870 19606 4922
rect 19606 4870 19636 4922
rect 19660 4870 19670 4922
rect 19670 4870 19716 4922
rect 19740 4870 19786 4922
rect 19786 4870 19796 4922
rect 19820 4870 19850 4922
rect 19850 4870 19876 4922
rect 19580 4868 19636 4870
rect 19660 4868 19716 4870
rect 19740 4868 19796 4870
rect 19820 4868 19876 4870
rect 21178 8608 21234 8664
rect 21822 7928 21878 7984
rect 23018 19916 23074 19952
rect 23018 19896 23020 19916
rect 23020 19896 23072 19916
rect 23072 19896 23074 19916
rect 23938 29008 23994 29064
rect 24214 29572 24270 29608
rect 24214 29552 24216 29572
rect 24216 29552 24268 29572
rect 24268 29552 24270 29572
rect 24674 29280 24730 29336
rect 25226 30796 25282 30832
rect 25226 30776 25228 30796
rect 25228 30776 25280 30796
rect 25280 30776 25282 30796
rect 25502 31728 25558 31784
rect 22650 8336 22706 8392
rect 23018 7928 23074 7984
rect 19580 3834 19636 3836
rect 19660 3834 19716 3836
rect 19740 3834 19796 3836
rect 19820 3834 19876 3836
rect 19580 3782 19606 3834
rect 19606 3782 19636 3834
rect 19660 3782 19670 3834
rect 19670 3782 19716 3834
rect 19740 3782 19786 3834
rect 19786 3782 19796 3834
rect 19820 3782 19850 3834
rect 19850 3782 19876 3834
rect 19580 3780 19636 3782
rect 19660 3780 19716 3782
rect 19740 3780 19796 3782
rect 19820 3780 19876 3782
rect 21730 3984 21786 4040
rect 19580 2746 19636 2748
rect 19660 2746 19716 2748
rect 19740 2746 19796 2748
rect 19820 2746 19876 2748
rect 19580 2694 19606 2746
rect 19606 2694 19636 2746
rect 19660 2694 19670 2746
rect 19670 2694 19716 2746
rect 19740 2694 19786 2746
rect 19786 2694 19796 2746
rect 19820 2694 19850 2746
rect 19850 2694 19876 2746
rect 19580 2692 19636 2694
rect 19660 2692 19716 2694
rect 19740 2692 19796 2694
rect 19820 2692 19876 2694
rect 23662 9460 23664 9480
rect 23664 9460 23716 9480
rect 23716 9460 23718 9480
rect 23662 9424 23718 9460
rect 24398 11192 24454 11248
rect 24950 9560 25006 9616
rect 23662 7928 23718 7984
rect 27066 30640 27122 30696
rect 25502 18944 25558 19000
rect 25318 18536 25374 18592
rect 27618 29008 27674 29064
rect 27526 28464 27582 28520
rect 26422 22516 26424 22536
rect 26424 22516 26476 22536
rect 26476 22516 26478 22536
rect 26422 22480 26478 22516
rect 26882 22480 26938 22536
rect 27802 28076 27858 28112
rect 27802 28056 27804 28076
rect 27804 28056 27856 28076
rect 27856 28056 27858 28076
rect 27158 18672 27214 18728
rect 25502 10784 25558 10840
rect 25410 9424 25466 9480
rect 27434 18536 27490 18592
rect 26238 7792 26294 7848
rect 27618 19080 27674 19136
rect 28262 18808 28318 18864
rect 28538 22480 28594 22536
rect 29182 32408 29238 32464
rect 28814 19216 28870 19272
rect 28906 19080 28962 19136
rect 28722 18808 28778 18864
rect 28906 18672 28962 18728
rect 28538 18420 28594 18456
rect 28538 18400 28540 18420
rect 28540 18400 28592 18420
rect 28592 18400 28594 18420
rect 29090 19488 29146 19544
rect 28630 14456 28686 14512
rect 29642 19080 29698 19136
rect 29734 18944 29790 19000
rect 28446 3984 28502 4040
rect 28078 3440 28134 3496
rect 29090 6196 29092 6216
rect 29092 6196 29144 6216
rect 29144 6196 29146 6216
rect 29090 6160 29146 6196
rect 29734 9016 29790 9072
rect 30286 19488 30342 19544
rect 30010 18400 30066 18456
rect 30378 18672 30434 18728
rect 30838 19080 30894 19136
rect 29918 9152 29974 9208
rect 34940 38106 34996 38108
rect 35020 38106 35076 38108
rect 35100 38106 35156 38108
rect 35180 38106 35236 38108
rect 34940 38054 34966 38106
rect 34966 38054 34996 38106
rect 35020 38054 35030 38106
rect 35030 38054 35076 38106
rect 35100 38054 35146 38106
rect 35146 38054 35156 38106
rect 35180 38054 35210 38106
rect 35210 38054 35236 38106
rect 34940 38052 34996 38054
rect 35020 38052 35076 38054
rect 35100 38052 35156 38054
rect 35180 38052 35236 38054
rect 35898 38664 35954 38720
rect 34940 37018 34996 37020
rect 35020 37018 35076 37020
rect 35100 37018 35156 37020
rect 35180 37018 35236 37020
rect 34940 36966 34966 37018
rect 34966 36966 34996 37018
rect 35020 36966 35030 37018
rect 35030 36966 35076 37018
rect 35100 36966 35146 37018
rect 35146 36966 35156 37018
rect 35180 36966 35210 37018
rect 35210 36966 35236 37018
rect 34940 36964 34996 36966
rect 35020 36964 35076 36966
rect 35100 36964 35156 36966
rect 35180 36964 35236 36966
rect 31390 19252 31392 19272
rect 31392 19252 31444 19272
rect 31444 19252 31446 19272
rect 31390 19216 31446 19252
rect 31574 19352 31630 19408
rect 31666 18808 31722 18864
rect 34940 35930 34996 35932
rect 35020 35930 35076 35932
rect 35100 35930 35156 35932
rect 35180 35930 35236 35932
rect 34940 35878 34966 35930
rect 34966 35878 34996 35930
rect 35020 35878 35030 35930
rect 35030 35878 35076 35930
rect 35100 35878 35146 35930
rect 35146 35878 35156 35930
rect 35180 35878 35210 35930
rect 35210 35878 35236 35930
rect 34940 35876 34996 35878
rect 35020 35876 35076 35878
rect 35100 35876 35156 35878
rect 35180 35876 35236 35878
rect 34940 34842 34996 34844
rect 35020 34842 35076 34844
rect 35100 34842 35156 34844
rect 35180 34842 35236 34844
rect 34940 34790 34966 34842
rect 34966 34790 34996 34842
rect 35020 34790 35030 34842
rect 35030 34790 35076 34842
rect 35100 34790 35146 34842
rect 35146 34790 35156 34842
rect 35180 34790 35210 34842
rect 35210 34790 35236 34842
rect 34940 34788 34996 34790
rect 35020 34788 35076 34790
rect 35100 34788 35156 34790
rect 35180 34788 35236 34790
rect 32126 19352 32182 19408
rect 32310 18300 32312 18320
rect 32312 18300 32364 18320
rect 32364 18300 32366 18320
rect 32310 18264 32366 18300
rect 33138 19080 33194 19136
rect 33690 18264 33746 18320
rect 31850 9560 31906 9616
rect 31574 8472 31630 8528
rect 29918 3304 29974 3360
rect 34940 33754 34996 33756
rect 35020 33754 35076 33756
rect 35100 33754 35156 33756
rect 35180 33754 35236 33756
rect 34940 33702 34966 33754
rect 34966 33702 34996 33754
rect 35020 33702 35030 33754
rect 35030 33702 35076 33754
rect 35100 33702 35146 33754
rect 35146 33702 35156 33754
rect 35180 33702 35210 33754
rect 35210 33702 35236 33754
rect 34940 33700 34996 33702
rect 35020 33700 35076 33702
rect 35100 33700 35156 33702
rect 35180 33700 35236 33702
rect 34940 32666 34996 32668
rect 35020 32666 35076 32668
rect 35100 32666 35156 32668
rect 35180 32666 35236 32668
rect 34940 32614 34966 32666
rect 34966 32614 34996 32666
rect 35020 32614 35030 32666
rect 35030 32614 35076 32666
rect 35100 32614 35146 32666
rect 35146 32614 35156 32666
rect 35180 32614 35210 32666
rect 35210 32614 35236 32666
rect 34940 32612 34996 32614
rect 35020 32612 35076 32614
rect 35100 32612 35156 32614
rect 35180 32612 35236 32614
rect 34940 31578 34996 31580
rect 35020 31578 35076 31580
rect 35100 31578 35156 31580
rect 35180 31578 35236 31580
rect 34940 31526 34966 31578
rect 34966 31526 34996 31578
rect 35020 31526 35030 31578
rect 35030 31526 35076 31578
rect 35100 31526 35146 31578
rect 35146 31526 35156 31578
rect 35180 31526 35210 31578
rect 35210 31526 35236 31578
rect 34940 31524 34996 31526
rect 35020 31524 35076 31526
rect 35100 31524 35156 31526
rect 35180 31524 35236 31526
rect 35898 35944 35954 36000
rect 34940 30490 34996 30492
rect 35020 30490 35076 30492
rect 35100 30490 35156 30492
rect 35180 30490 35236 30492
rect 34940 30438 34966 30490
rect 34966 30438 34996 30490
rect 35020 30438 35030 30490
rect 35030 30438 35076 30490
rect 35100 30438 35146 30490
rect 35146 30438 35156 30490
rect 35180 30438 35210 30490
rect 35210 30438 35236 30490
rect 34940 30436 34996 30438
rect 35020 30436 35076 30438
rect 35100 30436 35156 30438
rect 35180 30436 35236 30438
rect 34940 29402 34996 29404
rect 35020 29402 35076 29404
rect 35100 29402 35156 29404
rect 35180 29402 35236 29404
rect 34940 29350 34966 29402
rect 34966 29350 34996 29402
rect 35020 29350 35030 29402
rect 35030 29350 35076 29402
rect 35100 29350 35146 29402
rect 35146 29350 35156 29402
rect 35180 29350 35210 29402
rect 35210 29350 35236 29402
rect 34940 29348 34996 29350
rect 35020 29348 35076 29350
rect 35100 29348 35156 29350
rect 35180 29348 35236 29350
rect 34940 28314 34996 28316
rect 35020 28314 35076 28316
rect 35100 28314 35156 28316
rect 35180 28314 35236 28316
rect 34940 28262 34966 28314
rect 34966 28262 34996 28314
rect 35020 28262 35030 28314
rect 35030 28262 35076 28314
rect 35100 28262 35146 28314
rect 35146 28262 35156 28314
rect 35180 28262 35210 28314
rect 35210 28262 35236 28314
rect 34940 28260 34996 28262
rect 35020 28260 35076 28262
rect 35100 28260 35156 28262
rect 35180 28260 35236 28262
rect 34940 27226 34996 27228
rect 35020 27226 35076 27228
rect 35100 27226 35156 27228
rect 35180 27226 35236 27228
rect 34940 27174 34966 27226
rect 34966 27174 34996 27226
rect 35020 27174 35030 27226
rect 35030 27174 35076 27226
rect 35100 27174 35146 27226
rect 35146 27174 35156 27226
rect 35180 27174 35210 27226
rect 35210 27174 35236 27226
rect 34940 27172 34996 27174
rect 35020 27172 35076 27174
rect 35100 27172 35156 27174
rect 35180 27172 35236 27174
rect 34940 26138 34996 26140
rect 35020 26138 35076 26140
rect 35100 26138 35156 26140
rect 35180 26138 35236 26140
rect 34940 26086 34966 26138
rect 34966 26086 34996 26138
rect 35020 26086 35030 26138
rect 35030 26086 35076 26138
rect 35100 26086 35146 26138
rect 35146 26086 35156 26138
rect 35180 26086 35210 26138
rect 35210 26086 35236 26138
rect 34940 26084 34996 26086
rect 35020 26084 35076 26086
rect 35100 26084 35156 26086
rect 35180 26084 35236 26086
rect 34940 25050 34996 25052
rect 35020 25050 35076 25052
rect 35100 25050 35156 25052
rect 35180 25050 35236 25052
rect 34940 24998 34966 25050
rect 34966 24998 34996 25050
rect 35020 24998 35030 25050
rect 35030 24998 35076 25050
rect 35100 24998 35146 25050
rect 35146 24998 35156 25050
rect 35180 24998 35210 25050
rect 35210 24998 35236 25050
rect 34940 24996 34996 24998
rect 35020 24996 35076 24998
rect 35100 24996 35156 24998
rect 35180 24996 35236 24998
rect 34940 23962 34996 23964
rect 35020 23962 35076 23964
rect 35100 23962 35156 23964
rect 35180 23962 35236 23964
rect 34940 23910 34966 23962
rect 34966 23910 34996 23962
rect 35020 23910 35030 23962
rect 35030 23910 35076 23962
rect 35100 23910 35146 23962
rect 35146 23910 35156 23962
rect 35180 23910 35210 23962
rect 35210 23910 35236 23962
rect 34940 23908 34996 23910
rect 35020 23908 35076 23910
rect 35100 23908 35156 23910
rect 35180 23908 35236 23910
rect 34150 18808 34206 18864
rect 34940 22874 34996 22876
rect 35020 22874 35076 22876
rect 35100 22874 35156 22876
rect 35180 22874 35236 22876
rect 34940 22822 34966 22874
rect 34966 22822 34996 22874
rect 35020 22822 35030 22874
rect 35030 22822 35076 22874
rect 35100 22822 35146 22874
rect 35146 22822 35156 22874
rect 35180 22822 35210 22874
rect 35210 22822 35236 22874
rect 34940 22820 34996 22822
rect 35020 22820 35076 22822
rect 35100 22820 35156 22822
rect 35180 22820 35236 22822
rect 34940 21786 34996 21788
rect 35020 21786 35076 21788
rect 35100 21786 35156 21788
rect 35180 21786 35236 21788
rect 34940 21734 34966 21786
rect 34966 21734 34996 21786
rect 35020 21734 35030 21786
rect 35030 21734 35076 21786
rect 35100 21734 35146 21786
rect 35146 21734 35156 21786
rect 35180 21734 35210 21786
rect 35210 21734 35236 21786
rect 34940 21732 34996 21734
rect 35020 21732 35076 21734
rect 35100 21732 35156 21734
rect 35180 21732 35236 21734
rect 34940 20698 34996 20700
rect 35020 20698 35076 20700
rect 35100 20698 35156 20700
rect 35180 20698 35236 20700
rect 34940 20646 34966 20698
rect 34966 20646 34996 20698
rect 35020 20646 35030 20698
rect 35030 20646 35076 20698
rect 35100 20646 35146 20698
rect 35146 20646 35156 20698
rect 35180 20646 35210 20698
rect 35210 20646 35236 20698
rect 34940 20644 34996 20646
rect 35020 20644 35076 20646
rect 35100 20644 35156 20646
rect 35180 20644 35236 20646
rect 34940 19610 34996 19612
rect 35020 19610 35076 19612
rect 35100 19610 35156 19612
rect 35180 19610 35236 19612
rect 34940 19558 34966 19610
rect 34966 19558 34996 19610
rect 35020 19558 35030 19610
rect 35030 19558 35076 19610
rect 35100 19558 35146 19610
rect 35146 19558 35156 19610
rect 35180 19558 35210 19610
rect 35210 19558 35236 19610
rect 34940 19556 34996 19558
rect 35020 19556 35076 19558
rect 35100 19556 35156 19558
rect 35180 19556 35236 19558
rect 34940 18522 34996 18524
rect 35020 18522 35076 18524
rect 35100 18522 35156 18524
rect 35180 18522 35236 18524
rect 34940 18470 34966 18522
rect 34966 18470 34996 18522
rect 35020 18470 35030 18522
rect 35030 18470 35076 18522
rect 35100 18470 35146 18522
rect 35146 18470 35156 18522
rect 35180 18470 35210 18522
rect 35210 18470 35236 18522
rect 34940 18468 34996 18470
rect 35020 18468 35076 18470
rect 35100 18468 35156 18470
rect 35180 18468 35236 18470
rect 34940 17434 34996 17436
rect 35020 17434 35076 17436
rect 35100 17434 35156 17436
rect 35180 17434 35236 17436
rect 34940 17382 34966 17434
rect 34966 17382 34996 17434
rect 35020 17382 35030 17434
rect 35030 17382 35076 17434
rect 35100 17382 35146 17434
rect 35146 17382 35156 17434
rect 35180 17382 35210 17434
rect 35210 17382 35236 17434
rect 34940 17380 34996 17382
rect 35020 17380 35076 17382
rect 35100 17380 35156 17382
rect 35180 17380 35236 17382
rect 34940 16346 34996 16348
rect 35020 16346 35076 16348
rect 35100 16346 35156 16348
rect 35180 16346 35236 16348
rect 34940 16294 34966 16346
rect 34966 16294 34996 16346
rect 35020 16294 35030 16346
rect 35030 16294 35076 16346
rect 35100 16294 35146 16346
rect 35146 16294 35156 16346
rect 35180 16294 35210 16346
rect 35210 16294 35236 16346
rect 34940 16292 34996 16294
rect 35020 16292 35076 16294
rect 35100 16292 35156 16294
rect 35180 16292 35236 16294
rect 34940 15258 34996 15260
rect 35020 15258 35076 15260
rect 35100 15258 35156 15260
rect 35180 15258 35236 15260
rect 34940 15206 34966 15258
rect 34966 15206 34996 15258
rect 35020 15206 35030 15258
rect 35030 15206 35076 15258
rect 35100 15206 35146 15258
rect 35146 15206 35156 15258
rect 35180 15206 35210 15258
rect 35210 15206 35236 15258
rect 34940 15204 34996 15206
rect 35020 15204 35076 15206
rect 35100 15204 35156 15206
rect 35180 15204 35236 15206
rect 34940 14170 34996 14172
rect 35020 14170 35076 14172
rect 35100 14170 35156 14172
rect 35180 14170 35236 14172
rect 34940 14118 34966 14170
rect 34966 14118 34996 14170
rect 35020 14118 35030 14170
rect 35030 14118 35076 14170
rect 35100 14118 35146 14170
rect 35146 14118 35156 14170
rect 35180 14118 35210 14170
rect 35210 14118 35236 14170
rect 34940 14116 34996 14118
rect 35020 14116 35076 14118
rect 35100 14116 35156 14118
rect 35180 14116 35236 14118
rect 33138 9036 33194 9072
rect 34940 13082 34996 13084
rect 35020 13082 35076 13084
rect 35100 13082 35156 13084
rect 35180 13082 35236 13084
rect 34940 13030 34966 13082
rect 34966 13030 34996 13082
rect 35020 13030 35030 13082
rect 35030 13030 35076 13082
rect 35100 13030 35146 13082
rect 35146 13030 35156 13082
rect 35180 13030 35210 13082
rect 35210 13030 35236 13082
rect 34940 13028 34996 13030
rect 35020 13028 35076 13030
rect 35100 13028 35156 13030
rect 35180 13028 35236 13030
rect 34940 11994 34996 11996
rect 35020 11994 35076 11996
rect 35100 11994 35156 11996
rect 35180 11994 35236 11996
rect 34940 11942 34966 11994
rect 34966 11942 34996 11994
rect 35020 11942 35030 11994
rect 35030 11942 35076 11994
rect 35100 11942 35146 11994
rect 35146 11942 35156 11994
rect 35180 11942 35210 11994
rect 35210 11942 35236 11994
rect 34940 11940 34996 11942
rect 35020 11940 35076 11942
rect 35100 11940 35156 11942
rect 35180 11940 35236 11942
rect 34940 10906 34996 10908
rect 35020 10906 35076 10908
rect 35100 10906 35156 10908
rect 35180 10906 35236 10908
rect 34940 10854 34966 10906
rect 34966 10854 34996 10906
rect 35020 10854 35030 10906
rect 35030 10854 35076 10906
rect 35100 10854 35146 10906
rect 35146 10854 35156 10906
rect 35180 10854 35210 10906
rect 35210 10854 35236 10906
rect 34940 10852 34996 10854
rect 35020 10852 35076 10854
rect 35100 10852 35156 10854
rect 35180 10852 35236 10854
rect 34940 9818 34996 9820
rect 35020 9818 35076 9820
rect 35100 9818 35156 9820
rect 35180 9818 35236 9820
rect 34940 9766 34966 9818
rect 34966 9766 34996 9818
rect 35020 9766 35030 9818
rect 35030 9766 35076 9818
rect 35100 9766 35146 9818
rect 35146 9766 35156 9818
rect 35180 9766 35210 9818
rect 35210 9766 35236 9818
rect 34940 9764 34996 9766
rect 35020 9764 35076 9766
rect 35100 9764 35156 9766
rect 35180 9764 35236 9766
rect 37462 32408 37518 32464
rect 37738 32000 37794 32056
rect 35898 19080 35954 19136
rect 36266 19216 36322 19272
rect 36082 18808 36138 18864
rect 36358 18672 36414 18728
rect 36174 18284 36230 18320
rect 36174 18264 36176 18284
rect 36176 18264 36228 18284
rect 36228 18264 36230 18284
rect 35346 9152 35402 9208
rect 33138 9016 33140 9036
rect 33140 9016 33192 9036
rect 33192 9016 33194 9036
rect 34940 8730 34996 8732
rect 35020 8730 35076 8732
rect 35100 8730 35156 8732
rect 35180 8730 35236 8732
rect 34940 8678 34966 8730
rect 34966 8678 34996 8730
rect 35020 8678 35030 8730
rect 35030 8678 35076 8730
rect 35100 8678 35146 8730
rect 35146 8678 35156 8730
rect 35180 8678 35210 8730
rect 35210 8678 35236 8730
rect 34940 8676 34996 8678
rect 35020 8676 35076 8678
rect 35100 8676 35156 8678
rect 35180 8676 35236 8678
rect 31850 6160 31906 6216
rect 33690 3884 33692 3904
rect 33692 3884 33744 3904
rect 33744 3884 33746 3904
rect 33690 3848 33746 3884
rect 34940 7642 34996 7644
rect 35020 7642 35076 7644
rect 35100 7642 35156 7644
rect 35180 7642 35236 7644
rect 34940 7590 34966 7642
rect 34966 7590 34996 7642
rect 35020 7590 35030 7642
rect 35030 7590 35076 7642
rect 35100 7590 35146 7642
rect 35146 7590 35156 7642
rect 35180 7590 35210 7642
rect 35210 7590 35236 7642
rect 34940 7588 34996 7590
rect 35020 7588 35076 7590
rect 35100 7588 35156 7590
rect 35180 7588 35236 7590
rect 34940 6554 34996 6556
rect 35020 6554 35076 6556
rect 35100 6554 35156 6556
rect 35180 6554 35236 6556
rect 34940 6502 34966 6554
rect 34966 6502 34996 6554
rect 35020 6502 35030 6554
rect 35030 6502 35076 6554
rect 35100 6502 35146 6554
rect 35146 6502 35156 6554
rect 35180 6502 35210 6554
rect 35210 6502 35236 6554
rect 34940 6500 34996 6502
rect 35020 6500 35076 6502
rect 35100 6500 35156 6502
rect 35180 6500 35236 6502
rect 34940 5466 34996 5468
rect 35020 5466 35076 5468
rect 35100 5466 35156 5468
rect 35180 5466 35236 5468
rect 34940 5414 34966 5466
rect 34966 5414 34996 5466
rect 35020 5414 35030 5466
rect 35030 5414 35076 5466
rect 35100 5414 35146 5466
rect 35146 5414 35156 5466
rect 35180 5414 35210 5466
rect 35210 5414 35236 5466
rect 34940 5412 34996 5414
rect 35020 5412 35076 5414
rect 35100 5412 35156 5414
rect 35180 5412 35236 5414
rect 37922 21528 37978 21584
rect 37186 10124 37242 10160
rect 37186 10104 37188 10124
rect 37188 10104 37240 10124
rect 37240 10104 37242 10124
rect 39026 32952 39082 33008
rect 39118 30252 39174 30288
rect 39118 30232 39120 30252
rect 39120 30232 39172 30252
rect 39172 30232 39174 30252
rect 39946 27260 40002 27296
rect 39946 27240 39948 27260
rect 39948 27240 40000 27260
rect 40000 27240 40002 27260
rect 38290 24520 38346 24576
rect 38198 18944 38254 19000
rect 38474 15816 38530 15872
rect 38934 13096 38990 13152
rect 38566 7384 38622 7440
rect 35346 4392 35402 4448
rect 34940 4378 34996 4380
rect 35020 4378 35076 4380
rect 35100 4378 35156 4380
rect 35180 4378 35236 4380
rect 34940 4326 34966 4378
rect 34966 4326 34996 4378
rect 35020 4326 35030 4378
rect 35030 4326 35076 4378
rect 35100 4326 35146 4378
rect 35146 4326 35156 4378
rect 35180 4326 35210 4378
rect 35210 4326 35236 4378
rect 34940 4324 34996 4326
rect 35020 4324 35076 4326
rect 35100 4324 35156 4326
rect 35180 4324 35236 4326
rect 35898 3848 35954 3904
rect 34940 3290 34996 3292
rect 35020 3290 35076 3292
rect 35100 3290 35156 3292
rect 35180 3290 35236 3292
rect 34940 3238 34966 3290
rect 34966 3238 34996 3290
rect 35020 3238 35030 3290
rect 35030 3238 35076 3290
rect 35100 3238 35146 3290
rect 35146 3238 35156 3290
rect 35180 3238 35210 3290
rect 35210 3238 35236 3290
rect 34940 3236 34996 3238
rect 35020 3236 35076 3238
rect 35100 3236 35156 3238
rect 35180 3236 35236 3238
rect 34940 2202 34996 2204
rect 35020 2202 35076 2204
rect 35100 2202 35156 2204
rect 35180 2202 35236 2204
rect 34940 2150 34966 2202
rect 34966 2150 34996 2202
rect 35020 2150 35030 2202
rect 35030 2150 35076 2202
rect 35100 2150 35146 2202
rect 35146 2150 35156 2202
rect 35180 2150 35210 2202
rect 35210 2150 35236 2202
rect 34940 2148 34996 2150
rect 35020 2148 35076 2150
rect 35100 2148 35156 2150
rect 35180 2148 35236 2150
rect 37094 1672 37150 1728
<< metal3 >>
rect 35893 38722 35959 38725
rect 40200 38722 41000 38752
rect 35893 38720 41000 38722
rect 35893 38664 35898 38720
rect 35954 38664 41000 38720
rect 35893 38662 41000 38664
rect 35893 38659 35959 38662
rect 19568 38656 19888 38657
rect 19568 38592 19576 38656
rect 19640 38592 19656 38656
rect 19720 38592 19736 38656
rect 19800 38592 19816 38656
rect 19880 38592 19888 38656
rect 40200 38632 41000 38662
rect 19568 38591 19888 38592
rect 4208 38112 4528 38113
rect 4208 38048 4216 38112
rect 4280 38048 4296 38112
rect 4360 38048 4376 38112
rect 4440 38048 4456 38112
rect 4520 38048 4528 38112
rect 4208 38047 4528 38048
rect 34928 38112 35248 38113
rect 34928 38048 34936 38112
rect 35000 38048 35016 38112
rect 35080 38048 35096 38112
rect 35160 38048 35176 38112
rect 35240 38048 35248 38112
rect 34928 38047 35248 38048
rect 0 37906 800 37936
rect 2773 37906 2839 37909
rect 0 37904 2839 37906
rect 0 37848 2778 37904
rect 2834 37848 2839 37904
rect 0 37846 2839 37848
rect 0 37816 800 37846
rect 2773 37843 2839 37846
rect 19568 37568 19888 37569
rect 19568 37504 19576 37568
rect 19640 37504 19656 37568
rect 19720 37504 19736 37568
rect 19800 37504 19816 37568
rect 19880 37504 19888 37568
rect 19568 37503 19888 37504
rect 20897 37362 20963 37365
rect 22921 37362 22987 37365
rect 20897 37360 22987 37362
rect 20897 37304 20902 37360
rect 20958 37304 22926 37360
rect 22982 37304 22987 37360
rect 20897 37302 22987 37304
rect 20897 37299 20963 37302
rect 22921 37299 22987 37302
rect 4208 37024 4528 37025
rect 4208 36960 4216 37024
rect 4280 36960 4296 37024
rect 4360 36960 4376 37024
rect 4440 36960 4456 37024
rect 4520 36960 4528 37024
rect 4208 36959 4528 36960
rect 34928 37024 35248 37025
rect 34928 36960 34936 37024
rect 35000 36960 35016 37024
rect 35080 36960 35096 37024
rect 35160 36960 35176 37024
rect 35240 36960 35248 37024
rect 34928 36959 35248 36960
rect 10593 36682 10659 36685
rect 16573 36682 16639 36685
rect 10593 36680 16639 36682
rect 10593 36624 10598 36680
rect 10654 36624 16578 36680
rect 16634 36624 16639 36680
rect 10593 36622 16639 36624
rect 10593 36619 10659 36622
rect 16573 36619 16639 36622
rect 19793 36682 19859 36685
rect 21725 36682 21791 36685
rect 19793 36680 21791 36682
rect 19793 36624 19798 36680
rect 19854 36624 21730 36680
rect 21786 36624 21791 36680
rect 19793 36622 21791 36624
rect 19793 36619 19859 36622
rect 21725 36619 21791 36622
rect 19568 36480 19888 36481
rect 19568 36416 19576 36480
rect 19640 36416 19656 36480
rect 19720 36416 19736 36480
rect 19800 36416 19816 36480
rect 19880 36416 19888 36480
rect 19568 36415 19888 36416
rect 35893 36002 35959 36005
rect 40200 36002 41000 36032
rect 35893 36000 41000 36002
rect 35893 35944 35898 36000
rect 35954 35944 41000 36000
rect 35893 35942 41000 35944
rect 35893 35939 35959 35942
rect 4208 35936 4528 35937
rect 4208 35872 4216 35936
rect 4280 35872 4296 35936
rect 4360 35872 4376 35936
rect 4440 35872 4456 35936
rect 4520 35872 4528 35936
rect 4208 35871 4528 35872
rect 34928 35936 35248 35937
rect 34928 35872 34936 35936
rect 35000 35872 35016 35936
rect 35080 35872 35096 35936
rect 35160 35872 35176 35936
rect 35240 35872 35248 35936
rect 40200 35912 41000 35942
rect 34928 35871 35248 35872
rect 19568 35392 19888 35393
rect 19568 35328 19576 35392
rect 19640 35328 19656 35392
rect 19720 35328 19736 35392
rect 19800 35328 19816 35392
rect 19880 35328 19888 35392
rect 19568 35327 19888 35328
rect 0 34914 800 34944
rect 4061 34914 4127 34917
rect 0 34912 4127 34914
rect 0 34856 4066 34912
rect 4122 34856 4127 34912
rect 0 34854 4127 34856
rect 0 34824 800 34854
rect 4061 34851 4127 34854
rect 4208 34848 4528 34849
rect 4208 34784 4216 34848
rect 4280 34784 4296 34848
rect 4360 34784 4376 34848
rect 4440 34784 4456 34848
rect 4520 34784 4528 34848
rect 4208 34783 4528 34784
rect 34928 34848 35248 34849
rect 34928 34784 34936 34848
rect 35000 34784 35016 34848
rect 35080 34784 35096 34848
rect 35160 34784 35176 34848
rect 35240 34784 35248 34848
rect 34928 34783 35248 34784
rect 19568 34304 19888 34305
rect 19568 34240 19576 34304
rect 19640 34240 19656 34304
rect 19720 34240 19736 34304
rect 19800 34240 19816 34304
rect 19880 34240 19888 34304
rect 19568 34239 19888 34240
rect 4208 33760 4528 33761
rect 4208 33696 4216 33760
rect 4280 33696 4296 33760
rect 4360 33696 4376 33760
rect 4440 33696 4456 33760
rect 4520 33696 4528 33760
rect 4208 33695 4528 33696
rect 34928 33760 35248 33761
rect 34928 33696 34936 33760
rect 35000 33696 35016 33760
rect 35080 33696 35096 33760
rect 35160 33696 35176 33760
rect 35240 33696 35248 33760
rect 34928 33695 35248 33696
rect 19568 33216 19888 33217
rect 19568 33152 19576 33216
rect 19640 33152 19656 33216
rect 19720 33152 19736 33216
rect 19800 33152 19816 33216
rect 19880 33152 19888 33216
rect 19568 33151 19888 33152
rect 39021 33010 39087 33013
rect 40200 33010 41000 33040
rect 39021 33008 41000 33010
rect 39021 32952 39026 33008
rect 39082 32952 41000 33008
rect 39021 32950 41000 32952
rect 39021 32947 39087 32950
rect 40200 32920 41000 32950
rect 4208 32672 4528 32673
rect 4208 32608 4216 32672
rect 4280 32608 4296 32672
rect 4360 32608 4376 32672
rect 4440 32608 4456 32672
rect 4520 32608 4528 32672
rect 4208 32607 4528 32608
rect 34928 32672 35248 32673
rect 34928 32608 34936 32672
rect 35000 32608 35016 32672
rect 35080 32608 35096 32672
rect 35160 32608 35176 32672
rect 35240 32608 35248 32672
rect 34928 32607 35248 32608
rect 29177 32466 29243 32469
rect 37457 32466 37523 32469
rect 29177 32464 37523 32466
rect 29177 32408 29182 32464
rect 29238 32408 37462 32464
rect 37518 32408 37523 32464
rect 29177 32406 37523 32408
rect 29177 32403 29243 32406
rect 37457 32403 37523 32406
rect 0 32194 800 32224
rect 2957 32194 3023 32197
rect 0 32192 3023 32194
rect 0 32136 2962 32192
rect 3018 32136 3023 32192
rect 0 32134 3023 32136
rect 0 32104 800 32134
rect 2957 32131 3023 32134
rect 18413 32194 18479 32197
rect 19149 32194 19215 32197
rect 18413 32192 19215 32194
rect 18413 32136 18418 32192
rect 18474 32136 19154 32192
rect 19210 32136 19215 32192
rect 18413 32134 19215 32136
rect 18413 32131 18479 32134
rect 19149 32131 19215 32134
rect 19568 32128 19888 32129
rect 19568 32064 19576 32128
rect 19640 32064 19656 32128
rect 19720 32064 19736 32128
rect 19800 32064 19816 32128
rect 19880 32064 19888 32128
rect 19568 32063 19888 32064
rect 37733 32060 37799 32061
rect 37733 32056 37780 32060
rect 37844 32058 37850 32060
rect 37733 32000 37738 32056
rect 37733 31996 37780 32000
rect 37844 31998 37890 32058
rect 37844 31996 37850 31998
rect 37733 31995 37799 31996
rect 19333 31922 19399 31925
rect 20345 31922 20411 31925
rect 19333 31920 20411 31922
rect 19333 31864 19338 31920
rect 19394 31864 20350 31920
rect 20406 31864 20411 31920
rect 19333 31862 20411 31864
rect 19333 31859 19399 31862
rect 20345 31859 20411 31862
rect 23289 31786 23355 31789
rect 25497 31786 25563 31789
rect 23289 31784 25563 31786
rect 23289 31728 23294 31784
rect 23350 31728 25502 31784
rect 25558 31728 25563 31784
rect 23289 31726 25563 31728
rect 23289 31723 23355 31726
rect 25497 31723 25563 31726
rect 4208 31584 4528 31585
rect 4208 31520 4216 31584
rect 4280 31520 4296 31584
rect 4360 31520 4376 31584
rect 4440 31520 4456 31584
rect 4520 31520 4528 31584
rect 4208 31519 4528 31520
rect 34928 31584 35248 31585
rect 34928 31520 34936 31584
rect 35000 31520 35016 31584
rect 35080 31520 35096 31584
rect 35160 31520 35176 31584
rect 35240 31520 35248 31584
rect 34928 31519 35248 31520
rect 19568 31040 19888 31041
rect 19568 30976 19576 31040
rect 19640 30976 19656 31040
rect 19720 30976 19736 31040
rect 19800 30976 19816 31040
rect 19880 30976 19888 31040
rect 19568 30975 19888 30976
rect 13 30834 79 30837
rect 25221 30834 25287 30837
rect 13 30832 25287 30834
rect 13 30776 18 30832
rect 74 30776 25226 30832
rect 25282 30776 25287 30832
rect 13 30774 25287 30776
rect 13 30771 79 30774
rect 25221 30771 25287 30774
rect 27061 30700 27127 30701
rect 27061 30698 27108 30700
rect 27016 30696 27108 30698
rect 27016 30640 27066 30696
rect 27016 30638 27108 30640
rect 27061 30636 27108 30638
rect 27172 30636 27178 30700
rect 27061 30635 27127 30636
rect 4208 30496 4528 30497
rect 4208 30432 4216 30496
rect 4280 30432 4296 30496
rect 4360 30432 4376 30496
rect 4440 30432 4456 30496
rect 4520 30432 4528 30496
rect 4208 30431 4528 30432
rect 34928 30496 35248 30497
rect 34928 30432 34936 30496
rect 35000 30432 35016 30496
rect 35080 30432 35096 30496
rect 35160 30432 35176 30496
rect 35240 30432 35248 30496
rect 34928 30431 35248 30432
rect 39113 30290 39179 30293
rect 40200 30290 41000 30320
rect 39113 30288 41000 30290
rect 39113 30232 39118 30288
rect 39174 30232 41000 30288
rect 39113 30230 41000 30232
rect 39113 30227 39179 30230
rect 40200 30200 41000 30230
rect 19793 30154 19859 30157
rect 20713 30154 20779 30157
rect 19793 30152 20779 30154
rect 19793 30096 19798 30152
rect 19854 30096 20718 30152
rect 20774 30096 20779 30152
rect 19793 30094 20779 30096
rect 19793 30091 19859 30094
rect 20713 30091 20779 30094
rect 19568 29952 19888 29953
rect 19568 29888 19576 29952
rect 19640 29888 19656 29952
rect 19720 29888 19736 29952
rect 19800 29888 19816 29952
rect 19880 29888 19888 29952
rect 19568 29887 19888 29888
rect 10501 29746 10567 29749
rect 12617 29746 12683 29749
rect 10501 29744 12683 29746
rect 10501 29688 10506 29744
rect 10562 29688 12622 29744
rect 12678 29688 12683 29744
rect 10501 29686 12683 29688
rect 10501 29683 10567 29686
rect 12617 29683 12683 29686
rect 10041 29610 10107 29613
rect 10685 29610 10751 29613
rect 12893 29610 12959 29613
rect 10041 29608 12959 29610
rect 10041 29552 10046 29608
rect 10102 29552 10690 29608
rect 10746 29552 12898 29608
rect 12954 29552 12959 29608
rect 10041 29550 12959 29552
rect 10041 29547 10107 29550
rect 10685 29547 10751 29550
rect 12893 29547 12959 29550
rect 19609 29610 19675 29613
rect 19977 29610 20043 29613
rect 19609 29608 20043 29610
rect 19609 29552 19614 29608
rect 19670 29552 19982 29608
rect 20038 29552 20043 29608
rect 19609 29550 20043 29552
rect 19609 29547 19675 29550
rect 19977 29547 20043 29550
rect 22921 29610 22987 29613
rect 24209 29610 24275 29613
rect 22921 29608 24275 29610
rect 22921 29552 22926 29608
rect 22982 29552 24214 29608
rect 24270 29552 24275 29608
rect 22921 29550 24275 29552
rect 22921 29547 22987 29550
rect 24209 29547 24275 29550
rect 4208 29408 4528 29409
rect 4208 29344 4216 29408
rect 4280 29344 4296 29408
rect 4360 29344 4376 29408
rect 4440 29344 4456 29408
rect 4520 29344 4528 29408
rect 4208 29343 4528 29344
rect 34928 29408 35248 29409
rect 34928 29344 34936 29408
rect 35000 29344 35016 29408
rect 35080 29344 35096 29408
rect 35160 29344 35176 29408
rect 35240 29344 35248 29408
rect 34928 29343 35248 29344
rect 19793 29338 19859 29341
rect 20161 29338 20227 29341
rect 19793 29336 20227 29338
rect 19793 29280 19798 29336
rect 19854 29280 20166 29336
rect 20222 29280 20227 29336
rect 19793 29278 20227 29280
rect 19793 29275 19859 29278
rect 20161 29275 20227 29278
rect 23289 29338 23355 29341
rect 24669 29338 24735 29341
rect 23289 29336 24735 29338
rect 23289 29280 23294 29336
rect 23350 29280 24674 29336
rect 24730 29280 24735 29336
rect 23289 29278 24735 29280
rect 23289 29275 23355 29278
rect 24669 29275 24735 29278
rect 0 29202 800 29232
rect 9397 29202 9463 29205
rect 0 29200 9463 29202
rect 0 29144 9402 29200
rect 9458 29144 9463 29200
rect 0 29142 9463 29144
rect 0 29112 800 29142
rect 9397 29139 9463 29142
rect 18781 29202 18847 29205
rect 21817 29202 21883 29205
rect 18781 29200 21883 29202
rect 18781 29144 18786 29200
rect 18842 29144 21822 29200
rect 21878 29144 21883 29200
rect 18781 29142 21883 29144
rect 18781 29139 18847 29142
rect 21817 29139 21883 29142
rect 3969 29066 4035 29069
rect 3742 29064 4035 29066
rect 3742 29008 3974 29064
rect 4030 29008 4035 29064
rect 3742 29006 4035 29008
rect 3509 28794 3575 28797
rect 3742 28794 3802 29006
rect 3969 29003 4035 29006
rect 23933 29066 23999 29069
rect 27613 29066 27679 29069
rect 23933 29064 27679 29066
rect 23933 29008 23938 29064
rect 23994 29008 27618 29064
rect 27674 29008 27679 29064
rect 23933 29006 27679 29008
rect 23933 29003 23999 29006
rect 27613 29003 27679 29006
rect 19425 28932 19491 28933
rect 19374 28930 19380 28932
rect 19334 28870 19380 28930
rect 19444 28928 19491 28932
rect 19486 28872 19491 28928
rect 19374 28868 19380 28870
rect 19444 28868 19491 28872
rect 19425 28867 19491 28868
rect 19568 28864 19888 28865
rect 19568 28800 19576 28864
rect 19640 28800 19656 28864
rect 19720 28800 19736 28864
rect 19800 28800 19816 28864
rect 19880 28800 19888 28864
rect 19568 28799 19888 28800
rect 3509 28792 3802 28794
rect 3509 28736 3514 28792
rect 3570 28736 3802 28792
rect 3509 28734 3802 28736
rect 3509 28731 3575 28734
rect 19333 28522 19399 28525
rect 27521 28522 27587 28525
rect 19333 28520 27587 28522
rect 19333 28464 19338 28520
rect 19394 28464 27526 28520
rect 27582 28464 27587 28520
rect 19333 28462 27587 28464
rect 19333 28459 19399 28462
rect 27521 28459 27587 28462
rect 4208 28320 4528 28321
rect 4208 28256 4216 28320
rect 4280 28256 4296 28320
rect 4360 28256 4376 28320
rect 4440 28256 4456 28320
rect 4520 28256 4528 28320
rect 4208 28255 4528 28256
rect 34928 28320 35248 28321
rect 34928 28256 34936 28320
rect 35000 28256 35016 28320
rect 35080 28256 35096 28320
rect 35160 28256 35176 28320
rect 35240 28256 35248 28320
rect 34928 28255 35248 28256
rect 21541 28114 21607 28117
rect 27797 28114 27863 28117
rect 21541 28112 27863 28114
rect 21541 28056 21546 28112
rect 21602 28056 27802 28112
rect 27858 28056 27863 28112
rect 21541 28054 27863 28056
rect 21541 28051 21607 28054
rect 27797 28051 27863 28054
rect 19568 27776 19888 27777
rect 19568 27712 19576 27776
rect 19640 27712 19656 27776
rect 19720 27712 19736 27776
rect 19800 27712 19816 27776
rect 19880 27712 19888 27776
rect 19568 27711 19888 27712
rect 39941 27298 40007 27301
rect 40200 27298 41000 27328
rect 39941 27296 41000 27298
rect 39941 27240 39946 27296
rect 40002 27240 41000 27296
rect 39941 27238 41000 27240
rect 39941 27235 40007 27238
rect 4208 27232 4528 27233
rect 4208 27168 4216 27232
rect 4280 27168 4296 27232
rect 4360 27168 4376 27232
rect 4440 27168 4456 27232
rect 4520 27168 4528 27232
rect 4208 27167 4528 27168
rect 34928 27232 35248 27233
rect 34928 27168 34936 27232
rect 35000 27168 35016 27232
rect 35080 27168 35096 27232
rect 35160 27168 35176 27232
rect 35240 27168 35248 27232
rect 40200 27208 41000 27238
rect 34928 27167 35248 27168
rect 19568 26688 19888 26689
rect 19568 26624 19576 26688
rect 19640 26624 19656 26688
rect 19720 26624 19736 26688
rect 19800 26624 19816 26688
rect 19880 26624 19888 26688
rect 19568 26623 19888 26624
rect 0 26482 800 26512
rect 2865 26482 2931 26485
rect 0 26480 2931 26482
rect 0 26424 2870 26480
rect 2926 26424 2931 26480
rect 0 26422 2931 26424
rect 0 26392 800 26422
rect 2865 26419 2931 26422
rect 4208 26144 4528 26145
rect 4208 26080 4216 26144
rect 4280 26080 4296 26144
rect 4360 26080 4376 26144
rect 4440 26080 4456 26144
rect 4520 26080 4528 26144
rect 4208 26079 4528 26080
rect 34928 26144 35248 26145
rect 34928 26080 34936 26144
rect 35000 26080 35016 26144
rect 35080 26080 35096 26144
rect 35160 26080 35176 26144
rect 35240 26080 35248 26144
rect 34928 26079 35248 26080
rect 2313 25802 2379 25805
rect 6177 25802 6243 25805
rect 2313 25800 6243 25802
rect 2313 25744 2318 25800
rect 2374 25744 6182 25800
rect 6238 25744 6243 25800
rect 2313 25742 6243 25744
rect 2313 25739 2379 25742
rect 6177 25739 6243 25742
rect 19568 25600 19888 25601
rect 19568 25536 19576 25600
rect 19640 25536 19656 25600
rect 19720 25536 19736 25600
rect 19800 25536 19816 25600
rect 19880 25536 19888 25600
rect 19568 25535 19888 25536
rect 4208 25056 4528 25057
rect 4208 24992 4216 25056
rect 4280 24992 4296 25056
rect 4360 24992 4376 25056
rect 4440 24992 4456 25056
rect 4520 24992 4528 25056
rect 4208 24991 4528 24992
rect 34928 25056 35248 25057
rect 34928 24992 34936 25056
rect 35000 24992 35016 25056
rect 35080 24992 35096 25056
rect 35160 24992 35176 25056
rect 35240 24992 35248 25056
rect 34928 24991 35248 24992
rect 38285 24578 38351 24581
rect 40200 24578 41000 24608
rect 38285 24576 41000 24578
rect 38285 24520 38290 24576
rect 38346 24520 41000 24576
rect 38285 24518 41000 24520
rect 38285 24515 38351 24518
rect 19568 24512 19888 24513
rect 19568 24448 19576 24512
rect 19640 24448 19656 24512
rect 19720 24448 19736 24512
rect 19800 24448 19816 24512
rect 19880 24448 19888 24512
rect 40200 24488 41000 24518
rect 19568 24447 19888 24448
rect 4208 23968 4528 23969
rect 4208 23904 4216 23968
rect 4280 23904 4296 23968
rect 4360 23904 4376 23968
rect 4440 23904 4456 23968
rect 4520 23904 4528 23968
rect 4208 23903 4528 23904
rect 34928 23968 35248 23969
rect 34928 23904 34936 23968
rect 35000 23904 35016 23968
rect 35080 23904 35096 23968
rect 35160 23904 35176 23968
rect 35240 23904 35248 23968
rect 34928 23903 35248 23904
rect 0 23490 800 23520
rect 2773 23490 2839 23493
rect 0 23488 2839 23490
rect 0 23432 2778 23488
rect 2834 23432 2839 23488
rect 0 23430 2839 23432
rect 0 23400 800 23430
rect 2773 23427 2839 23430
rect 19568 23424 19888 23425
rect 19568 23360 19576 23424
rect 19640 23360 19656 23424
rect 19720 23360 19736 23424
rect 19800 23360 19816 23424
rect 19880 23360 19888 23424
rect 19568 23359 19888 23360
rect 19425 23356 19491 23357
rect 19374 23354 19380 23356
rect 19334 23294 19380 23354
rect 19444 23352 19491 23356
rect 19486 23296 19491 23352
rect 19374 23292 19380 23294
rect 19444 23292 19491 23296
rect 19425 23291 19491 23292
rect 4208 22880 4528 22881
rect 4208 22816 4216 22880
rect 4280 22816 4296 22880
rect 4360 22816 4376 22880
rect 4440 22816 4456 22880
rect 4520 22816 4528 22880
rect 4208 22815 4528 22816
rect 34928 22880 35248 22881
rect 34928 22816 34936 22880
rect 35000 22816 35016 22880
rect 35080 22816 35096 22880
rect 35160 22816 35176 22880
rect 35240 22816 35248 22880
rect 34928 22815 35248 22816
rect 26417 22538 26483 22541
rect 26877 22538 26943 22541
rect 28533 22538 28599 22541
rect 26417 22536 28599 22538
rect 26417 22480 26422 22536
rect 26478 22480 26882 22536
rect 26938 22480 28538 22536
rect 28594 22480 28599 22536
rect 26417 22478 28599 22480
rect 26417 22475 26483 22478
rect 26877 22475 26943 22478
rect 28533 22475 28599 22478
rect 19568 22336 19888 22337
rect 19568 22272 19576 22336
rect 19640 22272 19656 22336
rect 19720 22272 19736 22336
rect 19800 22272 19816 22336
rect 19880 22272 19888 22336
rect 19568 22271 19888 22272
rect 4208 21792 4528 21793
rect 4208 21728 4216 21792
rect 4280 21728 4296 21792
rect 4360 21728 4376 21792
rect 4440 21728 4456 21792
rect 4520 21728 4528 21792
rect 4208 21727 4528 21728
rect 34928 21792 35248 21793
rect 34928 21728 34936 21792
rect 35000 21728 35016 21792
rect 35080 21728 35096 21792
rect 35160 21728 35176 21792
rect 35240 21728 35248 21792
rect 34928 21727 35248 21728
rect 37917 21586 37983 21589
rect 40200 21586 41000 21616
rect 37917 21584 41000 21586
rect 37917 21528 37922 21584
rect 37978 21528 41000 21584
rect 37917 21526 41000 21528
rect 37917 21523 37983 21526
rect 40200 21496 41000 21526
rect 19568 21248 19888 21249
rect 19568 21184 19576 21248
rect 19640 21184 19656 21248
rect 19720 21184 19736 21248
rect 19800 21184 19816 21248
rect 19880 21184 19888 21248
rect 19568 21183 19888 21184
rect 0 20770 800 20800
rect 3417 20770 3483 20773
rect 0 20768 3483 20770
rect 0 20712 3422 20768
rect 3478 20712 3483 20768
rect 0 20710 3483 20712
rect 0 20680 800 20710
rect 3417 20707 3483 20710
rect 4208 20704 4528 20705
rect 4208 20640 4216 20704
rect 4280 20640 4296 20704
rect 4360 20640 4376 20704
rect 4440 20640 4456 20704
rect 4520 20640 4528 20704
rect 4208 20639 4528 20640
rect 34928 20704 35248 20705
rect 34928 20640 34936 20704
rect 35000 20640 35016 20704
rect 35080 20640 35096 20704
rect 35160 20640 35176 20704
rect 35240 20640 35248 20704
rect 34928 20639 35248 20640
rect 16297 20362 16363 20365
rect 37774 20362 37780 20364
rect 16297 20360 37780 20362
rect 16297 20304 16302 20360
rect 16358 20304 37780 20360
rect 16297 20302 37780 20304
rect 16297 20299 16363 20302
rect 37774 20300 37780 20302
rect 37844 20300 37850 20364
rect 19568 20160 19888 20161
rect 19568 20096 19576 20160
rect 19640 20096 19656 20160
rect 19720 20096 19736 20160
rect 19800 20096 19816 20160
rect 19880 20096 19888 20160
rect 19568 20095 19888 20096
rect 19425 19956 19491 19957
rect 19374 19954 19380 19956
rect 19334 19894 19380 19954
rect 19444 19952 19491 19956
rect 19486 19896 19491 19952
rect 19374 19892 19380 19894
rect 19444 19892 19491 19896
rect 19425 19891 19491 19892
rect 19701 19954 19767 19957
rect 23013 19954 23079 19957
rect 19701 19952 23079 19954
rect 19701 19896 19706 19952
rect 19762 19896 23018 19952
rect 23074 19896 23079 19952
rect 19701 19894 23079 19896
rect 19701 19891 19767 19894
rect 23013 19891 23079 19894
rect 4208 19616 4528 19617
rect 4208 19552 4216 19616
rect 4280 19552 4296 19616
rect 4360 19552 4376 19616
rect 4440 19552 4456 19616
rect 4520 19552 4528 19616
rect 4208 19551 4528 19552
rect 34928 19616 35248 19617
rect 34928 19552 34936 19616
rect 35000 19552 35016 19616
rect 35080 19552 35096 19616
rect 35160 19552 35176 19616
rect 35240 19552 35248 19616
rect 34928 19551 35248 19552
rect 19977 19546 20043 19549
rect 20161 19546 20227 19549
rect 19977 19544 20227 19546
rect 19977 19488 19982 19544
rect 20038 19488 20166 19544
rect 20222 19488 20227 19544
rect 19977 19486 20227 19488
rect 19977 19483 20043 19486
rect 20161 19483 20227 19486
rect 29085 19546 29151 19549
rect 30281 19546 30347 19549
rect 29085 19544 30347 19546
rect 29085 19488 29090 19544
rect 29146 19488 30286 19544
rect 30342 19488 30347 19544
rect 29085 19486 30347 19488
rect 29085 19483 29151 19486
rect 30281 19483 30347 19486
rect 21398 19348 21404 19412
rect 21468 19410 21474 19412
rect 21633 19410 21699 19413
rect 21468 19408 21699 19410
rect 21468 19352 21638 19408
rect 21694 19352 21699 19408
rect 21468 19350 21699 19352
rect 21468 19348 21474 19350
rect 21633 19347 21699 19350
rect 31569 19410 31635 19413
rect 32121 19410 32187 19413
rect 31569 19408 32187 19410
rect 31569 19352 31574 19408
rect 31630 19352 32126 19408
rect 32182 19352 32187 19408
rect 31569 19350 32187 19352
rect 31569 19347 31635 19350
rect 32121 19347 32187 19350
rect 28809 19276 28875 19277
rect 28758 19274 28764 19276
rect 28718 19214 28764 19274
rect 28828 19272 28875 19276
rect 28870 19216 28875 19272
rect 28758 19212 28764 19214
rect 28828 19212 28875 19216
rect 28809 19211 28875 19212
rect 31385 19274 31451 19277
rect 36261 19274 36327 19277
rect 31385 19272 36327 19274
rect 31385 19216 31390 19272
rect 31446 19216 36266 19272
rect 36322 19216 36327 19272
rect 31385 19214 36327 19216
rect 31385 19211 31451 19214
rect 36261 19211 36327 19214
rect 27613 19138 27679 19141
rect 28901 19138 28967 19141
rect 27613 19136 28967 19138
rect 27613 19080 27618 19136
rect 27674 19080 28906 19136
rect 28962 19080 28967 19136
rect 27613 19078 28967 19080
rect 27613 19075 27679 19078
rect 28901 19075 28967 19078
rect 29637 19138 29703 19141
rect 30833 19138 30899 19141
rect 33133 19138 33199 19141
rect 35893 19138 35959 19141
rect 29637 19136 35959 19138
rect 29637 19080 29642 19136
rect 29698 19080 30838 19136
rect 30894 19080 33138 19136
rect 33194 19080 35898 19136
rect 35954 19080 35959 19136
rect 29637 19078 35959 19080
rect 29637 19075 29703 19078
rect 30833 19075 30899 19078
rect 33133 19075 33199 19078
rect 35893 19075 35959 19078
rect 19568 19072 19888 19073
rect 19568 19008 19576 19072
rect 19640 19008 19656 19072
rect 19720 19008 19736 19072
rect 19800 19008 19816 19072
rect 19880 19008 19888 19072
rect 19568 19007 19888 19008
rect 25497 19002 25563 19005
rect 29729 19002 29795 19005
rect 38193 19002 38259 19005
rect 25497 19000 38259 19002
rect 25497 18944 25502 19000
rect 25558 18944 29734 19000
rect 29790 18944 38198 19000
rect 38254 18944 38259 19000
rect 25497 18942 38259 18944
rect 25497 18939 25563 18942
rect 29729 18939 29795 18942
rect 38193 18939 38259 18942
rect 19517 18866 19583 18869
rect 20529 18866 20595 18869
rect 19517 18864 20595 18866
rect 19517 18808 19522 18864
rect 19578 18808 20534 18864
rect 20590 18808 20595 18864
rect 19517 18806 20595 18808
rect 19517 18803 19583 18806
rect 20529 18803 20595 18806
rect 28257 18866 28323 18869
rect 28717 18866 28783 18869
rect 28257 18864 28783 18866
rect 28257 18808 28262 18864
rect 28318 18808 28722 18864
rect 28778 18808 28783 18864
rect 28257 18806 28783 18808
rect 28257 18803 28323 18806
rect 28717 18803 28783 18806
rect 31661 18866 31727 18869
rect 34145 18866 34211 18869
rect 31661 18864 34211 18866
rect 31661 18808 31666 18864
rect 31722 18808 34150 18864
rect 34206 18808 34211 18864
rect 31661 18806 34211 18808
rect 31661 18803 31727 18806
rect 34145 18803 34211 18806
rect 36077 18866 36143 18869
rect 40200 18866 41000 18896
rect 36077 18864 41000 18866
rect 36077 18808 36082 18864
rect 36138 18808 41000 18864
rect 36077 18806 41000 18808
rect 36077 18803 36143 18806
rect 40200 18776 41000 18806
rect 1945 18730 2011 18733
rect 9489 18730 9555 18733
rect 1945 18728 9555 18730
rect 1945 18672 1950 18728
rect 2006 18672 9494 18728
rect 9550 18672 9555 18728
rect 1945 18670 9555 18672
rect 1945 18667 2011 18670
rect 9489 18667 9555 18670
rect 19609 18730 19675 18733
rect 22093 18730 22159 18733
rect 19609 18728 22159 18730
rect 19609 18672 19614 18728
rect 19670 18672 22098 18728
rect 22154 18672 22159 18728
rect 19609 18670 22159 18672
rect 19609 18667 19675 18670
rect 22093 18667 22159 18670
rect 27153 18730 27219 18733
rect 28901 18730 28967 18733
rect 27153 18728 28967 18730
rect 27153 18672 27158 18728
rect 27214 18672 28906 18728
rect 28962 18672 28967 18728
rect 27153 18670 28967 18672
rect 27153 18667 27219 18670
rect 28901 18667 28967 18670
rect 30373 18730 30439 18733
rect 36353 18730 36419 18733
rect 30373 18728 36419 18730
rect 30373 18672 30378 18728
rect 30434 18672 36358 18728
rect 36414 18672 36419 18728
rect 30373 18670 36419 18672
rect 30373 18667 30439 18670
rect 36353 18667 36419 18670
rect 25313 18594 25379 18597
rect 27429 18594 27495 18597
rect 25313 18592 27495 18594
rect 25313 18536 25318 18592
rect 25374 18536 27434 18592
rect 27490 18536 27495 18592
rect 25313 18534 27495 18536
rect 25313 18531 25379 18534
rect 27429 18531 27495 18534
rect 4208 18528 4528 18529
rect 4208 18464 4216 18528
rect 4280 18464 4296 18528
rect 4360 18464 4376 18528
rect 4440 18464 4456 18528
rect 4520 18464 4528 18528
rect 4208 18463 4528 18464
rect 34928 18528 35248 18529
rect 34928 18464 34936 18528
rect 35000 18464 35016 18528
rect 35080 18464 35096 18528
rect 35160 18464 35176 18528
rect 35240 18464 35248 18528
rect 34928 18463 35248 18464
rect 28533 18458 28599 18461
rect 30005 18458 30071 18461
rect 28533 18456 30071 18458
rect 28533 18400 28538 18456
rect 28594 18400 30010 18456
rect 30066 18400 30071 18456
rect 28533 18398 30071 18400
rect 28533 18395 28599 18398
rect 30005 18395 30071 18398
rect 32305 18322 32371 18325
rect 33685 18322 33751 18325
rect 36169 18322 36235 18325
rect 32305 18320 36235 18322
rect 32305 18264 32310 18320
rect 32366 18264 33690 18320
rect 33746 18264 36174 18320
rect 36230 18264 36235 18320
rect 32305 18262 36235 18264
rect 32305 18259 32371 18262
rect 33685 18259 33751 18262
rect 36169 18259 36235 18262
rect 19149 18186 19215 18189
rect 19701 18186 19767 18189
rect 19149 18184 19767 18186
rect 19149 18128 19154 18184
rect 19210 18128 19706 18184
rect 19762 18128 19767 18184
rect 19149 18126 19767 18128
rect 19149 18123 19215 18126
rect 19701 18123 19767 18126
rect 19568 17984 19888 17985
rect 19568 17920 19576 17984
rect 19640 17920 19656 17984
rect 19720 17920 19736 17984
rect 19800 17920 19816 17984
rect 19880 17920 19888 17984
rect 19568 17919 19888 17920
rect 0 17778 800 17808
rect 1945 17778 2011 17781
rect 0 17776 2011 17778
rect 0 17720 1950 17776
rect 2006 17720 2011 17776
rect 0 17718 2011 17720
rect 0 17688 800 17718
rect 1945 17715 2011 17718
rect 4208 17440 4528 17441
rect 4208 17376 4216 17440
rect 4280 17376 4296 17440
rect 4360 17376 4376 17440
rect 4440 17376 4456 17440
rect 4520 17376 4528 17440
rect 4208 17375 4528 17376
rect 34928 17440 35248 17441
rect 34928 17376 34936 17440
rect 35000 17376 35016 17440
rect 35080 17376 35096 17440
rect 35160 17376 35176 17440
rect 35240 17376 35248 17440
rect 34928 17375 35248 17376
rect 19568 16896 19888 16897
rect 19568 16832 19576 16896
rect 19640 16832 19656 16896
rect 19720 16832 19736 16896
rect 19800 16832 19816 16896
rect 19880 16832 19888 16896
rect 19568 16831 19888 16832
rect 4208 16352 4528 16353
rect 4208 16288 4216 16352
rect 4280 16288 4296 16352
rect 4360 16288 4376 16352
rect 4440 16288 4456 16352
rect 4520 16288 4528 16352
rect 4208 16287 4528 16288
rect 34928 16352 35248 16353
rect 34928 16288 34936 16352
rect 35000 16288 35016 16352
rect 35080 16288 35096 16352
rect 35160 16288 35176 16352
rect 35240 16288 35248 16352
rect 34928 16287 35248 16288
rect 38469 15874 38535 15877
rect 40200 15874 41000 15904
rect 38469 15872 41000 15874
rect 38469 15816 38474 15872
rect 38530 15816 41000 15872
rect 38469 15814 41000 15816
rect 38469 15811 38535 15814
rect 19568 15808 19888 15809
rect 19568 15744 19576 15808
rect 19640 15744 19656 15808
rect 19720 15744 19736 15808
rect 19800 15744 19816 15808
rect 19880 15744 19888 15808
rect 40200 15784 41000 15814
rect 19568 15743 19888 15744
rect 4208 15264 4528 15265
rect 4208 15200 4216 15264
rect 4280 15200 4296 15264
rect 4360 15200 4376 15264
rect 4440 15200 4456 15264
rect 4520 15200 4528 15264
rect 4208 15199 4528 15200
rect 34928 15264 35248 15265
rect 34928 15200 34936 15264
rect 35000 15200 35016 15264
rect 35080 15200 35096 15264
rect 35160 15200 35176 15264
rect 35240 15200 35248 15264
rect 34928 15199 35248 15200
rect 0 15058 800 15088
rect 4061 15058 4127 15061
rect 0 15056 4127 15058
rect 0 15000 4066 15056
rect 4122 15000 4127 15056
rect 0 14998 4127 15000
rect 0 14968 800 14998
rect 4061 14995 4127 14998
rect 19568 14720 19888 14721
rect 19568 14656 19576 14720
rect 19640 14656 19656 14720
rect 19720 14656 19736 14720
rect 19800 14656 19816 14720
rect 19880 14656 19888 14720
rect 19568 14655 19888 14656
rect 3877 14650 3943 14653
rect 9489 14650 9555 14653
rect 3877 14648 9555 14650
rect 3877 14592 3882 14648
rect 3938 14592 9494 14648
rect 9550 14592 9555 14648
rect 3877 14590 9555 14592
rect 3877 14587 3943 14590
rect 9489 14587 9555 14590
rect 1669 14514 1735 14517
rect 5073 14514 5139 14517
rect 1669 14512 5139 14514
rect 1669 14456 1674 14512
rect 1730 14456 5078 14512
rect 5134 14456 5139 14512
rect 1669 14454 5139 14456
rect 1669 14451 1735 14454
rect 5073 14451 5139 14454
rect 28625 14514 28691 14517
rect 28758 14514 28764 14516
rect 28625 14512 28764 14514
rect 28625 14456 28630 14512
rect 28686 14456 28764 14512
rect 28625 14454 28764 14456
rect 28625 14451 28691 14454
rect 28758 14452 28764 14454
rect 28828 14452 28834 14516
rect 4208 14176 4528 14177
rect 4208 14112 4216 14176
rect 4280 14112 4296 14176
rect 4360 14112 4376 14176
rect 4440 14112 4456 14176
rect 4520 14112 4528 14176
rect 4208 14111 4528 14112
rect 34928 14176 35248 14177
rect 34928 14112 34936 14176
rect 35000 14112 35016 14176
rect 35080 14112 35096 14176
rect 35160 14112 35176 14176
rect 35240 14112 35248 14176
rect 34928 14111 35248 14112
rect 19568 13632 19888 13633
rect 19568 13568 19576 13632
rect 19640 13568 19656 13632
rect 19720 13568 19736 13632
rect 19800 13568 19816 13632
rect 19880 13568 19888 13632
rect 19568 13567 19888 13568
rect 38929 13154 38995 13157
rect 40200 13154 41000 13184
rect 38929 13152 41000 13154
rect 38929 13096 38934 13152
rect 38990 13096 41000 13152
rect 38929 13094 41000 13096
rect 38929 13091 38995 13094
rect 4208 13088 4528 13089
rect 4208 13024 4216 13088
rect 4280 13024 4296 13088
rect 4360 13024 4376 13088
rect 4440 13024 4456 13088
rect 4520 13024 4528 13088
rect 4208 13023 4528 13024
rect 34928 13088 35248 13089
rect 34928 13024 34936 13088
rect 35000 13024 35016 13088
rect 35080 13024 35096 13088
rect 35160 13024 35176 13088
rect 35240 13024 35248 13088
rect 40200 13064 41000 13094
rect 34928 13023 35248 13024
rect 19568 12544 19888 12545
rect 19568 12480 19576 12544
rect 19640 12480 19656 12544
rect 19720 12480 19736 12544
rect 19800 12480 19816 12544
rect 19880 12480 19888 12544
rect 19568 12479 19888 12480
rect 11513 12338 11579 12341
rect 16757 12338 16823 12341
rect 11513 12336 16823 12338
rect 11513 12280 11518 12336
rect 11574 12280 16762 12336
rect 16818 12280 16823 12336
rect 11513 12278 16823 12280
rect 11513 12275 11579 12278
rect 16757 12275 16823 12278
rect 0 12066 800 12096
rect 3049 12066 3115 12069
rect 0 12064 3115 12066
rect 0 12008 3054 12064
rect 3110 12008 3115 12064
rect 0 12006 3115 12008
rect 0 11976 800 12006
rect 3049 12003 3115 12006
rect 4208 12000 4528 12001
rect 4208 11936 4216 12000
rect 4280 11936 4296 12000
rect 4360 11936 4376 12000
rect 4440 11936 4456 12000
rect 4520 11936 4528 12000
rect 4208 11935 4528 11936
rect 34928 12000 35248 12001
rect 34928 11936 34936 12000
rect 35000 11936 35016 12000
rect 35080 11936 35096 12000
rect 35160 11936 35176 12000
rect 35240 11936 35248 12000
rect 34928 11935 35248 11936
rect 20253 11658 20319 11661
rect 20713 11658 20779 11661
rect 20253 11656 20779 11658
rect 20253 11600 20258 11656
rect 20314 11600 20718 11656
rect 20774 11600 20779 11656
rect 20253 11598 20779 11600
rect 20253 11595 20319 11598
rect 20713 11595 20779 11598
rect 19568 11456 19888 11457
rect 19568 11392 19576 11456
rect 19640 11392 19656 11456
rect 19720 11392 19736 11456
rect 19800 11392 19816 11456
rect 19880 11392 19888 11456
rect 19568 11391 19888 11392
rect 11237 11250 11303 11253
rect 24393 11250 24459 11253
rect 11237 11248 24459 11250
rect 11237 11192 11242 11248
rect 11298 11192 24398 11248
rect 24454 11192 24459 11248
rect 11237 11190 24459 11192
rect 11237 11187 11303 11190
rect 24393 11187 24459 11190
rect 4208 10912 4528 10913
rect 4208 10848 4216 10912
rect 4280 10848 4296 10912
rect 4360 10848 4376 10912
rect 4440 10848 4456 10912
rect 4520 10848 4528 10912
rect 4208 10847 4528 10848
rect 34928 10912 35248 10913
rect 34928 10848 34936 10912
rect 35000 10848 35016 10912
rect 35080 10848 35096 10912
rect 35160 10848 35176 10912
rect 35240 10848 35248 10912
rect 34928 10847 35248 10848
rect 19793 10842 19859 10845
rect 25497 10842 25563 10845
rect 19793 10840 25563 10842
rect 19793 10784 19798 10840
rect 19854 10784 25502 10840
rect 25558 10784 25563 10840
rect 19793 10782 25563 10784
rect 19793 10779 19859 10782
rect 25497 10779 25563 10782
rect 19568 10368 19888 10369
rect 19568 10304 19576 10368
rect 19640 10304 19656 10368
rect 19720 10304 19736 10368
rect 19800 10304 19816 10368
rect 19880 10304 19888 10368
rect 19568 10303 19888 10304
rect 37181 10162 37247 10165
rect 40200 10162 41000 10192
rect 37181 10160 41000 10162
rect 37181 10104 37186 10160
rect 37242 10104 41000 10160
rect 37181 10102 41000 10104
rect 37181 10099 37247 10102
rect 40200 10072 41000 10102
rect 11237 9890 11303 9893
rect 17401 9890 17467 9893
rect 11237 9888 17467 9890
rect 11237 9832 11242 9888
rect 11298 9832 17406 9888
rect 17462 9832 17467 9888
rect 11237 9830 17467 9832
rect 11237 9827 11303 9830
rect 17401 9827 17467 9830
rect 4208 9824 4528 9825
rect 4208 9760 4216 9824
rect 4280 9760 4296 9824
rect 4360 9760 4376 9824
rect 4440 9760 4456 9824
rect 4520 9760 4528 9824
rect 4208 9759 4528 9760
rect 34928 9824 35248 9825
rect 34928 9760 34936 9824
rect 35000 9760 35016 9824
rect 35080 9760 35096 9824
rect 35160 9760 35176 9824
rect 35240 9760 35248 9824
rect 34928 9759 35248 9760
rect 10041 9618 10107 9621
rect 12249 9618 12315 9621
rect 12525 9618 12591 9621
rect 10041 9616 12591 9618
rect 10041 9560 10046 9616
rect 10102 9560 12254 9616
rect 12310 9560 12530 9616
rect 12586 9560 12591 9616
rect 10041 9558 12591 9560
rect 10041 9555 10107 9558
rect 12249 9555 12315 9558
rect 12525 9555 12591 9558
rect 16665 9618 16731 9621
rect 24945 9618 25011 9621
rect 31845 9618 31911 9621
rect 16665 9616 31911 9618
rect 16665 9560 16670 9616
rect 16726 9560 24950 9616
rect 25006 9560 31850 9616
rect 31906 9560 31911 9616
rect 16665 9558 31911 9560
rect 16665 9555 16731 9558
rect 24945 9555 25011 9558
rect 31845 9555 31911 9558
rect 12525 9482 12591 9485
rect 12893 9482 12959 9485
rect 12525 9480 12959 9482
rect 12525 9424 12530 9480
rect 12586 9424 12898 9480
rect 12954 9424 12959 9480
rect 12525 9422 12959 9424
rect 12525 9419 12591 9422
rect 12893 9419 12959 9422
rect 19885 9482 19951 9485
rect 23657 9482 23723 9485
rect 25405 9482 25471 9485
rect 19885 9480 25471 9482
rect 19885 9424 19890 9480
rect 19946 9424 23662 9480
rect 23718 9424 25410 9480
rect 25466 9424 25471 9480
rect 19885 9422 25471 9424
rect 19885 9419 19951 9422
rect 23657 9419 23723 9422
rect 25405 9419 25471 9422
rect 0 9346 800 9376
rect 4061 9346 4127 9349
rect 0 9344 4127 9346
rect 0 9288 4066 9344
rect 4122 9288 4127 9344
rect 0 9286 4127 9288
rect 0 9256 800 9286
rect 4061 9283 4127 9286
rect 19568 9280 19888 9281
rect 19568 9216 19576 9280
rect 19640 9216 19656 9280
rect 19720 9216 19736 9280
rect 19800 9216 19816 9280
rect 19880 9216 19888 9280
rect 19568 9215 19888 9216
rect 29913 9210 29979 9213
rect 35341 9210 35407 9213
rect 29913 9208 35407 9210
rect 29913 9152 29918 9208
rect 29974 9152 35346 9208
rect 35402 9152 35407 9208
rect 29913 9150 35407 9152
rect 29913 9147 29979 9150
rect 35341 9147 35407 9150
rect 29729 9074 29795 9077
rect 33133 9074 33199 9077
rect 29729 9072 33199 9074
rect 29729 9016 29734 9072
rect 29790 9016 33138 9072
rect 33194 9016 33199 9072
rect 29729 9014 33199 9016
rect 29729 9011 29795 9014
rect 33133 9011 33199 9014
rect 4208 8736 4528 8737
rect 4208 8672 4216 8736
rect 4280 8672 4296 8736
rect 4360 8672 4376 8736
rect 4440 8672 4456 8736
rect 4520 8672 4528 8736
rect 4208 8671 4528 8672
rect 34928 8736 35248 8737
rect 34928 8672 34936 8736
rect 35000 8672 35016 8736
rect 35080 8672 35096 8736
rect 35160 8672 35176 8736
rect 35240 8672 35248 8736
rect 34928 8671 35248 8672
rect 19977 8666 20043 8669
rect 21173 8666 21239 8669
rect 19977 8664 21239 8666
rect 19977 8608 19982 8664
rect 20038 8608 21178 8664
rect 21234 8608 21239 8664
rect 19977 8606 21239 8608
rect 19977 8603 20043 8606
rect 21173 8603 21239 8606
rect 15101 8530 15167 8533
rect 31569 8530 31635 8533
rect 15101 8528 31635 8530
rect 15101 8472 15106 8528
rect 15162 8472 31574 8528
rect 31630 8472 31635 8528
rect 15101 8470 31635 8472
rect 15101 8467 15167 8470
rect 31569 8467 31635 8470
rect 19057 8394 19123 8397
rect 19241 8394 19307 8397
rect 22645 8394 22711 8397
rect 19057 8392 22711 8394
rect 19057 8336 19062 8392
rect 19118 8336 19246 8392
rect 19302 8336 22650 8392
rect 22706 8336 22711 8392
rect 19057 8334 22711 8336
rect 19057 8331 19123 8334
rect 19241 8331 19307 8334
rect 22645 8331 22711 8334
rect 19568 8192 19888 8193
rect 19568 8128 19576 8192
rect 19640 8128 19656 8192
rect 19720 8128 19736 8192
rect 19800 8128 19816 8192
rect 19880 8128 19888 8192
rect 19568 8127 19888 8128
rect 21817 7986 21883 7989
rect 23013 7986 23079 7989
rect 23657 7986 23723 7989
rect 21817 7984 23723 7986
rect 21817 7928 21822 7984
rect 21878 7928 23018 7984
rect 23074 7928 23662 7984
rect 23718 7928 23723 7984
rect 21817 7926 23723 7928
rect 21817 7923 21883 7926
rect 23013 7923 23079 7926
rect 23657 7923 23723 7926
rect 9857 7850 9923 7853
rect 26233 7850 26299 7853
rect 9857 7848 26299 7850
rect 9857 7792 9862 7848
rect 9918 7792 26238 7848
rect 26294 7792 26299 7848
rect 9857 7790 26299 7792
rect 9857 7787 9923 7790
rect 26233 7787 26299 7790
rect 4208 7648 4528 7649
rect 4208 7584 4216 7648
rect 4280 7584 4296 7648
rect 4360 7584 4376 7648
rect 4440 7584 4456 7648
rect 4520 7584 4528 7648
rect 4208 7583 4528 7584
rect 34928 7648 35248 7649
rect 34928 7584 34936 7648
rect 35000 7584 35016 7648
rect 35080 7584 35096 7648
rect 35160 7584 35176 7648
rect 35240 7584 35248 7648
rect 34928 7583 35248 7584
rect 10869 7442 10935 7445
rect 14457 7442 14523 7445
rect 10869 7440 14523 7442
rect 10869 7384 10874 7440
rect 10930 7384 14462 7440
rect 14518 7384 14523 7440
rect 10869 7382 14523 7384
rect 10869 7379 10935 7382
rect 14457 7379 14523 7382
rect 38561 7442 38627 7445
rect 40200 7442 41000 7472
rect 38561 7440 41000 7442
rect 38561 7384 38566 7440
rect 38622 7384 41000 7440
rect 38561 7382 41000 7384
rect 38561 7379 38627 7382
rect 40200 7352 41000 7382
rect 1577 7306 1643 7309
rect 21398 7306 21404 7308
rect 1577 7304 21404 7306
rect 1577 7248 1582 7304
rect 1638 7248 21404 7304
rect 1577 7246 21404 7248
rect 1577 7243 1643 7246
rect 21398 7244 21404 7246
rect 21468 7244 21474 7308
rect 19568 7104 19888 7105
rect 19568 7040 19576 7104
rect 19640 7040 19656 7104
rect 19720 7040 19736 7104
rect 19800 7040 19816 7104
rect 19880 7040 19888 7104
rect 19568 7039 19888 7040
rect 19241 6898 19307 6901
rect 19374 6898 19380 6900
rect 19241 6896 19380 6898
rect 19241 6840 19246 6896
rect 19302 6840 19380 6896
rect 19241 6838 19380 6840
rect 19241 6835 19307 6838
rect 19374 6836 19380 6838
rect 19444 6836 19450 6900
rect 4208 6560 4528 6561
rect 4208 6496 4216 6560
rect 4280 6496 4296 6560
rect 4360 6496 4376 6560
rect 4440 6496 4456 6560
rect 4520 6496 4528 6560
rect 4208 6495 4528 6496
rect 34928 6560 35248 6561
rect 34928 6496 34936 6560
rect 35000 6496 35016 6560
rect 35080 6496 35096 6560
rect 35160 6496 35176 6560
rect 35240 6496 35248 6560
rect 34928 6495 35248 6496
rect 0 6354 800 6384
rect 3969 6354 4035 6357
rect 0 6352 4035 6354
rect 0 6296 3974 6352
rect 4030 6296 4035 6352
rect 0 6294 4035 6296
rect 0 6264 800 6294
rect 3969 6291 4035 6294
rect 29085 6218 29151 6221
rect 31845 6218 31911 6221
rect 29085 6216 31911 6218
rect 29085 6160 29090 6216
rect 29146 6160 31850 6216
rect 31906 6160 31911 6216
rect 29085 6158 31911 6160
rect 29085 6155 29151 6158
rect 31845 6155 31911 6158
rect 19568 6016 19888 6017
rect 19568 5952 19576 6016
rect 19640 5952 19656 6016
rect 19720 5952 19736 6016
rect 19800 5952 19816 6016
rect 19880 5952 19888 6016
rect 19568 5951 19888 5952
rect 4208 5472 4528 5473
rect 4208 5408 4216 5472
rect 4280 5408 4296 5472
rect 4360 5408 4376 5472
rect 4440 5408 4456 5472
rect 4520 5408 4528 5472
rect 4208 5407 4528 5408
rect 34928 5472 35248 5473
rect 34928 5408 34936 5472
rect 35000 5408 35016 5472
rect 35080 5408 35096 5472
rect 35160 5408 35176 5472
rect 35240 5408 35248 5472
rect 34928 5407 35248 5408
rect 19568 4928 19888 4929
rect 19568 4864 19576 4928
rect 19640 4864 19656 4928
rect 19720 4864 19736 4928
rect 19800 4864 19816 4928
rect 19880 4864 19888 4928
rect 19568 4863 19888 4864
rect 35341 4450 35407 4453
rect 40200 4450 41000 4480
rect 35341 4448 41000 4450
rect 35341 4392 35346 4448
rect 35402 4392 41000 4448
rect 35341 4390 41000 4392
rect 35341 4387 35407 4390
rect 4208 4384 4528 4385
rect 4208 4320 4216 4384
rect 4280 4320 4296 4384
rect 4360 4320 4376 4384
rect 4440 4320 4456 4384
rect 4520 4320 4528 4384
rect 4208 4319 4528 4320
rect 34928 4384 35248 4385
rect 34928 4320 34936 4384
rect 35000 4320 35016 4384
rect 35080 4320 35096 4384
rect 35160 4320 35176 4384
rect 35240 4320 35248 4384
rect 40200 4360 41000 4390
rect 34928 4319 35248 4320
rect 21725 4042 21791 4045
rect 28441 4042 28507 4045
rect 21725 4040 28507 4042
rect 21725 3984 21730 4040
rect 21786 3984 28446 4040
rect 28502 3984 28507 4040
rect 21725 3982 28507 3984
rect 21725 3979 21791 3982
rect 28441 3979 28507 3982
rect 33685 3906 33751 3909
rect 35893 3906 35959 3909
rect 33685 3904 35959 3906
rect 33685 3848 33690 3904
rect 33746 3848 35898 3904
rect 35954 3848 35959 3904
rect 33685 3846 35959 3848
rect 33685 3843 33751 3846
rect 35893 3843 35959 3846
rect 19568 3840 19888 3841
rect 19568 3776 19576 3840
rect 19640 3776 19656 3840
rect 19720 3776 19736 3840
rect 19800 3776 19816 3840
rect 19880 3776 19888 3840
rect 19568 3775 19888 3776
rect 0 3634 800 3664
rect 3417 3634 3483 3637
rect 0 3632 3483 3634
rect 0 3576 3422 3632
rect 3478 3576 3483 3632
rect 0 3574 3483 3576
rect 0 3544 800 3574
rect 3417 3571 3483 3574
rect 17861 3634 17927 3637
rect 27102 3634 27108 3636
rect 17861 3632 27108 3634
rect 17861 3576 17866 3632
rect 17922 3576 27108 3632
rect 17861 3574 27108 3576
rect 17861 3571 17927 3574
rect 27102 3572 27108 3574
rect 27172 3572 27178 3636
rect 8109 3498 8175 3501
rect 28073 3498 28139 3501
rect 8109 3496 28139 3498
rect 8109 3440 8114 3496
rect 8170 3440 28078 3496
rect 28134 3440 28139 3496
rect 8109 3438 28139 3440
rect 8109 3435 8175 3438
rect 28073 3435 28139 3438
rect 6269 3362 6335 3365
rect 29913 3362 29979 3365
rect 6269 3360 29979 3362
rect 6269 3304 6274 3360
rect 6330 3304 29918 3360
rect 29974 3304 29979 3360
rect 6269 3302 29979 3304
rect 6269 3299 6335 3302
rect 29913 3299 29979 3302
rect 4208 3296 4528 3297
rect 4208 3232 4216 3296
rect 4280 3232 4296 3296
rect 4360 3232 4376 3296
rect 4440 3232 4456 3296
rect 4520 3232 4528 3296
rect 4208 3231 4528 3232
rect 34928 3296 35248 3297
rect 34928 3232 34936 3296
rect 35000 3232 35016 3296
rect 35080 3232 35096 3296
rect 35160 3232 35176 3296
rect 35240 3232 35248 3296
rect 34928 3231 35248 3232
rect 7281 2954 7347 2957
rect 9581 2954 9647 2957
rect 7281 2952 9647 2954
rect 7281 2896 7286 2952
rect 7342 2896 9586 2952
rect 9642 2896 9647 2952
rect 7281 2894 9647 2896
rect 7281 2891 7347 2894
rect 9581 2891 9647 2894
rect 19568 2752 19888 2753
rect 19568 2688 19576 2752
rect 19640 2688 19656 2752
rect 19720 2688 19736 2752
rect 19800 2688 19816 2752
rect 19880 2688 19888 2752
rect 19568 2687 19888 2688
rect 4208 2208 4528 2209
rect 4208 2144 4216 2208
rect 4280 2144 4296 2208
rect 4360 2144 4376 2208
rect 4440 2144 4456 2208
rect 4520 2144 4528 2208
rect 4208 2143 4528 2144
rect 34928 2208 35248 2209
rect 34928 2144 34936 2208
rect 35000 2144 35016 2208
rect 35080 2144 35096 2208
rect 35160 2144 35176 2208
rect 35240 2144 35248 2208
rect 34928 2143 35248 2144
rect 37089 1730 37155 1733
rect 40200 1730 41000 1760
rect 37089 1728 41000 1730
rect 37089 1672 37094 1728
rect 37150 1672 41000 1728
rect 37089 1670 41000 1672
rect 37089 1667 37155 1670
rect 40200 1640 41000 1670
<< via3 >>
rect 19576 38652 19640 38656
rect 19576 38596 19580 38652
rect 19580 38596 19636 38652
rect 19636 38596 19640 38652
rect 19576 38592 19640 38596
rect 19656 38652 19720 38656
rect 19656 38596 19660 38652
rect 19660 38596 19716 38652
rect 19716 38596 19720 38652
rect 19656 38592 19720 38596
rect 19736 38652 19800 38656
rect 19736 38596 19740 38652
rect 19740 38596 19796 38652
rect 19796 38596 19800 38652
rect 19736 38592 19800 38596
rect 19816 38652 19880 38656
rect 19816 38596 19820 38652
rect 19820 38596 19876 38652
rect 19876 38596 19880 38652
rect 19816 38592 19880 38596
rect 4216 38108 4280 38112
rect 4216 38052 4220 38108
rect 4220 38052 4276 38108
rect 4276 38052 4280 38108
rect 4216 38048 4280 38052
rect 4296 38108 4360 38112
rect 4296 38052 4300 38108
rect 4300 38052 4356 38108
rect 4356 38052 4360 38108
rect 4296 38048 4360 38052
rect 4376 38108 4440 38112
rect 4376 38052 4380 38108
rect 4380 38052 4436 38108
rect 4436 38052 4440 38108
rect 4376 38048 4440 38052
rect 4456 38108 4520 38112
rect 4456 38052 4460 38108
rect 4460 38052 4516 38108
rect 4516 38052 4520 38108
rect 4456 38048 4520 38052
rect 34936 38108 35000 38112
rect 34936 38052 34940 38108
rect 34940 38052 34996 38108
rect 34996 38052 35000 38108
rect 34936 38048 35000 38052
rect 35016 38108 35080 38112
rect 35016 38052 35020 38108
rect 35020 38052 35076 38108
rect 35076 38052 35080 38108
rect 35016 38048 35080 38052
rect 35096 38108 35160 38112
rect 35096 38052 35100 38108
rect 35100 38052 35156 38108
rect 35156 38052 35160 38108
rect 35096 38048 35160 38052
rect 35176 38108 35240 38112
rect 35176 38052 35180 38108
rect 35180 38052 35236 38108
rect 35236 38052 35240 38108
rect 35176 38048 35240 38052
rect 19576 37564 19640 37568
rect 19576 37508 19580 37564
rect 19580 37508 19636 37564
rect 19636 37508 19640 37564
rect 19576 37504 19640 37508
rect 19656 37564 19720 37568
rect 19656 37508 19660 37564
rect 19660 37508 19716 37564
rect 19716 37508 19720 37564
rect 19656 37504 19720 37508
rect 19736 37564 19800 37568
rect 19736 37508 19740 37564
rect 19740 37508 19796 37564
rect 19796 37508 19800 37564
rect 19736 37504 19800 37508
rect 19816 37564 19880 37568
rect 19816 37508 19820 37564
rect 19820 37508 19876 37564
rect 19876 37508 19880 37564
rect 19816 37504 19880 37508
rect 4216 37020 4280 37024
rect 4216 36964 4220 37020
rect 4220 36964 4276 37020
rect 4276 36964 4280 37020
rect 4216 36960 4280 36964
rect 4296 37020 4360 37024
rect 4296 36964 4300 37020
rect 4300 36964 4356 37020
rect 4356 36964 4360 37020
rect 4296 36960 4360 36964
rect 4376 37020 4440 37024
rect 4376 36964 4380 37020
rect 4380 36964 4436 37020
rect 4436 36964 4440 37020
rect 4376 36960 4440 36964
rect 4456 37020 4520 37024
rect 4456 36964 4460 37020
rect 4460 36964 4516 37020
rect 4516 36964 4520 37020
rect 4456 36960 4520 36964
rect 34936 37020 35000 37024
rect 34936 36964 34940 37020
rect 34940 36964 34996 37020
rect 34996 36964 35000 37020
rect 34936 36960 35000 36964
rect 35016 37020 35080 37024
rect 35016 36964 35020 37020
rect 35020 36964 35076 37020
rect 35076 36964 35080 37020
rect 35016 36960 35080 36964
rect 35096 37020 35160 37024
rect 35096 36964 35100 37020
rect 35100 36964 35156 37020
rect 35156 36964 35160 37020
rect 35096 36960 35160 36964
rect 35176 37020 35240 37024
rect 35176 36964 35180 37020
rect 35180 36964 35236 37020
rect 35236 36964 35240 37020
rect 35176 36960 35240 36964
rect 19576 36476 19640 36480
rect 19576 36420 19580 36476
rect 19580 36420 19636 36476
rect 19636 36420 19640 36476
rect 19576 36416 19640 36420
rect 19656 36476 19720 36480
rect 19656 36420 19660 36476
rect 19660 36420 19716 36476
rect 19716 36420 19720 36476
rect 19656 36416 19720 36420
rect 19736 36476 19800 36480
rect 19736 36420 19740 36476
rect 19740 36420 19796 36476
rect 19796 36420 19800 36476
rect 19736 36416 19800 36420
rect 19816 36476 19880 36480
rect 19816 36420 19820 36476
rect 19820 36420 19876 36476
rect 19876 36420 19880 36476
rect 19816 36416 19880 36420
rect 4216 35932 4280 35936
rect 4216 35876 4220 35932
rect 4220 35876 4276 35932
rect 4276 35876 4280 35932
rect 4216 35872 4280 35876
rect 4296 35932 4360 35936
rect 4296 35876 4300 35932
rect 4300 35876 4356 35932
rect 4356 35876 4360 35932
rect 4296 35872 4360 35876
rect 4376 35932 4440 35936
rect 4376 35876 4380 35932
rect 4380 35876 4436 35932
rect 4436 35876 4440 35932
rect 4376 35872 4440 35876
rect 4456 35932 4520 35936
rect 4456 35876 4460 35932
rect 4460 35876 4516 35932
rect 4516 35876 4520 35932
rect 4456 35872 4520 35876
rect 34936 35932 35000 35936
rect 34936 35876 34940 35932
rect 34940 35876 34996 35932
rect 34996 35876 35000 35932
rect 34936 35872 35000 35876
rect 35016 35932 35080 35936
rect 35016 35876 35020 35932
rect 35020 35876 35076 35932
rect 35076 35876 35080 35932
rect 35016 35872 35080 35876
rect 35096 35932 35160 35936
rect 35096 35876 35100 35932
rect 35100 35876 35156 35932
rect 35156 35876 35160 35932
rect 35096 35872 35160 35876
rect 35176 35932 35240 35936
rect 35176 35876 35180 35932
rect 35180 35876 35236 35932
rect 35236 35876 35240 35932
rect 35176 35872 35240 35876
rect 19576 35388 19640 35392
rect 19576 35332 19580 35388
rect 19580 35332 19636 35388
rect 19636 35332 19640 35388
rect 19576 35328 19640 35332
rect 19656 35388 19720 35392
rect 19656 35332 19660 35388
rect 19660 35332 19716 35388
rect 19716 35332 19720 35388
rect 19656 35328 19720 35332
rect 19736 35388 19800 35392
rect 19736 35332 19740 35388
rect 19740 35332 19796 35388
rect 19796 35332 19800 35388
rect 19736 35328 19800 35332
rect 19816 35388 19880 35392
rect 19816 35332 19820 35388
rect 19820 35332 19876 35388
rect 19876 35332 19880 35388
rect 19816 35328 19880 35332
rect 4216 34844 4280 34848
rect 4216 34788 4220 34844
rect 4220 34788 4276 34844
rect 4276 34788 4280 34844
rect 4216 34784 4280 34788
rect 4296 34844 4360 34848
rect 4296 34788 4300 34844
rect 4300 34788 4356 34844
rect 4356 34788 4360 34844
rect 4296 34784 4360 34788
rect 4376 34844 4440 34848
rect 4376 34788 4380 34844
rect 4380 34788 4436 34844
rect 4436 34788 4440 34844
rect 4376 34784 4440 34788
rect 4456 34844 4520 34848
rect 4456 34788 4460 34844
rect 4460 34788 4516 34844
rect 4516 34788 4520 34844
rect 4456 34784 4520 34788
rect 34936 34844 35000 34848
rect 34936 34788 34940 34844
rect 34940 34788 34996 34844
rect 34996 34788 35000 34844
rect 34936 34784 35000 34788
rect 35016 34844 35080 34848
rect 35016 34788 35020 34844
rect 35020 34788 35076 34844
rect 35076 34788 35080 34844
rect 35016 34784 35080 34788
rect 35096 34844 35160 34848
rect 35096 34788 35100 34844
rect 35100 34788 35156 34844
rect 35156 34788 35160 34844
rect 35096 34784 35160 34788
rect 35176 34844 35240 34848
rect 35176 34788 35180 34844
rect 35180 34788 35236 34844
rect 35236 34788 35240 34844
rect 35176 34784 35240 34788
rect 19576 34300 19640 34304
rect 19576 34244 19580 34300
rect 19580 34244 19636 34300
rect 19636 34244 19640 34300
rect 19576 34240 19640 34244
rect 19656 34300 19720 34304
rect 19656 34244 19660 34300
rect 19660 34244 19716 34300
rect 19716 34244 19720 34300
rect 19656 34240 19720 34244
rect 19736 34300 19800 34304
rect 19736 34244 19740 34300
rect 19740 34244 19796 34300
rect 19796 34244 19800 34300
rect 19736 34240 19800 34244
rect 19816 34300 19880 34304
rect 19816 34244 19820 34300
rect 19820 34244 19876 34300
rect 19876 34244 19880 34300
rect 19816 34240 19880 34244
rect 4216 33756 4280 33760
rect 4216 33700 4220 33756
rect 4220 33700 4276 33756
rect 4276 33700 4280 33756
rect 4216 33696 4280 33700
rect 4296 33756 4360 33760
rect 4296 33700 4300 33756
rect 4300 33700 4356 33756
rect 4356 33700 4360 33756
rect 4296 33696 4360 33700
rect 4376 33756 4440 33760
rect 4376 33700 4380 33756
rect 4380 33700 4436 33756
rect 4436 33700 4440 33756
rect 4376 33696 4440 33700
rect 4456 33756 4520 33760
rect 4456 33700 4460 33756
rect 4460 33700 4516 33756
rect 4516 33700 4520 33756
rect 4456 33696 4520 33700
rect 34936 33756 35000 33760
rect 34936 33700 34940 33756
rect 34940 33700 34996 33756
rect 34996 33700 35000 33756
rect 34936 33696 35000 33700
rect 35016 33756 35080 33760
rect 35016 33700 35020 33756
rect 35020 33700 35076 33756
rect 35076 33700 35080 33756
rect 35016 33696 35080 33700
rect 35096 33756 35160 33760
rect 35096 33700 35100 33756
rect 35100 33700 35156 33756
rect 35156 33700 35160 33756
rect 35096 33696 35160 33700
rect 35176 33756 35240 33760
rect 35176 33700 35180 33756
rect 35180 33700 35236 33756
rect 35236 33700 35240 33756
rect 35176 33696 35240 33700
rect 19576 33212 19640 33216
rect 19576 33156 19580 33212
rect 19580 33156 19636 33212
rect 19636 33156 19640 33212
rect 19576 33152 19640 33156
rect 19656 33212 19720 33216
rect 19656 33156 19660 33212
rect 19660 33156 19716 33212
rect 19716 33156 19720 33212
rect 19656 33152 19720 33156
rect 19736 33212 19800 33216
rect 19736 33156 19740 33212
rect 19740 33156 19796 33212
rect 19796 33156 19800 33212
rect 19736 33152 19800 33156
rect 19816 33212 19880 33216
rect 19816 33156 19820 33212
rect 19820 33156 19876 33212
rect 19876 33156 19880 33212
rect 19816 33152 19880 33156
rect 4216 32668 4280 32672
rect 4216 32612 4220 32668
rect 4220 32612 4276 32668
rect 4276 32612 4280 32668
rect 4216 32608 4280 32612
rect 4296 32668 4360 32672
rect 4296 32612 4300 32668
rect 4300 32612 4356 32668
rect 4356 32612 4360 32668
rect 4296 32608 4360 32612
rect 4376 32668 4440 32672
rect 4376 32612 4380 32668
rect 4380 32612 4436 32668
rect 4436 32612 4440 32668
rect 4376 32608 4440 32612
rect 4456 32668 4520 32672
rect 4456 32612 4460 32668
rect 4460 32612 4516 32668
rect 4516 32612 4520 32668
rect 4456 32608 4520 32612
rect 34936 32668 35000 32672
rect 34936 32612 34940 32668
rect 34940 32612 34996 32668
rect 34996 32612 35000 32668
rect 34936 32608 35000 32612
rect 35016 32668 35080 32672
rect 35016 32612 35020 32668
rect 35020 32612 35076 32668
rect 35076 32612 35080 32668
rect 35016 32608 35080 32612
rect 35096 32668 35160 32672
rect 35096 32612 35100 32668
rect 35100 32612 35156 32668
rect 35156 32612 35160 32668
rect 35096 32608 35160 32612
rect 35176 32668 35240 32672
rect 35176 32612 35180 32668
rect 35180 32612 35236 32668
rect 35236 32612 35240 32668
rect 35176 32608 35240 32612
rect 19576 32124 19640 32128
rect 19576 32068 19580 32124
rect 19580 32068 19636 32124
rect 19636 32068 19640 32124
rect 19576 32064 19640 32068
rect 19656 32124 19720 32128
rect 19656 32068 19660 32124
rect 19660 32068 19716 32124
rect 19716 32068 19720 32124
rect 19656 32064 19720 32068
rect 19736 32124 19800 32128
rect 19736 32068 19740 32124
rect 19740 32068 19796 32124
rect 19796 32068 19800 32124
rect 19736 32064 19800 32068
rect 19816 32124 19880 32128
rect 19816 32068 19820 32124
rect 19820 32068 19876 32124
rect 19876 32068 19880 32124
rect 19816 32064 19880 32068
rect 37780 32056 37844 32060
rect 37780 32000 37794 32056
rect 37794 32000 37844 32056
rect 37780 31996 37844 32000
rect 4216 31580 4280 31584
rect 4216 31524 4220 31580
rect 4220 31524 4276 31580
rect 4276 31524 4280 31580
rect 4216 31520 4280 31524
rect 4296 31580 4360 31584
rect 4296 31524 4300 31580
rect 4300 31524 4356 31580
rect 4356 31524 4360 31580
rect 4296 31520 4360 31524
rect 4376 31580 4440 31584
rect 4376 31524 4380 31580
rect 4380 31524 4436 31580
rect 4436 31524 4440 31580
rect 4376 31520 4440 31524
rect 4456 31580 4520 31584
rect 4456 31524 4460 31580
rect 4460 31524 4516 31580
rect 4516 31524 4520 31580
rect 4456 31520 4520 31524
rect 34936 31580 35000 31584
rect 34936 31524 34940 31580
rect 34940 31524 34996 31580
rect 34996 31524 35000 31580
rect 34936 31520 35000 31524
rect 35016 31580 35080 31584
rect 35016 31524 35020 31580
rect 35020 31524 35076 31580
rect 35076 31524 35080 31580
rect 35016 31520 35080 31524
rect 35096 31580 35160 31584
rect 35096 31524 35100 31580
rect 35100 31524 35156 31580
rect 35156 31524 35160 31580
rect 35096 31520 35160 31524
rect 35176 31580 35240 31584
rect 35176 31524 35180 31580
rect 35180 31524 35236 31580
rect 35236 31524 35240 31580
rect 35176 31520 35240 31524
rect 19576 31036 19640 31040
rect 19576 30980 19580 31036
rect 19580 30980 19636 31036
rect 19636 30980 19640 31036
rect 19576 30976 19640 30980
rect 19656 31036 19720 31040
rect 19656 30980 19660 31036
rect 19660 30980 19716 31036
rect 19716 30980 19720 31036
rect 19656 30976 19720 30980
rect 19736 31036 19800 31040
rect 19736 30980 19740 31036
rect 19740 30980 19796 31036
rect 19796 30980 19800 31036
rect 19736 30976 19800 30980
rect 19816 31036 19880 31040
rect 19816 30980 19820 31036
rect 19820 30980 19876 31036
rect 19876 30980 19880 31036
rect 19816 30976 19880 30980
rect 27108 30696 27172 30700
rect 27108 30640 27122 30696
rect 27122 30640 27172 30696
rect 27108 30636 27172 30640
rect 4216 30492 4280 30496
rect 4216 30436 4220 30492
rect 4220 30436 4276 30492
rect 4276 30436 4280 30492
rect 4216 30432 4280 30436
rect 4296 30492 4360 30496
rect 4296 30436 4300 30492
rect 4300 30436 4356 30492
rect 4356 30436 4360 30492
rect 4296 30432 4360 30436
rect 4376 30492 4440 30496
rect 4376 30436 4380 30492
rect 4380 30436 4436 30492
rect 4436 30436 4440 30492
rect 4376 30432 4440 30436
rect 4456 30492 4520 30496
rect 4456 30436 4460 30492
rect 4460 30436 4516 30492
rect 4516 30436 4520 30492
rect 4456 30432 4520 30436
rect 34936 30492 35000 30496
rect 34936 30436 34940 30492
rect 34940 30436 34996 30492
rect 34996 30436 35000 30492
rect 34936 30432 35000 30436
rect 35016 30492 35080 30496
rect 35016 30436 35020 30492
rect 35020 30436 35076 30492
rect 35076 30436 35080 30492
rect 35016 30432 35080 30436
rect 35096 30492 35160 30496
rect 35096 30436 35100 30492
rect 35100 30436 35156 30492
rect 35156 30436 35160 30492
rect 35096 30432 35160 30436
rect 35176 30492 35240 30496
rect 35176 30436 35180 30492
rect 35180 30436 35236 30492
rect 35236 30436 35240 30492
rect 35176 30432 35240 30436
rect 19576 29948 19640 29952
rect 19576 29892 19580 29948
rect 19580 29892 19636 29948
rect 19636 29892 19640 29948
rect 19576 29888 19640 29892
rect 19656 29948 19720 29952
rect 19656 29892 19660 29948
rect 19660 29892 19716 29948
rect 19716 29892 19720 29948
rect 19656 29888 19720 29892
rect 19736 29948 19800 29952
rect 19736 29892 19740 29948
rect 19740 29892 19796 29948
rect 19796 29892 19800 29948
rect 19736 29888 19800 29892
rect 19816 29948 19880 29952
rect 19816 29892 19820 29948
rect 19820 29892 19876 29948
rect 19876 29892 19880 29948
rect 19816 29888 19880 29892
rect 4216 29404 4280 29408
rect 4216 29348 4220 29404
rect 4220 29348 4276 29404
rect 4276 29348 4280 29404
rect 4216 29344 4280 29348
rect 4296 29404 4360 29408
rect 4296 29348 4300 29404
rect 4300 29348 4356 29404
rect 4356 29348 4360 29404
rect 4296 29344 4360 29348
rect 4376 29404 4440 29408
rect 4376 29348 4380 29404
rect 4380 29348 4436 29404
rect 4436 29348 4440 29404
rect 4376 29344 4440 29348
rect 4456 29404 4520 29408
rect 4456 29348 4460 29404
rect 4460 29348 4516 29404
rect 4516 29348 4520 29404
rect 4456 29344 4520 29348
rect 34936 29404 35000 29408
rect 34936 29348 34940 29404
rect 34940 29348 34996 29404
rect 34996 29348 35000 29404
rect 34936 29344 35000 29348
rect 35016 29404 35080 29408
rect 35016 29348 35020 29404
rect 35020 29348 35076 29404
rect 35076 29348 35080 29404
rect 35016 29344 35080 29348
rect 35096 29404 35160 29408
rect 35096 29348 35100 29404
rect 35100 29348 35156 29404
rect 35156 29348 35160 29404
rect 35096 29344 35160 29348
rect 35176 29404 35240 29408
rect 35176 29348 35180 29404
rect 35180 29348 35236 29404
rect 35236 29348 35240 29404
rect 35176 29344 35240 29348
rect 19380 28928 19444 28932
rect 19380 28872 19430 28928
rect 19430 28872 19444 28928
rect 19380 28868 19444 28872
rect 19576 28860 19640 28864
rect 19576 28804 19580 28860
rect 19580 28804 19636 28860
rect 19636 28804 19640 28860
rect 19576 28800 19640 28804
rect 19656 28860 19720 28864
rect 19656 28804 19660 28860
rect 19660 28804 19716 28860
rect 19716 28804 19720 28860
rect 19656 28800 19720 28804
rect 19736 28860 19800 28864
rect 19736 28804 19740 28860
rect 19740 28804 19796 28860
rect 19796 28804 19800 28860
rect 19736 28800 19800 28804
rect 19816 28860 19880 28864
rect 19816 28804 19820 28860
rect 19820 28804 19876 28860
rect 19876 28804 19880 28860
rect 19816 28800 19880 28804
rect 4216 28316 4280 28320
rect 4216 28260 4220 28316
rect 4220 28260 4276 28316
rect 4276 28260 4280 28316
rect 4216 28256 4280 28260
rect 4296 28316 4360 28320
rect 4296 28260 4300 28316
rect 4300 28260 4356 28316
rect 4356 28260 4360 28316
rect 4296 28256 4360 28260
rect 4376 28316 4440 28320
rect 4376 28260 4380 28316
rect 4380 28260 4436 28316
rect 4436 28260 4440 28316
rect 4376 28256 4440 28260
rect 4456 28316 4520 28320
rect 4456 28260 4460 28316
rect 4460 28260 4516 28316
rect 4516 28260 4520 28316
rect 4456 28256 4520 28260
rect 34936 28316 35000 28320
rect 34936 28260 34940 28316
rect 34940 28260 34996 28316
rect 34996 28260 35000 28316
rect 34936 28256 35000 28260
rect 35016 28316 35080 28320
rect 35016 28260 35020 28316
rect 35020 28260 35076 28316
rect 35076 28260 35080 28316
rect 35016 28256 35080 28260
rect 35096 28316 35160 28320
rect 35096 28260 35100 28316
rect 35100 28260 35156 28316
rect 35156 28260 35160 28316
rect 35096 28256 35160 28260
rect 35176 28316 35240 28320
rect 35176 28260 35180 28316
rect 35180 28260 35236 28316
rect 35236 28260 35240 28316
rect 35176 28256 35240 28260
rect 19576 27772 19640 27776
rect 19576 27716 19580 27772
rect 19580 27716 19636 27772
rect 19636 27716 19640 27772
rect 19576 27712 19640 27716
rect 19656 27772 19720 27776
rect 19656 27716 19660 27772
rect 19660 27716 19716 27772
rect 19716 27716 19720 27772
rect 19656 27712 19720 27716
rect 19736 27772 19800 27776
rect 19736 27716 19740 27772
rect 19740 27716 19796 27772
rect 19796 27716 19800 27772
rect 19736 27712 19800 27716
rect 19816 27772 19880 27776
rect 19816 27716 19820 27772
rect 19820 27716 19876 27772
rect 19876 27716 19880 27772
rect 19816 27712 19880 27716
rect 4216 27228 4280 27232
rect 4216 27172 4220 27228
rect 4220 27172 4276 27228
rect 4276 27172 4280 27228
rect 4216 27168 4280 27172
rect 4296 27228 4360 27232
rect 4296 27172 4300 27228
rect 4300 27172 4356 27228
rect 4356 27172 4360 27228
rect 4296 27168 4360 27172
rect 4376 27228 4440 27232
rect 4376 27172 4380 27228
rect 4380 27172 4436 27228
rect 4436 27172 4440 27228
rect 4376 27168 4440 27172
rect 4456 27228 4520 27232
rect 4456 27172 4460 27228
rect 4460 27172 4516 27228
rect 4516 27172 4520 27228
rect 4456 27168 4520 27172
rect 34936 27228 35000 27232
rect 34936 27172 34940 27228
rect 34940 27172 34996 27228
rect 34996 27172 35000 27228
rect 34936 27168 35000 27172
rect 35016 27228 35080 27232
rect 35016 27172 35020 27228
rect 35020 27172 35076 27228
rect 35076 27172 35080 27228
rect 35016 27168 35080 27172
rect 35096 27228 35160 27232
rect 35096 27172 35100 27228
rect 35100 27172 35156 27228
rect 35156 27172 35160 27228
rect 35096 27168 35160 27172
rect 35176 27228 35240 27232
rect 35176 27172 35180 27228
rect 35180 27172 35236 27228
rect 35236 27172 35240 27228
rect 35176 27168 35240 27172
rect 19576 26684 19640 26688
rect 19576 26628 19580 26684
rect 19580 26628 19636 26684
rect 19636 26628 19640 26684
rect 19576 26624 19640 26628
rect 19656 26684 19720 26688
rect 19656 26628 19660 26684
rect 19660 26628 19716 26684
rect 19716 26628 19720 26684
rect 19656 26624 19720 26628
rect 19736 26684 19800 26688
rect 19736 26628 19740 26684
rect 19740 26628 19796 26684
rect 19796 26628 19800 26684
rect 19736 26624 19800 26628
rect 19816 26684 19880 26688
rect 19816 26628 19820 26684
rect 19820 26628 19876 26684
rect 19876 26628 19880 26684
rect 19816 26624 19880 26628
rect 4216 26140 4280 26144
rect 4216 26084 4220 26140
rect 4220 26084 4276 26140
rect 4276 26084 4280 26140
rect 4216 26080 4280 26084
rect 4296 26140 4360 26144
rect 4296 26084 4300 26140
rect 4300 26084 4356 26140
rect 4356 26084 4360 26140
rect 4296 26080 4360 26084
rect 4376 26140 4440 26144
rect 4376 26084 4380 26140
rect 4380 26084 4436 26140
rect 4436 26084 4440 26140
rect 4376 26080 4440 26084
rect 4456 26140 4520 26144
rect 4456 26084 4460 26140
rect 4460 26084 4516 26140
rect 4516 26084 4520 26140
rect 4456 26080 4520 26084
rect 34936 26140 35000 26144
rect 34936 26084 34940 26140
rect 34940 26084 34996 26140
rect 34996 26084 35000 26140
rect 34936 26080 35000 26084
rect 35016 26140 35080 26144
rect 35016 26084 35020 26140
rect 35020 26084 35076 26140
rect 35076 26084 35080 26140
rect 35016 26080 35080 26084
rect 35096 26140 35160 26144
rect 35096 26084 35100 26140
rect 35100 26084 35156 26140
rect 35156 26084 35160 26140
rect 35096 26080 35160 26084
rect 35176 26140 35240 26144
rect 35176 26084 35180 26140
rect 35180 26084 35236 26140
rect 35236 26084 35240 26140
rect 35176 26080 35240 26084
rect 19576 25596 19640 25600
rect 19576 25540 19580 25596
rect 19580 25540 19636 25596
rect 19636 25540 19640 25596
rect 19576 25536 19640 25540
rect 19656 25596 19720 25600
rect 19656 25540 19660 25596
rect 19660 25540 19716 25596
rect 19716 25540 19720 25596
rect 19656 25536 19720 25540
rect 19736 25596 19800 25600
rect 19736 25540 19740 25596
rect 19740 25540 19796 25596
rect 19796 25540 19800 25596
rect 19736 25536 19800 25540
rect 19816 25596 19880 25600
rect 19816 25540 19820 25596
rect 19820 25540 19876 25596
rect 19876 25540 19880 25596
rect 19816 25536 19880 25540
rect 4216 25052 4280 25056
rect 4216 24996 4220 25052
rect 4220 24996 4276 25052
rect 4276 24996 4280 25052
rect 4216 24992 4280 24996
rect 4296 25052 4360 25056
rect 4296 24996 4300 25052
rect 4300 24996 4356 25052
rect 4356 24996 4360 25052
rect 4296 24992 4360 24996
rect 4376 25052 4440 25056
rect 4376 24996 4380 25052
rect 4380 24996 4436 25052
rect 4436 24996 4440 25052
rect 4376 24992 4440 24996
rect 4456 25052 4520 25056
rect 4456 24996 4460 25052
rect 4460 24996 4516 25052
rect 4516 24996 4520 25052
rect 4456 24992 4520 24996
rect 34936 25052 35000 25056
rect 34936 24996 34940 25052
rect 34940 24996 34996 25052
rect 34996 24996 35000 25052
rect 34936 24992 35000 24996
rect 35016 25052 35080 25056
rect 35016 24996 35020 25052
rect 35020 24996 35076 25052
rect 35076 24996 35080 25052
rect 35016 24992 35080 24996
rect 35096 25052 35160 25056
rect 35096 24996 35100 25052
rect 35100 24996 35156 25052
rect 35156 24996 35160 25052
rect 35096 24992 35160 24996
rect 35176 25052 35240 25056
rect 35176 24996 35180 25052
rect 35180 24996 35236 25052
rect 35236 24996 35240 25052
rect 35176 24992 35240 24996
rect 19576 24508 19640 24512
rect 19576 24452 19580 24508
rect 19580 24452 19636 24508
rect 19636 24452 19640 24508
rect 19576 24448 19640 24452
rect 19656 24508 19720 24512
rect 19656 24452 19660 24508
rect 19660 24452 19716 24508
rect 19716 24452 19720 24508
rect 19656 24448 19720 24452
rect 19736 24508 19800 24512
rect 19736 24452 19740 24508
rect 19740 24452 19796 24508
rect 19796 24452 19800 24508
rect 19736 24448 19800 24452
rect 19816 24508 19880 24512
rect 19816 24452 19820 24508
rect 19820 24452 19876 24508
rect 19876 24452 19880 24508
rect 19816 24448 19880 24452
rect 4216 23964 4280 23968
rect 4216 23908 4220 23964
rect 4220 23908 4276 23964
rect 4276 23908 4280 23964
rect 4216 23904 4280 23908
rect 4296 23964 4360 23968
rect 4296 23908 4300 23964
rect 4300 23908 4356 23964
rect 4356 23908 4360 23964
rect 4296 23904 4360 23908
rect 4376 23964 4440 23968
rect 4376 23908 4380 23964
rect 4380 23908 4436 23964
rect 4436 23908 4440 23964
rect 4376 23904 4440 23908
rect 4456 23964 4520 23968
rect 4456 23908 4460 23964
rect 4460 23908 4516 23964
rect 4516 23908 4520 23964
rect 4456 23904 4520 23908
rect 34936 23964 35000 23968
rect 34936 23908 34940 23964
rect 34940 23908 34996 23964
rect 34996 23908 35000 23964
rect 34936 23904 35000 23908
rect 35016 23964 35080 23968
rect 35016 23908 35020 23964
rect 35020 23908 35076 23964
rect 35076 23908 35080 23964
rect 35016 23904 35080 23908
rect 35096 23964 35160 23968
rect 35096 23908 35100 23964
rect 35100 23908 35156 23964
rect 35156 23908 35160 23964
rect 35096 23904 35160 23908
rect 35176 23964 35240 23968
rect 35176 23908 35180 23964
rect 35180 23908 35236 23964
rect 35236 23908 35240 23964
rect 35176 23904 35240 23908
rect 19576 23420 19640 23424
rect 19576 23364 19580 23420
rect 19580 23364 19636 23420
rect 19636 23364 19640 23420
rect 19576 23360 19640 23364
rect 19656 23420 19720 23424
rect 19656 23364 19660 23420
rect 19660 23364 19716 23420
rect 19716 23364 19720 23420
rect 19656 23360 19720 23364
rect 19736 23420 19800 23424
rect 19736 23364 19740 23420
rect 19740 23364 19796 23420
rect 19796 23364 19800 23420
rect 19736 23360 19800 23364
rect 19816 23420 19880 23424
rect 19816 23364 19820 23420
rect 19820 23364 19876 23420
rect 19876 23364 19880 23420
rect 19816 23360 19880 23364
rect 19380 23352 19444 23356
rect 19380 23296 19430 23352
rect 19430 23296 19444 23352
rect 19380 23292 19444 23296
rect 4216 22876 4280 22880
rect 4216 22820 4220 22876
rect 4220 22820 4276 22876
rect 4276 22820 4280 22876
rect 4216 22816 4280 22820
rect 4296 22876 4360 22880
rect 4296 22820 4300 22876
rect 4300 22820 4356 22876
rect 4356 22820 4360 22876
rect 4296 22816 4360 22820
rect 4376 22876 4440 22880
rect 4376 22820 4380 22876
rect 4380 22820 4436 22876
rect 4436 22820 4440 22876
rect 4376 22816 4440 22820
rect 4456 22876 4520 22880
rect 4456 22820 4460 22876
rect 4460 22820 4516 22876
rect 4516 22820 4520 22876
rect 4456 22816 4520 22820
rect 34936 22876 35000 22880
rect 34936 22820 34940 22876
rect 34940 22820 34996 22876
rect 34996 22820 35000 22876
rect 34936 22816 35000 22820
rect 35016 22876 35080 22880
rect 35016 22820 35020 22876
rect 35020 22820 35076 22876
rect 35076 22820 35080 22876
rect 35016 22816 35080 22820
rect 35096 22876 35160 22880
rect 35096 22820 35100 22876
rect 35100 22820 35156 22876
rect 35156 22820 35160 22876
rect 35096 22816 35160 22820
rect 35176 22876 35240 22880
rect 35176 22820 35180 22876
rect 35180 22820 35236 22876
rect 35236 22820 35240 22876
rect 35176 22816 35240 22820
rect 19576 22332 19640 22336
rect 19576 22276 19580 22332
rect 19580 22276 19636 22332
rect 19636 22276 19640 22332
rect 19576 22272 19640 22276
rect 19656 22332 19720 22336
rect 19656 22276 19660 22332
rect 19660 22276 19716 22332
rect 19716 22276 19720 22332
rect 19656 22272 19720 22276
rect 19736 22332 19800 22336
rect 19736 22276 19740 22332
rect 19740 22276 19796 22332
rect 19796 22276 19800 22332
rect 19736 22272 19800 22276
rect 19816 22332 19880 22336
rect 19816 22276 19820 22332
rect 19820 22276 19876 22332
rect 19876 22276 19880 22332
rect 19816 22272 19880 22276
rect 4216 21788 4280 21792
rect 4216 21732 4220 21788
rect 4220 21732 4276 21788
rect 4276 21732 4280 21788
rect 4216 21728 4280 21732
rect 4296 21788 4360 21792
rect 4296 21732 4300 21788
rect 4300 21732 4356 21788
rect 4356 21732 4360 21788
rect 4296 21728 4360 21732
rect 4376 21788 4440 21792
rect 4376 21732 4380 21788
rect 4380 21732 4436 21788
rect 4436 21732 4440 21788
rect 4376 21728 4440 21732
rect 4456 21788 4520 21792
rect 4456 21732 4460 21788
rect 4460 21732 4516 21788
rect 4516 21732 4520 21788
rect 4456 21728 4520 21732
rect 34936 21788 35000 21792
rect 34936 21732 34940 21788
rect 34940 21732 34996 21788
rect 34996 21732 35000 21788
rect 34936 21728 35000 21732
rect 35016 21788 35080 21792
rect 35016 21732 35020 21788
rect 35020 21732 35076 21788
rect 35076 21732 35080 21788
rect 35016 21728 35080 21732
rect 35096 21788 35160 21792
rect 35096 21732 35100 21788
rect 35100 21732 35156 21788
rect 35156 21732 35160 21788
rect 35096 21728 35160 21732
rect 35176 21788 35240 21792
rect 35176 21732 35180 21788
rect 35180 21732 35236 21788
rect 35236 21732 35240 21788
rect 35176 21728 35240 21732
rect 19576 21244 19640 21248
rect 19576 21188 19580 21244
rect 19580 21188 19636 21244
rect 19636 21188 19640 21244
rect 19576 21184 19640 21188
rect 19656 21244 19720 21248
rect 19656 21188 19660 21244
rect 19660 21188 19716 21244
rect 19716 21188 19720 21244
rect 19656 21184 19720 21188
rect 19736 21244 19800 21248
rect 19736 21188 19740 21244
rect 19740 21188 19796 21244
rect 19796 21188 19800 21244
rect 19736 21184 19800 21188
rect 19816 21244 19880 21248
rect 19816 21188 19820 21244
rect 19820 21188 19876 21244
rect 19876 21188 19880 21244
rect 19816 21184 19880 21188
rect 4216 20700 4280 20704
rect 4216 20644 4220 20700
rect 4220 20644 4276 20700
rect 4276 20644 4280 20700
rect 4216 20640 4280 20644
rect 4296 20700 4360 20704
rect 4296 20644 4300 20700
rect 4300 20644 4356 20700
rect 4356 20644 4360 20700
rect 4296 20640 4360 20644
rect 4376 20700 4440 20704
rect 4376 20644 4380 20700
rect 4380 20644 4436 20700
rect 4436 20644 4440 20700
rect 4376 20640 4440 20644
rect 4456 20700 4520 20704
rect 4456 20644 4460 20700
rect 4460 20644 4516 20700
rect 4516 20644 4520 20700
rect 4456 20640 4520 20644
rect 34936 20700 35000 20704
rect 34936 20644 34940 20700
rect 34940 20644 34996 20700
rect 34996 20644 35000 20700
rect 34936 20640 35000 20644
rect 35016 20700 35080 20704
rect 35016 20644 35020 20700
rect 35020 20644 35076 20700
rect 35076 20644 35080 20700
rect 35016 20640 35080 20644
rect 35096 20700 35160 20704
rect 35096 20644 35100 20700
rect 35100 20644 35156 20700
rect 35156 20644 35160 20700
rect 35096 20640 35160 20644
rect 35176 20700 35240 20704
rect 35176 20644 35180 20700
rect 35180 20644 35236 20700
rect 35236 20644 35240 20700
rect 35176 20640 35240 20644
rect 37780 20300 37844 20364
rect 19576 20156 19640 20160
rect 19576 20100 19580 20156
rect 19580 20100 19636 20156
rect 19636 20100 19640 20156
rect 19576 20096 19640 20100
rect 19656 20156 19720 20160
rect 19656 20100 19660 20156
rect 19660 20100 19716 20156
rect 19716 20100 19720 20156
rect 19656 20096 19720 20100
rect 19736 20156 19800 20160
rect 19736 20100 19740 20156
rect 19740 20100 19796 20156
rect 19796 20100 19800 20156
rect 19736 20096 19800 20100
rect 19816 20156 19880 20160
rect 19816 20100 19820 20156
rect 19820 20100 19876 20156
rect 19876 20100 19880 20156
rect 19816 20096 19880 20100
rect 19380 19952 19444 19956
rect 19380 19896 19430 19952
rect 19430 19896 19444 19952
rect 19380 19892 19444 19896
rect 4216 19612 4280 19616
rect 4216 19556 4220 19612
rect 4220 19556 4276 19612
rect 4276 19556 4280 19612
rect 4216 19552 4280 19556
rect 4296 19612 4360 19616
rect 4296 19556 4300 19612
rect 4300 19556 4356 19612
rect 4356 19556 4360 19612
rect 4296 19552 4360 19556
rect 4376 19612 4440 19616
rect 4376 19556 4380 19612
rect 4380 19556 4436 19612
rect 4436 19556 4440 19612
rect 4376 19552 4440 19556
rect 4456 19612 4520 19616
rect 4456 19556 4460 19612
rect 4460 19556 4516 19612
rect 4516 19556 4520 19612
rect 4456 19552 4520 19556
rect 34936 19612 35000 19616
rect 34936 19556 34940 19612
rect 34940 19556 34996 19612
rect 34996 19556 35000 19612
rect 34936 19552 35000 19556
rect 35016 19612 35080 19616
rect 35016 19556 35020 19612
rect 35020 19556 35076 19612
rect 35076 19556 35080 19612
rect 35016 19552 35080 19556
rect 35096 19612 35160 19616
rect 35096 19556 35100 19612
rect 35100 19556 35156 19612
rect 35156 19556 35160 19612
rect 35096 19552 35160 19556
rect 35176 19612 35240 19616
rect 35176 19556 35180 19612
rect 35180 19556 35236 19612
rect 35236 19556 35240 19612
rect 35176 19552 35240 19556
rect 21404 19348 21468 19412
rect 28764 19272 28828 19276
rect 28764 19216 28814 19272
rect 28814 19216 28828 19272
rect 28764 19212 28828 19216
rect 19576 19068 19640 19072
rect 19576 19012 19580 19068
rect 19580 19012 19636 19068
rect 19636 19012 19640 19068
rect 19576 19008 19640 19012
rect 19656 19068 19720 19072
rect 19656 19012 19660 19068
rect 19660 19012 19716 19068
rect 19716 19012 19720 19068
rect 19656 19008 19720 19012
rect 19736 19068 19800 19072
rect 19736 19012 19740 19068
rect 19740 19012 19796 19068
rect 19796 19012 19800 19068
rect 19736 19008 19800 19012
rect 19816 19068 19880 19072
rect 19816 19012 19820 19068
rect 19820 19012 19876 19068
rect 19876 19012 19880 19068
rect 19816 19008 19880 19012
rect 4216 18524 4280 18528
rect 4216 18468 4220 18524
rect 4220 18468 4276 18524
rect 4276 18468 4280 18524
rect 4216 18464 4280 18468
rect 4296 18524 4360 18528
rect 4296 18468 4300 18524
rect 4300 18468 4356 18524
rect 4356 18468 4360 18524
rect 4296 18464 4360 18468
rect 4376 18524 4440 18528
rect 4376 18468 4380 18524
rect 4380 18468 4436 18524
rect 4436 18468 4440 18524
rect 4376 18464 4440 18468
rect 4456 18524 4520 18528
rect 4456 18468 4460 18524
rect 4460 18468 4516 18524
rect 4516 18468 4520 18524
rect 4456 18464 4520 18468
rect 34936 18524 35000 18528
rect 34936 18468 34940 18524
rect 34940 18468 34996 18524
rect 34996 18468 35000 18524
rect 34936 18464 35000 18468
rect 35016 18524 35080 18528
rect 35016 18468 35020 18524
rect 35020 18468 35076 18524
rect 35076 18468 35080 18524
rect 35016 18464 35080 18468
rect 35096 18524 35160 18528
rect 35096 18468 35100 18524
rect 35100 18468 35156 18524
rect 35156 18468 35160 18524
rect 35096 18464 35160 18468
rect 35176 18524 35240 18528
rect 35176 18468 35180 18524
rect 35180 18468 35236 18524
rect 35236 18468 35240 18524
rect 35176 18464 35240 18468
rect 19576 17980 19640 17984
rect 19576 17924 19580 17980
rect 19580 17924 19636 17980
rect 19636 17924 19640 17980
rect 19576 17920 19640 17924
rect 19656 17980 19720 17984
rect 19656 17924 19660 17980
rect 19660 17924 19716 17980
rect 19716 17924 19720 17980
rect 19656 17920 19720 17924
rect 19736 17980 19800 17984
rect 19736 17924 19740 17980
rect 19740 17924 19796 17980
rect 19796 17924 19800 17980
rect 19736 17920 19800 17924
rect 19816 17980 19880 17984
rect 19816 17924 19820 17980
rect 19820 17924 19876 17980
rect 19876 17924 19880 17980
rect 19816 17920 19880 17924
rect 4216 17436 4280 17440
rect 4216 17380 4220 17436
rect 4220 17380 4276 17436
rect 4276 17380 4280 17436
rect 4216 17376 4280 17380
rect 4296 17436 4360 17440
rect 4296 17380 4300 17436
rect 4300 17380 4356 17436
rect 4356 17380 4360 17436
rect 4296 17376 4360 17380
rect 4376 17436 4440 17440
rect 4376 17380 4380 17436
rect 4380 17380 4436 17436
rect 4436 17380 4440 17436
rect 4376 17376 4440 17380
rect 4456 17436 4520 17440
rect 4456 17380 4460 17436
rect 4460 17380 4516 17436
rect 4516 17380 4520 17436
rect 4456 17376 4520 17380
rect 34936 17436 35000 17440
rect 34936 17380 34940 17436
rect 34940 17380 34996 17436
rect 34996 17380 35000 17436
rect 34936 17376 35000 17380
rect 35016 17436 35080 17440
rect 35016 17380 35020 17436
rect 35020 17380 35076 17436
rect 35076 17380 35080 17436
rect 35016 17376 35080 17380
rect 35096 17436 35160 17440
rect 35096 17380 35100 17436
rect 35100 17380 35156 17436
rect 35156 17380 35160 17436
rect 35096 17376 35160 17380
rect 35176 17436 35240 17440
rect 35176 17380 35180 17436
rect 35180 17380 35236 17436
rect 35236 17380 35240 17436
rect 35176 17376 35240 17380
rect 19576 16892 19640 16896
rect 19576 16836 19580 16892
rect 19580 16836 19636 16892
rect 19636 16836 19640 16892
rect 19576 16832 19640 16836
rect 19656 16892 19720 16896
rect 19656 16836 19660 16892
rect 19660 16836 19716 16892
rect 19716 16836 19720 16892
rect 19656 16832 19720 16836
rect 19736 16892 19800 16896
rect 19736 16836 19740 16892
rect 19740 16836 19796 16892
rect 19796 16836 19800 16892
rect 19736 16832 19800 16836
rect 19816 16892 19880 16896
rect 19816 16836 19820 16892
rect 19820 16836 19876 16892
rect 19876 16836 19880 16892
rect 19816 16832 19880 16836
rect 4216 16348 4280 16352
rect 4216 16292 4220 16348
rect 4220 16292 4276 16348
rect 4276 16292 4280 16348
rect 4216 16288 4280 16292
rect 4296 16348 4360 16352
rect 4296 16292 4300 16348
rect 4300 16292 4356 16348
rect 4356 16292 4360 16348
rect 4296 16288 4360 16292
rect 4376 16348 4440 16352
rect 4376 16292 4380 16348
rect 4380 16292 4436 16348
rect 4436 16292 4440 16348
rect 4376 16288 4440 16292
rect 4456 16348 4520 16352
rect 4456 16292 4460 16348
rect 4460 16292 4516 16348
rect 4516 16292 4520 16348
rect 4456 16288 4520 16292
rect 34936 16348 35000 16352
rect 34936 16292 34940 16348
rect 34940 16292 34996 16348
rect 34996 16292 35000 16348
rect 34936 16288 35000 16292
rect 35016 16348 35080 16352
rect 35016 16292 35020 16348
rect 35020 16292 35076 16348
rect 35076 16292 35080 16348
rect 35016 16288 35080 16292
rect 35096 16348 35160 16352
rect 35096 16292 35100 16348
rect 35100 16292 35156 16348
rect 35156 16292 35160 16348
rect 35096 16288 35160 16292
rect 35176 16348 35240 16352
rect 35176 16292 35180 16348
rect 35180 16292 35236 16348
rect 35236 16292 35240 16348
rect 35176 16288 35240 16292
rect 19576 15804 19640 15808
rect 19576 15748 19580 15804
rect 19580 15748 19636 15804
rect 19636 15748 19640 15804
rect 19576 15744 19640 15748
rect 19656 15804 19720 15808
rect 19656 15748 19660 15804
rect 19660 15748 19716 15804
rect 19716 15748 19720 15804
rect 19656 15744 19720 15748
rect 19736 15804 19800 15808
rect 19736 15748 19740 15804
rect 19740 15748 19796 15804
rect 19796 15748 19800 15804
rect 19736 15744 19800 15748
rect 19816 15804 19880 15808
rect 19816 15748 19820 15804
rect 19820 15748 19876 15804
rect 19876 15748 19880 15804
rect 19816 15744 19880 15748
rect 4216 15260 4280 15264
rect 4216 15204 4220 15260
rect 4220 15204 4276 15260
rect 4276 15204 4280 15260
rect 4216 15200 4280 15204
rect 4296 15260 4360 15264
rect 4296 15204 4300 15260
rect 4300 15204 4356 15260
rect 4356 15204 4360 15260
rect 4296 15200 4360 15204
rect 4376 15260 4440 15264
rect 4376 15204 4380 15260
rect 4380 15204 4436 15260
rect 4436 15204 4440 15260
rect 4376 15200 4440 15204
rect 4456 15260 4520 15264
rect 4456 15204 4460 15260
rect 4460 15204 4516 15260
rect 4516 15204 4520 15260
rect 4456 15200 4520 15204
rect 34936 15260 35000 15264
rect 34936 15204 34940 15260
rect 34940 15204 34996 15260
rect 34996 15204 35000 15260
rect 34936 15200 35000 15204
rect 35016 15260 35080 15264
rect 35016 15204 35020 15260
rect 35020 15204 35076 15260
rect 35076 15204 35080 15260
rect 35016 15200 35080 15204
rect 35096 15260 35160 15264
rect 35096 15204 35100 15260
rect 35100 15204 35156 15260
rect 35156 15204 35160 15260
rect 35096 15200 35160 15204
rect 35176 15260 35240 15264
rect 35176 15204 35180 15260
rect 35180 15204 35236 15260
rect 35236 15204 35240 15260
rect 35176 15200 35240 15204
rect 19576 14716 19640 14720
rect 19576 14660 19580 14716
rect 19580 14660 19636 14716
rect 19636 14660 19640 14716
rect 19576 14656 19640 14660
rect 19656 14716 19720 14720
rect 19656 14660 19660 14716
rect 19660 14660 19716 14716
rect 19716 14660 19720 14716
rect 19656 14656 19720 14660
rect 19736 14716 19800 14720
rect 19736 14660 19740 14716
rect 19740 14660 19796 14716
rect 19796 14660 19800 14716
rect 19736 14656 19800 14660
rect 19816 14716 19880 14720
rect 19816 14660 19820 14716
rect 19820 14660 19876 14716
rect 19876 14660 19880 14716
rect 19816 14656 19880 14660
rect 28764 14452 28828 14516
rect 4216 14172 4280 14176
rect 4216 14116 4220 14172
rect 4220 14116 4276 14172
rect 4276 14116 4280 14172
rect 4216 14112 4280 14116
rect 4296 14172 4360 14176
rect 4296 14116 4300 14172
rect 4300 14116 4356 14172
rect 4356 14116 4360 14172
rect 4296 14112 4360 14116
rect 4376 14172 4440 14176
rect 4376 14116 4380 14172
rect 4380 14116 4436 14172
rect 4436 14116 4440 14172
rect 4376 14112 4440 14116
rect 4456 14172 4520 14176
rect 4456 14116 4460 14172
rect 4460 14116 4516 14172
rect 4516 14116 4520 14172
rect 4456 14112 4520 14116
rect 34936 14172 35000 14176
rect 34936 14116 34940 14172
rect 34940 14116 34996 14172
rect 34996 14116 35000 14172
rect 34936 14112 35000 14116
rect 35016 14172 35080 14176
rect 35016 14116 35020 14172
rect 35020 14116 35076 14172
rect 35076 14116 35080 14172
rect 35016 14112 35080 14116
rect 35096 14172 35160 14176
rect 35096 14116 35100 14172
rect 35100 14116 35156 14172
rect 35156 14116 35160 14172
rect 35096 14112 35160 14116
rect 35176 14172 35240 14176
rect 35176 14116 35180 14172
rect 35180 14116 35236 14172
rect 35236 14116 35240 14172
rect 35176 14112 35240 14116
rect 19576 13628 19640 13632
rect 19576 13572 19580 13628
rect 19580 13572 19636 13628
rect 19636 13572 19640 13628
rect 19576 13568 19640 13572
rect 19656 13628 19720 13632
rect 19656 13572 19660 13628
rect 19660 13572 19716 13628
rect 19716 13572 19720 13628
rect 19656 13568 19720 13572
rect 19736 13628 19800 13632
rect 19736 13572 19740 13628
rect 19740 13572 19796 13628
rect 19796 13572 19800 13628
rect 19736 13568 19800 13572
rect 19816 13628 19880 13632
rect 19816 13572 19820 13628
rect 19820 13572 19876 13628
rect 19876 13572 19880 13628
rect 19816 13568 19880 13572
rect 4216 13084 4280 13088
rect 4216 13028 4220 13084
rect 4220 13028 4276 13084
rect 4276 13028 4280 13084
rect 4216 13024 4280 13028
rect 4296 13084 4360 13088
rect 4296 13028 4300 13084
rect 4300 13028 4356 13084
rect 4356 13028 4360 13084
rect 4296 13024 4360 13028
rect 4376 13084 4440 13088
rect 4376 13028 4380 13084
rect 4380 13028 4436 13084
rect 4436 13028 4440 13084
rect 4376 13024 4440 13028
rect 4456 13084 4520 13088
rect 4456 13028 4460 13084
rect 4460 13028 4516 13084
rect 4516 13028 4520 13084
rect 4456 13024 4520 13028
rect 34936 13084 35000 13088
rect 34936 13028 34940 13084
rect 34940 13028 34996 13084
rect 34996 13028 35000 13084
rect 34936 13024 35000 13028
rect 35016 13084 35080 13088
rect 35016 13028 35020 13084
rect 35020 13028 35076 13084
rect 35076 13028 35080 13084
rect 35016 13024 35080 13028
rect 35096 13084 35160 13088
rect 35096 13028 35100 13084
rect 35100 13028 35156 13084
rect 35156 13028 35160 13084
rect 35096 13024 35160 13028
rect 35176 13084 35240 13088
rect 35176 13028 35180 13084
rect 35180 13028 35236 13084
rect 35236 13028 35240 13084
rect 35176 13024 35240 13028
rect 19576 12540 19640 12544
rect 19576 12484 19580 12540
rect 19580 12484 19636 12540
rect 19636 12484 19640 12540
rect 19576 12480 19640 12484
rect 19656 12540 19720 12544
rect 19656 12484 19660 12540
rect 19660 12484 19716 12540
rect 19716 12484 19720 12540
rect 19656 12480 19720 12484
rect 19736 12540 19800 12544
rect 19736 12484 19740 12540
rect 19740 12484 19796 12540
rect 19796 12484 19800 12540
rect 19736 12480 19800 12484
rect 19816 12540 19880 12544
rect 19816 12484 19820 12540
rect 19820 12484 19876 12540
rect 19876 12484 19880 12540
rect 19816 12480 19880 12484
rect 4216 11996 4280 12000
rect 4216 11940 4220 11996
rect 4220 11940 4276 11996
rect 4276 11940 4280 11996
rect 4216 11936 4280 11940
rect 4296 11996 4360 12000
rect 4296 11940 4300 11996
rect 4300 11940 4356 11996
rect 4356 11940 4360 11996
rect 4296 11936 4360 11940
rect 4376 11996 4440 12000
rect 4376 11940 4380 11996
rect 4380 11940 4436 11996
rect 4436 11940 4440 11996
rect 4376 11936 4440 11940
rect 4456 11996 4520 12000
rect 4456 11940 4460 11996
rect 4460 11940 4516 11996
rect 4516 11940 4520 11996
rect 4456 11936 4520 11940
rect 34936 11996 35000 12000
rect 34936 11940 34940 11996
rect 34940 11940 34996 11996
rect 34996 11940 35000 11996
rect 34936 11936 35000 11940
rect 35016 11996 35080 12000
rect 35016 11940 35020 11996
rect 35020 11940 35076 11996
rect 35076 11940 35080 11996
rect 35016 11936 35080 11940
rect 35096 11996 35160 12000
rect 35096 11940 35100 11996
rect 35100 11940 35156 11996
rect 35156 11940 35160 11996
rect 35096 11936 35160 11940
rect 35176 11996 35240 12000
rect 35176 11940 35180 11996
rect 35180 11940 35236 11996
rect 35236 11940 35240 11996
rect 35176 11936 35240 11940
rect 19576 11452 19640 11456
rect 19576 11396 19580 11452
rect 19580 11396 19636 11452
rect 19636 11396 19640 11452
rect 19576 11392 19640 11396
rect 19656 11452 19720 11456
rect 19656 11396 19660 11452
rect 19660 11396 19716 11452
rect 19716 11396 19720 11452
rect 19656 11392 19720 11396
rect 19736 11452 19800 11456
rect 19736 11396 19740 11452
rect 19740 11396 19796 11452
rect 19796 11396 19800 11452
rect 19736 11392 19800 11396
rect 19816 11452 19880 11456
rect 19816 11396 19820 11452
rect 19820 11396 19876 11452
rect 19876 11396 19880 11452
rect 19816 11392 19880 11396
rect 4216 10908 4280 10912
rect 4216 10852 4220 10908
rect 4220 10852 4276 10908
rect 4276 10852 4280 10908
rect 4216 10848 4280 10852
rect 4296 10908 4360 10912
rect 4296 10852 4300 10908
rect 4300 10852 4356 10908
rect 4356 10852 4360 10908
rect 4296 10848 4360 10852
rect 4376 10908 4440 10912
rect 4376 10852 4380 10908
rect 4380 10852 4436 10908
rect 4436 10852 4440 10908
rect 4376 10848 4440 10852
rect 4456 10908 4520 10912
rect 4456 10852 4460 10908
rect 4460 10852 4516 10908
rect 4516 10852 4520 10908
rect 4456 10848 4520 10852
rect 34936 10908 35000 10912
rect 34936 10852 34940 10908
rect 34940 10852 34996 10908
rect 34996 10852 35000 10908
rect 34936 10848 35000 10852
rect 35016 10908 35080 10912
rect 35016 10852 35020 10908
rect 35020 10852 35076 10908
rect 35076 10852 35080 10908
rect 35016 10848 35080 10852
rect 35096 10908 35160 10912
rect 35096 10852 35100 10908
rect 35100 10852 35156 10908
rect 35156 10852 35160 10908
rect 35096 10848 35160 10852
rect 35176 10908 35240 10912
rect 35176 10852 35180 10908
rect 35180 10852 35236 10908
rect 35236 10852 35240 10908
rect 35176 10848 35240 10852
rect 19576 10364 19640 10368
rect 19576 10308 19580 10364
rect 19580 10308 19636 10364
rect 19636 10308 19640 10364
rect 19576 10304 19640 10308
rect 19656 10364 19720 10368
rect 19656 10308 19660 10364
rect 19660 10308 19716 10364
rect 19716 10308 19720 10364
rect 19656 10304 19720 10308
rect 19736 10364 19800 10368
rect 19736 10308 19740 10364
rect 19740 10308 19796 10364
rect 19796 10308 19800 10364
rect 19736 10304 19800 10308
rect 19816 10364 19880 10368
rect 19816 10308 19820 10364
rect 19820 10308 19876 10364
rect 19876 10308 19880 10364
rect 19816 10304 19880 10308
rect 4216 9820 4280 9824
rect 4216 9764 4220 9820
rect 4220 9764 4276 9820
rect 4276 9764 4280 9820
rect 4216 9760 4280 9764
rect 4296 9820 4360 9824
rect 4296 9764 4300 9820
rect 4300 9764 4356 9820
rect 4356 9764 4360 9820
rect 4296 9760 4360 9764
rect 4376 9820 4440 9824
rect 4376 9764 4380 9820
rect 4380 9764 4436 9820
rect 4436 9764 4440 9820
rect 4376 9760 4440 9764
rect 4456 9820 4520 9824
rect 4456 9764 4460 9820
rect 4460 9764 4516 9820
rect 4516 9764 4520 9820
rect 4456 9760 4520 9764
rect 34936 9820 35000 9824
rect 34936 9764 34940 9820
rect 34940 9764 34996 9820
rect 34996 9764 35000 9820
rect 34936 9760 35000 9764
rect 35016 9820 35080 9824
rect 35016 9764 35020 9820
rect 35020 9764 35076 9820
rect 35076 9764 35080 9820
rect 35016 9760 35080 9764
rect 35096 9820 35160 9824
rect 35096 9764 35100 9820
rect 35100 9764 35156 9820
rect 35156 9764 35160 9820
rect 35096 9760 35160 9764
rect 35176 9820 35240 9824
rect 35176 9764 35180 9820
rect 35180 9764 35236 9820
rect 35236 9764 35240 9820
rect 35176 9760 35240 9764
rect 19576 9276 19640 9280
rect 19576 9220 19580 9276
rect 19580 9220 19636 9276
rect 19636 9220 19640 9276
rect 19576 9216 19640 9220
rect 19656 9276 19720 9280
rect 19656 9220 19660 9276
rect 19660 9220 19716 9276
rect 19716 9220 19720 9276
rect 19656 9216 19720 9220
rect 19736 9276 19800 9280
rect 19736 9220 19740 9276
rect 19740 9220 19796 9276
rect 19796 9220 19800 9276
rect 19736 9216 19800 9220
rect 19816 9276 19880 9280
rect 19816 9220 19820 9276
rect 19820 9220 19876 9276
rect 19876 9220 19880 9276
rect 19816 9216 19880 9220
rect 4216 8732 4280 8736
rect 4216 8676 4220 8732
rect 4220 8676 4276 8732
rect 4276 8676 4280 8732
rect 4216 8672 4280 8676
rect 4296 8732 4360 8736
rect 4296 8676 4300 8732
rect 4300 8676 4356 8732
rect 4356 8676 4360 8732
rect 4296 8672 4360 8676
rect 4376 8732 4440 8736
rect 4376 8676 4380 8732
rect 4380 8676 4436 8732
rect 4436 8676 4440 8732
rect 4376 8672 4440 8676
rect 4456 8732 4520 8736
rect 4456 8676 4460 8732
rect 4460 8676 4516 8732
rect 4516 8676 4520 8732
rect 4456 8672 4520 8676
rect 34936 8732 35000 8736
rect 34936 8676 34940 8732
rect 34940 8676 34996 8732
rect 34996 8676 35000 8732
rect 34936 8672 35000 8676
rect 35016 8732 35080 8736
rect 35016 8676 35020 8732
rect 35020 8676 35076 8732
rect 35076 8676 35080 8732
rect 35016 8672 35080 8676
rect 35096 8732 35160 8736
rect 35096 8676 35100 8732
rect 35100 8676 35156 8732
rect 35156 8676 35160 8732
rect 35096 8672 35160 8676
rect 35176 8732 35240 8736
rect 35176 8676 35180 8732
rect 35180 8676 35236 8732
rect 35236 8676 35240 8732
rect 35176 8672 35240 8676
rect 19576 8188 19640 8192
rect 19576 8132 19580 8188
rect 19580 8132 19636 8188
rect 19636 8132 19640 8188
rect 19576 8128 19640 8132
rect 19656 8188 19720 8192
rect 19656 8132 19660 8188
rect 19660 8132 19716 8188
rect 19716 8132 19720 8188
rect 19656 8128 19720 8132
rect 19736 8188 19800 8192
rect 19736 8132 19740 8188
rect 19740 8132 19796 8188
rect 19796 8132 19800 8188
rect 19736 8128 19800 8132
rect 19816 8188 19880 8192
rect 19816 8132 19820 8188
rect 19820 8132 19876 8188
rect 19876 8132 19880 8188
rect 19816 8128 19880 8132
rect 4216 7644 4280 7648
rect 4216 7588 4220 7644
rect 4220 7588 4276 7644
rect 4276 7588 4280 7644
rect 4216 7584 4280 7588
rect 4296 7644 4360 7648
rect 4296 7588 4300 7644
rect 4300 7588 4356 7644
rect 4356 7588 4360 7644
rect 4296 7584 4360 7588
rect 4376 7644 4440 7648
rect 4376 7588 4380 7644
rect 4380 7588 4436 7644
rect 4436 7588 4440 7644
rect 4376 7584 4440 7588
rect 4456 7644 4520 7648
rect 4456 7588 4460 7644
rect 4460 7588 4516 7644
rect 4516 7588 4520 7644
rect 4456 7584 4520 7588
rect 34936 7644 35000 7648
rect 34936 7588 34940 7644
rect 34940 7588 34996 7644
rect 34996 7588 35000 7644
rect 34936 7584 35000 7588
rect 35016 7644 35080 7648
rect 35016 7588 35020 7644
rect 35020 7588 35076 7644
rect 35076 7588 35080 7644
rect 35016 7584 35080 7588
rect 35096 7644 35160 7648
rect 35096 7588 35100 7644
rect 35100 7588 35156 7644
rect 35156 7588 35160 7644
rect 35096 7584 35160 7588
rect 35176 7644 35240 7648
rect 35176 7588 35180 7644
rect 35180 7588 35236 7644
rect 35236 7588 35240 7644
rect 35176 7584 35240 7588
rect 21404 7244 21468 7308
rect 19576 7100 19640 7104
rect 19576 7044 19580 7100
rect 19580 7044 19636 7100
rect 19636 7044 19640 7100
rect 19576 7040 19640 7044
rect 19656 7100 19720 7104
rect 19656 7044 19660 7100
rect 19660 7044 19716 7100
rect 19716 7044 19720 7100
rect 19656 7040 19720 7044
rect 19736 7100 19800 7104
rect 19736 7044 19740 7100
rect 19740 7044 19796 7100
rect 19796 7044 19800 7100
rect 19736 7040 19800 7044
rect 19816 7100 19880 7104
rect 19816 7044 19820 7100
rect 19820 7044 19876 7100
rect 19876 7044 19880 7100
rect 19816 7040 19880 7044
rect 19380 6836 19444 6900
rect 4216 6556 4280 6560
rect 4216 6500 4220 6556
rect 4220 6500 4276 6556
rect 4276 6500 4280 6556
rect 4216 6496 4280 6500
rect 4296 6556 4360 6560
rect 4296 6500 4300 6556
rect 4300 6500 4356 6556
rect 4356 6500 4360 6556
rect 4296 6496 4360 6500
rect 4376 6556 4440 6560
rect 4376 6500 4380 6556
rect 4380 6500 4436 6556
rect 4436 6500 4440 6556
rect 4376 6496 4440 6500
rect 4456 6556 4520 6560
rect 4456 6500 4460 6556
rect 4460 6500 4516 6556
rect 4516 6500 4520 6556
rect 4456 6496 4520 6500
rect 34936 6556 35000 6560
rect 34936 6500 34940 6556
rect 34940 6500 34996 6556
rect 34996 6500 35000 6556
rect 34936 6496 35000 6500
rect 35016 6556 35080 6560
rect 35016 6500 35020 6556
rect 35020 6500 35076 6556
rect 35076 6500 35080 6556
rect 35016 6496 35080 6500
rect 35096 6556 35160 6560
rect 35096 6500 35100 6556
rect 35100 6500 35156 6556
rect 35156 6500 35160 6556
rect 35096 6496 35160 6500
rect 35176 6556 35240 6560
rect 35176 6500 35180 6556
rect 35180 6500 35236 6556
rect 35236 6500 35240 6556
rect 35176 6496 35240 6500
rect 19576 6012 19640 6016
rect 19576 5956 19580 6012
rect 19580 5956 19636 6012
rect 19636 5956 19640 6012
rect 19576 5952 19640 5956
rect 19656 6012 19720 6016
rect 19656 5956 19660 6012
rect 19660 5956 19716 6012
rect 19716 5956 19720 6012
rect 19656 5952 19720 5956
rect 19736 6012 19800 6016
rect 19736 5956 19740 6012
rect 19740 5956 19796 6012
rect 19796 5956 19800 6012
rect 19736 5952 19800 5956
rect 19816 6012 19880 6016
rect 19816 5956 19820 6012
rect 19820 5956 19876 6012
rect 19876 5956 19880 6012
rect 19816 5952 19880 5956
rect 4216 5468 4280 5472
rect 4216 5412 4220 5468
rect 4220 5412 4276 5468
rect 4276 5412 4280 5468
rect 4216 5408 4280 5412
rect 4296 5468 4360 5472
rect 4296 5412 4300 5468
rect 4300 5412 4356 5468
rect 4356 5412 4360 5468
rect 4296 5408 4360 5412
rect 4376 5468 4440 5472
rect 4376 5412 4380 5468
rect 4380 5412 4436 5468
rect 4436 5412 4440 5468
rect 4376 5408 4440 5412
rect 4456 5468 4520 5472
rect 4456 5412 4460 5468
rect 4460 5412 4516 5468
rect 4516 5412 4520 5468
rect 4456 5408 4520 5412
rect 34936 5468 35000 5472
rect 34936 5412 34940 5468
rect 34940 5412 34996 5468
rect 34996 5412 35000 5468
rect 34936 5408 35000 5412
rect 35016 5468 35080 5472
rect 35016 5412 35020 5468
rect 35020 5412 35076 5468
rect 35076 5412 35080 5468
rect 35016 5408 35080 5412
rect 35096 5468 35160 5472
rect 35096 5412 35100 5468
rect 35100 5412 35156 5468
rect 35156 5412 35160 5468
rect 35096 5408 35160 5412
rect 35176 5468 35240 5472
rect 35176 5412 35180 5468
rect 35180 5412 35236 5468
rect 35236 5412 35240 5468
rect 35176 5408 35240 5412
rect 19576 4924 19640 4928
rect 19576 4868 19580 4924
rect 19580 4868 19636 4924
rect 19636 4868 19640 4924
rect 19576 4864 19640 4868
rect 19656 4924 19720 4928
rect 19656 4868 19660 4924
rect 19660 4868 19716 4924
rect 19716 4868 19720 4924
rect 19656 4864 19720 4868
rect 19736 4924 19800 4928
rect 19736 4868 19740 4924
rect 19740 4868 19796 4924
rect 19796 4868 19800 4924
rect 19736 4864 19800 4868
rect 19816 4924 19880 4928
rect 19816 4868 19820 4924
rect 19820 4868 19876 4924
rect 19876 4868 19880 4924
rect 19816 4864 19880 4868
rect 4216 4380 4280 4384
rect 4216 4324 4220 4380
rect 4220 4324 4276 4380
rect 4276 4324 4280 4380
rect 4216 4320 4280 4324
rect 4296 4380 4360 4384
rect 4296 4324 4300 4380
rect 4300 4324 4356 4380
rect 4356 4324 4360 4380
rect 4296 4320 4360 4324
rect 4376 4380 4440 4384
rect 4376 4324 4380 4380
rect 4380 4324 4436 4380
rect 4436 4324 4440 4380
rect 4376 4320 4440 4324
rect 4456 4380 4520 4384
rect 4456 4324 4460 4380
rect 4460 4324 4516 4380
rect 4516 4324 4520 4380
rect 4456 4320 4520 4324
rect 34936 4380 35000 4384
rect 34936 4324 34940 4380
rect 34940 4324 34996 4380
rect 34996 4324 35000 4380
rect 34936 4320 35000 4324
rect 35016 4380 35080 4384
rect 35016 4324 35020 4380
rect 35020 4324 35076 4380
rect 35076 4324 35080 4380
rect 35016 4320 35080 4324
rect 35096 4380 35160 4384
rect 35096 4324 35100 4380
rect 35100 4324 35156 4380
rect 35156 4324 35160 4380
rect 35096 4320 35160 4324
rect 35176 4380 35240 4384
rect 35176 4324 35180 4380
rect 35180 4324 35236 4380
rect 35236 4324 35240 4380
rect 35176 4320 35240 4324
rect 19576 3836 19640 3840
rect 19576 3780 19580 3836
rect 19580 3780 19636 3836
rect 19636 3780 19640 3836
rect 19576 3776 19640 3780
rect 19656 3836 19720 3840
rect 19656 3780 19660 3836
rect 19660 3780 19716 3836
rect 19716 3780 19720 3836
rect 19656 3776 19720 3780
rect 19736 3836 19800 3840
rect 19736 3780 19740 3836
rect 19740 3780 19796 3836
rect 19796 3780 19800 3836
rect 19736 3776 19800 3780
rect 19816 3836 19880 3840
rect 19816 3780 19820 3836
rect 19820 3780 19876 3836
rect 19876 3780 19880 3836
rect 19816 3776 19880 3780
rect 27108 3572 27172 3636
rect 4216 3292 4280 3296
rect 4216 3236 4220 3292
rect 4220 3236 4276 3292
rect 4276 3236 4280 3292
rect 4216 3232 4280 3236
rect 4296 3292 4360 3296
rect 4296 3236 4300 3292
rect 4300 3236 4356 3292
rect 4356 3236 4360 3292
rect 4296 3232 4360 3236
rect 4376 3292 4440 3296
rect 4376 3236 4380 3292
rect 4380 3236 4436 3292
rect 4436 3236 4440 3292
rect 4376 3232 4440 3236
rect 4456 3292 4520 3296
rect 4456 3236 4460 3292
rect 4460 3236 4516 3292
rect 4516 3236 4520 3292
rect 4456 3232 4520 3236
rect 34936 3292 35000 3296
rect 34936 3236 34940 3292
rect 34940 3236 34996 3292
rect 34996 3236 35000 3292
rect 34936 3232 35000 3236
rect 35016 3292 35080 3296
rect 35016 3236 35020 3292
rect 35020 3236 35076 3292
rect 35076 3236 35080 3292
rect 35016 3232 35080 3236
rect 35096 3292 35160 3296
rect 35096 3236 35100 3292
rect 35100 3236 35156 3292
rect 35156 3236 35160 3292
rect 35096 3232 35160 3236
rect 35176 3292 35240 3296
rect 35176 3236 35180 3292
rect 35180 3236 35236 3292
rect 35236 3236 35240 3292
rect 35176 3232 35240 3236
rect 19576 2748 19640 2752
rect 19576 2692 19580 2748
rect 19580 2692 19636 2748
rect 19636 2692 19640 2748
rect 19576 2688 19640 2692
rect 19656 2748 19720 2752
rect 19656 2692 19660 2748
rect 19660 2692 19716 2748
rect 19716 2692 19720 2748
rect 19656 2688 19720 2692
rect 19736 2748 19800 2752
rect 19736 2692 19740 2748
rect 19740 2692 19796 2748
rect 19796 2692 19800 2748
rect 19736 2688 19800 2692
rect 19816 2748 19880 2752
rect 19816 2692 19820 2748
rect 19820 2692 19876 2748
rect 19876 2692 19880 2748
rect 19816 2688 19880 2692
rect 4216 2204 4280 2208
rect 4216 2148 4220 2204
rect 4220 2148 4276 2204
rect 4276 2148 4280 2204
rect 4216 2144 4280 2148
rect 4296 2204 4360 2208
rect 4296 2148 4300 2204
rect 4300 2148 4356 2204
rect 4356 2148 4360 2204
rect 4296 2144 4360 2148
rect 4376 2204 4440 2208
rect 4376 2148 4380 2204
rect 4380 2148 4436 2204
rect 4436 2148 4440 2204
rect 4376 2144 4440 2148
rect 4456 2204 4520 2208
rect 4456 2148 4460 2204
rect 4460 2148 4516 2204
rect 4516 2148 4520 2204
rect 4456 2144 4520 2148
rect 34936 2204 35000 2208
rect 34936 2148 34940 2204
rect 34940 2148 34996 2204
rect 34996 2148 35000 2204
rect 34936 2144 35000 2148
rect 35016 2204 35080 2208
rect 35016 2148 35020 2204
rect 35020 2148 35076 2204
rect 35076 2148 35080 2204
rect 35016 2144 35080 2148
rect 35096 2204 35160 2208
rect 35096 2148 35100 2204
rect 35100 2148 35156 2204
rect 35156 2148 35160 2204
rect 35096 2144 35160 2148
rect 35176 2204 35240 2208
rect 35176 2148 35180 2204
rect 35180 2148 35236 2204
rect 35236 2148 35240 2204
rect 35176 2144 35240 2148
<< metal4 >>
rect 4208 38112 4528 38672
rect 19568 38656 19888 38672
rect 4208 38048 4216 38112
rect 4280 38048 4296 38112
rect 4360 38048 4376 38112
rect 4440 38048 4456 38112
rect 4520 38048 4528 38112
rect 4208 37024 4528 38048
rect 4208 36960 4216 37024
rect 4280 36960 4296 37024
rect 4360 36960 4376 37024
rect 4440 36960 4456 37024
rect 4520 36960 4528 37024
rect 4208 35936 4528 36960
rect 4208 35872 4216 35936
rect 4280 35872 4296 35936
rect 4360 35872 4376 35936
rect 4440 35872 4456 35936
rect 4520 35872 4528 35936
rect 4208 34848 4528 35872
rect 4208 34784 4216 34848
rect 4280 34784 4296 34848
rect 4360 34784 4376 34848
rect 4440 34784 4456 34848
rect 4520 34784 4528 34848
rect 4208 33760 4528 34784
rect 4208 33696 4216 33760
rect 4280 33696 4296 33760
rect 4360 33696 4376 33760
rect 4440 33696 4456 33760
rect 4520 33696 4528 33760
rect 4208 32672 4528 33696
rect 4208 32608 4216 32672
rect 4280 32608 4296 32672
rect 4360 32608 4376 32672
rect 4440 32608 4456 32672
rect 4520 32608 4528 32672
rect 4208 31584 4528 32608
rect 4208 31520 4216 31584
rect 4280 31520 4296 31584
rect 4360 31520 4376 31584
rect 4440 31520 4456 31584
rect 4520 31520 4528 31584
rect 4208 30496 4528 31520
rect 4208 30432 4216 30496
rect 4280 30432 4296 30496
rect 4360 30432 4376 30496
rect 4440 30432 4456 30496
rect 4520 30432 4528 30496
rect 4208 29408 4528 30432
rect 4208 29344 4216 29408
rect 4280 29344 4296 29408
rect 4360 29344 4376 29408
rect 4440 29344 4456 29408
rect 4520 29344 4528 29408
rect 4208 28320 4528 29344
rect 4208 28256 4216 28320
rect 4280 28256 4296 28320
rect 4360 28256 4376 28320
rect 4440 28256 4456 28320
rect 4520 28256 4528 28320
rect 4208 27232 4528 28256
rect 4208 27168 4216 27232
rect 4280 27168 4296 27232
rect 4360 27168 4376 27232
rect 4440 27168 4456 27232
rect 4520 27168 4528 27232
rect 4208 26144 4528 27168
rect 4208 26080 4216 26144
rect 4280 26080 4296 26144
rect 4360 26080 4376 26144
rect 4440 26080 4456 26144
rect 4520 26080 4528 26144
rect 4208 25056 4528 26080
rect 4208 24992 4216 25056
rect 4280 24992 4296 25056
rect 4360 24992 4376 25056
rect 4440 24992 4456 25056
rect 4520 24992 4528 25056
rect 4208 23968 4528 24992
rect 4208 23904 4216 23968
rect 4280 23904 4296 23968
rect 4360 23904 4376 23968
rect 4440 23904 4456 23968
rect 4520 23904 4528 23968
rect 4208 22880 4528 23904
rect 4208 22816 4216 22880
rect 4280 22816 4296 22880
rect 4360 22816 4376 22880
rect 4440 22816 4456 22880
rect 4520 22816 4528 22880
rect 4208 21792 4528 22816
rect 4208 21728 4216 21792
rect 4280 21728 4296 21792
rect 4360 21728 4376 21792
rect 4440 21728 4456 21792
rect 4520 21728 4528 21792
rect 4208 20704 4528 21728
rect 4208 20640 4216 20704
rect 4280 20640 4296 20704
rect 4360 20640 4376 20704
rect 4440 20640 4456 20704
rect 4520 20640 4528 20704
rect 4208 19616 4528 20640
rect 4208 19552 4216 19616
rect 4280 19552 4296 19616
rect 4360 19552 4376 19616
rect 4440 19552 4456 19616
rect 4520 19552 4528 19616
rect 4208 18528 4528 19552
rect 4208 18464 4216 18528
rect 4280 18464 4296 18528
rect 4360 18464 4376 18528
rect 4440 18464 4456 18528
rect 4520 18464 4528 18528
rect 4208 17440 4528 18464
rect 4208 17376 4216 17440
rect 4280 17376 4296 17440
rect 4360 17376 4376 17440
rect 4440 17376 4456 17440
rect 4520 17376 4528 17440
rect 4208 16352 4528 17376
rect 4208 16288 4216 16352
rect 4280 16288 4296 16352
rect 4360 16288 4376 16352
rect 4440 16288 4456 16352
rect 4520 16288 4528 16352
rect 4208 15264 4528 16288
rect 4208 15200 4216 15264
rect 4280 15200 4296 15264
rect 4360 15200 4376 15264
rect 4440 15200 4456 15264
rect 4520 15200 4528 15264
rect 4208 14176 4528 15200
rect 4208 14112 4216 14176
rect 4280 14112 4296 14176
rect 4360 14112 4376 14176
rect 4440 14112 4456 14176
rect 4520 14112 4528 14176
rect 4208 13088 4528 14112
rect 4208 13024 4216 13088
rect 4280 13024 4296 13088
rect 4360 13024 4376 13088
rect 4440 13024 4456 13088
rect 4520 13024 4528 13088
rect 4208 12000 4528 13024
rect 4208 11936 4216 12000
rect 4280 11936 4296 12000
rect 4360 11936 4376 12000
rect 4440 11936 4456 12000
rect 4520 11936 4528 12000
rect 4208 10912 4528 11936
rect 4208 10848 4216 10912
rect 4280 10848 4296 10912
rect 4360 10848 4376 10912
rect 4440 10848 4456 10912
rect 4520 10848 4528 10912
rect 4208 9824 4528 10848
rect 4208 9760 4216 9824
rect 4280 9760 4296 9824
rect 4360 9760 4376 9824
rect 4440 9760 4456 9824
rect 4520 9760 4528 9824
rect 4208 8736 4528 9760
rect 4208 8672 4216 8736
rect 4280 8672 4296 8736
rect 4360 8672 4376 8736
rect 4440 8672 4456 8736
rect 4520 8672 4528 8736
rect 4208 7648 4528 8672
rect 4208 7584 4216 7648
rect 4280 7584 4296 7648
rect 4360 7584 4376 7648
rect 4440 7584 4456 7648
rect 4520 7584 4528 7648
rect 4208 6560 4528 7584
rect 4208 6496 4216 6560
rect 4280 6496 4296 6560
rect 4360 6496 4376 6560
rect 4440 6496 4456 6560
rect 4520 6496 4528 6560
rect 4208 5472 4528 6496
rect 4208 5408 4216 5472
rect 4280 5408 4296 5472
rect 4360 5408 4376 5472
rect 4440 5408 4456 5472
rect 4520 5408 4528 5472
rect 4208 4384 4528 5408
rect 4208 4320 4216 4384
rect 4280 4320 4296 4384
rect 4360 4320 4376 4384
rect 4440 4320 4456 4384
rect 4520 4320 4528 4384
rect 4208 3296 4528 4320
rect 4208 3232 4216 3296
rect 4280 3232 4296 3296
rect 4360 3232 4376 3296
rect 4440 3232 4456 3296
rect 4520 3232 4528 3296
rect 4208 2208 4528 3232
rect 4208 2144 4216 2208
rect 4280 2144 4296 2208
rect 4360 2144 4376 2208
rect 4440 2144 4456 2208
rect 4520 2144 4528 2208
rect 4868 2176 5188 38624
rect 5528 2176 5848 38624
rect 6188 2176 6508 38624
rect 19568 38592 19576 38656
rect 19640 38592 19656 38656
rect 19720 38592 19736 38656
rect 19800 38592 19816 38656
rect 19880 38592 19888 38656
rect 19568 37568 19888 38592
rect 19568 37504 19576 37568
rect 19640 37504 19656 37568
rect 19720 37504 19736 37568
rect 19800 37504 19816 37568
rect 19880 37504 19888 37568
rect 19568 36480 19888 37504
rect 19568 36416 19576 36480
rect 19640 36416 19656 36480
rect 19720 36416 19736 36480
rect 19800 36416 19816 36480
rect 19880 36416 19888 36480
rect 19568 35392 19888 36416
rect 19568 35328 19576 35392
rect 19640 35328 19656 35392
rect 19720 35328 19736 35392
rect 19800 35328 19816 35392
rect 19880 35328 19888 35392
rect 19568 34304 19888 35328
rect 19568 34240 19576 34304
rect 19640 34240 19656 34304
rect 19720 34240 19736 34304
rect 19800 34240 19816 34304
rect 19880 34240 19888 34304
rect 19568 33216 19888 34240
rect 19568 33152 19576 33216
rect 19640 33152 19656 33216
rect 19720 33152 19736 33216
rect 19800 33152 19816 33216
rect 19880 33152 19888 33216
rect 19568 32128 19888 33152
rect 19568 32064 19576 32128
rect 19640 32064 19656 32128
rect 19720 32064 19736 32128
rect 19800 32064 19816 32128
rect 19880 32064 19888 32128
rect 19568 31040 19888 32064
rect 19568 30976 19576 31040
rect 19640 30976 19656 31040
rect 19720 30976 19736 31040
rect 19800 30976 19816 31040
rect 19880 30976 19888 31040
rect 19568 29952 19888 30976
rect 19568 29888 19576 29952
rect 19640 29888 19656 29952
rect 19720 29888 19736 29952
rect 19800 29888 19816 29952
rect 19880 29888 19888 29952
rect 19379 28932 19445 28933
rect 19379 28868 19380 28932
rect 19444 28868 19445 28932
rect 19379 28867 19445 28868
rect 19382 23357 19442 28867
rect 19568 28864 19888 29888
rect 19568 28800 19576 28864
rect 19640 28800 19656 28864
rect 19720 28800 19736 28864
rect 19800 28800 19816 28864
rect 19880 28800 19888 28864
rect 19568 27776 19888 28800
rect 19568 27712 19576 27776
rect 19640 27712 19656 27776
rect 19720 27712 19736 27776
rect 19800 27712 19816 27776
rect 19880 27712 19888 27776
rect 19568 26688 19888 27712
rect 19568 26624 19576 26688
rect 19640 26624 19656 26688
rect 19720 26624 19736 26688
rect 19800 26624 19816 26688
rect 19880 26624 19888 26688
rect 19568 25600 19888 26624
rect 19568 25536 19576 25600
rect 19640 25536 19656 25600
rect 19720 25536 19736 25600
rect 19800 25536 19816 25600
rect 19880 25536 19888 25600
rect 19568 24512 19888 25536
rect 19568 24448 19576 24512
rect 19640 24448 19656 24512
rect 19720 24448 19736 24512
rect 19800 24448 19816 24512
rect 19880 24448 19888 24512
rect 19568 23424 19888 24448
rect 19568 23360 19576 23424
rect 19640 23360 19656 23424
rect 19720 23360 19736 23424
rect 19800 23360 19816 23424
rect 19880 23360 19888 23424
rect 19379 23356 19445 23357
rect 19379 23292 19380 23356
rect 19444 23292 19445 23356
rect 19379 23291 19445 23292
rect 19568 22336 19888 23360
rect 19568 22272 19576 22336
rect 19640 22272 19656 22336
rect 19720 22272 19736 22336
rect 19800 22272 19816 22336
rect 19880 22272 19888 22336
rect 19568 21248 19888 22272
rect 19568 21184 19576 21248
rect 19640 21184 19656 21248
rect 19720 21184 19736 21248
rect 19800 21184 19816 21248
rect 19880 21184 19888 21248
rect 19568 20160 19888 21184
rect 19568 20096 19576 20160
rect 19640 20096 19656 20160
rect 19720 20096 19736 20160
rect 19800 20096 19816 20160
rect 19880 20096 19888 20160
rect 19379 19956 19445 19957
rect 19379 19892 19380 19956
rect 19444 19892 19445 19956
rect 19379 19891 19445 19892
rect 19382 6901 19442 19891
rect 19568 19072 19888 20096
rect 19568 19008 19576 19072
rect 19640 19008 19656 19072
rect 19720 19008 19736 19072
rect 19800 19008 19816 19072
rect 19880 19008 19888 19072
rect 19568 17984 19888 19008
rect 19568 17920 19576 17984
rect 19640 17920 19656 17984
rect 19720 17920 19736 17984
rect 19800 17920 19816 17984
rect 19880 17920 19888 17984
rect 19568 16896 19888 17920
rect 19568 16832 19576 16896
rect 19640 16832 19656 16896
rect 19720 16832 19736 16896
rect 19800 16832 19816 16896
rect 19880 16832 19888 16896
rect 19568 15808 19888 16832
rect 19568 15744 19576 15808
rect 19640 15744 19656 15808
rect 19720 15744 19736 15808
rect 19800 15744 19816 15808
rect 19880 15744 19888 15808
rect 19568 14720 19888 15744
rect 19568 14656 19576 14720
rect 19640 14656 19656 14720
rect 19720 14656 19736 14720
rect 19800 14656 19816 14720
rect 19880 14656 19888 14720
rect 19568 13632 19888 14656
rect 19568 13568 19576 13632
rect 19640 13568 19656 13632
rect 19720 13568 19736 13632
rect 19800 13568 19816 13632
rect 19880 13568 19888 13632
rect 19568 12544 19888 13568
rect 19568 12480 19576 12544
rect 19640 12480 19656 12544
rect 19720 12480 19736 12544
rect 19800 12480 19816 12544
rect 19880 12480 19888 12544
rect 19568 11456 19888 12480
rect 19568 11392 19576 11456
rect 19640 11392 19656 11456
rect 19720 11392 19736 11456
rect 19800 11392 19816 11456
rect 19880 11392 19888 11456
rect 19568 10368 19888 11392
rect 19568 10304 19576 10368
rect 19640 10304 19656 10368
rect 19720 10304 19736 10368
rect 19800 10304 19816 10368
rect 19880 10304 19888 10368
rect 19568 9280 19888 10304
rect 19568 9216 19576 9280
rect 19640 9216 19656 9280
rect 19720 9216 19736 9280
rect 19800 9216 19816 9280
rect 19880 9216 19888 9280
rect 19568 8192 19888 9216
rect 19568 8128 19576 8192
rect 19640 8128 19656 8192
rect 19720 8128 19736 8192
rect 19800 8128 19816 8192
rect 19880 8128 19888 8192
rect 19568 7104 19888 8128
rect 19568 7040 19576 7104
rect 19640 7040 19656 7104
rect 19720 7040 19736 7104
rect 19800 7040 19816 7104
rect 19880 7040 19888 7104
rect 19379 6900 19445 6901
rect 19379 6836 19380 6900
rect 19444 6836 19445 6900
rect 19379 6835 19445 6836
rect 19568 6016 19888 7040
rect 19568 5952 19576 6016
rect 19640 5952 19656 6016
rect 19720 5952 19736 6016
rect 19800 5952 19816 6016
rect 19880 5952 19888 6016
rect 19568 4928 19888 5952
rect 19568 4864 19576 4928
rect 19640 4864 19656 4928
rect 19720 4864 19736 4928
rect 19800 4864 19816 4928
rect 19880 4864 19888 4928
rect 19568 3840 19888 4864
rect 19568 3776 19576 3840
rect 19640 3776 19656 3840
rect 19720 3776 19736 3840
rect 19800 3776 19816 3840
rect 19880 3776 19888 3840
rect 19568 2752 19888 3776
rect 19568 2688 19576 2752
rect 19640 2688 19656 2752
rect 19720 2688 19736 2752
rect 19800 2688 19816 2752
rect 19880 2688 19888 2752
rect 4208 2128 4528 2144
rect 19568 2128 19888 2688
rect 20228 2176 20548 38624
rect 20888 2176 21208 38624
rect 21403 19412 21469 19413
rect 21403 19348 21404 19412
rect 21468 19348 21469 19412
rect 21403 19347 21469 19348
rect 21406 7309 21466 19347
rect 21403 7308 21469 7309
rect 21403 7244 21404 7308
rect 21468 7244 21469 7308
rect 21403 7243 21469 7244
rect 21548 2176 21868 38624
rect 34928 38112 35248 38672
rect 34928 38048 34936 38112
rect 35000 38048 35016 38112
rect 35080 38048 35096 38112
rect 35160 38048 35176 38112
rect 35240 38048 35248 38112
rect 34928 37024 35248 38048
rect 34928 36960 34936 37024
rect 35000 36960 35016 37024
rect 35080 36960 35096 37024
rect 35160 36960 35176 37024
rect 35240 36960 35248 37024
rect 34928 35936 35248 36960
rect 34928 35872 34936 35936
rect 35000 35872 35016 35936
rect 35080 35872 35096 35936
rect 35160 35872 35176 35936
rect 35240 35872 35248 35936
rect 34928 34848 35248 35872
rect 34928 34784 34936 34848
rect 35000 34784 35016 34848
rect 35080 34784 35096 34848
rect 35160 34784 35176 34848
rect 35240 34784 35248 34848
rect 34928 33760 35248 34784
rect 34928 33696 34936 33760
rect 35000 33696 35016 33760
rect 35080 33696 35096 33760
rect 35160 33696 35176 33760
rect 35240 33696 35248 33760
rect 34928 32672 35248 33696
rect 34928 32608 34936 32672
rect 35000 32608 35016 32672
rect 35080 32608 35096 32672
rect 35160 32608 35176 32672
rect 35240 32608 35248 32672
rect 34928 31584 35248 32608
rect 34928 31520 34936 31584
rect 35000 31520 35016 31584
rect 35080 31520 35096 31584
rect 35160 31520 35176 31584
rect 35240 31520 35248 31584
rect 27107 30700 27173 30701
rect 27107 30636 27108 30700
rect 27172 30636 27173 30700
rect 27107 30635 27173 30636
rect 27110 3637 27170 30635
rect 34928 30496 35248 31520
rect 34928 30432 34936 30496
rect 35000 30432 35016 30496
rect 35080 30432 35096 30496
rect 35160 30432 35176 30496
rect 35240 30432 35248 30496
rect 34928 29408 35248 30432
rect 34928 29344 34936 29408
rect 35000 29344 35016 29408
rect 35080 29344 35096 29408
rect 35160 29344 35176 29408
rect 35240 29344 35248 29408
rect 34928 28320 35248 29344
rect 34928 28256 34936 28320
rect 35000 28256 35016 28320
rect 35080 28256 35096 28320
rect 35160 28256 35176 28320
rect 35240 28256 35248 28320
rect 34928 27232 35248 28256
rect 34928 27168 34936 27232
rect 35000 27168 35016 27232
rect 35080 27168 35096 27232
rect 35160 27168 35176 27232
rect 35240 27168 35248 27232
rect 34928 26144 35248 27168
rect 34928 26080 34936 26144
rect 35000 26080 35016 26144
rect 35080 26080 35096 26144
rect 35160 26080 35176 26144
rect 35240 26080 35248 26144
rect 34928 25056 35248 26080
rect 34928 24992 34936 25056
rect 35000 24992 35016 25056
rect 35080 24992 35096 25056
rect 35160 24992 35176 25056
rect 35240 24992 35248 25056
rect 34928 23968 35248 24992
rect 34928 23904 34936 23968
rect 35000 23904 35016 23968
rect 35080 23904 35096 23968
rect 35160 23904 35176 23968
rect 35240 23904 35248 23968
rect 34928 22880 35248 23904
rect 34928 22816 34936 22880
rect 35000 22816 35016 22880
rect 35080 22816 35096 22880
rect 35160 22816 35176 22880
rect 35240 22816 35248 22880
rect 34928 21792 35248 22816
rect 34928 21728 34936 21792
rect 35000 21728 35016 21792
rect 35080 21728 35096 21792
rect 35160 21728 35176 21792
rect 35240 21728 35248 21792
rect 34928 20704 35248 21728
rect 34928 20640 34936 20704
rect 35000 20640 35016 20704
rect 35080 20640 35096 20704
rect 35160 20640 35176 20704
rect 35240 20640 35248 20704
rect 34928 19616 35248 20640
rect 34928 19552 34936 19616
rect 35000 19552 35016 19616
rect 35080 19552 35096 19616
rect 35160 19552 35176 19616
rect 35240 19552 35248 19616
rect 28763 19276 28829 19277
rect 28763 19212 28764 19276
rect 28828 19212 28829 19276
rect 28763 19211 28829 19212
rect 28766 14517 28826 19211
rect 34928 18528 35248 19552
rect 34928 18464 34936 18528
rect 35000 18464 35016 18528
rect 35080 18464 35096 18528
rect 35160 18464 35176 18528
rect 35240 18464 35248 18528
rect 34928 17440 35248 18464
rect 34928 17376 34936 17440
rect 35000 17376 35016 17440
rect 35080 17376 35096 17440
rect 35160 17376 35176 17440
rect 35240 17376 35248 17440
rect 34928 16352 35248 17376
rect 34928 16288 34936 16352
rect 35000 16288 35016 16352
rect 35080 16288 35096 16352
rect 35160 16288 35176 16352
rect 35240 16288 35248 16352
rect 34928 15264 35248 16288
rect 34928 15200 34936 15264
rect 35000 15200 35016 15264
rect 35080 15200 35096 15264
rect 35160 15200 35176 15264
rect 35240 15200 35248 15264
rect 28763 14516 28829 14517
rect 28763 14452 28764 14516
rect 28828 14452 28829 14516
rect 28763 14451 28829 14452
rect 34928 14176 35248 15200
rect 34928 14112 34936 14176
rect 35000 14112 35016 14176
rect 35080 14112 35096 14176
rect 35160 14112 35176 14176
rect 35240 14112 35248 14176
rect 34928 13088 35248 14112
rect 34928 13024 34936 13088
rect 35000 13024 35016 13088
rect 35080 13024 35096 13088
rect 35160 13024 35176 13088
rect 35240 13024 35248 13088
rect 34928 12000 35248 13024
rect 34928 11936 34936 12000
rect 35000 11936 35016 12000
rect 35080 11936 35096 12000
rect 35160 11936 35176 12000
rect 35240 11936 35248 12000
rect 34928 10912 35248 11936
rect 34928 10848 34936 10912
rect 35000 10848 35016 10912
rect 35080 10848 35096 10912
rect 35160 10848 35176 10912
rect 35240 10848 35248 10912
rect 34928 9824 35248 10848
rect 34928 9760 34936 9824
rect 35000 9760 35016 9824
rect 35080 9760 35096 9824
rect 35160 9760 35176 9824
rect 35240 9760 35248 9824
rect 34928 8736 35248 9760
rect 34928 8672 34936 8736
rect 35000 8672 35016 8736
rect 35080 8672 35096 8736
rect 35160 8672 35176 8736
rect 35240 8672 35248 8736
rect 34928 7648 35248 8672
rect 34928 7584 34936 7648
rect 35000 7584 35016 7648
rect 35080 7584 35096 7648
rect 35160 7584 35176 7648
rect 35240 7584 35248 7648
rect 34928 6560 35248 7584
rect 34928 6496 34936 6560
rect 35000 6496 35016 6560
rect 35080 6496 35096 6560
rect 35160 6496 35176 6560
rect 35240 6496 35248 6560
rect 34928 5472 35248 6496
rect 34928 5408 34936 5472
rect 35000 5408 35016 5472
rect 35080 5408 35096 5472
rect 35160 5408 35176 5472
rect 35240 5408 35248 5472
rect 34928 4384 35248 5408
rect 34928 4320 34936 4384
rect 35000 4320 35016 4384
rect 35080 4320 35096 4384
rect 35160 4320 35176 4384
rect 35240 4320 35248 4384
rect 27107 3636 27173 3637
rect 27107 3572 27108 3636
rect 27172 3572 27173 3636
rect 27107 3571 27173 3572
rect 34928 3296 35248 4320
rect 34928 3232 34936 3296
rect 35000 3232 35016 3296
rect 35080 3232 35096 3296
rect 35160 3232 35176 3296
rect 35240 3232 35248 3296
rect 34928 2208 35248 3232
rect 34928 2144 34936 2208
rect 35000 2144 35016 2208
rect 35080 2144 35096 2208
rect 35160 2144 35176 2208
rect 35240 2144 35248 2208
rect 35588 2176 35908 38624
rect 36248 2176 36568 38624
rect 36908 2176 37228 38624
rect 37779 32060 37845 32061
rect 37779 31996 37780 32060
rect 37844 31996 37845 32060
rect 37779 31995 37845 31996
rect 37782 20365 37842 31995
rect 37779 20364 37845 20365
rect 37779 20300 37780 20364
rect 37844 20300 37845 20364
rect 37779 20299 37845 20300
rect 34928 2128 35248 2144
use sky130_fd_sc_hd__fill_1  FILLER_1_21 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 3036 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_15 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 2484 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 1380 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_15
timestamp 1608254825
transform 1 0 2484 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_3
timestamp 1608254825
transform 1 0 1380 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1608254825
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _2557_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 3128 0 1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_1_41
timestamp 1608254825
transform 1 0 4876 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_44
timestamp 1608254825
transform 1 0 5152 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_32
timestamp 1608254825
transform 1 0 4048 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_66
timestamp 1608254825
transform 1 0 7176 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_62
timestamp 1608254825
transform 1 0 6808 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_53 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 5980 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_63
timestamp 1608254825
transform 1 0 6900 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56
timestamp 1608254825
transform 1 0 6256 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1608254825
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1608254825
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2576_
timestamp 1608254825
transform 1 0 7176 0 -1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__and2_4  _1916_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 7268 0 1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_1_87
timestamp 1608254825
transform 1 0 9108 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_74
timestamp 1608254825
transform 1 0 7912 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_85
timestamp 1608254825
transform 1 0 8924 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _2580_
timestamp 1608254825
transform 1 0 9476 0 1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__nor2_4  _1908_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 8280 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_1_114
timestamp 1608254825
transform 1 0 11592 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_110
timestamp 1608254825
transform 1 0 11224 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_100
timestamp 1608254825
transform 1 0 10304 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_94
timestamp 1608254825
transform 1 0 9752 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1608254825
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2574_
timestamp 1608254825
transform 1 0 10396 0 -1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_1_118
timestamp 1608254825
transform 1 0 11960 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_134
timestamp 1608254825
transform 1 0 13432 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_120
timestamp 1608254825
transform 1 0 12144 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1608254825
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1608254825
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2570_
timestamp 1608254825
transform 1 0 12420 0 1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_2  _1922_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 11684 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_4  _1910_
timestamp 1608254825
transform 1 0 12604 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_1_156
timestamp 1608254825
transform 1 0 15456 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_148
timestamp 1608254825
transform 1 0 14720 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_142
timestamp 1608254825
transform 1 0 14168 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_147
timestamp 1608254825
transform 1 0 14628 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1608254825
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2573_
timestamp 1608254825
transform 1 0 15456 0 -1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__and2_4  _1917_
timestamp 1608254825
transform 1 0 13984 0 -1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _1911_
timestamp 1608254825
transform 1 0 14812 0 1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_1_179
timestamp 1608254825
transform 1 0 17572 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_175
timestamp 1608254825
transform 1 0 17204 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _2565_
timestamp 1608254825
transform 1 0 15824 0 1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_1_191
timestamp 1608254825
transform 1 0 18676 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_187
timestamp 1608254825
transform 1 0 18308 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_183
timestamp 1608254825
transform 1 0 17940 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1608254825
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1608254825
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _1943_
timestamp 1608254825
transform 1 0 18032 0 1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_1_204
timestamp 1608254825
transform 1 0 19872 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_4  _1928_
timestamp 1608254825
transform 1 0 19044 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_0_205
timestamp 1608254825
transform 1 0 19964 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__o21a_4  _2388_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 18860 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_228
timestamp 1608254825
transform 1 0 22080 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_208
timestamp 1608254825
transform 1 0 20240 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_227
timestamp 1608254825
transform 1 0 21988 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1608254825
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2566_
timestamp 1608254825
transform 1 0 20332 0 1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__nand2_4  _2387_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 21160 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_1_239
timestamp 1608254825
transform 1 0 23092 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_231
timestamp 1608254825
transform 1 0 22356 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _1940_
timestamp 1608254825
transform 1 0 22448 0 1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_1_251
timestamp 1608254825
transform 1 0 24196 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_245
timestamp 1608254825
transform 1 0 23644 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_243
timestamp 1608254825
transform 1 0 23460 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_244
timestamp 1608254825
transform 1 0 23552 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1608254825
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1608254825
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _1942_
timestamp 1608254825
transform 1 0 24012 0 -1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_4  _1803_
timestamp 1608254825
transform 1 0 22448 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_271
timestamp 1608254825
transform 1 0 26036 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_273
timestamp 1608254825
transform 1 0 26220 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_260
timestamp 1608254825
transform 1 0 25024 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_256
timestamp 1608254825
transform 1 0 24656 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2636_
timestamp 1608254825
transform 1 0 24288 0 1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__o21a_4  _1800_
timestamp 1608254825
transform 1 0 25116 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_294
timestamp 1608254825
transform 1 0 28152 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_292
timestamp 1608254825
transform 1 0 27968 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1608254825
transform 1 0 26772 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2634_
timestamp 1608254825
transform 1 0 26404 0 1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  _2406_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 28336 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_4  _1802_
timestamp 1608254825
transform 1 0 26864 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_318
timestamp 1608254825
transform 1 0 30360 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_302
timestamp 1608254825
transform 1 0 28888 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_308 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 29440 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_300
timestamp 1608254825
transform 1 0 28704 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1608254825
transform 1 0 29164 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1608254825
transform 1 0 29624 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2562_
timestamp 1608254825
transform 1 0 29716 0 -1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__o21a_4  _1805_
timestamp 1608254825
transform 1 0 29256 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_330
timestamp 1608254825
transform 1 0 31464 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_340
timestamp 1608254825
transform 1 0 32384 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_332
timestamp 1608254825
transform 1 0 31648 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_5 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 31464 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1608254825
transform 1 0 32476 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2558_
timestamp 1608254825
transform 1 0 31556 0 1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__o21a_4  _1807_
timestamp 1608254825
transform 1 0 32568 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_358
timestamp 1608254825
transform 1 0 34040 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_350
timestamp 1608254825
transform 1 0 33304 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_354
timestamp 1608254825
transform 1 0 33672 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _1799_
timestamp 1608254825
transform 1 0 33672 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_387
timestamp 1608254825
transform 1 0 36708 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_379
timestamp 1608254825
transform 1 0 35972 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_366
timestamp 1608254825
transform 1 0 34776 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1608254825
transform 1 0 34776 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1608254825
transform 1 0 35328 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2560_
timestamp 1608254825
transform 1 0 35420 0 -1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _2549_
timestamp 1608254825
transform 1 0 36800 0 1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__o21a_4  _1809_
timestamp 1608254825
transform 1 0 34868 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_407
timestamp 1608254825
transform 1 0 38548 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_0_404
timestamp 1608254825
transform 1 0 38272 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_400
timestamp 1608254825
transform 1 0 37904 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_392
timestamp 1608254825
transform 1 0 37168 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1608254825
transform 1 0 38180 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_415
timestamp 1608254825
transform 1 0 39284 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_416
timestamp 1608254825
transform 1 0 39376 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1608254825
transform -1 0 39836 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1608254825
transform -1 0 39836 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_15
timestamp 1608254825
transform 1 0 2484 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1608254825
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1608254825
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_44
timestamp 1608254825
transform 1 0 5152 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_32
timestamp 1608254825
transform 1 0 4048 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_27
timestamp 1608254825
transform 1 0 3588 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1608254825
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_64
timestamp 1608254825
transform 1 0 6992 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_56
timestamp 1608254825
transform 1 0 6256 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _2591_
timestamp 1608254825
transform 1 0 7176 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_2_91
timestamp 1608254825
transform 1 0 9476 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_85
timestamp 1608254825
transform 1 0 8924 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_2_114
timestamp 1608254825
transform 1 0 11592 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_104
timestamp 1608254825
transform 1 0 10672 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_100
timestamp 1608254825
transform 1 0 10304 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1608254825
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _1903_
timestamp 1608254825
transform 1 0 10764 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__and2_4  _1897_
timestamp 1608254825
transform 1 0 9660 0 -1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_2_122
timestamp 1608254825
transform 1 0 12328 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2579_
timestamp 1608254825
transform 1 0 12420 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  FILLER_2_150
timestamp 1608254825
transform 1 0 14904 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_142
timestamp 1608254825
transform 1 0 14168 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1608254825
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2584_
timestamp 1608254825
transform 1 0 15272 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_2_173
timestamp 1608254825
transform 1 0 17020 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  _2463_
timestamp 1608254825
transform 1 0 17572 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_2_205
timestamp 1608254825
transform 1 0 19964 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_198
timestamp 1608254825
transform 1 0 19320 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1933_
timestamp 1608254825
transform 1 0 19688 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_213
timestamp 1608254825
transform 1 0 20700 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1608254825
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2568_
timestamp 1608254825
transform 1 0 20884 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_2_234
timestamp 1608254825
transform 1 0 22632 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2635_
timestamp 1608254825
transform 1 0 23000 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  FILLER_2_272
timestamp 1608254825
transform 1 0 26128 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_264
timestamp 1608254825
transform 1 0 25392 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_257
timestamp 1608254825
transform 1 0 24748 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2386_
timestamp 1608254825
transform 1 0 25116 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_292
timestamp 1608254825
transform 1 0 27968 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_288
timestamp 1608254825
transform 1 0 27600 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1608254825
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2633_
timestamp 1608254825
transform 1 0 28060 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__o21a_4  _1801_
timestamp 1608254825
transform 1 0 26496 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_312
timestamp 1608254825
transform 1 0 29808 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_4  _1806_
timestamp 1608254825
transform 1 0 30176 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_342
timestamp 1608254825
transform 1 0 32568 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_337
timestamp 1608254825
transform 1 0 32108 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_328
timestamp 1608254825
transform 1 0 31280 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1608254825
transform 1 0 32016 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1798_
timestamp 1608254825
transform 1 0 32200 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_365
timestamp 1608254825
transform 1 0 34684 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _2631_
timestamp 1608254825
transform 1 0 32936 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_2_373
timestamp 1608254825
transform 1 0 35420 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2578_
timestamp 1608254825
transform 1 0 35512 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_2_410
timestamp 1608254825
transform 1 0 38824 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_2_398
timestamp 1608254825
transform 1 0 37720 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_393
timestamp 1608254825
transform 1 0 37260 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1608254825
transform 1 0 37628 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1608254825
transform -1 0 39836 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_15
timestamp 1608254825
transform 1 0 2484 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1608254825
transform 1 0 1380 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1608254825
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_44
timestamp 1608254825
transform 1 0 5152 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_27
timestamp 1608254825
transform 1 0 3588 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__and3_4  _1971_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 4324 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_3_68
timestamp 1608254825
transform 1 0 7360 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_62
timestamp 1608254825
transform 1 0 6808 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_57
timestamp 1608254825
transform 1 0 6348 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1608254825
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__and3_4  _1973_
timestamp 1608254825
transform 1 0 5520 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_3_76
timestamp 1608254825
transform 1 0 8096 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2585_
timestamp 1608254825
transform 1 0 8464 0 1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__and2_4  _1913_
timestamp 1608254825
transform 1 0 7452 0 1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_3_114
timestamp 1608254825
transform 1 0 11592 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_3_99
timestamp 1608254825
transform 1 0 10212 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_4  _1888_
timestamp 1608254825
transform 1 0 10764 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_3_136
timestamp 1608254825
transform 1 0 13616 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_123
timestamp 1608254825
transform 1 0 12420 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1608254825
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _1899_
timestamp 1608254825
transform 1 0 12788 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_3_159
timestamp 1608254825
transform 1 0 15732 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _2460_
timestamp 1608254825
transform 1 0 13984 0 1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_3_182
timestamp 1608254825
transform 1 0 17848 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_176
timestamp 1608254825
transform 1 0 17296 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_4  _1934_
timestamp 1608254825
transform 1 0 16468 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_3_201
timestamp 1608254825
transform 1 0 19596 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_191
timestamp 1608254825
transform 1 0 18676 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_187
timestamp 1608254825
transform 1 0 18308 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1608254825
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2569_
timestamp 1608254825
transform 1 0 19964 0 1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__nor2_4  _1932_
timestamp 1608254825
transform 1 0 18768 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1925_
timestamp 1608254825
transform 1 0 18032 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_224
timestamp 1608254825
transform 1 0 21712 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__and2_4  _1939_
timestamp 1608254825
transform 1 0 22080 0 1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_3_243
timestamp 1608254825
transform 1 0 23460 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_235
timestamp 1608254825
transform 1 0 22724 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1608254825
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_4  _1781_
timestamp 1608254825
transform 1 0 23644 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_273
timestamp 1608254825
transform 1 0 26220 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_257
timestamp 1608254825
transform 1 0 24748 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_4  _1783_
timestamp 1608254825
transform 1 0 25116 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_289
timestamp 1608254825
transform 1 0 27692 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__o21a_4  _1786_
timestamp 1608254825
transform 1 0 26588 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_319
timestamp 1608254825
transform 1 0 30452 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_311
timestamp 1608254825
transform 1 0 29716 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_306
timestamp 1608254825
transform 1 0 29256 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_301
timestamp 1608254825
transform 1 0 28796 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1608254825
transform 1 0 29164 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1773_
timestamp 1608254825
transform 1 0 29440 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_339
timestamp 1608254825
transform 1 0 32292 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2632_
timestamp 1608254825
transform 1 0 30544 0 1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_3_362
timestamp 1608254825
transform 1 0 34408 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_355
timestamp 1608254825
transform 1 0 33764 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_4  _1808_
timestamp 1608254825
transform 1 0 32660 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1797_
timestamp 1608254825
transform 1 0 34132 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_379
timestamp 1608254825
transform 1 0 35972 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1608254825
transform 1 0 34776 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_4  _1811_
timestamp 1608254825
transform 1 0 34868 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_391
timestamp 1608254825
transform 1 0 37076 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2561_
timestamp 1608254825
transform 1 0 37444 0 1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_3_414
timestamp 1608254825
transform 1 0 39192 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1608254825
transform -1 0 39836 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1608254825
transform 1 0 2484 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1608254825
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1608254825
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_36
timestamp 1608254825
transform 1 0 4416 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_32
timestamp 1608254825
transform 1 0 4048 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_27
timestamp 1608254825
transform 1 0 3588 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1608254825
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_4  _1834_
timestamp 1608254825
transform 1 0 4508 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_4_58
timestamp 1608254825
transform 1 0 6440 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_46
timestamp 1608254825
transform 1 0 5336 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _2582_
timestamp 1608254825
transform 1 0 6808 0 -1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  FILLER_4_89
timestamp 1608254825
transform 1 0 9292 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_4_81
timestamp 1608254825
transform 1 0 8556 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_114
timestamp 1608254825
transform 1 0 11592 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_97
timestamp 1608254825
transform 1 0 10028 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_93
timestamp 1608254825
transform 1 0 9660 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1608254825
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _2311_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 10120 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_4_137
timestamp 1608254825
transform 1 0 13708 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2468_
timestamp 1608254825
transform 1 0 11960 0 -1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  FILLER_4_154
timestamp 1608254825
transform 1 0 15272 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_152
timestamp 1608254825
transform 1 0 15088 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_148
timestamp 1608254825
transform 1 0 14720 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1608254825
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _2308_
timestamp 1608254825
transform 1 0 15548 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__and2_4  _1937_
timestamp 1608254825
transform 1 0 14076 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_4_161
timestamp 1608254825
transform 1 0 15916 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2467_
timestamp 1608254825
transform 1 0 16284 0 -1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_4_203
timestamp 1608254825
transform 1 0 19780 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_192
timestamp 1608254825
transform 1 0 18768 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_184
timestamp 1608254825
transform 1 0 18032 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_4  _1926_
timestamp 1608254825
transform 1 0 18952 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_4_215
timestamp 1608254825
transform 1 0 20884 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_210
timestamp 1608254825
transform 1 0 20424 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1608254825
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2643_
timestamp 1608254825
transform 1 0 21252 0 -1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_2  _2296_
timestamp 1608254825
transform 1 0 20148 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_246
timestamp 1608254825
transform 1 0 23736 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_238
timestamp 1608254825
transform 1 0 23000 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_4  _1780_
timestamp 1608254825
transform 1 0 23828 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_271
timestamp 1608254825
transform 1 0 26036 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_259
timestamp 1608254825
transform 1 0 24932 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_292
timestamp 1608254825
transform 1 0 27968 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_288
timestamp 1608254825
transform 1 0 27600 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1608254825
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2640_
timestamp 1608254825
transform 1 0 28060 0 -1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__o21a_4  _1785_
timestamp 1608254825
transform 1 0 26496 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_312
timestamp 1608254825
transform 1 0 29808 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_4  _1788_
timestamp 1608254825
transform 1 0 30176 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_328
timestamp 1608254825
transform 1 0 31280 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1608254825
transform 1 0 32016 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_4  _1791_
timestamp 1608254825
transform 1 0 32108 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_365
timestamp 1608254825
transform 1 0 34684 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_349
timestamp 1608254825
transform 1 0 33212 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_4  _1810_
timestamp 1608254825
transform 1 0 33580 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_381
timestamp 1608254825
transform 1 0 36156 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_4  _1812_
timestamp 1608254825
transform 1 0 35052 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_410
timestamp 1608254825
transform 1 0 38824 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_4_398
timestamp 1608254825
transform 1 0 37720 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_396
timestamp 1608254825
transform 1 0 37536 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_392
timestamp 1608254825
transform 1 0 37168 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1608254825
transform 1 0 37628 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1749_
timestamp 1608254825
transform 1 0 36892 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1608254825
transform -1 0 39836 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_3
timestamp 1608254825
transform 1 0 1380 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1608254825
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _2543_
timestamp 1608254825
transform 1 0 1472 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_5_31
timestamp 1608254825
transform 1 0 3956 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_23
timestamp 1608254825
transform 1 0 3220 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__nand3_4  _1965_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 4048 0 1 4896
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_5_62
timestamp 1608254825
transform 1 0 6808 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_57
timestamp 1608254825
transform 1 0 6348 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_46
timestamp 1608254825
transform 1 0 5336 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1608254825
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _1972_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 5704 0 1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_5_74
timestamp 1608254825
transform 1 0 7912 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _2466_
timestamp 1608254825
transform 1 0 8096 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_5_95
timestamp 1608254825
transform 1 0 9844 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_4  _2313_
timestamp 1608254825
transform 1 0 10212 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_5_132
timestamp 1608254825
transform 1 0 13248 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_121
timestamp 1608254825
transform 1 0 12236 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_115
timestamp 1608254825
transform 1 0 11684 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1608254825
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__o32ai_4  _2327_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 13616 0 1 4896
box -38 -48 2062 592
use sky130_fd_sc_hd__nor2_4  _1923_
timestamp 1608254825
transform 1 0 12420 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_5_158
timestamp 1608254825
transform 1 0 15640 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_182
timestamp 1608254825
transform 1 0 17848 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_178
timestamp 1608254825
transform 1 0 17480 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_4  _2312_
timestamp 1608254825
transform 1 0 16008 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_5_188
timestamp 1608254825
transform 1 0 18400 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_184
timestamp 1608254825
transform 1 0 18032 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1608254825
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2464_
timestamp 1608254825
transform 1 0 18492 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1608254825
transform 1 0 21620 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_215
timestamp 1608254825
transform 1 0 20884 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_5_208
timestamp 1608254825
transform 1 0 20240 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_4  _2131_
timestamp 1608254825
transform 1 0 21712 0 1 4896
box -38 -48 1326 592
use sky130_fd_sc_hd__inv_2  _1931_
timestamp 1608254825
transform 1 0 20608 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_249
timestamp 1608254825
transform 1 0 24012 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_238
timestamp 1608254825
transform 1 0 23000 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1608254825
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1468_
timestamp 1608254825
transform 1 0 23644 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_265
timestamp 1608254825
transform 1 0 25484 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2641_
timestamp 1608254825
transform 1 0 25852 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__o21a_4  _1779_
timestamp 1608254825
transform 1 0 24380 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_296
timestamp 1608254825
transform 1 0 28336 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_288
timestamp 1608254825
transform 1 0 27600 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_5_310
timestamp 1608254825
transform 1 0 29624 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_5_301
timestamp 1608254825
transform 1 0 28796 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1608254825
transform 1 0 29164 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2639_
timestamp 1608254825
transform 1 0 30360 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  _1775_
timestamp 1608254825
transform 1 0 28428 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1502_
timestamp 1608254825
transform 1 0 29256 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_337
timestamp 1608254825
transform 1 0 32108 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_4  _1790_
timestamp 1608254825
transform 1 0 32476 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_365
timestamp 1608254825
transform 1 0 34684 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_353
timestamp 1608254825
transform 1 0 33580 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_374
timestamp 1608254825
transform 1 0 35512 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1608254825
transform 1 0 34776 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2507_
timestamp 1608254825
transform 1 0 36064 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__and2_4  _2102_
timestamp 1608254825
transform 1 0 34868 0 1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_5_399
timestamp 1608254825
transform 1 0 37812 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_4  _1820_
timestamp 1608254825
transform 1 0 38180 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_5_412
timestamp 1608254825
transform 1 0 39008 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1608254825
transform -1 0 39836 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_7
timestamp 1608254825
transform 1 0 1748 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_3
timestamp 1608254825
transform 1 0 1380 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_6_11
timestamp 1608254825
transform 1 0 2116 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_6_3
timestamp 1608254825
transform 1 0 1380 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1608254825
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1608254825
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_4  _1969_
timestamp 1608254825
transform 1 0 1840 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_7_17
timestamp 1608254825
transform 1 0 2668 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_4  _1967_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 2392 0 -1 5984
box -38 -48 1234 592
use sky130_fd_sc_hd__nor3_4  _1835_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 3036 0 1 5984
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_7_34
timestamp 1608254825
transform 1 0 4232 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_45
timestamp 1608254825
transform 1 0 5244 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_41
timestamp 1608254825
transform 1 0 4876 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_27
timestamp 1608254825
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1608254825
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2542_
timestamp 1608254825
transform 1 0 4600 0 1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__nor2_4  _1966_
timestamp 1608254825
transform 1 0 4048 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_7_62
timestamp 1608254825
transform 1 0 6808 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_57
timestamp 1608254825
transform 1 0 6348 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_65
timestamp 1608254825
transform 1 0 7084 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1608254825
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2541_
timestamp 1608254825
transform 1 0 5336 0 -1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_6_88
timestamp 1608254825
transform 1 0 9200 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_77
timestamp 1608254825
transform 1 0 8188 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _2470_
timestamp 1608254825
transform 1 0 7912 0 1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_2  _1927_
timestamp 1608254825
transform 1 0 8924 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_7_93
timestamp 1608254825
transform 1 0 9660 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_6_109
timestamp 1608254825
transform 1 0 11132 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1608254825
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2458_
timestamp 1608254825
transform 1 0 10212 0 1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__a2bb2o_4  _2309_
timestamp 1608254825
transform 1 0 9660 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_7_137
timestamp 1608254825
transform 1 0 13708 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_126
timestamp 1608254825
transform 1 0 12696 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_7_118
timestamp 1608254825
transform 1 0 11960 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_134
timestamp 1608254825
transform 1 0 13432 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1608254825
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2469_
timestamp 1608254825
transform 1 0 11684 0 -1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_2  _1902_
timestamp 1608254825
transform 1 0 12420 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1638_
timestamp 1608254825
transform 1 0 13432 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_157
timestamp 1608254825
transform 1 0 15548 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_141
timestamp 1608254825
transform 1 0 14076 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1608254825
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__o32ai_4  _2325_
timestamp 1608254825
transform 1 0 14076 0 1 5984
box -38 -48 2062 592
use sky130_fd_sc_hd__inv_2  _1920_
timestamp 1608254825
transform 1 0 13800 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1898_
timestamp 1608254825
transform 1 0 15272 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_179
timestamp 1608254825
transform 1 0 17572 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_171
timestamp 1608254825
transform 1 0 16836 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_163
timestamp 1608254825
transform 1 0 16100 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_177
timestamp 1608254825
transform 1 0 17388 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_4  _2316_
timestamp 1608254825
transform 1 0 15916 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__a2bb2o_4  _2315_
timestamp 1608254825
transform 1 0 17756 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  _2306_
timestamp 1608254825
transform 1 0 17204 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1924_
timestamp 1608254825
transform 1 0 16468 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_187
timestamp 1608254825
transform 1 0 18308 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_204
timestamp 1608254825
transform 1 0 19872 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_197
timestamp 1608254825
transform 1 0 19228 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_188
timestamp 1608254825
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2492_
timestamp 1608254825
transform 1 0 18676 0 1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_2  _1929_
timestamp 1608254825
transform 1 0 19596 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1909_
timestamp 1608254825
transform 1 0 18032 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_7_228
timestamp 1608254825
transform 1 0 22080 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_7_210
timestamp 1608254825
transform 1 0 20424 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_212
timestamp 1608254825
transform 1 0 20608 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1608254825
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__nand3_4  _2129_
timestamp 1608254825
transform 1 0 20792 0 1 5984
box -38 -48 1326 592
use sky130_fd_sc_hd__nand3_4  _2125_
timestamp 1608254825
transform 1 0 20884 0 -1 5984
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_2  FILLER_7_245
timestamp 1608254825
transform 1 0 23644 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_240
timestamp 1608254825
transform 1 0 23184 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_236
timestamp 1608254825
transform 1 0 22816 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_237
timestamp 1608254825
transform 1 0 22908 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_229
timestamp 1608254825
transform 1 0 22172 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_189
timestamp 1608254825
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2642_
timestamp 1608254825
transform 1 0 23000 0 -1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__o21a_4  _1782_
timestamp 1608254825
transform 1 0 23828 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1700_
timestamp 1608254825
transform 1 0 22908 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_259
timestamp 1608254825
transform 1 0 24932 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_273
timestamp 1608254825
transform 1 0 26220 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_265
timestamp 1608254825
transform 1 0 25484 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_257
timestamp 1608254825
transform 1 0 24748 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2644_
timestamp 1608254825
transform 1 0 25300 0 1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  _1777_
timestamp 1608254825
transform 1 0 25116 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_282
timestamp 1608254825
transform 1 0 27048 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_292
timestamp 1608254825
transform 1 0 27968 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_288
timestamp 1608254825
transform 1 0 27600 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_4_0_addressalyzerBlock.SPI_CLK $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 27416 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1608254825
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_4  _1795_
timestamp 1608254825
transform 1 0 27692 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__o21a_4  _1787_
timestamp 1608254825
transform 1 0 28060 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__o21a_4  _1778_
timestamp 1608254825
transform 1 0 26496 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_301
timestamp 1608254825
transform 1 0 28796 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_305
timestamp 1608254825
transform 1 0 29164 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_190
timestamp 1608254825
transform 1 0 29164 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1804_
timestamp 1608254825
transform 1 0 29256 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_310
timestamp 1608254825
transform 1 0 29624 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_319
timestamp 1608254825
transform 1 0 30452 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_313
timestamp 1608254825
transform 1 0 29900 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_addressalyzerBlock.SPI_CLK
timestamp 1608254825
transform 1 0 29992 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1774_
timestamp 1608254825
transform 1 0 29532 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2638_
timestamp 1608254825
transform 1 0 30268 0 1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_7_336
timestamp 1608254825
transform 1 0 32016 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_332
timestamp 1608254825
transform 1 0 31648 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1608254825
transform 1 0 32016 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2630_
timestamp 1608254825
transform 1 0 32384 0 1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__o21a_4  _1793_
timestamp 1608254825
transform 1 0 32108 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__o21a_4  _1792_
timestamp 1608254825
transform 1 0 30544 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_365
timestamp 1608254825
transform 1 0 34684 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_359
timestamp 1608254825
transform 1 0 34132 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_357
timestamp 1608254825
transform 1 0 33948 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_349
timestamp 1608254825
transform 1 0 33212 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _2629_
timestamp 1608254825
transform 1 0 34040 0 -1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_7_371
timestamp 1608254825
transform 1 0 35236 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_367
timestamp 1608254825
transform 1 0 34868 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_377
timestamp 1608254825
transform 1 0 35788 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_191
timestamp 1608254825
transform 1 0 34776 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2647_
timestamp 1608254825
transform 1 0 35328 0 1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__o21a_4  _1816_
timestamp 1608254825
transform 1 0 36156 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_391
timestamp 1608254825
transform 1 0 37076 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_407
timestamp 1608254825
transform 1 0 38548 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_393
timestamp 1608254825
transform 1 0 37260 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1608254825
transform 1 0 37628 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2628_
timestamp 1608254825
transform 1 0 37444 0 1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_2  _1818_
timestamp 1608254825
transform 1 0 38916 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_4  _1750_
timestamp 1608254825
transform 1 0 37720 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_7_414
timestamp 1608254825
transform 1 0 39192 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_414
timestamp 1608254825
transform 1 0 39192 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1608254825
transform -1 0 39836 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1608254825
transform -1 0 39836 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_3
timestamp 1608254825
transform 1 0 1380 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1608254825
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_4  _1968_
timestamp 1608254825
transform 1 0 2116 0 -1 7072
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_6  FILLER_8_32
timestamp 1608254825
transform 1 0 4048 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_30
timestamp 1608254825
transform 1 0 3864 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_24
timestamp 1608254825
transform 1 0 3312 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_192
timestamp 1608254825
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__a21o_4  _1970_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 4600 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_50
timestamp 1608254825
transform 1 0 5704 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  _2453_
timestamp 1608254825
transform 1 0 6256 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_8_88
timestamp 1608254825
transform 1 0 9200 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_83
timestamp 1608254825
transform 1 0 8740 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_75
timestamp 1608254825
transform 1 0 8004 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1918_
timestamp 1608254825
transform 1 0 8924 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_102
timestamp 1608254825
transform 1 0 10488 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_193
timestamp 1608254825
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _2310_
timestamp 1608254825
transform 1 0 11224 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__nor2_4  _1919_
timestamp 1608254825
transform 1 0 9660 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_8_126
timestamp 1608254825
transform 1 0 12696 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2462_
timestamp 1608254825
transform 1 0 13064 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_8_157
timestamp 1608254825
transform 1 0 15548 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_8_149
timestamp 1608254825
transform 1 0 14812 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_194
timestamp 1608254825
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1550_
timestamp 1608254825
transform 1 0 15272 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_165
timestamp 1608254825
transform 1 0 16284 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _2465_
timestamp 1608254825
transform 1 0 16468 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_8_194
timestamp 1608254825
transform 1 0 18952 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_186
timestamp 1608254825
transform 1 0 18216 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__nand3_4  _2118_
timestamp 1608254825
transform 1 0 19136 0 -1 7072
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_2  FILLER_8_215
timestamp 1608254825
transform 1 0 20884 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_210
timestamp 1608254825
transform 1 0 20424 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_195
timestamp 1608254825
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__nand3_4  _2133_
timestamp 1608254825
transform 1 0 21068 0 -1 7072
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_1  FILLER_8_235
timestamp 1608254825
transform 1 0 22724 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_231
timestamp 1608254825
transform 1 0 22356 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_4  _2355_
timestamp 1608254825
transform 1 0 22816 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_8_274
timestamp 1608254825
transform 1 0 26312 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_268
timestamp 1608254825
transform 1 0 25760 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_260
timestamp 1608254825
transform 1 0 25024 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_252
timestamp 1608254825
transform 1 0 24288 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1789_
timestamp 1608254825
transform 1 0 25392 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1481_
timestamp 1608254825
transform 1 0 24656 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_285
timestamp 1608254825
transform 1 0 27324 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_280
timestamp 1608254825
transform 1 0 26864 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_276
timestamp 1608254825
transform 1 0 26496 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_196
timestamp 1608254825
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2637_
timestamp 1608254825
transform 1 0 27692 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  _1784_
timestamp 1608254825
transform 1 0 26956 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_308
timestamp 1608254825
transform 1 0 29440 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_4  _1796_
timestamp 1608254825
transform 1 0 29808 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_342
timestamp 1608254825
transform 1 0 32568 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_337
timestamp 1608254825
transform 1 0 32108 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_335
timestamp 1608254825
transform 1 0 31924 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_331
timestamp 1608254825
transform 1 0 31556 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_324
timestamp 1608254825
transform 1 0 30912 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_5_0_addressalyzerBlock.SPI_CLK
timestamp 1608254825
transform 1 0 31280 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_197
timestamp 1608254825
transform 1 0 32016 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1826_
timestamp 1608254825
transform 1 0 32292 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_358
timestamp 1608254825
transform 1 0 34040 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_4  _1814_
timestamp 1608254825
transform 1 0 34408 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__o21a_4  _1813_
timestamp 1608254825
transform 1 0 32936 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_374
timestamp 1608254825
transform 1 0 35512 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_4  _1817_
timestamp 1608254825
transform 1 0 35880 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_398
timestamp 1608254825
transform 1 0 37720 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_396
timestamp 1608254825
transform 1 0 37536 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_390
timestamp 1608254825
transform 1 0 36984 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_198
timestamp 1608254825
transform 1 0 37628 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_4  _1821_
timestamp 1608254825
transform 1 0 37812 0 -1 7072
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_6  FILLER_8_412
timestamp 1608254825
transform 1 0 39008 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1608254825
transform -1 0 39836 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_17
timestamp 1608254825
transform 1 0 2668 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_3
timestamp 1608254825
transform 1 0 1380 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1608254825
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_4  _2391_
timestamp 1608254825
transform 1 0 1564 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _2389_
timestamp 1608254825
transform 1 0 3036 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_28
timestamp 1608254825
transform 1 0 3680 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_24
timestamp 1608254825
transform 1 0 3312 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2540_
timestamp 1608254825
transform 1 0 3772 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_9_60
timestamp 1608254825
transform 1 0 6624 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_48
timestamp 1608254825
transform 1 0 5520 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_199
timestamp 1608254825
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_4  _2338_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 6808 0 1 7072
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_1  FILLER_9_81
timestamp 1608254825
transform 1 0 8556 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_75
timestamp 1608254825
transform 1 0 8004 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_4  _2335_
timestamp 1608254825
transform 1 0 8648 0 1 7072
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_9_109
timestamp 1608254825
transform 1 0 11132 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_96
timestamp 1608254825
transform 1 0 9936 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1906_
timestamp 1608254825
transform 1 0 11500 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_4  _1551_
timestamp 1608254825
transform 1 0 10304 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_9_132
timestamp 1608254825
transform 1 0 13248 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_121
timestamp 1608254825
transform 1 0 12236 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_117
timestamp 1608254825
transform 1 0 11868 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_1_0_addressalyzerBlock.SPI_CLK
timestamp 1608254825
transform 1 0 13616 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_200
timestamp 1608254825
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _1921_
timestamp 1608254825
transform 1 0 12420 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__o32ai_4  _2323_
timestamp 1608254825
transform 1 0 13892 0 1 7072
box -38 -48 2062 592
use sky130_fd_sc_hd__decap_8  FILLER_9_175
timestamp 1608254825
transform 1 0 17204 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_165
timestamp 1608254825
transform 1 0 16284 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_161
timestamp 1608254825
transform 1 0 15916 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_4  _1930_
timestamp 1608254825
transform 1 0 16376 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_9_197
timestamp 1608254825
transform 1 0 19228 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_201
timestamp 1608254825
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__nand3_4  _2121_
timestamp 1608254825
transform 1 0 19596 0 1 7072
box -38 -48 1326 592
use sky130_fd_sc_hd__o21ai_4  _2119_
timestamp 1608254825
transform 1 0 18032 0 1 7072
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_6  FILLER_9_215
timestamp 1608254825
transform 1 0 20884 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_4  _2358_
timestamp 1608254825
transform 1 0 21436 0 1 7072
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_3  FILLER_9_241
timestamp 1608254825
transform 1 0 23276 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_234
timestamp 1608254825
transform 1 0 22632 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_2_0_m1_clk_local
timestamp 1608254825
transform 1 0 23000 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_202
timestamp 1608254825
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2446_
timestamp 1608254825
transform 1 0 23644 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_9_264
timestamp 1608254825
transform 1 0 25392 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1672_
timestamp 1608254825
transform 1 0 26128 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_290
timestamp 1608254825
transform 1 0 27784 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_283
timestamp 1608254825
transform 1 0 27140 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_275
timestamp 1608254825
transform 1 0 26404 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__and2_4  _2087_
timestamp 1608254825
transform 1 0 28152 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1489_
timestamp 1608254825
transform 1 0 27508 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1452_
timestamp 1608254825
transform 1 0 26772 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_309
timestamp 1608254825
transform 1 0 29532 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_301
timestamp 1608254825
transform 1 0 28796 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_203
timestamp 1608254825
transform 1 0 29164 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2511_
timestamp 1608254825
transform 1 0 29900 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_2  _1532_
timestamp 1608254825
transform 1 0 29256 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_9_332
timestamp 1608254825
transform 1 0 31648 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  _2500_
timestamp 1608254825
transform 1 0 32200 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_9_365
timestamp 1608254825
transform 1 0 34684 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_357
timestamp 1608254825
transform 1 0 33948 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_367
timestamp 1608254825
transform 1 0 34868 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_204
timestamp 1608254825
transform 1 0 34776 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2627_
timestamp 1608254825
transform 1 0 35144 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_9_395
timestamp 1608254825
transform 1 0 37444 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_389
timestamp 1608254825
transform 1 0 36892 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__nand4_4  _1747_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 37536 0 1 7072
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_1  FILLER_9_417
timestamp 1608254825
transform 1 0 39468 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_413
timestamp 1608254825
transform 1 0 39100 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1608254825
transform -1 0 39836 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_7
timestamp 1608254825
transform 1 0 1748 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_3
timestamp 1608254825
transform 1 0 1380 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1608254825
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _2625_
timestamp 1608254825
transform 1 0 1840 0 -1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_10_42
timestamp 1608254825
transform 1 0 4968 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_36
timestamp 1608254825
transform 1 0 4416 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_32
timestamp 1608254825
transform 1 0 4048 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_27
timestamp 1608254825
transform 1 0 3588 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_205
timestamp 1608254825
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2452_
timestamp 1608254825
transform 1 0 5060 0 -1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_2  _1975_
timestamp 1608254825
transform 1 0 4140 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_10_62
timestamp 1608254825
transform 1 0 6808 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_4  _2337_
timestamp 1608254825
transform 1 0 7360 0 -1 8160
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_2  FILLER_10_90
timestamp 1608254825
transform 1 0 9384 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_82
timestamp 1608254825
transform 1 0 8648 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_112
timestamp 1608254825
transform 1 0 11408 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_106
timestamp 1608254825
transform 1 0 10856 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_206
timestamp 1608254825
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_4  _2336_
timestamp 1608254825
transform 1 0 9660 0 -1 8160
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_4  _2141_
timestamp 1608254825
transform 1 0 11500 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_10_122
timestamp 1608254825
transform 1 0 12328 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2461_
timestamp 1608254825
transform 1 0 12696 0 -1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_10_158
timestamp 1608254825
transform 1 0 15640 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_145
timestamp 1608254825
transform 1 0 14444 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_207
timestamp 1608254825
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _2320_
timestamp 1608254825
transform 1 0 15272 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_182
timestamp 1608254825
transform 1 0 17848 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_165
timestamp 1608254825
transform 1 0 16284 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_0_0_m1_clk_local
timestamp 1608254825
transform 1 0 16008 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_4  _2314_
timestamp 1608254825
transform 1 0 16376 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_10_200
timestamp 1608254825
transform 1 0 19504 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _2117_
timestamp 1608254825
transform 1 0 19872 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_4  _2116_
timestamp 1608254825
transform 1 0 18216 0 -1 8160
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_10_221
timestamp 1608254825
transform 1 0 21436 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_10_215
timestamp 1608254825
transform 1 0 20884 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_10_208
timestamp 1608254825
transform 1 0 20240 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_208
timestamp 1608254825
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2445_
timestamp 1608254825
transform 1 0 21804 0 -1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_2  _2356_
timestamp 1608254825
transform 1 0 21160 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_251
timestamp 1608254825
transform 1 0 24196 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_244
timestamp 1608254825
transform 1 0 23552 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1564_
timestamp 1608254825
transform 1 0 23920 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_271
timestamp 1608254825
transform 1 0 26036 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_4  _2360_
timestamp 1608254825
transform 1 0 24564 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_10_295
timestamp 1608254825
transform 1 0 28244 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_209
timestamp 1608254825
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2443_
timestamp 1608254825
transform 1 0 26496 0 -1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp 1608254825
transform 1 0 29348 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_303
timestamp 1608254825
transform 1 0 28980 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1794_
timestamp 1608254825
transform 1 0 28612 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_4  _1741_
timestamp 1608254825
transform 1 0 29440 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_340
timestamp 1608254825
transform 1 0 32384 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_332
timestamp 1608254825
transform 1 0 31648 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_324
timestamp 1608254825
transform 1 0 30912 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_320
timestamp 1608254825
transform 1 0 30544 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_210
timestamp 1608254825
transform 1 0 32016 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _2086_
timestamp 1608254825
transform 1 0 31004 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1737_
timestamp 1608254825
transform 1 0 32108 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_351
timestamp 1608254825
transform 1 0 33396 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2501_
timestamp 1608254825
transform 1 0 33764 0 -1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__and2_4  _2100_
timestamp 1608254825
transform 1 0 32752 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_10_374
timestamp 1608254825
transform 1 0 35512 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_4  _1824_
timestamp 1608254825
transform 1 0 36064 0 -1 8160
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_10_393
timestamp 1608254825
transform 1 0 37260 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_211
timestamp 1608254825
transform 1 0 37628 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__nand3_4  _1819_
timestamp 1608254825
transform 1 0 37720 0 -1 8160
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_6  FILLER_10_412
timestamp 1608254825
transform 1 0 39008 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1608254825
transform -1 0 39836 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_11
timestamp 1608254825
transform 1 0 2116 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_3
timestamp 1608254825
transform 1 0 1380 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1608254825
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_4  _1836_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 2208 0 1 8160
box -38 -48 2062 592
use sky130_fd_sc_hd__decap_12  FILLER_11_34
timestamp 1608254825
transform 1 0 4232 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_62
timestamp 1608254825
transform 1 0 6808 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_58
timestamp 1608254825
transform 1 0 6440 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_46
timestamp 1608254825
transform 1 0 5336 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_212
timestamp 1608254825
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__nand3_4  _2339_
timestamp 1608254825
transform 1 0 6900 0 1 8160
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_11_77
timestamp 1608254825
transform 1 0 8188 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2454_
timestamp 1608254825
transform 1 0 8556 0 1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_11_100
timestamp 1608254825
transform 1 0 10304 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_4  _2142_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 10672 0 1 8160
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_11_132
timestamp 1608254825
transform 1 0 13248 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_118
timestamp 1608254825
transform 1 0 11960 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_213
timestamp 1608254825
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__o32ai_4  _2324_
timestamp 1608254825
transform 1 0 13616 0 1 8160
box -38 -48 2062 592
use sky130_fd_sc_hd__nor2_4  _1639_
timestamp 1608254825
transform 1 0 12420 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_11_158
timestamp 1608254825
transform 1 0 15640 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_181
timestamp 1608254825
transform 1 0 17756 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_174
timestamp 1608254825
transform 1 0 17112 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_166
timestamp 1608254825
transform 1 0 16376 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_m1_clk_local
timestamp 1608254825
transform 1 0 17480 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _2322_
timestamp 1608254825
transform 1 0 16744 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _2317_
timestamp 1608254825
transform 1 0 16008 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_198
timestamp 1608254825
transform 1 0 19320 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_214
timestamp 1608254825
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2491_
timestamp 1608254825
transform 1 0 19688 0 1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__nand3_4  _2120_
timestamp 1608254825
transform 1 0 18032 0 1 8160
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_11_221
timestamp 1608254825
transform 1 0 21436 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_4  _2357_
timestamp 1608254825
transform 1 0 21804 0 1 8160
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_11_245
timestamp 1608254825
transform 1 0 23644 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_243
timestamp 1608254825
transform 1 0 23460 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_239
timestamp 1608254825
transform 1 0 23092 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_215
timestamp 1608254825
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1761_
timestamp 1608254825
transform 1 0 24012 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_252
timestamp 1608254825
transform 1 0 24288 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2441_
timestamp 1608254825
transform 1 0 24656 0 1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_11_293
timestamp 1608254825
transform 1 0 28060 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_285
timestamp 1608254825
transform 1 0 27324 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_281
timestamp 1608254825
transform 1 0 26956 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_275
timestamp 1608254825
transform 1 0 26404 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _1827_
timestamp 1608254825
transform 1 0 27692 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1760_
timestamp 1608254825
transform 1 0 27048 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_301
timestamp 1608254825
transform 1 0 28796 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_216
timestamp 1608254825
transform 1 0 29164 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2649_
timestamp 1608254825
transform 1 0 29256 0 1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  _1815_
timestamp 1608254825
transform 1 0 28428 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_337
timestamp 1608254825
transform 1 0 32108 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_329
timestamp 1608254825
transform 1 0 31372 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_325
timestamp 1608254825
transform 1 0 31004 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2502_
timestamp 1608254825
transform 1 0 32476 0 1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__and2_4  _2101_
timestamp 1608254825
transform 1 0 31464 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_11_360
timestamp 1608254825
transform 1 0 34224 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_11_381
timestamp 1608254825
transform 1 0 36156 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_367
timestamp 1608254825
transform 1 0 34868 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_217
timestamp 1608254825
transform 1 0 34776 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2626_
timestamp 1608254825
transform 1 0 36524 0 1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__a21o_4  _1825_
timestamp 1608254825
transform 1 0 35052 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_411
timestamp 1608254825
transform 1 0 38916 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_11_404
timestamp 1608254825
transform 1 0 38272 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1823_
timestamp 1608254825
transform 1 0 38640 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_417
timestamp 1608254825
transform 1 0 39468 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1608254825
transform -1 0 39836 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_12_17
timestamp 1608254825
transform 1 0 2668 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_13
timestamp 1608254825
transform 1 0 2300 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_3
timestamp 1608254825
transform 1 0 1380 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1608254825
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_4  _2390_
timestamp 1608254825
transform 1 0 1472 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_4  _1837_
timestamp 1608254825
transform 1 0 2760 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_12_45
timestamp 1608254825
transform 1 0 5244 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_41
timestamp 1608254825
transform 1 0 4876 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_27
timestamp 1608254825
transform 1 0 3588 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_218
timestamp 1608254825
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__or3_4  _1974_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 4048 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_12_68
timestamp 1608254825
transform 1 0 7360 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__o32ai_4  _2297_
timestamp 1608254825
transform 1 0 5336 0 -1 9248
box -38 -48 2062 592
use sky130_fd_sc_hd__fill_2  FILLER_12_87
timestamp 1608254825
transform 1 0 9108 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_12_75
timestamp 1608254825
transform 1 0 8004 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_0_0_addressalyzerBlock.SPI_CLK
timestamp 1608254825
transform 1 0 9292 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1642_
timestamp 1608254825
transform 1 0 7728 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_12_107
timestamp 1608254825
transform 1 0 10948 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_219
timestamp 1608254825
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__a211o_4  _1640_
timestamp 1608254825
transform 1 0 11500 0 -1 9248
box -38 -48 1326 592
use sky130_fd_sc_hd__a211o_4  _1552_
timestamp 1608254825
transform 1 0 9660 0 -1 9248
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_3  FILLER_12_134
timestamp 1608254825
transform 1 0 13432 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_127
timestamp 1608254825
transform 1 0 12788 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_addressalyzerBlock.SPI_CLK
timestamp 1608254825
transform 1 0 13156 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_4  _2251_
timestamp 1608254825
transform 1 0 13708 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_12_154
timestamp 1608254825
transform 1 0 15272 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_152
timestamp 1608254825
transform 1 0 15088 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_146
timestamp 1608254825
transform 1 0 14536 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_220
timestamp 1608254825
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_179
timestamp 1608254825
transform 1 0 17572 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2455_
timestamp 1608254825
transform 1 0 15824 0 -1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_12_197
timestamp 1608254825
transform 1 0 19228 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_4  _2137_
timestamp 1608254825
transform 1 0 17940 0 -1 9248
box -38 -48 1326 592
use sky130_fd_sc_hd__nor2_4  _1565_
timestamp 1608254825
transform 1 0 19596 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_12_228
timestamp 1608254825
transform 1 0 22080 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_210
timestamp 1608254825
transform 1 0 20424 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_221
timestamp 1608254825
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_4  _2122_
timestamp 1608254825
transform 1 0 20884 0 -1 9248
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_6  FILLER_12_244
timestamp 1608254825
transform 1 0 23552 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_236
timestamp 1608254825
transform 1 0 22816 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_4  _2362_
timestamp 1608254825
transform 1 0 24104 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  _2354_
timestamp 1608254825
transform 1 0 23184 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _2343_
timestamp 1608254825
transform 1 0 22448 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_274
timestamp 1608254825
transform 1 0 26312 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_266
timestamp 1608254825
transform 1 0 25576 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_12_296
timestamp 1608254825
transform 1 0 28336 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_283
timestamp 1608254825
transform 1 0 27140 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_279
timestamp 1608254825
transform 1 0 26772 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_222
timestamp 1608254825
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1752_
timestamp 1608254825
transform 1 0 26496 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_4  _1711_
timestamp 1608254825
transform 1 0 27232 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_312
timestamp 1608254825
transform 1 0 29808 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_308
timestamp 1608254825
transform 1 0 29440 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_304
timestamp 1608254825
transform 1 0 29072 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_addressalyzerBlock.SPI_CLK
timestamp 1608254825
transform 1 0 29532 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_4  _1740_
timestamp 1608254825
transform 1 0 29900 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _1697_
timestamp 1608254825
transform 1 0 28704 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_337
timestamp 1608254825
transform 1 0 32108 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_332
timestamp 1608254825
transform 1 0 31648 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_325
timestamp 1608254825
transform 1 0 31004 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_223
timestamp 1608254825
transform 1 0 32016 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__a21o_4  _1734_
timestamp 1608254825
transform 1 0 32292 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1729_
timestamp 1608254825
transform 1 0 31372 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_359
timestamp 1608254825
transform 1 0 34132 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_351
timestamp 1608254825
transform 1 0 33396 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _2503_
timestamp 1608254825
transform 1 0 34316 0 -1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_12_380
timestamp 1608254825
transform 1 0 36064 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__and2_4  _2085_
timestamp 1608254825
transform 1 0 36432 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_12_410
timestamp 1608254825
transform 1 0 38824 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_12_391
timestamp 1608254825
transform 1 0 37076 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_224
timestamp 1608254825
transform 1 0 37628 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_4  _1831_
timestamp 1608254825
transform 1 0 37720 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1608254825
transform -1 0 39836 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_22
timestamp 1608254825
transform 1 0 3128 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_11
timestamp 1608254825
transform 1 0 2116 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_3
timestamp 1608254825
transform 1 0 1380 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1608254825
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1608254825
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _2411_
timestamp 1608254825
transform 1 0 2300 0 1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _2409_
timestamp 1608254825
transform 1 0 1380 0 -1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_14_32
timestamp 1608254825
transform 1 0 4048 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_30
timestamp 1608254825
transform 1 0 3864 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_26
timestamp 1608254825
transform 1 0 3496 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_32
timestamp 1608254825
transform 1 0 4048 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_4_0_m1_clk_local
timestamp 1608254825
transform 1 0 3588 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_231
timestamp 1608254825
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2477_
timestamp 1608254825
transform 1 0 4600 0 1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _2476_
timestamp 1608254825
transform 1 0 4416 0 -1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_14_55
timestamp 1608254825
transform 1 0 6164 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_57
timestamp 1608254825
transform 1 0 6348 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_225
timestamp 1608254825
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_4  _2340_
timestamp 1608254825
transform 1 0 6808 0 1 9248
box -38 -48 1234 592
use sky130_fd_sc_hd__o32ai_4  _2295_
timestamp 1608254825
transform 1 0 6532 0 -1 10336
box -38 -48 2062 592
use sky130_fd_sc_hd__decap_4  FILLER_14_88
timestamp 1608254825
transform 1 0 9200 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_81
timestamp 1608254825
transform 1 0 8556 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_84
timestamp 1608254825
transform 1 0 8832 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_75
timestamp 1608254825
transform 1 0 8004 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1907_
timestamp 1608254825
transform 1 0 8556 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_4  _1556_
timestamp 1608254825
transform 1 0 9200 0 1 9248
box -38 -48 1326 592
use sky130_fd_sc_hd__inv_2  _1554_
timestamp 1608254825
transform 1 0 8924 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_102
timestamp 1608254825
transform 1 0 10488 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_102
timestamp 1608254825
transform 1 0 10488 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_232
timestamp 1608254825
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__a21o_4  _2145_
timestamp 1608254825
transform 1 0 10856 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__a211o_4  _1644_
timestamp 1608254825
transform 1 0 11224 0 -1 10336
box -38 -48 1326 592
use sky130_fd_sc_hd__nor2_4  _1555_
timestamp 1608254825
transform 1 0 9660 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_14_124
timestamp 1608254825
transform 1 0 12512 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_135
timestamp 1608254825
transform 1 0 13524 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_127
timestamp 1608254825
transform 1 0 12788 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_118
timestamp 1608254825
transform 1 0 11960 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_226
timestamp 1608254825
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2456_
timestamp 1608254825
transform 1 0 12880 0 -1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  _1553_
timestamp 1608254825
transform 1 0 13156 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1549_
timestamp 1608254825
transform 1 0 12420 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_154
timestamp 1608254825
transform 1 0 15272 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_14_147
timestamp 1608254825
transform 1 0 14628 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_141
timestamp 1608254825
transform 1 0 14076 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_233
timestamp 1608254825
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__o32ai_4  _2326_
timestamp 1608254825
transform 1 0 14168 0 1 9248
box -38 -48 2062 592
use sky130_fd_sc_hd__decap_4  FILLER_14_182
timestamp 1608254825
transform 1 0 17848 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_179
timestamp 1608254825
transform 1 0 17572 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_171
timestamp 1608254825
transform 1 0 16836 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_164
timestamp 1608254825
transform 1 0 16192 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__o32ai_4  _2330_
timestamp 1608254825
transform 1 0 15824 0 -1 10336
box -38 -48 2062 592
use sky130_fd_sc_hd__buf_2  _1563_
timestamp 1608254825
transform 1 0 17204 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1517_
timestamp 1608254825
transform 1 0 16560 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_190
timestamp 1608254825
transform 1 0 18584 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_200
timestamp 1608254825
transform 1 0 19504 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_184
timestamp 1608254825
transform 1 0 18032 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_227
timestamp 1608254825
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__nand3_4  _2135_
timestamp 1608254825
transform 1 0 18216 0 1 9248
box -38 -48 1326 592
use sky130_fd_sc_hd__a211o_4  _1566_
timestamp 1608254825
transform 1 0 18952 0 -1 10336
box -38 -48 1326 592
use sky130_fd_sc_hd__buf_2  _1561_
timestamp 1608254825
transform 1 0 18216 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1522_
timestamp 1608254825
transform 1 0 19872 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_14_228
timestamp 1608254825
transform 1 0 22080 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_224
timestamp 1608254825
transform 1 0 21712 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_208
timestamp 1608254825
transform 1 0 20240 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_224
timestamp 1608254825
transform 1 0 21712 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_207
timestamp 1608254825
transform 1 0 20148 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_234
timestamp 1608254825
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_4  _1651_
timestamp 1608254825
transform 1 0 22080 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_4  _1650_
timestamp 1608254825
transform 1 0 20516 0 1 9248
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_4  _1649_
timestamp 1608254825
transform 1 0 20884 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_14_248
timestamp 1608254825
transform 1 0 23920 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_237
timestamp 1608254825
transform 1 0 22908 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_m1_clk_local
timestamp 1608254825
transform 1 0 23276 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_228
timestamp 1608254825
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2442_
timestamp 1608254825
transform 1 0 22172 0 -1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__a2bb2o_4  _2361_
timestamp 1608254825
transform 1 0 23644 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_14_271
timestamp 1608254825
transform 1 0 26036 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_261
timestamp 1608254825
transform 1 0 25116 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2444_
timestamp 1608254825
transform 1 0 25484 0 1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _2440_
timestamp 1608254825
transform 1 0 24288 0 -1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_14_276
timestamp 1608254825
transform 1 0 26496 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_284
timestamp 1608254825
transform 1 0 27232 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_235
timestamp 1608254825
transform 1 0 26404 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2653_
timestamp 1608254825
transform 1 0 26864 0 -1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__o21ai_4  _1701_
timestamp 1608254825
transform 1 0 27600 0 1 9248
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_14_312
timestamp 1608254825
transform 1 0 29808 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_299
timestamp 1608254825
transform 1 0 28612 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_319
timestamp 1608254825
transform 1 0 30452 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_301
timestamp 1608254825
transform 1 0 28796 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_229
timestamp 1608254825
transform 1 0 29164 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__and4_4  _1765_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 28980 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_4  _1739_
timestamp 1608254825
transform 1 0 30176 0 -1 10336
box -38 -48 1234 592
use sky130_fd_sc_hd__o21ai_4  _1736_
timestamp 1608254825
transform 1 0 29256 0 1 9248
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_1  FILLER_14_335
timestamp 1608254825
transform 1 0 31924 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_329
timestamp 1608254825
transform 1 0 31372 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_330
timestamp 1608254825
transform 1 0 31464 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_addressalyzerBlock.SPI_CLK
timestamp 1608254825
transform 1 0 30820 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_236
timestamp 1608254825
transform 1 0 32016 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _2103_
timestamp 1608254825
transform 1 0 32108 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_4  _1731_
timestamp 1608254825
transform 1 0 31832 0 1 9248
box -38 -48 1234 592
use sky130_fd_sc_hd__buf_2  _1695_
timestamp 1608254825
transform 1 0 31096 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_344
timestamp 1608254825
transform 1 0 32752 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_360
timestamp 1608254825
transform 1 0 34224 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_347
timestamp 1608254825
transform 1 0 33028 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_7_0_addressalyzerBlock.SPI_CLK
timestamp 1608254825
transform 1 0 33120 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _2650_
timestamp 1608254825
transform 1 0 33396 0 -1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__nand2_4  _1732_
timestamp 1608254825
transform 1 0 33396 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_14_370
timestamp 1608254825
transform 1 0 35144 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_371
timestamp 1608254825
transform 1 0 35236 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_230
timestamp 1608254825
transform 1 0 34776 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2548_
timestamp 1608254825
transform 1 0 35512 0 -1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__nand3_4  _1829_
timestamp 1608254825
transform 1 0 35788 0 1 9248
box -38 -48 1326 592
use sky130_fd_sc_hd__buf_2  _1716_
timestamp 1608254825
transform 1 0 34868 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_407
timestamp 1608254825
transform 1 0 38548 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_393
timestamp 1608254825
transform 1 0 37260 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_391
timestamp 1608254825
transform 1 0 37076 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_4
timestamp 1608254825
transform 1 0 37260 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_237
timestamp 1608254825
transform 1 0 37628 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2539_
timestamp 1608254825
transform 1 0 37444 0 1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_2  _1830_
timestamp 1608254825
transform 1 0 38916 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_4  _1822_
timestamp 1608254825
transform 1 0 37720 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_14_414
timestamp 1608254825
transform 1 0 39192 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_414
timestamp 1608254825
transform 1 0 39192 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1608254825
transform -1 0 39836 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1608254825
transform -1 0 39836 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_22
timestamp 1608254825
transform 1 0 3128 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1608254825
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _2410_
timestamp 1608254825
transform 1 0 1380 0 1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_15_45
timestamp 1608254825
transform 1 0 5244 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  _2412_
timestamp 1608254825
transform 1 0 3496 0 1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_15_55
timestamp 1608254825
transform 1 0 6164 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_51
timestamp 1608254825
transform 1 0 5796 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_238
timestamp 1608254825
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2478_
timestamp 1608254825
transform 1 0 6808 0 1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_2  _1876_
timestamp 1608254825
transform 1 0 5888 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_15_81
timestamp 1608254825
transform 1 0 8556 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_4  _1557_
timestamp 1608254825
transform 1 0 9292 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_15_98
timestamp 1608254825
transform 1 0 10120 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_4  _1645_
timestamp 1608254825
transform 1 0 10856 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_132
timestamp 1608254825
transform 1 0 13248 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_118
timestamp 1608254825
transform 1 0 11960 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_239
timestamp 1608254825
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_4  _2199_
timestamp 1608254825
transform 1 0 12420 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__o32ai_4  _2329_
timestamp 1608254825
transform 1 0 13800 0 1 10336
box -38 -48 2062 592
use sky130_fd_sc_hd__fill_1  FILLER_15_182
timestamp 1608254825
transform 1 0 17848 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_178
timestamp 1608254825
transform 1 0 17480 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_167
timestamp 1608254825
transform 1 0 16468 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_160
timestamp 1608254825
transform 1 0 15824 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_1_0_m1_clk_local
timestamp 1608254825
transform 1 0 16192 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_4  _2223_
timestamp 1608254825
transform 1 0 16652 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_15_192
timestamp 1608254825
transform 1 0 18768 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_188
timestamp 1608254825
transform 1 0 18400 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_240
timestamp 1608254825
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__a21boi_4  _1567_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 18860 0 1 10336
box -38 -48 1418 592
use sky130_fd_sc_hd__buf_2  _1545_
timestamp 1608254825
transform 1 0 18032 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_215
timestamp 1608254825
transform 1 0 20884 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_208
timestamp 1608254825
transform 1 0 20240 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_m1_clk_local
timestamp 1608254825
transform 1 0 20608 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_4  _1648_
timestamp 1608254825
transform 1 0 20976 0 1 10336
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_15_250
timestamp 1608254825
transform 1 0 24104 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_245
timestamp 1608254825
transform 1 0 23644 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_240
timestamp 1608254825
transform 1 0 23184 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_233
timestamp 1608254825
transform 1 0 22540 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_229
timestamp 1608254825
transform 1 0 22172 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_3_0_m1_clk_local
timestamp 1608254825
transform 1 0 22632 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_241
timestamp 1608254825
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _2352_
timestamp 1608254825
transform 1 0 23736 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1758_
timestamp 1608254825
transform 1 0 22908 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_15_273
timestamp 1608254825
transform 1 0 26220 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_addressalyzerBlock.SPI_CLK
timestamp 1608254825
transform 1 0 24472 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_4  _2359_
timestamp 1608254825
transform 1 0 24748 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_15_285
timestamp 1608254825
transform 1 0 27324 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_4  _1710_
timestamp 1608254825
transform 1 0 27692 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _1679_
timestamp 1608254825
transform 1 0 26956 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_306
timestamp 1608254825
transform 1 0 29256 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_301
timestamp 1608254825
transform 1 0 28796 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_242
timestamp 1608254825
transform 1 0 29164 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__a22oi_4  _1764_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 29624 0 1 10336
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_6  FILLER_15_327
timestamp 1608254825
transform 1 0 31188 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__nand4_4  _1730_
timestamp 1608254825
transform 1 0 31740 0 1 10336
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_8  FILLER_15_358
timestamp 1608254825
transform 1 0 34040 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_15_350
timestamp 1608254825
transform 1 0 33304 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1686_
timestamp 1608254825
transform 1 0 33672 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_380
timestamp 1608254825
transform 1 0 36064 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_376
timestamp 1608254825
transform 1 0 35696 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_243
timestamp 1608254825
transform 1 0 34776 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2513_
timestamp 1608254825
transform 1 0 36156 0 1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__nand2_4  _1719_
timestamp 1608254825
transform 1 0 34868 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_15_400
timestamp 1608254825
transform 1 0 37904 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_412
timestamp 1608254825
transform 1 0 39008 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1608254825
transform -1 0 39836 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_22
timestamp 1608254825
transform 1 0 3128 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_16_3
timestamp 1608254825
transform 1 0 1380 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1608254825
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_4  _1833_
timestamp 1608254825
transform 1 0 1932 0 -1 11424
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_1  FILLER_16_44
timestamp 1608254825
transform 1 0 5152 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_32
timestamp 1608254825
transform 1 0 4048 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_30
timestamp 1608254825
transform 1 0 3864 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_244
timestamp 1608254825
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__o32ai_4  _2298_
timestamp 1608254825
transform 1 0 5244 0 -1 11424
box -38 -48 2062 592
use sky130_fd_sc_hd__decap_4  FILLER_16_67
timestamp 1608254825
transform 1 0 7268 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_88
timestamp 1608254825
transform 1 0 9200 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_75
timestamp 1608254825
transform 1 0 8004 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_71
timestamp 1608254825
transform 1 0 7636 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _2300_
timestamp 1608254825
transform 1 0 7728 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_4  _1643_
timestamp 1608254825
transform 1 0 8372 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_16_102
timestamp 1608254825
transform 1 0 10488 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_addressalyzerBlock.SPI_CLK
timestamp 1608254825
transform 1 0 11040 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_245
timestamp 1608254825
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__a211o_4  _2144_
timestamp 1608254825
transform 1 0 11316 0 -1 11424
box -38 -48 1326 592
use sky130_fd_sc_hd__nor2_4  _2143_
timestamp 1608254825
transform 1 0 9660 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_16_125
timestamp 1608254825
transform 1 0 12604 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_4  _2225_
timestamp 1608254825
transform 1 0 12972 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_16_152
timestamp 1608254825
transform 1 0 15088 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_146
timestamp 1608254825
transform 1 0 14536 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_138
timestamp 1608254825
transform 1 0 13800 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_246
timestamp 1608254825
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2459_
timestamp 1608254825
transform 1 0 15272 0 -1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  _2173_
timestamp 1608254825
transform 1 0 14168 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_179
timestamp 1608254825
transform 1 0 17572 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_173
timestamp 1608254825
transform 1 0 17020 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_4  _2249_
timestamp 1608254825
transform 1 0 17664 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_16_202
timestamp 1608254825
transform 1 0 19688 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_189
timestamp 1608254825
transform 1 0 18492 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_4  _2177_
timestamp 1608254825
transform 1 0 18860 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_16_215
timestamp 1608254825
transform 1 0 20884 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_210
timestamp 1608254825
transform 1 0 20424 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_247
timestamp 1608254825
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_4  _2146_
timestamp 1608254825
transform 1 0 20976 0 -1 11424
box -38 -48 1234 592
use sky130_fd_sc_hd__buf_2  _1562_
timestamp 1608254825
transform 1 0 20056 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_240
timestamp 1608254825
transform 1 0 23184 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_236
timestamp 1608254825
transform 1 0 22816 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_229
timestamp 1608254825
transform 1 0 22172 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_4  _2363_
timestamp 1608254825
transform 1 0 23276 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  _1558_
timestamp 1608254825
transform 1 0 22540 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_271
timestamp 1608254825
transform 1 0 26036 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_264
timestamp 1608254825
transform 1 0 25392 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_257
timestamp 1608254825
transform 1 0 24748 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1751_
timestamp 1608254825
transform 1 0 25116 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1702_
timestamp 1608254825
transform 1 0 25760 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_16_291
timestamp 1608254825
transform 1 0 27876 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_285
timestamp 1608254825
transform 1 0 27324 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_6_0_addressalyzerBlock.SPI_CLK
timestamp 1608254825
transform 1 0 27968 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_248
timestamp 1608254825
transform 1 0 26404 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_4  _1759_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 28244 0 -1 11424
box -38 -48 1326 592
use sky130_fd_sc_hd__nor2_4  _1753_
timestamp 1608254825
transform 1 0 26496 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_16_309
timestamp 1608254825
transform 1 0 29532 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_4  _1762_
timestamp 1608254825
transform 1 0 29900 0 -1 11424
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_1  FILLER_16_335
timestamp 1608254825
transform 1 0 31924 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_327
timestamp 1608254825
transform 1 0 31188 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_249
timestamp 1608254825
transform 1 0 32016 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_4  _1684_
timestamp 1608254825
transform 1 0 32108 0 -1 11424
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_16_350
timestamp 1608254825
transform 1 0 33304 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_4  _1735_
timestamp 1608254825
transform 1 0 33672 0 -1 11424
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_1  FILLER_16_373
timestamp 1608254825
transform 1 0 35420 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_367
timestamp 1608254825
transform 1 0 34868 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  _2497_
timestamp 1608254825
transform 1 0 35512 0 -1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_16_405
timestamp 1608254825
transform 1 0 38364 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_393
timestamp 1608254825
transform 1 0 37260 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_250
timestamp 1608254825
transform 1 0 37628 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _2106_
timestamp 1608254825
transform 1 0 37720 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _2083_
timestamp 1608254825
transform 1 0 38732 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_16_412
timestamp 1608254825
transform 1 0 39008 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1608254825
transform -1 0 39836 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_20
timestamp 1608254825
transform 1 0 2944 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_15
timestamp 1608254825
transform 1 0 2484 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1608254825
transform 1 0 1380 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1608254825
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1832_
timestamp 1608254825
transform 1 0 2668 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_43
timestamp 1608254825
transform 1 0 5060 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _2413_
timestamp 1608254825
transform 1 0 3312 0 1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_17_55
timestamp 1608254825
transform 1 0 6164 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_251
timestamp 1608254825
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2474_
timestamp 1608254825
transform 1 0 6808 0 1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_17_91
timestamp 1608254825
transform 1 0 9476 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_87
timestamp 1608254825
transform 1 0 9108 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_81
timestamp 1608254825
transform 1 0 8556 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _2332_
timestamp 1608254825
transform 1 0 9200 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_109
timestamp 1608254825
transform 1 0 11132 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_4  _2197_
timestamp 1608254825
transform 1 0 9844 0 1 11424
box -38 -48 1326 592
use sky130_fd_sc_hd__buf_2  _1641_
timestamp 1608254825
transform 1 0 11500 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_127
timestamp 1608254825
transform 1 0 12788 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_121
timestamp 1608254825
transform 1 0 12236 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_117
timestamp 1608254825
transform 1 0 11868 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_252
timestamp 1608254825
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__nand3_4  _2250_
timestamp 1608254825
transform 1 0 13340 0 1 11424
box -38 -48 1326 592
use sky130_fd_sc_hd__buf_2  _1548_
timestamp 1608254825
transform 1 0 12420 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_155
timestamp 1608254825
transform 1 0 15364 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_147
timestamp 1608254825
transform 1 0 14628 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_4  _2171_
timestamp 1608254825
transform 1 0 15456 0 1 11424
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_17_179
timestamp 1608254825
transform 1 0 17572 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_169
timestamp 1608254825
transform 1 0 16652 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _1560_
timestamp 1608254825
transform 1 0 17204 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_192
timestamp 1608254825
transform 1 0 18768 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_188
timestamp 1608254825
transform 1 0 18400 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_253
timestamp 1608254825
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_4  _2244_
timestamp 1608254825
transform 1 0 18860 0 1 11424
box -38 -48 1234 592
use sky130_fd_sc_hd__buf_2  _1546_
timestamp 1608254825
transform 1 0 18032 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_223
timestamp 1608254825
transform 1 0 21620 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_206
timestamp 1608254825
transform 1 0 20056 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_4  _2226_
timestamp 1608254825
transform 1 0 20424 0 1 11424
box -38 -48 1234 592
use sky130_fd_sc_hd__a21oi_4  _2202_
timestamp 1608254825
transform 1 0 21988 0 1 11424
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_12  FILLER_17_245
timestamp 1608254825
transform 1 0 23644 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_240
timestamp 1608254825
transform 1 0 23184 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_254
timestamp 1608254825
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__xor2_4  _1755_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 24748 0 1 11424
box -38 -48 2062 592
use sky130_fd_sc_hd__decap_4  FILLER_17_279
timestamp 1608254825
transform 1 0 26772 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__a2111o_4  _1756_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 27140 0 1 11424
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_1  FILLER_17_306
timestamp 1608254825
transform 1 0 29256 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_304
timestamp 1608254825
transform 1 0 29072 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_300
timestamp 1608254825
transform 1 0 28704 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_255
timestamp 1608254825
transform 1 0 29164 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__a22oi_4  _1763_
timestamp 1608254825
transform 1 0 29348 0 1 11424
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_17_332
timestamp 1608254825
transform 1 0 31648 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_324
timestamp 1608254825
transform 1 0 30912 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1715_
timestamp 1608254825
transform 1 0 31280 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_4  _1687_
timestamp 1608254825
transform 1 0 32016 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_17_362
timestamp 1608254825
transform 1 0 34408 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_345
timestamp 1608254825
transform 1 0 32844 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_4  _1723_
timestamp 1608254825
transform 1 0 33212 0 1 11424
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_8  FILLER_17_384
timestamp 1608254825
transform 1 0 36432 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_371
timestamp 1608254825
transform 1 0 35236 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_367
timestamp 1608254825
transform 1 0 34868 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_256
timestamp 1608254825
transform 1 0 34776 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__a21o_4  _1766_
timestamp 1608254825
transform 1 0 35328 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_17_392
timestamp 1608254825
transform 1 0 37168 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _2496_
timestamp 1608254825
transform 1 0 37444 0 1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_17_414
timestamp 1608254825
transform 1 0 39192 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1608254825
transform -1 0 39836 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_18_7
timestamp 1608254825
transform 1 0 1748 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_3
timestamp 1608254825
transform 1 0 1380 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1608254825
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _2414_
timestamp 1608254825
transform 1 0 1840 0 -1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_18_45
timestamp 1608254825
transform 1 0 5244 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_39
timestamp 1608254825
transform 1 0 4692 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_32
timestamp 1608254825
transform 1 0 4048 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_27
timestamp 1608254825
transform 1 0 3588 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_m1_clk_local
timestamp 1608254825
transform 1 0 4416 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_257
timestamp 1608254825
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_68
timestamp 1608254825
transform 1 0 7360 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__o32ai_4  _2301_
timestamp 1608254825
transform 1 0 5336 0 -1 12512
box -38 -48 2062 592
use sky130_fd_sc_hd__decap_6  FILLER_18_86
timestamp 1608254825
transform 1 0 9016 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_4  _2344_
timestamp 1608254825
transform 1 0 7728 0 -1 12512
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_18_107
timestamp 1608254825
transform 1 0 10948 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_258
timestamp 1608254825
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__nand3_4  _2224_
timestamp 1608254825
transform 1 0 11316 0 -1 12512
box -38 -48 1326 592
use sky130_fd_sc_hd__nand3_4  _2200_
timestamp 1608254825
transform 1 0 9660 0 -1 12512
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_18_125
timestamp 1608254825
transform 1 0 12604 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_4  _2247_
timestamp 1608254825
transform 1 0 12972 0 -1 12512
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_2  FILLER_18_151
timestamp 1608254825
transform 1 0 14996 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_143
timestamp 1608254825
transform 1 0 14260 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_259
timestamp 1608254825
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_4  _2245_
timestamp 1608254825
transform 1 0 15272 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_18_169
timestamp 1608254825
transform 1 0 16652 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_163
timestamp 1608254825
transform 1 0 16100 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_4  _2273_
timestamp 1608254825
transform 1 0 16744 0 -1 12512
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_18_202
timestamp 1608254825
transform 1 0 19688 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_184
timestamp 1608254825
transform 1 0 18032 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_4  _2178_
timestamp 1608254825
transform 1 0 18400 0 -1 12512
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_6  FILLER_18_224
timestamp 1608254825
transform 1 0 21712 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_210
timestamp 1608254825
transform 1 0 20424 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_260
timestamp 1608254825
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_4  _2243_
timestamp 1608254825
transform 1 0 20884 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _1559_
timestamp 1608254825
transform 1 0 20056 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_246
timestamp 1608254825
transform 1 0 23736 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2439_
timestamp 1608254825
transform 1 0 24104 0 -1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__a2bb2o_4  _2364_
timestamp 1608254825
transform 1 0 22264 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_18_269
timestamp 1608254825
transform 1 0 25852 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_284
timestamp 1608254825
transform 1 0 27232 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_280
timestamp 1608254825
transform 1 0 26864 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_276
timestamp 1608254825
transform 1 0 26496 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_261
timestamp 1608254825
transform 1 0 26404 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_4  _1709_
timestamp 1608254825
transform 1 0 27600 0 -1 12512
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _1705_
timestamp 1608254825
transform 1 0 26956 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_18_313
timestamp 1608254825
transform 1 0 29900 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_309
timestamp 1608254825
transform 1 0 29532 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_301
timestamp 1608254825
transform 1 0 28796 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1706_
timestamp 1608254825
transform 1 0 29164 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__and4_4  _1678_
timestamp 1608254825
transform 1 0 29992 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_18_330
timestamp 1608254825
transform 1 0 31464 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_323
timestamp 1608254825
transform 1 0 30820 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_262
timestamp 1608254825
transform 1 0 32016 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1738_
timestamp 1608254825
transform 1 0 31188 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__o32ai_4  _1718_
timestamp 1608254825
transform 1 0 32108 0 -1 12512
box -38 -48 2062 592
use sky130_fd_sc_hd__decap_4  FILLER_18_359
timestamp 1608254825
transform 1 0 34132 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2652_
timestamp 1608254825
transform 1 0 34500 0 -1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_18_382
timestamp 1608254825
transform 1 0 36248 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_402
timestamp 1608254825
transform 1 0 38088 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_398
timestamp 1608254825
transform 1 0 37720 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_393
timestamp 1608254825
transform 1 0 37260 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_263
timestamp 1608254825
transform 1 0 37628 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_4  _1771_
timestamp 1608254825
transform 1 0 38180 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1616_
timestamp 1608254825
transform 1 0 36984 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_18_412
timestamp 1608254825
transform 1 0 39008 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1608254825
transform -1 0 39836 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_20_22
timestamp 1608254825
transform 1 0 3128 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_22
timestamp 1608254825
transform 1 0 3128 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1608254825
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1608254825
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _2416_
timestamp 1608254825
transform 1 0 1380 0 -1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _2415_
timestamp 1608254825
transform 1 0 1380 0 1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_20_30
timestamp 1608254825
transform 1 0 3864 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_45
timestamp 1608254825
transform 1 0 5244 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_270
timestamp 1608254825
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2419_
timestamp 1608254825
transform 1 0 4048 0 -1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _2417_
timestamp 1608254825
transform 1 0 3496 0 1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_20_55
timestamp 1608254825
transform 1 0 6164 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_51
timestamp 1608254825
transform 1 0 5796 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_57
timestamp 1608254825
transform 1 0 6348 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_53
timestamp 1608254825
transform 1 0 5980 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1880_
timestamp 1608254825
transform 1 0 6072 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1878_
timestamp 1608254825
transform 1 0 6256 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_59
timestamp 1608254825
transform 1 0 6532 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_62
timestamp 1608254825
transform 1 0 6808 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_264
timestamp 1608254825
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2450_
timestamp 1608254825
transform 1 0 6992 0 1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__o21ai_4  _2345_
timestamp 1608254825
transform 1 0 6900 0 -1 13600
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_20_88
timestamp 1608254825
transform 1 0 9200 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_76
timestamp 1608254825
transform 1 0 8096 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_83
timestamp 1608254825
transform 1 0 8740 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _2333_
timestamp 1608254825
transform 1 0 8832 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_4  _2196_
timestamp 1608254825
transform 1 0 9108 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_20_106
timestamp 1608254825
transform 1 0 10856 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_93
timestamp 1608254825
transform 1 0 9660 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_109
timestamp 1608254825
transform 1 0 11132 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_96
timestamp 1608254825
transform 1 0 9936 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_271
timestamp 1608254825
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__nand3_4  _2221_
timestamp 1608254825
transform 1 0 11408 0 -1 13600
box -38 -48 1326 592
use sky130_fd_sc_hd__nand2_4  _2201_
timestamp 1608254825
transform 1 0 10028 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  _2198_
timestamp 1608254825
transform 1 0 10304 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_20_126
timestamp 1608254825
transform 1 0 12696 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_132
timestamp 1608254825
transform 1 0 13248 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_118
timestamp 1608254825
transform 1 0 11960 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_265
timestamp 1608254825
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_4  _2219_
timestamp 1608254825
transform 1 0 13064 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  _2195_
timestamp 1608254825
transform 1 0 12420 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1547_
timestamp 1608254825
transform 1 0 11684 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_149
timestamp 1608254825
transform 1 0 14812 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_139
timestamp 1608254825
transform 1 0 13892 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_143
timestamp 1608254825
transform 1 0 14260 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_138
timestamp 1608254825
transform 1 0 13800 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_272
timestamp 1608254825
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_4  _2267_
timestamp 1608254825
transform 1 0 14628 0 1 12512
box -38 -48 1234 592
use sky130_fd_sc_hd__o21ai_4  _2172_
timestamp 1608254825
transform 1 0 15272 0 -1 13600
box -38 -48 1234 592
use sky130_fd_sc_hd__buf_2  _2170_
timestamp 1608254825
transform 1 0 13892 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1647_
timestamp 1608254825
transform 1 0 14444 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_181
timestamp 1608254825
transform 1 0 17756 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_175
timestamp 1608254825
transform 1 0 17204 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_167
timestamp 1608254825
transform 1 0 16468 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_177
timestamp 1608254825
transform 1 0 17388 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_160
timestamp 1608254825
transform 1 0 15824 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_4  _2266_
timestamp 1608254825
transform 1 0 16192 0 1 12512
box -38 -48 1234 592
use sky130_fd_sc_hd__buf_2  _2194_
timestamp 1608254825
transform 1 0 16836 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__a21boi_4  _2179_
timestamp 1608254825
transform 1 0 17848 0 -1 13600
box -38 -48 1418 592
use sky130_fd_sc_hd__decap_4  FILLER_20_197
timestamp 1608254825
transform 1 0 19228 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_203
timestamp 1608254825
transform 1 0 19780 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_199
timestamp 1608254825
transform 1 0 19412 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_266
timestamp 1608254825
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__a21boi_4  _2274_
timestamp 1608254825
transform 1 0 18032 0 1 12512
box -38 -48 1418 592
use sky130_fd_sc_hd__a22oi_4  _2252_
timestamp 1608254825
transform 1 0 19872 0 1 12512
box -38 -48 1602 592
use sky130_fd_sc_hd__nand2_4  _2147_
timestamp 1608254825
transform 1 0 19596 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_20_228
timestamp 1608254825
transform 1 0 22080 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_210
timestamp 1608254825
transform 1 0 20424 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_221
timestamp 1608254825
transform 1 0 21436 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_273
timestamp 1608254825
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_4  _2203_
timestamp 1608254825
transform 1 0 21804 0 1 12512
box -38 -48 1234 592
use sky130_fd_sc_hd__a21oi_4  _2148_
timestamp 1608254825
transform 1 0 20884 0 -1 13600
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_20_247
timestamp 1608254825
transform 1 0 23828 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_245
timestamp 1608254825
transform 1 0 23644 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_19_238
timestamp 1608254825
transform 1 0 23000 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_267
timestamp 1608254825
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_4  _2227_
timestamp 1608254825
transform 1 0 24196 0 -1 13600
box -38 -48 1234 592
use sky130_fd_sc_hd__a21boi_4  _2204_
timestamp 1608254825
transform 1 0 22448 0 -1 13600
box -38 -48 1418 592
use sky130_fd_sc_hd__decap_3  FILLER_20_272
timestamp 1608254825
transform 1 0 26128 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_20_264
timestamp 1608254825
transform 1 0 25392 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_257
timestamp 1608254825
transform 1 0 24748 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_253
timestamp 1608254825
transform 1 0 24380 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _2271_
timestamp 1608254825
transform 1 0 24472 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_4  _1754_
timestamp 1608254825
transform 1 0 25116 0 1 12512
box -38 -48 2062 592
use sky130_fd_sc_hd__fill_1  FILLER_20_280
timestamp 1608254825
transform 1 0 26864 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_276
timestamp 1608254825
transform 1 0 26496 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_287
timestamp 1608254825
transform 1 0 27508 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_283
timestamp 1608254825
transform 1 0 27140 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_274
timestamp 1608254825
transform 1 0 26404 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__a41o_4  _1733_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 26956 0 -1 13600
box -38 -48 1602 592
use sky130_fd_sc_hd__and4_4  _1704_
timestamp 1608254825
transform 1 0 27600 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_20_298
timestamp 1608254825
transform 1 0 28520 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_19_297
timestamp 1608254825
transform 1 0 28428 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_268
timestamp 1608254825
transform 1 0 29164 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__and4_4  _1681_
timestamp 1608254825
transform 1 0 29072 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _1680_
timestamp 1608254825
transform 1 0 29256 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_313
timestamp 1608254825
transform 1 0 29900 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_314
timestamp 1608254825
transform 1 0 29992 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_310
timestamp 1608254825
transform 1 0 29624 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__and4_4  _1724_
timestamp 1608254825
transform 1 0 30084 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_4  _1725_
timestamp 1608254825
transform 1 0 30452 0 -1 13600
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_6  FILLER_20_341
timestamp 1608254825
transform 1 0 32476 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_332
timestamp 1608254825
transform 1 0 31648 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_324
timestamp 1608254825
transform 1 0 30912 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_275
timestamp 1608254825
transform 1 0 32016 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__nand4_4  _1717_
timestamp 1608254825
transform 1 0 31280 0 1 12512
box -38 -48 1602 592
use sky130_fd_sc_hd__buf_2  _1682_
timestamp 1608254825
transform 1 0 32108 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_365
timestamp 1608254825
transform 1 0 34684 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_361
timestamp 1608254825
transform 1 0 34316 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_347
timestamp 1608254825
transform 1 0 33028 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_362
timestamp 1608254825
transform 1 0 34408 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_345
timestamp 1608254825
transform 1 0 32844 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_4  _1721_
timestamp 1608254825
transform 1 0 33212 0 1 12512
box -38 -48 1234 592
use sky130_fd_sc_hd__a21oi_4  _1691_
timestamp 1608254825
transform 1 0 33120 0 -1 13600
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_1  FILLER_20_378
timestamp 1608254825
transform 1 0 35880 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_370
timestamp 1608254825
transform 1 0 35144 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_370
timestamp 1608254825
transform 1 0 35144 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_269
timestamp 1608254825
transform 1 0 34776 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _2099_
timestamp 1608254825
transform 1 0 34776 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__nand4_4  _1770_
timestamp 1608254825
transform 1 0 35512 0 1 12512
box -38 -48 1602 592
use sky130_fd_sc_hd__nand3_4  _1767_
timestamp 1608254825
transform 1 0 35972 0 -1 13600
box -38 -48 1326 592
use sky130_fd_sc_hd__inv_2  _1757_
timestamp 1608254825
transform 1 0 34868 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_20_411
timestamp 1608254825
transform 1 0 38916 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_393
timestamp 1608254825
transform 1 0 37260 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_391
timestamp 1608254825
transform 1 0 37076 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_276
timestamp 1608254825
transform 1 0 37628 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2645_
timestamp 1608254825
transform 1 0 37444 0 1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__a21oi_4  _1772_
timestamp 1608254825
transform 1 0 37720 0 -1 13600
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_1  FILLER_20_417
timestamp 1608254825
transform 1 0 39468 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_414
timestamp 1608254825
transform 1 0 39192 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1608254825
transform -1 0 39836 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1608254825
transform -1 0 39836 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_18
timestamp 1608254825
transform 1 0 2760 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1608254825
transform 1 0 1380 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_5_0_m1_clk_local
timestamp 1608254825
transform 1 0 2484 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1608254825
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _2418_
timestamp 1608254825
transform 1 0 3128 0 1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_21_41
timestamp 1608254825
transform 1 0 4876 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_57
timestamp 1608254825
transform 1 0 6348 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_277
timestamp 1608254825
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__o32ai_4  _2299_
timestamp 1608254825
transform 1 0 6808 0 1 13600
box -38 -48 2062 592
use sky130_fd_sc_hd__buf_2  _2294_
timestamp 1608254825
transform 1 0 5980 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_84
timestamp 1608254825
transform 1 0 8832 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2448_
timestamp 1608254825
transform 1 0 9200 0 1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_21_107
timestamp 1608254825
transform 1 0 10948 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _2334_
timestamp 1608254825
transform 1 0 11316 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_127
timestamp 1608254825
transform 1 0 12788 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_123
timestamp 1608254825
transform 1 0 12420 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_115
timestamp 1608254825
transform 1 0 11684 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_addressalyzerBlock.SPI_CLK
timestamp 1608254825
transform 1 0 12052 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_278
timestamp 1608254825
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_4  _2174_
timestamp 1608254825
transform 1 0 13156 0 1 13600
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _1646_
timestamp 1608254825
transform 1 0 12512 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_21_151
timestamp 1608254825
transform 1 0 14996 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_144
timestamp 1608254825
transform 1 0 14352 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_3_0_addressalyzerBlock.SPI_CLK
timestamp 1608254825
transform 1 0 14720 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_4  _2175_
timestamp 1608254825
transform 1 0 15088 0 1 13600
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_1  FILLER_21_182
timestamp 1608254825
transform 1 0 17848 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_178
timestamp 1608254825
transform 1 0 17480 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_165
timestamp 1608254825
transform 1 0 16284 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_4  _2176_
timestamp 1608254825
transform 1 0 16652 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_21_193
timestamp 1608254825
transform 1 0 18860 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_279
timestamp 1608254825
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2486_
timestamp 1608254825
transform 1 0 19412 0 1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__nand2_4  _2270_
timestamp 1608254825
transform 1 0 18032 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_21_224
timestamp 1608254825
transform 1 0 21712 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_218
timestamp 1608254825
transform 1 0 21160 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__a21boi_4  _2228_
timestamp 1608254825
transform 1 0 21804 0 1 13600
box -38 -48 1418 592
use sky130_fd_sc_hd__decap_4  FILLER_21_240
timestamp 1608254825
transform 1 0 23184 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_280
timestamp 1608254825
transform 1 0 23552 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _1948_
timestamp 1608254825
transform 1 0 23644 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_21_266
timestamp 1608254825
transform 1 0 25576 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_258
timestamp 1608254825
transform 1 0 24840 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_254
timestamp 1608254825
transform 1 0 24472 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__and2_4  _1960_
timestamp 1608254825
transform 1 0 24932 0 1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_4  _1708_
timestamp 1608254825
transform 1 0 25944 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_21_296
timestamp 1608254825
transform 1 0 28336 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_21_279
timestamp 1608254825
transform 1 0 26772 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_4  _1742_
timestamp 1608254825
transform 1 0 27140 0 1 13600
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_8  FILLER_21_315
timestamp 1608254825
transform 1 0 30084 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_304
timestamp 1608254825
transform 1 0 29072 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_281
timestamp 1608254825
transform 1 0 29164 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__and4_4  _1692_
timestamp 1608254825
transform 1 0 29256 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__a41oi_4  _1720_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 30820 0 1 13600
box -38 -48 2062 592
use sky130_fd_sc_hd__decap_4  FILLER_21_362
timestamp 1608254825
transform 1 0 34408 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_345
timestamp 1608254825
transform 1 0 32844 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_4  _1690_
timestamp 1608254825
transform 1 0 33212 0 1 13600
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_1  FILLER_21_373
timestamp 1608254825
transform 1 0 35420 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_367
timestamp 1608254825
transform 1 0 34868 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_282
timestamp 1608254825
transform 1 0 34776 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2659_
timestamp 1608254825
transform 1 0 35512 0 1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_21_409
timestamp 1608254825
transform 1 0 38732 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_399
timestamp 1608254825
transform 1 0 37812 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_393
timestamp 1608254825
transform 1 0 37260 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_4  _1768_
timestamp 1608254825
transform 1 0 37904 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_21_417
timestamp 1608254825
transform 1 0 39468 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1608254825
transform -1 0 39836 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_22_22
timestamp 1608254825
transform 1 0 3128 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1608254825
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _2421_
timestamp 1608254825
transform 1 0 1380 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_m1_clk_local
timestamp 1608254825
transform 1 0 3680 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_283
timestamp 1608254825
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2420_
timestamp 1608254825
transform 1 0 4048 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_22_51
timestamp 1608254825
transform 1 0 5796 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2475_
timestamp 1608254825
transform 1 0 6164 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_22_88
timestamp 1608254825
transform 1 0 9200 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_78
timestamp 1608254825
transform 1 0 8280 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_74
timestamp 1608254825
transform 1 0 7912 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_4  _2246_
timestamp 1608254825
transform 1 0 8372 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_22_107
timestamp 1608254825
transform 1 0 10948 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_284
timestamp 1608254825
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2471_
timestamp 1608254825
transform 1 0 11316 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__nand3_4  _2348_
timestamp 1608254825
transform 1 0 9660 0 -1 14688
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_22_130
timestamp 1608254825
transform 1 0 13064 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_4  _2268_
timestamp 1608254825
transform 1 0 13432 0 -1 14688
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_6  FILLER_22_147
timestamp 1608254825
transform 1 0 14628 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_285
timestamp 1608254825
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _2342_
timestamp 1608254825
transform 1 0 15272 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_22_177
timestamp 1608254825
transform 1 0 17388 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_170
timestamp 1608254825
transform 1 0 16744 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2169_
timestamp 1608254825
transform 1 0 17112 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_203
timestamp 1608254825
transform 1 0 19780 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_183
timestamp 1608254825
transform 1 0 17940 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2489_
timestamp 1608254825
transform 1 0 18032 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  FILLER_22_223
timestamp 1608254825
transform 1 0 21620 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_22_215
timestamp 1608254825
transform 1 0 20884 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_22_210
timestamp 1608254825
transform 1 0 20424 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_286
timestamp 1608254825
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2488_
timestamp 1608254825
transform 1 0 21896 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_2  _1947_
timestamp 1608254825
transform 1 0 20148 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_22_249
timestamp 1608254825
transform 1 0 24012 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_245
timestamp 1608254825
transform 1 0 23644 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2554_
timestamp 1608254825
transform 1 0 24104 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_22_269
timestamp 1608254825
transform 1 0 25852 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_289
timestamp 1608254825
transform 1 0 27692 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_283
timestamp 1608254825
transform 1 0 27140 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_287
timestamp 1608254825
transform 1 0 26404 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _1959_
timestamp 1608254825
transform 1 0 26496 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__nand4_4  _1707_
timestamp 1608254825
transform 1 0 27784 0 -1 14688
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_22_307
timestamp 1608254825
transform 1 0 29348 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_4  _1693_
timestamp 1608254825
transform 1 0 29716 0 -1 14688
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_22_341
timestamp 1608254825
transform 1 0 32476 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_332
timestamp 1608254825
transform 1 0 31648 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_324
timestamp 1608254825
transform 1 0 30912 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_288
timestamp 1608254825
transform 1 0 32016 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1677_
timestamp 1608254825
transform 1 0 31280 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1674_
timestamp 1608254825
transform 1 0 32108 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_349
timestamp 1608254825
transform 1 0 33212 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_345
timestamp 1608254825
transform 1 0 32844 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2655_
timestamp 1608254825
transform 1 0 33580 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_2  _1688_
timestamp 1608254825
transform 1 0 32936 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_372
timestamp 1608254825
transform 1 0 35328 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_4  _1621_
timestamp 1608254825
transform 1 0 35696 0 -1 14688
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_6  FILLER_22_411
timestamp 1608254825
transform 1 0 38916 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_22_389
timestamp 1608254825
transform 1 0 36892 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_289
timestamp 1608254825
transform 1 0 37628 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_4  _1769_
timestamp 1608254825
transform 1 0 37720 0 -1 14688
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_1  FILLER_22_417
timestamp 1608254825
transform 1 0 39468 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1608254825
transform -1 0 39836 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_23_3
timestamp 1608254825
transform 1 0 1380 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1608254825
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _2422_
timestamp 1608254825
transform 1 0 1656 0 1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_23_25
timestamp 1608254825
transform 1 0 3404 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2423_
timestamp 1608254825
transform 1 0 3772 0 1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_23_57
timestamp 1608254825
transform 1 0 6348 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_52
timestamp 1608254825
transform 1 0 5888 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_48
timestamp 1608254825
transform 1 0 5520 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_290
timestamp 1608254825
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2473_
timestamp 1608254825
transform 1 0 6808 0 1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  _2292_
timestamp 1608254825
transform 1 0 5980 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_81
timestamp 1608254825
transform 1 0 8556 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_4  _2349_
timestamp 1608254825
transform 1 0 8924 0 1 14688
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_23_113
timestamp 1608254825
transform 1 0 11500 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_98
timestamp 1608254825
transform 1 0 10120 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_4  _2220_
timestamp 1608254825
transform 1 0 10672 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_23_126
timestamp 1608254825
transform 1 0 12696 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_120
timestamp 1608254825
transform 1 0 12144 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_2_0_addressalyzerBlock.SPI_CLK
timestamp 1608254825
transform 1 0 11868 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_291
timestamp 1608254825
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_4  _2248_
timestamp 1608254825
transform 1 0 13064 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1887_
timestamp 1608254825
transform 1 0 12420 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_139
timestamp 1608254825
transform 1 0 13892 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2451_
timestamp 1608254825
transform 1 0 14260 0 1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_23_179
timestamp 1608254825
transform 1 0 17572 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_162
timestamp 1608254825
transform 1 0 16008 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_4  _2269_
timestamp 1608254825
transform 1 0 16376 0 1 14688
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_23_194
timestamp 1608254825
transform 1 0 18952 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_184
timestamp 1608254825
transform 1 0 18032 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_292
timestamp 1608254825
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _2272_
timestamp 1608254825
transform 1 0 18124 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__o32ai_4  _2130_
timestamp 1608254825
transform 1 0 19320 0 1 14688
box -38 -48 2062 592
use sky130_fd_sc_hd__decap_8  FILLER_23_227
timestamp 1608254825
transform 1 0 21988 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_23_220
timestamp 1608254825
transform 1 0 21344 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1953_
timestamp 1608254825
transform 1 0 21712 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_23_249
timestamp 1608254825
transform 1 0 24012 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_245
timestamp 1608254825
transform 1 0 23644 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_240
timestamp 1608254825
transform 1 0 23184 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_235
timestamp 1608254825
transform 1 0 22724 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_293
timestamp 1608254825
transform 1 0 23552 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2555_
timestamp 1608254825
transform 1 0 24104 0 1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_2  _1949_
timestamp 1608254825
transform 1 0 22908 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_269
timestamp 1608254825
transform 1 0 25852 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2648_
timestamp 1608254825
transform 1 0 26220 0 1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_23_292
timestamp 1608254825
transform 1 0 27968 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_306
timestamp 1608254825
transform 1 0 29256 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_304
timestamp 1608254825
transform 1 0 29072 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_294
timestamp 1608254825
transform 1 0 29164 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_4  _1745_
timestamp 1608254825
transform 1 0 29440 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_332
timestamp 1608254825
transform 1 0 31648 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_320
timestamp 1608254825
transform 1 0 30544 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1712_
timestamp 1608254825
transform 1 0 31280 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__nand4_4  _1683_
timestamp 1608254825
transform 1 0 32016 0 1 14688
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_6  FILLER_23_360
timestamp 1608254825
transform 1 0 34224 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_353
timestamp 1608254825
transform 1 0 33580 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2377_
timestamp 1608254825
transform 1 0 33948 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_23_385
timestamp 1608254825
transform 1 0 36524 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_23_367
timestamp 1608254825
transform 1 0 34868 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_295
timestamp 1608254825
transform 1 0 34776 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__a21o_4  _1617_
timestamp 1608254825
transform 1 0 35420 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_393
timestamp 1608254825
transform 1 0 37260 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _2646_
timestamp 1608254825
transform 1 0 37444 0 1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_23_414
timestamp 1608254825
transform 1 0 39192 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1608254825
transform -1 0 39836 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_24_22
timestamp 1608254825
transform 1 0 3128 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1608254825
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _2408_
timestamp 1608254825
transform 1 0 1380 0 -1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_24_30
timestamp 1608254825
transform 1 0 3864 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_296
timestamp 1608254825
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2424_
timestamp 1608254825
transform 1 0 4048 0 -1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_24_51
timestamp 1608254825
transform 1 0 5796 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2425_
timestamp 1608254825
transform 1 0 6164 0 -1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_24_90
timestamp 1608254825
transform 1 0 9384 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_82
timestamp 1608254825
transform 1 0 8648 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_24_74
timestamp 1608254825
transform 1 0 7912 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _2289_
timestamp 1608254825
transform 1 0 8280 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_107
timestamp 1608254825
transform 1 0 10948 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_97
timestamp 1608254825
transform 1 0 10028 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_93
timestamp 1608254825
transform 1 0 9660 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_297
timestamp 1608254825
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__o32ai_4  _2304_
timestamp 1608254825
transform 1 0 11316 0 -1 15776
box -38 -48 2062 592
use sky130_fd_sc_hd__nand2_4  _2222_
timestamp 1608254825
transform 1 0 10120 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_24_133
timestamp 1608254825
transform 1 0 13340 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_m1_clk_local
timestamp 1608254825
transform 1 0 13708 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_157
timestamp 1608254825
transform 1 0 15548 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_149
timestamp 1608254825
transform 1 0 14812 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_298
timestamp 1608254825
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _1901_
timestamp 1608254825
transform 1 0 13984 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1900_
timestamp 1608254825
transform 1 0 15272 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_24_164
timestamp 1608254825
transform 1 0 16192 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  _2447_
timestamp 1608254825
transform 1 0 16744 0 -1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_2  _1904_
timestamp 1608254825
transform 1 0 15916 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_189
timestamp 1608254825
transform 1 0 18492 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_4  _2350_
timestamp 1608254825
transform 1 0 18860 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_24_215
timestamp 1608254825
transform 1 0 20884 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_213
timestamp 1608254825
transform 1 0 20700 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_209
timestamp 1608254825
transform 1 0 20332 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_299
timestamp 1608254825
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__o32ai_4  _2132_
timestamp 1608254825
transform 1 0 21252 0 -1 15776
box -38 -48 2062 592
use sky130_fd_sc_hd__decap_4  FILLER_24_241
timestamp 1608254825
transform 1 0 23276 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_4  _1950_
timestamp 1608254825
transform 1 0 23644 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_24_274
timestamp 1608254825
transform 1 0 26312 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_266
timestamp 1608254825
transform 1 0 25576 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_24_254
timestamp 1608254825
transform 1 0 24472 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_283
timestamp 1608254825
transform 1 0 27140 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_300
timestamp 1608254825
transform 1 0 26404 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _1962_
timestamp 1608254825
transform 1 0 26496 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_4  _1698_
timestamp 1608254825
transform 1 0 27876 0 -1 15776
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_6  FILLER_24_304
timestamp 1608254825
transform 1 0 29072 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_4  _1727_
timestamp 1608254825
transform 1 0 29624 0 -1 15776
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_24_332
timestamp 1608254825
transform 1 0 31648 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_327
timestamp 1608254825
transform 1 0 31188 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_323
timestamp 1608254825
transform 1 0 30820 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_301
timestamp 1608254825
transform 1 0 32016 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_4  _1689_
timestamp 1608254825
transform 1 0 32108 0 -1 15776
box -38 -48 1234 592
use sky130_fd_sc_hd__buf_2  _1449_
timestamp 1608254825
transform 1 0 31280 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_359
timestamp 1608254825
transform 1 0 34132 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_350
timestamp 1608254825
transform 1 0 33304 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__or2_4  _2098_
timestamp 1608254825
transform 1 0 34500 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1675_
timestamp 1608254825
transform 1 0 33856 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_370
timestamp 1608254825
transform 1 0 35144 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2504_
timestamp 1608254825
transform 1 0 35512 0 -1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_24_401
timestamp 1608254825
transform 1 0 37996 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_393
timestamp 1608254825
transform 1 0 37260 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_302
timestamp 1608254825
transform 1 0 37628 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _2402_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 37720 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__and2_4  _2107_
timestamp 1608254825
transform 1 0 38364 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_24_412
timestamp 1608254825
transform 1 0 39008 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1608254825
transform -1 0 39836 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_25_19
timestamp 1608254825
transform 1 0 2852 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_15
timestamp 1608254825
transform 1 0 2484 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_3
timestamp 1608254825
transform 1 0 1380 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1608254825
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _2596_
timestamp 1608254825
transform 1 0 2944 0 1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_25_43
timestamp 1608254825
transform 1 0 5060 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_39
timestamp 1608254825
transform 1 0 4692 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_4  _1881_
timestamp 1608254825
transform 1 0 5152 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_25_53
timestamp 1608254825
transform 1 0 5980 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_303
timestamp 1608254825
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__o32ai_4  _2302_
timestamp 1608254825
transform 1 0 6808 0 1 15776
box -38 -48 2062 592
use sky130_fd_sc_hd__decap_6  FILLER_25_84
timestamp 1608254825
transform 1 0 8832 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  _2449_
timestamp 1608254825
transform 1 0 9384 0 1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_25_109
timestamp 1608254825
transform 1 0 11132 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1886_
timestamp 1608254825
transform 1 0 11500 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_135
timestamp 1608254825
transform 1 0 13524 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_25_123
timestamp 1608254825
transform 1 0 12420 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_25_121
timestamp 1608254825
transform 1 0 12236 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_117
timestamp 1608254825
transform 1 0 11868 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_304
timestamp 1608254825
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _1905_
timestamp 1608254825
transform 1 0 12696 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__o32ai_4  _2328_
timestamp 1608254825
transform 1 0 13892 0 1 15776
box -38 -48 2062 592
use sky130_fd_sc_hd__fill_2  FILLER_25_181
timestamp 1608254825
transform 1 0 17756 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_173
timestamp 1608254825
transform 1 0 17020 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_25_161
timestamp 1608254825
transform 1 0 15916 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1944_
timestamp 1608254825
transform 1 0 16652 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_198
timestamp 1608254825
transform 1 0 19320 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_194
timestamp 1608254825
transform 1 0 18952 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_187
timestamp 1608254825
transform 1 0 18308 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_305
timestamp 1608254825
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__o32ai_4  _2136_
timestamp 1608254825
transform 1 0 19412 0 1 15776
box -38 -48 2062 592
use sky130_fd_sc_hd__inv_2  _1977_
timestamp 1608254825
transform 1 0 18676 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1955_
timestamp 1608254825
transform 1 0 18032 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_25_221
timestamp 1608254825
transform 1 0 21436 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_25_240
timestamp 1608254825
transform 1 0 23184 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_229
timestamp 1608254825
transform 1 0 22172 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_306
timestamp 1608254825
transform 1 0 23552 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _1954_
timestamp 1608254825
transform 1 0 22356 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_4  _1952_
timestamp 1608254825
transform 1 0 23644 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_25_266
timestamp 1608254825
transform 1 0 25576 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_254
timestamp 1608254825
transform 1 0 24472 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__o21a_4  _1746_
timestamp 1608254825
transform 1 0 25760 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_296
timestamp 1608254825
transform 1 0 28336 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_25_280
timestamp 1608254825
transform 1 0 26864 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_4  _1744_
timestamp 1608254825
transform 1 0 27232 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_25_314
timestamp 1608254825
transform 1 0 29992 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_25_306
timestamp 1608254825
transform 1 0 29256 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_304
timestamp 1608254825
transform 1 0 29072 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_307
timestamp 1608254825
transform 1 0 29164 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2651_
timestamp 1608254825
transform 1 0 30268 0 1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_25_336
timestamp 1608254825
transform 1 0 32016 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1448_
timestamp 1608254825
transform 1 0 32384 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_362
timestamp 1608254825
transform 1 0 34408 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_347
timestamp 1608254825
transform 1 0 33028 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_343
timestamp 1608254825
transform 1 0 32660 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_4  _2369_
timestamp 1608254825
transform 1 0 33120 0 1 15776
box -38 -48 1326 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_308
timestamp 1608254825
transform 1 0 34776 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__o41ai_4  _2370_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 34868 0 1 15776
box -38 -48 2062 592
use sky130_fd_sc_hd__decap_4  FILLER_25_389
timestamp 1608254825
transform 1 0 36892 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2505_
timestamp 1608254825
transform 1 0 37260 0 1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_25_412
timestamp 1608254825
transform 1 0 39008 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1608254825
transform -1 0 39836 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_22
timestamp 1608254825
transform 1 0 3128 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_18
timestamp 1608254825
transform 1 0 2760 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_11
timestamp 1608254825
transform 1 0 2116 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_3
timestamp 1608254825
transform 1 0 1380 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_6_0_m1_clk_local
timestamp 1608254825
transform 1 0 2484 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1608254825
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1608254825
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _2588_
timestamp 1608254825
transform 1 0 1380 0 1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  _2405_
timestamp 1608254825
transform 1 0 1748 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_45
timestamp 1608254825
transform 1 0 5244 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_43
timestamp 1608254825
transform 1 0 5060 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_39
timestamp 1608254825
transform 1 0 4692 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_30
timestamp 1608254825
transform 1 0 3864 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_309
timestamp 1608254825
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2594_
timestamp 1608254825
transform 1 0 3496 0 1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__and2_4  _1891_
timestamp 1608254825
transform 1 0 4048 0 -1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_4  _1877_
timestamp 1608254825
transform 1 0 5152 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_27_56
timestamp 1608254825
transform 1 0 6256 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_53
timestamp 1608254825
transform 1 0 5980 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_m1_clk_local
timestamp 1608254825
transform 1 0 6348 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__and2_4  _1893_
timestamp 1608254825
transform 1 0 5612 0 1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_27_66
timestamp 1608254825
transform 1 0 7176 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_62
timestamp 1608254825
transform 1 0 6808 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_60
timestamp 1608254825
transform 1 0 6624 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_316
timestamp 1608254825
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _1879_
timestamp 1608254825
transform 1 0 6624 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_4  _2595_
timestamp 1608254825
transform 1 0 7268 0 1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_27_86
timestamp 1608254825
transform 1 0 9016 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_88
timestamp 1608254825
transform 1 0 9200 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_69
timestamp 1608254825
transform 1 0 7452 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_4  _2347_
timestamp 1608254825
transform 1 0 8004 0 -1 16864
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_1  FILLER_27_100
timestamp 1608254825
transform 1 0 10304 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_96
timestamp 1608254825
transform 1 0 9936 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_310
timestamp 1608254825
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _1885_
timestamp 1608254825
transform 1 0 10396 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _1874_
timestamp 1608254825
transform 1 0 9568 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_110
timestamp 1608254825
transform 1 0 11224 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_107
timestamp 1608254825
transform 1 0 10948 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1875_
timestamp 1608254825
transform 1 0 11592 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1425_
timestamp 1608254825
transform 1 0 11316 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_4  _2346_
timestamp 1608254825
transform 1 0 9660 0 -1 16864
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_27_118
timestamp 1608254825
transform 1 0 11960 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_115
timestamp 1608254825
transform 1 0 11684 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_317
timestamp 1608254825
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2472_
timestamp 1608254825
transform 1 0 12420 0 1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _2457_
timestamp 1608254825
transform 1 0 12420 0 -1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_27_142
timestamp 1608254825
transform 1 0 14168 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_158
timestamp 1608254825
transform 1 0 15640 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_149
timestamp 1608254825
transform 1 0 14812 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_142
timestamp 1608254825
transform 1 0 14168 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_311
timestamp 1608254825
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2567_
timestamp 1608254825
transform 1 0 14720 0 1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  _1938_
timestamp 1608254825
transform 1 0 15272 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1884_
timestamp 1608254825
transform 1 0 14536 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_179
timestamp 1608254825
transform 1 0 17572 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_175
timestamp 1608254825
transform 1 0 17204 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_167
timestamp 1608254825
transform 1 0 16468 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_166
timestamp 1608254825
transform 1 0 16376 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2485_
timestamp 1608254825
transform 1 0 16744 0 -1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  _1957_
timestamp 1608254825
transform 1 0 16008 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1210_
timestamp 1608254825
transform 1 0 17296 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_27_193
timestamp 1608254825
transform 1 0 18860 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_26_200
timestamp 1608254825
transform 1 0 19504 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp 1608254825
transform 1 0 19044 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_189
timestamp 1608254825
transform 1 0 18492 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_318
timestamp 1608254825
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__o32ai_4  _2128_
timestamp 1608254825
transform 1 0 19412 0 1 16864
box -38 -48 2062 592
use sky130_fd_sc_hd__buf_2  _2127_
timestamp 1608254825
transform 1 0 19136 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_4  _1946_
timestamp 1608254825
transform 1 0 18032 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_27_221
timestamp 1608254825
transform 1 0 21436 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_215
timestamp 1608254825
transform 1 0 20884 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_210
timestamp 1608254825
transform 1 0 20424 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_206
timestamp 1608254825
transform 1 0 20056 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_312
timestamp 1608254825
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__o32ai_4  _2134_
timestamp 1608254825
transform 1 0 20976 0 -1 16864
box -38 -48 2062 592
use sky130_fd_sc_hd__buf_2  _2123_
timestamp 1608254825
transform 1 0 21988 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1945_
timestamp 1608254825
transform 1 0 20148 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_27_235
timestamp 1608254825
transform 1 0 22724 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_231
timestamp 1608254825
transform 1 0 22356 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_238
timestamp 1608254825
transform 1 0 23000 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1776_
timestamp 1608254825
transform 1 0 22816 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_245
timestamp 1608254825
transform 1 0 23644 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_240
timestamp 1608254825
transform 1 0 23184 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_245
timestamp 1608254825
transform 1 0 23644 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_319
timestamp 1608254825
transform 1 0 23552 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1951_
timestamp 1608254825
transform 1 0 23368 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _2553_
timestamp 1608254825
transform 1 0 24012 0 1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _2552_
timestamp 1608254825
transform 1 0 24012 0 -1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_27_268
timestamp 1608254825
transform 1 0 25760 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_274
timestamp 1608254825
transform 1 0 26312 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_268
timestamp 1608254825
transform 1 0 25760 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__and2_4  _1961_
timestamp 1608254825
transform 1 0 26128 0 1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_27_295
timestamp 1608254825
transform 1 0 28244 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_285
timestamp 1608254825
transform 1 0 27324 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_279
timestamp 1608254825
transform 1 0 26772 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_313
timestamp 1608254825
transform 1 0 26404 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__a41oi_4  _1743_
timestamp 1608254825
transform 1 0 26496 0 -1 16864
box -38 -48 2062 592
use sky130_fd_sc_hd__and4_4  _1713_
timestamp 1608254825
transform 1 0 27416 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_27_311
timestamp 1608254825
transform 1 0 29716 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_306
timestamp 1608254825
transform 1 0 29256 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_303
timestamp 1608254825
transform 1 0 28980 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_298
timestamp 1608254825
transform 1 0 28520 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_320
timestamp 1608254825
transform 1 0 29164 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2654_
timestamp 1608254825
transform 1 0 28888 0 -1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__a41oi_4  _1728_
timestamp 1608254825
transform 1 0 30084 0 1 16864
box -38 -48 2062 592
use sky130_fd_sc_hd__inv_2  _1673_
timestamp 1608254825
transform 1 0 29440 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_27_337
timestamp 1608254825
transform 1 0 32108 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_341
timestamp 1608254825
transform 1 0 32476 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_335
timestamp 1608254825
transform 1 0 31924 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_329
timestamp 1608254825
transform 1 0 31372 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_321
timestamp 1608254825
transform 1 0 30636 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_314
timestamp 1608254825
transform 1 0 32016 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1714_
timestamp 1608254825
transform 1 0 31004 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1488_
timestamp 1608254825
transform 1 0 32108 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_362
timestamp 1608254825
transform 1 0 34408 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_349
timestamp 1608254825
transform 1 0 33212 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_345
timestamp 1608254825
transform 1 0 32844 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_350
timestamp 1608254825
transform 1 0 33304 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_345
timestamp 1608254825
transform 1 0 32844 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2431_
timestamp 1608254825
transform 1 0 33672 0 -1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  _1722_
timestamp 1608254825
transform 1 0 32936 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1619_
timestamp 1608254825
transform 1 0 32936 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_4  _1611_
timestamp 1608254825
transform 1 0 33580 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_27_370
timestamp 1608254825
transform 1 0 35144 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_385
timestamp 1608254825
transform 1 0 36524 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_381
timestamp 1608254825
transform 1 0 36156 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_373
timestamp 1608254825
transform 1 0 35420 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_321
timestamp 1608254825
transform 1 0 34776 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _2097_
timestamp 1608254825
transform 1 0 36616 0 -1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__nor4_4  _2093_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 35512 0 1 16864
box -38 -48 1602 592
use sky130_fd_sc_hd__inv_2  _1613_
timestamp 1608254825
transform 1 0 34868 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1492_
timestamp 1608254825
transform 1 0 35788 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_391
timestamp 1608254825
transform 1 0 37076 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_408
timestamp 1608254825
transform 1 0 38640 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_398
timestamp 1608254825
transform 1 0 37720 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_393
timestamp 1608254825
transform 1 0 37260 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_315
timestamp 1608254825
transform 1 0 37628 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2506_
timestamp 1608254825
transform 1 0 37444 0 1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__and4_4  _2095_
timestamp 1608254825
transform 1 0 37812 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_27_414
timestamp 1608254825
transform 1 0 39192 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_416
timestamp 1608254825
transform 1 0 39376 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1608254825
transform -1 0 39836 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1608254825
transform -1 0 39836 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_28_22
timestamp 1608254825
transform 1 0 3128 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1608254825
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _2590_
timestamp 1608254825
transform 1 0 1380 0 -1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_28_40
timestamp 1608254825
transform 1 0 4784 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_32
timestamp 1608254825
transform 1 0 4048 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_30
timestamp 1608254825
transform 1 0 3864 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_322
timestamp 1608254825
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _1883_
timestamp 1608254825
transform 1 0 4876 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_28_50
timestamp 1608254825
transform 1 0 5704 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2427_
timestamp 1608254825
transform 1 0 6072 0 -1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_28_91
timestamp 1608254825
transform 1 0 9476 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_83
timestamp 1608254825
transform 1 0 8740 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_28_73
timestamp 1608254825
transform 1 0 7820 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _1292_
timestamp 1608254825
transform 1 0 8372 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_108
timestamp 1608254825
transform 1 0 11040 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_100
timestamp 1608254825
transform 1 0 10304 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_323
timestamp 1608254825
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__o32ai_4  _2303_
timestamp 1608254825
transform 1 0 11224 0 -1 17952
box -38 -48 2062 592
use sky130_fd_sc_hd__and2_4  _1892_
timestamp 1608254825
transform 1 0 9660 0 -1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_28_132
timestamp 1608254825
transform 1 0 13248 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_158
timestamp 1608254825
transform 1 0 15640 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_154
timestamp 1608254825
transform 1 0 15272 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_149
timestamp 1608254825
transform 1 0 14812 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_140
timestamp 1608254825
transform 1 0 13984 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_324
timestamp 1608254825
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _1958_
timestamp 1608254825
transform 1 0 14168 0 -1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _1941_
timestamp 1608254825
transform 1 0 15732 0 -1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_28_166
timestamp 1608254825
transform 1 0 16376 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__o32ai_4  _2138_
timestamp 1608254825
transform 1 0 17112 0 -1 17952
box -38 -48 2062 592
use sky130_fd_sc_hd__decap_4  FILLER_28_196
timestamp 1608254825
transform 1 0 19136 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_4  _2126_
timestamp 1608254825
transform 1 0 19504 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_28_215
timestamp 1608254825
transform 1 0 20884 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_213
timestamp 1608254825
transform 1 0 20700 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_209
timestamp 1608254825
transform 1 0 20332 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_325
timestamp 1608254825
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2487_
timestamp 1608254825
transform 1 0 21436 0 -1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_28_240
timestamp 1608254825
transform 1 0 23184 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2495_
timestamp 1608254825
transform 1 0 23552 0 -1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_28_271
timestamp 1608254825
transform 1 0 26036 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_263
timestamp 1608254825
transform 1 0 25300 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1521_
timestamp 1608254825
transform 1 0 25668 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_294
timestamp 1608254825
transform 1 0 28152 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_288
timestamp 1608254825
transform 1 0 27600 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_326
timestamp 1608254825
transform 1 0 26404 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__a41oi_4  _1699_
timestamp 1608254825
transform 1 0 28244 0 -1 17952
box -38 -48 2062 592
use sky130_fd_sc_hd__a21o_4  _1519_
timestamp 1608254825
transform 1 0 26496 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_317
timestamp 1608254825
transform 1 0 30268 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_28_337
timestamp 1608254825
transform 1 0 32108 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_332
timestamp 1608254825
transform 1 0 31648 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_327
timestamp 1608254825
transform 1 0 32016 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2433_
timestamp 1608254825
transform 1 0 32292 0 -1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__nand2_4  _1726_
timestamp 1608254825
transform 1 0 30820 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_28_358
timestamp 1608254825
transform 1 0 34040 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_4  _1610_
timestamp 1608254825
transform 1 0 34408 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_383
timestamp 1608254825
transform 1 0 36340 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_378
timestamp 1608254825
transform 1 0 35880 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_374
timestamp 1608254825
transform 1 0 35512 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1451_
timestamp 1608254825
transform 1 0 36708 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1244_
timestamp 1608254825
transform 1 0 35972 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_407
timestamp 1608254825
transform 1 0 38548 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_391
timestamp 1608254825
transform 1 0 37076 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_328
timestamp 1608254825
transform 1 0 37628 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _2094_
timestamp 1608254825
transform 1 0 38916 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_4  _2084_
timestamp 1608254825
transform 1 0 37720 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_28_414
timestamp 1608254825
transform 1 0 39192 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1608254825
transform -1 0 39836 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_29_19
timestamp 1608254825
transform 1 0 2852 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_15
timestamp 1608254825
transform 1 0 2484 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_3
timestamp 1608254825
transform 1 0 1380 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1608254825
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_4  _2081_
timestamp 1608254825
transform 1 0 2944 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_36
timestamp 1608254825
transform 1 0 4416 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_32
timestamp 1608254825
transform 1 0 4048 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2593_
timestamp 1608254825
transform 1 0 4508 0 1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_29_68
timestamp 1608254825
transform 1 0 7360 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_29_62
timestamp 1608254825
transform 1 0 6808 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_29_60
timestamp 1608254825
transform 1 0 6624 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_56
timestamp 1608254825
transform 1 0 6256 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_329
timestamp 1608254825
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1882_
timestamp 1608254825
transform 1 0 7084 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_91
timestamp 1608254825
transform 1 0 9476 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2428_
timestamp 1608254825
transform 1 0 7728 0 1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_29_114
timestamp 1608254825
transform 1 0 11592 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _2572_
timestamp 1608254825
transform 1 0 9844 0 1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_29_130
timestamp 1608254825
transform 1 0 13064 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_330
timestamp 1608254825
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _1895_
timestamp 1608254825
transform 1 0 12420 0 1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_29_157
timestamp 1608254825
transform 1 0 15548 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2556_
timestamp 1608254825
transform 1 0 13800 0 1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_29_179
timestamp 1608254825
transform 1 0 17572 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_166
timestamp 1608254825
transform 1 0 16376 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_161
timestamp 1608254825
transform 1 0 15916 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__and3_4  _2307_
timestamp 1608254825
transform 1 0 16744 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _1241_
timestamp 1608254825
transform 1 0 16008 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_194
timestamp 1608254825
transform 1 0 18952 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_184
timestamp 1608254825
transform 1 0 18032 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_331
timestamp 1608254825
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2490_
timestamp 1608254825
transform 1 0 19320 0 1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  _1516_
timestamp 1608254825
transform 1 0 18584 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_217
timestamp 1608254825
transform 1 0 21068 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_4  _2110_
timestamp 1608254825
transform 1 0 21436 0 1 17952
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_1  FILLER_29_249
timestamp 1608254825
transform 1 0 24012 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_245
timestamp 1608254825
transform 1 0 23644 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_242
timestamp 1608254825
transform 1 0 23368 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_234
timestamp 1608254825
transform 1 0 22632 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_332
timestamp 1608254825
transform 1 0 23552 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__o32a_4  _1518_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 24104 0 1 17952
box -38 -48 1694 592
use sky130_fd_sc_hd__fill_1  FILLER_29_274
timestamp 1608254825
transform 1 0 26312 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_268
timestamp 1608254825
transform 1 0 25760 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_296
timestamp 1608254825
transform 1 0 28336 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_292
timestamp 1608254825
transform 1 0 27968 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__a22oi_4  _1473_
timestamp 1608254825
transform 1 0 26404 0 1 17952
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_6  FILLER_29_315
timestamp 1608254825
transform 1 0 30084 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_301
timestamp 1608254825
transform 1 0 28796 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_333
timestamp 1608254825
transform 1 0 29164 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_4  _1694_
timestamp 1608254825
transform 1 0 29256 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _1211_
timestamp 1608254825
transform 1 0 28428 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_338
timestamp 1608254825
transform 1 0 32200 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_334
timestamp 1608254825
transform 1 0 31832 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_12_0_addressalyzerBlock.SPI_CLK
timestamp 1608254825
transform 1 0 32292 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_4  _2379_
timestamp 1608254825
transform 1 0 32568 0 1 17952
box -38 -48 1234 592
use sky130_fd_sc_hd__a21oi_4  _1685_
timestamp 1608254825
transform 1 0 30636 0 1 17952
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_29_362
timestamp 1608254825
transform 1 0 34408 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_355
timestamp 1608254825
transform 1 0 33764 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1607_
timestamp 1608254825
transform 1 0 34132 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_386
timestamp 1608254825
transform 1 0 36616 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_367
timestamp 1608254825
transform 1 0 34868 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_334
timestamp 1608254825
transform 1 0 34776 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__nand4_4  _1615_
timestamp 1608254825
transform 1 0 35052 0 1 17952
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_1  FILLER_29_393
timestamp 1608254825
transform 1 0 37260 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_13_0_addressalyzerBlock.SPI_CLK
timestamp 1608254825
transform 1 0 36984 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _2514_
timestamp 1608254825
transform 1 0 37352 0 1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_29_417
timestamp 1608254825
transform 1 0 39468 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_413
timestamp 1608254825
transform 1 0 39100 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1608254825
transform -1 0 39836 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_30_22
timestamp 1608254825
transform 1 0 3128 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1608254825
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _2587_
timestamp 1608254825
transform 1 0 1380 0 -1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_30_35
timestamp 1608254825
transform 1 0 4324 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_30
timestamp 1608254825
transform 1 0 3864 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_335
timestamp 1608254825
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _2075_
timestamp 1608254825
transform 1 0 4048 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__and2_4  _1894_
timestamp 1608254825
transform 1 0 5060 0 -1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_30_61
timestamp 1608254825
transform 1 0 6716 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_57
timestamp 1608254825
transform 1 0 6348 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_50
timestamp 1608254825
transform 1 0 5704 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_7_0_m1_clk_local
timestamp 1608254825
transform 1 0 6072 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _2407_
timestamp 1608254825
transform 1 0 6808 0 -1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_30_88
timestamp 1608254825
transform 1 0 9200 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_81
timestamp 1608254825
transform 1 0 8556 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1273_
timestamp 1608254825
transform 1 0 8924 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_96
timestamp 1608254825
transform 1 0 9936 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_336
timestamp 1608254825
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2592_
timestamp 1608254825
transform 1 0 10304 0 -1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_2  _2291_
timestamp 1608254825
transform 1 0 9660 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_119
timestamp 1608254825
transform 1 0 12052 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2494_
timestamp 1608254825
transform 1 0 12420 0 -1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_30_149
timestamp 1608254825
transform 1 0 14812 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_142
timestamp 1608254825
transform 1 0 14168 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_337
timestamp 1608254825
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2493_
timestamp 1608254825
transform 1 0 15272 0 -1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_2  _2288_
timestamp 1608254825
transform 1 0 14536 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_30_179
timestamp 1608254825
transform 1 0 17572 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_173
timestamp 1608254825
transform 1 0 17020 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__nor4_4  _2331_
timestamp 1608254825
transform 1 0 17664 0 -1 19040
box -38 -48 1602 592
use sky130_fd_sc_hd__and4_4  _2290_
timestamp 1608254825
transform 1 0 19596 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _1630_
timestamp 1608254825
transform 1 0 19228 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_228
timestamp 1608254825
transform 1 0 22080 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_210
timestamp 1608254825
transform 1 0 20424 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_338
timestamp 1608254825
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_4  _1537_
timestamp 1608254825
transform 1 0 20884 0 -1 19040
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_1  FILLER_30_242
timestamp 1608254825
transform 1 0 23368 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_236
timestamp 1608254825
transform 1 0 22816 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _2124_
timestamp 1608254825
transform 1 0 22448 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_4  _2108_
timestamp 1608254825
transform 1 0 23460 0 -1 19040
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_30_271
timestamp 1608254825
transform 1 0 26036 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_263
timestamp 1608254825
transform 1 0 25300 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_256
timestamp 1608254825
transform 1 0 24656 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2385_
timestamp 1608254825
transform 1 0 25024 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1696_
timestamp 1608254825
transform 1 0 25668 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_293
timestamp 1608254825
transform 1 0 28060 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_339
timestamp 1608254825
transform 1 0 26404 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__a22oi_4  _1482_
timestamp 1608254825
transform 1 0 26496 0 -1 19040
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_30_300
timestamp 1608254825
transform 1 0 28704 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2544_
timestamp 1608254825
transform 1 0 29072 0 -1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_2  _1470_
timestamp 1608254825
transform 1 0 28428 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_30_335
timestamp 1608254825
transform 1 0 31924 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_331
timestamp 1608254825
transform 1 0 31556 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_323
timestamp 1608254825
transform 1 0 30820 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_340
timestamp 1608254825
transform 1 0 32016 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1469_
timestamp 1608254825
transform 1 0 31188 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_4  _1454_
timestamp 1608254825
transform 1 0 32108 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_30_363
timestamp 1608254825
transform 1 0 34500 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_350
timestamp 1608254825
transform 1 0 33304 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_346
timestamp 1608254825
transform 1 0 32936 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_addressalyzerBlock.SPI_CLK
timestamp 1608254825
transform 1 0 33396 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_4  _1608_
timestamp 1608254825
transform 1 0 33672 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_30_385
timestamp 1608254825
transform 1 0 36524 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_367
timestamp 1608254825
transform 1 0 34868 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__nand4_4  _1620_
timestamp 1608254825
transform 1 0 34960 0 -1 19040
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_30_407
timestamp 1608254825
transform 1 0 38548 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_393
timestamp 1608254825
transform 1 0 37260 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_341
timestamp 1608254825
transform 1 0 37628 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _1748_
timestamp 1608254825
transform 1 0 37720 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1614_
timestamp 1608254825
transform 1 0 38916 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1243_
timestamp 1608254825
transform 1 0 36892 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_414
timestamp 1608254825
transform 1 0 39192 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1608254825
transform -1 0 39836 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_14
timestamp 1608254825
transform 1 0 2392 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_3
timestamp 1608254825
transform 1 0 1380 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1608254825
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _2516_
timestamp 1608254825
transform 1 0 2760 0 1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__and3_4  _2079_
timestamp 1608254825
transform 1 0 1564 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_31_37
timestamp 1608254825
transform 1 0 4508 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_60
timestamp 1608254825
transform 1 0 6624 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_56
timestamp 1608254825
transform 1 0 6256 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_31_49
timestamp 1608254825
transform 1 0 5612 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_342
timestamp 1608254825
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _2082_
timestamp 1608254825
transform 1 0 6808 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _2073_
timestamp 1608254825
transform 1 0 5888 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_91
timestamp 1608254825
transform 1 0 9476 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_83
timestamp 1608254825
transform 1 0 8740 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_31_71
timestamp 1608254825
transform 1 0 7636 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1408_
timestamp 1608254825
transform 1 0 8372 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_109
timestamp 1608254825
transform 1 0 11132 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_101
timestamp 1608254825
transform 1 0 10396 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_97
timestamp 1608254825
transform 1 0 10028 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__and2_4  _1935_
timestamp 1608254825
transform 1 0 10488 0 1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _1890_
timestamp 1608254825
transform 1 0 11500 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1889_
timestamp 1608254825
transform 1 0 9660 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_121
timestamp 1608254825
transform 1 0 12236 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_117
timestamp 1608254825
transform 1 0 11868 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_343
timestamp 1608254825
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2571_
timestamp 1608254825
transform 1 0 12420 0 1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_31_158
timestamp 1608254825
transform 1 0 15640 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_150
timestamp 1608254825
transform 1 0 14904 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_142
timestamp 1608254825
transform 1 0 14168 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__and2_4  _1914_
timestamp 1608254825
transform 1 0 14996 0 1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_31_179
timestamp 1608254825
transform 1 0 17572 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__a41o_4  _2305_
timestamp 1608254825
transform 1 0 16008 0 1 19040
box -38 -48 1602 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_344
timestamp 1608254825
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__a41o_4  _2351_
timestamp 1608254825
transform 1 0 18860 0 1 19040
box -38 -48 1602 592
use sky130_fd_sc_hd__nor2_4  _2287_
timestamp 1608254825
transform 1 0 18032 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_31_223
timestamp 1608254825
transform 1 0 21620 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__a21oi_4  _2109_
timestamp 1608254825
transform 1 0 20424 0 1 19040
box -38 -48 1234 592
use sky130_fd_sc_hd__o22a_4  _1524_
timestamp 1608254825
transform 1 0 21804 0 1 19040
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_1  FILLER_31_243
timestamp 1608254825
transform 1 0 23460 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_239
timestamp 1608254825
transform 1 0 23092 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_345
timestamp 1608254825
transform 1 0 23552 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_4  _1520_
timestamp 1608254825
transform 1 0 23644 0 1 19040
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_2  FILLER_31_266
timestamp 1608254825
transform 1 0 25576 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_258
timestamp 1608254825
transform 1 0 24840 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__a22oi_4  _1503_
timestamp 1608254825
transform 1 0 25760 0 1 19040
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_1  FILLER_31_291
timestamp 1608254825
transform 1 0 27876 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_285
timestamp 1608254825
transform 1 0 27324 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_4  _1964_
timestamp 1608254825
transform 1 0 27968 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_31_319
timestamp 1608254825
transform 1 0 30452 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_31_301
timestamp 1608254825
transform 1 0 28796 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_346
timestamp 1608254825
transform 1 0 29164 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_4  _1453_
timestamp 1608254825
transform 1 0 29256 0 1 19040
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_31_341
timestamp 1608254825
transform 1 0 32476 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_4  _1456_
timestamp 1608254825
transform 1 0 31188 0 1 19040
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_31_362
timestamp 1608254825
transform 1 0 34408 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_355
timestamp 1608254825
transform 1 0 33764 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_345
timestamp 1608254825
transform 1 0 32844 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_4  _2378_
timestamp 1608254825
transform 1 0 32936 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1205_
timestamp 1608254825
transform 1 0 34132 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_378
timestamp 1608254825
transform 1 0 35880 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_371
timestamp 1608254825
transform 1 0 35236 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_347
timestamp 1608254825
transform 1 0 34776 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _2375_
timestamp 1608254825
transform 1 0 36248 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1612_
timestamp 1608254825
transform 1 0 35604 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1239_
timestamp 1608254825
transform 1 0 34868 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_391
timestamp 1608254825
transform 1 0 37076 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2434_
timestamp 1608254825
transform 1 0 37444 0 1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_31_414
timestamp 1608254825
transform 1 0 39192 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1608254825
transform -1 0 39836 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_11
timestamp 1608254825
transform 1 0 2116 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_3
timestamp 1608254825
transform 1 0 1380 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1608254825
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_4  _2074_
timestamp 1608254825
transform 1 0 2300 0 -1 20128
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_32_45
timestamp 1608254825
transform 1 0 5244 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_27
timestamp 1608254825
transform 1 0 3588 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_348
timestamp 1608254825
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_4  _2080_
timestamp 1608254825
transform 1 0 4048 0 -1 20128
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_1  FILLER_32_49
timestamp 1608254825
transform 1 0 5612 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2426_
timestamp 1608254825
transform 1 0 5704 0 -1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_32_88
timestamp 1608254825
transform 1 0 9200 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_75
timestamp 1608254825
transform 1 0 8004 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_69
timestamp 1608254825
transform 1 0 7452 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_4  _1436_
timestamp 1608254825
transform 1 0 8096 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_112
timestamp 1608254825
transform 1 0 11408 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_108
timestamp 1608254825
transform 1 0 11040 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_100
timestamp 1608254825
transform 1 0 10304 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_32_93
timestamp 1608254825
transform 1 0 9660 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_349
timestamp 1608254825
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2670_
timestamp 1608254825
transform 1 0 11500 0 -1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  _1896_
timestamp 1608254825
transform 1 0 10672 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1426_
timestamp 1608254825
transform 1 0 9936 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_132
timestamp 1608254825
transform 1 0 13248 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_32_158
timestamp 1608254825
transform 1 0 15640 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_152
timestamp 1608254825
transform 1 0 15088 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_148
timestamp 1608254825
transform 1 0 14720 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_140
timestamp 1608254825
transform 1 0 13984 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_350
timestamp 1608254825
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _1936_
timestamp 1608254825
transform 1 0 14076 0 -1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _1915_
timestamp 1608254825
transform 1 0 15272 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_162
timestamp 1608254825
transform 1 0 16008 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__a41o_4  _2293_
timestamp 1608254825
transform 1 0 16100 0 -1 20128
box -38 -48 1602 592
use sky130_fd_sc_hd__buf_2  _1242_
timestamp 1608254825
transform 1 0 17664 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_201
timestamp 1608254825
transform 1 0 19596 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__a41o_4  _2341_
timestamp 1608254825
transform 1 0 18032 0 -1 20128
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_1  FILLER_32_225
timestamp 1608254825
transform 1 0 21804 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_219
timestamp 1608254825
transform 1 0 21252 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_32_211
timestamp 1608254825
transform 1 0 20516 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_351
timestamp 1608254825
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1631_
timestamp 1608254825
transform 1 0 20884 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1629_
timestamp 1608254825
transform 1 0 20148 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_4  _1533_
timestamp 1608254825
transform 1 0 21896 0 -1 20128
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_6  FILLER_32_240
timestamp 1608254825
transform 1 0 23184 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_4  _1513_
timestamp 1608254825
transform 1 0 23736 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_271
timestamp 1608254825
transform 1 0 26036 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_266
timestamp 1608254825
transform 1 0 25576 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_258
timestamp 1608254825
transform 1 0 24840 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1440_
timestamp 1608254825
transform 1 0 25760 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_32_295
timestamp 1608254825
transform 1 0 28244 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_32_276
timestamp 1608254825
transform 1 0 26496 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_352
timestamp 1608254825
transform 1 0 26404 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_4  _1480_
timestamp 1608254825
transform 1 0 27048 0 -1 20128
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_32_317
timestamp 1608254825
transform 1 0 30268 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_303
timestamp 1608254825
transform 1 0 28980 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_4  _1509_
timestamp 1608254825
transform 1 0 29072 0 -1 20128
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_6  FILLER_32_330
timestamp 1608254825
transform 1 0 31464 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_353
timestamp 1608254825
transform 1 0 32016 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_4  _1618_
timestamp 1608254825
transform 1 0 30636 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__and2_4  _1457_
timestamp 1608254825
transform 1 0 32108 0 -1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_32_348
timestamp 1608254825
transform 1 0 33120 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_344
timestamp 1608254825
transform 1 0 32752 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__o32ai_4  _2380_
timestamp 1608254825
transform 1 0 33212 0 -1 20128
box -38 -48 2062 592
use sky130_fd_sc_hd__fill_1  FILLER_32_375
timestamp 1608254825
transform 1 0 35604 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_371
timestamp 1608254825
transform 1 0 35236 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__a22oi_4  _2374_
timestamp 1608254825
transform 1 0 35696 0 -1 20128
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_32_393
timestamp 1608254825
transform 1 0 37260 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_354
timestamp 1608254825
transform 1 0 37628 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__a211o_4  _2383_
timestamp 1608254825
transform 1 0 37720 0 -1 20128
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_6  FILLER_32_412
timestamp 1608254825
transform 1 0 39008 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1608254825
transform -1 0 39836 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_11
timestamp 1608254825
transform 1 0 2116 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_7
timestamp 1608254825
transform 1 0 1748 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_3
timestamp 1608254825
transform 1 0 1380 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_22
timestamp 1608254825
transform 1 0 3128 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1608254825
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1608254825
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _2517_
timestamp 1608254825
transform 1 0 1380 0 1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__a21o_4  _2078_
timestamp 1608254825
transform 1 0 2484 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _2065_
timestamp 1608254825
transform 1 0 1840 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_34_32
timestamp 1608254825
transform 1 0 4048 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_27
timestamp 1608254825
transform 1 0 3588 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_34
timestamp 1608254825
transform 1 0 4232 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_26
timestamp 1608254825
transform 1 0 3496 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_361
timestamp 1608254825
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2518_
timestamp 1608254825
transform 1 0 4600 0 1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__and3_4  _2077_
timestamp 1608254825
transform 1 0 4600 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__or2_4  _2076_
timestamp 1608254825
transform 1 0 3588 0 1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_34_47
timestamp 1608254825
transform 1 0 5428 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_62
timestamp 1608254825
transform 1 0 6808 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_57
timestamp 1608254825
transform 1 0 6348 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_355
timestamp 1608254825
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2515_
timestamp 1608254825
transform 1 0 5796 0 -1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_34_88
timestamp 1608254825
transform 1 0 9200 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_74
timestamp 1608254825
transform 1 0 7912 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_70
timestamp 1608254825
transform 1 0 7544 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2669_
timestamp 1608254825
transform 1 0 7912 0 1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__a21oi_4  _1435_
timestamp 1608254825
transform 1 0 8004 0 -1 21216
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_33_111
timestamp 1608254825
transform 1 0 11316 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_93
timestamp 1608254825
transform 1 0 9660 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_362
timestamp 1608254825
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__nand3_4  _1432_
timestamp 1608254825
transform 1 0 10028 0 1 20128
box -38 -48 1326 592
use sky130_fd_sc_hd__a41oi_4  _1427_
timestamp 1608254825
transform 1 0 9660 0 -1 21216
box -38 -48 2062 592
use sky130_fd_sc_hd__decap_8  FILLER_34_115
timestamp 1608254825
transform 1 0 11684 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_33_135
timestamp 1608254825
transform 1 0 13524 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_118
timestamp 1608254825
transform 1 0 11960 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_356
timestamp 1608254825
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1434_
timestamp 1608254825
transform 1 0 11684 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_4  _1431_
timestamp 1608254825
transform 1 0 12420 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__nand4_4  _1253_
timestamp 1608254825
transform 1 0 12420 0 -1 21216
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_6  FILLER_34_157
timestamp 1608254825
transform 1 0 15548 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_152
timestamp 1608254825
transform 1 0 15088 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_148
timestamp 1608254825
transform 1 0 14720 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_140
timestamp 1608254825
transform 1 0 13984 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_158
timestamp 1608254825
transform 1 0 15640 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_363
timestamp 1608254825
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2581_
timestamp 1608254825
transform 1 0 13892 0 1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_2  _1421_
timestamp 1608254825
transform 1 0 15272 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1413_
timestamp 1608254825
transform 1 0 14352 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_181
timestamp 1608254825
transform 1 0 17756 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_163
timestamp 1608254825
transform 1 0 16100 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_179
timestamp 1608254825
transform 1 0 17572 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_169
timestamp 1608254825
transform 1 0 16652 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__a41o_4  _2321_
timestamp 1608254825
transform 1 0 16192 0 -1 21216
box -38 -48 1602 592
use sky130_fd_sc_hd__buf_2  _2115_
timestamp 1608254825
transform 1 0 17204 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__and2_4  _1912_
timestamp 1608254825
transform 1 0 16008 0 1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_34_200
timestamp 1608254825
transform 1 0 19504 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_34_194
timestamp 1608254825
transform 1 0 18952 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_33_196
timestamp 1608254825
transform 1 0 19136 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_33_184
timestamp 1608254825
transform 1 0 18032 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_m1_clk_local $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 19412 0 1 20128
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_357
timestamp 1608254825
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__and4_4  _2353_
timestamp 1608254825
transform 1 0 19596 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_4  _1978_
timestamp 1608254825
transform 1 0 18124 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_34_215
timestamp 1608254825
transform 1 0 20884 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_210
timestamp 1608254825
transform 1 0 20424 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_219
timestamp 1608254825
transform 1 0 21252 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_addressalyzerBlock.SPI_CLK
timestamp 1608254825
transform 1 0 21620 0 1 20128
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_364
timestamp 1608254825
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_4  _1529_
timestamp 1608254825
transform 1 0 21068 0 -1 21216
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_2  FILLER_34_230
timestamp 1608254825
transform 1 0 22264 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_243
timestamp 1608254825
transform 1 0 23460 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_358
timestamp 1608254825
transform 1 0 23552 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _1976_
timestamp 1608254825
transform 1 0 22448 0 -1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_4  _1491_
timestamp 1608254825
transform 1 0 23736 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__o32ai_4  _1490_
timestamp 1608254825
transform 1 0 23644 0 1 20128
box -38 -48 2062 592
use sky130_fd_sc_hd__buf_2  _1474_
timestamp 1608254825
transform 1 0 23092 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1441_
timestamp 1608254825
transform 1 0 23460 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_271
timestamp 1608254825
transform 1 0 26036 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_255
timestamp 1608254825
transform 1 0 24564 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_267
timestamp 1608254825
transform 1 0 25668 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_4  _1483_
timestamp 1608254825
transform 1 0 24932 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_283
timestamp 1608254825
transform 1 0 27140 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_34_276
timestamp 1608254825
transform 1 0 26496 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_294
timestamp 1608254825
transform 1 0 28152 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_365
timestamp 1608254825
transform 1 0 26404 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2666_
timestamp 1608254825
transform 1 0 26404 0 1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__a21oi_4  _1479_
timestamp 1608254825
transform 1 0 27508 0 -1 21216
box -38 -48 1234 592
use sky130_fd_sc_hd__buf_2  _1458_
timestamp 1608254825
transform 1 0 26772 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_300
timestamp 1608254825
transform 1 0 28704 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_33_306
timestamp 1608254825
transform 1 0 29256 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_301
timestamp 1608254825
transform 1 0 28796 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_359
timestamp 1608254825
transform 1 0 29164 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__and4_4  _1676_
timestamp 1608254825
transform 1 0 29072 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1485_
timestamp 1608254825
transform 1 0 28520 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_34_319
timestamp 1608254825
transform 1 0 30452 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_34_313
timestamp 1608254825
transform 1 0 29900 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_313
timestamp 1608254825
transform 1 0 29900 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1472_
timestamp 1608254825
transform 1 0 29532 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_4  _1627_
timestamp 1608254825
transform 1 0 30268 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_34_337
timestamp 1608254825
transform 1 0 32108 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_332
timestamp 1608254825
transform 1 0 31648 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_324
timestamp 1608254825
transform 1 0 30912 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_333
timestamp 1608254825
transform 1 0 31740 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_366
timestamp 1608254825
transform 1 0 32016 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1471_
timestamp 1608254825
transform 1 0 30544 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_4  _1455_
timestamp 1608254825
transform 1 0 32108 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _1447_
timestamp 1608254825
transform 1 0 31280 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1206_
timestamp 1608254825
transform 1 0 32384 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_344
timestamp 1608254825
transform 1 0 32752 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_362
timestamp 1608254825
transform 1 0 34408 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_349
timestamp 1608254825
transform 1 0 33212 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2432_
timestamp 1608254825
transform 1 0 33120 0 -1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__nor2_4  _1446_
timestamp 1608254825
transform 1 0 33580 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_34_373
timestamp 1608254825
transform 1 0 35420 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_34_367
timestamp 1608254825
transform 1 0 34868 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_33_376
timestamp 1608254825
transform 1 0 35696 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_360
timestamp 1608254825
transform 1 0 34776 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2509_
timestamp 1608254825
transform 1 0 35512 0 -1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _2429_
timestamp 1608254825
transform 1 0 36432 0 1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__nor2_4  _1609_
timestamp 1608254825
transform 1 0 34868 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_34_393
timestamp 1608254825
transform 1 0 37260 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_410
timestamp 1608254825
transform 1 0 38824 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_33_403
timestamp 1608254825
transform 1 0 38180 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_367
timestamp 1608254825
transform 1 0 37628 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__nand3_4  _2381_
timestamp 1608254825
transform 1 0 37720 0 -1 21216
box -38 -48 1326 592
use sky130_fd_sc_hd__inv_2  _1828_
timestamp 1608254825
transform 1 0 38548 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_34_412
timestamp 1608254825
transform 1 0 39008 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1608254825
transform -1 0 39836 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1608254825
transform -1 0 39836 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_35_22
timestamp 1608254825
transform 1 0 3128 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1608254825
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _2521_
timestamp 1608254825
transform 1 0 1380 0 1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_35_30
timestamp 1608254825
transform 1 0 3864 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__nand4_4  _1986_
timestamp 1608254825
transform 1 0 3956 0 1 21216
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_1  FILLER_35_60
timestamp 1608254825
transform 1 0 6624 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_56
timestamp 1608254825
transform 1 0 6256 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_48
timestamp 1608254825
transform 1 0 5520 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_368
timestamp 1608254825
transform 1 0 6716 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_4  _2072_
timestamp 1608254825
transform 1 0 6808 0 1 21216
box -38 -48 1234 592
use sky130_fd_sc_hd__buf_2  _2054_
timestamp 1608254825
transform 1 0 5888 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_87
timestamp 1608254825
transform 1 0 9108 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_75
timestamp 1608254825
transform 1 0 8004 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_99
timestamp 1608254825
transform 1 0 10212 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__nand3_4  _1433_
timestamp 1608254825
transform 1 0 10396 0 1 21216
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_1  FILLER_35_123
timestamp 1608254825
transform 1 0 12420 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_35_121
timestamp 1608254825
transform 1 0 12236 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_115
timestamp 1608254825
transform 1 0 11684 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_369
timestamp 1608254825
transform 1 0 12328 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__nand3_4  _1414_
timestamp 1608254825
transform 1 0 12512 0 1 21216
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_35_138
timestamp 1608254825
transform 1 0 13800 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2583_
timestamp 1608254825
transform 1 0 14168 0 1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_35_182
timestamp 1608254825
transform 1 0 17848 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_174
timestamp 1608254825
transform 1 0 17112 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_35_161
timestamp 1608254825
transform 1 0 15916 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_4  _2318_
timestamp 1608254825
transform 1 0 16284 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_35_187
timestamp 1608254825
transform 1 0 18308 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_370
timestamp 1608254825
transform 1 0 17940 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2538_
timestamp 1608254825
transform 1 0 18860 0 1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_2  _2157_
timestamp 1608254825
transform 1 0 18032 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_212
timestamp 1608254825
transform 1 0 20608 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_4  _1536_
timestamp 1608254825
transform 1 0 22080 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__a21o_4  _1528_
timestamp 1608254825
transform 1 0 20976 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_243
timestamp 1608254825
transform 1 0 23460 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_371
timestamp 1608254825
transform 1 0 23552 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2665_
timestamp 1608254825
transform 1 0 23644 0 1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_2  _2319_
timestamp 1608254825
transform 1 0 23184 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_35_264
timestamp 1608254825
transform 1 0 25392 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_4  _1484_
timestamp 1608254825
transform 1 0 26128 0 1 21216
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_35_285
timestamp 1608254825
transform 1 0 27324 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_4  _1477_
timestamp 1608254825
transform 1 0 27692 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_35_304
timestamp 1608254825
transform 1 0 29072 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_298
timestamp 1608254825
transform 1 0 28520 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_372
timestamp 1608254825
transform 1 0 29164 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2658_
timestamp 1608254825
transform 1 0 29256 0 1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_35_342
timestamp 1608254825
transform 1 0 32568 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_325
timestamp 1608254825
transform 1 0 31004 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_4  _1634_
timestamp 1608254825
transform 1 0 31372 0 1 21216
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_35_362
timestamp 1608254825
transform 1 0 34408 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_346
timestamp 1608254825
transform 1 0 32936 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_addressalyzerBlock.SPI_CLK
timestamp 1608254825
transform 1 0 33028 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_4  _2372_
timestamp 1608254825
transform 1 0 33304 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_373
timestamp 1608254825
transform 1 0 34776 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__o32ai_4  _2373_
timestamp 1608254825
transform 1 0 34868 0 1 21216
box -38 -48 2062 592
use sky130_fd_sc_hd__decap_6  FILLER_35_389
timestamp 1608254825
transform 1 0 36892 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  _2508_
timestamp 1608254825
transform 1 0 37444 0 1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_35_414
timestamp 1608254825
transform 1 0 39192 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1608254825
transform -1 0 39836 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_7
timestamp 1608254825
transform 1 0 1748 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1608254825
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_4  _2064_
timestamp 1608254825
transform 1 0 2116 0 -1 22304
box -38 -48 1234 592
use sky130_fd_sc_hd__buf_2  _2053_
timestamp 1608254825
transform 1 0 1380 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_43
timestamp 1608254825
transform 1 0 5060 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_32
timestamp 1608254825
transform 1 0 4048 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_36_30
timestamp 1608254825
transform 1 0 3864 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_24
timestamp 1608254825
transform 1 0 3312 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_374
timestamp 1608254825
transform 1 0 3956 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _2055_
timestamp 1608254825
transform 1 0 4232 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_4  _2519_
timestamp 1608254825
transform 1 0 5796 0 -1 22304
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_36_88
timestamp 1608254825
transform 1 0 9200 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_74
timestamp 1608254825
transform 1 0 7912 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_70
timestamp 1608254825
transform 1 0 7544 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_4  _1428_
timestamp 1608254825
transform 1 0 8004 0 -1 22304
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_8  FILLER_36_114
timestamp 1608254825
transform 1 0 11592 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_36_106
timestamp 1608254825
transform 1 0 10856 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_102
timestamp 1608254825
transform 1 0 10488 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_96
timestamp 1608254825
transform 1 0 9936 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_375
timestamp 1608254825
transform 1 0 9568 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1424_
timestamp 1608254825
transform 1 0 9660 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1416_
timestamp 1608254825
transform 1 0 11224 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1251_
timestamp 1608254825
transform 1 0 10580 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_136
timestamp 1608254825
transform 1 0 13616 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_4  _1420_
timestamp 1608254825
transform 1 0 12328 0 -1 22304
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_6  FILLER_36_157
timestamp 1608254825
transform 1 0 15548 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_36_147
timestamp 1608254825
transform 1 0 14628 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_376
timestamp 1608254825
transform 1 0 15180 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _1429_
timestamp 1608254825
transform 1 0 13984 0 -1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1415_
timestamp 1608254825
transform 1 0 15272 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_180
timestamp 1608254825
transform 1 0 17664 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__a2111o_4  _2280_
timestamp 1608254825
transform 1 0 16100 0 -1 22304
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_36_202
timestamp 1608254825
transform 1 0 19688 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_184
timestamp 1608254825
transform 1 0 18032 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__nand4_4  _2114_
timestamp 1608254825
transform 1 0 18124 0 -1 22304
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_36_210
timestamp 1608254825
transform 1 0 20424 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_377
timestamp 1608254825
transform 1 0 20792 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2661_
timestamp 1608254825
transform 1 0 20884 0 -1 22304
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  _2112_
timestamp 1608254825
transform 1 0 20056 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_242
timestamp 1608254825
transform 1 0 23368 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_234
timestamp 1608254825
transform 1 0 22632 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_4  _1493_
timestamp 1608254825
transform 1 0 23552 0 -1 22304
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_36_271
timestamp 1608254825
transform 1 0 26036 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_261
timestamp 1608254825
transform 1 0 25116 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_257
timestamp 1608254825
transform 1 0 24748 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_4  _1541_
timestamp 1608254825
transform 1 0 25208 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_36_295
timestamp 1608254825
transform 1 0 28244 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_36_276
timestamp 1608254825
transform 1 0 26496 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_378
timestamp 1608254825
transform 1 0 26404 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__nor4_4  _1703_
timestamp 1608254825
transform 1 0 26680 0 -1 22304
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_36_315
timestamp 1608254825
transform 1 0 30084 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_301
timestamp 1608254825
transform 1 0 28796 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__nor3_4  _2384_
timestamp 1608254825
transform 1 0 28888 0 -1 22304
box -38 -48 1234 592
use sky130_fd_sc_hd__o21ai_4  _1628_
timestamp 1608254825
transform 1 0 30452 0 -1 22304
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_2  FILLER_36_337
timestamp 1608254825
transform 1 0 32108 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_332
timestamp 1608254825
transform 1 0 31648 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_379
timestamp 1608254825
transform 1 0 32016 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1478_
timestamp 1608254825
transform 1 0 32292 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_360
timestamp 1608254825
transform 1 0 34224 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_36_343
timestamp 1608254825
transform 1 0 32660 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_4  _1665_
timestamp 1608254825
transform 1 0 33028 0 -1 22304
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_2  FILLER_36_368
timestamp 1608254825
transform 1 0 34960 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _2430_
timestamp 1608254825
transform 1 0 35144 0 -1 22304
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_36_411
timestamp 1608254825
transform 1 0 38916 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_36_389
timestamp 1608254825
transform 1 0 36892 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_380
timestamp 1608254825
transform 1 0 37628 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__nor3_4  _2092_
timestamp 1608254825
transform 1 0 37720 0 -1 22304
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_1  FILLER_36_417
timestamp 1608254825
transform 1 0 39468 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1608254825
transform -1 0 39836 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_22
timestamp 1608254825
transform 1 0 3128 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_3
timestamp 1608254825
transform 1 0 1380 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1608254825
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_4  _2063_
timestamp 1608254825
transform 1 0 1932 0 1 22304
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_37_43
timestamp 1608254825
transform 1 0 5060 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__nor4_4  _1987_
timestamp 1608254825
transform 1 0 3496 0 1 22304
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_37_57
timestamp 1608254825
transform 1 0 6348 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_47
timestamp 1608254825
transform 1 0 5428 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_381
timestamp 1608254825
transform 1 0 6716 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _2067_
timestamp 1608254825
transform 1 0 5520 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  _1985_
timestamp 1608254825
transform 1 0 6808 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_37_71
timestamp 1608254825
transform 1 0 7636 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2672_
timestamp 1608254825
transform 1 0 8004 0 1 22304
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_37_94
timestamp 1608254825
transform 1 0 9752 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2673_
timestamp 1608254825
transform 1 0 10120 0 1 22304
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_37_132
timestamp 1608254825
transform 1 0 13248 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_121
timestamp 1608254825
transform 1 0 12236 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_117
timestamp 1608254825
transform 1 0 11868 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_382
timestamp 1608254825
transform 1 0 12328 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _1418_
timestamp 1608254825
transform 1 0 12420 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_37_157
timestamp 1608254825
transform 1 0 15548 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2674_
timestamp 1608254825
transform 1 0 13800 0 1 22304
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_37_179
timestamp 1608254825
transform 1 0 17572 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_161
timestamp 1608254825
transform 1 0 15916 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__a2111o_4  _2185_
timestamp 1608254825
transform 1 0 16008 0 1 22304
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_1  FILLER_37_202
timestamp 1608254825
transform 1 0 19688 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_37_196
timestamp 1608254825
transform 1 0 19136 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_37_188
timestamp 1608254825
transform 1 0 18400 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_383
timestamp 1608254825
transform 1 0 17940 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_4  _2151_
timestamp 1608254825
transform 1 0 19780 0 1 22304
box -38 -48 1234 592
use sky130_fd_sc_hd__buf_2  _1656_
timestamp 1608254825
transform 1 0 18032 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1512_
timestamp 1608254825
transform 1 0 18768 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_216
timestamp 1608254825
transform 1 0 20976 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2662_
timestamp 1608254825
transform 1 0 21344 0 1 22304
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_37_249
timestamp 1608254825
transform 1 0 24012 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_243
timestamp 1608254825
transform 1 0 23460 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_239
timestamp 1608254825
transform 1 0 23092 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_384
timestamp 1608254825
transform 1 0 23552 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1461_
timestamp 1608254825
transform 1 0 23644 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_265
timestamp 1608254825
transform 1 0 25484 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_4  _1487_
timestamp 1608254825
transform 1 0 24380 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__o41a_4  _1462_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 25852 0 1 22304
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_6  FILLER_37_296
timestamp 1608254825
transform 1 0 28336 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_37_286
timestamp 1608254825
transform 1 0 27416 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _1445_
timestamp 1608254825
transform 1 0 27968 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_37_306
timestamp 1608254825
transform 1 0 29256 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_14_0_addressalyzerBlock.SPI_CLK
timestamp 1608254825
transform 1 0 28888 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_385
timestamp 1608254825
transform 1 0 29164 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2437_
timestamp 1608254825
transform 1 0 29532 0 1 22304
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_37_328
timestamp 1608254825
transform 1 0 31280 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__nand4_4  _1633_
timestamp 1608254825
transform 1 0 31648 0 1 22304
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_1  FILLER_37_365
timestamp 1608254825
transform 1 0 34684 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_357
timestamp 1608254825
transform 1 0 33948 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_37_349
timestamp 1608254825
transform 1 0 33212 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1506_
timestamp 1608254825
transform 1 0 33580 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_387
timestamp 1608254825
transform 1 0 36708 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_377
timestamp 1608254825
transform 1 0 35788 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_37_371
timestamp 1608254825
transform 1 0 35236 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_386
timestamp 1608254825
transform 1 0 34776 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__and3_4  _2382_
timestamp 1608254825
transform 1 0 35880 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _1507_
timestamp 1608254825
transform 1 0 34868 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_409
timestamp 1608254825
transform 1 0 38732 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_399
timestamp 1608254825
transform 1 0 37812 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_395
timestamp 1608254825
transform 1 0 37444 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _2091_
timestamp 1608254825
transform 1 0 37076 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__and3_4  _2090_
timestamp 1608254825
transform 1 0 37904 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_37_417
timestamp 1608254825
transform 1 0 39468 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1608254825
transform -1 0 39836 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_38_3
timestamp 1608254825
transform 1 0 1380 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1608254825
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _2522_
timestamp 1608254825
transform 1 0 1472 0 -1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_38_45
timestamp 1608254825
transform 1 0 5244 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_23
timestamp 1608254825
transform 1 0 3220 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_387
timestamp 1608254825
transform 1 0 3956 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__nor3_4  _2048_
timestamp 1608254825
transform 1 0 4048 0 -1 23392
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_38_62
timestamp 1608254825
transform 1 0 6808 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_4  _2071_
timestamp 1608254825
transform 1 0 5612 0 -1 23392
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _2066_
timestamp 1608254825
transform 1 0 7176 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_38_91
timestamp 1608254825
transform 1 0 9476 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_85
timestamp 1608254825
transform 1 0 8924 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_38_77
timestamp 1608254825
transform 1 0 8188 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_69
timestamp 1608254825
transform 1 0 7452 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1299_
timestamp 1608254825
transform 1 0 7820 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1298_
timestamp 1608254825
transform 1 0 8556 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_112
timestamp 1608254825
transform 1 0 11408 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_106
timestamp 1608254825
transform 1 0 10856 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_388
timestamp 1608254825
transform 1 0 9568 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_4  _1422_
timestamp 1608254825
transform 1 0 9660 0 -1 23392
box -38 -48 1234 592
use sky130_fd_sc_hd__nand3_4  _1419_
timestamp 1608254825
transform 1 0 11500 0 -1 23392
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_38_127
timestamp 1608254825
transform 1 0 12788 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__a41o_4  _1417_
timestamp 1608254825
transform 1 0 13156 0 -1 23392
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_38_159
timestamp 1608254825
transform 1 0 15732 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_154
timestamp 1608254825
transform 1 0 15272 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_38_152
timestamp 1608254825
transform 1 0 15088 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_148
timestamp 1608254825
transform 1 0 14720 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_389
timestamp 1608254825
transform 1 0 15180 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _2158_
timestamp 1608254825
transform 1 0 15364 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_180
timestamp 1608254825
transform 1 0 17664 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__a2111o_4  _2159_
timestamp 1608254825
transform 1 0 16100 0 -1 23392
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_38_203
timestamp 1608254825
transform 1 0 19780 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__a2111o_4  _2210_
timestamp 1608254825
transform 1 0 18216 0 -1 23392
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_38_226
timestamp 1608254825
transform 1 0 21896 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_215
timestamp 1608254825
transform 1 0 20884 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_210
timestamp 1608254825
transform 1 0 20424 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_390
timestamp 1608254825
transform 1 0 20792 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _1538_
timestamp 1608254825
transform 1 0 21068 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1534_
timestamp 1608254825
transform 1 0 20148 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_233
timestamp 1608254825
transform 1 0 22540 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2663_
timestamp 1608254825
transform 1 0 22908 0 -1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_2  _1525_
timestamp 1608254825
transform 1 0 22264 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_271
timestamp 1608254825
transform 1 0 26036 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_256
timestamp 1608254825
transform 1 0 24656 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_4  _1486_
timestamp 1608254825
transform 1 0 25208 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_38_289
timestamp 1608254825
transform 1 0 27692 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_391
timestamp 1608254825
transform 1 0 26404 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_4  _1476_
timestamp 1608254825
transform 1 0 28060 0 -1 23392
box -38 -48 1234 592
use sky130_fd_sc_hd__nor3_4  _1444_
timestamp 1608254825
transform 1 0 26496 0 -1 23392
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_1  FILLER_38_312
timestamp 1608254825
transform 1 0 29808 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_306
timestamp 1608254825
transform 1 0 29256 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_4  _1623_
timestamp 1608254825
transform 1 0 29900 0 -1 23392
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_1  FILLER_38_332
timestamp 1608254825
transform 1 0 31648 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_326
timestamp 1608254825
transform 1 0 31096 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_addressalyzerBlock.SPI_CLK
timestamp 1608254825
transform 1 0 31740 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_392
timestamp 1608254825
transform 1 0 32016 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__nor3_4  _1625_
timestamp 1608254825
transform 1 0 32108 0 -1 23392
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_2  FILLER_38_357
timestamp 1608254825
transform 1 0 33948 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_350
timestamp 1608254825
transform 1 0 33304 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_15_0_addressalyzerBlock.SPI_CLK
timestamp 1608254825
transform 1 0 33672 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_4  _2376_
timestamp 1608254825
transform 1 0 34132 0 -1 23392
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_38_373
timestamp 1608254825
transform 1 0 35420 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_4  _2366_
timestamp 1608254825
transform 1 0 35788 0 -1 23392
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_38_407
timestamp 1608254825
transform 1 0 38548 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_396
timestamp 1608254825
transform 1 0 37536 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_390
timestamp 1608254825
transform 1 0 36984 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_393
timestamp 1608254825
transform 1 0 37628 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _2371_
timestamp 1608254825
transform 1 0 38916 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_4  _2105_
timestamp 1608254825
transform 1 0 37720 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_38_414
timestamp 1608254825
transform 1 0 39192 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1608254825
transform -1 0 39836 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_20
timestamp 1608254825
transform 1 0 2944 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_3
timestamp 1608254825
transform 1 0 1380 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_3
timestamp 1608254825
transform 1 0 1380 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1608254825
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1608254825
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_4  _2062_
timestamp 1608254825
transform 1 0 1748 0 -1 24480
box -38 -48 1234 592
use sky130_fd_sc_hd__a21oi_4  _2061_
timestamp 1608254825
transform 1 0 2484 0 1 23392
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_40_27
timestamp 1608254825
transform 1 0 3588 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_28
timestamp 1608254825
transform 1 0 3680 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_400
timestamp 1608254825
transform 1 0 3956 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _2049_
timestamp 1608254825
transform 1 0 4048 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1984_
timestamp 1608254825
transform 1 0 4048 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1983_
timestamp 1608254825
transform 1 0 3312 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_40_41
timestamp 1608254825
transform 1 0 4876 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_40_35
timestamp 1608254825
transform 1 0 4324 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_44
timestamp 1608254825
transform 1 0 5152 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_36
timestamp 1608254825
transform 1 0 4416 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _2520_
timestamp 1608254825
transform 1 0 4968 0 -1 24480
box -38 -48 1786 592
use sky130_fd_sc_hd__a21o_4  _2069_
timestamp 1608254825
transform 1 0 5244 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_68
timestamp 1608254825
transform 1 0 7360 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_40_61
timestamp 1608254825
transform 1 0 6716 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_62
timestamp 1608254825
transform 1 0 6808 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_39_57
timestamp 1608254825
transform 1 0 6348 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_394
timestamp 1608254825
transform 1 0 6716 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _2070_
timestamp 1608254825
transform 1 0 7084 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_88
timestamp 1608254825
transform 1 0 9200 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_74
timestamp 1608254825
transform 1 0 7912 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_39_82
timestamp 1608254825
transform 1 0 8648 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_74
timestamp 1608254825
transform 1 0 7912 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_4  _1423_
timestamp 1608254825
transform 1 0 8740 0 1 23392
box -38 -48 1234 592
use sky130_fd_sc_hd__nor3_4  _1412_
timestamp 1608254825
transform 1 0 8004 0 -1 24480
box -38 -48 1234 592
use sky130_fd_sc_hd__buf_2  _1405_
timestamp 1608254825
transform 1 0 7544 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_102
timestamp 1608254825
transform 1 0 10488 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_104
timestamp 1608254825
transform 1 0 10672 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_96
timestamp 1608254825
transform 1 0 9936 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_401
timestamp 1608254825
transform 1 0 9568 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _1411_
timestamp 1608254825
transform 1 0 9660 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__nor3_4  _1380_
timestamp 1608254825
transform 1 0 10764 0 1 23392
box -38 -48 1234 592
use sky130_fd_sc_hd__nor4_4  _1254_
timestamp 1608254825
transform 1 0 10856 0 -1 24480
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_2  FILLER_40_131
timestamp 1608254825
transform 1 0 13156 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_40_123
timestamp 1608254825
transform 1 0 12420 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_39_132
timestamp 1608254825
transform 1 0 13248 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_39_118
timestamp 1608254825
transform 1 0 11960 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_395
timestamp 1608254825
transform 1 0 12328 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_4  _1392_
timestamp 1608254825
transform 1 0 13340 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  _1252_
timestamp 1608254825
transform 1 0 12420 0 1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_40_157
timestamp 1608254825
transform 1 0 15548 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_149
timestamp 1608254825
transform 1 0 14812 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_142
timestamp 1608254825
transform 1 0 14168 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_159
timestamp 1608254825
transform 1 0 15732 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_402
timestamp 1608254825
transform 1 0 15180 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2671_
timestamp 1608254825
transform 1 0 13984 0 1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_2  _1393_
timestamp 1608254825
transform 1 0 15272 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1250_
timestamp 1608254825
transform 1 0 14536 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_179
timestamp 1608254825
transform 1 0 17572 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_172
timestamp 1608254825
transform 1 0 16928 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__a2111oi_4  _1660_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 15916 0 -1 24480
box -38 -48 2062 592
use sky130_fd_sc_hd__and3_4  _1430_
timestamp 1608254825
transform 1 0 16100 0 1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1395_
timestamp 1608254825
transform 1 0 17296 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_40_204
timestamp 1608254825
transform 1 0 19872 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_40_183
timestamp 1608254825
transform 1 0 17940 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_204
timestamp 1608254825
transform 1 0 19872 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_39_184
timestamp 1608254825
transform 1 0 18032 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_396
timestamp 1608254825
transform 1 0 17940 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__a2111o_4  _2258_
timestamp 1608254825
transform 1 0 18308 0 -1 24480
box -38 -48 1602 592
use sky130_fd_sc_hd__a2111o_4  _2234_
timestamp 1608254825
transform 1 0 18308 0 1 23392
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_1  FILLER_40_223
timestamp 1608254825
transform 1 0 21620 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_219
timestamp 1608254825
transform 1 0 21252 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_212
timestamp 1608254825
transform 1 0 20608 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_217
timestamp 1608254825
transform 1 0 21068 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_403
timestamp 1608254825
transform 1 0 20792 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__nand3_4  _1598_
timestamp 1608254825
transform 1 0 21712 0 -1 24480
box -38 -48 1326 592
use sky130_fd_sc_hd__nor2_4  _1523_
timestamp 1608254825
transform 1 0 21436 0 1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  _1508_
timestamp 1608254825
transform 1 0 20240 0 1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _1497_
timestamp 1608254825
transform 1 0 20884 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_238
timestamp 1608254825
transform 1 0 23000 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_238
timestamp 1608254825
transform 1 0 23000 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_230
timestamp 1608254825
transform 1 0 22264 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_397
timestamp 1608254825
transform 1 0 23552 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__nor3_4  _1571_
timestamp 1608254825
transform 1 0 23368 0 -1 24480
box -38 -48 1234 592
use sky130_fd_sc_hd__nand4_4  _1443_
timestamp 1608254825
transform 1 0 23644 0 1 23392
box -38 -48 1602 592
use sky130_fd_sc_hd__buf_2  _1442_
timestamp 1608254825
transform 1 0 22632 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_271
timestamp 1608254825
transform 1 0 26036 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_255
timestamp 1608254825
transform 1 0 24564 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_266
timestamp 1608254825
transform 1 0 25576 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_262
timestamp 1608254825
transform 1 0 25208 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_4  _1475_
timestamp 1608254825
transform 1 0 24932 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__o21ai_4  _1467_
timestamp 1608254825
transform 1 0 25668 0 1 23392
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_40_285
timestamp 1608254825
transform 1 0 27324 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_276
timestamp 1608254825
transform 1 0 26496 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_280
timestamp 1608254825
transform 1 0 26864 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_404
timestamp 1608254825
transform 1 0 26404 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_4  _1466_
timestamp 1608254825
transform 1 0 27692 0 -1 24480
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _1460_
timestamp 1608254825
transform 1 0 27048 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__nand4_4  _1450_
timestamp 1608254825
transform 1 0 27232 0 1 23392
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_8  FILLER_40_302
timestamp 1608254825
transform 1 0 28888 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_306
timestamp 1608254825
transform 1 0 29256 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_301
timestamp 1608254825
transform 1 0 28796 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_398
timestamp 1608254825
transform 1 0 29164 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_310
timestamp 1608254825
transform 1 0 29624 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_319
timestamp 1608254825
transform 1 0 30452 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_312
timestamp 1608254825
transform 1 0 29808 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1624_
timestamp 1608254825
transform 1 0 29532 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1622_
timestamp 1608254825
transform 1 0 30176 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _2438_
timestamp 1608254825
transform 1 0 29808 0 -1 24480
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_40_337
timestamp 1608254825
transform 1 0 32108 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_335
timestamp 1608254825
transform 1 0 31924 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_331
timestamp 1608254825
transform 1 0 31556 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_335
timestamp 1608254825
transform 1 0 31924 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_405
timestamp 1608254825
transform 1 0 32016 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_4  _2367_
timestamp 1608254825
transform 1 0 30820 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__a211o_4  _1666_
timestamp 1608254825
transform 1 0 32292 0 1 23392
box -38 -48 1326 592
use sky130_fd_sc_hd__nor3_4  _1664_
timestamp 1608254825
transform 1 0 32292 0 -1 24480
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_1  FILLER_40_356
timestamp 1608254825
transform 1 0 33856 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_352
timestamp 1608254825
transform 1 0 33488 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_365
timestamp 1608254825
transform 1 0 34684 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_361
timestamp 1608254825
transform 1 0 34316 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_353
timestamp 1608254825
transform 1 0 33580 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2435_
timestamp 1608254825
transform 1 0 33948 0 -1 24480
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  _1668_
timestamp 1608254825
transform 1 0 33948 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_376
timestamp 1608254825
transform 1 0 35696 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_388
timestamp 1608254825
transform 1 0 36800 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_39_367
timestamp 1608254825
transform 1 0 34868 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_399
timestamp 1608254825
transform 1 0 34776 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2436_
timestamp 1608254825
transform 1 0 35052 0 1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__nand2_4  _2365_
timestamp 1608254825
transform 1 0 36064 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_40_407
timestamp 1608254825
transform 1 0 38548 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_389
timestamp 1608254825
transform 1 0 36892 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_394
timestamp 1608254825
transform 1 0 37352 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_406
timestamp 1608254825
transform 1 0 37628 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2498_
timestamp 1608254825
transform 1 0 37444 0 1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__nand2_4  _2104_
timestamp 1608254825
transform 1 0 37720 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _2089_
timestamp 1608254825
transform 1 0 38916 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_414
timestamp 1608254825
transform 1 0 39192 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_414
timestamp 1608254825
transform 1 0 39192 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1608254825
transform -1 0 39836 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1608254825
transform -1 0 39836 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_41_11
timestamp 1608254825
transform 1 0 2116 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_3
timestamp 1608254825
transform 1 0 1380 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1608254825
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__a41oi_4  _2056_
timestamp 1608254825
transform 1 0 2208 0 1 24480
box -38 -48 2062 592
use sky130_fd_sc_hd__fill_2  FILLER_41_42
timestamp 1608254825
transform 1 0 4968 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_41_34
timestamp 1608254825
transform 1 0 4232 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_4  _2068_
timestamp 1608254825
transform 1 0 5152 0 1 24480
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_41_57
timestamp 1608254825
transform 1 0 6348 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_407
timestamp 1608254825
transform 1 0 6716 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__nor3_4  _1407_
timestamp 1608254825
transform 1 0 6808 0 1 24480
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_1  FILLER_41_79
timestamp 1608254825
transform 1 0 8372 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_75
timestamp 1608254825
transform 1 0 8004 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2675_
timestamp 1608254825
transform 1 0 8464 0 1 24480
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_41_112
timestamp 1608254825
transform 1 0 11408 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_41_99
timestamp 1608254825
transform 1 0 10212 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__and4_4  _1399_
timestamp 1608254825
transform 1 0 10580 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_41_132
timestamp 1608254825
transform 1 0 13248 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_120
timestamp 1608254825
transform 1 0 12144 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_408
timestamp 1608254825
transform 1 0 12328 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__and4_4  _1389_
timestamp 1608254825
transform 1 0 12420 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_41_159
timestamp 1608254825
transform 1 0 15732 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _2680_
timestamp 1608254825
transform 1 0 13984 0 1 24480
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_41_181
timestamp 1608254825
transform 1 0 17756 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_41_173
timestamp 1608254825
transform 1 0 17020 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_167
timestamp 1608254825
transform 1 0 16468 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _1588_
timestamp 1608254825
transform 1 0 16652 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_203
timestamp 1608254825
transform 1 0 19780 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_198
timestamp 1608254825
transform 1 0 19320 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_194
timestamp 1608254825
transform 1 0 18952 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_184
timestamp 1608254825
transform 1 0 18032 0 1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_409
timestamp 1608254825
transform 1 0 17940 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1530_
timestamp 1608254825
transform 1 0 19412 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1511_
timestamp 1608254825
transform 1 0 18584 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_219
timestamp 1608254825
transform 1 0 21252 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_41_211
timestamp 1608254825
transform 1 0 20516 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1527_
timestamp 1608254825
transform 1 0 20148 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1526_
timestamp 1608254825
transform 1 0 21988 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1498_
timestamp 1608254825
transform 1 0 20884 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_249
timestamp 1608254825
transform 1 0 24012 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_243
timestamp 1608254825
transform 1 0 23460 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_239
timestamp 1608254825
transform 1 0 23092 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_231
timestamp 1608254825
transform 1 0 22356 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_410
timestamp 1608254825
transform 1 0 23552 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1535_
timestamp 1608254825
transform 1 0 22724 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1496_
timestamp 1608254825
transform 1 0 23644 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_273
timestamp 1608254825
transform 1 0 26220 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_253
timestamp 1608254825
transform 1 0 24380 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2664_
timestamp 1608254825
transform 1 0 24472 0 1 24480
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_41_281
timestamp 1608254825
transform 1 0 26956 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _2161_
timestamp 1608254825
transform 1 0 26588 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_4  _1465_
timestamp 1608254825
transform 1 0 27324 0 1 24480
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_41_311
timestamp 1608254825
transform 1 0 29716 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_306
timestamp 1608254825
transform 1 0 29256 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_298
timestamp 1608254825
transform 1 0 28520 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_addressalyzerBlock.SPI_CLK
timestamp 1608254825
transform 1 0 28888 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_411
timestamp 1608254825
transform 1 0 29164 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_4  _2368_
timestamp 1608254825
transform 1 0 30084 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1626_
timestamp 1608254825
transform 1 0 29440 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_41_327
timestamp 1608254825
transform 1 0 31188 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__nor3_4  _1667_
timestamp 1608254825
transform 1 0 31924 0 1 24480
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_41_362
timestamp 1608254825
transform 1 0 34408 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_356
timestamp 1608254825
transform 1 0 33856 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_41_348
timestamp 1608254825
transform 1 0 33120 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _2096_
timestamp 1608254825
transform 1 0 34040 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_388
timestamp 1608254825
transform 1 0 36800 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_380
timestamp 1608254825
transform 1 0 36064 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_376
timestamp 1608254825
transform 1 0 35696 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_412
timestamp 1608254825
transform 1 0 34776 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _2088_
timestamp 1608254825
transform 1 0 36156 0 1 24480
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_4  _1240_
timestamp 1608254825
transform 1 0 34868 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_41_411
timestamp 1608254825
transform 1 0 38916 0 1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  _2499_
timestamp 1608254825
transform 1 0 37168 0 1 24480
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_41_417
timestamp 1608254825
transform 1 0 39468 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1608254825
transform -1 0 39836 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_42_22
timestamp 1608254825
transform 1 0 3128 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1608254825
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _2524_
timestamp 1608254825
transform 1 0 1380 0 -1 25568
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_42_44
timestamp 1608254825
transform 1 0 5152 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_30
timestamp 1608254825
transform 1 0 3864 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_413
timestamp 1608254825
transform 1 0 3956 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_4  _2060_
timestamp 1608254825
transform 1 0 4048 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_58
timestamp 1608254825
transform 1 0 6440 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_52
timestamp 1608254825
transform 1 0 5888 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  _2677_
timestamp 1608254825
transform 1 0 6532 0 -1 25568
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  _2050_
timestamp 1608254825
transform 1 0 5520 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_88
timestamp 1608254825
transform 1 0 9200 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_78
timestamp 1608254825
transform 1 0 8280 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _1401_
timestamp 1608254825
transform 1 0 8832 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_110
timestamp 1608254825
transform 1 0 11224 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_106
timestamp 1608254825
transform 1 0 10856 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_414
timestamp 1608254825
transform 1 0 9568 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_4  _1409_
timestamp 1608254825
transform 1 0 9660 0 -1 25568
box -38 -48 1234 592
use sky130_fd_sc_hd__and4_4  _1382_
timestamp 1608254825
transform 1 0 11316 0 -1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_42_128
timestamp 1608254825
transform 1 0 12880 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_120
timestamp 1608254825
transform 1 0 12144 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__nand3_4  _1391_
timestamp 1608254825
transform 1 0 12972 0 -1 25568
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_2  FILLER_42_154
timestamp 1608254825
transform 1 0 15272 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_151
timestamp 1608254825
transform 1 0 14996 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_42_143
timestamp 1608254825
transform 1 0 14260 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_415
timestamp 1608254825
transform 1 0 15180 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _2113_
timestamp 1608254825
transform 1 0 15456 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_172
timestamp 1608254825
transform 1 0 16928 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_168
timestamp 1608254825
transform 1 0 16560 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_160
timestamp 1608254825
transform 1 0 15824 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_4  _2193_
timestamp 1608254825
transform 1 0 17020 0 -1 25568
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  _1589_
timestamp 1608254825
transform 1 0 16192 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_195
timestamp 1608254825
transform 1 0 19044 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_189
timestamp 1608254825
transform 1 0 18492 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_4  _1499_
timestamp 1608254825
transform 1 0 19136 0 -1 25568
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_42_210
timestamp 1608254825
transform 1 0 20424 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_416
timestamp 1608254825
transform 1 0 20792 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__nand3_4  _1595_
timestamp 1608254825
transform 1 0 20884 0 -1 25568
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_42_247
timestamp 1608254825
transform 1 0 23828 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_237
timestamp 1608254825
transform 1 0 22908 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_229
timestamp 1608254825
transform 1 0 22172 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__or3_4  _1602_
timestamp 1608254825
transform 1 0 23000 0 -1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1510_
timestamp 1608254825
transform 1 0 24196 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_271
timestamp 1608254825
transform 1 0 26036 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_254
timestamp 1608254825
transform 1 0 24472 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_4  _1505_
timestamp 1608254825
transform 1 0 24840 0 -1 25568
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_42_296
timestamp 1608254825
transform 1 0 28336 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_276
timestamp 1608254825
transform 1 0 26496 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_417
timestamp 1608254825
transform 1 0 26404 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2667_
timestamp 1608254825
transform 1 0 26588 0 -1 25568
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_42_312
timestamp 1608254825
transform 1 0 29808 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_4  _2212_
timestamp 1608254825
transform 1 0 30176 0 -1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_4  _1459_
timestamp 1608254825
transform 1 0 28704 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_332
timestamp 1608254825
transform 1 0 31648 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_325
timestamp 1608254825
transform 1 0 31004 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_418
timestamp 1608254825
transform 1 0 32016 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_4  _1669_
timestamp 1608254825
transform 1 0 32108 0 -1 25568
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _1632_
timestamp 1608254825
transform 1 0 31372 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_350
timestamp 1608254825
transform 1 0 33304 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_4  _1670_
timestamp 1608254825
transform 1 0 33672 0 -1 25568
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_42_385
timestamp 1608254825
transform 1 0 36524 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_371
timestamp 1608254825
transform 1 0 35236 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_367
timestamp 1608254825
transform 1 0 34868 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_4  _1245_
timestamp 1608254825
transform 1 0 35328 0 -1 25568
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_3  FILLER_42_398
timestamp 1608254825
transform 1 0 37720 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_393
timestamp 1608254825
transform 1 0 37260 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_419
timestamp 1608254825
transform 1 0 37628 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_4  _2394_
timestamp 1608254825
transform 1 0 37996 0 -1 25568
box -38 -48 1234 592
use sky130_fd_sc_hd__buf_2  _1202_
timestamp 1608254825
transform 1 0 36892 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_414
timestamp 1608254825
transform 1 0 39192 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1608254825
transform -1 0 39836 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_17
timestamp 1608254825
transform 1 0 2668 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_3
timestamp 1608254825
transform 1 0 1380 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1608254825
transform 1 0 1104 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__a41oi_4  _2059_
timestamp 1608254825
transform 1 0 3036 0 1 25568
box -38 -48 2062 592
use sky130_fd_sc_hd__nor3_4  _2058_
timestamp 1608254825
transform 1 0 1472 0 1 25568
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_43_43
timestamp 1608254825
transform 1 0 5060 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_62
timestamp 1608254825
transform 1 0 6808 0 1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_60
timestamp 1608254825
transform 1 0 6624 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_56
timestamp 1608254825
transform 1 0 6256 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_420
timestamp 1608254825
transform 1 0 6716 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__and4_4  _2057_
timestamp 1608254825
transform 1 0 5428 0 1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_4  _1406_
timestamp 1608254825
transform 1 0 7360 0 1 25568
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_43_81
timestamp 1608254825
transform 1 0 8556 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_4  _1410_
timestamp 1608254825
transform 1 0 8924 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_97
timestamp 1608254825
transform 1 0 10028 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__a41o_4  _1397_
timestamp 1608254825
transform 1 0 10396 0 1 25568
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_43_123
timestamp 1608254825
transform 1 0 12420 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_118
timestamp 1608254825
transform 1 0 11960 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_421
timestamp 1608254825
transform 1 0 12328 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_4  _1390_
timestamp 1608254825
transform 1 0 12788 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_153
timestamp 1608254825
transform 1 0 15180 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_43_147
timestamp 1608254825
transform 1 0 14628 0 1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_139
timestamp 1608254825
transform 1 0 13892 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_4  _2265_
timestamp 1608254825
transform 1 0 15272 0 1 25568
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  _1383_
timestamp 1608254825
transform 1 0 14260 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_182
timestamp 1608254825
transform 1 0 17848 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_178
timestamp 1608254825
transform 1 0 17480 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_170
timestamp 1608254825
transform 1 0 16744 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1592_
timestamp 1608254825
transform 1 0 17112 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_195
timestamp 1608254825
transform 1 0 19044 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_191
timestamp 1608254825
transform 1 0 18676 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_422
timestamp 1608254825
transform 1 0 17940 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_4  _2211_
timestamp 1608254825
transform 1 0 19136 0 1 25568
box -38 -48 1234 592
use sky130_fd_sc_hd__or2_4  _2167_
timestamp 1608254825
transform 1 0 18032 0 1 25568
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_43_223
timestamp 1608254825
transform 1 0 21620 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_43_217
timestamp 1608254825
transform 1 0 21068 0 1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_209
timestamp 1608254825
transform 1 0 20332 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_4  _1596_
timestamp 1608254825
transform 1 0 21712 0 1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _1500_
timestamp 1608254825
transform 1 0 20700 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_240
timestamp 1608254825
transform 1 0 23184 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_233
timestamp 1608254825
transform 1 0 22540 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_423
timestamp 1608254825
transform 1 0 23552 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _1600_
timestamp 1608254825
transform 1 0 23644 0 1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1590_
timestamp 1608254825
transform 1 0 22908 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_271
timestamp 1608254825
transform 1 0 26036 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_258
timestamp 1608254825
transform 1 0 24840 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_254
timestamp 1608254825
transform 1 0 24472 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_4  _1501_
timestamp 1608254825
transform 1 0 24932 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_287
timestamp 1608254825
transform 1 0 27508 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_4  _1540_
timestamp 1608254825
transform 1 0 27876 0 1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_4  _1504_
timestamp 1608254825
transform 1 0 26404 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_306
timestamp 1608254825
transform 1 0 29256 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_304
timestamp 1608254825
transform 1 0 29072 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_300
timestamp 1608254825
transform 1 0 28704 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_424
timestamp 1608254825
transform 1 0 29164 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_4  _2213_
timestamp 1608254825
transform 1 0 29624 0 1 25568
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_43_331
timestamp 1608254825
transform 1 0 31556 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_327
timestamp 1608254825
transform 1 0 31188 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_323
timestamp 1608254825
transform 1 0 30820 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2656_
timestamp 1608254825
transform 1 0 31924 0 1 25568
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_2  _1671_
timestamp 1608254825
transform 1 0 31280 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_362
timestamp 1608254825
transform 1 0 34408 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_354
timestamp 1608254825
transform 1 0 33672 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1212_
timestamp 1608254825
transform 1 0 34040 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_43_367
timestamp 1608254825
transform 1 0 34868 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_425
timestamp 1608254825
transform 1 0 34776 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2701_
timestamp 1608254825
transform 1 0 35144 0 1 25568
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_43_389
timestamp 1608254825
transform 1 0 36892 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2510_
timestamp 1608254825
transform 1 0 37260 0 1 25568
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_43_412
timestamp 1608254825
transform 1 0 39008 0 1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1608254825
transform -1 0 39836 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_44_9
timestamp 1608254825
transform 1 0 1932 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_44_3
timestamp 1608254825
transform 1 0 1380 0 -1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1608254825
transform 1 0 1104 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__a41o_4  _2051_
timestamp 1608254825
transform 1 0 2024 0 -1 26656
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_44_27
timestamp 1608254825
transform 1 0 3588 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_426
timestamp 1608254825
transform 1 0 3956 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2523_
timestamp 1608254825
transform 1 0 4048 0 -1 26656
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_44_59
timestamp 1608254825
transform 1 0 6532 0 -1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_44_51
timestamp 1608254825
transform 1 0 5796 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _2022_
timestamp 1608254825
transform 1 0 6164 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__nand4_4  _1402_
timestamp 1608254825
transform 1 0 7084 0 -1 26656
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_2  FILLER_44_90
timestamp 1608254825
transform 1 0 9384 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_44_82
timestamp 1608254825
transform 1 0 8648 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_44_112
timestamp 1608254825
transform 1 0 11408 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_427
timestamp 1608254825
transform 1 0 9568 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2676_
timestamp 1608254825
transform 1 0 9660 0 -1 26656
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_44_133
timestamp 1608254825
transform 1 0 13340 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__nand4_4  _1259_
timestamp 1608254825
transform 1 0 11776 0 -1 26656
box -38 -48 1602 592
use sky130_fd_sc_hd__nand2_4  _1257_
timestamp 1608254825
transform 1 0 13708 0 -1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_44_146
timestamp 1608254825
transform 1 0 14536 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_m1_clk_local
timestamp 1608254825
transform 1 0 14904 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_428
timestamp 1608254825
transform 1 0 15180 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__nor3_4  _1594_
timestamp 1608254825
transform 1 0 15272 0 -1 26656
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_1  FILLER_44_175
timestamp 1608254825
transform 1 0 17204 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_167
timestamp 1608254825
transform 1 0 16468 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_4  _2242_
timestamp 1608254825
transform 1 0 17296 0 -1 26656
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_44_205
timestamp 1608254825
transform 1 0 19964 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_44_192
timestamp 1608254825
transform 1 0 18768 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_4  _1591_
timestamp 1608254825
transform 1 0 19136 0 -1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_44_226
timestamp 1608254825
transform 1 0 21896 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_219
timestamp 1608254825
transform 1 0 21252 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_213
timestamp 1608254825
transform 1 0 20700 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_429
timestamp 1608254825
transform 1 0 20792 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1539_
timestamp 1608254825
transform 1 0 21620 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1514_
timestamp 1608254825
transform 1 0 20884 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_250
timestamp 1608254825
transform 1 0 24104 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_243
timestamp 1608254825
transform 1 0 23460 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1601_
timestamp 1608254825
transform 1 0 23828 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_4  _1599_
timestamp 1608254825
transform 1 0 22264 0 -1 26656
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_44_271
timestamp 1608254825
transform 1 0 26036 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__nand4_4  _1542_
timestamp 1608254825
transform 1 0 24472 0 -1 26656
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_44_280
timestamp 1608254825
transform 1 0 26864 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_430
timestamp 1608254825
transform 1 0 26404 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2668_
timestamp 1608254825
transform 1 0 27232 0 -1 26656
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  _1437_
timestamp 1608254825
transform 1 0 26496 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_309
timestamp 1608254825
transform 1 0 29532 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_44_303
timestamp 1608254825
transform 1 0 28980 0 -1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_4  _2282_
timestamp 1608254825
transform 1 0 29624 0 -1 26656
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_2  FILLER_44_337
timestamp 1608254825
transform 1 0 32108 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_332
timestamp 1608254825
transform 1 0 31648 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_44_323
timestamp 1608254825
transform 1 0 30820 0 -1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_431
timestamp 1608254825
transform 1 0 32016 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _2392_
timestamp 1608254825
transform 1 0 31372 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_4  _2285_
timestamp 1608254825
transform 1 0 32292 0 -1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_44_348
timestamp 1608254825
transform 1 0 33120 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2479_
timestamp 1608254825
transform 1 0 33488 0 -1 26656
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_44_371
timestamp 1608254825
transform 1 0 35236 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__nand3_4  _1238_
timestamp 1608254825
transform 1 0 35972 0 -1 26656
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_44_401
timestamp 1608254825
transform 1 0 37996 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_393
timestamp 1608254825
transform 1 0 37260 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_432
timestamp 1608254825
transform 1 0 37628 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _2393_
timestamp 1608254825
transform 1 0 38364 0 -1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1200_
timestamp 1608254825
transform 1 0 37720 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_44_414
timestamp 1608254825
transform 1 0 39192 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1608254825
transform -1 0 39836 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_45_3
timestamp 1608254825
transform 1 0 1380 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1608254825
transform 1 0 1104 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _2525_
timestamp 1608254825
transform 1 0 1564 0 1 26656
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_45_45
timestamp 1608254825
transform 1 0 5244 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_45_24
timestamp 1608254825
transform 1 0 3312 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__nand4_4  _1988_
timestamp 1608254825
transform 1 0 3680 0 1 26656
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_45_57
timestamp 1608254825
transform 1 0 6348 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_433
timestamp 1608254825
transform 1 0 6716 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2678_
timestamp 1608254825
transform 1 0 6808 0 1 26656
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  _1362_
timestamp 1608254825
transform 1 0 5980 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_89
timestamp 1608254825
transform 1 0 9292 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_81
timestamp 1608254825
transform 1 0 8556 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1275_
timestamp 1608254825
transform 1 0 9384 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_105
timestamp 1608254825
transform 1 0 10764 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_94
timestamp 1608254825
transform 1 0 9752 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_10_0_m1_clk_local
timestamp 1608254825
transform 1 0 10120 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1396_
timestamp 1608254825
transform 1 0 10396 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_4  _1255_
timestamp 1608254825
transform 1 0 11132 0 1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_45_134
timestamp 1608254825
transform 1 0 13432 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_126
timestamp 1608254825
transform 1 0 12696 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_45_118
timestamp 1608254825
transform 1 0 11960 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_434
timestamp 1608254825
transform 1 0 12328 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2679_
timestamp 1608254825
transform 1 0 13524 0 1 26656
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_2  _1256_
timestamp 1608254825
transform 1 0 12420 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_45_154
timestamp 1608254825
transform 1 0 15272 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _2154_
timestamp 1608254825
transform 1 0 15640 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_179
timestamp 1608254825
transform 1 0 17572 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_162
timestamp 1608254825
transform 1 0 16008 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_4  _2281_
timestamp 1608254825
transform 1 0 16376 0 1 26656
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_45_202
timestamp 1608254825
transform 1 0 19688 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_435
timestamp 1608254825
transform 1 0 17940 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__o32a_4  _2155_
timestamp 1608254825
transform 1 0 18032 0 1 26656
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_8  FILLER_45_215
timestamp 1608254825
transform 1 0 20884 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_4  _2156_
timestamp 1608254825
transform 1 0 20056 0 1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_4  _1543_
timestamp 1608254825
transform 1 0 21620 0 1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_45_245
timestamp 1608254825
transform 1 0 23644 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_240
timestamp 1608254825
transform 1 0 23184 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_232
timestamp 1608254825
transform 1 0 22448 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_436
timestamp 1608254825
transform 1 0 23552 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2657_
timestamp 1608254825
transform 1 0 23736 0 1 26656
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  _1531_
timestamp 1608254825
transform 1 0 22816 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_265
timestamp 1608254825
transform 1 0 25484 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_4  _1586_
timestamp 1608254825
transform 1 0 25852 0 1 26656
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_6  FILLER_45_283
timestamp 1608254825
transform 1 0 27140 0 1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_4  _2284_
timestamp 1608254825
transform 1 0 27692 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_317
timestamp 1608254825
transform 1 0 30268 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_306
timestamp 1608254825
transform 1 0 29256 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_301
timestamp 1608254825
transform 1 0 28796 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_437
timestamp 1608254825
transform 1 0 29164 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__or4_4  _2396_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 29440 0 1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_45_340
timestamp 1608254825
transform 1 0 32384 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _2512_
timestamp 1608254825
transform 1 0 30636 0 1 26656
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_45_365
timestamp 1608254825
transform 1 0 34684 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_361
timestamp 1608254825
transform 1 0 34316 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_4  _2286_
timestamp 1608254825
transform 1 0 33120 0 1 26656
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_6  FILLER_45_372
timestamp 1608254825
transform 1 0 35328 0 1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_367
timestamp 1608254825
transform 1 0 34868 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_438
timestamp 1608254825
transform 1 0 34776 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1872_
timestamp 1608254825
transform 1 0 34960 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_4  _1214_
timestamp 1608254825
transform 1 0 35880 0 1 26656
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_8  FILLER_45_408
timestamp 1608254825
transform 1 0 38640 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_399
timestamp 1608254825
transform 1 0 37812 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_45_391
timestamp 1608254825
transform 1 0 37076 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__or2_4  _1203_
timestamp 1608254825
transform 1 0 37996 0 1 26656
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_45_416
timestamp 1608254825
transform 1 0 39376 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1608254825
transform -1 0 39836 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_47_8
timestamp 1608254825
transform 1 0 1840 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_3
timestamp 1608254825
transform 1 0 1380 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_9
timestamp 1608254825
transform 1 0 1932 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_46_3
timestamp 1608254825
transform 1 0 1380 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1608254825
transform 1 0 1104 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1608254825
transform 1 0 1104 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2045_
timestamp 1608254825
transform 1 0 1656 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2036_
timestamp 1608254825
transform 1 0 1564 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_47_15
timestamp 1608254825
transform 1 0 2484 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_22
timestamp 1608254825
transform 1 0 3128 0 -1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__and3_4  _2052_
timestamp 1608254825
transform 1 0 2300 0 -1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1980_
timestamp 1608254825
transform 1 0 2208 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_4  _2046_
timestamp 1608254825
transform 1 0 2852 0 1 27744
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_47_32
timestamp 1608254825
transform 1 0 4048 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_45
timestamp 1608254825
transform 1 0 5244 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_8_0_m1_clk_local
timestamp 1608254825
transform 1 0 3680 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_439
timestamp 1608254825
transform 1 0 3956 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_4  _2047_
timestamp 1608254825
transform 1 0 4048 0 -1 27744
box -38 -48 1234 592
use sky130_fd_sc_hd__o21ai_4  _2043_
timestamp 1608254825
transform 1 0 4416 0 1 27744
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_47_57
timestamp 1608254825
transform 1 0 6348 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_49
timestamp 1608254825
transform 1 0 5612 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_52
timestamp 1608254825
transform 1 0 5888 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _2035_
timestamp 1608254825
transform 1 0 5980 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1404_
timestamp 1608254825
transform 1 0 5612 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1287_
timestamp 1608254825
transform 1 0 6256 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_64
timestamp 1608254825
transform 1 0 6992 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_60
timestamp 1608254825
transform 1 0 6624 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_446
timestamp 1608254825
transform 1 0 6716 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_4  _1403_
timestamp 1608254825
transform 1 0 6808 0 1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_4  _1400_
timestamp 1608254825
transform 1 0 7084 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_71
timestamp 1608254825
transform 1 0 7636 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_m1_clk_local
timestamp 1608254825
transform 1 0 8004 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_47_82
timestamp 1608254825
transform 1 0 8648 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_77
timestamp 1608254825
transform 1 0 8188 0 -1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _1328_
timestamp 1608254825
transform 1 0 8280 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_88
timestamp 1608254825
transform 1 0 9200 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 1608254825
transform 1 0 8740 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1311_
timestamp 1608254825
transform 1 0 9016 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1274_
timestamp 1608254825
transform 1 0 8832 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_90
timestamp 1608254825
transform 1 0 9384 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_114
timestamp 1608254825
transform 1 0 11592 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_107
timestamp 1608254825
transform 1 0 10948 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_107
timestamp 1608254825
transform 1 0 10948 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_93
timestamp 1608254825
transform 1 0 9660 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_m1_clk_local
timestamp 1608254825
transform 1 0 11316 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_440
timestamp 1608254825
transform 1 0 9568 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_4  _1387_
timestamp 1608254825
transform 1 0 9752 0 -1 27744
box -38 -48 1234 592
use sky130_fd_sc_hd__buf_2  _1381_
timestamp 1608254825
transform 1 0 11316 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_4  _1373_
timestamp 1608254825
transform 1 0 9752 0 1 27744
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_8  FILLER_47_127
timestamp 1608254825
transform 1 0 12788 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_47_118
timestamp 1608254825
transform 1 0 11960 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_136
timestamp 1608254825
transform 1 0 13616 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_115
timestamp 1608254825
transform 1 0 11684 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_447
timestamp 1608254825
transform 1 0 12328 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_4  _1398_
timestamp 1608254825
transform 1 0 13524 0 1 27744
box -38 -48 1234 592
use sky130_fd_sc_hd__nand4_4  _1384_
timestamp 1608254825
transform 1 0 12052 0 -1 27744
box -38 -48 1602 592
use sky130_fd_sc_hd__buf_2  _1366_
timestamp 1608254825
transform 1 0 12420 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1258_
timestamp 1608254825
transform 1 0 11684 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_47_159
timestamp 1608254825
transform 1 0 15732 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_155
timestamp 1608254825
transform 1 0 15364 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_148
timestamp 1608254825
transform 1 0 14720 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_157
timestamp 1608254825
transform 1 0 15548 0 -1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_46_149
timestamp 1608254825
transform 1 0 14812 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_441
timestamp 1608254825
transform 1 0 15180 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1394_
timestamp 1608254825
transform 1 0 15272 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1386_
timestamp 1608254825
transform 1 0 15088 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_4  _1385_
timestamp 1608254825
transform 1 0 13984 0 -1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_47_181
timestamp 1608254825
transform 1 0 17756 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_47_173
timestamp 1608254825
transform 1 0 17020 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_46_177
timestamp 1608254825
transform 1 0 17388 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_4  _1661_
timestamp 1608254825
transform 1 0 15824 0 1 27744
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_4  _1658_
timestamp 1608254825
transform 1 0 17756 0 -1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_4  _1657_
timestamp 1608254825
transform 1 0 16100 0 -1 27744
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_1  FILLER_46_196
timestamp 1608254825
transform 1 0 19136 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_46_190
timestamp 1608254825
transform 1 0 18584 0 -1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_448
timestamp 1608254825
transform 1 0 17940 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__o41ai_4  _2218_
timestamp 1608254825
transform 1 0 18032 0 1 27744
box -38 -48 2062 592
use sky130_fd_sc_hd__o21ai_4  _2153_
timestamp 1608254825
transform 1 0 19228 0 -1 27744
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_1  FILLER_47_210
timestamp 1608254825
transform 1 0 20424 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_206
timestamp 1608254825
transform 1 0 20056 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_228
timestamp 1608254825
transform 1 0 22080 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_210
timestamp 1608254825
transform 1 0 20424 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_442
timestamp 1608254825
transform 1 0 20792 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__o32ai_4  _1655_
timestamp 1608254825
transform 1 0 20516 0 1 27744
box -38 -48 2062 592
use sky130_fd_sc_hd__a21oi_4  _1654_
timestamp 1608254825
transform 1 0 20884 0 -1 27744
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_47_233
timestamp 1608254825
transform 1 0 22540 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_236
timestamp 1608254825
transform 1 0 22816 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1583_
timestamp 1608254825
transform 1 0 22448 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1494_
timestamp 1608254825
transform 1 0 22908 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_47_245
timestamp 1608254825
transform 1 0 23644 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_47_240
timestamp 1608254825
transform 1 0 23184 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_240
timestamp 1608254825
transform 1 0 23184 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_449
timestamp 1608254825
transform 1 0 23552 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _2139_
timestamp 1608254825
transform 1 0 23920 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_4  _1663_
timestamp 1608254825
transform 1 0 23276 0 -1 27744
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_47_260
timestamp 1608254825
transform 1 0 25024 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_252
timestamp 1608254825
transform 1 0 24288 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_267
timestamp 1608254825
transform 1 0 25668 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_46_254
timestamp 1608254825
transform 1 0 24472 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_4  _1662_
timestamp 1608254825
transform 1 0 24840 0 -1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _1636_
timestamp 1608254825
transform 1 0 24656 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_4  _1570_
timestamp 1608254825
transform 1 0 25392 0 1 27744
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_6  FILLER_47_291
timestamp 1608254825
transform 1 0 27876 0 1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_47_278
timestamp 1608254825
transform 1 0 26680 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_295
timestamp 1608254825
transform 1 0 28244 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_282
timestamp 1608254825
transform 1 0 27048 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_276
timestamp 1608254825
transform 1 0 26496 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_443
timestamp 1608254825
transform 1 0 26404 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__and4_4  _2163_
timestamp 1608254825
transform 1 0 27416 0 -1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__and4_4  _1637_
timestamp 1608254825
transform 1 0 27048 0 1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _1495_
timestamp 1608254825
transform 1 0 26680 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_313
timestamp 1608254825
transform 1 0 29900 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_301
timestamp 1608254825
transform 1 0 28796 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_312
timestamp 1608254825
transform 1 0 29808 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_450
timestamp 1608254825
transform 1 0 29164 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2597_
timestamp 1608254825
transform 1 0 30268 0 1 27744
box -38 -48 1786 592
use sky130_fd_sc_hd__nor3_4  _2283_
timestamp 1608254825
transform 1 0 28612 0 -1 27744
box -38 -48 1234 592
use sky130_fd_sc_hd__and2_4  _1868_
timestamp 1608254825
transform 1 0 29256 0 1 27744
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _1866_
timestamp 1608254825
transform 1 0 28428 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_336
timestamp 1608254825
transform 1 0 32016 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_46_337
timestamp 1608254825
transform 1 0 32108 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_46_330
timestamp 1608254825
transform 1 0 31464 0 -1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_320
timestamp 1608254825
transform 1 0 30544 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_444
timestamp 1608254825
transform 1 0 32016 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__or4_4  _2395_
timestamp 1608254825
transform 1 0 30636 0 -1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_4  _2166_
timestamp 1608254825
transform 1 0 32384 0 1 27744
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _1597_
timestamp 1608254825
transform 1 0 32384 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_47_365
timestamp 1608254825
transform 1 0 34684 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_361
timestamp 1608254825
transform 1 0 34316 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_353
timestamp 1608254825
transform 1 0 33580 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_364
timestamp 1608254825
transform 1 0 34592 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_356
timestamp 1608254825
transform 1 0 33856 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_343
timestamp 1608254825
transform 1 0 32660 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _2189_
timestamp 1608254825
transform 1 0 34224 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_4  _2165_
timestamp 1608254825
transform 1 0 33028 0 -1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _1604_
timestamp 1608254825
transform 1 0 33948 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_47_367
timestamp 1608254825
transform 1 0 34868 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_46_385
timestamp 1608254825
transform 1 0 36524 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_381
timestamp 1608254825
transform 1 0 36156 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_451
timestamp 1608254825
transform 1 0 34776 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2707_
timestamp 1608254825
transform 1 0 35144 0 1 27744
box -38 -48 1786 592
use sky130_fd_sc_hd__or2_4  _1215_
timestamp 1608254825
transform 1 0 36616 0 -1 27744
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_4  _1213_
timestamp 1608254825
transform 1 0 34960 0 -1 27744
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_47_389
timestamp 1608254825
transform 1 0 36892 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_398
timestamp 1608254825
transform 1 0 37720 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_393
timestamp 1608254825
transform 1 0 37260 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_445
timestamp 1608254825
transform 1 0 37628 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2706_
timestamp 1608254825
transform 1 0 37260 0 1 27744
box -38 -48 1786 592
use sky130_fd_sc_hd__o21ai_4  _1204_
timestamp 1608254825
transform 1 0 37812 0 -1 27744
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_6  FILLER_47_412
timestamp 1608254825
transform 1 0 39008 0 1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_46_412
timestamp 1608254825
transform 1 0 39008 0 -1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1608254825
transform -1 0 39836 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1608254825
transform -1 0 39836 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_48_3
timestamp 1608254825
transform 1 0 1380 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1608254825
transform 1 0 1104 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _2526_
timestamp 1608254825
transform 1 0 1656 0 -1 28832
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_48_36
timestamp 1608254825
transform 1 0 4416 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_32
timestamp 1608254825
transform 1 0 4048 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_25
timestamp 1608254825
transform 1 0 3404 0 -1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_452
timestamp 1608254825
transform 1 0 3956 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__nor3_4  _2010_
timestamp 1608254825
transform 1 0 4508 0 -1 28832
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_48_50
timestamp 1608254825
transform 1 0 5704 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2527_
timestamp 1608254825
transform 1 0 6072 0 -1 28832
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_48_88
timestamp 1608254825
transform 1 0 9200 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_84
timestamp 1608254825
transform 1 0 8832 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_80
timestamp 1608254825
transform 1 0 8464 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_73
timestamp 1608254825
transform 1 0 7820 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1375_
timestamp 1608254825
transform 1 0 8188 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1372_
timestamp 1608254825
transform 1 0 8924 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_48_97
timestamp 1608254825
transform 1 0 10028 0 -1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_453
timestamp 1608254825
transform 1 0 9568 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2681_
timestamp 1608254825
transform 1 0 10580 0 -1 28832
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  _1378_
timestamp 1608254825
transform 1 0 9660 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_122
timestamp 1608254825
transform 1 0 12328 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _2682_
timestamp 1608254825
transform 1 0 13064 0 -1 28832
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_48_149
timestamp 1608254825
transform 1 0 14812 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_454
timestamp 1608254825
transform 1 0 15180 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2oi_4  _1659_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608254825
transform 1 0 15272 0 -1 28832
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_4  FILLER_48_175
timestamp 1608254825
transform 1 0 17204 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__o41ai_4  _2168_
timestamp 1608254825
transform 1 0 17572 0 -1 28832
box -38 -48 2062 592
use sky130_fd_sc_hd__decap_4  FILLER_48_201
timestamp 1608254825
transform 1 0 19596 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _2111_
timestamp 1608254825
transform 1 0 19964 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_219
timestamp 1608254825
transform 1 0 21252 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_213
timestamp 1608254825
transform 1 0 20700 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_209
timestamp 1608254825
transform 1 0 20332 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_455
timestamp 1608254825
transform 1 0 20792 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__o32ai_4  _2140_
timestamp 1608254825
transform 1 0 21620 0 -1 28832
box -38 -48 2062 592
use sky130_fd_sc_hd__buf_2  _1587_
timestamp 1608254825
transform 1 0 20884 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_245
timestamp 1608254825
transform 1 0 23644 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_4  _1603_
timestamp 1608254825
transform 1 0 24012 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_271
timestamp 1608254825
transform 1 0 26036 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_261
timestamp 1608254825
transform 1 0 25116 0 -1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _1464_
timestamp 1608254825
transform 1 0 25668 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_289
timestamp 1608254825
transform 1 0 27692 0 -1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_456
timestamp 1608254825
transform 1 0 26404 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_4  _2164_
timestamp 1608254825
transform 1 0 28244 0 -1 28832
box -38 -48 1234 592
use sky130_fd_sc_hd__o21ai_4  _1569_
timestamp 1608254825
transform 1 0 26496 0 -1 28832
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_48_308
timestamp 1608254825
transform 1 0 29440 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_4  _2187_
timestamp 1608254825
transform 1 0 29808 0 -1 28832
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_48_332
timestamp 1608254825
transform 1 0 31648 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_325
timestamp 1608254825
transform 1 0 31004 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_457
timestamp 1608254825
transform 1 0 32016 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _2162_
timestamp 1608254825
transform 1 0 31372 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__and2_4  _1873_
timestamp 1608254825
transform 1 0 32108 0 -1 28832
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_48_344
timestamp 1608254825
transform 1 0 32752 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2484_
timestamp 1608254825
transform 1 0 33120 0 -1 28832
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_48_384
timestamp 1608254825
transform 1 0 36432 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_367
timestamp 1608254825
transform 1 0 34868 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_4  _1217_
timestamp 1608254825
transform 1 0 35236 0 -1 28832
box -38 -48 1234 592
use sky130_fd_sc_hd__buf_2  _1209_
timestamp 1608254825
transform 1 0 36800 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_398
timestamp 1608254825
transform 1 0 37720 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_48_396
timestamp 1608254825
transform 1 0 37536 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_392
timestamp 1608254825
transform 1 0 37168 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_458
timestamp 1608254825
transform 1 0 37628 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_4  _1216_
timestamp 1608254825
transform 1 0 37904 0 -1 28832
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_1  FILLER_48_417
timestamp 1608254825
transform 1 0 39468 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_413
timestamp 1608254825
transform 1 0 39100 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1608254825
transform -1 0 39836 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_49_13
timestamp 1608254825
transform 1 0 2300 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_3
timestamp 1608254825
transform 1 0 1380 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1608254825
transform 1 0 1104 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__and3_4  _2039_
timestamp 1608254825
transform 1 0 1472 0 1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__and4_4  _2030_
timestamp 1608254825
transform 1 0 2668 0 1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_49_39
timestamp 1608254825
transform 1 0 4692 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_26
timestamp 1608254825
transform 1 0 3496 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_4  _2044_
timestamp 1608254825
transform 1 0 5060 0 1 28832
box -38 -48 1326 592
use sky130_fd_sc_hd__nor2_4  _2024_
timestamp 1608254825
transform 1 0 3864 0 1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_49_66
timestamp 1608254825
transform 1 0 7176 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_57
timestamp 1608254825
transform 1 0 6348 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_459
timestamp 1608254825
transform 1 0 6716 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _2025_
timestamp 1608254825
transform 1 0 6808 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_89
timestamp 1608254825
transform 1 0 9292 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2683_
timestamp 1608254825
transform 1 0 7544 0 1 28832
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_49_114
timestamp 1608254825
transform 1 0 11592 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_49_107
timestamp 1608254825
transform 1 0 10948 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_4  _1374_
timestamp 1608254825
transform 1 0 9660 0 1 28832
box -38 -48 1326 592
use sky130_fd_sc_hd__inv_2  _1365_
timestamp 1608254825
transform 1 0 11316 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_49_123
timestamp 1608254825
transform 1 0 12420 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_460
timestamp 1608254825
transform 1 0 12328 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_4  _1379_
timestamp 1608254825
transform 1 0 12696 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_49_149
timestamp 1608254825
transform 1 0 14812 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_145
timestamp 1608254825
transform 1 0 14444 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_138
timestamp 1608254825
transform 1 0 13800 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2oi_4  _1593_
timestamp 1608254825
transform 1 0 14904 0 1 28832
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_2  _1376_
timestamp 1608254825
transform 1 0 14168 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_49_179
timestamp 1608254825
transform 1 0 17572 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_171
timestamp 1608254825
transform 1 0 16836 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1582_
timestamp 1608254825
transform 1 0 17204 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_197
timestamp 1608254825
transform 1 0 19228 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_461
timestamp 1608254825
transform 1 0 17940 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_4  _2186_
timestamp 1608254825
transform 1 0 18032 0 1 28832
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_4  _2160_
timestamp 1608254825
transform 1 0 19596 0 1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_49_216
timestamp 1608254825
transform 1 0 20976 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_49_210
timestamp 1608254825
transform 1 0 20424 0 1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_4  _1584_
timestamp 1608254825
transform 1 0 21068 0 1 28832
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_49_240
timestamp 1608254825
transform 1 0 23184 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_231
timestamp 1608254825
transform 1 0 22356 0 1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_462
timestamp 1608254825
transform 1 0 23552 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__nor3_4  _1579_
timestamp 1608254825
transform 1 0 23644 0 1 28832
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _1572_
timestamp 1608254825
transform 1 0 22908 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_49_267
timestamp 1608254825
transform 1 0 25668 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_262
timestamp 1608254825
transform 1 0 25208 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_258
timestamp 1608254825
transform 1 0 24840 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__and2_4  _1635_
timestamp 1608254825
transform 1 0 26036 0 1 28832
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _1578_
timestamp 1608254825
transform 1 0 25300 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_285
timestamp 1608254825
transform 1 0 27324 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_278
timestamp 1608254825
transform 1 0 26680 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_4  _2188_
timestamp 1608254825
transform 1 0 27692 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1438_
timestamp 1608254825
transform 1 0 27048 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_49_301
timestamp 1608254825
transform 1 0 28796 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_463
timestamp 1608254825
transform 1 0 29164 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2601_
timestamp 1608254825
transform 1 0 29256 0 1 28832
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_49_340
timestamp 1608254825
transform 1 0 32384 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_325
timestamp 1608254825
transform 1 0 31004 0 1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_4  _2190_
timestamp 1608254825
transform 1 0 31556 0 1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_49_365
timestamp 1608254825
transform 1 0 34684 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_357
timestamp 1608254825
transform 1 0 33948 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_4  _2191_
timestamp 1608254825
transform 1 0 32752 0 1 28832
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_49_386
timestamp 1608254825
transform 1 0 36616 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_367
timestamp 1608254825
transform 1 0 34868 0 1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_464
timestamp 1608254825
transform 1 0 34776 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_4  _2400_
timestamp 1608254825
transform 1 0 35420 0 1 28832
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_6  FILLER_49_411
timestamp 1608254825
transform 1 0 38916 0 1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_49_403
timestamp 1608254825
transform 1 0 38180 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1219_
timestamp 1608254825
transform 1 0 38548 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_4  _1218_
timestamp 1608254825
transform 1 0 36984 0 1 28832
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_1  FILLER_49_417
timestamp 1608254825
transform 1 0 39468 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1608254825
transform -1 0 39836 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_50_22
timestamp 1608254825
transform 1 0 3128 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1608254825
transform 1 0 1104 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _2529_
timestamp 1608254825
transform 1 0 1380 0 -1 29920
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_50_36
timestamp 1608254825
transform 1 0 4416 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_30
timestamp 1608254825
transform 1 0 3864 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_465
timestamp 1608254825
transform 1 0 3956 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _2009_
timestamp 1608254825
transform 1 0 4048 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__nor4_4  _1989_
timestamp 1608254825
transform 1 0 4784 0 -1 29920
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_50_64
timestamp 1608254825
transform 1 0 6992 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_57
timestamp 1608254825
transform 1 0 6348 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2042_
timestamp 1608254825
transform 1 0 7360 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1981_
timestamp 1608254825
transform 1 0 6716 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_50_88
timestamp 1608254825
transform 1 0 9200 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_75
timestamp 1608254825
transform 1 0 8004 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_71
timestamp 1608254825
transform 1 0 7636 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_4  _1368_
timestamp 1608254825
transform 1 0 8096 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_106
timestamp 1608254825
transform 1 0 10856 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_466
timestamp 1608254825
transform 1 0 9568 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_4  _1388_
timestamp 1608254825
transform 1 0 11224 0 -1 29920
box -38 -48 1234 592
use sky130_fd_sc_hd__nor3_4  _1367_
timestamp 1608254825
transform 1 0 9660 0 -1 29920
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_50_136
timestamp 1608254825
transform 1 0 13616 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_123
timestamp 1608254825
transform 1 0 12420 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_4  _1249_
timestamp 1608254825
transform 1 0 12788 0 -1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_50_149
timestamp 1608254825
transform 1 0 14812 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_467
timestamp 1608254825
transform 1 0 15180 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _1377_
timestamp 1608254825
transform 1 0 13984 0 -1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  _1353_
timestamp 1608254825
transform 1 0 15272 0 -1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_50_182
timestamp 1608254825
transform 1 0 17848 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_50_163
timestamp 1608254825
transform 1 0 16100 0 -1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_4  _2152_
timestamp 1608254825
transform 1 0 16652 0 -1 29920
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_50_199
timestamp 1608254825
transform 1 0 19412 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_4  _2184_
timestamp 1608254825
transform 1 0 18216 0 -1 29920
box -38 -48 1234 592
use sky130_fd_sc_hd__buf_2  _1515_
timestamp 1608254825
transform 1 0 19780 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_227
timestamp 1608254825
transform 1 0 21988 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_223
timestamp 1608254825
transform 1 0 21620 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_219
timestamp 1608254825
transform 1 0 21252 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_213
timestamp 1608254825
transform 1 0 20700 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_50_207
timestamp 1608254825
transform 1 0 20148 0 -1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_468
timestamp 1608254825
transform 1 0 20792 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1581_
timestamp 1608254825
transform 1 0 20884 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1575_
timestamp 1608254825
transform 1 0 21712 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_50_244
timestamp 1608254825
transform 1 0 23552 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_4  _1585_
timestamp 1608254825
transform 1 0 22356 0 -1 29920
box -38 -48 1234 592
use sky130_fd_sc_hd__a21oi_4  _1580_
timestamp 1608254825
transform 1 0 23920 0 -1 29920
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_6  FILLER_50_269
timestamp 1608254825
transform 1 0 25852 0 -1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_50_261
timestamp 1608254825
transform 1 0 25116 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1576_
timestamp 1608254825
transform 1 0 25484 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_284
timestamp 1608254825
transform 1 0 27232 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_280
timestamp 1608254825
transform 1 0 26864 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_469
timestamp 1608254825
transform 1 0 26404 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2607_
timestamp 1608254825
transform 1 0 27324 0 -1 29920
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  _1463_
timestamp 1608254825
transform 1 0 26496 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_315
timestamp 1608254825
transform 1 0 30084 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_304
timestamp 1608254825
transform 1 0 29072 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__and4_4  _2192_
timestamp 1608254825
transform 1 0 30452 0 -1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__and2_4  _1863_
timestamp 1608254825
transform 1 0 29440 0 -1 29920
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_50_342
timestamp 1608254825
transform 1 0 32568 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_337
timestamp 1608254825
transform 1 0 32108 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_328
timestamp 1608254825
transform 1 0 31280 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_470
timestamp 1608254825
transform 1 0 32016 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1235_
timestamp 1608254825
transform 1 0 32200 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_50_365
timestamp 1608254825
transform 1 0 34684 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _2483_
timestamp 1608254825
transform 1 0 32936 0 -1 29920
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_50_373
timestamp 1608254825
transform 1 0 35420 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2708_
timestamp 1608254825
transform 1 0 35512 0 -1 29920
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_50_411
timestamp 1608254825
transform 1 0 38916 0 -1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_50_393
timestamp 1608254825
transform 1 0 37260 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_471
timestamp 1608254825
transform 1 0 37628 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_4  _2398_
timestamp 1608254825
transform 1 0 37720 0 -1 29920
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_1  FILLER_50_417
timestamp 1608254825
transform 1 0 39468 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1608254825
transform -1 0 39836 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_51_11
timestamp 1608254825
transform 1 0 2116 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_51_3
timestamp 1608254825
transform 1 0 1380 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1608254825
transform 1 0 1104 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__a41o_4  _2037_
timestamp 1608254825
transform 1 0 2300 0 1 29920
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_51_30
timestamp 1608254825
transform 1 0 3864 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__nand4_4  _2038_
timestamp 1608254825
transform 1 0 4232 0 1 29920
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_51_67
timestamp 1608254825
transform 1 0 7268 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_51_62
timestamp 1608254825
transform 1 0 6808 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_51_58
timestamp 1608254825
transform 1 0 6440 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_51_51
timestamp 1608254825
transform 1 0 5796 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_m1_clk_local
timestamp 1608254825
transform 1 0 6164 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_472
timestamp 1608254825
transform 1 0 6716 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1371_
timestamp 1608254825
transform 1 0 6992 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_51_80
timestamp 1608254825
transform 1 0 8464 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_4  _1369_
timestamp 1608254825
transform 1 0 8832 0 1 29920
box -38 -48 1326 592
use sky130_fd_sc_hd__nand2_4  _1261_
timestamp 1608254825
transform 1 0 7636 0 1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_51_114
timestamp 1608254825
transform 1 0 11592 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_51_98
timestamp 1608254825
transform 1 0 10120 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_4  _1360_
timestamp 1608254825
transform 1 0 10488 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_473
timestamp 1608254825
transform 1 0 12328 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2686_
timestamp 1608254825
transform 1 0 12420 0 1 29920
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_51_156
timestamp 1608254825
transform 1 0 15456 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_146
timestamp 1608254825
transform 1 0 14536 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_142
timestamp 1608254825
transform 1 0 14168 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__and4_4  _1347_
timestamp 1608254825
transform 1 0 14628 0 1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_51_179
timestamp 1608254825
transform 1 0 17572 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_51_164
timestamp 1608254825
transform 1 0 16192 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__o21ai_4  _2259_
timestamp 1608254825
transform 1 0 16376 0 1 29920
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_2  FILLER_51_196
timestamp 1608254825
transform 1 0 19136 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_51_184
timestamp 1608254825
transform 1 0 18032 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_474
timestamp 1608254825
transform 1 0 17940 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__a2111oi_4  _2256_
timestamp 1608254825
transform 1 0 19320 0 1 29920
box -38 -48 2062 592
use sky130_fd_sc_hd__decap_4  FILLER_51_220
timestamp 1608254825
transform 1 0 21344 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_4  _2235_
timestamp 1608254825
transform 1 0 21712 0 1 29920
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_1  FILLER_51_243
timestamp 1608254825
transform 1 0 23460 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_51_237
timestamp 1608254825
transform 1 0 22908 0 1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_475
timestamp 1608254825
transform 1 0 23552 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_4  _2257_
timestamp 1608254825
transform 1 0 23644 0 1 29920
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_6  FILLER_51_258
timestamp 1608254825
transform 1 0 24840 0 1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_4  _2253_
timestamp 1608254825
transform 1 0 25392 0 1 29920
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_51_293
timestamp 1608254825
transform 1 0 28060 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_282
timestamp 1608254825
transform 1 0 27048 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_278
timestamp 1608254825
transform 1 0 26680 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_8_0_addressalyzerBlock.SPI_CLK
timestamp 1608254825
transform 1 0 27140 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__or2_4  _1568_
timestamp 1608254825
transform 1 0 27416 0 1 29920
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_51_306
timestamp 1608254825
transform 1 0 29256 0 1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_51_301
timestamp 1608254825
transform 1 0 28796 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_476
timestamp 1608254825
transform 1 0 29164 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__and4_4  _2217_
timestamp 1608254825
transform 1 0 29808 0 1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _1652_
timestamp 1608254825
transform 1 0 28428 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_338
timestamp 1608254825
transform 1 0 32200 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_321
timestamp 1608254825
transform 1 0 30636 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_9_0_addressalyzerBlock.SPI_CLK
timestamp 1608254825
transform 1 0 32568 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_4  _2214_
timestamp 1608254825
transform 1 0 31004 0 1 29920
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_51_362
timestamp 1608254825
transform 1 0 34408 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_354
timestamp 1608254825
transform 1 0 33672 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_4  _1605_
timestamp 1608254825
transform 1 0 32844 0 1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _1207_
timestamp 1608254825
transform 1 0 34040 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_380
timestamp 1608254825
transform 1 0 36064 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_477
timestamp 1608254825
transform 1 0 34776 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _2397_
timestamp 1608254825
transform 1 0 36432 0 1 29920
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_4  _1223_
timestamp 1608254825
transform 1 0 34868 0 1 29920
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_51_391
timestamp 1608254825
transform 1 0 37076 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2547_
timestamp 1608254825
transform 1 0 37444 0 1 29920
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_51_414
timestamp 1608254825
transform 1 0 39192 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1608254825
transform -1 0 39836 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_53_8
timestamp 1608254825
transform 1 0 1840 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_53_3
timestamp 1608254825
transform 1 0 1380 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_52_3
timestamp 1608254825
transform 1 0 1380 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1608254825
transform 1 0 1104 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1608254825
transform 1 0 1104 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2034_
timestamp 1608254825
transform 1 0 1564 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__nand4_4  _2032_
timestamp 1608254825
transform 1 0 2208 0 1 31008
box -38 -48 1602 592
use sky130_fd_sc_hd__o21a_4  _2031_
timestamp 1608254825
transform 1 0 2484 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_29
timestamp 1608254825
transform 1 0 3772 0 1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_52_45
timestamp 1608254825
transform 1 0 5244 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_27
timestamp 1608254825
transform 1 0 3588 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_478
timestamp 1608254825
transform 1 0 3956 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__nor3_4  _2041_
timestamp 1608254825
transform 1 0 4048 0 -1 31008
box -38 -48 1234 592
use sky130_fd_sc_hd__a21oi_4  _2040_
timestamp 1608254825
transform 1 0 4324 0 1 31008
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_53_65
timestamp 1608254825
transform 1 0 7084 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_57
timestamp 1608254825
transform 1 0 6348 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_52
timestamp 1608254825
transform 1 0 5888 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_48
timestamp 1608254825
transform 1 0 5520 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_52_68
timestamp 1608254825
transform 1 0 7360 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_485
timestamp 1608254825
transform 1 0 6716 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2528_
timestamp 1608254825
transform 1 0 5612 0 -1 31008
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  _2011_
timestamp 1608254825
transform 1 0 5980 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1982_
timestamp 1608254825
transform 1 0 6808 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_53_88
timestamp 1608254825
transform 1 0 9200 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_85
timestamp 1608254825
transform 1 0 8924 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_11_0_m1_clk_local
timestamp 1608254825
transform 1 0 9292 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _2684_
timestamp 1608254825
transform 1 0 7452 0 1 31008
box -38 -48 1786 592
use sky130_fd_sc_hd__nand2_4  _1370_
timestamp 1608254825
transform 1 0 8096 0 -1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_53_101
timestamp 1608254825
transform 1 0 10396 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_96
timestamp 1608254825
transform 1 0 9936 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_479
timestamp 1608254825
transform 1 0 9568 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__nor4_4  _1350_
timestamp 1608254825
transform 1 0 10304 0 -1 31008
box -38 -48 1602 592
use sky130_fd_sc_hd__inv_2  _1349_
timestamp 1608254825
transform 1 0 9660 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_4  _1277_
timestamp 1608254825
transform 1 0 10764 0 1 31008
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_4  _1260_
timestamp 1608254825
transform 1 0 9568 0 1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_53_135
timestamp 1608254825
transform 1 0 13524 0 1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_53_118
timestamp 1608254825
transform 1 0 11960 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_52_124
timestamp 1608254825
transform 1 0 12512 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_52_117
timestamp 1608254825
transform 1 0 11868 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_486
timestamp 1608254825
transform 1 0 12328 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_4  _1359_
timestamp 1608254825
transform 1 0 12420 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__nand4_4  _1352_
timestamp 1608254825
transform 1 0 13248 0 -1 31008
box -38 -48 1602 592
use sky130_fd_sc_hd__inv_2  _1262_
timestamp 1608254825
transform 1 0 12236 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_53_150
timestamp 1608254825
transform 1 0 14904 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_146
timestamp 1608254825
transform 1 0 14536 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_141
timestamp 1608254825
transform 1 0 14076 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_149
timestamp 1608254825
transform 1 0 14812 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_480
timestamp 1608254825
transform 1 0 15180 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2688_
timestamp 1608254825
transform 1 0 14996 0 1 31008
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  _1351_
timestamp 1608254825
transform 1 0 14168 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_4  _1348_
timestamp 1608254825
transform 1 0 15272 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_177
timestamp 1608254825
transform 1 0 17388 0 1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_53_170
timestamp 1608254825
transform 1 0 16744 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_166
timestamp 1608254825
transform 1 0 16376 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_12_0_m1_clk_local
timestamp 1608254825
transform 1 0 17112 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__a2111oi_4  _2183_
timestamp 1608254825
transform 1 0 16744 0 -1 31008
box -38 -48 2062 592
use sky130_fd_sc_hd__decap_12  FILLER_53_184
timestamp 1608254825
transform 1 0 18032 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_192
timestamp 1608254825
transform 1 0 18768 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_487
timestamp 1608254825
transform 1 0 17940 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__a2111oi_4  _2232_
timestamp 1608254825
transform 1 0 19136 0 1 31008
box -38 -48 2062 592
use sky130_fd_sc_hd__o21ai_4  _2181_
timestamp 1608254825
transform 1 0 19136 0 -1 31008
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_1  FILLER_53_226
timestamp 1608254825
transform 1 0 21896 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_218
timestamp 1608254825
transform 1 0 21160 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_52_215
timestamp 1608254825
transform 1 0 20884 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_213
timestamp 1608254825
transform 1 0 20700 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_209
timestamp 1608254825
transform 1 0 20332 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_481
timestamp 1608254825
transform 1 0 20792 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_4  _2233_
timestamp 1608254825
transform 1 0 21620 0 -1 31008
box -38 -48 1234 592
use sky130_fd_sc_hd__o21ai_4  _2230_
timestamp 1608254825
transform 1 0 21988 0 1 31008
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_53_240
timestamp 1608254825
transform 1 0 23184 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_244
timestamp 1608254825
transform 1 0 23552 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_236
timestamp 1608254825
transform 1 0 22816 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_488
timestamp 1608254825
transform 1 0 23552 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_4  _2261_
timestamp 1608254825
transform 1 0 23644 0 1 31008
box -38 -48 1234 592
use sky130_fd_sc_hd__a21oi_4  _2237_
timestamp 1608254825
transform 1 0 23644 0 -1 31008
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_53_271
timestamp 1608254825
transform 1 0 26036 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_258
timestamp 1608254825
transform 1 0 24840 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_271
timestamp 1608254825
transform 1 0 26036 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_258
timestamp 1608254825
transform 1 0 24840 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_4  _2260_
timestamp 1608254825
transform 1 0 25208 0 1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  _2236_
timestamp 1608254825
transform 1 0 25208 0 -1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_53_275
timestamp 1608254825
transform 1 0 26404 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_52_276
timestamp 1608254825
transform 1 0 26496 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_0
timestamp 1608254825
transform 1 0 26772 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_482
timestamp 1608254825
transform 1 0 26404 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _1861_
timestamp 1608254825
transform 1 0 26956 0 -1 31008
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_53_292
timestamp 1608254825
transform 1 0 27968 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_288
timestamp 1608254825
transform 1 0 27600 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1439_
timestamp 1608254825
transform 1 0 28336 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2605_
timestamp 1608254825
transform 1 0 27968 0 -1 31008
box -38 -48 1786 592
use sky130_fd_sc_hd__a2bb2o_4  _2150_
timestamp 1608254825
transform 1 0 26496 0 1 31008
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_53_306
timestamp 1608254825
transform 1 0 29256 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_53_304
timestamp 1608254825
transform 1 0 29072 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_300
timestamp 1608254825
transform 1 0 28704 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_315
timestamp 1608254825
transform 1 0 30084 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_311
timestamp 1608254825
transform 1 0 29716 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_addressalyzerBlock.SPI_CLK
timestamp 1608254825
transform 1 0 30176 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_489
timestamp 1608254825
transform 1 0 29164 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2599_
timestamp 1608254825
transform 1 0 29440 0 1 31008
box -38 -48 1786 592
use sky130_fd_sc_hd__o21ai_4  _2238_
timestamp 1608254825
transform 1 0 30452 0 -1 31008
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_53_327
timestamp 1608254825
transform 1 0 31188 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_52_337
timestamp 1608254825
transform 1 0 32108 0 -1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_52_332
timestamp 1608254825
transform 1 0 31648 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_483
timestamp 1608254825
transform 1 0 32016 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_4  _2262_
timestamp 1608254825
transform 1 0 31556 0 1 31008
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_53_362
timestamp 1608254825
transform 1 0 34408 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_348
timestamp 1608254825
transform 1 0 33120 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_344
timestamp 1608254825
transform 1 0 32752 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_52_362
timestamp 1608254825
transform 1 0 34408 0 -1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  _2660_
timestamp 1608254825
transform 1 0 32660 0 -1 31008
box -38 -48 1786 592
use sky130_fd_sc_hd__o21ai_4  _2399_
timestamp 1608254825
transform 1 0 33212 0 1 31008
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_6  FILLER_53_372
timestamp 1608254825
transform 1 0 35328 0 1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_367
timestamp 1608254825
transform 1 0 34868 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_52_385
timestamp 1608254825
transform 1 0 36524 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_381
timestamp 1608254825
transform 1 0 36156 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_490
timestamp 1608254825
transform 1 0 34776 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_4  _1237_
timestamp 1608254825
transform 1 0 34960 0 -1 31008
box -38 -48 1234 592
use sky130_fd_sc_hd__o21ai_4  _1234_
timestamp 1608254825
transform 1 0 35880 0 1 31008
box -38 -48 1234 592
use sky130_fd_sc_hd__or2_4  _1233_
timestamp 1608254825
transform 1 0 36616 0 -1 31008
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _1222_
timestamp 1608254825
transform 1 0 34960 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_391
timestamp 1608254825
transform 1 0 37076 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_52_411
timestamp 1608254825
transform 1 0 38916 0 -1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_52_393
timestamp 1608254825
transform 1 0 37260 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_484
timestamp 1608254825
transform 1 0 37628 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2705_
timestamp 1608254825
transform 1 0 37444 0 1 31008
box -38 -48 1786 592
use sky130_fd_sc_hd__a21oi_4  _1224_
timestamp 1608254825
transform 1 0 37720 0 -1 31008
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_53_414
timestamp 1608254825
transform 1 0 39192 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_417
timestamp 1608254825
transform 1 0 39468 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1608254825
transform -1 0 39836 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1608254825
transform -1 0 39836 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_54_22
timestamp 1608254825
transform 1 0 3128 0 -1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1608254825
transform 1 0 1104 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _2530_
timestamp 1608254825
transform 1 0 1380 0 -1 32096
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  FILLER_54_32
timestamp 1608254825
transform 1 0 4048 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_9_0_m1_clk_local
timestamp 1608254825
transform 1 0 3680 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_491
timestamp 1608254825
transform 1 0 3956 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__a41o_4  _2021_
timestamp 1608254825
transform 1 0 4324 0 -1 32096
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_54_52
timestamp 1608254825
transform 1 0 5888 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_4  _2014_
timestamp 1608254825
transform 1 0 6256 0 -1 32096
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_54_88
timestamp 1608254825
transform 1 0 9200 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_80
timestamp 1608254825
transform 1 0 8464 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_69
timestamp 1608254825
transform 1 0 7452 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1361_
timestamp 1608254825
transform 1 0 8188 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1346_
timestamp 1608254825
transform 1 0 8832 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_107
timestamp 1608254825
transform 1 0 10948 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_492
timestamp 1608254825
transform 1 0 9568 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__nand3_4  _1363_
timestamp 1608254825
transform 1 0 9660 0 -1 32096
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_8  FILLER_54_137
timestamp 1608254825
transform 1 0 13708 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__a41oi_4  _1358_
timestamp 1608254825
transform 1 0 11684 0 -1 32096
box -38 -48 2062 592
use sky130_fd_sc_hd__decap_4  FILLER_54_158
timestamp 1608254825
transform 1 0 15640 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_149
timestamp 1608254825
transform 1 0 14812 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_145
timestamp 1608254825
transform 1 0 14444 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_493
timestamp 1608254825
transform 1 0 15180 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1354_
timestamp 1608254825
transform 1 0 14536 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1345_
timestamp 1608254825
transform 1 0 15272 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__a2111oi_4  _2278_
timestamp 1608254825
transform 1 0 16008 0 -1 32096
box -38 -48 2062 592
use sky130_fd_sc_hd__decap_4  FILLER_54_184
timestamp 1608254825
transform 1 0 18032 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__a2111oi_4  _2208_
timestamp 1608254825
transform 1 0 18400 0 -1 32096
box -38 -48 2062 592
use sky130_fd_sc_hd__decap_4  FILLER_54_228
timestamp 1608254825
transform 1 0 22080 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_210
timestamp 1608254825
transform 1 0 20424 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_494
timestamp 1608254825
transform 1 0 20792 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_4  _2254_
timestamp 1608254825
transform 1 0 20884 0 -1 32096
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_54_235
timestamp 1608254825
transform 1 0 22724 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_4  _2206_
timestamp 1608254825
transform 1 0 23092 0 -1 32096
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _1297_
timestamp 1608254825
transform 1 0 22448 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_54_271
timestamp 1608254825
transform 1 0 26036 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_256
timestamp 1608254825
transform 1 0 24656 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_252
timestamp 1608254825
transform 1 0 24288 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_4  _2229_
timestamp 1608254825
transform 1 0 24748 0 -1 32096
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_54_290
timestamp 1608254825
transform 1 0 27784 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_495
timestamp 1608254825
transform 1 0 26404 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_4  _2180_
timestamp 1608254825
transform 1 0 26496 0 -1 32096
box -38 -48 1326 592
use sky130_fd_sc_hd__and2_4  _1859_
timestamp 1608254825
transform 1 0 28152 0 -1 32096
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_54_315
timestamp 1608254825
transform 1 0 30084 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_305
timestamp 1608254825
transform 1 0 29164 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_301
timestamp 1608254825
transform 1 0 28796 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_4  _2263_
timestamp 1608254825
transform 1 0 29256 0 -1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__and4_4  _2241_
timestamp 1608254825
transform 1 0 30452 0 -1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_54_337
timestamp 1608254825
transform 1 0 32108 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_328
timestamp 1608254825
transform 1 0 31280 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_496
timestamp 1608254825
transform 1 0 32016 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2480_
timestamp 1608254825
transform 1 0 32200 0 -1 32096
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  FILLER_54_365
timestamp 1608254825
transform 1 0 34684 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_54_357
timestamp 1608254825
transform 1 0 33948 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_54_387
timestamp 1608254825
transform 1 0 36708 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _2702_
timestamp 1608254825
transform 1 0 34960 0 -1 32096
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_54_398
timestamp 1608254825
transform 1 0 37720 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_54_395
timestamp 1608254825
transform 1 0 37444 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_497
timestamp 1608254825
transform 1 0 37628 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_4  _1221_
timestamp 1608254825
transform 1 0 37812 0 -1 32096
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_6  FILLER_54_412
timestamp 1608254825
transform 1 0 39008 0 -1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1608254825
transform -1 0 39836 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_55_16
timestamp 1608254825
transform 1 0 2576 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_3
timestamp 1608254825
transform 1 0 1380 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1608254825
transform 1 0 1104 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__and4_4  _2027_
timestamp 1608254825
transform 1 0 1748 0 1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  _1990_
timestamp 1608254825
transform 1 0 2944 0 1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_55_36
timestamp 1608254825
transform 1 0 4416 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_29
timestamp 1608254825
transform 1 0 3772 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__nand4_4  _1992_
timestamp 1608254825
transform 1 0 4784 0 1 32096
box -38 -48 1602 592
use sky130_fd_sc_hd__inv_2  _1991_
timestamp 1608254825
transform 1 0 4140 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_55_57
timestamp 1608254825
transform 1 0 6348 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_498
timestamp 1608254825
transform 1 0 6716 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2535_
timestamp 1608254825
transform 1 0 6808 0 1 32096
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_55_81
timestamp 1608254825
transform 1 0 8556 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2685_
timestamp 1608254825
transform 1 0 8924 0 1 32096
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_55_112
timestamp 1608254825
transform 1 0 11408 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_55_104
timestamp 1608254825
transform 1 0 10672 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1341_
timestamp 1608254825
transform 1 0 11592 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_128
timestamp 1608254825
transform 1 0 12880 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_123
timestamp 1608254825
transform 1 0 12420 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_118
timestamp 1608254825
transform 1 0 11960 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_499
timestamp 1608254825
transform 1 0 12328 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__a41oi_4  _1356_
timestamp 1608254825
transform 1 0 13248 0 1 32096
box -38 -48 2062 592
use sky130_fd_sc_hd__buf_2  _1338_
timestamp 1608254825
transform 1 0 12512 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_154
timestamp 1608254825
transform 1 0 15272 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2687_
timestamp 1608254825
transform 1 0 15640 0 1 32096
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_55_177
timestamp 1608254825
transform 1 0 17388 0 1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_55_197
timestamp 1608254825
transform 1 0 19228 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_500
timestamp 1608254825
transform 1 0 17940 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_4  _2276_
timestamp 1608254825
transform 1 0 18032 0 1 32096
box -38 -48 1234 592
use sky130_fd_sc_hd__a21oi_4  _2209_
timestamp 1608254825
transform 1 0 19596 0 1 32096
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_2  FILLER_55_222
timestamp 1608254825
transform 1 0 21528 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_55_214
timestamp 1608254825
transform 1 0 20792 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_4  _2231_
timestamp 1608254825
transform 1 0 21712 0 1 32096
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_55_249
timestamp 1608254825
transform 1 0 24012 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_243
timestamp 1608254825
transform 1 0 23460 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_55_237
timestamp 1608254825
transform 1 0 22908 0 1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_501
timestamp 1608254825
transform 1 0 23552 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1544_
timestamp 1608254825
transform 1 0 23644 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_55_269
timestamp 1608254825
transform 1 0 25852 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_55_256
timestamp 1608254825
transform 1 0 24656 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_4  _1573_
timestamp 1608254825
transform 1 0 25024 0 1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1291_
timestamp 1608254825
transform 1 0 24380 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_55_292
timestamp 1608254825
transform 1 0 27968 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_277
timestamp 1608254825
transform 1 0 26588 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_4  _2205_
timestamp 1608254825
transform 1 0 26680 0 1 32096
box -38 -48 1326 592
use sky130_fd_sc_hd__buf_2  _2149_
timestamp 1608254825
transform 1 0 28336 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_55_306
timestamp 1608254825
transform 1 0 29256 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_55_304
timestamp 1608254825
transform 1 0 29072 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_300
timestamp 1608254825
transform 1 0 28704 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_502
timestamp 1608254825
transform 1 0 29164 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2602_
timestamp 1608254825
transform 1 0 29440 0 1 32096
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_55_338
timestamp 1608254825
transform 1 0 32200 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_327
timestamp 1608254825
transform 1 0 31188 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__and2_4  _1867_
timestamp 1608254825
transform 1 0 31556 0 1 32096
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_4  _1606_
timestamp 1608254825
transform 1 0 32568 0 1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_55_363
timestamp 1608254825
transform 1 0 34500 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_55_351
timestamp 1608254825
transform 1 0 33396 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_380
timestamp 1608254825
transform 1 0 36064 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_503
timestamp 1608254825
transform 1 0 34776 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_4  _1236_
timestamp 1608254825
transform 1 0 34868 0 1 32096
box -38 -48 1234 592
use sky130_fd_sc_hd__or2_4  _1229_
timestamp 1608254825
transform 1 0 36432 0 1 32096
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_55_391
timestamp 1608254825
transform 1 0 37076 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2577_
timestamp 1608254825
transform 1 0 37444 0 1 32096
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_55_414
timestamp 1608254825
transform 1 0 39192 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1608254825
transform -1 0 39836 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_56_11
timestamp 1608254825
transform 1 0 2116 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_56_3
timestamp 1608254825
transform 1 0 1380 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1608254825
transform 1 0 1104 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_4  _2029_
timestamp 1608254825
transform 1 0 2300 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_38
timestamp 1608254825
transform 1 0 4600 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_56_32
timestamp 1608254825
transform 1 0 4048 0 -1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_56_25
timestamp 1608254825
transform 1 0 3404 0 -1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_504
timestamp 1608254825
transform 1 0 3956 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__and4_4  _2012_
timestamp 1608254825
transform 1 0 4692 0 -1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_56_48
timestamp 1608254825
transform 1 0 5520 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__a41oi_4  _2013_
timestamp 1608254825
transform 1 0 5888 0 -1 33184
box -38 -48 2062 592
use sky130_fd_sc_hd__fill_1  FILLER_56_91
timestamp 1608254825
transform 1 0 9476 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_56_85
timestamp 1608254825
transform 1 0 8924 0 -1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_80
timestamp 1608254825
transform 1 0 8464 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_56_74
timestamp 1608254825
transform 1 0 7912 0 -1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _1293_
timestamp 1608254825
transform 1 0 8556 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_505
timestamp 1608254825
transform 1 0 9568 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__a41oi_4  _1342_
timestamp 1608254825
transform 1 0 9660 0 -1 33184
box -38 -48 2062 592
use sky130_fd_sc_hd__decap_4  FILLER_56_128
timestamp 1608254825
transform 1 0 12880 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_115
timestamp 1608254825
transform 1 0 11684 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_4  _1357_
timestamp 1608254825
transform 1 0 13248 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__and4_4  _1355_
timestamp 1608254825
transform 1 0 12052 0 -1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_56_152
timestamp 1608254825
transform 1 0 15088 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_144
timestamp 1608254825
transform 1 0 14352 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_506
timestamp 1608254825
transform 1 0 15180 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__and4_4  _1263_
timestamp 1608254825
transform 1 0 15272 0 -1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_56_163
timestamp 1608254825
transform 1 0 16100 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_m1_clk_local
timestamp 1608254825
transform 1 0 16468 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_4  _2279_
timestamp 1608254825
transform 1 0 16744 0 -1 33184
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_56_200
timestamp 1608254825
transform 1 0 19504 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_183
timestamp 1608254825
transform 1 0 17940 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_4  _2182_
timestamp 1608254825
transform 1 0 18308 0 -1 33184
box -38 -48 1234 592
use sky130_fd_sc_hd__buf_2  _1269_
timestamp 1608254825
transform 1 0 19872 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_219
timestamp 1608254825
transform 1 0 21252 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_215
timestamp 1608254825
transform 1 0 20884 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_56_208
timestamp 1608254825
transform 1 0 20240 0 -1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_507
timestamp 1608254825
transform 1 0 20792 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_4  _2255_
timestamp 1608254825
transform 1 0 21344 0 -1 33184
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_8  FILLER_56_246
timestamp 1608254825
transform 1 0 23736 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_56_233
timestamp 1608254825
transform 1 0 22540 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_4  _1296_
timestamp 1608254825
transform 1 0 22908 0 -1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_56_273
timestamp 1608254825
transform 1 0 26220 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_56_265
timestamp 1608254825
transform 1 0 25484 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_254
timestamp 1608254825
transform 1 0 24472 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__nand2_4  _1653_
timestamp 1608254825
transform 1 0 24656 0 -1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_56_280
timestamp 1608254825
transform 1 0 26864 0 -1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_508
timestamp 1608254825
transform 1 0 26404 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2608_
timestamp 1608254825
transform 1 0 27416 0 -1 33184
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  _1577_
timestamp 1608254825
transform 1 0 26496 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_309
timestamp 1608254825
transform 1 0 29532 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_305
timestamp 1608254825
transform 1 0 29164 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2612_
timestamp 1608254825
transform 1 0 29624 0 -1 33184
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_56_337
timestamp 1608254825
transform 1 0 32108 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_329
timestamp 1608254825
transform 1 0 31372 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_addressalyzerBlock.SPI_CLK
timestamp 1608254825
transform 1 0 31740 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_509
timestamp 1608254825
transform 1 0 32016 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_4  _2215_
timestamp 1608254825
transform 1 0 32200 0 -1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_56_359
timestamp 1608254825
transform 1 0 34132 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_347
timestamp 1608254825
transform 1 0 33028 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__o21ai_4  _1231_
timestamp 1608254825
transform 1 0 34224 0 -1 33184
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_1  FILLER_56_379
timestamp 1608254825
transform 1 0 35972 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_56_373
timestamp 1608254825
transform 1 0 35420 0 -1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_4  _1230_
timestamp 1608254825
transform 1 0 36064 0 -1 33184
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_6  FILLER_56_411
timestamp 1608254825
transform 1 0 38916 0 -1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_56_398
timestamp 1608254825
transform 1 0 37720 0 -1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_56_393
timestamp 1608254825
transform 1 0 37260 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_510
timestamp 1608254825
transform 1 0 37628 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _1220_
timestamp 1608254825
transform 1 0 38272 0 -1 33184
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_56_417
timestamp 1608254825
transform 1 0 39468 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1608254825
transform -1 0 39836 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_57_12
timestamp 1608254825
transform 1 0 2208 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1608254825
transform 1 0 1104 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_4  _2033_
timestamp 1608254825
transform 1 0 1380 0 1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__a41oi_4  _2028_
timestamp 1608254825
transform 1 0 2576 0 1 33184
box -38 -48 2062 592
use sky130_fd_sc_hd__decap_4  FILLER_57_38
timestamp 1608254825
transform 1 0 4600 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__and3_4  _2023_
timestamp 1608254825
transform 1 0 4968 0 1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_57_62
timestamp 1608254825
transform 1 0 6808 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_57_59
timestamp 1608254825
transform 1 0 6532 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_57_51
timestamp 1608254825
transform 1 0 5796 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_511
timestamp 1608254825
transform 1 0 6716 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _2006_
timestamp 1608254825
transform 1 0 7176 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_57_83
timestamp 1608254825
transform 1 0 8740 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_57_77
timestamp 1608254825
transform 1 0 8188 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_57_69
timestamp 1608254825
transform 1 0 7452 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1364_
timestamp 1608254825
transform 1 0 8464 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_4  _1343_
timestamp 1608254825
transform 1 0 9108 0 1 33184
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_57_100
timestamp 1608254825
transform 1 0 10304 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_4  _1339_
timestamp 1608254825
transform 1 0 10672 0 1 33184
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_57_132
timestamp 1608254825
transform 1 0 13248 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_118
timestamp 1608254825
transform 1 0 11960 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_512
timestamp 1608254825
transform 1 0 12328 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__and4_4  _1333_
timestamp 1608254825
transform 1 0 12420 0 1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _1278_
timestamp 1608254825
transform 1 0 13616 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_154
timestamp 1608254825
transform 1 0 15272 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_144
timestamp 1608254825
transform 1 0 14352 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_140
timestamp 1608254825
transform 1 0 13984 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2694_
timestamp 1608254825
transform 1 0 15640 0 1 33184
box -38 -48 1786 592
use sky130_fd_sc_hd__nand2_4  _1315_
timestamp 1608254825
transform 1 0 14444 0 1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_57_177
timestamp 1608254825
transform 1 0 17388 0 1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_204
timestamp 1608254825
transform 1 0 19872 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_197
timestamp 1608254825
transform 1 0 19228 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_m1_clk_local
timestamp 1608254825
transform 1 0 19596 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_513
timestamp 1608254825
transform 1 0 17940 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_4  _2277_
timestamp 1608254825
transform 1 0 18032 0 1 33184
box -38 -48 1234 592
use sky130_fd_sc_hd__a21oi_4  _2207_
timestamp 1608254825
transform 1 0 19964 0 1 33184
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_57_218
timestamp 1608254825
transform 1 0 21160 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_m1_clk_local
timestamp 1608254825
transform 1 0 21528 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_4  _1294_
timestamp 1608254825
transform 1 0 21804 0 1 33184
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_6  FILLER_57_238
timestamp 1608254825
transform 1 0 23000 0 1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_514
timestamp 1608254825
transform 1 0 23552 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2698_
timestamp 1608254825
transform 1 0 23644 0 1 33184
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_57_264
timestamp 1608254825
transform 1 0 25392 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_2
timestamp 1608254825
transform 1 0 25576 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _1843_
timestamp 1608254825
transform 1 0 25760 0 1 33184
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_57_293
timestamp 1608254825
transform 1 0 28060 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_275
timestamp 1608254825
transform 1 0 26404 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_4  _2275_
timestamp 1608254825
transform 1 0 26772 0 1 33184
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_2  FILLER_57_315
timestamp 1608254825
transform 1 0 30084 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_301
timestamp 1608254825
transform 1 0 28796 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_1
timestamp 1608254825
transform 1 0 29900 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_515
timestamp 1608254825
transform 1 0 29164 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1860_
timestamp 1608254825
transform 1 0 28428 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__and2_4  _1855_
timestamp 1608254825
transform 1 0 30268 0 1 33184
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _1845_
timestamp 1608254825
transform 1 0 29256 0 1 33184
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_57_342
timestamp 1608254825
transform 1 0 32568 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_338
timestamp 1608254825
transform 1 0 32200 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_328
timestamp 1608254825
transform 1 0 31280 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_324
timestamp 1608254825
transform 1 0 30912 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_4  _2216_
timestamp 1608254825
transform 1 0 31372 0 1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_57_362
timestamp 1608254825
transform 1 0 34408 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2481_
timestamp 1608254825
transform 1 0 32660 0 1 33184
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_57_388
timestamp 1608254825
transform 1 0 36800 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_380
timestamp 1608254825
transform 1 0 36064 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_516
timestamp 1608254825
transform 1 0 34776 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_4  _1227_
timestamp 1608254825
transform 1 0 34868 0 1 33184
box -38 -48 1234 592
use sky130_fd_sc_hd__buf_2  _1208_
timestamp 1608254825
transform 1 0 36432 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_405
timestamp 1608254825
transform 1 0 38364 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_4  _1226_
timestamp 1608254825
transform 1 0 37168 0 1 33184
box -38 -48 1234 592
use sky130_fd_sc_hd__buf_2  _1201_
timestamp 1608254825
transform 1 0 38732 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_417
timestamp 1608254825
transform 1 0 39468 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_413
timestamp 1608254825
transform 1 0 39100 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1608254825
transform -1 0 39836 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_58_3
timestamp 1608254825
transform 1 0 1380 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1608254825
transform 1 0 1104 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _2531_
timestamp 1608254825
transform 1 0 1564 0 -1 34272
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_58_30
timestamp 1608254825
transform 1 0 3864 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_58_24
timestamp 1608254825
transform 1 0 3312 0 -1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_517
timestamp 1608254825
transform 1 0 3956 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2532_
timestamp 1608254825
transform 1 0 4048 0 -1 34272
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_58_57
timestamp 1608254825
transform 1 0 6348 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_58_51
timestamp 1608254825
transform 1 0 5796 0 -1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_4  _1999_
timestamp 1608254825
transform 1 0 6440 0 -1 34272
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_58_88
timestamp 1608254825
transform 1 0 9200 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_84
timestamp 1608254825
transform 1 0 8832 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_58_78
timestamp 1608254825
transform 1 0 8280 0 -1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_58_71
timestamp 1608254825
transform 1 0 7636 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1998_
timestamp 1608254825
transform 1 0 8004 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1344_
timestamp 1608254825
transform 1 0 8924 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_58_98
timestamp 1608254825
transform 1 0 10120 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_58_93
timestamp 1608254825
transform 1 0 9660 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_518
timestamp 1608254825
transform 1 0 9568 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1340_
timestamp 1608254825
transform 1 0 9844 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__nand4_4  _1335_
timestamp 1608254825
transform 1 0 10488 0 -1 34272
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_58_119
timestamp 1608254825
transform 1 0 12052 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__nand4_4  _1266_
timestamp 1608254825
transform 1 0 12420 0 -1 34272
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_2  FILLER_58_154
timestamp 1608254825
transform 1 0 15272 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_58_152
timestamp 1608254825
transform 1 0 15088 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_140
timestamp 1608254825
transform 1 0 13984 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_519
timestamp 1608254825
transform 1 0 15180 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_4  _1312_
timestamp 1608254825
transform 1 0 15456 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_182
timestamp 1608254825
transform 1 0 17848 0 -1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_58_175
timestamp 1608254825
transform 1 0 17204 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_168
timestamp 1608254825
transform 1 0 16560 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1320_
timestamp 1608254825
transform 1 0 17572 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1316_
timestamp 1608254825
transform 1 0 16928 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _2697_
timestamp 1608254825
transform 1 0 18400 0 -1 34272
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_58_213
timestamp 1608254825
transform 1 0 20700 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_58_207
timestamp 1608254825
transform 1 0 20148 0 -1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_520
timestamp 1608254825
transform 1 0 20792 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__nand4_4  _1290_
timestamp 1608254825
transform 1 0 20884 0 -1 34272
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_58_245
timestamp 1608254825
transform 1 0 23644 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_232
timestamp 1608254825
transform 1 0 22448 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_14_0_m1_clk_local
timestamp 1608254825
transform 1 0 24012 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_4  _1270_
timestamp 1608254825
transform 1 0 22816 0 -1 34272
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_58_271
timestamp 1608254825
transform 1 0 26036 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2622_
timestamp 1608254825
transform 1 0 24288 0 -1 34272
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_58_295
timestamp 1608254825
transform 1 0 28244 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_521
timestamp 1608254825
transform 1 0 26404 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2614_
timestamp 1608254825
transform 1 0 26496 0 -1 34272
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_58_318
timestamp 1608254825
transform 1 0 30360 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2620_
timestamp 1608254825
transform 1 0 28612 0 -1 34272
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_58_335
timestamp 1608254825
transform 1 0 31924 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_58_329
timestamp 1608254825
transform 1 0 31372 0 -1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_522
timestamp 1608254825
transform 1 0 32016 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2482_
timestamp 1608254825
transform 1 0 32108 0 -1 34272
box -38 -48 1786 592
use sky130_fd_sc_hd__and2_4  _1870_
timestamp 1608254825
transform 1 0 30728 0 -1 34272
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_58_356
timestamp 1608254825
transform 1 0 33856 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_4  _2240_
timestamp 1608254825
transform 1 0 34224 0 -1 34272
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_58_369
timestamp 1608254825
transform 1 0 35052 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2703_
timestamp 1608254825
transform 1 0 35420 0 -1 34272
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_58_411
timestamp 1608254825
transform 1 0 38916 0 -1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_396
timestamp 1608254825
transform 1 0 37536 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_392
timestamp 1608254825
transform 1 0 37168 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_523
timestamp 1608254825
transform 1 0 37628 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_4  _1228_
timestamp 1608254825
transform 1 0 37720 0 -1 34272
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_1  FILLER_58_417
timestamp 1608254825
transform 1 0 39468 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1608254825
transform -1 0 39836 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_60_15
timestamp 1608254825
transform 1 0 2484 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_3
timestamp 1608254825
transform 1 0 1380 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_15
timestamp 1608254825
transform 1 0 2484 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_3
timestamp 1608254825
transform 1 0 1380 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1608254825
transform 1 0 1104 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1608254825
transform 1 0 1104 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_60_27
timestamp 1608254825
transform 1 0 3588 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_59_42
timestamp 1608254825
transform 1 0 4968 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_59_34
timestamp 1608254825
transform 1 0 4232 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_59_27
timestamp 1608254825
transform 1 0 3588 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_530
timestamp 1608254825
transform 1 0 3956 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2533_
timestamp 1608254825
transform 1 0 4048 0 -1 35360
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  _2026_
timestamp 1608254825
transform 1 0 3864 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_4  _2016_
timestamp 1608254825
transform 1 0 5152 0 1 34272
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_1  FILLER_60_67
timestamp 1608254825
transform 1 0 7268 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_60_59
timestamp 1608254825
transform 1 0 6532 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_60_51
timestamp 1608254825
transform 1 0 5796 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_57
timestamp 1608254825
transform 1 0 6348 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_524
timestamp 1608254825
transform 1 0 6716 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__nand3_4  _2017_
timestamp 1608254825
transform 1 0 7360 0 -1 35360
box -38 -48 1326 592
use sky130_fd_sc_hd__nor4_4  _2008_
timestamp 1608254825
transform 1 0 6808 0 1 34272
box -38 -48 1602 592
use sky130_fd_sc_hd__buf_2  _1997_
timestamp 1608254825
transform 1 0 6164 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_60_90
timestamp 1608254825
transform 1 0 9384 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_60_82
timestamp 1608254825
transform 1 0 8648 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_59_87
timestamp 1608254825
transform 1 0 9108 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_79
timestamp 1608254825
transform 1 0 8372 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _2689_
timestamp 1608254825
transform 1 0 9200 0 1 34272
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_60_103
timestamp 1608254825
transform 1 0 10580 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_96
timestamp 1608254825
transform 1 0 9936 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_107
timestamp 1608254825
transform 1 0 10948 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_531
timestamp 1608254825
transform 1 0 9568 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2690_
timestamp 1608254825
transform 1 0 10948 0 -1 35360
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_2  _2018_
timestamp 1608254825
transform 1 0 10304 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2015_
timestamp 1608254825
transform 1 0 9660 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1332_
timestamp 1608254825
transform 1 0 11316 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_126
timestamp 1608254825
transform 1 0 12696 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_126
timestamp 1608254825
transform 1 0 12696 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_121
timestamp 1608254825
transform 1 0 12236 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_59_115
timestamp 1608254825
transform 1 0 11684 0 1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_525
timestamp 1608254825
transform 1 0 12328 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__nand4_4  _1280_
timestamp 1608254825
transform 1 0 13064 0 1 34272
box -38 -48 1602 592
use sky130_fd_sc_hd__inv_2  _1265_
timestamp 1608254825
transform 1 0 12420 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_4  _1264_
timestamp 1608254825
transform 1 0 13064 0 -1 35360
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_60_154
timestamp 1608254825
transform 1 0 15272 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_60_147
timestamp 1608254825
transform 1 0 14628 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_60_139
timestamp 1608254825
transform 1 0 13892 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_59_147
timestamp 1608254825
transform 1 0 14628 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_13_0_m1_clk_local
timestamp 1608254825
transform 1 0 14904 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_532
timestamp 1608254825
transform 1 0 15180 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__nand4_4  _1314_
timestamp 1608254825
transform 1 0 14996 0 1 34272
box -38 -48 1602 592
use sky130_fd_sc_hd__nor2_4  _1310_
timestamp 1608254825
transform 1 0 15640 0 -1 35360
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_60_167
timestamp 1608254825
transform 1 0 16468 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_59_175
timestamp 1608254825
transform 1 0 17204 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_59_168
timestamp 1608254825
transform 1 0 16560 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2693_
timestamp 1608254825
transform 1 0 16836 0 -1 35360
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_2  _1309_
timestamp 1608254825
transform 1 0 16928 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_60_203
timestamp 1608254825
transform 1 0 19780 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_60_190
timestamp 1608254825
transform 1 0 18584 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_200
timestamp 1608254825
transform 1 0 19504 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_59_184
timestamp 1608254825
transform 1 0 18032 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_526
timestamp 1608254825
transform 1 0 17940 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__nor3_4  _1302_
timestamp 1608254825
transform 1 0 18308 0 1 34272
box -38 -48 1234 592
use sky130_fd_sc_hd__a21oi_4  _1301_
timestamp 1608254825
transform 1 0 19872 0 1 34272
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_4  _1248_
timestamp 1608254825
transform 1 0 18952 0 -1 35360
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_60_224
timestamp 1608254825
transform 1 0 21712 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_60_211
timestamp 1608254825
transform 1 0 20516 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_59_217
timestamp 1608254825
transform 1 0 21068 0 1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_15_0_m1_clk_local
timestamp 1608254825
transform 1 0 22080 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_533
timestamp 1608254825
transform 1 0 20792 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__and4_4  _1300_
timestamp 1608254825
transform 1 0 20884 0 -1 35360
box -38 -48 866 592
use sky130_fd_sc_hd__nand4_4  _1295_
timestamp 1608254825
transform 1 0 21620 0 1 34272
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_60_248
timestamp 1608254825
transform 1 0 23920 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_249
timestamp 1608254825
transform 1 0 24012 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_240
timestamp 1608254825
transform 1 0 23184 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_527
timestamp 1608254825
transform 1 0 23552 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1574_
timestamp 1608254825
transform 1 0 23644 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__nand4_4  _1288_
timestamp 1608254825
transform 1 0 22356 0 -1 35360
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_60_271
timestamp 1608254825
transform 1 0 26036 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_263
timestamp 1608254825
transform 1 0 25300 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_60_255
timestamp 1608254825
transform 1 0 24564 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_272
timestamp 1608254825
transform 1 0 26128 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_59_260
timestamp 1608254825
transform 1 0 25024 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _2611_
timestamp 1608254825
transform 1 0 26312 0 1 34272
box -38 -48 1786 592
use sky130_fd_sc_hd__and2_4  _1856_
timestamp 1608254825
transform 1 0 25392 0 -1 35360
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _1846_
timestamp 1608254825
transform 1 0 24380 0 1 34272
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1271_
timestamp 1608254825
transform 1 0 24288 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_60_292
timestamp 1608254825
transform 1 0 27968 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_287
timestamp 1608254825
transform 1 0 27508 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_283
timestamp 1608254825
transform 1 0 27140 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_293
timestamp 1608254825
transform 1 0 28060 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_534
timestamp 1608254825
transform 1 0 26404 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _1871_
timestamp 1608254825
transform 1 0 28336 0 -1 35360
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _1852_
timestamp 1608254825
transform 1 0 26496 0 -1 35360
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _1848_
timestamp 1608254825
transform 1 0 27600 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_303
timestamp 1608254825
transform 1 0 28980 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_319
timestamp 1608254825
transform 1 0 30452 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_59_306
timestamp 1608254825
transform 1 0 29256 0 1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_59_301
timestamp 1608254825
transform 1 0 28796 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_528
timestamp 1608254825
transform 1 0 29164 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2598_
timestamp 1608254825
transform 1 0 29348 0 -1 35360
box -38 -48 1786 592
use sky130_fd_sc_hd__and2_4  _1869_
timestamp 1608254825
transform 1 0 29808 0 1 34272
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _1838_
timestamp 1608254825
transform 1 0 28428 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_332
timestamp 1608254825
transform 1 0 31648 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_60_326
timestamp 1608254825
transform 1 0 31096 0 -1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_59_340
timestamp 1608254825
transform 1 0 32384 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_327
timestamp 1608254825
transform 1 0 31188 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_11_0_addressalyzerBlock.SPI_CLK
timestamp 1608254825
transform 1 0 31740 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_535
timestamp 1608254825
transform 1 0 32016 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2615_
timestamp 1608254825
transform 1 0 32108 0 -1 35360
box -38 -48 1786 592
use sky130_fd_sc_hd__nand2_4  _2264_
timestamp 1608254825
transform 1 0 31556 0 1 34272
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _1839_
timestamp 1608254825
transform 1 0 30820 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_356
timestamp 1608254825
transform 1 0 33856 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_365
timestamp 1608254825
transform 1 0 34684 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_353
timestamp 1608254825
transform 1 0 33580 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _2616_
timestamp 1608254825
transform 1 0 34224 0 -1 35360
box -38 -48 1786 592
use sky130_fd_sc_hd__nand2_4  _2239_
timestamp 1608254825
transform 1 0 32752 0 1 34272
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_60_379
timestamp 1608254825
transform 1 0 35972 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_385
timestamp 1608254825
transform 1 0 36524 0 1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_371
timestamp 1608254825
transform 1 0 35236 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_367
timestamp 1608254825
transform 1 0 34868 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_529
timestamp 1608254825
transform 1 0 34776 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_4  _1232_
timestamp 1608254825
transform 1 0 35328 0 1 34272
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_8  FILLER_60_408
timestamp 1608254825
transform 1 0 38640 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_60_398
timestamp 1608254825
transform 1 0 37720 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_60_391
timestamp 1608254825
transform 1 0 37076 0 -1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_59_410
timestamp 1608254825
transform 1 0 38824 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_536
timestamp 1608254825
transform 1 0 37628 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2704_
timestamp 1608254825
transform 1 0 37076 0 1 34272
box -38 -48 1786 592
use sky130_fd_sc_hd__or2_4  _1225_
timestamp 1608254825
transform 1 0 37996 0 -1 35360
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_60_416
timestamp 1608254825
transform 1 0 39376 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1608254825
transform -1 0 39836 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1608254825
transform -1 0 39836 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_61_15
timestamp 1608254825
transform 1 0 2484 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_3
timestamp 1608254825
transform 1 0 1380 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1608254825
transform 1 0 1104 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_61_43
timestamp 1608254825
transform 1 0 5060 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_61_27
timestamp 1608254825
transform 1 0 3588 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_4  _2019_
timestamp 1608254825
transform 1 0 3864 0 1 35360
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_6  FILLER_61_66
timestamp 1608254825
transform 1 0 7176 0 1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_61_57
timestamp 1608254825
transform 1 0 6348 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_47
timestamp 1608254825
transform 1 0 5428 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_537
timestamp 1608254825
transform 1 0 6716 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _2007_
timestamp 1608254825
transform 1 0 6808 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_4  _1993_
timestamp 1608254825
transform 1 0 5520 0 1 35360
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_61_72
timestamp 1608254825
transform 1 0 7728 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2534_
timestamp 1608254825
transform 1 0 7820 0 1 35360
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_61_105
timestamp 1608254825
transform 1 0 10764 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_61_100
timestamp 1608254825
transform 1 0 10304 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_61_92
timestamp 1608254825
transform 1 0 9568 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1337_
timestamp 1608254825
transform 1 0 10488 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_4  _1336_
timestamp 1608254825
transform 1 0 11132 0 1 35360
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_61_135
timestamp 1608254825
transform 1 0 13524 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_118
timestamp 1608254825
transform 1 0 11960 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_538
timestamp 1608254825
transform 1 0 12328 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_4  _1334_
timestamp 1608254825
transform 1 0 12420 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_61_147
timestamp 1608254825
transform 1 0 14628 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_4  _1317_
timestamp 1608254825
transform 1 0 14904 0 1 35360
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_6  FILLER_61_177
timestamp 1608254825
transform 1 0 17388 0 1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_61_164
timestamp 1608254825
transform 1 0 16192 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_4  _1318_
timestamp 1608254825
transform 1 0 16560 0 1 35360
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_61_197
timestamp 1608254825
transform 1 0 19228 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_539
timestamp 1608254825
transform 1 0 17940 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__nor3_4  _1304_
timestamp 1608254825
transform 1 0 18032 0 1 35360
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_4  _1285_
timestamp 1608254825
transform 1 0 19596 0 1 35360
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_61_210
timestamp 1608254825
transform 1 0 20424 0 1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__a41o_4  _1286_
timestamp 1608254825
transform 1 0 20976 0 1 35360
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_8  FILLER_61_249
timestamp 1608254825
transform 1 0 24012 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_61_241
timestamp 1608254825
transform 1 0 23276 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_61_233
timestamp 1608254825
transform 1 0 22540 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_540
timestamp 1608254825
transform 1 0 23552 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1268_
timestamp 1608254825
transform 1 0 23644 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2619_
timestamp 1608254825
transform 1 0 24748 0 1 35360
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_61_291
timestamp 1608254825
transform 1 0 27876 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_61_276
timestamp 1608254825
transform 1 0 26496 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_10_0_addressalyzerBlock.SPI_CLK
timestamp 1608254825
transform 1 0 27232 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1854_
timestamp 1608254825
transform 1 0 27508 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1842_
timestamp 1608254825
transform 1 0 28244 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_306
timestamp 1608254825
transform 1 0 29256 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_61_299
timestamp 1608254825
transform 1 0 28612 0 1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_addressalyzerBlock.SPI_CLK
timestamp 1608254825
transform 1 0 29624 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_541
timestamp 1608254825
transform 1 0 29164 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2600_
timestamp 1608254825
transform 1 0 29900 0 1 35360
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_61_332
timestamp 1608254825
transform 1 0 31648 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2623_
timestamp 1608254825
transform 1 0 32016 0 1 35360
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  FILLER_61_363
timestamp 1608254825
transform 1 0 34500 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_61_355
timestamp 1608254825
transform 1 0 33764 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_61_386
timestamp 1608254825
transform 1 0 36616 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_542
timestamp 1608254825
transform 1 0 34776 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2624_
timestamp 1608254825
transform 1 0 34868 0 1 35360
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_61_410
timestamp 1608254825
transform 1 0 38824 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_61_398
timestamp 1608254825
transform 1 0 37720 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1608254825
transform -1 0 39836 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_62_15
timestamp 1608254825
transform 1 0 2484 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_3
timestamp 1608254825
transform 1 0 1380 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1608254825
transform 1 0 1104 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_62_45
timestamp 1608254825
transform 1 0 5244 0 -1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_62_27
timestamp 1608254825
transform 1 0 3588 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_543
timestamp 1608254825
transform 1 0 3956 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_4  _2020_
timestamp 1608254825
transform 1 0 4048 0 -1 36448
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_1  FILLER_62_51
timestamp 1608254825
transform 1 0 5796 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__nand4_4  _1994_
timestamp 1608254825
transform 1 0 5888 0 -1 36448
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_1  FILLER_62_91
timestamp 1608254825
transform 1 0 9476 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_83
timestamp 1608254825
transform 1 0 8740 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_62_76
timestamp 1608254825
transform 1 0 8096 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_69
timestamp 1608254825
transform 1 0 7452 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2003_
timestamp 1608254825
transform 1 0 8464 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1979_
timestamp 1608254825
transform 1 0 7820 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_62_112
timestamp 1608254825
transform 1 0 11408 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_544
timestamp 1608254825
transform 1 0 9568 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2551_
timestamp 1608254825
transform 1 0 9660 0 -1 36448
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_62_133
timestamp 1608254825
transform 1 0 13340 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_4  _1323_
timestamp 1608254825
transform 1 0 13708 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_4  _1322_
timestamp 1608254825
transform 1 0 12512 0 -1 36448
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_62_157
timestamp 1608254825
transform 1 0 15548 0 -1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_62_149
timestamp 1608254825
transform 1 0 14812 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_545
timestamp 1608254825
transform 1 0 15180 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1279_
timestamp 1608254825
transform 1 0 15272 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_62_177
timestamp 1608254825
transform 1 0 17388 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__nand3_4  _1319_
timestamp 1608254825
transform 1 0 16100 0 -1 36448
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_62_188
timestamp 1608254825
transform 1 0 18400 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1276_
timestamp 1608254825
transform 1 0 18124 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__nor4_4  _1267_
timestamp 1608254825
transform 1 0 18768 0 -1 36448
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_62_228
timestamp 1608254825
transform 1 0 22080 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_213
timestamp 1608254825
transform 1 0 20700 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_209
timestamp 1608254825
transform 1 0 20332 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_546
timestamp 1608254825
transform 1 0 20792 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_4  _1306_
timestamp 1608254825
transform 1 0 20884 0 -1 36448
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_62_242
timestamp 1608254825
transform 1 0 23368 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_232
timestamp 1608254825
transform 1 0 22448 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2699_
timestamp 1608254825
transform 1 0 23736 0 -1 36448
box -38 -48 1786 592
use sky130_fd_sc_hd__and3_4  _1289_
timestamp 1608254825
transform 1 0 22540 0 -1 36448
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_62_273
timestamp 1608254825
transform 1 0 26220 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_62_265
timestamp 1608254825
transform 1 0 25484 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_62_283
timestamp 1608254825
transform 1 0 27140 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_547
timestamp 1608254825
transform 1 0 26404 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2609_
timestamp 1608254825
transform 1 0 27508 0 -1 36448
box -38 -48 1786 592
use sky130_fd_sc_hd__and2_4  _1857_
timestamp 1608254825
transform 1 0 26496 0 -1 36448
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  FILLER_62_314
timestamp 1608254825
transform 1 0 29992 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_62_306
timestamp 1608254825
transform 1 0 29256 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__and2_4  _1841_
timestamp 1608254825
transform 1 0 30268 0 -1 36448
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_62_337
timestamp 1608254825
transform 1 0 32108 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_62_324
timestamp 1608254825
transform 1 0 30912 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_548
timestamp 1608254825
transform 1 0 32016 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_363
timestamp 1608254825
transform 1 0 34500 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_352
timestamp 1608254825
transform 1 0 33488 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__and2_4  _1851_
timestamp 1608254825
transform 1 0 33856 0 -1 36448
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _1850_
timestamp 1608254825
transform 1 0 32844 0 -1 36448
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_62_387
timestamp 1608254825
transform 1 0 36708 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_62_375
timestamp 1608254825
transform 1 0 35604 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_367
timestamp 1608254825
transform 1 0 34868 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _1840_
timestamp 1608254825
transform 1 0 34960 0 -1 36448
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_62_410
timestamp 1608254825
transform 1 0 38824 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_62_398
timestamp 1608254825
transform 1 0 37720 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_62_395
timestamp 1608254825
transform 1 0 37444 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_549
timestamp 1608254825
transform 1 0 37628 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1608254825
transform -1 0 39836 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_63_22
timestamp 1608254825
transform 1 0 3128 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1608254825
transform 1 0 1104 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _2550_
timestamp 1608254825
transform 1 0 1380 0 1 36448
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_63_34
timestamp 1608254825
transform 1 0 4232 0 1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__a41o_4  _2004_
timestamp 1608254825
transform 1 0 4784 0 1 36448
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_3  FILLER_63_62
timestamp 1608254825
transform 1 0 6808 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_63_57
timestamp 1608254825
transform 1 0 6348 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_550
timestamp 1608254825
transform 1 0 6716 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__nand4_4  _2000_
timestamp 1608254825
transform 1 0 7084 0 1 36448
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_2  FILLER_63_90
timestamp 1608254825
transform 1 0 9384 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_63_82
timestamp 1608254825
transform 1 0 8648 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_63_101
timestamp 1608254825
transform 1 0 10396 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_4  _1956_
timestamp 1608254825
transform 1 0 9568 0 1 36448
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  _1329_
timestamp 1608254825
transform 1 0 11132 0 1 36448
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_63_137
timestamp 1608254825
transform 1 0 13708 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_63_118
timestamp 1608254825
transform 1 0 11960 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_551
timestamp 1608254825
transform 1 0 12328 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__nand3_4  _1330_
timestamp 1608254825
transform 1 0 12420 0 1 36448
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_2  FILLER_63_145
timestamp 1608254825
transform 1 0 14444 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _2692_
timestamp 1608254825
transform 1 0 14628 0 1 36448
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_63_179
timestamp 1608254825
transform 1 0 17572 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_166
timestamp 1608254825
transform 1 0 16376 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_4  _1247_
timestamp 1608254825
transform 1 0 16744 0 1 36448
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_63_203
timestamp 1608254825
transform 1 0 19780 0 1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_552
timestamp 1608254825
transform 1 0 17940 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2696_
timestamp 1608254825
transform 1 0 18032 0 1 36448
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_63_220
timestamp 1608254825
transform 1 0 21344 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_212
timestamp 1608254825
transform 1 0 20608 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__nand4_4  _1282_
timestamp 1608254825
transform 1 0 21436 0 1 36448
box -38 -48 1602 592
use sky130_fd_sc_hd__inv_2  _1246_
timestamp 1608254825
transform 1 0 20332 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_63_251
timestamp 1608254825
transform 1 0 24196 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_63_245
timestamp 1608254825
transform 1 0 23644 0 1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_63_238
timestamp 1608254825
transform 1 0 23000 0 1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_553
timestamp 1608254825
transform 1 0 23552 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_63_267
timestamp 1608254825
transform 1 0 25668 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_259
timestamp 1608254825
transform 1 0 24932 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _2610_
timestamp 1608254825
transform 1 0 25760 0 1 36448
box -38 -48 1786 592
use sky130_fd_sc_hd__and2_4  _1844_
timestamp 1608254825
transform 1 0 24288 0 1 36448
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_63_293
timestamp 1608254825
transform 1 0 28060 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_63_287
timestamp 1608254825
transform 1 0 27508 0 1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__and2_4  _1858_
timestamp 1608254825
transform 1 0 28152 0 1 36448
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_63_301
timestamp 1608254825
transform 1 0 28796 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_554
timestamp 1608254825
transform 1 0 29164 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2606_
timestamp 1608254825
transform 1 0 29256 0 1 36448
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_63_337
timestamp 1608254825
transform 1 0 32108 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_63_325
timestamp 1608254825
transform 1 0 31004 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__and2_4  _1849_
timestamp 1608254825
transform 1 0 32476 0 1 36448
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_63_360
timestamp 1608254825
transform 1 0 34224 0 1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_63_348
timestamp 1608254825
transform 1 0 33120 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_379
timestamp 1608254825
transform 1 0 35972 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_367
timestamp 1608254825
transform 1 0 34868 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_555
timestamp 1608254825
transform 1 0 34776 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_403
timestamp 1608254825
transform 1 0 38180 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_391
timestamp 1608254825
transform 1 0 37076 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_63_415
timestamp 1608254825
transform 1 0 39284 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1608254825
transform -1 0 39836 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_15
timestamp 1608254825
transform 1 0 2484 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_3
timestamp 1608254825
transform 1 0 1380 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1608254825
transform 1 0 1104 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_64_45
timestamp 1608254825
transform 1 0 5244 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_32
timestamp 1608254825
transform 1 0 4048 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_27
timestamp 1608254825
transform 1 0 3588 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_556
timestamp 1608254825
transform 1 0 3956 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__and3_4  _2005_
timestamp 1608254825
transform 1 0 4416 0 -1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_64_68
timestamp 1608254825
transform 1 0 7360 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  _2536_
timestamp 1608254825
transform 1 0 5612 0 -1 37536
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_64_88
timestamp 1608254825
transform 1 0 9200 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_4  _2001_
timestamp 1608254825
transform 1 0 7912 0 -1 37536
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_64_96
timestamp 1608254825
transform 1 0 9936 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_557
timestamp 1608254825
transform 1 0 9568 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2589_
timestamp 1608254825
transform 1 0 10304 0 -1 37536
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_2  _1995_
timestamp 1608254825
transform 1 0 9660 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_64_131
timestamp 1608254825
transform 1 0 13156 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_127
timestamp 1608254825
transform 1 0 12788 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_119
timestamp 1608254825
transform 1 0 12052 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1327_
timestamp 1608254825
transform 1 0 12880 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_4  _1324_
timestamp 1608254825
transform 1 0 13524 0 -1 37536
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_64_159
timestamp 1608254825
transform 1 0 15732 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_154
timestamp 1608254825
transform 1 0 15272 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_149
timestamp 1608254825
transform 1 0 14812 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_558
timestamp 1608254825
transform 1 0 15180 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1313_
timestamp 1608254825
transform 1 0 15456 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_64_163
timestamp 1608254825
transform 1 0 16100 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2575_
timestamp 1608254825
transform 1 0 16192 0 -1 37536
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_64_183
timestamp 1608254825
transform 1 0 17940 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__nor4_4  _1281_
timestamp 1608254825
transform 1 0 18492 0 -1 37536
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_64_226
timestamp 1608254825
transform 1 0 21896 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_222
timestamp 1608254825
transform 1 0 21528 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_218
timestamp 1608254825
transform 1 0 21160 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_206
timestamp 1608254825
transform 1 0 20056 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_559
timestamp 1608254825
transform 1 0 20792 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1305_
timestamp 1608254825
transform 1 0 20884 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1284_
timestamp 1608254825
transform 1 0 21620 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_64_251
timestamp 1608254825
transform 1 0 24196 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_247
timestamp 1608254825
transform 1 0 23828 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__a41o_4  _1272_
timestamp 1608254825
transform 1 0 22264 0 -1 37536
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_64_271
timestamp 1608254825
transform 1 0 26036 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2618_
timestamp 1608254825
transform 1 0 24288 0 -1 37536
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_64_284
timestamp 1608254825
transform 1 0 27232 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_276
timestamp 1608254825
transform 1 0 26496 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_560
timestamp 1608254825
transform 1 0 26404 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2604_
timestamp 1608254825
transform 1 0 27324 0 -1 37536
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_64_304
timestamp 1608254825
transform 1 0 29072 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2603_
timestamp 1608254825
transform 1 0 29440 0 -1 37536
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_64_335
timestamp 1608254825
transform 1 0 31924 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_327
timestamp 1608254825
transform 1 0 31188 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_561
timestamp 1608254825
transform 1 0 32016 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2546_
timestamp 1608254825
transform 1 0 32108 0 -1 37536
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_64_356
timestamp 1608254825
transform 1 0 33856 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2586_
timestamp 1608254825
transform 1 0 34224 0 -1 37536
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_64_379
timestamp 1608254825
transform 1 0 35972 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_410
timestamp 1608254825
transform 1 0 38824 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_64_398
timestamp 1608254825
transform 1 0 37720 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_391
timestamp 1608254825
transform 1 0 37076 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_562
timestamp 1608254825
transform 1 0 37628 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1608254825
transform -1 0 39836 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_65_15
timestamp 1608254825
transform 1 0 2484 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_3
timestamp 1608254825
transform 1 0 1380 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1608254825
transform 1 0 1104 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _2564_
timestamp 1608254825
transform 1 0 3588 0 1 37536
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_65_65
timestamp 1608254825
transform 1 0 7084 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_65_58
timestamp 1608254825
transform 1 0 6440 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_65_46
timestamp 1608254825
transform 1 0 5336 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_563
timestamp 1608254825
transform 1 0 6716 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _2401_
timestamp 1608254825
transform 1 0 6808 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_65_76
timestamp 1608254825
transform 1 0 8096 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2537_
timestamp 1608254825
transform 1 0 8464 0 1 37536
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_2  _2002_
timestamp 1608254825
transform 1 0 7820 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_65_110
timestamp 1608254825
transform 1 0 11224 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_99
timestamp 1608254825
transform 1 0 10212 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__and2_4  _1963_
timestamp 1608254825
transform 1 0 10580 0 1 37536
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_564
timestamp 1608254825
transform 1 0 12328 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2691_
timestamp 1608254825
transform 1 0 12420 0 1 37536
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_65_155
timestamp 1608254825
transform 1 0 15364 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_65_149
timestamp 1608254825
transform 1 0 14812 0 1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_65_142
timestamp 1608254825
transform 1 0 14168 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2559_
timestamp 1608254825
transform 1 0 15456 0 1 37536
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_2  _1321_
timestamp 1608254825
transform 1 0 14536 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_65_175
timestamp 1608254825
transform 1 0 17204 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_65_201
timestamp 1608254825
transform 1 0 19596 0 1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_565
timestamp 1608254825
transform 1 0 17940 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__o41a_4  _1303_
timestamp 1608254825
transform 1 0 18032 0 1 37536
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_6  FILLER_65_227
timestamp 1608254825
transform 1 0 21988 0 1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_207
timestamp 1608254825
transform 1 0 20148 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2695_
timestamp 1608254825
transform 1 0 20240 0 1 37536
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_65_240
timestamp 1608254825
transform 1 0 23184 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_566
timestamp 1608254825
transform 1 0 23552 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2700_
timestamp 1608254825
transform 1 0 23644 0 1 37536
box -38 -48 1786 592
use sky130_fd_sc_hd__and2_4  _1847_
timestamp 1608254825
transform 1 0 22540 0 1 37536
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_65_264
timestamp 1608254825
transform 1 0 25392 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _2613_
timestamp 1608254825
transform 1 0 26128 0 1 37536
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_65_291
timestamp 1608254825
transform 1 0 27876 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _2404_
timestamp 1608254825
transform 1 0 28244 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_65_306
timestamp 1608254825
transform 1 0 29256 0 1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_65_299
timestamp 1608254825
transform 1 0 28612 0 1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_6
timestamp 1608254825
transform 1 0 29808 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_567
timestamp 1608254825
transform 1 0 29164 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2563_
timestamp 1608254825
transform 1 0 29992 0 1 37536
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_65_337
timestamp 1608254825
transform 1 0 32108 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_333
timestamp 1608254825
transform 1 0 31740 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _2617_
timestamp 1608254825
transform 1 0 32200 0 1 37536
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_65_365
timestamp 1608254825
transform 1 0 34684 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_65_357
timestamp 1608254825
transform 1 0 33948 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_65_379
timestamp 1608254825
transform 1 0 35972 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_367
timestamp 1608254825
transform 1 0 34868 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_568
timestamp 1608254825
transform 1 0 34776 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_65_403
timestamp 1608254825
transform 1 0 38180 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_65_391
timestamp 1608254825
transform 1 0 37076 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_3
timestamp 1608254825
transform 1 0 38456 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _2403_
timestamp 1608254825
transform 1 0 38640 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_65_412
timestamp 1608254825
transform 1 0 39008 0 1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1608254825
transform -1 0 39836 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_66_15
timestamp 1608254825
transform 1 0 2484 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_3
timestamp 1608254825
transform 1 0 1380 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1608254825
transform 1 0 1104 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_66_44
timestamp 1608254825
transform 1 0 5152 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_32
timestamp 1608254825
transform 1 0 4048 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_66_27
timestamp 1608254825
transform 1 0 3588 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_569
timestamp 1608254825
transform 1 0 3956 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_63
timestamp 1608254825
transform 1 0 6900 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_56
timestamp 1608254825
transform 1 0 6256 0 -1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_570
timestamp 1608254825
transform 1 0 6808 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_66_84
timestamp 1608254825
transform 1 0 8832 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_4  _1996_
timestamp 1608254825
transform 1 0 8004 0 -1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_66_94
timestamp 1608254825
transform 1 0 9752 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_66_92
timestamp 1608254825
transform 1 0 9568 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_571
timestamp 1608254825
transform 1 0 9660 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2545_
timestamp 1608254825
transform 1 0 9936 0 -1 38624
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_66_130
timestamp 1608254825
transform 1 0 13064 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_66_125
timestamp 1608254825
transform 1 0 12604 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_66_123
timestamp 1608254825
transform 1 0 12420 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_66_115
timestamp 1608254825
transform 1 0 11684 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_572
timestamp 1608254825
transform 1 0 12512 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1331_
timestamp 1608254825
transform 1 0 12788 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_66_159
timestamp 1608254825
transform 1 0 15732 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_66_151
timestamp 1608254825
transform 1 0 14996 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_573
timestamp 1608254825
transform 1 0 15364 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1326_
timestamp 1608254825
transform 1 0 15456 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_4  _1325_
timestamp 1608254825
transform 1 0 14168 0 -1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_66_171
timestamp 1608254825
transform 1 0 16836 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_66_195
timestamp 1608254825
transform 1 0 19044 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_191
timestamp 1608254825
transform 1 0 18676 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_187
timestamp 1608254825
transform 1 0 18308 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_66_183
timestamp 1608254825
transform 1 0 17940 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_574
timestamp 1608254825
transform 1 0 18216 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1308_
timestamp 1608254825
transform 1 0 18768 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_4  _1307_
timestamp 1608254825
transform 1 0 19412 0 -1 38624
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_1  FILLER_66_222
timestamp 1608254825
transform 1 0 21528 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_218
timestamp 1608254825
transform 1 0 21160 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_213
timestamp 1608254825
transform 1 0 20700 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_575
timestamp 1608254825
transform 1 0 21068 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__nand3_4  _1283_
timestamp 1608254825
transform 1 0 21620 0 -1 38624
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_6  FILLER_66_249
timestamp 1608254825
transform 1 0 24012 0 -1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_66_245
timestamp 1608254825
transform 1 0 23644 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_66_237
timestamp 1608254825
transform 1 0 22908 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_576
timestamp 1608254825
transform 1 0 23920 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_66_255
timestamp 1608254825
transform 1 0 24564 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _2621_
timestamp 1608254825
transform 1 0 24656 0 -1 38624
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_66_287
timestamp 1608254825
transform 1 0 27508 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_275
timestamp 1608254825
transform 1 0 26404 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_577
timestamp 1608254825
transform 1 0 26772 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _1864_
timestamp 1608254825
transform 1 0 27876 0 -1 38624
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _1853_
timestamp 1608254825
transform 1 0 26864 0 -1 38624
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_66_318
timestamp 1608254825
transform 1 0 30360 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_66_298
timestamp 1608254825
transform 1 0 28520 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_578
timestamp 1608254825
transform 1 0 29624 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _1862_
timestamp 1608254825
transform 1 0 29716 0 -1 38624
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_66_342
timestamp 1608254825
transform 1 0 32568 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_329
timestamp 1608254825
transform 1 0 31372 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_579
timestamp 1608254825
transform 1 0 32476 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _1865_
timestamp 1608254825
transform 1 0 30728 0 -1 38624
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_66_354
timestamp 1608254825
transform 1 0 33672 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_385
timestamp 1608254825
transform 1 0 36524 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_373
timestamp 1608254825
transform 1 0 35420 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_366
timestamp 1608254825
transform 1 0 34776 0 -1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_580
timestamp 1608254825
transform 1 0 35328 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_404
timestamp 1608254825
transform 1 0 38272 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_397
timestamp 1608254825
transform 1 0 37628 0 -1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_581
timestamp 1608254825
transform 1 0 38180 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_66_416
timestamp 1608254825
transform 1 0 39376 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1608254825
transform -1 0 39836 0 -1 38624
box -38 -48 314 592
<< labels >>
rlabel metal2 s 12346 40200 12402 41000 6 CLK_LED
port 0 nsew signal tristate
rlabel metal2 s 29826 40200 29882 41000 6 DATA_AVAILABLE[0]
port 1 nsew signal input
rlabel metal2 s 25962 40200 26018 41000 6 DATA_AVAILABLE[1]
port 2 nsew signal input
rlabel metal3 s 0 29112 800 29232 6 DATA_AVAILABLE[2]
port 3 nsew signal input
rlabel metal3 s 40200 38632 41000 38752 6 DATA_AVAILABLE[3]
port 4 nsew signal input
rlabel metal2 s 17866 0 17922 800 6 DATA_AVAILABLE[4]
port 5 nsew signal input
rlabel metal2 s 21730 0 21786 800 6 DATA_AVAILABLE[5]
port 6 nsew signal input
rlabel metal2 s 37554 40200 37610 41000 6 DATA_FROM_HASH[0]
port 7 nsew signal input
rlabel metal2 s 14370 40200 14426 41000 6 DATA_FROM_HASH[1]
port 8 nsew signal input
rlabel metal3 s 0 34824 800 34944 6 DATA_FROM_HASH[2]
port 9 nsew signal input
rlabel metal3 s 40200 4360 41000 4480 6 DATA_FROM_HASH[3]
port 10 nsew signal input
rlabel metal2 s 23938 40200 23994 41000 6 DATA_FROM_HASH[4]
port 11 nsew signal input
rlabel metal2 s 23570 0 23626 800 6 DATA_FROM_HASH[5]
port 12 nsew signal input
rlabel metal2 s 2778 40200 2834 41000 6 DATA_FROM_HASH[6]
port 13 nsew signal input
rlabel metal3 s 40200 35912 41000 36032 6 DATA_FROM_HASH[7]
port 14 nsew signal input
rlabel metal2 s 4250 0 4306 800 6 DATA_TO_HASH[0]
port 15 nsew signal tristate
rlabel metal2 s 33322 0 33378 800 6 DATA_TO_HASH[1]
port 16 nsew signal tristate
rlabel metal2 s 16210 40200 16266 41000 6 DATA_TO_HASH[2]
port 17 nsew signal tristate
rlabel metal2 s 37186 0 37242 800 6 DATA_TO_HASH[3]
port 18 nsew signal tristate
rlabel metal3 s 40200 13064 41000 13184 6 DATA_TO_HASH[4]
port 19 nsew signal tristate
rlabel metal2 s 31298 0 31354 800 6 DATA_TO_HASH[5]
port 20 nsew signal tristate
rlabel metal2 s 31666 40200 31722 41000 6 DATA_TO_HASH[6]
port 21 nsew signal tristate
rlabel metal2 s 4618 40200 4674 41000 6 DATA_TO_HASH[7]
port 22 nsew signal tristate
rlabel metal2 s 29458 0 29514 800 6 EXT_RESET_N_fromHost
port 23 nsew signal input
rlabel metal2 s 39394 40200 39450 41000 6 EXT_RESET_N_toClient
port 24 nsew signal tristate
rlabel metal2 s 10138 0 10194 800 6 HASH_ADDR[0]
port 25 nsew signal tristate
rlabel metal2 s 35530 40200 35586 41000 6 HASH_ADDR[1]
port 26 nsew signal tristate
rlabel metal3 s 0 23400 800 23520 6 HASH_ADDR[2]
port 27 nsew signal tristate
rlabel metal3 s 0 26392 800 26512 6 HASH_ADDR[3]
port 28 nsew signal tristate
rlabel metal2 s 22098 40200 22154 41000 6 HASH_ADDR[4]
port 29 nsew signal tristate
rlabel metal3 s 0 32104 800 32224 6 HASH_ADDR[5]
port 30 nsew signal tristate
rlabel metal3 s 40200 7352 41000 7472 6 HASH_EN
port 31 nsew signal tristate
rlabel metal3 s 0 9256 800 9376 6 HASH_LED
port 32 nsew signal tristate
rlabel metal3 s 40200 15784 41000 15904 6 ID_fromClient
port 33 nsew signal input
rlabel metal3 s 0 20680 800 20800 6 ID_toHost
port 34 nsew signal tristate
rlabel metal2 s 8114 0 8170 800 6 IRQ_OUT_fromClient
port 35 nsew signal input
rlabel metal2 s 6274 0 6330 800 6 IRQ_OUT_toHost
port 36 nsew signal tristate
rlabel metal2 s 25594 0 25650 800 6 M1_CLK_IN
port 37 nsew signal input
rlabel metal2 s 19706 0 19762 800 6 M1_CLK_SELECT
port 38 nsew signal input
rlabel metal2 s 15842 0 15898 800 6 MACRO_RD_SELECT[0]
port 39 nsew signal tristate
rlabel metal2 s 11978 0 12034 800 6 MACRO_RD_SELECT[1]
port 40 nsew signal tristate
rlabel metal2 s 18234 40200 18290 41000 6 MACRO_RD_SELECT[2]
port 41 nsew signal tristate
rlabel metal2 s 2410 0 2466 800 6 MACRO_RD_SELECT[3]
port 42 nsew signal tristate
rlabel metal3 s 40200 32920 41000 33040 6 MACRO_RD_SELECT[4]
port 43 nsew signal tristate
rlabel metal3 s 40200 1640 41000 1760 6 MACRO_RD_SELECT[5]
port 44 nsew signal tristate
rlabel metal2 s 10506 40200 10562 41000 6 MACRO_WR_SELECT[0]
port 45 nsew signal tristate
rlabel metal2 s 33690 40200 33746 41000 6 MACRO_WR_SELECT[1]
port 46 nsew signal tristate
rlabel metal3 s 40200 30200 41000 30320 6 MACRO_WR_SELECT[2]
port 47 nsew signal tristate
rlabel metal3 s 40200 10072 41000 10192 6 MACRO_WR_SELECT[3]
port 48 nsew signal tristate
rlabel metal2 s 39026 0 39082 800 6 MACRO_WR_SELECT[4]
port 49 nsew signal tristate
rlabel metal3 s 0 37816 800 37936 6 MACRO_WR_SELECT[5]
port 50 nsew signal tristate
rlabel metal3 s 40200 27208 41000 27328 6 MISO_fromClient
port 51 nsew signal input
rlabel metal3 s 40200 24488 41000 24608 6 MISO_toHost
port 52 nsew signal tristate
rlabel metal2 s 8482 40200 8538 41000 6 MOSI_fromHost
port 53 nsew signal input
rlabel metal2 s 27802 40200 27858 41000 6 MOSI_toClient
port 54 nsew signal tristate
rlabel metal3 s 0 3544 800 3664 6 PLL_INPUT
port 55 nsew signal input
rlabel metal2 s 570 0 626 800 6 S1_CLK_IN
port 56 nsew signal input
rlabel metal3 s 0 11976 800 12096 6 S1_CLK_SELECT
port 57 nsew signal input
rlabel metal2 s 14002 0 14058 800 6 SCLK_fromHost
port 58 nsew signal input
rlabel metal3 s 0 17688 800 17808 6 SCLK_toClient
port 59 nsew signal tristate
rlabel metal3 s 0 14968 800 15088 6 SCSN_fromHost
port 60 nsew signal input
rlabel metal2 s 27434 0 27490 800 6 SCSN_toClient
port 61 nsew signal tristate
rlabel metal2 s 35162 0 35218 800 6 THREAD_COUNT[0]
port 62 nsew signal input
rlabel metal2 s 20074 40200 20130 41000 6 THREAD_COUNT[1]
port 63 nsew signal input
rlabel metal2 s 754 40200 810 41000 6 THREAD_COUNT[2]
port 64 nsew signal input
rlabel metal3 s 40200 18776 41000 18896 6 THREAD_COUNT[3]
port 65 nsew signal input
rlabel metal3 s 0 6264 800 6384 6 m1_clk_local
port 66 nsew signal tristate
rlabel metal2 s 6642 40200 6698 41000 6 one
port 67 nsew signal tristate
rlabel metal3 s 40200 21496 41000 21616 6 zero
port 68 nsew signal tristate
rlabel metal4 s 34928 2128 35248 38672 6 vccd1
port 69 nsew power bidirectional
rlabel metal4 s 4208 2128 4528 38672 6 vccd1
port 70 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 38672 6 vssd1
port 71 nsew ground bidirectional
rlabel metal4 s 35588 2176 35908 38624 6 vccd2
port 72 nsew power bidirectional
rlabel metal4 s 4868 2176 5188 38624 6 vccd2
port 73 nsew power bidirectional
rlabel metal4 s 20228 2176 20548 38624 6 vssd2
port 74 nsew ground bidirectional
rlabel metal4 s 36248 2176 36568 38624 6 vdda1
port 75 nsew power bidirectional
rlabel metal4 s 5528 2176 5848 38624 6 vdda1
port 76 nsew power bidirectional
rlabel metal4 s 20888 2176 21208 38624 6 vssa1
port 77 nsew ground bidirectional
rlabel metal4 s 36908 2176 37228 38624 6 vdda2
port 78 nsew power bidirectional
rlabel metal4 s 6188 2176 6508 38624 6 vdda2
port 79 nsew power bidirectional
rlabel metal4 s 21548 2176 21868 38624 6 vssa2
port 80 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 41000 41000
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1608271489
<< obsli1 >>
rect 1104 85 238832 197489
<< obsm1 >>
rect 566 8 238832 197520
<< metal2 >>
rect 10690 199200 10746 200000
rect 34794 199200 34850 200000
rect 58898 199200 58954 200000
rect 82818 199200 82874 200000
rect 106922 199200 106978 200000
rect 131026 199200 131082 200000
rect 155130 199200 155186 200000
rect 179234 199200 179290 200000
rect 203154 199200 203210 200000
rect 227258 199200 227314 200000
rect 570 0 626 800
rect 24490 0 24546 800
rect 48594 0 48650 800
rect 72698 0 72754 800
rect 96802 0 96858 800
rect 120722 0 120778 800
rect 144826 0 144882 800
rect 168930 0 168986 800
rect 193034 0 193090 800
rect 216954 0 217010 800
<< obsm2 >>
rect 18 199144 10634 199200
rect 10802 199144 34738 199200
rect 34906 199144 58842 199200
rect 59010 199144 82762 199200
rect 82930 199144 106866 199200
rect 107034 199144 130970 199200
rect 131138 199144 155074 199200
rect 155242 199144 179178 199200
rect 179346 199144 203098 199200
rect 203266 199144 227202 199200
rect 227370 199144 238444 199200
rect 18 856 238444 199144
rect 18 2 514 856
rect 682 2 24434 856
rect 24602 2 48538 856
rect 48706 2 72642 856
rect 72810 2 96746 856
rect 96914 2 120666 856
rect 120834 2 144770 856
rect 144938 2 168874 856
rect 169042 2 192978 856
rect 193146 2 216898 856
rect 217066 2 238444 856
<< metal3 >>
rect 239200 181160 240000 181280
rect 0 178440 800 178560
rect 239200 145528 240000 145648
rect 0 143080 800 143200
rect 239200 110168 240000 110288
rect 0 107448 800 107568
rect 239200 74536 240000 74656
rect 0 71816 800 71936
rect 239200 38904 240000 39024
rect 0 36184 800 36304
rect 239200 3272 240000 3392
<< obsm3 >>
rect 13 181360 239200 197505
rect 13 181080 239120 181360
rect 13 178640 239200 181080
rect 880 178360 239200 178640
rect 13 145728 239200 178360
rect 13 145448 239120 145728
rect 13 143280 239200 145448
rect 880 143000 239200 143280
rect 13 110368 239200 143000
rect 13 110088 239120 110368
rect 13 107648 239200 110088
rect 880 107368 239200 107648
rect 13 74736 239200 107368
rect 13 74456 239120 74736
rect 13 72016 239200 74456
rect 880 71736 239200 72016
rect 13 39104 239200 71736
rect 13 38824 239120 39104
rect 13 36384 239200 38824
rect 880 36104 239200 36384
rect 13 3472 239200 36104
rect 13 3192 239120 3472
rect 13 35 239200 3192
<< metal4 >>
rect 4208 2128 4528 197520
rect 19568 2128 19888 197520
rect 34928 2128 35248 197520
rect 50288 2128 50608 197520
rect 65648 2128 65968 197520
rect 81008 2128 81328 197520
rect 96368 2128 96688 197520
rect 111728 2128 112048 197520
rect 127088 2128 127408 197520
rect 142448 2128 142768 197520
rect 157808 2128 158128 197520
rect 173168 2128 173488 197520
rect 188528 2128 188848 197520
rect 203888 2128 204208 197520
rect 219248 2128 219568 197520
rect 234608 2128 234928 197520
<< obsm4 >>
rect 2819 2048 4128 197165
rect 4608 2048 19488 197165
rect 19968 2048 34848 197165
rect 35328 2048 50208 197165
rect 50688 2048 65568 197165
rect 66048 2048 80928 197165
rect 81408 2048 96288 197165
rect 96768 2048 111648 197165
rect 112128 2048 127008 197165
rect 127488 2048 142368 197165
rect 142848 2048 157728 197165
rect 158208 2048 173088 197165
rect 173568 2048 188448 197165
rect 188928 2048 203808 197165
rect 204288 2048 219168 197165
rect 219648 2048 234528 197165
rect 235008 2048 235645 197165
rect 2819 307 235645 2048
<< obsm5 >>
rect 61572 17180 189588 121540
<< labels >>
rlabel metal2 s 131026 199200 131082 200000 6 CLK
port 1 nsew signal input
rlabel metal2 s 144826 0 144882 800 6 DATA_AVAILABLE
port 2 nsew signal output
rlabel metal2 s 24490 0 24546 800 6 DATA_FROM_HASH[0]
port 3 nsew signal output
rlabel metal2 s 570 0 626 800 6 DATA_FROM_HASH[1]
port 4 nsew signal output
rlabel metal2 s 179234 199200 179290 200000 6 DATA_FROM_HASH[2]
port 5 nsew signal output
rlabel metal2 s 216954 0 217010 800 6 DATA_FROM_HASH[3]
port 6 nsew signal output
rlabel metal3 s 239200 38904 240000 39024 6 DATA_FROM_HASH[4]
port 7 nsew signal output
rlabel metal2 s 72698 0 72754 800 6 DATA_FROM_HASH[5]
port 8 nsew signal output
rlabel metal2 s 34794 199200 34850 200000 6 DATA_FROM_HASH[6]
port 9 nsew signal output
rlabel metal3 s 0 143080 800 143200 6 DATA_FROM_HASH[7]
port 10 nsew signal output
rlabel metal2 s 82818 199200 82874 200000 6 DATA_TO_HASH[0]
port 11 nsew signal input
rlabel metal3 s 0 71816 800 71936 6 DATA_TO_HASH[1]
port 12 nsew signal input
rlabel metal3 s 239200 74536 240000 74656 6 DATA_TO_HASH[2]
port 13 nsew signal input
rlabel metal3 s 239200 3272 240000 3392 6 DATA_TO_HASH[3]
port 14 nsew signal input
rlabel metal3 s 0 178440 800 178560 6 DATA_TO_HASH[4]
port 15 nsew signal input
rlabel metal2 s 48594 0 48650 800 6 DATA_TO_HASH[5]
port 16 nsew signal input
rlabel metal2 s 203154 199200 203210 200000 6 DATA_TO_HASH[6]
port 17 nsew signal input
rlabel metal2 s 58898 199200 58954 200000 6 DATA_TO_HASH[7]
port 18 nsew signal input
rlabel metal2 s 155130 199200 155186 200000 6 HASH_ADDR[0]
port 19 nsew signal input
rlabel metal2 s 10690 199200 10746 200000 6 HASH_ADDR[1]
port 20 nsew signal input
rlabel metal2 s 227258 199200 227314 200000 6 HASH_ADDR[2]
port 21 nsew signal input
rlabel metal2 s 193034 0 193090 800 6 HASH_ADDR[3]
port 22 nsew signal input
rlabel metal3 s 0 36184 800 36304 6 HASH_ADDR[4]
port 23 nsew signal input
rlabel metal3 s 239200 181160 240000 181280 6 HASH_ADDR[5]
port 24 nsew signal input
rlabel metal2 s 96802 0 96858 800 6 HASH_EN
port 25 nsew signal input
rlabel metal2 s 120722 0 120778 800 6 MACRO_RD_SELECT
port 26 nsew signal input
rlabel metal3 s 239200 110168 240000 110288 6 MACRO_WR_SELECT
port 27 nsew signal input
rlabel metal3 s 239200 145528 240000 145648 6 THREAD_COUNT[0]
port 28 nsew signal output
rlabel metal3 s 0 107448 800 107568 6 THREAD_COUNT[1]
port 29 nsew signal output
rlabel metal2 s 106922 199200 106978 200000 6 THREAD_COUNT[2]
port 30 nsew signal output
rlabel metal2 s 168930 0 168986 800 6 THREAD_COUNT[3]
port 31 nsew signal output
rlabel metal4 s 219248 2128 219568 197520 6 VPWR
port 32 nsew power bidirectional
rlabel metal4 s 188528 2128 188848 197520 6 VPWR
port 33 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 197520 6 VPWR
port 34 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 197520 6 VPWR
port 35 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 197520 6 VPWR
port 36 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 197520 6 VPWR
port 37 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 197520 6 VPWR
port 38 nsew power bidirectional
rlabel metal4 s 4208 2128 4528 197520 6 VPWR
port 39 nsew power bidirectional
rlabel metal4 s 234608 2128 234928 197520 6 VGND
port 40 nsew ground bidirectional
rlabel metal4 s 203888 2128 204208 197520 6 VGND
port 41 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 197520 6 VGND
port 42 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 197520 6 VGND
port 43 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 197520 6 VGND
port 44 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 197520 6 VGND
port 45 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 197520 6 VGND
port 46 nsew ground bidirectional
rlabel metal4 s 19568 2128 19888 197520 6 VGND
port 47 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 240000 200000
string LEFview TRUE
<< end >>
